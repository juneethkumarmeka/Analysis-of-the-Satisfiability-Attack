module basic_1500_15000_2000_5_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_450,In_412);
and U1 (N_1,In_214,In_380);
or U2 (N_2,In_1416,In_1454);
xor U3 (N_3,In_196,In_1066);
nand U4 (N_4,In_612,In_1043);
nand U5 (N_5,In_1242,In_276);
nand U6 (N_6,In_983,In_1208);
or U7 (N_7,In_1136,In_742);
nand U8 (N_8,In_705,In_40);
or U9 (N_9,In_530,In_1426);
nand U10 (N_10,In_476,In_625);
nor U11 (N_11,In_1305,In_1435);
nor U12 (N_12,In_367,In_1108);
nor U13 (N_13,In_349,In_200);
or U14 (N_14,In_782,In_956);
xor U15 (N_15,In_206,In_925);
or U16 (N_16,In_108,In_644);
or U17 (N_17,In_1004,In_109);
and U18 (N_18,In_697,In_18);
xnor U19 (N_19,In_41,In_991);
xor U20 (N_20,In_1332,In_1476);
xnor U21 (N_21,In_418,In_970);
or U22 (N_22,In_185,In_1339);
nor U23 (N_23,In_1433,In_1440);
nand U24 (N_24,In_1079,In_1163);
and U25 (N_25,In_313,In_753);
or U26 (N_26,In_1458,In_219);
or U27 (N_27,In_518,In_519);
and U28 (N_28,In_718,In_700);
nor U29 (N_29,In_482,In_298);
xor U30 (N_30,In_842,In_536);
nor U31 (N_31,In_657,In_791);
or U32 (N_32,In_1463,In_49);
nor U33 (N_33,In_894,In_14);
or U34 (N_34,In_436,In_480);
or U35 (N_35,In_977,In_233);
xor U36 (N_36,In_1159,In_1289);
xnor U37 (N_37,In_998,In_578);
nor U38 (N_38,In_356,In_391);
nand U39 (N_39,In_580,In_1457);
xnor U40 (N_40,In_247,In_346);
nor U41 (N_41,In_169,In_211);
nor U42 (N_42,In_1116,In_1177);
xnor U43 (N_43,In_432,In_966);
nor U44 (N_44,In_881,In_1414);
nand U45 (N_45,In_1491,In_1037);
and U46 (N_46,In_145,In_25);
and U47 (N_47,In_1232,In_735);
xnor U48 (N_48,In_1376,In_904);
nand U49 (N_49,In_309,In_1248);
nand U50 (N_50,In_1386,In_408);
and U51 (N_51,In_938,In_318);
xnor U52 (N_52,In_301,In_1);
nor U53 (N_53,In_484,In_1373);
nor U54 (N_54,In_57,In_290);
and U55 (N_55,In_1156,In_996);
xnor U56 (N_56,In_382,In_148);
or U57 (N_57,In_443,In_74);
and U58 (N_58,In_1175,In_926);
and U59 (N_59,In_328,In_1234);
or U60 (N_60,In_1383,In_260);
and U61 (N_61,In_902,In_610);
and U62 (N_62,In_725,In_1205);
nand U63 (N_63,In_1410,In_638);
nand U64 (N_64,In_22,In_1132);
xnor U65 (N_65,In_101,In_766);
or U66 (N_66,In_815,In_1387);
or U67 (N_67,In_682,In_497);
and U68 (N_68,In_1231,In_469);
or U69 (N_69,In_32,In_854);
xnor U70 (N_70,In_872,In_361);
nand U71 (N_71,In_331,In_559);
nand U72 (N_72,In_68,In_634);
nand U73 (N_73,In_188,In_1046);
nand U74 (N_74,In_957,In_66);
and U75 (N_75,In_603,In_447);
xor U76 (N_76,In_707,In_2);
nor U77 (N_77,In_1460,In_543);
xor U78 (N_78,In_969,In_359);
or U79 (N_79,In_1478,In_776);
or U80 (N_80,In_1169,In_319);
nand U81 (N_81,In_781,In_964);
nand U82 (N_82,In_245,In_943);
nor U83 (N_83,In_1298,In_726);
nand U84 (N_84,In_581,In_106);
and U85 (N_85,In_680,In_237);
xnor U86 (N_86,In_263,In_1093);
nor U87 (N_87,In_236,In_1192);
and U88 (N_88,In_1388,In_647);
nand U89 (N_89,In_1183,In_1041);
xnor U90 (N_90,In_1214,In_793);
nand U91 (N_91,In_118,In_900);
nand U92 (N_92,In_761,In_1436);
or U93 (N_93,In_927,In_997);
and U94 (N_94,In_1449,In_466);
nor U95 (N_95,In_656,In_1134);
and U96 (N_96,In_661,In_558);
xnor U97 (N_97,In_1350,In_48);
nor U98 (N_98,In_1385,In_394);
or U99 (N_99,In_1210,In_453);
nor U100 (N_100,In_336,In_75);
xor U101 (N_101,In_917,In_1431);
or U102 (N_102,In_215,In_1085);
nand U103 (N_103,In_660,In_590);
and U104 (N_104,In_732,In_712);
nand U105 (N_105,In_857,In_1001);
nand U106 (N_106,In_459,In_1178);
nor U107 (N_107,In_1455,In_1328);
nor U108 (N_108,In_327,In_1076);
nor U109 (N_109,In_841,In_929);
nand U110 (N_110,In_351,In_1061);
nand U111 (N_111,In_566,In_69);
nand U112 (N_112,In_151,In_1228);
xor U113 (N_113,In_181,In_796);
nor U114 (N_114,In_1258,In_15);
nand U115 (N_115,In_401,In_93);
nand U116 (N_116,In_993,In_863);
nor U117 (N_117,In_639,In_640);
xor U118 (N_118,In_1171,In_172);
xnor U119 (N_119,In_1086,In_468);
xnor U120 (N_120,In_1400,In_867);
nor U121 (N_121,In_1196,In_1408);
nand U122 (N_122,In_1212,In_873);
xnor U123 (N_123,In_887,In_375);
xor U124 (N_124,In_1427,In_921);
xor U125 (N_125,In_1225,In_345);
xor U126 (N_126,In_84,In_1027);
nor U127 (N_127,In_1009,In_344);
nand U128 (N_128,In_1052,In_176);
or U129 (N_129,In_315,In_1166);
nand U130 (N_130,In_1187,In_187);
nor U131 (N_131,In_64,In_579);
or U132 (N_132,In_42,In_940);
and U133 (N_133,In_1343,In_242);
nand U134 (N_134,In_175,In_1073);
and U135 (N_135,In_1493,In_1124);
nor U136 (N_136,In_458,In_1444);
nor U137 (N_137,In_811,In_475);
and U138 (N_138,In_968,In_686);
xor U139 (N_139,In_704,In_1346);
or U140 (N_140,In_504,In_365);
and U141 (N_141,In_1301,In_1285);
or U142 (N_142,In_1084,In_958);
and U143 (N_143,In_90,In_850);
or U144 (N_144,In_1068,In_522);
or U145 (N_145,In_950,In_1390);
nand U146 (N_146,In_292,In_1157);
and U147 (N_147,In_960,In_893);
and U148 (N_148,In_1302,In_147);
xor U149 (N_149,In_990,In_483);
nand U150 (N_150,In_995,In_801);
xor U151 (N_151,In_1000,In_160);
or U152 (N_152,In_944,In_1135);
or U153 (N_153,In_1259,In_238);
nor U154 (N_154,In_103,In_249);
and U155 (N_155,In_370,In_1303);
and U156 (N_156,In_1424,In_560);
nand U157 (N_157,In_892,In_1054);
nand U158 (N_158,In_1103,In_212);
xor U159 (N_159,In_561,In_875);
or U160 (N_160,In_1468,In_1217);
or U161 (N_161,In_1353,In_271);
xnor U162 (N_162,In_1481,In_554);
nand U163 (N_163,In_163,In_687);
or U164 (N_164,In_73,In_1310);
nor U165 (N_165,In_422,In_743);
and U166 (N_166,In_1280,In_144);
or U167 (N_167,In_1405,In_912);
xor U168 (N_168,In_1490,In_1415);
and U169 (N_169,In_728,In_1437);
and U170 (N_170,In_1391,In_643);
or U171 (N_171,In_1226,In_906);
nand U172 (N_172,In_501,In_976);
and U173 (N_173,In_1271,In_737);
nand U174 (N_174,In_794,In_1221);
xor U175 (N_175,In_859,In_722);
nor U176 (N_176,In_39,In_1282);
nand U177 (N_177,In_646,In_767);
nor U178 (N_178,In_821,In_1083);
or U179 (N_179,In_589,In_355);
xnor U180 (N_180,In_1198,In_903);
nand U181 (N_181,In_1201,In_1125);
nor U182 (N_182,In_777,In_12);
nor U183 (N_183,In_1397,In_651);
nand U184 (N_184,In_227,In_1030);
xor U185 (N_185,In_823,In_514);
or U186 (N_186,In_348,In_243);
nand U187 (N_187,In_43,In_1233);
nand U188 (N_188,In_556,In_257);
or U189 (N_189,In_1112,In_673);
xor U190 (N_190,In_1260,In_445);
and U191 (N_191,In_1399,In_462);
and U192 (N_192,In_204,In_878);
nand U193 (N_193,In_54,In_1380);
nand U194 (N_194,In_547,In_528);
or U195 (N_195,In_114,In_305);
xnor U196 (N_196,In_1266,In_282);
xnor U197 (N_197,In_748,In_1456);
nand U198 (N_198,In_296,In_652);
nand U199 (N_199,In_322,In_202);
and U200 (N_200,In_936,In_749);
and U201 (N_201,In_414,In_1174);
and U202 (N_202,In_895,In_1360);
nand U203 (N_203,In_1011,In_789);
and U204 (N_204,In_133,In_542);
xnor U205 (N_205,In_1074,In_496);
and U206 (N_206,In_1056,In_416);
nor U207 (N_207,In_324,In_283);
nor U208 (N_208,In_1355,In_222);
and U209 (N_209,In_21,In_1209);
nor U210 (N_210,In_107,In_1296);
nand U211 (N_211,In_511,In_802);
xor U212 (N_212,In_540,In_916);
nand U213 (N_213,In_1315,In_810);
and U214 (N_214,In_223,In_78);
or U215 (N_215,In_303,In_617);
nor U216 (N_216,In_24,In_509);
and U217 (N_217,In_1077,In_1247);
nor U218 (N_218,In_383,In_1498);
and U219 (N_219,In_410,In_1019);
or U220 (N_220,In_1281,In_930);
nor U221 (N_221,In_493,In_1092);
nor U222 (N_222,In_783,In_1459);
xor U223 (N_223,In_1176,In_464);
nor U224 (N_224,In_633,In_350);
and U225 (N_225,In_404,In_491);
and U226 (N_226,In_494,In_1106);
or U227 (N_227,In_369,In_439);
xnor U228 (N_228,In_937,In_645);
nor U229 (N_229,In_1269,In_1143);
xnor U230 (N_230,In_465,In_232);
nor U231 (N_231,In_1200,In_1039);
nor U232 (N_232,In_862,In_193);
and U233 (N_233,In_96,In_1487);
or U234 (N_234,In_562,In_548);
nand U235 (N_235,In_1138,In_374);
nand U236 (N_236,In_1291,In_1155);
and U237 (N_237,In_860,In_979);
or U238 (N_238,In_81,In_1434);
nand U239 (N_239,In_1401,In_190);
and U240 (N_240,In_675,In_325);
nor U241 (N_241,In_1477,In_846);
or U242 (N_242,In_1229,In_61);
and U243 (N_243,In_773,In_339);
nand U244 (N_244,In_433,In_387);
xnor U245 (N_245,In_827,In_88);
nand U246 (N_246,In_1420,In_1145);
or U247 (N_247,In_1133,In_935);
xor U248 (N_248,In_1186,In_1382);
xor U249 (N_249,In_914,In_1307);
or U250 (N_250,In_658,In_472);
and U251 (N_251,In_1294,In_601);
and U252 (N_252,In_122,In_648);
nand U253 (N_253,In_1115,In_573);
nor U254 (N_254,In_1341,In_905);
and U255 (N_255,In_775,In_1097);
nor U256 (N_256,In_1264,In_1423);
or U257 (N_257,In_1216,In_134);
nand U258 (N_258,In_490,In_963);
xnor U259 (N_259,In_877,In_272);
and U260 (N_260,In_759,In_941);
xor U261 (N_261,In_533,In_1015);
xnor U262 (N_262,In_1241,In_779);
nand U263 (N_263,In_994,In_498);
and U264 (N_264,In_220,In_138);
or U265 (N_265,In_89,In_97);
and U266 (N_266,In_1031,In_539);
nand U267 (N_267,In_1497,In_839);
nor U268 (N_268,In_911,In_812);
or U269 (N_269,In_70,In_140);
xnor U270 (N_270,In_816,In_250);
and U271 (N_271,In_758,In_1101);
or U272 (N_272,In_1309,In_128);
nand U273 (N_273,In_1150,In_1368);
xnor U274 (N_274,In_1203,In_1014);
and U275 (N_275,In_654,In_524);
xnor U276 (N_276,In_1121,In_901);
xor U277 (N_277,In_285,In_1235);
xnor U278 (N_278,In_701,In_461);
or U279 (N_279,In_931,In_1238);
and U280 (N_280,In_1049,In_745);
xor U281 (N_281,In_1158,In_596);
nand U282 (N_282,In_664,In_959);
or U283 (N_283,In_951,In_1377);
or U284 (N_284,In_570,In_1075);
xor U285 (N_285,In_53,In_1044);
nor U286 (N_286,In_865,In_1185);
and U287 (N_287,In_198,In_507);
and U288 (N_288,In_1189,In_891);
nor U289 (N_289,In_1236,In_479);
and U290 (N_290,In_731,In_1010);
or U291 (N_291,In_487,In_999);
and U292 (N_292,In_588,In_764);
nand U293 (N_293,In_1202,In_83);
or U294 (N_294,In_534,In_520);
and U295 (N_295,In_180,In_1372);
or U296 (N_296,In_1114,In_1336);
or U297 (N_297,In_314,In_844);
xnor U298 (N_298,In_517,In_440);
nor U299 (N_299,In_535,In_289);
nor U300 (N_300,In_388,In_378);
nand U301 (N_301,In_830,In_618);
and U302 (N_302,In_919,In_1317);
or U303 (N_303,In_1167,In_1421);
or U304 (N_304,In_1467,In_1105);
or U305 (N_305,In_636,In_826);
xor U306 (N_306,In_692,In_1363);
and U307 (N_307,In_1117,In_218);
and U308 (N_308,In_1293,In_1495);
nand U309 (N_309,In_1219,In_270);
or U310 (N_310,In_164,In_577);
or U311 (N_311,In_785,In_1499);
xor U312 (N_312,In_1334,In_33);
nand U313 (N_313,In_11,In_591);
and U314 (N_314,In_1439,In_455);
nor U315 (N_315,In_795,In_1365);
and U316 (N_316,In_1256,In_946);
or U317 (N_317,In_699,In_199);
xor U318 (N_318,In_111,In_1329);
nand U319 (N_319,In_438,In_442);
or U320 (N_320,In_441,In_168);
nor U321 (N_321,In_1398,In_368);
or U322 (N_322,In_105,In_1139);
nor U323 (N_323,In_1218,In_321);
nor U324 (N_324,In_1412,In_1072);
nor U325 (N_325,In_1411,In_31);
nor U326 (N_326,In_741,In_619);
nor U327 (N_327,In_628,In_209);
or U328 (N_328,In_347,In_400);
or U329 (N_329,In_843,In_311);
nor U330 (N_330,In_550,In_332);
nor U331 (N_331,In_1040,In_828);
nand U332 (N_332,In_1288,In_1038);
xor U333 (N_333,In_832,In_1206);
and U334 (N_334,In_304,In_130);
xor U335 (N_335,In_91,In_788);
nand U336 (N_336,In_76,In_463);
nor U337 (N_337,In_1022,In_281);
nand U338 (N_338,In_756,In_1181);
nor U339 (N_339,In_1240,In_677);
xor U340 (N_340,In_165,In_470);
xor U341 (N_341,In_112,In_869);
and U342 (N_342,In_1126,In_273);
nand U343 (N_343,In_1274,In_653);
or U344 (N_344,In_1070,In_0);
and U345 (N_345,In_593,In_17);
or U346 (N_346,In_703,In_973);
and U347 (N_347,In_564,In_829);
nor U348 (N_348,In_1149,In_545);
or U349 (N_349,In_655,In_121);
xor U350 (N_350,In_306,In_505);
and U351 (N_351,In_800,In_254);
xor U352 (N_352,In_1062,In_1348);
or U353 (N_353,In_1028,In_79);
nand U354 (N_354,In_553,In_626);
nand U355 (N_355,In_797,In_240);
nand U356 (N_356,In_510,In_477);
xnor U357 (N_357,In_586,In_294);
and U358 (N_358,In_609,In_861);
and U359 (N_359,In_1462,In_373);
nand U360 (N_360,In_399,In_495);
xnor U361 (N_361,In_1252,In_1419);
nand U362 (N_362,In_771,In_104);
xnor U363 (N_363,In_635,In_616);
nand U364 (N_364,In_1013,In_36);
nand U365 (N_365,In_1170,In_1162);
xor U366 (N_366,In_814,In_1131);
nand U367 (N_367,In_228,In_606);
or U368 (N_368,In_155,In_690);
or U369 (N_369,In_1479,In_1223);
nand U370 (N_370,In_1127,In_1335);
nand U371 (N_371,In_451,In_672);
nor U372 (N_372,In_1017,In_1403);
xnor U373 (N_373,In_1033,In_203);
nand U374 (N_374,In_293,In_642);
xnor U375 (N_375,In_984,In_1306);
nor U376 (N_376,In_264,In_736);
or U377 (N_377,In_1316,In_774);
nand U378 (N_378,In_809,In_1057);
nor U379 (N_379,In_473,In_1267);
and U380 (N_380,In_47,In_1120);
nand U381 (N_381,In_421,In_965);
nand U382 (N_382,In_1250,In_702);
nor U383 (N_383,In_286,In_1195);
nand U384 (N_384,In_723,In_1286);
nand U385 (N_385,In_267,In_1110);
xnor U386 (N_386,In_913,In_1445);
and U387 (N_387,In_1448,In_1331);
xnor U388 (N_388,In_825,In_51);
nand U389 (N_389,In_1026,In_149);
and U390 (N_390,In_1297,In_1006);
xnor U391 (N_391,In_1482,In_110);
nor U392 (N_392,In_768,In_786);
nor U393 (N_393,In_713,In_1313);
xnor U394 (N_394,In_398,In_523);
nand U395 (N_395,In_1058,In_157);
nor U396 (N_396,In_607,In_711);
nor U397 (N_397,In_424,In_123);
and U398 (N_398,In_158,In_343);
nand U399 (N_399,In_225,In_1230);
nand U400 (N_400,In_1165,In_605);
nor U401 (N_401,In_7,In_978);
nor U402 (N_402,In_627,In_1404);
and U403 (N_403,In_1194,In_288);
or U404 (N_404,In_1064,In_953);
nand U405 (N_405,In_909,In_1249);
nor U406 (N_406,In_615,In_258);
nor U407 (N_407,In_1193,In_1244);
nor U408 (N_408,In_256,In_437);
and U409 (N_409,In_1094,In_478);
or U410 (N_410,In_55,In_407);
nor U411 (N_411,In_734,In_1344);
nand U412 (N_412,In_1224,In_1107);
xor U413 (N_413,In_1299,In_1474);
or U414 (N_414,In_952,In_329);
or U415 (N_415,In_1204,In_419);
or U416 (N_416,In_874,In_72);
or U417 (N_417,In_972,In_1428);
xor U418 (N_418,In_770,In_1413);
and U419 (N_419,In_52,In_113);
xor U420 (N_420,In_1374,In_1489);
nand U421 (N_421,In_727,In_954);
nand U422 (N_422,In_799,In_141);
nand U423 (N_423,In_674,In_598);
nand U424 (N_424,In_326,In_908);
nand U425 (N_425,In_1333,In_576);
xnor U426 (N_426,In_161,In_765);
and U427 (N_427,In_1263,In_1442);
nand U428 (N_428,In_221,In_23);
nor U429 (N_429,In_1323,In_526);
nand U430 (N_430,In_226,In_1304);
nor U431 (N_431,In_710,In_557);
and U432 (N_432,In_77,In_30);
nor U433 (N_433,In_502,In_847);
nor U434 (N_434,In_132,In_915);
nand U435 (N_435,In_817,In_1067);
nor U436 (N_436,In_4,In_721);
nor U437 (N_437,In_1087,In_486);
and U438 (N_438,In_156,In_415);
xnor U439 (N_439,In_1364,In_420);
xnor U440 (N_440,In_531,In_435);
and U441 (N_441,In_621,In_1464);
or U442 (N_442,In_274,In_244);
xnor U443 (N_443,In_1102,In_1409);
or U444 (N_444,In_569,In_183);
nor U445 (N_445,In_1262,In_864);
nor U446 (N_446,In_201,In_131);
nand U447 (N_447,In_760,In_1160);
or U448 (N_448,In_898,In_116);
and U449 (N_449,In_928,In_1213);
nor U450 (N_450,In_1091,In_948);
or U451 (N_451,In_932,In_44);
xor U452 (N_452,In_335,In_1308);
xnor U453 (N_453,In_173,In_813);
xor U454 (N_454,In_572,In_955);
and U455 (N_455,In_159,In_397);
nand U456 (N_456,In_688,In_1290);
xor U457 (N_457,In_259,In_592);
nor U458 (N_458,In_1432,In_879);
and U459 (N_459,In_992,In_1227);
xor U460 (N_460,In_546,In_503);
or U461 (N_461,In_769,In_352);
and U462 (N_462,In_922,In_1441);
nor U463 (N_463,In_334,In_95);
and U464 (N_464,In_681,In_1425);
xor U465 (N_465,In_402,In_279);
xnor U466 (N_466,In_1361,In_449);
and U467 (N_467,In_624,In_529);
xor U468 (N_468,In_757,In_308);
nor U469 (N_469,In_357,In_1351);
xor U470 (N_470,In_751,In_207);
or U471 (N_471,In_1366,In_755);
xnor U472 (N_472,In_689,In_428);
xnor U473 (N_473,In_255,In_818);
nor U474 (N_474,In_239,In_1023);
nor U475 (N_475,In_384,In_582);
or U476 (N_476,In_630,In_1008);
nand U477 (N_477,In_323,In_571);
nor U478 (N_478,In_693,In_235);
or U479 (N_479,In_287,In_379);
xor U480 (N_480,In_974,In_241);
and U481 (N_481,In_822,In_971);
nand U482 (N_482,In_537,In_166);
nand U483 (N_483,In_853,In_772);
nand U484 (N_484,In_1345,In_268);
or U485 (N_485,In_280,In_583);
nor U486 (N_486,In_708,In_85);
xnor U487 (N_487,In_231,In_360);
nand U488 (N_488,In_1471,In_277);
nor U489 (N_489,In_1443,In_87);
nand U490 (N_490,In_65,In_1246);
nand U491 (N_491,In_1480,In_595);
and U492 (N_492,In_716,In_143);
and U493 (N_493,In_525,In_587);
or U494 (N_494,In_427,In_933);
nand U495 (N_495,In_1325,In_1020);
and U496 (N_496,In_641,In_385);
xnor U497 (N_497,In_1319,In_1142);
or U498 (N_498,In_137,In_907);
and U499 (N_499,In_457,In_9);
xor U500 (N_500,In_154,In_1123);
and U501 (N_501,In_62,In_1347);
and U502 (N_502,In_1453,In_848);
xor U503 (N_503,In_1050,In_195);
and U504 (N_504,In_1469,In_358);
and U505 (N_505,In_1254,In_856);
xor U506 (N_506,In_338,In_837);
nand U507 (N_507,In_890,In_1024);
nand U508 (N_508,In_488,In_1287);
and U509 (N_509,In_448,In_481);
or U510 (N_510,In_1154,In_386);
nor U511 (N_511,In_806,In_1140);
and U512 (N_512,In_1211,In_186);
and U513 (N_513,In_208,In_1168);
nor U514 (N_514,In_1379,In_597);
and U515 (N_515,In_1389,In_1096);
or U516 (N_516,In_429,In_1395);
nor U517 (N_517,In_659,In_310);
nand U518 (N_518,In_1438,In_1342);
nand U519 (N_519,In_563,In_1327);
xnor U520 (N_520,In_1320,In_1257);
xnor U521 (N_521,In_189,In_1340);
nand U522 (N_522,In_541,In_1311);
or U523 (N_523,In_120,In_840);
nand U524 (N_524,In_19,In_452);
nor U525 (N_525,In_1255,In_986);
and U526 (N_526,In_182,In_1370);
nor U527 (N_527,In_527,In_67);
or U528 (N_528,In_1007,In_1393);
nand U529 (N_529,In_127,In_35);
nand U530 (N_530,In_1349,In_317);
nand U531 (N_531,In_1378,In_1191);
nor U532 (N_532,In_1318,In_1078);
and U533 (N_533,In_396,In_831);
or U534 (N_534,In_614,In_499);
and U535 (N_535,In_1089,In_670);
nor U536 (N_536,In_629,In_1082);
nor U537 (N_537,In_1407,In_1251);
nand U538 (N_538,In_299,In_623);
xor U539 (N_539,In_178,In_126);
nand U540 (N_540,In_1059,In_506);
and U541 (N_541,In_835,In_1002);
or U542 (N_542,In_600,In_975);
or U543 (N_543,In_1314,In_37);
xor U544 (N_544,In_80,In_763);
nor U545 (N_545,In_706,In_1180);
nor U546 (N_546,In_1279,In_192);
nor U547 (N_547,In_730,In_1016);
or U548 (N_548,In_1275,In_8);
nor U549 (N_549,In_552,In_229);
nor U550 (N_550,In_434,In_1021);
xor U551 (N_551,In_38,In_1222);
and U552 (N_552,In_1080,In_1100);
xor U553 (N_553,In_284,In_1312);
or U554 (N_554,In_150,In_16);
and U555 (N_555,In_1485,In_142);
nor U556 (N_556,In_1104,In_939);
xor U557 (N_557,In_26,In_885);
xnor U558 (N_558,In_82,In_733);
or U559 (N_559,In_585,In_1113);
and U560 (N_560,In_1450,In_883);
xnor U561 (N_561,In_1283,In_790);
or U562 (N_562,In_500,In_1277);
or U563 (N_563,In_836,In_278);
nor U564 (N_564,In_1470,In_1130);
nand U565 (N_565,In_60,In_1473);
xnor U566 (N_566,In_1122,In_316);
and U567 (N_567,In_744,In_162);
or U568 (N_568,In_1472,In_403);
nor U569 (N_569,In_1099,In_63);
and U570 (N_570,In_714,In_337);
or U571 (N_571,In_234,In_1243);
xor U572 (N_572,In_1447,In_1375);
nor U573 (N_573,In_197,In_389);
nor U574 (N_574,In_1109,In_631);
or U575 (N_575,In_620,In_1352);
xnor U576 (N_576,In_1475,In_513);
xnor U577 (N_577,In_1063,In_870);
nor U578 (N_578,In_45,In_982);
nand U579 (N_579,In_333,In_599);
or U580 (N_580,In_662,In_516);
and U581 (N_581,In_1053,In_393);
nand U582 (N_582,In_666,In_320);
nand U583 (N_583,In_217,In_1496);
nor U584 (N_584,In_1090,In_5);
and U585 (N_585,In_213,In_819);
and U586 (N_586,In_1446,In_947);
and U587 (N_587,In_532,In_1005);
xor U588 (N_588,In_1179,In_34);
or U589 (N_589,In_803,In_678);
xor U590 (N_590,In_780,In_981);
xnor U591 (N_591,In_1237,In_899);
nor U592 (N_592,In_544,In_94);
nor U593 (N_593,In_1245,In_1465);
xnor U594 (N_594,In_102,In_594);
and U595 (N_595,In_1147,In_1354);
xor U596 (N_596,In_833,In_882);
xnor U597 (N_597,In_1190,In_353);
xnor U598 (N_598,In_471,In_1119);
nand U599 (N_599,In_184,In_460);
nor U600 (N_600,In_1369,In_1484);
and U601 (N_601,In_967,In_1396);
nor U602 (N_602,In_6,In_1418);
nor U603 (N_603,In_58,In_1273);
or U604 (N_604,In_454,In_515);
xor U605 (N_605,In_312,In_417);
and U606 (N_606,In_411,In_1359);
or U607 (N_607,In_622,In_858);
xnor U608 (N_608,In_679,In_456);
xnor U609 (N_609,In_119,In_538);
or U610 (N_610,In_1161,In_1172);
and U611 (N_611,In_521,In_740);
nand U612 (N_612,In_1095,In_13);
or U613 (N_613,In_739,In_253);
xnor U614 (N_614,In_307,In_1042);
nor U615 (N_615,In_549,In_988);
and U616 (N_616,In_98,In_778);
nor U617 (N_617,In_362,In_663);
xor U618 (N_618,In_71,In_179);
nand U619 (N_619,In_1461,In_1276);
nor U620 (N_620,In_1422,In_124);
nand U621 (N_621,In_784,In_300);
or U622 (N_622,In_676,In_430);
or U623 (N_623,In_275,In_1430);
nand U624 (N_624,In_1207,In_1451);
nor U625 (N_625,In_866,In_613);
nor U626 (N_626,In_1486,In_1268);
and U627 (N_627,In_604,In_792);
nor U628 (N_628,In_1321,In_934);
and U629 (N_629,In_117,In_1394);
xnor U630 (N_630,In_1417,In_426);
or U631 (N_631,In_918,In_746);
and U632 (N_632,In_1129,In_1337);
xnor U633 (N_633,In_889,In_1048);
xnor U634 (N_634,In_1111,In_100);
nand U635 (N_635,In_1384,In_1272);
xor U636 (N_636,In_1088,In_1069);
nand U637 (N_637,In_942,In_1356);
nor U638 (N_638,In_980,In_949);
and U639 (N_639,In_787,In_565);
and U640 (N_640,In_210,In_99);
or U641 (N_641,In_423,In_174);
or U642 (N_642,In_551,In_667);
or U643 (N_643,In_880,In_171);
nor U644 (N_644,In_291,In_1045);
or U645 (N_645,In_724,In_251);
nor U646 (N_646,In_489,In_876);
nor U647 (N_647,In_897,In_302);
or U648 (N_648,In_1051,In_265);
xor U649 (N_649,In_671,In_1338);
nor U650 (N_650,In_1035,In_135);
and U651 (N_651,In_1494,In_56);
nand U652 (N_652,In_747,In_668);
nor U653 (N_653,In_86,In_413);
and U654 (N_654,In_719,In_834);
or U655 (N_655,In_1118,In_555);
xnor U656 (N_656,In_390,In_341);
nand U657 (N_657,In_405,In_10);
nor U658 (N_658,In_1153,In_266);
xor U659 (N_659,In_444,In_896);
or U660 (N_660,In_1358,In_1300);
nand U661 (N_661,In_1184,In_1292);
or U662 (N_662,In_431,In_252);
xnor U663 (N_663,In_824,In_611);
or U664 (N_664,In_297,In_152);
nand U665 (N_665,In_92,In_752);
or U666 (N_666,In_584,In_665);
and U667 (N_667,In_492,In_669);
xor U668 (N_668,In_129,In_849);
nand U669 (N_669,In_170,In_381);
or U670 (N_670,In_224,In_1330);
nor U671 (N_671,In_146,In_1197);
nor U672 (N_672,In_798,In_1151);
and U673 (N_673,In_602,In_46);
or U674 (N_674,In_695,In_50);
nor U675 (N_675,In_406,In_910);
xnor U676 (N_676,In_709,In_1367);
and U677 (N_677,In_246,In_1483);
xnor U678 (N_678,In_720,In_29);
nor U679 (N_679,In_1322,In_261);
nand U680 (N_680,In_696,In_567);
nand U681 (N_681,In_1492,In_376);
xnor U682 (N_682,In_139,In_342);
xnor U683 (N_683,In_1173,In_194);
nor U684 (N_684,In_750,In_762);
or U685 (N_685,In_136,In_685);
nor U686 (N_686,In_715,In_923);
xor U687 (N_687,In_1261,In_1371);
or U688 (N_688,In_987,In_637);
nor U689 (N_689,In_1253,In_177);
nor U690 (N_690,In_1098,In_1220);
or U691 (N_691,In_684,In_485);
xnor U692 (N_692,In_1141,In_989);
xor U693 (N_693,In_1452,In_409);
or U694 (N_694,In_1071,In_924);
or U695 (N_695,In_1146,In_1278);
and U696 (N_696,In_1003,In_807);
xor U697 (N_697,In_377,In_804);
xnor U698 (N_698,In_1148,In_1188);
nor U699 (N_699,In_364,In_698);
and U700 (N_700,In_205,In_372);
nor U701 (N_701,In_855,In_1164);
xnor U702 (N_702,In_1270,In_683);
or U703 (N_703,In_961,In_295);
and U704 (N_704,In_1144,In_945);
or U705 (N_705,In_27,In_467);
nand U706 (N_706,In_1295,In_392);
or U707 (N_707,In_608,In_1284);
nand U708 (N_708,In_216,In_738);
and U709 (N_709,In_1215,In_1047);
nand U710 (N_710,In_1199,In_754);
or U711 (N_711,In_395,In_632);
nor U712 (N_712,In_1012,In_3);
nand U713 (N_713,In_1488,In_153);
nor U714 (N_714,In_354,In_1357);
nor U715 (N_715,In_1055,In_28);
nand U716 (N_716,In_852,In_446);
and U717 (N_717,In_888,In_1402);
or U718 (N_718,In_1025,In_1060);
or U719 (N_719,In_1381,In_167);
or U720 (N_720,In_1182,In_886);
nor U721 (N_721,In_568,In_871);
nand U722 (N_722,In_191,In_269);
xor U723 (N_723,In_1081,In_1065);
or U724 (N_724,In_1429,In_474);
or U725 (N_725,In_1324,In_851);
xor U726 (N_726,In_1036,In_363);
or U727 (N_727,In_1326,In_1239);
nand U728 (N_728,In_884,In_115);
xnor U729 (N_729,In_1137,In_366);
xnor U730 (N_730,In_694,In_1034);
xor U731 (N_731,In_508,In_248);
or U732 (N_732,In_1128,In_729);
nand U733 (N_733,In_262,In_691);
nand U734 (N_734,In_845,In_717);
nand U735 (N_735,In_985,In_575);
or U736 (N_736,In_650,In_808);
nand U737 (N_737,In_1362,In_230);
and U738 (N_738,In_1029,In_920);
xor U739 (N_739,In_125,In_962);
or U740 (N_740,In_512,In_1406);
xor U741 (N_741,In_1466,In_330);
or U742 (N_742,In_425,In_805);
and U743 (N_743,In_340,In_1032);
nand U744 (N_744,In_20,In_820);
nand U745 (N_745,In_838,In_649);
nand U746 (N_746,In_1265,In_868);
nand U747 (N_747,In_59,In_1392);
or U748 (N_748,In_1018,In_371);
nand U749 (N_749,In_1152,In_574);
xnor U750 (N_750,In_1323,In_763);
and U751 (N_751,In_89,In_1334);
nor U752 (N_752,In_1451,In_233);
or U753 (N_753,In_305,In_888);
nor U754 (N_754,In_753,In_1078);
and U755 (N_755,In_638,In_260);
nand U756 (N_756,In_1465,In_427);
nand U757 (N_757,In_927,In_217);
xor U758 (N_758,In_771,In_949);
or U759 (N_759,In_1401,In_1013);
nand U760 (N_760,In_790,In_695);
or U761 (N_761,In_372,In_698);
xor U762 (N_762,In_742,In_1419);
nand U763 (N_763,In_565,In_511);
or U764 (N_764,In_715,In_742);
nand U765 (N_765,In_361,In_737);
nor U766 (N_766,In_1229,In_365);
or U767 (N_767,In_1277,In_753);
nor U768 (N_768,In_1185,In_495);
nand U769 (N_769,In_435,In_1004);
and U770 (N_770,In_531,In_1087);
nand U771 (N_771,In_1124,In_1432);
xnor U772 (N_772,In_38,In_610);
nor U773 (N_773,In_57,In_1194);
nand U774 (N_774,In_41,In_632);
and U775 (N_775,In_1258,In_686);
and U776 (N_776,In_1223,In_1454);
and U777 (N_777,In_1299,In_1296);
nor U778 (N_778,In_804,In_564);
nor U779 (N_779,In_223,In_1008);
and U780 (N_780,In_1431,In_151);
nor U781 (N_781,In_633,In_212);
nor U782 (N_782,In_15,In_845);
nor U783 (N_783,In_1191,In_172);
nor U784 (N_784,In_870,In_1140);
or U785 (N_785,In_1273,In_261);
xor U786 (N_786,In_335,In_485);
nor U787 (N_787,In_222,In_14);
nand U788 (N_788,In_1443,In_595);
or U789 (N_789,In_1216,In_671);
or U790 (N_790,In_150,In_1482);
and U791 (N_791,In_1199,In_307);
nand U792 (N_792,In_330,In_1365);
or U793 (N_793,In_1448,In_1234);
or U794 (N_794,In_479,In_507);
and U795 (N_795,In_163,In_1054);
nand U796 (N_796,In_173,In_241);
and U797 (N_797,In_1118,In_837);
nand U798 (N_798,In_961,In_262);
and U799 (N_799,In_81,In_321);
or U800 (N_800,In_1078,In_1487);
nor U801 (N_801,In_928,In_1376);
or U802 (N_802,In_1267,In_415);
nor U803 (N_803,In_1265,In_154);
or U804 (N_804,In_1237,In_1030);
nor U805 (N_805,In_261,In_1359);
and U806 (N_806,In_978,In_956);
or U807 (N_807,In_320,In_921);
xor U808 (N_808,In_502,In_910);
and U809 (N_809,In_248,In_1395);
and U810 (N_810,In_1130,In_453);
xor U811 (N_811,In_576,In_519);
xnor U812 (N_812,In_1115,In_1285);
and U813 (N_813,In_183,In_193);
nor U814 (N_814,In_1115,In_502);
nor U815 (N_815,In_908,In_1365);
nor U816 (N_816,In_373,In_206);
and U817 (N_817,In_788,In_575);
and U818 (N_818,In_525,In_1325);
and U819 (N_819,In_223,In_1070);
nor U820 (N_820,In_630,In_988);
and U821 (N_821,In_268,In_943);
nand U822 (N_822,In_103,In_699);
nor U823 (N_823,In_397,In_963);
or U824 (N_824,In_1048,In_109);
and U825 (N_825,In_756,In_914);
nor U826 (N_826,In_718,In_1044);
nor U827 (N_827,In_1121,In_1226);
or U828 (N_828,In_1000,In_574);
and U829 (N_829,In_950,In_1027);
or U830 (N_830,In_1437,In_402);
and U831 (N_831,In_1321,In_467);
xnor U832 (N_832,In_1306,In_1399);
xnor U833 (N_833,In_107,In_591);
xor U834 (N_834,In_850,In_655);
nor U835 (N_835,In_506,In_1477);
nor U836 (N_836,In_174,In_1022);
nand U837 (N_837,In_723,In_356);
and U838 (N_838,In_604,In_631);
and U839 (N_839,In_479,In_960);
and U840 (N_840,In_1193,In_316);
nand U841 (N_841,In_625,In_1488);
nand U842 (N_842,In_182,In_1221);
nand U843 (N_843,In_926,In_1350);
or U844 (N_844,In_1212,In_1136);
nor U845 (N_845,In_923,In_438);
nor U846 (N_846,In_105,In_451);
nor U847 (N_847,In_500,In_862);
nand U848 (N_848,In_1409,In_1202);
or U849 (N_849,In_487,In_365);
or U850 (N_850,In_604,In_832);
xnor U851 (N_851,In_255,In_714);
and U852 (N_852,In_796,In_915);
and U853 (N_853,In_22,In_288);
and U854 (N_854,In_134,In_166);
or U855 (N_855,In_825,In_107);
xnor U856 (N_856,In_1149,In_52);
nor U857 (N_857,In_471,In_37);
nand U858 (N_858,In_555,In_115);
and U859 (N_859,In_1256,In_602);
and U860 (N_860,In_680,In_478);
nand U861 (N_861,In_513,In_1291);
nand U862 (N_862,In_135,In_271);
nor U863 (N_863,In_587,In_125);
xnor U864 (N_864,In_1246,In_742);
or U865 (N_865,In_1244,In_601);
or U866 (N_866,In_495,In_326);
nand U867 (N_867,In_854,In_199);
xor U868 (N_868,In_85,In_778);
xor U869 (N_869,In_1180,In_1235);
xor U870 (N_870,In_1332,In_216);
and U871 (N_871,In_940,In_1123);
nand U872 (N_872,In_1457,In_60);
xnor U873 (N_873,In_452,In_422);
xnor U874 (N_874,In_464,In_144);
nand U875 (N_875,In_1335,In_1086);
or U876 (N_876,In_1395,In_1451);
and U877 (N_877,In_326,In_981);
or U878 (N_878,In_1188,In_1027);
or U879 (N_879,In_712,In_46);
xnor U880 (N_880,In_1344,In_1299);
and U881 (N_881,In_1436,In_769);
and U882 (N_882,In_1177,In_714);
nor U883 (N_883,In_405,In_717);
nor U884 (N_884,In_1009,In_627);
or U885 (N_885,In_1272,In_491);
or U886 (N_886,In_45,In_1390);
xor U887 (N_887,In_1232,In_125);
or U888 (N_888,In_1164,In_1445);
nor U889 (N_889,In_1183,In_1486);
or U890 (N_890,In_186,In_874);
nand U891 (N_891,In_927,In_1158);
xnor U892 (N_892,In_474,In_464);
and U893 (N_893,In_773,In_1381);
xor U894 (N_894,In_1466,In_47);
or U895 (N_895,In_116,In_98);
or U896 (N_896,In_1454,In_401);
nand U897 (N_897,In_48,In_773);
xor U898 (N_898,In_1269,In_183);
nand U899 (N_899,In_496,In_425);
and U900 (N_900,In_135,In_548);
or U901 (N_901,In_284,In_439);
nand U902 (N_902,In_77,In_553);
nand U903 (N_903,In_617,In_409);
xnor U904 (N_904,In_305,In_493);
or U905 (N_905,In_622,In_745);
and U906 (N_906,In_730,In_998);
and U907 (N_907,In_996,In_519);
or U908 (N_908,In_1222,In_328);
nor U909 (N_909,In_505,In_423);
or U910 (N_910,In_1232,In_1487);
nor U911 (N_911,In_263,In_188);
or U912 (N_912,In_1122,In_353);
nand U913 (N_913,In_491,In_512);
or U914 (N_914,In_354,In_724);
and U915 (N_915,In_129,In_915);
xnor U916 (N_916,In_1009,In_230);
or U917 (N_917,In_334,In_1296);
nor U918 (N_918,In_273,In_26);
nor U919 (N_919,In_65,In_1474);
and U920 (N_920,In_1423,In_708);
or U921 (N_921,In_1227,In_1465);
nor U922 (N_922,In_960,In_1220);
xnor U923 (N_923,In_485,In_1320);
nand U924 (N_924,In_680,In_1307);
and U925 (N_925,In_61,In_111);
or U926 (N_926,In_1123,In_1139);
xor U927 (N_927,In_161,In_191);
nand U928 (N_928,In_1125,In_137);
nor U929 (N_929,In_260,In_367);
or U930 (N_930,In_1372,In_953);
nand U931 (N_931,In_179,In_604);
or U932 (N_932,In_759,In_318);
xnor U933 (N_933,In_281,In_719);
xnor U934 (N_934,In_1352,In_1495);
nand U935 (N_935,In_1212,In_377);
xnor U936 (N_936,In_1393,In_1427);
or U937 (N_937,In_310,In_876);
and U938 (N_938,In_1056,In_1119);
or U939 (N_939,In_270,In_985);
nor U940 (N_940,In_538,In_19);
and U941 (N_941,In_260,In_797);
or U942 (N_942,In_479,In_934);
nor U943 (N_943,In_459,In_167);
nand U944 (N_944,In_539,In_1002);
or U945 (N_945,In_590,In_1039);
nand U946 (N_946,In_652,In_1019);
nand U947 (N_947,In_744,In_595);
and U948 (N_948,In_812,In_1071);
xnor U949 (N_949,In_111,In_541);
nor U950 (N_950,In_1499,In_377);
or U951 (N_951,In_177,In_233);
or U952 (N_952,In_1306,In_1362);
xor U953 (N_953,In_473,In_122);
nand U954 (N_954,In_112,In_237);
xnor U955 (N_955,In_274,In_429);
xnor U956 (N_956,In_890,In_675);
nand U957 (N_957,In_704,In_100);
nor U958 (N_958,In_1243,In_768);
nor U959 (N_959,In_954,In_610);
or U960 (N_960,In_836,In_727);
xnor U961 (N_961,In_631,In_111);
nand U962 (N_962,In_1316,In_626);
nand U963 (N_963,In_590,In_237);
and U964 (N_964,In_1151,In_228);
xnor U965 (N_965,In_351,In_1320);
and U966 (N_966,In_368,In_274);
or U967 (N_967,In_80,In_1497);
nand U968 (N_968,In_279,In_1432);
or U969 (N_969,In_1302,In_197);
xnor U970 (N_970,In_559,In_185);
nand U971 (N_971,In_171,In_965);
nand U972 (N_972,In_780,In_1278);
or U973 (N_973,In_1103,In_860);
and U974 (N_974,In_1456,In_1450);
xor U975 (N_975,In_565,In_216);
nor U976 (N_976,In_989,In_275);
and U977 (N_977,In_911,In_1251);
and U978 (N_978,In_1405,In_550);
nand U979 (N_979,In_530,In_399);
and U980 (N_980,In_532,In_695);
and U981 (N_981,In_1027,In_990);
or U982 (N_982,In_496,In_116);
or U983 (N_983,In_612,In_406);
nor U984 (N_984,In_1285,In_211);
nand U985 (N_985,In_1285,In_1192);
and U986 (N_986,In_1290,In_113);
xnor U987 (N_987,In_359,In_635);
nor U988 (N_988,In_151,In_732);
nand U989 (N_989,In_658,In_1124);
or U990 (N_990,In_287,In_1416);
xnor U991 (N_991,In_1025,In_102);
nor U992 (N_992,In_1422,In_1033);
and U993 (N_993,In_537,In_575);
nand U994 (N_994,In_268,In_153);
nand U995 (N_995,In_771,In_45);
and U996 (N_996,In_1184,In_1063);
nand U997 (N_997,In_476,In_1371);
or U998 (N_998,In_439,In_142);
nor U999 (N_999,In_359,In_1396);
xnor U1000 (N_1000,In_72,In_1298);
xnor U1001 (N_1001,In_1334,In_452);
nor U1002 (N_1002,In_530,In_1174);
or U1003 (N_1003,In_1315,In_922);
nor U1004 (N_1004,In_1376,In_109);
nor U1005 (N_1005,In_1378,In_229);
nor U1006 (N_1006,In_1177,In_663);
nand U1007 (N_1007,In_237,In_549);
or U1008 (N_1008,In_63,In_657);
or U1009 (N_1009,In_378,In_1165);
nor U1010 (N_1010,In_1223,In_1335);
xor U1011 (N_1011,In_827,In_1104);
xor U1012 (N_1012,In_983,In_1313);
nor U1013 (N_1013,In_230,In_237);
xnor U1014 (N_1014,In_258,In_1458);
xnor U1015 (N_1015,In_277,In_1252);
nor U1016 (N_1016,In_879,In_788);
nand U1017 (N_1017,In_839,In_233);
xor U1018 (N_1018,In_406,In_127);
and U1019 (N_1019,In_1472,In_708);
and U1020 (N_1020,In_1200,In_474);
or U1021 (N_1021,In_399,In_1466);
and U1022 (N_1022,In_468,In_489);
nor U1023 (N_1023,In_361,In_574);
or U1024 (N_1024,In_970,In_300);
nor U1025 (N_1025,In_1123,In_1135);
or U1026 (N_1026,In_637,In_78);
or U1027 (N_1027,In_587,In_716);
and U1028 (N_1028,In_1396,In_1462);
and U1029 (N_1029,In_516,In_846);
xnor U1030 (N_1030,In_949,In_1362);
or U1031 (N_1031,In_317,In_380);
or U1032 (N_1032,In_1027,In_1061);
nand U1033 (N_1033,In_510,In_932);
xor U1034 (N_1034,In_228,In_491);
or U1035 (N_1035,In_1013,In_539);
and U1036 (N_1036,In_1245,In_356);
and U1037 (N_1037,In_1390,In_1401);
and U1038 (N_1038,In_1293,In_1095);
and U1039 (N_1039,In_305,In_174);
nand U1040 (N_1040,In_1420,In_1325);
nor U1041 (N_1041,In_1170,In_895);
and U1042 (N_1042,In_1391,In_1399);
or U1043 (N_1043,In_750,In_1197);
and U1044 (N_1044,In_748,In_63);
or U1045 (N_1045,In_235,In_580);
and U1046 (N_1046,In_749,In_923);
xor U1047 (N_1047,In_798,In_648);
or U1048 (N_1048,In_1338,In_1187);
nor U1049 (N_1049,In_1234,In_560);
nor U1050 (N_1050,In_1063,In_326);
nor U1051 (N_1051,In_184,In_598);
and U1052 (N_1052,In_1432,In_636);
nor U1053 (N_1053,In_1378,In_639);
and U1054 (N_1054,In_928,In_1410);
nand U1055 (N_1055,In_269,In_626);
nor U1056 (N_1056,In_376,In_1013);
and U1057 (N_1057,In_438,In_322);
nand U1058 (N_1058,In_1270,In_1187);
xnor U1059 (N_1059,In_137,In_538);
and U1060 (N_1060,In_1200,In_1105);
nor U1061 (N_1061,In_717,In_926);
and U1062 (N_1062,In_276,In_793);
xor U1063 (N_1063,In_1051,In_568);
nand U1064 (N_1064,In_851,In_723);
and U1065 (N_1065,In_178,In_47);
xnor U1066 (N_1066,In_79,In_331);
nand U1067 (N_1067,In_344,In_1447);
or U1068 (N_1068,In_295,In_1097);
xor U1069 (N_1069,In_903,In_1163);
xor U1070 (N_1070,In_762,In_1156);
and U1071 (N_1071,In_903,In_1479);
and U1072 (N_1072,In_1009,In_1378);
xnor U1073 (N_1073,In_799,In_661);
and U1074 (N_1074,In_2,In_1147);
or U1075 (N_1075,In_962,In_673);
xnor U1076 (N_1076,In_180,In_733);
xor U1077 (N_1077,In_742,In_544);
and U1078 (N_1078,In_1118,In_729);
xor U1079 (N_1079,In_332,In_62);
nand U1080 (N_1080,In_834,In_57);
nand U1081 (N_1081,In_297,In_35);
and U1082 (N_1082,In_59,In_1130);
xnor U1083 (N_1083,In_517,In_542);
or U1084 (N_1084,In_635,In_953);
nand U1085 (N_1085,In_264,In_1059);
nor U1086 (N_1086,In_245,In_39);
xor U1087 (N_1087,In_718,In_1372);
or U1088 (N_1088,In_207,In_224);
and U1089 (N_1089,In_1288,In_1460);
nor U1090 (N_1090,In_686,In_1012);
nor U1091 (N_1091,In_68,In_1344);
or U1092 (N_1092,In_956,In_1481);
nor U1093 (N_1093,In_1467,In_843);
xnor U1094 (N_1094,In_569,In_1198);
or U1095 (N_1095,In_1365,In_173);
nor U1096 (N_1096,In_1233,In_926);
or U1097 (N_1097,In_638,In_1441);
nor U1098 (N_1098,In_627,In_92);
or U1099 (N_1099,In_638,In_632);
nor U1100 (N_1100,In_496,In_18);
nand U1101 (N_1101,In_1098,In_1000);
nor U1102 (N_1102,In_679,In_1385);
or U1103 (N_1103,In_667,In_1143);
nor U1104 (N_1104,In_741,In_219);
and U1105 (N_1105,In_166,In_1047);
or U1106 (N_1106,In_839,In_40);
nor U1107 (N_1107,In_123,In_1010);
and U1108 (N_1108,In_338,In_377);
or U1109 (N_1109,In_111,In_198);
xnor U1110 (N_1110,In_1270,In_801);
and U1111 (N_1111,In_792,In_54);
xor U1112 (N_1112,In_1175,In_85);
nor U1113 (N_1113,In_472,In_883);
xnor U1114 (N_1114,In_1253,In_153);
xnor U1115 (N_1115,In_1175,In_946);
xor U1116 (N_1116,In_1231,In_1362);
nor U1117 (N_1117,In_349,In_567);
xnor U1118 (N_1118,In_365,In_1445);
xor U1119 (N_1119,In_1301,In_1312);
xnor U1120 (N_1120,In_822,In_1312);
and U1121 (N_1121,In_1322,In_675);
or U1122 (N_1122,In_1082,In_654);
nand U1123 (N_1123,In_13,In_1491);
nor U1124 (N_1124,In_1216,In_911);
nor U1125 (N_1125,In_405,In_418);
nand U1126 (N_1126,In_9,In_272);
nand U1127 (N_1127,In_916,In_181);
and U1128 (N_1128,In_946,In_553);
nor U1129 (N_1129,In_1301,In_1061);
xor U1130 (N_1130,In_679,In_129);
nor U1131 (N_1131,In_1181,In_513);
nand U1132 (N_1132,In_1214,In_1036);
xnor U1133 (N_1133,In_1150,In_1059);
or U1134 (N_1134,In_723,In_974);
and U1135 (N_1135,In_344,In_915);
nor U1136 (N_1136,In_970,In_440);
or U1137 (N_1137,In_417,In_1302);
nand U1138 (N_1138,In_524,In_1359);
or U1139 (N_1139,In_1092,In_717);
or U1140 (N_1140,In_717,In_736);
and U1141 (N_1141,In_475,In_932);
nand U1142 (N_1142,In_1198,In_1285);
nor U1143 (N_1143,In_46,In_257);
and U1144 (N_1144,In_447,In_1031);
nand U1145 (N_1145,In_23,In_1096);
xnor U1146 (N_1146,In_85,In_1321);
nand U1147 (N_1147,In_679,In_37);
and U1148 (N_1148,In_1113,In_685);
xor U1149 (N_1149,In_438,In_586);
nor U1150 (N_1150,In_464,In_633);
nand U1151 (N_1151,In_1318,In_105);
nor U1152 (N_1152,In_809,In_511);
xnor U1153 (N_1153,In_1258,In_210);
nor U1154 (N_1154,In_909,In_400);
nand U1155 (N_1155,In_1378,In_31);
nor U1156 (N_1156,In_577,In_1107);
and U1157 (N_1157,In_331,In_1223);
nand U1158 (N_1158,In_753,In_1190);
or U1159 (N_1159,In_546,In_1130);
or U1160 (N_1160,In_342,In_1128);
and U1161 (N_1161,In_163,In_685);
xor U1162 (N_1162,In_1059,In_470);
nor U1163 (N_1163,In_907,In_424);
or U1164 (N_1164,In_75,In_164);
or U1165 (N_1165,In_628,In_1455);
nand U1166 (N_1166,In_1076,In_318);
nor U1167 (N_1167,In_572,In_865);
nand U1168 (N_1168,In_455,In_852);
nor U1169 (N_1169,In_1186,In_1128);
nand U1170 (N_1170,In_677,In_1307);
nor U1171 (N_1171,In_917,In_660);
xor U1172 (N_1172,In_3,In_530);
xnor U1173 (N_1173,In_900,In_309);
and U1174 (N_1174,In_935,In_1151);
xor U1175 (N_1175,In_402,In_859);
and U1176 (N_1176,In_786,In_1472);
nor U1177 (N_1177,In_1443,In_736);
and U1178 (N_1178,In_1449,In_276);
and U1179 (N_1179,In_488,In_1373);
nand U1180 (N_1180,In_146,In_570);
xnor U1181 (N_1181,In_867,In_998);
or U1182 (N_1182,In_950,In_1206);
and U1183 (N_1183,In_1359,In_214);
nor U1184 (N_1184,In_1073,In_166);
nor U1185 (N_1185,In_150,In_1419);
or U1186 (N_1186,In_490,In_950);
nand U1187 (N_1187,In_1454,In_1392);
xnor U1188 (N_1188,In_1363,In_1388);
xnor U1189 (N_1189,In_26,In_84);
nand U1190 (N_1190,In_540,In_1459);
nand U1191 (N_1191,In_1387,In_495);
nor U1192 (N_1192,In_1303,In_434);
nor U1193 (N_1193,In_1071,In_1063);
and U1194 (N_1194,In_378,In_734);
nor U1195 (N_1195,In_270,In_1009);
xor U1196 (N_1196,In_516,In_974);
xor U1197 (N_1197,In_220,In_751);
or U1198 (N_1198,In_453,In_1022);
nor U1199 (N_1199,In_50,In_1428);
xnor U1200 (N_1200,In_1344,In_159);
or U1201 (N_1201,In_1353,In_16);
nand U1202 (N_1202,In_212,In_674);
nor U1203 (N_1203,In_1119,In_1245);
and U1204 (N_1204,In_1461,In_917);
nand U1205 (N_1205,In_575,In_211);
xnor U1206 (N_1206,In_1155,In_1037);
nand U1207 (N_1207,In_888,In_442);
nor U1208 (N_1208,In_719,In_1400);
or U1209 (N_1209,In_7,In_235);
nor U1210 (N_1210,In_783,In_980);
nor U1211 (N_1211,In_404,In_853);
xor U1212 (N_1212,In_456,In_1113);
xor U1213 (N_1213,In_998,In_748);
nor U1214 (N_1214,In_554,In_313);
or U1215 (N_1215,In_1465,In_789);
nand U1216 (N_1216,In_1041,In_1414);
and U1217 (N_1217,In_1278,In_274);
nor U1218 (N_1218,In_289,In_700);
and U1219 (N_1219,In_760,In_273);
nand U1220 (N_1220,In_434,In_903);
xor U1221 (N_1221,In_535,In_774);
nor U1222 (N_1222,In_557,In_128);
nor U1223 (N_1223,In_1419,In_730);
xor U1224 (N_1224,In_293,In_1312);
nand U1225 (N_1225,In_261,In_276);
nand U1226 (N_1226,In_1125,In_1488);
or U1227 (N_1227,In_941,In_777);
nor U1228 (N_1228,In_396,In_139);
or U1229 (N_1229,In_935,In_527);
nor U1230 (N_1230,In_316,In_147);
nor U1231 (N_1231,In_267,In_817);
nor U1232 (N_1232,In_705,In_391);
or U1233 (N_1233,In_567,In_1406);
and U1234 (N_1234,In_1378,In_1172);
xor U1235 (N_1235,In_1404,In_1476);
nor U1236 (N_1236,In_137,In_1083);
xnor U1237 (N_1237,In_221,In_1327);
xnor U1238 (N_1238,In_98,In_747);
nor U1239 (N_1239,In_307,In_1132);
and U1240 (N_1240,In_729,In_277);
or U1241 (N_1241,In_412,In_1177);
nand U1242 (N_1242,In_1307,In_905);
nor U1243 (N_1243,In_1076,In_534);
xor U1244 (N_1244,In_524,In_1430);
or U1245 (N_1245,In_193,In_398);
or U1246 (N_1246,In_799,In_1487);
nand U1247 (N_1247,In_1328,In_881);
and U1248 (N_1248,In_646,In_977);
nor U1249 (N_1249,In_556,In_192);
and U1250 (N_1250,In_793,In_964);
xor U1251 (N_1251,In_319,In_1362);
nand U1252 (N_1252,In_1344,In_406);
or U1253 (N_1253,In_44,In_632);
nand U1254 (N_1254,In_472,In_598);
or U1255 (N_1255,In_1153,In_556);
or U1256 (N_1256,In_826,In_442);
xnor U1257 (N_1257,In_511,In_828);
or U1258 (N_1258,In_845,In_678);
xor U1259 (N_1259,In_767,In_564);
or U1260 (N_1260,In_1022,In_529);
and U1261 (N_1261,In_1245,In_153);
or U1262 (N_1262,In_964,In_328);
and U1263 (N_1263,In_966,In_30);
and U1264 (N_1264,In_1060,In_1191);
nor U1265 (N_1265,In_552,In_6);
xnor U1266 (N_1266,In_1319,In_587);
nand U1267 (N_1267,In_596,In_917);
and U1268 (N_1268,In_1149,In_363);
nand U1269 (N_1269,In_1349,In_1109);
and U1270 (N_1270,In_1151,In_281);
xor U1271 (N_1271,In_1492,In_91);
nand U1272 (N_1272,In_789,In_1498);
nand U1273 (N_1273,In_163,In_29);
nand U1274 (N_1274,In_924,In_768);
xnor U1275 (N_1275,In_328,In_534);
nor U1276 (N_1276,In_337,In_841);
nor U1277 (N_1277,In_691,In_719);
nor U1278 (N_1278,In_816,In_371);
nand U1279 (N_1279,In_419,In_771);
and U1280 (N_1280,In_626,In_1213);
nand U1281 (N_1281,In_882,In_96);
xor U1282 (N_1282,In_1444,In_672);
xor U1283 (N_1283,In_688,In_1091);
or U1284 (N_1284,In_302,In_1409);
or U1285 (N_1285,In_607,In_998);
xnor U1286 (N_1286,In_69,In_1315);
nor U1287 (N_1287,In_1042,In_1252);
and U1288 (N_1288,In_838,In_249);
and U1289 (N_1289,In_1092,In_385);
nand U1290 (N_1290,In_1496,In_1411);
nor U1291 (N_1291,In_985,In_818);
nand U1292 (N_1292,In_141,In_1120);
xnor U1293 (N_1293,In_377,In_332);
xnor U1294 (N_1294,In_1361,In_293);
or U1295 (N_1295,In_440,In_1386);
nor U1296 (N_1296,In_447,In_1010);
and U1297 (N_1297,In_972,In_388);
and U1298 (N_1298,In_325,In_1013);
nor U1299 (N_1299,In_1345,In_1006);
or U1300 (N_1300,In_609,In_206);
and U1301 (N_1301,In_936,In_495);
and U1302 (N_1302,In_1271,In_950);
nor U1303 (N_1303,In_922,In_79);
or U1304 (N_1304,In_759,In_243);
and U1305 (N_1305,In_888,In_1388);
and U1306 (N_1306,In_979,In_146);
nand U1307 (N_1307,In_207,In_1061);
and U1308 (N_1308,In_1262,In_1069);
or U1309 (N_1309,In_1130,In_367);
nor U1310 (N_1310,In_630,In_979);
nor U1311 (N_1311,In_201,In_1133);
nor U1312 (N_1312,In_1255,In_846);
and U1313 (N_1313,In_29,In_571);
nand U1314 (N_1314,In_446,In_1439);
xnor U1315 (N_1315,In_490,In_1487);
xnor U1316 (N_1316,In_1184,In_1047);
or U1317 (N_1317,In_765,In_208);
and U1318 (N_1318,In_890,In_77);
or U1319 (N_1319,In_523,In_21);
nand U1320 (N_1320,In_73,In_804);
nand U1321 (N_1321,In_324,In_764);
xnor U1322 (N_1322,In_652,In_818);
or U1323 (N_1323,In_626,In_221);
and U1324 (N_1324,In_239,In_808);
xor U1325 (N_1325,In_938,In_94);
nor U1326 (N_1326,In_1434,In_1231);
xor U1327 (N_1327,In_1171,In_784);
nand U1328 (N_1328,In_1098,In_814);
and U1329 (N_1329,In_1433,In_182);
xnor U1330 (N_1330,In_681,In_215);
nor U1331 (N_1331,In_1474,In_1217);
xor U1332 (N_1332,In_974,In_840);
nor U1333 (N_1333,In_1178,In_302);
and U1334 (N_1334,In_80,In_358);
or U1335 (N_1335,In_355,In_655);
or U1336 (N_1336,In_856,In_1479);
and U1337 (N_1337,In_853,In_103);
nand U1338 (N_1338,In_900,In_507);
nand U1339 (N_1339,In_92,In_1207);
xor U1340 (N_1340,In_85,In_627);
and U1341 (N_1341,In_1059,In_987);
nand U1342 (N_1342,In_50,In_404);
and U1343 (N_1343,In_730,In_1428);
or U1344 (N_1344,In_54,In_1266);
nand U1345 (N_1345,In_1324,In_129);
nor U1346 (N_1346,In_546,In_418);
or U1347 (N_1347,In_1029,In_1472);
or U1348 (N_1348,In_223,In_779);
nand U1349 (N_1349,In_26,In_956);
or U1350 (N_1350,In_1274,In_1432);
xor U1351 (N_1351,In_1001,In_125);
or U1352 (N_1352,In_19,In_1281);
nor U1353 (N_1353,In_923,In_870);
and U1354 (N_1354,In_984,In_114);
xnor U1355 (N_1355,In_833,In_1146);
or U1356 (N_1356,In_428,In_911);
nand U1357 (N_1357,In_696,In_1426);
or U1358 (N_1358,In_649,In_602);
or U1359 (N_1359,In_946,In_629);
or U1360 (N_1360,In_1188,In_2);
nand U1361 (N_1361,In_71,In_463);
nand U1362 (N_1362,In_1064,In_1357);
and U1363 (N_1363,In_1047,In_660);
nand U1364 (N_1364,In_173,In_1345);
nor U1365 (N_1365,In_169,In_1267);
xnor U1366 (N_1366,In_1398,In_1455);
nor U1367 (N_1367,In_1167,In_899);
xnor U1368 (N_1368,In_1297,In_223);
nor U1369 (N_1369,In_851,In_447);
nand U1370 (N_1370,In_339,In_1378);
or U1371 (N_1371,In_662,In_816);
xor U1372 (N_1372,In_229,In_817);
or U1373 (N_1373,In_49,In_1342);
xnor U1374 (N_1374,In_1048,In_943);
or U1375 (N_1375,In_988,In_1142);
nand U1376 (N_1376,In_285,In_343);
or U1377 (N_1377,In_243,In_104);
and U1378 (N_1378,In_1136,In_1060);
and U1379 (N_1379,In_1148,In_1133);
nand U1380 (N_1380,In_765,In_16);
and U1381 (N_1381,In_467,In_833);
xnor U1382 (N_1382,In_559,In_356);
or U1383 (N_1383,In_1343,In_1226);
nor U1384 (N_1384,In_291,In_189);
or U1385 (N_1385,In_570,In_536);
nand U1386 (N_1386,In_183,In_741);
nor U1387 (N_1387,In_922,In_847);
or U1388 (N_1388,In_979,In_1019);
nand U1389 (N_1389,In_328,In_720);
xor U1390 (N_1390,In_534,In_1020);
nand U1391 (N_1391,In_877,In_75);
nand U1392 (N_1392,In_249,In_1466);
or U1393 (N_1393,In_1283,In_354);
and U1394 (N_1394,In_1499,In_1117);
or U1395 (N_1395,In_638,In_258);
and U1396 (N_1396,In_83,In_1480);
nor U1397 (N_1397,In_761,In_145);
nor U1398 (N_1398,In_101,In_1340);
nor U1399 (N_1399,In_506,In_818);
nor U1400 (N_1400,In_1171,In_481);
xor U1401 (N_1401,In_1491,In_1337);
nor U1402 (N_1402,In_174,In_705);
nor U1403 (N_1403,In_986,In_71);
nor U1404 (N_1404,In_1024,In_317);
xnor U1405 (N_1405,In_438,In_1041);
xnor U1406 (N_1406,In_603,In_296);
or U1407 (N_1407,In_472,In_753);
nand U1408 (N_1408,In_1353,In_1377);
or U1409 (N_1409,In_1209,In_647);
nand U1410 (N_1410,In_323,In_1117);
xor U1411 (N_1411,In_1107,In_1204);
or U1412 (N_1412,In_1481,In_514);
nand U1413 (N_1413,In_496,In_1333);
xor U1414 (N_1414,In_476,In_907);
or U1415 (N_1415,In_333,In_66);
nand U1416 (N_1416,In_1064,In_307);
and U1417 (N_1417,In_968,In_824);
nand U1418 (N_1418,In_746,In_97);
and U1419 (N_1419,In_253,In_1334);
nand U1420 (N_1420,In_1368,In_845);
or U1421 (N_1421,In_966,In_842);
xor U1422 (N_1422,In_1155,In_352);
xor U1423 (N_1423,In_1097,In_714);
or U1424 (N_1424,In_268,In_64);
or U1425 (N_1425,In_868,In_1041);
nand U1426 (N_1426,In_207,In_854);
or U1427 (N_1427,In_606,In_1156);
nand U1428 (N_1428,In_1446,In_1398);
xnor U1429 (N_1429,In_1481,In_406);
or U1430 (N_1430,In_1204,In_123);
xor U1431 (N_1431,In_126,In_870);
nand U1432 (N_1432,In_445,In_372);
nor U1433 (N_1433,In_543,In_110);
or U1434 (N_1434,In_1050,In_105);
xor U1435 (N_1435,In_159,In_976);
or U1436 (N_1436,In_980,In_217);
or U1437 (N_1437,In_98,In_193);
nor U1438 (N_1438,In_334,In_1037);
nand U1439 (N_1439,In_214,In_531);
nand U1440 (N_1440,In_156,In_1009);
nand U1441 (N_1441,In_851,In_1089);
nand U1442 (N_1442,In_674,In_670);
xor U1443 (N_1443,In_30,In_232);
xor U1444 (N_1444,In_913,In_468);
or U1445 (N_1445,In_665,In_613);
xnor U1446 (N_1446,In_724,In_1055);
nor U1447 (N_1447,In_1313,In_266);
and U1448 (N_1448,In_1426,In_997);
and U1449 (N_1449,In_357,In_101);
or U1450 (N_1450,In_414,In_888);
and U1451 (N_1451,In_742,In_402);
nor U1452 (N_1452,In_854,In_1451);
nand U1453 (N_1453,In_1398,In_363);
and U1454 (N_1454,In_1357,In_899);
nand U1455 (N_1455,In_1311,In_304);
nor U1456 (N_1456,In_996,In_399);
xor U1457 (N_1457,In_337,In_1465);
and U1458 (N_1458,In_180,In_1351);
nor U1459 (N_1459,In_1173,In_550);
xor U1460 (N_1460,In_224,In_852);
nand U1461 (N_1461,In_1455,In_377);
and U1462 (N_1462,In_572,In_553);
nand U1463 (N_1463,In_127,In_435);
nor U1464 (N_1464,In_887,In_655);
or U1465 (N_1465,In_21,In_638);
xor U1466 (N_1466,In_71,In_670);
or U1467 (N_1467,In_333,In_1408);
and U1468 (N_1468,In_478,In_598);
and U1469 (N_1469,In_1208,In_326);
and U1470 (N_1470,In_945,In_927);
or U1471 (N_1471,In_146,In_1434);
and U1472 (N_1472,In_1414,In_314);
or U1473 (N_1473,In_485,In_470);
or U1474 (N_1474,In_1306,In_679);
xnor U1475 (N_1475,In_768,In_232);
or U1476 (N_1476,In_720,In_321);
xor U1477 (N_1477,In_241,In_1470);
and U1478 (N_1478,In_302,In_454);
nor U1479 (N_1479,In_1347,In_1100);
or U1480 (N_1480,In_744,In_314);
xnor U1481 (N_1481,In_537,In_1253);
nand U1482 (N_1482,In_1158,In_672);
nand U1483 (N_1483,In_501,In_11);
and U1484 (N_1484,In_719,In_1340);
xor U1485 (N_1485,In_543,In_370);
and U1486 (N_1486,In_1234,In_836);
nand U1487 (N_1487,In_902,In_688);
or U1488 (N_1488,In_1129,In_539);
nor U1489 (N_1489,In_148,In_1130);
nor U1490 (N_1490,In_107,In_285);
and U1491 (N_1491,In_364,In_1470);
nand U1492 (N_1492,In_386,In_523);
nand U1493 (N_1493,In_456,In_928);
or U1494 (N_1494,In_378,In_1004);
nor U1495 (N_1495,In_213,In_1280);
or U1496 (N_1496,In_1447,In_470);
and U1497 (N_1497,In_684,In_566);
nand U1498 (N_1498,In_273,In_1241);
nor U1499 (N_1499,In_511,In_191);
nand U1500 (N_1500,In_1300,In_1131);
nor U1501 (N_1501,In_1423,In_1393);
or U1502 (N_1502,In_579,In_368);
xor U1503 (N_1503,In_781,In_1272);
xnor U1504 (N_1504,In_655,In_1230);
or U1505 (N_1505,In_61,In_643);
nor U1506 (N_1506,In_78,In_272);
nand U1507 (N_1507,In_991,In_740);
xnor U1508 (N_1508,In_1232,In_831);
and U1509 (N_1509,In_400,In_100);
xor U1510 (N_1510,In_800,In_1168);
nor U1511 (N_1511,In_1198,In_172);
xor U1512 (N_1512,In_205,In_566);
nand U1513 (N_1513,In_138,In_1066);
nand U1514 (N_1514,In_1357,In_1038);
nand U1515 (N_1515,In_338,In_1454);
xor U1516 (N_1516,In_665,In_113);
nor U1517 (N_1517,In_714,In_1270);
nor U1518 (N_1518,In_1420,In_131);
nand U1519 (N_1519,In_682,In_1197);
nand U1520 (N_1520,In_385,In_888);
and U1521 (N_1521,In_501,In_759);
or U1522 (N_1522,In_1173,In_312);
xor U1523 (N_1523,In_938,In_1462);
and U1524 (N_1524,In_325,In_828);
nor U1525 (N_1525,In_64,In_820);
nor U1526 (N_1526,In_123,In_498);
xor U1527 (N_1527,In_921,In_495);
nor U1528 (N_1528,In_117,In_526);
nand U1529 (N_1529,In_1152,In_703);
xnor U1530 (N_1530,In_311,In_618);
nand U1531 (N_1531,In_1137,In_204);
xor U1532 (N_1532,In_730,In_359);
and U1533 (N_1533,In_1121,In_99);
xnor U1534 (N_1534,In_207,In_233);
and U1535 (N_1535,In_504,In_245);
nand U1536 (N_1536,In_447,In_404);
nor U1537 (N_1537,In_172,In_977);
nand U1538 (N_1538,In_1479,In_1165);
xor U1539 (N_1539,In_776,In_1351);
xor U1540 (N_1540,In_944,In_1465);
and U1541 (N_1541,In_1132,In_239);
and U1542 (N_1542,In_421,In_1182);
nand U1543 (N_1543,In_1048,In_513);
or U1544 (N_1544,In_870,In_1066);
xor U1545 (N_1545,In_321,In_951);
and U1546 (N_1546,In_826,In_70);
nand U1547 (N_1547,In_1012,In_310);
nand U1548 (N_1548,In_777,In_1061);
nor U1549 (N_1549,In_1253,In_879);
xnor U1550 (N_1550,In_393,In_283);
nand U1551 (N_1551,In_1161,In_933);
nand U1552 (N_1552,In_49,In_896);
and U1553 (N_1553,In_1188,In_550);
and U1554 (N_1554,In_164,In_48);
nand U1555 (N_1555,In_759,In_154);
nor U1556 (N_1556,In_1025,In_1053);
and U1557 (N_1557,In_954,In_655);
xnor U1558 (N_1558,In_669,In_1381);
nand U1559 (N_1559,In_242,In_760);
nand U1560 (N_1560,In_1457,In_674);
and U1561 (N_1561,In_216,In_1409);
and U1562 (N_1562,In_588,In_433);
and U1563 (N_1563,In_496,In_1123);
or U1564 (N_1564,In_1092,In_1314);
nand U1565 (N_1565,In_484,In_664);
nand U1566 (N_1566,In_199,In_1253);
or U1567 (N_1567,In_600,In_1395);
xor U1568 (N_1568,In_29,In_1030);
or U1569 (N_1569,In_783,In_1400);
xor U1570 (N_1570,In_898,In_394);
nor U1571 (N_1571,In_134,In_970);
xnor U1572 (N_1572,In_558,In_1417);
nand U1573 (N_1573,In_571,In_970);
or U1574 (N_1574,In_855,In_124);
nand U1575 (N_1575,In_314,In_480);
nand U1576 (N_1576,In_254,In_1321);
nand U1577 (N_1577,In_439,In_851);
nand U1578 (N_1578,In_88,In_972);
xor U1579 (N_1579,In_465,In_841);
xor U1580 (N_1580,In_1007,In_867);
or U1581 (N_1581,In_601,In_623);
nor U1582 (N_1582,In_296,In_1392);
xor U1583 (N_1583,In_77,In_296);
nor U1584 (N_1584,In_29,In_1489);
or U1585 (N_1585,In_1146,In_266);
or U1586 (N_1586,In_165,In_0);
or U1587 (N_1587,In_597,In_93);
xor U1588 (N_1588,In_665,In_1169);
nor U1589 (N_1589,In_516,In_955);
or U1590 (N_1590,In_1112,In_1478);
or U1591 (N_1591,In_360,In_371);
xnor U1592 (N_1592,In_159,In_911);
nand U1593 (N_1593,In_591,In_930);
xor U1594 (N_1594,In_624,In_1152);
nor U1595 (N_1595,In_1098,In_568);
or U1596 (N_1596,In_440,In_1470);
nand U1597 (N_1597,In_412,In_889);
or U1598 (N_1598,In_1364,In_872);
or U1599 (N_1599,In_568,In_804);
nor U1600 (N_1600,In_1260,In_326);
and U1601 (N_1601,In_797,In_643);
xnor U1602 (N_1602,In_1365,In_766);
or U1603 (N_1603,In_251,In_285);
xnor U1604 (N_1604,In_532,In_1013);
and U1605 (N_1605,In_478,In_893);
nor U1606 (N_1606,In_913,In_397);
nor U1607 (N_1607,In_551,In_1466);
or U1608 (N_1608,In_715,In_31);
nor U1609 (N_1609,In_966,In_346);
and U1610 (N_1610,In_132,In_40);
nor U1611 (N_1611,In_1149,In_827);
xnor U1612 (N_1612,In_1333,In_445);
nor U1613 (N_1613,In_333,In_1022);
or U1614 (N_1614,In_639,In_1432);
nor U1615 (N_1615,In_1414,In_471);
and U1616 (N_1616,In_1066,In_715);
nor U1617 (N_1617,In_1457,In_1456);
or U1618 (N_1618,In_779,In_747);
or U1619 (N_1619,In_525,In_1349);
nand U1620 (N_1620,In_748,In_825);
or U1621 (N_1621,In_1255,In_439);
and U1622 (N_1622,In_255,In_308);
and U1623 (N_1623,In_687,In_700);
xor U1624 (N_1624,In_841,In_873);
and U1625 (N_1625,In_729,In_544);
nor U1626 (N_1626,In_539,In_188);
nand U1627 (N_1627,In_1135,In_1035);
or U1628 (N_1628,In_612,In_978);
nand U1629 (N_1629,In_231,In_661);
or U1630 (N_1630,In_1399,In_355);
nor U1631 (N_1631,In_965,In_915);
and U1632 (N_1632,In_1300,In_1408);
nand U1633 (N_1633,In_1136,In_1093);
xnor U1634 (N_1634,In_303,In_1335);
xnor U1635 (N_1635,In_494,In_1030);
nand U1636 (N_1636,In_657,In_182);
nand U1637 (N_1637,In_1153,In_1315);
xor U1638 (N_1638,In_1247,In_296);
nand U1639 (N_1639,In_832,In_128);
and U1640 (N_1640,In_1204,In_847);
and U1641 (N_1641,In_200,In_546);
and U1642 (N_1642,In_29,In_879);
xnor U1643 (N_1643,In_1139,In_231);
and U1644 (N_1644,In_490,In_732);
and U1645 (N_1645,In_1251,In_1089);
xnor U1646 (N_1646,In_1144,In_1472);
xnor U1647 (N_1647,In_686,In_903);
nor U1648 (N_1648,In_1176,In_494);
xor U1649 (N_1649,In_433,In_42);
xor U1650 (N_1650,In_728,In_479);
xnor U1651 (N_1651,In_419,In_1470);
and U1652 (N_1652,In_621,In_896);
xnor U1653 (N_1653,In_1096,In_315);
nor U1654 (N_1654,In_1188,In_1211);
nor U1655 (N_1655,In_331,In_261);
nor U1656 (N_1656,In_1328,In_958);
and U1657 (N_1657,In_297,In_1110);
nand U1658 (N_1658,In_488,In_831);
or U1659 (N_1659,In_429,In_823);
and U1660 (N_1660,In_784,In_366);
nand U1661 (N_1661,In_65,In_1356);
nor U1662 (N_1662,In_358,In_1424);
and U1663 (N_1663,In_578,In_760);
nand U1664 (N_1664,In_1129,In_1285);
xor U1665 (N_1665,In_381,In_313);
nor U1666 (N_1666,In_1040,In_394);
or U1667 (N_1667,In_1008,In_578);
xnor U1668 (N_1668,In_927,In_1480);
and U1669 (N_1669,In_950,In_920);
nand U1670 (N_1670,In_852,In_762);
and U1671 (N_1671,In_1416,In_946);
and U1672 (N_1672,In_588,In_1057);
or U1673 (N_1673,In_284,In_569);
xnor U1674 (N_1674,In_705,In_1088);
and U1675 (N_1675,In_58,In_186);
nand U1676 (N_1676,In_1047,In_1397);
nand U1677 (N_1677,In_579,In_1174);
and U1678 (N_1678,In_705,In_106);
or U1679 (N_1679,In_576,In_831);
nand U1680 (N_1680,In_458,In_359);
xor U1681 (N_1681,In_51,In_56);
or U1682 (N_1682,In_618,In_1378);
nand U1683 (N_1683,In_997,In_84);
and U1684 (N_1684,In_1188,In_380);
nand U1685 (N_1685,In_1440,In_1477);
nand U1686 (N_1686,In_662,In_183);
and U1687 (N_1687,In_1267,In_84);
nor U1688 (N_1688,In_981,In_1078);
and U1689 (N_1689,In_755,In_249);
nor U1690 (N_1690,In_622,In_422);
or U1691 (N_1691,In_535,In_682);
xor U1692 (N_1692,In_183,In_943);
xor U1693 (N_1693,In_1371,In_1069);
xor U1694 (N_1694,In_22,In_1337);
or U1695 (N_1695,In_178,In_6);
or U1696 (N_1696,In_836,In_1344);
and U1697 (N_1697,In_844,In_409);
nor U1698 (N_1698,In_1011,In_829);
nand U1699 (N_1699,In_773,In_167);
and U1700 (N_1700,In_492,In_1421);
or U1701 (N_1701,In_632,In_1158);
nor U1702 (N_1702,In_50,In_444);
and U1703 (N_1703,In_1321,In_808);
nand U1704 (N_1704,In_1358,In_256);
xnor U1705 (N_1705,In_520,In_1065);
nand U1706 (N_1706,In_1352,In_277);
or U1707 (N_1707,In_923,In_200);
nand U1708 (N_1708,In_1233,In_706);
or U1709 (N_1709,In_661,In_527);
nor U1710 (N_1710,In_146,In_578);
nand U1711 (N_1711,In_176,In_995);
nor U1712 (N_1712,In_88,In_392);
nor U1713 (N_1713,In_113,In_991);
and U1714 (N_1714,In_560,In_1482);
nand U1715 (N_1715,In_62,In_108);
and U1716 (N_1716,In_1386,In_566);
or U1717 (N_1717,In_708,In_864);
nand U1718 (N_1718,In_993,In_117);
xor U1719 (N_1719,In_309,In_643);
nor U1720 (N_1720,In_741,In_618);
nand U1721 (N_1721,In_1276,In_1013);
xnor U1722 (N_1722,In_1243,In_56);
or U1723 (N_1723,In_1029,In_1007);
and U1724 (N_1724,In_982,In_135);
or U1725 (N_1725,In_772,In_1437);
nand U1726 (N_1726,In_1344,In_206);
nand U1727 (N_1727,In_718,In_1264);
or U1728 (N_1728,In_551,In_288);
xnor U1729 (N_1729,In_1116,In_403);
nand U1730 (N_1730,In_838,In_834);
nor U1731 (N_1731,In_375,In_511);
nand U1732 (N_1732,In_1249,In_49);
nand U1733 (N_1733,In_50,In_691);
or U1734 (N_1734,In_1187,In_728);
or U1735 (N_1735,In_837,In_48);
or U1736 (N_1736,In_910,In_1141);
nand U1737 (N_1737,In_860,In_506);
or U1738 (N_1738,In_1307,In_945);
or U1739 (N_1739,In_1234,In_308);
nor U1740 (N_1740,In_1369,In_939);
xor U1741 (N_1741,In_1145,In_1371);
xor U1742 (N_1742,In_1335,In_1013);
xnor U1743 (N_1743,In_62,In_945);
and U1744 (N_1744,In_1330,In_1263);
nor U1745 (N_1745,In_1404,In_635);
nor U1746 (N_1746,In_1262,In_291);
or U1747 (N_1747,In_158,In_510);
nor U1748 (N_1748,In_1408,In_250);
and U1749 (N_1749,In_1148,In_1226);
nand U1750 (N_1750,In_1131,In_1035);
xnor U1751 (N_1751,In_402,In_1159);
xor U1752 (N_1752,In_1004,In_294);
and U1753 (N_1753,In_1157,In_281);
xnor U1754 (N_1754,In_1161,In_454);
and U1755 (N_1755,In_787,In_107);
nor U1756 (N_1756,In_516,In_486);
or U1757 (N_1757,In_1247,In_1302);
nor U1758 (N_1758,In_126,In_722);
or U1759 (N_1759,In_464,In_26);
nand U1760 (N_1760,In_1362,In_1199);
nand U1761 (N_1761,In_443,In_1378);
xnor U1762 (N_1762,In_401,In_795);
or U1763 (N_1763,In_899,In_1315);
or U1764 (N_1764,In_889,In_506);
or U1765 (N_1765,In_523,In_1051);
xor U1766 (N_1766,In_155,In_899);
or U1767 (N_1767,In_10,In_1469);
nor U1768 (N_1768,In_185,In_877);
nand U1769 (N_1769,In_1261,In_304);
nor U1770 (N_1770,In_744,In_428);
nor U1771 (N_1771,In_685,In_1455);
or U1772 (N_1772,In_431,In_367);
nand U1773 (N_1773,In_565,In_1482);
xnor U1774 (N_1774,In_593,In_741);
and U1775 (N_1775,In_221,In_947);
nand U1776 (N_1776,In_76,In_1371);
and U1777 (N_1777,In_642,In_761);
or U1778 (N_1778,In_313,In_915);
or U1779 (N_1779,In_775,In_1200);
nor U1780 (N_1780,In_1413,In_72);
or U1781 (N_1781,In_1036,In_67);
nand U1782 (N_1782,In_168,In_744);
and U1783 (N_1783,In_789,In_846);
nand U1784 (N_1784,In_352,In_1476);
and U1785 (N_1785,In_327,In_235);
nor U1786 (N_1786,In_658,In_1010);
xnor U1787 (N_1787,In_689,In_889);
or U1788 (N_1788,In_1060,In_1182);
nand U1789 (N_1789,In_1124,In_554);
nand U1790 (N_1790,In_360,In_471);
xnor U1791 (N_1791,In_81,In_341);
and U1792 (N_1792,In_596,In_710);
nand U1793 (N_1793,In_1015,In_450);
and U1794 (N_1794,In_1266,In_1038);
and U1795 (N_1795,In_1199,In_932);
or U1796 (N_1796,In_408,In_1397);
nor U1797 (N_1797,In_813,In_37);
or U1798 (N_1798,In_1364,In_1181);
nor U1799 (N_1799,In_938,In_1341);
and U1800 (N_1800,In_98,In_756);
and U1801 (N_1801,In_675,In_1410);
and U1802 (N_1802,In_289,In_186);
and U1803 (N_1803,In_936,In_553);
or U1804 (N_1804,In_561,In_1087);
nor U1805 (N_1805,In_1224,In_1248);
xnor U1806 (N_1806,In_899,In_781);
nand U1807 (N_1807,In_1034,In_896);
and U1808 (N_1808,In_1077,In_707);
nor U1809 (N_1809,In_55,In_789);
xor U1810 (N_1810,In_1027,In_809);
nand U1811 (N_1811,In_486,In_850);
xnor U1812 (N_1812,In_1327,In_777);
nor U1813 (N_1813,In_531,In_107);
xor U1814 (N_1814,In_1141,In_1087);
nand U1815 (N_1815,In_202,In_343);
nor U1816 (N_1816,In_1473,In_525);
xor U1817 (N_1817,In_376,In_269);
nand U1818 (N_1818,In_1007,In_147);
xor U1819 (N_1819,In_720,In_150);
nand U1820 (N_1820,In_1305,In_71);
or U1821 (N_1821,In_1015,In_40);
nor U1822 (N_1822,In_1312,In_490);
nor U1823 (N_1823,In_573,In_1284);
or U1824 (N_1824,In_453,In_136);
nand U1825 (N_1825,In_1438,In_1023);
xor U1826 (N_1826,In_289,In_1273);
nand U1827 (N_1827,In_745,In_216);
or U1828 (N_1828,In_575,In_1343);
and U1829 (N_1829,In_354,In_284);
xor U1830 (N_1830,In_957,In_452);
nand U1831 (N_1831,In_1481,In_213);
nand U1832 (N_1832,In_510,In_735);
nor U1833 (N_1833,In_158,In_960);
nor U1834 (N_1834,In_603,In_1168);
nor U1835 (N_1835,In_1211,In_221);
nand U1836 (N_1836,In_469,In_255);
xor U1837 (N_1837,In_395,In_951);
nor U1838 (N_1838,In_801,In_901);
xnor U1839 (N_1839,In_99,In_1332);
nand U1840 (N_1840,In_1466,In_329);
xor U1841 (N_1841,In_1426,In_197);
nor U1842 (N_1842,In_780,In_345);
and U1843 (N_1843,In_424,In_713);
nand U1844 (N_1844,In_1019,In_425);
nor U1845 (N_1845,In_997,In_502);
xnor U1846 (N_1846,In_201,In_1223);
nand U1847 (N_1847,In_1386,In_289);
nand U1848 (N_1848,In_549,In_1486);
and U1849 (N_1849,In_1458,In_862);
nand U1850 (N_1850,In_880,In_292);
xor U1851 (N_1851,In_788,In_420);
nand U1852 (N_1852,In_1405,In_509);
nor U1853 (N_1853,In_601,In_1270);
nor U1854 (N_1854,In_1079,In_125);
xor U1855 (N_1855,In_113,In_367);
and U1856 (N_1856,In_1212,In_1372);
or U1857 (N_1857,In_661,In_494);
and U1858 (N_1858,In_188,In_455);
nand U1859 (N_1859,In_1490,In_336);
and U1860 (N_1860,In_648,In_564);
and U1861 (N_1861,In_711,In_1015);
xnor U1862 (N_1862,In_112,In_174);
nor U1863 (N_1863,In_359,In_407);
and U1864 (N_1864,In_617,In_1262);
nand U1865 (N_1865,In_1070,In_1257);
nor U1866 (N_1866,In_36,In_44);
or U1867 (N_1867,In_1145,In_1036);
and U1868 (N_1868,In_1352,In_1047);
nor U1869 (N_1869,In_171,In_40);
or U1870 (N_1870,In_998,In_684);
nor U1871 (N_1871,In_1080,In_157);
xnor U1872 (N_1872,In_1481,In_809);
or U1873 (N_1873,In_310,In_1068);
xor U1874 (N_1874,In_716,In_1213);
and U1875 (N_1875,In_137,In_672);
and U1876 (N_1876,In_1452,In_4);
nor U1877 (N_1877,In_918,In_409);
and U1878 (N_1878,In_466,In_1245);
and U1879 (N_1879,In_134,In_456);
or U1880 (N_1880,In_1388,In_1465);
nand U1881 (N_1881,In_508,In_290);
nand U1882 (N_1882,In_1342,In_1324);
xor U1883 (N_1883,In_1134,In_1472);
nand U1884 (N_1884,In_1443,In_191);
xor U1885 (N_1885,In_327,In_1247);
or U1886 (N_1886,In_753,In_562);
and U1887 (N_1887,In_797,In_117);
nor U1888 (N_1888,In_456,In_1148);
nor U1889 (N_1889,In_738,In_585);
nand U1890 (N_1890,In_368,In_1288);
nor U1891 (N_1891,In_1184,In_886);
or U1892 (N_1892,In_863,In_230);
xor U1893 (N_1893,In_1007,In_360);
and U1894 (N_1894,In_124,In_869);
or U1895 (N_1895,In_540,In_829);
or U1896 (N_1896,In_1178,In_152);
xor U1897 (N_1897,In_1038,In_7);
nor U1898 (N_1898,In_638,In_837);
and U1899 (N_1899,In_1091,In_475);
or U1900 (N_1900,In_440,In_923);
nor U1901 (N_1901,In_148,In_1370);
or U1902 (N_1902,In_762,In_1331);
nor U1903 (N_1903,In_183,In_444);
nand U1904 (N_1904,In_1360,In_114);
or U1905 (N_1905,In_795,In_577);
xor U1906 (N_1906,In_650,In_640);
and U1907 (N_1907,In_1247,In_620);
nor U1908 (N_1908,In_1277,In_436);
nand U1909 (N_1909,In_481,In_618);
or U1910 (N_1910,In_910,In_144);
or U1911 (N_1911,In_601,In_447);
xnor U1912 (N_1912,In_264,In_1148);
nand U1913 (N_1913,In_1294,In_785);
and U1914 (N_1914,In_86,In_1201);
xor U1915 (N_1915,In_453,In_694);
nand U1916 (N_1916,In_117,In_998);
or U1917 (N_1917,In_28,In_1122);
xor U1918 (N_1918,In_280,In_1219);
or U1919 (N_1919,In_1475,In_825);
xor U1920 (N_1920,In_1170,In_711);
nor U1921 (N_1921,In_431,In_921);
nor U1922 (N_1922,In_1410,In_346);
nand U1923 (N_1923,In_1155,In_496);
and U1924 (N_1924,In_985,In_976);
nor U1925 (N_1925,In_93,In_97);
or U1926 (N_1926,In_806,In_1314);
or U1927 (N_1927,In_898,In_1323);
xor U1928 (N_1928,In_146,In_1483);
and U1929 (N_1929,In_800,In_1479);
nand U1930 (N_1930,In_361,In_111);
nor U1931 (N_1931,In_395,In_255);
and U1932 (N_1932,In_723,In_295);
nor U1933 (N_1933,In_969,In_268);
nor U1934 (N_1934,In_840,In_367);
nor U1935 (N_1935,In_1017,In_1364);
or U1936 (N_1936,In_922,In_18);
nor U1937 (N_1937,In_849,In_1450);
nor U1938 (N_1938,In_307,In_678);
or U1939 (N_1939,In_1332,In_526);
nor U1940 (N_1940,In_750,In_1201);
nand U1941 (N_1941,In_730,In_1207);
or U1942 (N_1942,In_605,In_642);
or U1943 (N_1943,In_990,In_1462);
xnor U1944 (N_1944,In_766,In_899);
nor U1945 (N_1945,In_1076,In_880);
nor U1946 (N_1946,In_1433,In_173);
and U1947 (N_1947,In_239,In_940);
or U1948 (N_1948,In_291,In_1001);
nand U1949 (N_1949,In_1416,In_706);
xor U1950 (N_1950,In_568,In_1016);
and U1951 (N_1951,In_720,In_71);
or U1952 (N_1952,In_1033,In_1009);
and U1953 (N_1953,In_297,In_107);
nor U1954 (N_1954,In_417,In_189);
nor U1955 (N_1955,In_1428,In_768);
xor U1956 (N_1956,In_1047,In_1167);
or U1957 (N_1957,In_937,In_612);
nand U1958 (N_1958,In_101,In_254);
and U1959 (N_1959,In_983,In_1072);
nor U1960 (N_1960,In_606,In_1130);
nand U1961 (N_1961,In_11,In_164);
xnor U1962 (N_1962,In_260,In_1242);
xor U1963 (N_1963,In_832,In_730);
nor U1964 (N_1964,In_168,In_394);
and U1965 (N_1965,In_380,In_196);
xnor U1966 (N_1966,In_1248,In_133);
xnor U1967 (N_1967,In_1255,In_1412);
xor U1968 (N_1968,In_512,In_511);
or U1969 (N_1969,In_1470,In_1112);
nor U1970 (N_1970,In_562,In_228);
nor U1971 (N_1971,In_519,In_602);
xor U1972 (N_1972,In_1380,In_938);
nand U1973 (N_1973,In_252,In_404);
nor U1974 (N_1974,In_1268,In_754);
and U1975 (N_1975,In_1283,In_414);
nand U1976 (N_1976,In_721,In_1254);
nand U1977 (N_1977,In_496,In_1238);
xnor U1978 (N_1978,In_362,In_315);
xnor U1979 (N_1979,In_512,In_1475);
xnor U1980 (N_1980,In_1189,In_1420);
nand U1981 (N_1981,In_1003,In_1164);
nor U1982 (N_1982,In_484,In_673);
nor U1983 (N_1983,In_136,In_1396);
nor U1984 (N_1984,In_1351,In_739);
xnor U1985 (N_1985,In_343,In_930);
or U1986 (N_1986,In_1433,In_448);
and U1987 (N_1987,In_1258,In_1238);
or U1988 (N_1988,In_660,In_909);
nor U1989 (N_1989,In_732,In_1414);
nand U1990 (N_1990,In_1084,In_58);
nor U1991 (N_1991,In_52,In_1254);
xor U1992 (N_1992,In_1351,In_152);
xor U1993 (N_1993,In_300,In_1039);
nand U1994 (N_1994,In_144,In_1227);
and U1995 (N_1995,In_377,In_897);
nand U1996 (N_1996,In_691,In_1242);
and U1997 (N_1997,In_276,In_543);
or U1998 (N_1998,In_514,In_411);
or U1999 (N_1999,In_472,In_776);
and U2000 (N_2000,In_768,In_115);
and U2001 (N_2001,In_1300,In_683);
or U2002 (N_2002,In_630,In_335);
xor U2003 (N_2003,In_1124,In_47);
nor U2004 (N_2004,In_345,In_946);
xnor U2005 (N_2005,In_867,In_1473);
and U2006 (N_2006,In_1,In_560);
and U2007 (N_2007,In_983,In_728);
or U2008 (N_2008,In_1370,In_1122);
nand U2009 (N_2009,In_858,In_1343);
xor U2010 (N_2010,In_90,In_1410);
and U2011 (N_2011,In_1311,In_788);
nor U2012 (N_2012,In_1179,In_820);
or U2013 (N_2013,In_164,In_212);
or U2014 (N_2014,In_366,In_979);
nor U2015 (N_2015,In_1079,In_188);
nand U2016 (N_2016,In_832,In_1469);
nand U2017 (N_2017,In_174,In_1168);
nor U2018 (N_2018,In_665,In_642);
nand U2019 (N_2019,In_1351,In_1480);
xor U2020 (N_2020,In_1192,In_615);
or U2021 (N_2021,In_147,In_862);
and U2022 (N_2022,In_881,In_22);
nor U2023 (N_2023,In_1473,In_945);
and U2024 (N_2024,In_780,In_1374);
nor U2025 (N_2025,In_12,In_1330);
xnor U2026 (N_2026,In_1353,In_454);
or U2027 (N_2027,In_397,In_1348);
nand U2028 (N_2028,In_853,In_263);
nor U2029 (N_2029,In_592,In_1128);
and U2030 (N_2030,In_272,In_216);
nor U2031 (N_2031,In_940,In_997);
and U2032 (N_2032,In_704,In_680);
xor U2033 (N_2033,In_476,In_1476);
nor U2034 (N_2034,In_130,In_671);
or U2035 (N_2035,In_876,In_725);
nor U2036 (N_2036,In_773,In_124);
nor U2037 (N_2037,In_1494,In_1321);
nor U2038 (N_2038,In_561,In_536);
xor U2039 (N_2039,In_74,In_774);
nand U2040 (N_2040,In_539,In_803);
or U2041 (N_2041,In_1354,In_1180);
nand U2042 (N_2042,In_1013,In_1191);
or U2043 (N_2043,In_33,In_1236);
or U2044 (N_2044,In_924,In_483);
xor U2045 (N_2045,In_743,In_1225);
or U2046 (N_2046,In_350,In_9);
nor U2047 (N_2047,In_1003,In_648);
nor U2048 (N_2048,In_775,In_953);
or U2049 (N_2049,In_455,In_425);
xnor U2050 (N_2050,In_476,In_1120);
and U2051 (N_2051,In_480,In_457);
nand U2052 (N_2052,In_760,In_244);
or U2053 (N_2053,In_526,In_83);
nand U2054 (N_2054,In_1272,In_451);
nand U2055 (N_2055,In_378,In_1025);
and U2056 (N_2056,In_221,In_577);
nand U2057 (N_2057,In_1321,In_790);
and U2058 (N_2058,In_1355,In_990);
or U2059 (N_2059,In_981,In_1086);
nor U2060 (N_2060,In_141,In_409);
nor U2061 (N_2061,In_872,In_1261);
xor U2062 (N_2062,In_745,In_1038);
nand U2063 (N_2063,In_502,In_425);
xnor U2064 (N_2064,In_1485,In_1321);
nor U2065 (N_2065,In_234,In_269);
nand U2066 (N_2066,In_434,In_801);
and U2067 (N_2067,In_192,In_152);
and U2068 (N_2068,In_810,In_649);
and U2069 (N_2069,In_461,In_1013);
or U2070 (N_2070,In_482,In_185);
nor U2071 (N_2071,In_1229,In_1212);
xor U2072 (N_2072,In_915,In_904);
nor U2073 (N_2073,In_1181,In_1147);
or U2074 (N_2074,In_728,In_408);
xnor U2075 (N_2075,In_536,In_207);
nand U2076 (N_2076,In_450,In_304);
nand U2077 (N_2077,In_932,In_409);
and U2078 (N_2078,In_432,In_827);
and U2079 (N_2079,In_1431,In_1048);
nand U2080 (N_2080,In_630,In_611);
or U2081 (N_2081,In_1374,In_650);
or U2082 (N_2082,In_1396,In_1112);
xor U2083 (N_2083,In_23,In_153);
and U2084 (N_2084,In_570,In_205);
and U2085 (N_2085,In_569,In_688);
or U2086 (N_2086,In_858,In_1434);
and U2087 (N_2087,In_1396,In_827);
and U2088 (N_2088,In_1142,In_466);
and U2089 (N_2089,In_65,In_298);
or U2090 (N_2090,In_280,In_758);
and U2091 (N_2091,In_1326,In_43);
and U2092 (N_2092,In_1281,In_853);
nand U2093 (N_2093,In_1276,In_503);
and U2094 (N_2094,In_138,In_1241);
and U2095 (N_2095,In_657,In_1356);
nand U2096 (N_2096,In_1460,In_408);
and U2097 (N_2097,In_411,In_1063);
xor U2098 (N_2098,In_1101,In_406);
or U2099 (N_2099,In_429,In_1274);
nor U2100 (N_2100,In_120,In_699);
xnor U2101 (N_2101,In_1209,In_879);
and U2102 (N_2102,In_1144,In_207);
or U2103 (N_2103,In_260,In_1331);
or U2104 (N_2104,In_14,In_1199);
nand U2105 (N_2105,In_1389,In_543);
xor U2106 (N_2106,In_910,In_274);
nand U2107 (N_2107,In_313,In_1290);
nand U2108 (N_2108,In_945,In_384);
nor U2109 (N_2109,In_412,In_695);
or U2110 (N_2110,In_43,In_520);
and U2111 (N_2111,In_916,In_354);
xor U2112 (N_2112,In_293,In_712);
nand U2113 (N_2113,In_669,In_1098);
nand U2114 (N_2114,In_1368,In_1371);
and U2115 (N_2115,In_750,In_752);
or U2116 (N_2116,In_1236,In_782);
and U2117 (N_2117,In_87,In_192);
xnor U2118 (N_2118,In_976,In_686);
xor U2119 (N_2119,In_377,In_80);
and U2120 (N_2120,In_253,In_132);
or U2121 (N_2121,In_1320,In_1353);
or U2122 (N_2122,In_1413,In_644);
xor U2123 (N_2123,In_371,In_617);
nand U2124 (N_2124,In_262,In_175);
nand U2125 (N_2125,In_1029,In_1182);
nor U2126 (N_2126,In_1075,In_871);
xnor U2127 (N_2127,In_1390,In_567);
xor U2128 (N_2128,In_1130,In_1473);
nor U2129 (N_2129,In_412,In_1393);
or U2130 (N_2130,In_1033,In_1134);
nand U2131 (N_2131,In_1497,In_765);
xor U2132 (N_2132,In_1262,In_276);
or U2133 (N_2133,In_314,In_335);
xor U2134 (N_2134,In_289,In_1023);
nor U2135 (N_2135,In_1392,In_466);
nor U2136 (N_2136,In_447,In_1001);
nor U2137 (N_2137,In_71,In_1417);
xor U2138 (N_2138,In_1243,In_1416);
nor U2139 (N_2139,In_320,In_929);
xnor U2140 (N_2140,In_633,In_774);
nor U2141 (N_2141,In_334,In_583);
and U2142 (N_2142,In_122,In_775);
xnor U2143 (N_2143,In_1235,In_734);
nand U2144 (N_2144,In_1287,In_199);
nor U2145 (N_2145,In_1259,In_13);
or U2146 (N_2146,In_456,In_306);
and U2147 (N_2147,In_5,In_726);
or U2148 (N_2148,In_1315,In_1190);
xnor U2149 (N_2149,In_502,In_399);
or U2150 (N_2150,In_1158,In_1440);
nor U2151 (N_2151,In_1359,In_917);
xor U2152 (N_2152,In_743,In_1430);
and U2153 (N_2153,In_1205,In_952);
xor U2154 (N_2154,In_870,In_816);
nand U2155 (N_2155,In_838,In_980);
xnor U2156 (N_2156,In_284,In_846);
and U2157 (N_2157,In_165,In_1416);
nand U2158 (N_2158,In_614,In_1497);
nand U2159 (N_2159,In_1456,In_381);
nand U2160 (N_2160,In_7,In_120);
or U2161 (N_2161,In_930,In_426);
nor U2162 (N_2162,In_1444,In_478);
and U2163 (N_2163,In_616,In_1400);
and U2164 (N_2164,In_721,In_1472);
nand U2165 (N_2165,In_942,In_169);
and U2166 (N_2166,In_690,In_202);
and U2167 (N_2167,In_207,In_1221);
and U2168 (N_2168,In_414,In_274);
and U2169 (N_2169,In_240,In_1383);
nand U2170 (N_2170,In_1383,In_927);
xor U2171 (N_2171,In_776,In_186);
nor U2172 (N_2172,In_1428,In_938);
or U2173 (N_2173,In_272,In_1442);
nand U2174 (N_2174,In_652,In_1189);
nor U2175 (N_2175,In_1466,In_1191);
xnor U2176 (N_2176,In_1311,In_634);
xor U2177 (N_2177,In_330,In_901);
nand U2178 (N_2178,In_727,In_135);
nand U2179 (N_2179,In_796,In_1383);
or U2180 (N_2180,In_460,In_225);
nor U2181 (N_2181,In_1357,In_4);
xnor U2182 (N_2182,In_496,In_616);
xor U2183 (N_2183,In_1351,In_880);
or U2184 (N_2184,In_508,In_500);
nand U2185 (N_2185,In_417,In_823);
nand U2186 (N_2186,In_1292,In_1268);
xnor U2187 (N_2187,In_266,In_1453);
nand U2188 (N_2188,In_274,In_743);
or U2189 (N_2189,In_1079,In_1453);
or U2190 (N_2190,In_274,In_53);
nor U2191 (N_2191,In_143,In_448);
nor U2192 (N_2192,In_386,In_528);
or U2193 (N_2193,In_338,In_1372);
xor U2194 (N_2194,In_425,In_1393);
xnor U2195 (N_2195,In_587,In_250);
xnor U2196 (N_2196,In_61,In_1249);
and U2197 (N_2197,In_1054,In_545);
and U2198 (N_2198,In_1040,In_728);
xor U2199 (N_2199,In_784,In_1173);
or U2200 (N_2200,In_1232,In_927);
nor U2201 (N_2201,In_48,In_198);
or U2202 (N_2202,In_213,In_643);
or U2203 (N_2203,In_1497,In_769);
and U2204 (N_2204,In_796,In_1407);
or U2205 (N_2205,In_470,In_127);
or U2206 (N_2206,In_19,In_1158);
xnor U2207 (N_2207,In_976,In_1368);
xnor U2208 (N_2208,In_441,In_842);
nor U2209 (N_2209,In_1432,In_421);
and U2210 (N_2210,In_406,In_1356);
nor U2211 (N_2211,In_147,In_1060);
or U2212 (N_2212,In_1389,In_366);
nand U2213 (N_2213,In_29,In_1420);
xnor U2214 (N_2214,In_1326,In_1120);
or U2215 (N_2215,In_544,In_475);
nand U2216 (N_2216,In_1272,In_1037);
xor U2217 (N_2217,In_89,In_24);
nand U2218 (N_2218,In_225,In_1143);
xor U2219 (N_2219,In_486,In_1162);
nor U2220 (N_2220,In_190,In_1499);
nand U2221 (N_2221,In_148,In_1338);
nand U2222 (N_2222,In_883,In_328);
nor U2223 (N_2223,In_903,In_412);
and U2224 (N_2224,In_22,In_1009);
nand U2225 (N_2225,In_611,In_777);
xor U2226 (N_2226,In_1437,In_353);
xnor U2227 (N_2227,In_998,In_75);
or U2228 (N_2228,In_1099,In_1421);
or U2229 (N_2229,In_472,In_656);
xnor U2230 (N_2230,In_890,In_558);
nand U2231 (N_2231,In_1354,In_1267);
or U2232 (N_2232,In_1288,In_260);
nor U2233 (N_2233,In_1497,In_588);
or U2234 (N_2234,In_770,In_549);
and U2235 (N_2235,In_38,In_278);
xnor U2236 (N_2236,In_1155,In_445);
xnor U2237 (N_2237,In_1090,In_21);
nor U2238 (N_2238,In_730,In_767);
xnor U2239 (N_2239,In_1213,In_695);
and U2240 (N_2240,In_264,In_432);
nand U2241 (N_2241,In_301,In_1140);
or U2242 (N_2242,In_1114,In_785);
or U2243 (N_2243,In_369,In_1391);
or U2244 (N_2244,In_112,In_708);
xnor U2245 (N_2245,In_1298,In_850);
nand U2246 (N_2246,In_769,In_500);
nor U2247 (N_2247,In_1290,In_1064);
nor U2248 (N_2248,In_1411,In_498);
nor U2249 (N_2249,In_1181,In_653);
nor U2250 (N_2250,In_213,In_440);
or U2251 (N_2251,In_1031,In_775);
nand U2252 (N_2252,In_38,In_1319);
nor U2253 (N_2253,In_1412,In_1448);
nor U2254 (N_2254,In_126,In_886);
or U2255 (N_2255,In_1312,In_902);
nand U2256 (N_2256,In_1057,In_1026);
nor U2257 (N_2257,In_1318,In_1183);
nand U2258 (N_2258,In_1447,In_1120);
xor U2259 (N_2259,In_531,In_1066);
or U2260 (N_2260,In_1170,In_239);
xnor U2261 (N_2261,In_1443,In_311);
nor U2262 (N_2262,In_972,In_689);
or U2263 (N_2263,In_986,In_364);
nand U2264 (N_2264,In_646,In_797);
nor U2265 (N_2265,In_383,In_613);
nor U2266 (N_2266,In_866,In_532);
xnor U2267 (N_2267,In_1356,In_868);
or U2268 (N_2268,In_1090,In_1058);
and U2269 (N_2269,In_1045,In_1456);
or U2270 (N_2270,In_1292,In_600);
or U2271 (N_2271,In_427,In_51);
nand U2272 (N_2272,In_1142,In_628);
and U2273 (N_2273,In_430,In_1120);
and U2274 (N_2274,In_1335,In_553);
or U2275 (N_2275,In_459,In_1171);
and U2276 (N_2276,In_946,In_1376);
xor U2277 (N_2277,In_1045,In_435);
nand U2278 (N_2278,In_959,In_31);
nand U2279 (N_2279,In_1087,In_490);
and U2280 (N_2280,In_874,In_192);
or U2281 (N_2281,In_1134,In_619);
or U2282 (N_2282,In_151,In_1384);
nor U2283 (N_2283,In_914,In_162);
and U2284 (N_2284,In_1098,In_878);
nand U2285 (N_2285,In_416,In_1199);
nor U2286 (N_2286,In_1363,In_1205);
nor U2287 (N_2287,In_496,In_10);
or U2288 (N_2288,In_540,In_1160);
and U2289 (N_2289,In_989,In_366);
nand U2290 (N_2290,In_891,In_738);
or U2291 (N_2291,In_161,In_513);
or U2292 (N_2292,In_687,In_936);
nand U2293 (N_2293,In_1049,In_471);
and U2294 (N_2294,In_989,In_516);
nand U2295 (N_2295,In_184,In_1048);
nor U2296 (N_2296,In_506,In_867);
xnor U2297 (N_2297,In_1122,In_335);
nor U2298 (N_2298,In_627,In_1094);
nor U2299 (N_2299,In_1076,In_773);
nand U2300 (N_2300,In_1314,In_14);
xnor U2301 (N_2301,In_1206,In_1236);
nand U2302 (N_2302,In_1019,In_1338);
xor U2303 (N_2303,In_846,In_201);
and U2304 (N_2304,In_1481,In_1425);
nor U2305 (N_2305,In_448,In_470);
and U2306 (N_2306,In_147,In_1089);
xor U2307 (N_2307,In_688,In_74);
nand U2308 (N_2308,In_1021,In_1225);
and U2309 (N_2309,In_827,In_286);
or U2310 (N_2310,In_110,In_414);
or U2311 (N_2311,In_1256,In_1077);
xnor U2312 (N_2312,In_791,In_161);
or U2313 (N_2313,In_1017,In_869);
nor U2314 (N_2314,In_870,In_896);
nand U2315 (N_2315,In_328,In_1396);
or U2316 (N_2316,In_44,In_1388);
or U2317 (N_2317,In_936,In_638);
and U2318 (N_2318,In_850,In_93);
nor U2319 (N_2319,In_181,In_923);
xor U2320 (N_2320,In_79,In_1034);
or U2321 (N_2321,In_961,In_508);
nor U2322 (N_2322,In_867,In_533);
nor U2323 (N_2323,In_167,In_1148);
and U2324 (N_2324,In_188,In_1456);
xor U2325 (N_2325,In_1394,In_660);
nand U2326 (N_2326,In_51,In_144);
nand U2327 (N_2327,In_364,In_328);
and U2328 (N_2328,In_782,In_18);
and U2329 (N_2329,In_200,In_8);
nor U2330 (N_2330,In_663,In_465);
nand U2331 (N_2331,In_390,In_599);
nand U2332 (N_2332,In_294,In_503);
nand U2333 (N_2333,In_1117,In_14);
nor U2334 (N_2334,In_1324,In_1066);
xnor U2335 (N_2335,In_729,In_350);
nor U2336 (N_2336,In_863,In_266);
or U2337 (N_2337,In_1494,In_1153);
nor U2338 (N_2338,In_1489,In_256);
or U2339 (N_2339,In_1167,In_220);
and U2340 (N_2340,In_789,In_284);
or U2341 (N_2341,In_1088,In_1386);
nand U2342 (N_2342,In_236,In_1193);
xor U2343 (N_2343,In_656,In_1038);
or U2344 (N_2344,In_978,In_873);
xnor U2345 (N_2345,In_950,In_476);
or U2346 (N_2346,In_587,In_1363);
nand U2347 (N_2347,In_260,In_524);
nand U2348 (N_2348,In_1254,In_84);
nor U2349 (N_2349,In_479,In_426);
nor U2350 (N_2350,In_257,In_611);
or U2351 (N_2351,In_345,In_529);
xor U2352 (N_2352,In_95,In_1304);
nor U2353 (N_2353,In_531,In_450);
nor U2354 (N_2354,In_1011,In_97);
and U2355 (N_2355,In_477,In_1267);
nand U2356 (N_2356,In_324,In_528);
xnor U2357 (N_2357,In_665,In_441);
nor U2358 (N_2358,In_204,In_357);
nand U2359 (N_2359,In_830,In_274);
or U2360 (N_2360,In_770,In_1030);
xnor U2361 (N_2361,In_710,In_1047);
and U2362 (N_2362,In_744,In_431);
nor U2363 (N_2363,In_1154,In_1066);
and U2364 (N_2364,In_232,In_896);
nor U2365 (N_2365,In_82,In_17);
or U2366 (N_2366,In_726,In_1333);
and U2367 (N_2367,In_1348,In_1156);
nor U2368 (N_2368,In_418,In_1469);
and U2369 (N_2369,In_1193,In_146);
xnor U2370 (N_2370,In_1419,In_287);
xnor U2371 (N_2371,In_573,In_466);
or U2372 (N_2372,In_464,In_552);
and U2373 (N_2373,In_779,In_1030);
xnor U2374 (N_2374,In_879,In_31);
or U2375 (N_2375,In_819,In_748);
xnor U2376 (N_2376,In_535,In_989);
nand U2377 (N_2377,In_828,In_1427);
nor U2378 (N_2378,In_1169,In_1173);
or U2379 (N_2379,In_940,In_268);
nand U2380 (N_2380,In_721,In_347);
or U2381 (N_2381,In_91,In_1402);
and U2382 (N_2382,In_648,In_212);
nand U2383 (N_2383,In_470,In_1486);
nor U2384 (N_2384,In_597,In_1182);
xnor U2385 (N_2385,In_807,In_902);
or U2386 (N_2386,In_1024,In_82);
and U2387 (N_2387,In_1043,In_398);
nor U2388 (N_2388,In_20,In_951);
xnor U2389 (N_2389,In_1381,In_1250);
xor U2390 (N_2390,In_1426,In_1387);
xor U2391 (N_2391,In_1223,In_257);
and U2392 (N_2392,In_1003,In_833);
xnor U2393 (N_2393,In_1036,In_125);
nand U2394 (N_2394,In_1227,In_1133);
and U2395 (N_2395,In_1340,In_983);
xnor U2396 (N_2396,In_1094,In_1273);
xnor U2397 (N_2397,In_335,In_863);
and U2398 (N_2398,In_1155,In_127);
nor U2399 (N_2399,In_67,In_832);
xnor U2400 (N_2400,In_1254,In_274);
nand U2401 (N_2401,In_1221,In_288);
and U2402 (N_2402,In_685,In_149);
or U2403 (N_2403,In_1239,In_437);
nor U2404 (N_2404,In_1343,In_1208);
nor U2405 (N_2405,In_1480,In_326);
xor U2406 (N_2406,In_1204,In_526);
nor U2407 (N_2407,In_659,In_275);
xor U2408 (N_2408,In_56,In_1149);
and U2409 (N_2409,In_1070,In_1485);
nand U2410 (N_2410,In_90,In_976);
xor U2411 (N_2411,In_1370,In_156);
nand U2412 (N_2412,In_972,In_258);
nor U2413 (N_2413,In_635,In_297);
nor U2414 (N_2414,In_466,In_5);
nor U2415 (N_2415,In_664,In_746);
xnor U2416 (N_2416,In_129,In_1124);
and U2417 (N_2417,In_1230,In_1040);
nand U2418 (N_2418,In_277,In_1102);
nand U2419 (N_2419,In_1268,In_802);
nand U2420 (N_2420,In_216,In_195);
nor U2421 (N_2421,In_1363,In_105);
or U2422 (N_2422,In_870,In_519);
xor U2423 (N_2423,In_511,In_712);
xnor U2424 (N_2424,In_341,In_1235);
or U2425 (N_2425,In_608,In_96);
nand U2426 (N_2426,In_302,In_666);
nand U2427 (N_2427,In_175,In_665);
or U2428 (N_2428,In_690,In_80);
nand U2429 (N_2429,In_310,In_657);
and U2430 (N_2430,In_950,In_917);
xor U2431 (N_2431,In_790,In_453);
and U2432 (N_2432,In_889,In_900);
nor U2433 (N_2433,In_1409,In_599);
nand U2434 (N_2434,In_1466,In_369);
and U2435 (N_2435,In_642,In_615);
and U2436 (N_2436,In_583,In_1426);
nand U2437 (N_2437,In_782,In_251);
nand U2438 (N_2438,In_874,In_421);
and U2439 (N_2439,In_442,In_1061);
or U2440 (N_2440,In_113,In_424);
xor U2441 (N_2441,In_1125,In_1280);
and U2442 (N_2442,In_221,In_895);
xor U2443 (N_2443,In_63,In_653);
nand U2444 (N_2444,In_697,In_3);
or U2445 (N_2445,In_1297,In_1383);
xor U2446 (N_2446,In_241,In_4);
xnor U2447 (N_2447,In_104,In_732);
nor U2448 (N_2448,In_1293,In_1124);
and U2449 (N_2449,In_1229,In_535);
xor U2450 (N_2450,In_9,In_1208);
and U2451 (N_2451,In_693,In_781);
or U2452 (N_2452,In_421,In_719);
and U2453 (N_2453,In_807,In_1385);
nor U2454 (N_2454,In_1057,In_845);
or U2455 (N_2455,In_566,In_381);
xor U2456 (N_2456,In_279,In_821);
nor U2457 (N_2457,In_496,In_1312);
nor U2458 (N_2458,In_502,In_445);
nand U2459 (N_2459,In_283,In_157);
or U2460 (N_2460,In_918,In_173);
xnor U2461 (N_2461,In_1309,In_158);
nor U2462 (N_2462,In_1326,In_1420);
and U2463 (N_2463,In_238,In_452);
nor U2464 (N_2464,In_887,In_952);
or U2465 (N_2465,In_766,In_1436);
nor U2466 (N_2466,In_1223,In_169);
or U2467 (N_2467,In_952,In_163);
nor U2468 (N_2468,In_1014,In_15);
nor U2469 (N_2469,In_1318,In_996);
nor U2470 (N_2470,In_61,In_1412);
and U2471 (N_2471,In_896,In_704);
or U2472 (N_2472,In_245,In_992);
xnor U2473 (N_2473,In_907,In_21);
nor U2474 (N_2474,In_1448,In_1257);
xor U2475 (N_2475,In_1337,In_1080);
and U2476 (N_2476,In_909,In_887);
xnor U2477 (N_2477,In_216,In_1118);
and U2478 (N_2478,In_89,In_1080);
nor U2479 (N_2479,In_1,In_294);
nand U2480 (N_2480,In_860,In_823);
nor U2481 (N_2481,In_1182,In_129);
xnor U2482 (N_2482,In_1327,In_28);
or U2483 (N_2483,In_1029,In_91);
or U2484 (N_2484,In_921,In_266);
and U2485 (N_2485,In_1022,In_1484);
xnor U2486 (N_2486,In_1380,In_710);
or U2487 (N_2487,In_1366,In_1061);
xor U2488 (N_2488,In_815,In_623);
nand U2489 (N_2489,In_117,In_1486);
or U2490 (N_2490,In_811,In_1140);
and U2491 (N_2491,In_1392,In_1316);
and U2492 (N_2492,In_1175,In_591);
nor U2493 (N_2493,In_428,In_476);
and U2494 (N_2494,In_960,In_1149);
nor U2495 (N_2495,In_497,In_1425);
nand U2496 (N_2496,In_778,In_1386);
and U2497 (N_2497,In_949,In_160);
and U2498 (N_2498,In_1368,In_902);
and U2499 (N_2499,In_447,In_945);
nor U2500 (N_2500,In_1163,In_1337);
xor U2501 (N_2501,In_288,In_82);
nor U2502 (N_2502,In_130,In_377);
nand U2503 (N_2503,In_1148,In_1127);
and U2504 (N_2504,In_1294,In_671);
and U2505 (N_2505,In_919,In_1476);
nand U2506 (N_2506,In_167,In_338);
or U2507 (N_2507,In_999,In_1020);
xnor U2508 (N_2508,In_643,In_1059);
nand U2509 (N_2509,In_625,In_877);
nor U2510 (N_2510,In_826,In_178);
and U2511 (N_2511,In_606,In_1084);
and U2512 (N_2512,In_665,In_1073);
and U2513 (N_2513,In_857,In_1388);
nor U2514 (N_2514,In_1204,In_132);
xor U2515 (N_2515,In_1017,In_1023);
and U2516 (N_2516,In_1232,In_991);
xnor U2517 (N_2517,In_576,In_1101);
and U2518 (N_2518,In_157,In_986);
or U2519 (N_2519,In_435,In_371);
nand U2520 (N_2520,In_1398,In_623);
or U2521 (N_2521,In_905,In_399);
nor U2522 (N_2522,In_691,In_1378);
nand U2523 (N_2523,In_467,In_568);
and U2524 (N_2524,In_1273,In_295);
nand U2525 (N_2525,In_1145,In_720);
nand U2526 (N_2526,In_1313,In_770);
xnor U2527 (N_2527,In_305,In_568);
or U2528 (N_2528,In_918,In_451);
or U2529 (N_2529,In_1460,In_1096);
or U2530 (N_2530,In_186,In_589);
and U2531 (N_2531,In_1438,In_1333);
or U2532 (N_2532,In_586,In_1445);
or U2533 (N_2533,In_724,In_797);
and U2534 (N_2534,In_1366,In_740);
xnor U2535 (N_2535,In_610,In_1088);
and U2536 (N_2536,In_463,In_376);
nor U2537 (N_2537,In_678,In_11);
nand U2538 (N_2538,In_528,In_1403);
nor U2539 (N_2539,In_199,In_168);
nand U2540 (N_2540,In_695,In_62);
xnor U2541 (N_2541,In_1110,In_1058);
xnor U2542 (N_2542,In_662,In_236);
xor U2543 (N_2543,In_260,In_937);
or U2544 (N_2544,In_1051,In_722);
or U2545 (N_2545,In_97,In_553);
nand U2546 (N_2546,In_585,In_1080);
nor U2547 (N_2547,In_93,In_159);
nand U2548 (N_2548,In_914,In_489);
and U2549 (N_2549,In_739,In_1444);
xor U2550 (N_2550,In_1306,In_433);
xnor U2551 (N_2551,In_1109,In_1103);
xor U2552 (N_2552,In_249,In_88);
nor U2553 (N_2553,In_366,In_450);
nor U2554 (N_2554,In_476,In_269);
nand U2555 (N_2555,In_1259,In_783);
or U2556 (N_2556,In_698,In_128);
or U2557 (N_2557,In_468,In_760);
or U2558 (N_2558,In_645,In_602);
nand U2559 (N_2559,In_993,In_1214);
xnor U2560 (N_2560,In_1253,In_336);
nand U2561 (N_2561,In_454,In_766);
nor U2562 (N_2562,In_185,In_292);
and U2563 (N_2563,In_374,In_355);
and U2564 (N_2564,In_904,In_814);
or U2565 (N_2565,In_570,In_179);
or U2566 (N_2566,In_901,In_787);
or U2567 (N_2567,In_17,In_1425);
nor U2568 (N_2568,In_1254,In_627);
and U2569 (N_2569,In_907,In_1159);
nand U2570 (N_2570,In_746,In_578);
xor U2571 (N_2571,In_1222,In_399);
and U2572 (N_2572,In_1259,In_544);
and U2573 (N_2573,In_1106,In_756);
xnor U2574 (N_2574,In_478,In_231);
xor U2575 (N_2575,In_499,In_1133);
and U2576 (N_2576,In_812,In_27);
nand U2577 (N_2577,In_1230,In_383);
nand U2578 (N_2578,In_949,In_1290);
nor U2579 (N_2579,In_909,In_1097);
nor U2580 (N_2580,In_1436,In_1130);
and U2581 (N_2581,In_155,In_1367);
and U2582 (N_2582,In_435,In_869);
xnor U2583 (N_2583,In_1247,In_658);
nand U2584 (N_2584,In_1442,In_641);
xnor U2585 (N_2585,In_258,In_733);
and U2586 (N_2586,In_553,In_877);
or U2587 (N_2587,In_80,In_1183);
nor U2588 (N_2588,In_1254,In_875);
xor U2589 (N_2589,In_633,In_47);
nand U2590 (N_2590,In_456,In_899);
and U2591 (N_2591,In_1063,In_1490);
and U2592 (N_2592,In_1481,In_468);
nor U2593 (N_2593,In_1388,In_1412);
nor U2594 (N_2594,In_123,In_1353);
nand U2595 (N_2595,In_1229,In_1457);
nand U2596 (N_2596,In_965,In_653);
and U2597 (N_2597,In_968,In_807);
and U2598 (N_2598,In_481,In_543);
nand U2599 (N_2599,In_434,In_32);
and U2600 (N_2600,In_1030,In_724);
nor U2601 (N_2601,In_986,In_296);
and U2602 (N_2602,In_1103,In_1228);
nor U2603 (N_2603,In_546,In_982);
and U2604 (N_2604,In_851,In_681);
or U2605 (N_2605,In_304,In_545);
xnor U2606 (N_2606,In_330,In_940);
or U2607 (N_2607,In_187,In_873);
xor U2608 (N_2608,In_591,In_547);
or U2609 (N_2609,In_763,In_758);
or U2610 (N_2610,In_1095,In_201);
nand U2611 (N_2611,In_617,In_505);
xor U2612 (N_2612,In_1131,In_1007);
xnor U2613 (N_2613,In_605,In_328);
nand U2614 (N_2614,In_1160,In_534);
or U2615 (N_2615,In_506,In_1065);
nor U2616 (N_2616,In_914,In_1265);
xnor U2617 (N_2617,In_1315,In_1304);
nand U2618 (N_2618,In_1461,In_1426);
nand U2619 (N_2619,In_1211,In_29);
or U2620 (N_2620,In_75,In_1421);
or U2621 (N_2621,In_667,In_59);
and U2622 (N_2622,In_466,In_1285);
and U2623 (N_2623,In_899,In_1244);
xnor U2624 (N_2624,In_1273,In_1282);
xnor U2625 (N_2625,In_1360,In_1117);
or U2626 (N_2626,In_579,In_8);
nor U2627 (N_2627,In_1327,In_951);
nor U2628 (N_2628,In_1411,In_673);
nor U2629 (N_2629,In_899,In_1340);
xor U2630 (N_2630,In_176,In_931);
nand U2631 (N_2631,In_486,In_1233);
and U2632 (N_2632,In_791,In_235);
and U2633 (N_2633,In_947,In_1047);
nand U2634 (N_2634,In_238,In_99);
or U2635 (N_2635,In_83,In_1);
or U2636 (N_2636,In_399,In_323);
nand U2637 (N_2637,In_1299,In_456);
or U2638 (N_2638,In_1462,In_1135);
and U2639 (N_2639,In_561,In_1148);
xnor U2640 (N_2640,In_325,In_1319);
nor U2641 (N_2641,In_1263,In_1038);
nand U2642 (N_2642,In_1220,In_150);
xor U2643 (N_2643,In_28,In_734);
nand U2644 (N_2644,In_559,In_1289);
or U2645 (N_2645,In_160,In_1160);
xor U2646 (N_2646,In_801,In_896);
and U2647 (N_2647,In_638,In_879);
and U2648 (N_2648,In_283,In_565);
or U2649 (N_2649,In_1073,In_113);
or U2650 (N_2650,In_1209,In_125);
xnor U2651 (N_2651,In_1300,In_1378);
and U2652 (N_2652,In_131,In_308);
or U2653 (N_2653,In_114,In_934);
nand U2654 (N_2654,In_228,In_1490);
and U2655 (N_2655,In_1396,In_1496);
or U2656 (N_2656,In_756,In_57);
nor U2657 (N_2657,In_1423,In_227);
xnor U2658 (N_2658,In_760,In_1205);
nand U2659 (N_2659,In_430,In_253);
nand U2660 (N_2660,In_1101,In_325);
and U2661 (N_2661,In_825,In_804);
or U2662 (N_2662,In_295,In_873);
nand U2663 (N_2663,In_788,In_672);
and U2664 (N_2664,In_915,In_1394);
xor U2665 (N_2665,In_1147,In_1432);
nor U2666 (N_2666,In_969,In_843);
nor U2667 (N_2667,In_67,In_1468);
nand U2668 (N_2668,In_337,In_1486);
nand U2669 (N_2669,In_60,In_309);
and U2670 (N_2670,In_492,In_1004);
and U2671 (N_2671,In_1027,In_333);
nand U2672 (N_2672,In_543,In_1388);
xor U2673 (N_2673,In_509,In_1193);
and U2674 (N_2674,In_1467,In_1159);
and U2675 (N_2675,In_729,In_1177);
nor U2676 (N_2676,In_284,In_291);
xor U2677 (N_2677,In_123,In_136);
nor U2678 (N_2678,In_475,In_1229);
or U2679 (N_2679,In_24,In_1176);
or U2680 (N_2680,In_62,In_951);
nor U2681 (N_2681,In_1064,In_1072);
or U2682 (N_2682,In_1039,In_151);
xnor U2683 (N_2683,In_1485,In_1079);
nor U2684 (N_2684,In_1106,In_966);
nand U2685 (N_2685,In_130,In_520);
xnor U2686 (N_2686,In_1102,In_627);
or U2687 (N_2687,In_714,In_712);
nor U2688 (N_2688,In_670,In_976);
nor U2689 (N_2689,In_287,In_161);
or U2690 (N_2690,In_865,In_667);
or U2691 (N_2691,In_612,In_1436);
or U2692 (N_2692,In_561,In_1204);
nor U2693 (N_2693,In_91,In_647);
and U2694 (N_2694,In_375,In_1008);
and U2695 (N_2695,In_1070,In_333);
nor U2696 (N_2696,In_280,In_104);
nand U2697 (N_2697,In_600,In_779);
or U2698 (N_2698,In_17,In_164);
nand U2699 (N_2699,In_1045,In_574);
nor U2700 (N_2700,In_213,In_1070);
nor U2701 (N_2701,In_1127,In_456);
nor U2702 (N_2702,In_1305,In_771);
and U2703 (N_2703,In_396,In_1444);
nand U2704 (N_2704,In_148,In_446);
or U2705 (N_2705,In_250,In_82);
nor U2706 (N_2706,In_1025,In_330);
or U2707 (N_2707,In_1394,In_728);
nand U2708 (N_2708,In_258,In_151);
nand U2709 (N_2709,In_177,In_1381);
nor U2710 (N_2710,In_24,In_50);
and U2711 (N_2711,In_1183,In_1465);
and U2712 (N_2712,In_1406,In_1196);
and U2713 (N_2713,In_446,In_155);
nand U2714 (N_2714,In_1405,In_48);
and U2715 (N_2715,In_903,In_1054);
xor U2716 (N_2716,In_1049,In_312);
nor U2717 (N_2717,In_80,In_1428);
xnor U2718 (N_2718,In_776,In_729);
nand U2719 (N_2719,In_435,In_609);
or U2720 (N_2720,In_500,In_869);
nor U2721 (N_2721,In_368,In_114);
nor U2722 (N_2722,In_130,In_646);
or U2723 (N_2723,In_1374,In_1028);
and U2724 (N_2724,In_410,In_1194);
xor U2725 (N_2725,In_1179,In_851);
and U2726 (N_2726,In_690,In_388);
nand U2727 (N_2727,In_1366,In_1418);
and U2728 (N_2728,In_215,In_281);
and U2729 (N_2729,In_1197,In_389);
nand U2730 (N_2730,In_198,In_1246);
and U2731 (N_2731,In_549,In_1041);
nor U2732 (N_2732,In_1146,In_152);
nor U2733 (N_2733,In_825,In_738);
or U2734 (N_2734,In_1005,In_392);
nor U2735 (N_2735,In_711,In_487);
xnor U2736 (N_2736,In_890,In_781);
nand U2737 (N_2737,In_29,In_444);
nand U2738 (N_2738,In_1058,In_1341);
nor U2739 (N_2739,In_780,In_953);
or U2740 (N_2740,In_970,In_1334);
or U2741 (N_2741,In_1218,In_605);
xor U2742 (N_2742,In_709,In_352);
or U2743 (N_2743,In_1473,In_287);
nand U2744 (N_2744,In_1126,In_664);
xor U2745 (N_2745,In_1381,In_1129);
xnor U2746 (N_2746,In_1000,In_881);
xnor U2747 (N_2747,In_542,In_1270);
nand U2748 (N_2748,In_707,In_14);
nor U2749 (N_2749,In_894,In_949);
nor U2750 (N_2750,In_514,In_227);
and U2751 (N_2751,In_456,In_1466);
xor U2752 (N_2752,In_1391,In_379);
xor U2753 (N_2753,In_770,In_490);
nor U2754 (N_2754,In_318,In_1209);
or U2755 (N_2755,In_782,In_1129);
xor U2756 (N_2756,In_1221,In_1236);
nor U2757 (N_2757,In_365,In_667);
nor U2758 (N_2758,In_849,In_307);
or U2759 (N_2759,In_1206,In_531);
nand U2760 (N_2760,In_545,In_1248);
xnor U2761 (N_2761,In_1497,In_1111);
or U2762 (N_2762,In_87,In_66);
nor U2763 (N_2763,In_277,In_243);
nand U2764 (N_2764,In_360,In_264);
nand U2765 (N_2765,In_494,In_1137);
nor U2766 (N_2766,In_13,In_1013);
nand U2767 (N_2767,In_143,In_216);
or U2768 (N_2768,In_1066,In_1373);
and U2769 (N_2769,In_1484,In_1493);
and U2770 (N_2770,In_628,In_247);
nor U2771 (N_2771,In_1279,In_86);
nor U2772 (N_2772,In_1128,In_1367);
and U2773 (N_2773,In_526,In_582);
nand U2774 (N_2774,In_328,In_1224);
or U2775 (N_2775,In_731,In_971);
nand U2776 (N_2776,In_1330,In_740);
and U2777 (N_2777,In_593,In_1344);
or U2778 (N_2778,In_886,In_1264);
nor U2779 (N_2779,In_1082,In_701);
or U2780 (N_2780,In_924,In_559);
and U2781 (N_2781,In_1323,In_834);
nand U2782 (N_2782,In_94,In_227);
nor U2783 (N_2783,In_507,In_43);
or U2784 (N_2784,In_276,In_640);
nor U2785 (N_2785,In_152,In_1473);
or U2786 (N_2786,In_1011,In_1457);
nor U2787 (N_2787,In_1316,In_1231);
xor U2788 (N_2788,In_560,In_1477);
or U2789 (N_2789,In_887,In_1369);
nand U2790 (N_2790,In_1069,In_831);
nand U2791 (N_2791,In_269,In_701);
and U2792 (N_2792,In_970,In_1306);
and U2793 (N_2793,In_254,In_919);
or U2794 (N_2794,In_1237,In_1355);
or U2795 (N_2795,In_1005,In_594);
nand U2796 (N_2796,In_1478,In_1169);
nand U2797 (N_2797,In_418,In_1193);
nand U2798 (N_2798,In_256,In_112);
nand U2799 (N_2799,In_884,In_813);
xnor U2800 (N_2800,In_13,In_1280);
or U2801 (N_2801,In_384,In_1219);
xnor U2802 (N_2802,In_223,In_844);
nand U2803 (N_2803,In_260,In_553);
and U2804 (N_2804,In_77,In_998);
xnor U2805 (N_2805,In_925,In_139);
or U2806 (N_2806,In_674,In_637);
xor U2807 (N_2807,In_966,In_591);
nand U2808 (N_2808,In_408,In_853);
or U2809 (N_2809,In_1436,In_1496);
xnor U2810 (N_2810,In_276,In_51);
nor U2811 (N_2811,In_1359,In_36);
xnor U2812 (N_2812,In_860,In_1081);
and U2813 (N_2813,In_366,In_83);
xor U2814 (N_2814,In_1186,In_1038);
nor U2815 (N_2815,In_1188,In_1002);
nor U2816 (N_2816,In_270,In_183);
nand U2817 (N_2817,In_319,In_1171);
and U2818 (N_2818,In_1024,In_112);
and U2819 (N_2819,In_695,In_508);
or U2820 (N_2820,In_103,In_1103);
xnor U2821 (N_2821,In_220,In_126);
xnor U2822 (N_2822,In_1179,In_551);
and U2823 (N_2823,In_1187,In_392);
and U2824 (N_2824,In_156,In_669);
nand U2825 (N_2825,In_169,In_919);
xor U2826 (N_2826,In_107,In_585);
nor U2827 (N_2827,In_748,In_567);
nor U2828 (N_2828,In_1006,In_312);
or U2829 (N_2829,In_1039,In_1441);
xnor U2830 (N_2830,In_167,In_412);
or U2831 (N_2831,In_1314,In_1391);
and U2832 (N_2832,In_1261,In_22);
nand U2833 (N_2833,In_248,In_1245);
and U2834 (N_2834,In_800,In_572);
nor U2835 (N_2835,In_648,In_108);
xor U2836 (N_2836,In_849,In_589);
and U2837 (N_2837,In_761,In_897);
and U2838 (N_2838,In_746,In_360);
nand U2839 (N_2839,In_171,In_667);
nor U2840 (N_2840,In_501,In_248);
xnor U2841 (N_2841,In_550,In_287);
and U2842 (N_2842,In_183,In_1428);
nand U2843 (N_2843,In_802,In_982);
nor U2844 (N_2844,In_1134,In_503);
nand U2845 (N_2845,In_1007,In_118);
xnor U2846 (N_2846,In_596,In_634);
nand U2847 (N_2847,In_1059,In_1243);
nand U2848 (N_2848,In_1321,In_130);
or U2849 (N_2849,In_610,In_254);
xor U2850 (N_2850,In_326,In_1264);
nor U2851 (N_2851,In_955,In_31);
and U2852 (N_2852,In_785,In_498);
nand U2853 (N_2853,In_167,In_791);
xor U2854 (N_2854,In_71,In_1151);
or U2855 (N_2855,In_1309,In_596);
nand U2856 (N_2856,In_1393,In_415);
and U2857 (N_2857,In_385,In_527);
and U2858 (N_2858,In_1215,In_1400);
or U2859 (N_2859,In_456,In_247);
xnor U2860 (N_2860,In_1157,In_214);
and U2861 (N_2861,In_963,In_472);
xor U2862 (N_2862,In_815,In_520);
nor U2863 (N_2863,In_309,In_307);
nand U2864 (N_2864,In_1116,In_133);
xor U2865 (N_2865,In_85,In_1444);
and U2866 (N_2866,In_1007,In_1104);
or U2867 (N_2867,In_1492,In_38);
and U2868 (N_2868,In_209,In_1010);
or U2869 (N_2869,In_277,In_806);
nor U2870 (N_2870,In_1183,In_474);
nand U2871 (N_2871,In_216,In_202);
and U2872 (N_2872,In_758,In_340);
nor U2873 (N_2873,In_233,In_306);
or U2874 (N_2874,In_393,In_411);
xor U2875 (N_2875,In_592,In_1277);
nor U2876 (N_2876,In_1471,In_298);
and U2877 (N_2877,In_235,In_312);
xor U2878 (N_2878,In_453,In_573);
or U2879 (N_2879,In_684,In_833);
or U2880 (N_2880,In_1199,In_790);
or U2881 (N_2881,In_748,In_1472);
nand U2882 (N_2882,In_630,In_1014);
nand U2883 (N_2883,In_1373,In_16);
xor U2884 (N_2884,In_1217,In_651);
and U2885 (N_2885,In_1271,In_930);
and U2886 (N_2886,In_704,In_1420);
xnor U2887 (N_2887,In_844,In_1061);
xor U2888 (N_2888,In_840,In_1127);
xor U2889 (N_2889,In_1150,In_1166);
and U2890 (N_2890,In_896,In_622);
or U2891 (N_2891,In_1480,In_928);
xnor U2892 (N_2892,In_1051,In_727);
nand U2893 (N_2893,In_411,In_310);
xor U2894 (N_2894,In_680,In_1079);
and U2895 (N_2895,In_382,In_1048);
nand U2896 (N_2896,In_241,In_945);
nor U2897 (N_2897,In_453,In_627);
and U2898 (N_2898,In_1457,In_520);
xor U2899 (N_2899,In_387,In_823);
and U2900 (N_2900,In_499,In_127);
xnor U2901 (N_2901,In_568,In_831);
nand U2902 (N_2902,In_1306,In_1307);
nand U2903 (N_2903,In_306,In_343);
xnor U2904 (N_2904,In_1355,In_1037);
nand U2905 (N_2905,In_1091,In_1114);
and U2906 (N_2906,In_599,In_1223);
xnor U2907 (N_2907,In_1476,In_123);
xnor U2908 (N_2908,In_299,In_253);
nor U2909 (N_2909,In_375,In_22);
xor U2910 (N_2910,In_826,In_11);
xor U2911 (N_2911,In_1431,In_1391);
nor U2912 (N_2912,In_907,In_1408);
and U2913 (N_2913,In_761,In_567);
or U2914 (N_2914,In_1014,In_297);
xor U2915 (N_2915,In_474,In_1374);
xnor U2916 (N_2916,In_843,In_607);
or U2917 (N_2917,In_999,In_305);
nor U2918 (N_2918,In_409,In_1289);
nand U2919 (N_2919,In_539,In_120);
nand U2920 (N_2920,In_408,In_1093);
nor U2921 (N_2921,In_868,In_1164);
nor U2922 (N_2922,In_1236,In_414);
or U2923 (N_2923,In_1050,In_80);
nand U2924 (N_2924,In_1431,In_1436);
or U2925 (N_2925,In_443,In_379);
xor U2926 (N_2926,In_1257,In_788);
nor U2927 (N_2927,In_627,In_1378);
xnor U2928 (N_2928,In_1412,In_1422);
nand U2929 (N_2929,In_156,In_1391);
or U2930 (N_2930,In_569,In_230);
xor U2931 (N_2931,In_76,In_205);
or U2932 (N_2932,In_1419,In_1417);
nand U2933 (N_2933,In_1403,In_525);
nand U2934 (N_2934,In_1396,In_1286);
or U2935 (N_2935,In_812,In_1186);
xor U2936 (N_2936,In_460,In_1095);
nand U2937 (N_2937,In_1000,In_1467);
or U2938 (N_2938,In_170,In_1058);
nand U2939 (N_2939,In_255,In_1278);
and U2940 (N_2940,In_219,In_1164);
nor U2941 (N_2941,In_896,In_666);
xnor U2942 (N_2942,In_748,In_1140);
nand U2943 (N_2943,In_1154,In_912);
nand U2944 (N_2944,In_37,In_189);
xor U2945 (N_2945,In_1023,In_543);
or U2946 (N_2946,In_575,In_100);
xnor U2947 (N_2947,In_456,In_285);
and U2948 (N_2948,In_1395,In_198);
nand U2949 (N_2949,In_1037,In_226);
or U2950 (N_2950,In_583,In_772);
nor U2951 (N_2951,In_474,In_174);
xnor U2952 (N_2952,In_426,In_1116);
nand U2953 (N_2953,In_1293,In_28);
or U2954 (N_2954,In_1127,In_1340);
and U2955 (N_2955,In_120,In_9);
nand U2956 (N_2956,In_1352,In_1371);
xor U2957 (N_2957,In_301,In_454);
nand U2958 (N_2958,In_740,In_640);
and U2959 (N_2959,In_979,In_692);
nor U2960 (N_2960,In_52,In_1270);
xnor U2961 (N_2961,In_496,In_2);
nor U2962 (N_2962,In_18,In_1083);
or U2963 (N_2963,In_778,In_146);
nand U2964 (N_2964,In_1385,In_576);
and U2965 (N_2965,In_1480,In_228);
and U2966 (N_2966,In_450,In_431);
xor U2967 (N_2967,In_486,In_1115);
and U2968 (N_2968,In_1080,In_536);
or U2969 (N_2969,In_86,In_1067);
nor U2970 (N_2970,In_1053,In_954);
nor U2971 (N_2971,In_734,In_873);
and U2972 (N_2972,In_522,In_1238);
nor U2973 (N_2973,In_1271,In_886);
and U2974 (N_2974,In_470,In_547);
nand U2975 (N_2975,In_1486,In_555);
and U2976 (N_2976,In_1443,In_1417);
or U2977 (N_2977,In_861,In_592);
nor U2978 (N_2978,In_855,In_32);
and U2979 (N_2979,In_871,In_562);
or U2980 (N_2980,In_1264,In_702);
or U2981 (N_2981,In_1355,In_1084);
xnor U2982 (N_2982,In_1488,In_88);
and U2983 (N_2983,In_1115,In_1272);
nor U2984 (N_2984,In_84,In_225);
xnor U2985 (N_2985,In_1295,In_246);
nor U2986 (N_2986,In_516,In_217);
nand U2987 (N_2987,In_226,In_683);
nand U2988 (N_2988,In_301,In_1280);
or U2989 (N_2989,In_1184,In_1296);
or U2990 (N_2990,In_307,In_972);
or U2991 (N_2991,In_186,In_1236);
xnor U2992 (N_2992,In_716,In_700);
nor U2993 (N_2993,In_1385,In_396);
nor U2994 (N_2994,In_876,In_1190);
xnor U2995 (N_2995,In_1466,In_1216);
xor U2996 (N_2996,In_18,In_791);
xnor U2997 (N_2997,In_1420,In_987);
xor U2998 (N_2998,In_1452,In_271);
nand U2999 (N_2999,In_554,In_982);
nand U3000 (N_3000,N_2512,N_1490);
nand U3001 (N_3001,N_738,N_477);
nor U3002 (N_3002,N_1639,N_2339);
nand U3003 (N_3003,N_2154,N_1778);
nor U3004 (N_3004,N_692,N_906);
or U3005 (N_3005,N_1954,N_145);
or U3006 (N_3006,N_1578,N_374);
or U3007 (N_3007,N_1846,N_383);
xor U3008 (N_3008,N_45,N_1467);
nor U3009 (N_3009,N_1617,N_1154);
nor U3010 (N_3010,N_798,N_1050);
nand U3011 (N_3011,N_1461,N_19);
or U3012 (N_3012,N_861,N_1269);
or U3013 (N_3013,N_1263,N_2521);
or U3014 (N_3014,N_1933,N_1260);
or U3015 (N_3015,N_155,N_1322);
nor U3016 (N_3016,N_1828,N_923);
and U3017 (N_3017,N_2249,N_1953);
or U3018 (N_3018,N_1730,N_766);
nand U3019 (N_3019,N_874,N_1091);
nor U3020 (N_3020,N_2586,N_110);
or U3021 (N_3021,N_2106,N_2258);
nor U3022 (N_3022,N_1297,N_1818);
nand U3023 (N_3023,N_2053,N_2368);
xor U3024 (N_3024,N_2729,N_39);
xnor U3025 (N_3025,N_2322,N_1536);
nand U3026 (N_3026,N_1149,N_2202);
and U3027 (N_3027,N_1148,N_70);
nor U3028 (N_3028,N_870,N_35);
nand U3029 (N_3029,N_2359,N_224);
xnor U3030 (N_3030,N_2735,N_2244);
xor U3031 (N_3031,N_2019,N_1298);
nand U3032 (N_3032,N_2127,N_1176);
nor U3033 (N_3033,N_1039,N_77);
nor U3034 (N_3034,N_799,N_206);
and U3035 (N_3035,N_592,N_1463);
and U3036 (N_3036,N_220,N_2495);
nor U3037 (N_3037,N_1078,N_2924);
xor U3038 (N_3038,N_1669,N_598);
xor U3039 (N_3039,N_287,N_1040);
xor U3040 (N_3040,N_1371,N_1546);
nand U3041 (N_3041,N_1679,N_415);
and U3042 (N_3042,N_2403,N_118);
and U3043 (N_3043,N_2045,N_2354);
nor U3044 (N_3044,N_191,N_1480);
and U3045 (N_3045,N_1034,N_2835);
and U3046 (N_3046,N_2808,N_770);
nand U3047 (N_3047,N_2948,N_673);
nor U3048 (N_3048,N_697,N_108);
nor U3049 (N_3049,N_227,N_1093);
xor U3050 (N_3050,N_1376,N_2736);
nand U3051 (N_3051,N_714,N_1698);
nor U3052 (N_3052,N_307,N_2073);
or U3053 (N_3053,N_2259,N_2724);
xor U3054 (N_3054,N_777,N_258);
and U3055 (N_3055,N_638,N_1887);
xor U3056 (N_3056,N_90,N_195);
or U3057 (N_3057,N_61,N_1518);
xor U3058 (N_3058,N_1006,N_194);
or U3059 (N_3059,N_2913,N_2270);
nand U3060 (N_3060,N_857,N_2183);
nand U3061 (N_3061,N_1700,N_214);
nand U3062 (N_3062,N_2556,N_959);
nand U3063 (N_3063,N_2875,N_541);
and U3064 (N_3064,N_2666,N_1080);
xnor U3065 (N_3065,N_2885,N_103);
xor U3066 (N_3066,N_1513,N_1549);
nand U3067 (N_3067,N_2429,N_1843);
nand U3068 (N_3068,N_866,N_2993);
or U3069 (N_3069,N_208,N_555);
and U3070 (N_3070,N_1787,N_1280);
xor U3071 (N_3071,N_705,N_1731);
nand U3072 (N_3072,N_2380,N_719);
xor U3073 (N_3073,N_2461,N_1147);
nand U3074 (N_3074,N_325,N_2109);
nor U3075 (N_3075,N_1898,N_2225);
and U3076 (N_3076,N_1950,N_1916);
nor U3077 (N_3077,N_2230,N_1164);
nand U3078 (N_3078,N_776,N_449);
or U3079 (N_3079,N_1305,N_512);
xor U3080 (N_3080,N_1524,N_221);
xor U3081 (N_3081,N_382,N_936);
nand U3082 (N_3082,N_368,N_335);
or U3083 (N_3083,N_838,N_1345);
nor U3084 (N_3084,N_2162,N_2925);
or U3085 (N_3085,N_628,N_1509);
xnor U3086 (N_3086,N_2803,N_2854);
and U3087 (N_3087,N_899,N_920);
nor U3088 (N_3088,N_877,N_2123);
xor U3089 (N_3089,N_2800,N_2907);
xnor U3090 (N_3090,N_599,N_16);
nor U3091 (N_3091,N_1014,N_1876);
nand U3092 (N_3092,N_97,N_1842);
nor U3093 (N_3093,N_1388,N_1226);
nand U3094 (N_3094,N_2003,N_872);
nand U3095 (N_3095,N_497,N_167);
nand U3096 (N_3096,N_1794,N_1047);
xnor U3097 (N_3097,N_925,N_2166);
nor U3098 (N_3098,N_728,N_1563);
or U3099 (N_3099,N_402,N_1606);
nor U3100 (N_3100,N_2767,N_800);
nor U3101 (N_3101,N_352,N_1009);
nand U3102 (N_3102,N_2066,N_2099);
xnor U3103 (N_3103,N_20,N_2028);
or U3104 (N_3104,N_759,N_192);
or U3105 (N_3105,N_2132,N_93);
and U3106 (N_3106,N_1429,N_2761);
xor U3107 (N_3107,N_422,N_687);
nor U3108 (N_3108,N_2231,N_1835);
and U3109 (N_3109,N_2366,N_2916);
xnor U3110 (N_3110,N_515,N_2604);
nor U3111 (N_3111,N_33,N_1740);
nand U3112 (N_3112,N_819,N_2638);
nor U3113 (N_3113,N_1935,N_2242);
and U3114 (N_3114,N_2320,N_2237);
nand U3115 (N_3115,N_124,N_988);
xnor U3116 (N_3116,N_1455,N_2509);
xor U3117 (N_3117,N_2549,N_1663);
and U3118 (N_3118,N_904,N_1443);
and U3119 (N_3119,N_150,N_1003);
nand U3120 (N_3120,N_2575,N_583);
nand U3121 (N_3121,N_359,N_672);
xor U3122 (N_3122,N_2864,N_606);
nand U3123 (N_3123,N_1087,N_1348);
or U3124 (N_3124,N_740,N_387);
or U3125 (N_3125,N_722,N_2603);
xnor U3126 (N_3126,N_1688,N_2542);
xor U3127 (N_3127,N_101,N_212);
nand U3128 (N_3128,N_2213,N_657);
and U3129 (N_3129,N_865,N_2457);
xor U3130 (N_3130,N_641,N_1032);
nor U3131 (N_3131,N_755,N_827);
nand U3132 (N_3132,N_2409,N_466);
and U3133 (N_3133,N_426,N_2896);
and U3134 (N_3134,N_1210,N_475);
nand U3135 (N_3135,N_2086,N_2677);
nand U3136 (N_3136,N_2517,N_297);
xnor U3137 (N_3137,N_1988,N_1083);
and U3138 (N_3138,N_1121,N_1572);
or U3139 (N_3139,N_1676,N_1433);
nor U3140 (N_3140,N_2945,N_2006);
nand U3141 (N_3141,N_1364,N_806);
and U3142 (N_3142,N_1718,N_1444);
and U3143 (N_3143,N_1355,N_1253);
or U3144 (N_3144,N_1508,N_1943);
or U3145 (N_3145,N_586,N_2500);
nand U3146 (N_3146,N_1105,N_1271);
nor U3147 (N_3147,N_2927,N_1293);
or U3148 (N_3148,N_468,N_3);
nor U3149 (N_3149,N_363,N_2937);
nor U3150 (N_3150,N_1715,N_1761);
or U3151 (N_3151,N_1754,N_1379);
xor U3152 (N_3152,N_1870,N_1707);
nand U3153 (N_3153,N_286,N_660);
and U3154 (N_3154,N_1519,N_198);
nand U3155 (N_3155,N_2141,N_2034);
or U3156 (N_3156,N_811,N_1108);
or U3157 (N_3157,N_2817,N_1431);
xor U3158 (N_3158,N_2718,N_743);
and U3159 (N_3159,N_1928,N_1523);
xor U3160 (N_3160,N_2007,N_663);
nor U3161 (N_3161,N_2962,N_447);
xnor U3162 (N_3162,N_2210,N_903);
nor U3163 (N_3163,N_1960,N_2918);
or U3164 (N_3164,N_1276,N_2867);
nor U3165 (N_3165,N_342,N_260);
and U3166 (N_3166,N_1425,N_1408);
or U3167 (N_3167,N_2682,N_2195);
xnor U3168 (N_3168,N_1879,N_2250);
xor U3169 (N_3169,N_2621,N_726);
nor U3170 (N_3170,N_652,N_364);
xor U3171 (N_3171,N_1247,N_532);
xnor U3172 (N_3172,N_480,N_381);
and U3173 (N_3173,N_1945,N_825);
xor U3174 (N_3174,N_2633,N_979);
or U3175 (N_3175,N_2506,N_1535);
nand U3176 (N_3176,N_546,N_876);
or U3177 (N_3177,N_1330,N_1144);
nor U3178 (N_3178,N_2528,N_1011);
or U3179 (N_3179,N_2274,N_1368);
and U3180 (N_3180,N_971,N_614);
nor U3181 (N_3181,N_2544,N_2869);
nand U3182 (N_3182,N_1178,N_2358);
and U3183 (N_3183,N_1206,N_1805);
nand U3184 (N_3184,N_233,N_1094);
or U3185 (N_3185,N_2441,N_1837);
nand U3186 (N_3186,N_2773,N_2292);
and U3187 (N_3187,N_2135,N_1495);
xor U3188 (N_3188,N_1106,N_2827);
or U3189 (N_3189,N_1932,N_1325);
or U3190 (N_3190,N_322,N_1815);
xor U3191 (N_3191,N_2858,N_2049);
nor U3192 (N_3192,N_2806,N_2485);
or U3193 (N_3193,N_2752,N_618);
nand U3194 (N_3194,N_593,N_1249);
nor U3195 (N_3195,N_1030,N_2238);
nor U3196 (N_3196,N_1044,N_626);
nand U3197 (N_3197,N_2969,N_1346);
or U3198 (N_3198,N_1162,N_905);
nor U3199 (N_3199,N_289,N_397);
xnor U3200 (N_3200,N_313,N_622);
or U3201 (N_3201,N_303,N_684);
xor U3202 (N_3202,N_717,N_2727);
nor U3203 (N_3203,N_55,N_1079);
nand U3204 (N_3204,N_2093,N_1602);
xor U3205 (N_3205,N_2856,N_434);
and U3206 (N_3206,N_2092,N_711);
nor U3207 (N_3207,N_2702,N_2932);
nand U3208 (N_3208,N_419,N_1415);
xor U3209 (N_3209,N_1258,N_758);
or U3210 (N_3210,N_281,N_339);
nor U3211 (N_3211,N_247,N_1151);
or U3212 (N_3212,N_938,N_2828);
xnor U3213 (N_3213,N_2012,N_1021);
and U3214 (N_3214,N_1802,N_1385);
and U3215 (N_3215,N_1442,N_1278);
nor U3216 (N_3216,N_1333,N_1387);
nand U3217 (N_3217,N_1634,N_2190);
and U3218 (N_3218,N_2963,N_2487);
nor U3219 (N_3219,N_1062,N_829);
nand U3220 (N_3220,N_709,N_1274);
xor U3221 (N_3221,N_2928,N_1741);
xnor U3222 (N_3222,N_2017,N_2988);
and U3223 (N_3223,N_2921,N_276);
and U3224 (N_3224,N_1059,N_2656);
xnor U3225 (N_3225,N_2934,N_2079);
nor U3226 (N_3226,N_954,N_2389);
and U3227 (N_3227,N_2795,N_520);
and U3228 (N_3228,N_601,N_1375);
and U3229 (N_3229,N_1643,N_1214);
xor U3230 (N_3230,N_2583,N_2745);
or U3231 (N_3231,N_251,N_2164);
nor U3232 (N_3232,N_430,N_196);
nor U3233 (N_3233,N_2505,N_2033);
nor U3234 (N_3234,N_265,N_2236);
and U3235 (N_3235,N_1252,N_311);
nor U3236 (N_3236,N_2031,N_1315);
nand U3237 (N_3237,N_1008,N_1589);
xor U3238 (N_3238,N_2206,N_892);
and U3239 (N_3239,N_1073,N_981);
or U3240 (N_3240,N_886,N_908);
nand U3241 (N_3241,N_160,N_1165);
xnor U3242 (N_3242,N_230,N_737);
nand U3243 (N_3243,N_804,N_1581);
and U3244 (N_3244,N_1358,N_1931);
xor U3245 (N_3245,N_72,N_1290);
nand U3246 (N_3246,N_186,N_760);
or U3247 (N_3247,N_1028,N_69);
and U3248 (N_3248,N_1714,N_189);
or U3249 (N_3249,N_1808,N_1940);
nand U3250 (N_3250,N_1584,N_1613);
nand U3251 (N_3251,N_944,N_772);
nor U3252 (N_3252,N_26,N_2104);
nor U3253 (N_3253,N_1789,N_2900);
or U3254 (N_3254,N_2475,N_1357);
nand U3255 (N_3255,N_2965,N_510);
xnor U3256 (N_3256,N_365,N_79);
nor U3257 (N_3257,N_2943,N_837);
and U3258 (N_3258,N_200,N_2791);
or U3259 (N_3259,N_1347,N_389);
xor U3260 (N_3260,N_1129,N_1488);
nor U3261 (N_3261,N_1025,N_1246);
nor U3262 (N_3262,N_2632,N_587);
nor U3263 (N_3263,N_1880,N_2440);
and U3264 (N_3264,N_2699,N_2116);
xnor U3265 (N_3265,N_2272,N_831);
or U3266 (N_3266,N_1853,N_361);
nand U3267 (N_3267,N_1962,N_2645);
nor U3268 (N_3268,N_2118,N_782);
nand U3269 (N_3269,N_2406,N_2443);
or U3270 (N_3270,N_2836,N_2563);
and U3271 (N_3271,N_1575,N_620);
xnor U3272 (N_3272,N_2911,N_2484);
or U3273 (N_3273,N_2121,N_1155);
or U3274 (N_3274,N_282,N_348);
xor U3275 (N_3275,N_552,N_2862);
nand U3276 (N_3276,N_1955,N_1288);
xnor U3277 (N_3277,N_2744,N_527);
and U3278 (N_3278,N_1307,N_1185);
xnor U3279 (N_3279,N_2321,N_1595);
nor U3280 (N_3280,N_949,N_1324);
nor U3281 (N_3281,N_2407,N_459);
and U3282 (N_3282,N_1235,N_2514);
and U3283 (N_3283,N_1990,N_1830);
or U3284 (N_3284,N_1102,N_2878);
and U3285 (N_3285,N_1396,N_600);
nand U3286 (N_3286,N_1560,N_2762);
or U3287 (N_3287,N_156,N_1746);
nor U3288 (N_3288,N_2282,N_1294);
or U3289 (N_3289,N_159,N_1506);
or U3290 (N_3290,N_830,N_2103);
nor U3291 (N_3291,N_2305,N_2284);
xnor U3292 (N_3292,N_1958,N_788);
nand U3293 (N_3293,N_1066,N_2383);
nand U3294 (N_3294,N_2470,N_2749);
nand U3295 (N_3295,N_1732,N_203);
nor U3296 (N_3296,N_99,N_438);
xor U3297 (N_3297,N_636,N_958);
nor U3298 (N_3298,N_508,N_2035);
and U3299 (N_3299,N_1555,N_1769);
nor U3300 (N_3300,N_1365,N_2560);
or U3301 (N_3301,N_184,N_1114);
and U3302 (N_3302,N_1825,N_2071);
nand U3303 (N_3303,N_37,N_2765);
nand U3304 (N_3304,N_2941,N_2629);
nor U3305 (N_3305,N_1614,N_1196);
xnor U3306 (N_3306,N_655,N_1194);
xor U3307 (N_3307,N_1976,N_2208);
xor U3308 (N_3308,N_2480,N_581);
and U3309 (N_3309,N_2929,N_589);
or U3310 (N_3310,N_972,N_683);
nor U3311 (N_3311,N_1735,N_1781);
nor U3312 (N_3312,N_2692,N_1734);
nand U3313 (N_3313,N_1076,N_471);
nand U3314 (N_3314,N_2551,N_1085);
nor U3315 (N_3315,N_499,N_967);
and U3316 (N_3316,N_314,N_1845);
and U3317 (N_3317,N_249,N_2748);
nor U3318 (N_3318,N_2091,N_1666);
or U3319 (N_3319,N_1267,N_573);
or U3320 (N_3320,N_1042,N_2655);
or U3321 (N_3321,N_795,N_1948);
or U3322 (N_3322,N_2136,N_2920);
nor U3323 (N_3323,N_46,N_2573);
nand U3324 (N_3324,N_2823,N_1435);
and U3325 (N_3325,N_775,N_2311);
and U3326 (N_3326,N_1860,N_1636);
xor U3327 (N_3327,N_1137,N_22);
nand U3328 (N_3328,N_994,N_2165);
and U3329 (N_3329,N_2599,N_1970);
and U3330 (N_3330,N_2014,N_130);
nor U3331 (N_3331,N_403,N_1166);
xnor U3332 (N_3332,N_2138,N_1122);
xor U3333 (N_3333,N_1604,N_1938);
nand U3334 (N_3334,N_1097,N_65);
xnor U3335 (N_3335,N_1022,N_1213);
nor U3336 (N_3336,N_1233,N_823);
nand U3337 (N_3337,N_469,N_2652);
or U3338 (N_3338,N_1138,N_531);
or U3339 (N_3339,N_2764,N_2851);
and U3340 (N_3340,N_539,N_960);
nor U3341 (N_3341,N_2490,N_1370);
xor U3342 (N_3342,N_1107,N_183);
and U3343 (N_3343,N_2353,N_2535);
nor U3344 (N_3344,N_2508,N_619);
nor U3345 (N_3345,N_631,N_2126);
or U3346 (N_3346,N_2788,N_602);
xnor U3347 (N_3347,N_1564,N_1986);
and U3348 (N_3348,N_2408,N_351);
xnor U3349 (N_3349,N_2115,N_1055);
xor U3350 (N_3350,N_1559,N_437);
nand U3351 (N_3351,N_2482,N_1646);
xor U3352 (N_3352,N_2690,N_2847);
and U3353 (N_3353,N_373,N_1470);
and U3354 (N_3354,N_1018,N_1332);
nand U3355 (N_3355,N_178,N_1542);
or U3356 (N_3356,N_1302,N_100);
and U3357 (N_3357,N_1631,N_1979);
xnor U3358 (N_3358,N_654,N_1456);
or U3359 (N_3359,N_2679,N_1775);
nand U3360 (N_3360,N_318,N_1343);
nand U3361 (N_3361,N_835,N_2531);
nand U3362 (N_3362,N_1354,N_1497);
or U3363 (N_3363,N_417,N_179);
nand U3364 (N_3364,N_2192,N_143);
xnor U3365 (N_3365,N_237,N_98);
or U3366 (N_3366,N_2108,N_2248);
and U3367 (N_3367,N_2774,N_1693);
or U3368 (N_3368,N_1321,N_2515);
nand U3369 (N_3369,N_1854,N_2285);
xor U3370 (N_3370,N_2820,N_794);
nand U3371 (N_3371,N_817,N_2152);
nand U3372 (N_3372,N_689,N_771);
or U3373 (N_3373,N_2193,N_1476);
xnor U3374 (N_3374,N_2469,N_2615);
xor U3375 (N_3375,N_302,N_1483);
and U3376 (N_3376,N_1386,N_170);
or U3377 (N_3377,N_1472,N_2356);
nor U3378 (N_3378,N_343,N_1531);
and U3379 (N_3379,N_2362,N_2898);
xnor U3380 (N_3380,N_1098,N_885);
xnor U3381 (N_3381,N_2568,N_2614);
xnor U3382 (N_3382,N_1309,N_1996);
xor U3383 (N_3383,N_1677,N_1193);
or U3384 (N_3384,N_2704,N_1172);
or U3385 (N_3385,N_142,N_1793);
and U3386 (N_3386,N_1684,N_1974);
nand U3387 (N_3387,N_1096,N_561);
and U3388 (N_3388,N_125,N_91);
xor U3389 (N_3389,N_2239,N_316);
and U3390 (N_3390,N_340,N_1699);
xor U3391 (N_3391,N_1720,N_677);
and U3392 (N_3392,N_85,N_239);
xnor U3393 (N_3393,N_2426,N_1556);
nor U3394 (N_3394,N_752,N_907);
or U3395 (N_3395,N_2959,N_1882);
nor U3396 (N_3396,N_2961,N_919);
nand U3397 (N_3397,N_2060,N_1132);
and U3398 (N_3398,N_801,N_2566);
nor U3399 (N_3399,N_2792,N_2693);
or U3400 (N_3400,N_439,N_2063);
or U3401 (N_3401,N_1587,N_2785);
and U3402 (N_3402,N_2289,N_1349);
or U3403 (N_3403,N_2223,N_1770);
and U3404 (N_3404,N_973,N_1339);
and U3405 (N_3405,N_2290,N_245);
and U3406 (N_3406,N_2578,N_2177);
nand U3407 (N_3407,N_1250,N_346);
nand U3408 (N_3408,N_2589,N_168);
nand U3409 (N_3409,N_1123,N_1141);
nor U3410 (N_3410,N_24,N_2709);
nor U3411 (N_3411,N_1806,N_1822);
xnor U3412 (N_3412,N_1736,N_1458);
nand U3413 (N_3413,N_112,N_2228);
and U3414 (N_3414,N_2799,N_2314);
or U3415 (N_3415,N_1627,N_691);
nor U3416 (N_3416,N_2131,N_544);
or U3417 (N_3417,N_2734,N_1514);
and U3418 (N_3418,N_2390,N_21);
or U3419 (N_3419,N_918,N_2468);
nand U3420 (N_3420,N_2020,N_651);
xnor U3421 (N_3421,N_1146,N_1817);
or U3422 (N_3422,N_27,N_187);
nand U3423 (N_3423,N_2554,N_2462);
xor U3424 (N_3424,N_241,N_1539);
nor U3425 (N_3425,N_190,N_2149);
nor U3426 (N_3426,N_1160,N_2985);
nor U3427 (N_3427,N_2,N_2931);
or U3428 (N_3428,N_1993,N_94);
xnor U3429 (N_3429,N_152,N_1527);
nor U3430 (N_3430,N_379,N_2215);
and U3431 (N_3431,N_1204,N_188);
xnor U3432 (N_3432,N_1020,N_2395);
nor U3433 (N_3433,N_420,N_1703);
or U3434 (N_3434,N_1074,N_306);
and U3435 (N_3435,N_1464,N_2871);
and U3436 (N_3436,N_977,N_2618);
or U3437 (N_3437,N_2891,N_850);
and U3438 (N_3438,N_25,N_1101);
nor U3439 (N_3439,N_2876,N_310);
and U3440 (N_3440,N_1867,N_1521);
nor U3441 (N_3441,N_219,N_1115);
nand U3442 (N_3442,N_12,N_1067);
nand U3443 (N_3443,N_336,N_1981);
nand U3444 (N_3444,N_2897,N_490);
nor U3445 (N_3445,N_1543,N_1173);
xor U3446 (N_3446,N_669,N_1682);
xor U3447 (N_3447,N_240,N_707);
or U3448 (N_3448,N_1336,N_217);
nand U3449 (N_3449,N_1209,N_2981);
nor U3450 (N_3450,N_467,N_2597);
nor U3451 (N_3451,N_613,N_1601);
nand U3452 (N_3452,N_40,N_2872);
xor U3453 (N_3453,N_2606,N_2720);
and U3454 (N_3454,N_580,N_2902);
nand U3455 (N_3455,N_78,N_1446);
and U3456 (N_3456,N_119,N_1767);
xnor U3457 (N_3457,N_957,N_2779);
xor U3458 (N_3458,N_2341,N_2453);
nand U3459 (N_3459,N_0,N_1363);
xnor U3460 (N_3460,N_1623,N_2899);
xnor U3461 (N_3461,N_412,N_2770);
and U3462 (N_3462,N_1850,N_407);
nand U3463 (N_3463,N_2030,N_935);
and U3464 (N_3464,N_2393,N_378);
and U3465 (N_3465,N_1747,N_2279);
nand U3466 (N_3466,N_1914,N_174);
nor U3467 (N_3467,N_2780,N_354);
nor U3468 (N_3468,N_2098,N_32);
nand U3469 (N_3469,N_173,N_893);
or U3470 (N_3470,N_1439,N_2413);
nand U3471 (N_3471,N_1051,N_2302);
or U3472 (N_3472,N_523,N_1855);
or U3473 (N_3473,N_2975,N_2529);
nor U3474 (N_3474,N_128,N_2841);
nand U3475 (N_3475,N_1551,N_1749);
nor U3476 (N_3476,N_848,N_229);
nor U3477 (N_3477,N_1896,N_2392);
nand U3478 (N_3478,N_2846,N_914);
nand U3479 (N_3479,N_264,N_1200);
nand U3480 (N_3480,N_732,N_329);
nand U3481 (N_3481,N_1190,N_680);
and U3482 (N_3482,N_1580,N_2686);
xnor U3483 (N_3483,N_643,N_2807);
xnor U3484 (N_3484,N_1743,N_2502);
or U3485 (N_3485,N_597,N_828);
nand U3486 (N_3486,N_1199,N_165);
nand U3487 (N_3487,N_1434,N_942);
and U3488 (N_3488,N_1571,N_1216);
xor U3489 (N_3489,N_1489,N_1187);
nor U3490 (N_3490,N_1565,N_23);
and U3491 (N_3491,N_1265,N_774);
nor U3492 (N_3492,N_1283,N_1525);
nor U3493 (N_3493,N_571,N_2719);
and U3494 (N_3494,N_1485,N_259);
nand U3495 (N_3495,N_2658,N_731);
and U3496 (N_3496,N_2175,N_915);
and U3497 (N_3497,N_2660,N_2478);
xor U3498 (N_3498,N_2750,N_2967);
nand U3499 (N_3499,N_441,N_1785);
and U3500 (N_3500,N_2796,N_2609);
nor U3501 (N_3501,N_575,N_2608);
xnor U3502 (N_3502,N_485,N_2960);
xor U3503 (N_3503,N_1393,N_940);
or U3504 (N_3504,N_987,N_2155);
nand U3505 (N_3505,N_2246,N_2338);
xor U3506 (N_3506,N_502,N_2915);
xnor U3507 (N_3507,N_844,N_778);
or U3508 (N_3508,N_1765,N_498);
nor U3509 (N_3509,N_1275,N_1616);
and U3510 (N_3510,N_48,N_1877);
nor U3511 (N_3511,N_551,N_1925);
nor U3512 (N_3512,N_2200,N_1900);
nor U3513 (N_3513,N_73,N_616);
nor U3514 (N_3514,N_5,N_2663);
xnor U3515 (N_3515,N_1306,N_2318);
xor U3516 (N_3516,N_1174,N_662);
and U3517 (N_3517,N_315,N_2802);
nor U3518 (N_3518,N_370,N_1600);
or U3519 (N_3519,N_1236,N_2445);
nor U3520 (N_3520,N_369,N_1756);
nor U3521 (N_3521,N_116,N_2584);
or U3522 (N_3522,N_2574,N_2634);
and U3523 (N_3523,N_1398,N_2895);
xor U3524 (N_3524,N_854,N_2067);
nor U3525 (N_3525,N_1314,N_401);
xnor U3526 (N_3526,N_1462,N_2619);
or U3527 (N_3527,N_2772,N_666);
xnor U3528 (N_3528,N_1657,N_748);
nand U3529 (N_3529,N_1961,N_2798);
and U3530 (N_3530,N_2486,N_2074);
and U3531 (N_3531,N_1410,N_2998);
and U3532 (N_3532,N_513,N_2949);
nor U3533 (N_3533,N_2170,N_136);
xnor U3534 (N_3534,N_2685,N_1254);
and U3535 (N_3535,N_2254,N_715);
or U3536 (N_3536,N_134,N_745);
nand U3537 (N_3537,N_1820,N_1501);
xnor U3538 (N_3538,N_172,N_2731);
nor U3539 (N_3539,N_444,N_1655);
nor U3540 (N_3540,N_712,N_894);
or U3541 (N_3541,N_2151,N_9);
nor U3542 (N_3542,N_2569,N_2843);
and U3543 (N_3543,N_1019,N_1374);
and U3544 (N_3544,N_948,N_2378);
xnor U3545 (N_3545,N_1068,N_1624);
or U3546 (N_3546,N_2794,N_1015);
xor U3547 (N_3547,N_1277,N_95);
and U3548 (N_3548,N_2328,N_1897);
nand U3549 (N_3549,N_1936,N_1871);
or U3550 (N_3550,N_700,N_360);
or U3551 (N_3551,N_1430,N_2661);
or U3552 (N_3552,N_2111,N_269);
or U3553 (N_3553,N_2624,N_222);
nand U3554 (N_3554,N_395,N_410);
and U3555 (N_3555,N_146,N_545);
or U3556 (N_3556,N_1728,N_141);
nand U3557 (N_3557,N_2759,N_1341);
xnor U3558 (N_3558,N_2078,N_1859);
xor U3559 (N_3559,N_1351,N_1710);
and U3560 (N_3560,N_1134,N_4);
xor U3561 (N_3561,N_2369,N_2159);
or U3562 (N_3562,N_478,N_38);
nand U3563 (N_3563,N_2973,N_2421);
nor U3564 (N_3564,N_182,N_272);
nor U3565 (N_3565,N_863,N_2174);
xor U3566 (N_3566,N_1507,N_2728);
nand U3567 (N_3567,N_1266,N_2579);
nor U3568 (N_3568,N_769,N_852);
or U3569 (N_3569,N_1757,N_2550);
xor U3570 (N_3570,N_1255,N_2013);
xnor U3571 (N_3571,N_1413,N_2630);
or U3572 (N_3572,N_501,N_2387);
nor U3573 (N_3573,N_749,N_2261);
nand U3574 (N_3574,N_137,N_2315);
xnor U3575 (N_3575,N_13,N_809);
xor U3576 (N_3576,N_2068,N_1759);
nand U3577 (N_3577,N_1956,N_2805);
nor U3578 (N_3578,N_1474,N_1484);
and U3579 (N_3579,N_2601,N_67);
and U3580 (N_3580,N_999,N_2075);
and U3581 (N_3581,N_2379,N_1997);
xnor U3582 (N_3582,N_2783,N_1554);
and U3583 (N_3583,N_1344,N_2562);
or U3584 (N_3584,N_2600,N_1320);
nor U3585 (N_3585,N_849,N_2958);
xnor U3586 (N_3586,N_859,N_347);
nor U3587 (N_3587,N_2412,N_2002);
nor U3588 (N_3588,N_493,N_974);
or U3589 (N_3589,N_1329,N_1576);
nand U3590 (N_3590,N_1675,N_2784);
nand U3591 (N_3591,N_1372,N_1662);
and U3592 (N_3592,N_670,N_718);
or U3593 (N_3593,N_2781,N_1412);
nor U3594 (N_3594,N_2883,N_2654);
or U3595 (N_3595,N_2094,N_236);
xnor U3596 (N_3596,N_80,N_2229);
nand U3597 (N_3597,N_2414,N_1681);
and U3598 (N_3598,N_151,N_1026);
xor U3599 (N_3599,N_1251,N_751);
or U3600 (N_3600,N_1594,N_2893);
and U3601 (N_3601,N_2113,N_699);
or U3602 (N_3602,N_2904,N_2051);
xor U3603 (N_3603,N_588,N_1660);
or U3604 (N_3604,N_2038,N_1796);
or U3605 (N_3605,N_982,N_47);
or U3606 (N_3606,N_910,N_1826);
nor U3607 (N_3607,N_2473,N_1689);
nor U3608 (N_3608,N_1218,N_279);
or U3609 (N_3609,N_702,N_1899);
or U3610 (N_3610,N_1670,N_2423);
or U3611 (N_3611,N_1366,N_2570);
nand U3612 (N_3612,N_912,N_1460);
and U3613 (N_3613,N_2072,N_2052);
nand U3614 (N_3614,N_2273,N_2865);
nor U3615 (N_3615,N_529,N_2919);
and U3616 (N_3616,N_431,N_2097);
and U3617 (N_3617,N_1145,N_122);
nor U3618 (N_3618,N_2324,N_1592);
or U3619 (N_3619,N_2565,N_1110);
nor U3620 (N_3620,N_2757,N_2947);
and U3621 (N_3621,N_2046,N_284);
nor U3622 (N_3622,N_1378,N_2860);
and U3623 (N_3623,N_2148,N_1127);
xnor U3624 (N_3624,N_1864,N_2343);
and U3625 (N_3625,N_2288,N_1126);
xor U3626 (N_3626,N_1473,N_2234);
nor U3627 (N_3627,N_1980,N_1240);
or U3628 (N_3628,N_465,N_1272);
and U3629 (N_3629,N_2553,N_996);
nand U3630 (N_3630,N_1834,N_2110);
xnor U3631 (N_3631,N_2247,N_2687);
nor U3632 (N_3632,N_2399,N_2346);
xnor U3633 (N_3633,N_2541,N_2438);
nor U3634 (N_3634,N_1529,N_1803);
and U3635 (N_3635,N_517,N_2327);
xnor U3636 (N_3636,N_2137,N_978);
and U3637 (N_3637,N_1664,N_1777);
nand U3638 (N_3638,N_2187,N_1125);
and U3639 (N_3639,N_2105,N_540);
xnor U3640 (N_3640,N_953,N_163);
nand U3641 (N_3641,N_2350,N_1478);
xnor U3642 (N_3642,N_1424,N_783);
or U3643 (N_3643,N_2435,N_2220);
xor U3644 (N_3644,N_1745,N_2298);
nor U3645 (N_3645,N_1722,N_295);
nor U3646 (N_3646,N_2232,N_2592);
and U3647 (N_3647,N_2460,N_659);
or U3648 (N_3648,N_1285,N_2363);
nor U3649 (N_3649,N_1984,N_891);
xnor U3650 (N_3650,N_2001,N_149);
or U3651 (N_3651,N_2494,N_2737);
or U3652 (N_3652,N_1419,N_140);
xnor U3653 (N_3653,N_2555,N_1242);
or U3654 (N_3654,N_1208,N_1784);
and U3655 (N_3655,N_2539,N_2420);
and U3656 (N_3656,N_786,N_2268);
xor U3657 (N_3657,N_2427,N_964);
or U3658 (N_3658,N_621,N_169);
nor U3659 (N_3659,N_292,N_1992);
or U3660 (N_3660,N_1821,N_2277);
or U3661 (N_3661,N_2504,N_1002);
nor U3662 (N_3662,N_319,N_661);
or U3663 (N_3663,N_2886,N_2880);
xor U3664 (N_3664,N_1709,N_2507);
xnor U3665 (N_3665,N_1048,N_2868);
and U3666 (N_3666,N_2986,N_780);
and U3667 (N_3667,N_2956,N_2740);
or U3668 (N_3668,N_1502,N_761);
nand U3669 (N_3669,N_1888,N_779);
nand U3670 (N_3670,N_129,N_1373);
nor U3671 (N_3671,N_1586,N_1856);
nand U3672 (N_3672,N_2084,N_2826);
nand U3673 (N_3673,N_559,N_2989);
nor U3674 (N_3674,N_1232,N_2042);
xnor U3675 (N_3675,N_980,N_950);
nand U3676 (N_3676,N_928,N_326);
nand U3677 (N_3677,N_1776,N_1886);
or U3678 (N_3678,N_492,N_243);
or U3679 (N_3679,N_2590,N_2160);
nor U3680 (N_3680,N_6,N_926);
xor U3681 (N_3681,N_1783,N_2616);
or U3682 (N_3682,N_991,N_308);
nor U3683 (N_3683,N_2041,N_2455);
and U3684 (N_3684,N_2483,N_911);
xnor U3685 (N_3685,N_139,N_2776);
or U3686 (N_3686,N_1081,N_554);
or U3687 (N_3687,N_84,N_2142);
and U3688 (N_3688,N_946,N_2161);
and U3689 (N_3689,N_2571,N_608);
nand U3690 (N_3690,N_1755,N_1453);
nor U3691 (N_3691,N_582,N_1095);
xor U3692 (N_3692,N_634,N_1450);
nor U3693 (N_3693,N_1550,N_330);
or U3694 (N_3694,N_205,N_408);
nor U3695 (N_3695,N_1702,N_2697);
xnor U3696 (N_3696,N_2209,N_2884);
and U3697 (N_3697,N_210,N_1739);
nor U3698 (N_3698,N_2769,N_888);
or U3699 (N_3699,N_2683,N_2610);
nor U3700 (N_3700,N_2382,N_2169);
xnor U3701 (N_3701,N_1186,N_2198);
and U3702 (N_3702,N_385,N_1243);
nand U3703 (N_3703,N_2437,N_2199);
xnor U3704 (N_3704,N_432,N_674);
nand U3705 (N_3705,N_724,N_2914);
nor U3706 (N_3706,N_562,N_76);
xnor U3707 (N_3707,N_576,N_1316);
nor U3708 (N_3708,N_1628,N_2552);
and U3709 (N_3709,N_538,N_304);
xnor U3710 (N_3710,N_74,N_650);
or U3711 (N_3711,N_2523,N_256);
or U3712 (N_3712,N_2628,N_2901);
nor U3713 (N_3713,N_1432,N_2545);
nand U3714 (N_3714,N_1526,N_565);
xor U3715 (N_3715,N_2857,N_864);
nand U3716 (N_3716,N_428,N_1911);
xnor U3717 (N_3717,N_2117,N_2793);
nor U3718 (N_3718,N_2778,N_1640);
or U3719 (N_3719,N_2102,N_2994);
nor U3720 (N_3720,N_223,N_511);
xnor U3721 (N_3721,N_1852,N_1947);
nor U3722 (N_3722,N_667,N_983);
or U3723 (N_3723,N_1104,N_1500);
and U3724 (N_3724,N_1326,N_2452);
nand U3725 (N_3725,N_916,N_1189);
nand U3726 (N_3726,N_2214,N_1065);
or U3727 (N_3727,N_409,N_1438);
nand U3728 (N_3728,N_1528,N_362);
or U3729 (N_3729,N_768,N_1848);
or U3730 (N_3730,N_665,N_747);
nand U3731 (N_3731,N_695,N_2221);
xor U3732 (N_3732,N_1626,N_2185);
nand U3733 (N_3733,N_1459,N_1494);
nand U3734 (N_3734,N_2029,N_2401);
nor U3735 (N_3735,N_1452,N_2280);
or U3736 (N_3736,N_1465,N_1401);
and U3737 (N_3737,N_1654,N_1667);
nor U3738 (N_3738,N_1000,N_1975);
or U3739 (N_3739,N_1651,N_753);
nand U3740 (N_3740,N_1827,N_404);
or U3741 (N_3741,N_2890,N_1762);
xor U3742 (N_3742,N_1695,N_2707);
nand U3743 (N_3743,N_2830,N_1140);
nor U3744 (N_3744,N_2525,N_1904);
nand U3745 (N_3745,N_887,N_2212);
xor U3746 (N_3746,N_2675,N_484);
and U3747 (N_3747,N_1840,N_386);
or U3748 (N_3748,N_433,N_496);
or U3749 (N_3749,N_1691,N_2715);
xor U3750 (N_3750,N_487,N_1704);
xor U3751 (N_3751,N_1245,N_1404);
xnor U3752 (N_3752,N_2491,N_1168);
xnor U3753 (N_3753,N_2725,N_388);
nor U3754 (N_3754,N_2703,N_1971);
xnor U3755 (N_3755,N_1023,N_1912);
nand U3756 (N_3756,N_832,N_2526);
nor U3757 (N_3757,N_44,N_1967);
nor U3758 (N_3758,N_1228,N_2122);
nor U3759 (N_3759,N_2056,N_1838);
xor U3760 (N_3760,N_851,N_2997);
nor U3761 (N_3761,N_2979,N_2004);
and U3762 (N_3762,N_2524,N_1338);
nor U3763 (N_3763,N_1583,N_2184);
and U3764 (N_3764,N_1915,N_1717);
and U3765 (N_3765,N_53,N_446);
xnor U3766 (N_3766,N_682,N_881);
and U3767 (N_3767,N_595,N_2219);
and U3768 (N_3768,N_1807,N_2755);
and U3769 (N_3769,N_2317,N_1753);
or U3770 (N_3770,N_290,N_1052);
xnor U3771 (N_3771,N_266,N_1447);
and U3772 (N_3772,N_2347,N_1649);
nor U3773 (N_3773,N_158,N_2319);
nand U3774 (N_3774,N_1570,N_596);
or U3775 (N_3775,N_2385,N_1645);
or U3776 (N_3776,N_2205,N_1117);
or U3777 (N_3777,N_2669,N_2153);
nor U3778 (N_3778,N_1923,N_2577);
nand U3779 (N_3779,N_826,N_1865);
xnor U3780 (N_3780,N_1772,N_462);
nor U3781 (N_3781,N_1908,N_2849);
and U3782 (N_3782,N_2361,N_1920);
or U3783 (N_3783,N_14,N_483);
nand U3784 (N_3784,N_560,N_1619);
and U3785 (N_3785,N_1103,N_1319);
and U3786 (N_3786,N_2245,N_1790);
nand U3787 (N_3787,N_1045,N_1946);
xnor U3788 (N_3788,N_500,N_1532);
and U3789 (N_3789,N_1811,N_1049);
xnor U3790 (N_3790,N_144,N_8);
and U3791 (N_3791,N_328,N_2332);
or U3792 (N_3792,N_566,N_1027);
nor U3793 (N_3793,N_63,N_1175);
nand U3794 (N_3794,N_2838,N_2467);
xor U3795 (N_3795,N_2576,N_235);
xnor U3796 (N_3796,N_639,N_1635);
nor U3797 (N_3797,N_1471,N_563);
nor U3798 (N_3798,N_2371,N_1959);
xor U3799 (N_3799,N_1701,N_474);
or U3800 (N_3800,N_1792,N_1130);
nand U3801 (N_3801,N_642,N_2978);
and U3802 (N_3802,N_2516,N_824);
xnor U3803 (N_3803,N_1360,N_464);
nor U3804 (N_3804,N_2832,N_2124);
and U3805 (N_3805,N_2351,N_2887);
or U3806 (N_3806,N_2308,N_2812);
and U3807 (N_3807,N_1672,N_966);
or U3808 (N_3808,N_572,N_757);
nand U3809 (N_3809,N_797,N_425);
and U3810 (N_3810,N_856,N_1630);
nor U3811 (N_3811,N_1758,N_2218);
and U3812 (N_3812,N_2732,N_693);
and U3813 (N_3813,N_1906,N_1395);
xnor U3814 (N_3814,N_875,N_1422);
xnor U3815 (N_3815,N_2101,N_1530);
or U3816 (N_3816,N_1768,N_913);
xnor U3817 (N_3817,N_564,N_2342);
nand U3818 (N_3818,N_202,N_1440);
nor U3819 (N_3819,N_2442,N_1468);
nor U3820 (N_3820,N_1177,N_2181);
and U3821 (N_3821,N_1591,N_2678);
nand U3822 (N_3822,N_2023,N_2950);
xnor U3823 (N_3823,N_2580,N_1894);
or U3824 (N_3824,N_1621,N_380);
nand U3825 (N_3825,N_1256,N_107);
xor U3826 (N_3826,N_1427,N_275);
nand U3827 (N_3827,N_1873,N_416);
nand U3828 (N_3828,N_2513,N_1726);
nand U3829 (N_3829,N_2039,N_218);
xor U3830 (N_3830,N_533,N_578);
nor U3831 (N_3831,N_2814,N_706);
xor U3832 (N_3832,N_1399,N_884);
and U3833 (N_3833,N_1139,N_1544);
and U3834 (N_3834,N_257,N_2710);
nor U3835 (N_3835,N_261,N_2983);
nand U3836 (N_3836,N_1381,N_2639);
nor U3837 (N_3837,N_1511,N_2309);
xnor U3838 (N_3838,N_1181,N_762);
and U3839 (N_3839,N_2422,N_1647);
nor U3840 (N_3840,N_1585,N_2459);
nand U3841 (N_3841,N_2201,N_2594);
or U3842 (N_3842,N_2266,N_476);
xnor U3843 (N_3843,N_2712,N_1449);
nand U3844 (N_3844,N_2204,N_2432);
or U3845 (N_3845,N_623,N_1383);
nand U3846 (N_3846,N_605,N_2472);
nor U3847 (N_3847,N_2617,N_2536);
nor U3848 (N_3848,N_1353,N_1437);
nor U3849 (N_3849,N_847,N_842);
and U3850 (N_3850,N_344,N_2954);
nand U3851 (N_3851,N_1949,N_2511);
and U3852 (N_3852,N_1183,N_2026);
nand U3853 (N_3853,N_1451,N_2964);
nand U3854 (N_3854,N_1498,N_1694);
xnor U3855 (N_3855,N_1801,N_228);
or U3856 (N_3856,N_1286,N_1737);
xnor U3857 (N_3857,N_2957,N_1868);
or U3858 (N_3858,N_1426,N_921);
nand U3859 (N_3859,N_924,N_1963);
nor U3860 (N_3860,N_2476,N_2048);
and U3861 (N_3861,N_2415,N_989);
and U3862 (N_3862,N_2635,N_2892);
nor U3863 (N_3863,N_2464,N_2211);
or U3864 (N_3864,N_1257,N_1612);
and U3865 (N_3865,N_2968,N_2448);
and U3866 (N_3866,N_1804,N_2503);
and U3867 (N_3867,N_50,N_2171);
xor U3868 (N_3868,N_1198,N_516);
xor U3869 (N_3869,N_2595,N_2375);
or U3870 (N_3870,N_166,N_896);
and U3871 (N_3871,N_2647,N_2058);
nand U3872 (N_3872,N_2434,N_2984);
xnor U3873 (N_3873,N_1060,N_1905);
nand U3874 (N_3874,N_1832,N_1522);
or U3875 (N_3875,N_28,N_1487);
xor U3876 (N_3876,N_2990,N_2163);
and U3877 (N_3877,N_2620,N_574);
nand U3878 (N_3878,N_2065,N_2062);
xnor U3879 (N_3879,N_2564,N_1061);
or U3880 (N_3880,N_1671,N_2360);
and U3881 (N_3881,N_2520,N_1063);
nand U3882 (N_3882,N_1318,N_1418);
or U3883 (N_3883,N_250,N_296);
nor U3884 (N_3884,N_2227,N_341);
or U3885 (N_3885,N_2723,N_2933);
or U3886 (N_3886,N_2287,N_488);
and U3887 (N_3887,N_2644,N_2240);
xor U3888 (N_3888,N_1515,N_1405);
nor U3889 (N_3889,N_1922,N_427);
xnor U3890 (N_3890,N_1367,N_30);
or U3891 (N_3891,N_518,N_2746);
or U3892 (N_3892,N_442,N_522);
nor U3893 (N_3893,N_1152,N_2833);
nand U3894 (N_3894,N_2253,N_653);
nor U3895 (N_3895,N_2510,N_2301);
and U3896 (N_3896,N_356,N_1244);
and U3897 (N_3897,N_479,N_2196);
nand U3898 (N_3898,N_1352,N_1482);
and U3899 (N_3899,N_1615,N_1579);
nand U3900 (N_3900,N_1391,N_1119);
or U3901 (N_3901,N_1012,N_2275);
nor U3902 (N_3902,N_1510,N_2271);
xnor U3903 (N_3903,N_1350,N_2680);
xor U3904 (N_3904,N_2477,N_1118);
or U3905 (N_3905,N_2255,N_2096);
nand U3906 (N_3906,N_157,N_1929);
and U3907 (N_3907,N_2158,N_1420);
or U3908 (N_3908,N_802,N_735);
xnor U3909 (N_3909,N_2766,N_1071);
or U3910 (N_3910,N_392,N_1157);
xnor U3911 (N_3911,N_1409,N_2786);
and U3912 (N_3912,N_1179,N_2926);
nor U3913 (N_3913,N_453,N_2372);
nand U3914 (N_3914,N_489,N_2257);
and U3915 (N_3915,N_1977,N_2992);
or U3916 (N_3916,N_1659,N_1810);
nor U3917 (N_3917,N_270,N_207);
xor U3918 (N_3918,N_377,N_231);
nand U3919 (N_3919,N_96,N_1);
or U3920 (N_3920,N_127,N_1328);
or U3921 (N_3921,N_327,N_1917);
or U3922 (N_3922,N_716,N_1406);
nand U3923 (N_3923,N_2821,N_2125);
nand U3924 (N_3924,N_2649,N_2701);
xor U3925 (N_3925,N_690,N_1362);
and U3926 (N_3926,N_624,N_1202);
nor U3927 (N_3927,N_394,N_1661);
xnor U3928 (N_3928,N_1207,N_1217);
xor U3929 (N_3929,N_2295,N_2365);
nor U3930 (N_3930,N_2044,N_969);
and U3931 (N_3931,N_2444,N_2818);
and U3932 (N_3932,N_1596,N_472);
nand U3933 (N_3933,N_2400,N_2070);
xnor U3934 (N_3934,N_2010,N_1361);
and U3935 (N_3935,N_615,N_1169);
nand U3936 (N_3936,N_64,N_664);
or U3937 (N_3937,N_2294,N_132);
xor U3938 (N_3938,N_2016,N_2217);
nand U3939 (N_3939,N_263,N_2451);
or U3940 (N_3940,N_1952,N_62);
and U3941 (N_3941,N_2043,N_2036);
xor U3942 (N_3942,N_635,N_556);
and U3943 (N_3943,N_2930,N_785);
and U3944 (N_3944,N_584,N_2756);
and U3945 (N_3945,N_1237,N_2714);
and U3946 (N_3946,N_357,N_1469);
or U3947 (N_3947,N_810,N_285);
nand U3948 (N_3948,N_932,N_1128);
or U3949 (N_3949,N_1171,N_1964);
or U3950 (N_3950,N_1901,N_1192);
nor U3951 (N_3951,N_2411,N_1072);
xor U3952 (N_3952,N_2233,N_2167);
and U3953 (N_3953,N_1394,N_2825);
or U3954 (N_3954,N_1224,N_1496);
xor U3955 (N_3955,N_2446,N_121);
xor U3956 (N_3956,N_790,N_2559);
xnor U3957 (N_3957,N_2405,N_29);
nor U3958 (N_3958,N_754,N_2386);
or U3959 (N_3959,N_1678,N_524);
or U3960 (N_3960,N_2384,N_445);
and U3961 (N_3961,N_1384,N_1303);
nor U3962 (N_3962,N_1423,N_1836);
xnor U3963 (N_3963,N_1013,N_2894);
nor U3964 (N_3964,N_66,N_399);
and U3965 (N_3965,N_1454,N_2543);
or U3966 (N_3966,N_123,N_2180);
xor U3967 (N_3967,N_1597,N_1742);
xnor U3968 (N_3968,N_880,N_1159);
and U3969 (N_3969,N_2938,N_840);
nor U3970 (N_3970,N_2018,N_836);
or U3971 (N_3971,N_2310,N_1705);
xor U3972 (N_3972,N_813,N_2623);
and U3973 (N_3973,N_1881,N_1327);
nor U3974 (N_3974,N_1641,N_321);
and U3975 (N_3975,N_2582,N_727);
nand U3976 (N_3976,N_1642,N_2376);
nor U3977 (N_3977,N_2130,N_750);
or U3978 (N_3978,N_721,N_1738);
xnor U3979 (N_3979,N_2057,N_2863);
and U3980 (N_3980,N_2681,N_986);
nand U3981 (N_3981,N_2050,N_126);
xor U3982 (N_3982,N_1262,N_1301);
and U3983 (N_3983,N_2810,N_2397);
or U3984 (N_3984,N_860,N_2844);
nor U3985 (N_3985,N_2456,N_1723);
and U3986 (N_3986,N_1552,N_2760);
or U3987 (N_3987,N_1359,N_375);
and U3988 (N_3988,N_89,N_1637);
and U3989 (N_3989,N_413,N_2581);
xor U3990 (N_3990,N_1774,N_1725);
and U3991 (N_3991,N_1310,N_393);
or U3992 (N_3992,N_2593,N_1229);
xor U3993 (N_3993,N_1082,N_482);
and U3994 (N_3994,N_1885,N_567);
or U3995 (N_3995,N_2107,N_2598);
xor U3996 (N_3996,N_637,N_470);
nand U3997 (N_3997,N_15,N_2674);
nand U3998 (N_3998,N_997,N_1665);
and U3999 (N_3999,N_739,N_1203);
xnor U4000 (N_4000,N_543,N_2855);
nor U4001 (N_4001,N_2492,N_548);
nand U4002 (N_4002,N_252,N_1878);
and U4003 (N_4003,N_2842,N_317);
nand U4004 (N_4004,N_2747,N_791);
and U4005 (N_4005,N_742,N_2146);
and U4006 (N_4006,N_1941,N_1182);
and U4007 (N_4007,N_2498,N_1504);
xor U4008 (N_4008,N_193,N_2691);
or U4009 (N_4009,N_1304,N_473);
xnor U4010 (N_4010,N_1448,N_1116);
xnor U4011 (N_4011,N_1814,N_337);
and U4012 (N_4012,N_2742,N_992);
xor U4013 (N_4013,N_299,N_763);
and U4014 (N_4014,N_371,N_273);
xor U4015 (N_4015,N_2917,N_2312);
xor U4016 (N_4016,N_58,N_1590);
or U4017 (N_4017,N_2207,N_2357);
or U4018 (N_4018,N_525,N_1603);
nand U4019 (N_4019,N_1849,N_345);
xnor U4020 (N_4020,N_1998,N_1883);
nand U4021 (N_4021,N_1823,N_1212);
nor U4022 (N_4022,N_1077,N_2667);
or U4023 (N_4023,N_435,N_1031);
nor U4024 (N_4024,N_2995,N_2186);
or U4025 (N_4025,N_2532,N_324);
nor U4026 (N_4026,N_216,N_10);
nor U4027 (N_4027,N_1273,N_1937);
or U4028 (N_4028,N_1445,N_909);
nand U4029 (N_4029,N_2653,N_2497);
and U4030 (N_4030,N_2533,N_1697);
xnor U4031 (N_4031,N_2047,N_2518);
nand U4032 (N_4032,N_730,N_820);
and U4033 (N_4033,N_161,N_2722);
nand U4034 (N_4034,N_1167,N_1751);
or U4035 (N_4035,N_1120,N_1223);
xnor U4036 (N_4036,N_1004,N_43);
or U4037 (N_4037,N_367,N_2143);
nor U4038 (N_4038,N_2874,N_812);
or U4039 (N_4039,N_34,N_2853);
nor U4040 (N_4040,N_2612,N_481);
nor U4041 (N_4041,N_2815,N_625);
nor U4042 (N_4042,N_503,N_2022);
and U4043 (N_4043,N_1605,N_833);
or U4044 (N_4044,N_2463,N_720);
xor U4045 (N_4045,N_2262,N_2133);
and U4046 (N_4046,N_1752,N_951);
nor U4047 (N_4047,N_1566,N_542);
and U4048 (N_4048,N_1833,N_331);
xor U4049 (N_4049,N_590,N_2120);
nand U4050 (N_4050,N_1632,N_1491);
nand U4051 (N_4051,N_1197,N_577);
xor U4052 (N_4052,N_528,N_2751);
or U4053 (N_4053,N_1788,N_781);
xor U4054 (N_4054,N_897,N_2419);
nand U4055 (N_4055,N_1041,N_729);
xor U4056 (N_4056,N_2797,N_2519);
or U4057 (N_4057,N_1289,N_2267);
nor U4058 (N_4058,N_185,N_1599);
xor U4059 (N_4059,N_2333,N_504);
nor U4060 (N_4060,N_332,N_1402);
and U4061 (N_4061,N_2176,N_1582);
nor U4062 (N_4062,N_2191,N_2721);
nand U4063 (N_4063,N_933,N_1112);
nor U4064 (N_4064,N_1577,N_649);
xnor U4065 (N_4065,N_1331,N_2173);
and U4066 (N_4066,N_2627,N_2055);
nor U4067 (N_4067,N_922,N_1421);
nand U4068 (N_4068,N_929,N_1831);
xnor U4069 (N_4069,N_1512,N_215);
xor U4070 (N_4070,N_2140,N_1968);
and U4071 (N_4071,N_1017,N_1457);
xor U4072 (N_4072,N_491,N_1942);
nor U4073 (N_4073,N_507,N_2499);
nor U4074 (N_4074,N_1400,N_1692);
xor U4075 (N_4075,N_1086,N_2178);
nor U4076 (N_4076,N_1819,N_105);
xnor U4077 (N_4077,N_2976,N_1668);
and U4078 (N_4078,N_1337,N_2428);
nand U4079 (N_4079,N_2971,N_2813);
and U4080 (N_4080,N_301,N_1234);
or U4081 (N_4081,N_2054,N_1567);
nor U4082 (N_4082,N_349,N_2188);
nand U4083 (N_4083,N_1844,N_2189);
nor U4084 (N_4084,N_1239,N_376);
nand U4085 (N_4085,N_733,N_2296);
nand U4086 (N_4086,N_869,N_2561);
and U4087 (N_4087,N_834,N_2416);
and U4088 (N_4088,N_902,N_2905);
and U4089 (N_4089,N_736,N_164);
nand U4090 (N_4090,N_955,N_1142);
or U4091 (N_4091,N_1441,N_2852);
nand U4092 (N_4092,N_2935,N_2970);
or U4093 (N_4093,N_2588,N_2522);
or U4094 (N_4094,N_1493,N_2861);
and U4095 (N_4095,N_1939,N_2953);
or U4096 (N_4096,N_1436,N_254);
xor U4097 (N_4097,N_703,N_2596);
nand U4098 (N_4098,N_2291,N_1092);
xor U4099 (N_4099,N_450,N_2625);
xnor U4100 (N_4100,N_789,N_268);
nor U4101 (N_4101,N_1113,N_1046);
xnor U4102 (N_4102,N_2758,N_2402);
or U4103 (N_4103,N_1557,N_277);
xnor U4104 (N_4104,N_2394,N_1816);
and U4105 (N_4105,N_333,N_1317);
or U4106 (N_4106,N_1517,N_2431);
xnor U4107 (N_4107,N_2352,N_889);
or U4108 (N_4108,N_2648,N_2763);
and U4109 (N_4109,N_1889,N_746);
xnor U4110 (N_4110,N_2657,N_133);
or U4111 (N_4111,N_2753,N_2888);
nand U4112 (N_4112,N_1099,N_734);
or U4113 (N_4113,N_176,N_1131);
nand U4114 (N_4114,N_1869,N_2955);
or U4115 (N_4115,N_2804,N_2640);
or U4116 (N_4116,N_878,N_411);
nor U4117 (N_4117,N_2611,N_2493);
nor U4118 (N_4118,N_2283,N_1771);
nor U4119 (N_4119,N_2424,N_2040);
nor U4120 (N_4120,N_366,N_2256);
or U4121 (N_4121,N_81,N_853);
nand U4122 (N_4122,N_1069,N_309);
nand U4123 (N_4123,N_460,N_696);
or U4124 (N_4124,N_1038,N_2299);
and U4125 (N_4125,N_610,N_1153);
xor U4126 (N_4126,N_2695,N_114);
xor U4127 (N_4127,N_1088,N_962);
xnor U4128 (N_4128,N_267,N_686);
nor U4129 (N_4129,N_1696,N_1180);
xnor U4130 (N_4130,N_1568,N_1972);
or U4131 (N_4131,N_456,N_569);
xnor U4132 (N_4132,N_2069,N_2881);
nor U4133 (N_4133,N_609,N_984);
nand U4134 (N_4134,N_232,N_1261);
nand U4135 (N_4135,N_2077,N_2304);
nand U4136 (N_4136,N_1417,N_1356);
nor U4137 (N_4137,N_1227,N_305);
nand U4138 (N_4138,N_1987,N_530);
nand U4139 (N_4139,N_568,N_2425);
or U4140 (N_4140,N_509,N_814);
nand U4141 (N_4141,N_454,N_1537);
and U4142 (N_4142,N_59,N_845);
or U4143 (N_4143,N_1890,N_109);
or U4144 (N_4144,N_1625,N_1706);
xor U4145 (N_4145,N_2064,N_756);
nand U4146 (N_4146,N_2809,N_2364);
and U4147 (N_4147,N_2433,N_1279);
or U4148 (N_4148,N_895,N_1043);
nand U4149 (N_4149,N_1163,N_353);
nor U4150 (N_4150,N_629,N_2391);
or U4151 (N_4151,N_68,N_519);
nor U4152 (N_4152,N_2313,N_505);
xnor U4153 (N_4153,N_2790,N_2673);
xnor U4154 (N_4154,N_1652,N_2370);
or U4155 (N_4155,N_1919,N_839);
and U4156 (N_4156,N_2037,N_2534);
xnor U4157 (N_4157,N_1520,N_1797);
or U4158 (N_4158,N_1609,N_452);
xor U4159 (N_4159,N_1547,N_2150);
nor U4160 (N_4160,N_2194,N_1035);
or U4161 (N_4161,N_630,N_1411);
nand U4162 (N_4162,N_197,N_1541);
nand U4163 (N_4163,N_31,N_120);
or U4164 (N_4164,N_2637,N_440);
nor U4165 (N_4165,N_1486,N_2908);
and U4166 (N_4166,N_293,N_1033);
nor U4167 (N_4167,N_1721,N_1607);
nand U4168 (N_4168,N_495,N_2711);
and U4169 (N_4169,N_2059,N_594);
nor U4170 (N_4170,N_2754,N_1622);
xnor U4171 (N_4171,N_585,N_1892);
nand U4172 (N_4172,N_2636,N_271);
or U4173 (N_4173,N_2605,N_579);
or U4174 (N_4174,N_741,N_406);
nor U4175 (N_4175,N_2011,N_995);
and U4176 (N_4176,N_1927,N_2373);
nand U4177 (N_4177,N_2265,N_550);
nor U4178 (N_4178,N_2912,N_767);
nor U4179 (N_4179,N_2726,N_1763);
or U4180 (N_4180,N_2946,N_2903);
xor U4181 (N_4181,N_1648,N_71);
nand U4182 (N_4182,N_280,N_1862);
xnor U4183 (N_4183,N_1799,N_2548);
or U4184 (N_4184,N_961,N_2537);
or U4185 (N_4185,N_547,N_424);
nor U4186 (N_4186,N_1170,N_2782);
or U4187 (N_4187,N_1653,N_2388);
nand U4188 (N_4188,N_2730,N_1610);
nand U4189 (N_4189,N_1323,N_1477);
or U4190 (N_4190,N_927,N_1184);
and U4191 (N_4191,N_2787,N_255);
and U4192 (N_4192,N_2330,N_1007);
xor U4193 (N_4193,N_2337,N_274);
nor U4194 (N_4194,N_1010,N_1957);
xor U4195 (N_4195,N_822,N_632);
xnor U4196 (N_4196,N_1211,N_1658);
nor U4197 (N_4197,N_2222,N_2987);
nand U4198 (N_4198,N_1918,N_536);
nor U4199 (N_4199,N_177,N_2848);
nor U4200 (N_4200,N_204,N_1951);
and U4201 (N_4201,N_2090,N_41);
nand U4202 (N_4202,N_1492,N_2458);
and U4203 (N_4203,N_1829,N_2951);
and U4204 (N_4204,N_1281,N_2024);
or U4205 (N_4205,N_2689,N_2367);
nand U4206 (N_4206,N_1499,N_2980);
or U4207 (N_4207,N_2771,N_1686);
nand U4208 (N_4208,N_1150,N_2659);
xor U4209 (N_4209,N_2145,N_1874);
xor U4210 (N_4210,N_1416,N_2741);
nand U4211 (N_4211,N_2276,N_2471);
or U4212 (N_4212,N_1397,N_2114);
and U4213 (N_4213,N_418,N_2870);
xor U4214 (N_4214,N_113,N_54);
xnor U4215 (N_4215,N_943,N_773);
nand U4216 (N_4216,N_2297,N_49);
xnor U4217 (N_4217,N_2404,N_2670);
and U4218 (N_4218,N_2591,N_1851);
xnor U4219 (N_4219,N_1683,N_2496);
or U4220 (N_4220,N_278,N_846);
nand U4221 (N_4221,N_2777,N_713);
xor U4222 (N_4222,N_1893,N_1545);
xor U4223 (N_4223,N_1308,N_1995);
and U4224 (N_4224,N_1534,N_2665);
nand U4225 (N_4225,N_1291,N_2293);
and U4226 (N_4226,N_213,N_521);
nand U4227 (N_4227,N_725,N_1053);
or U4228 (N_4228,N_945,N_2840);
and U4229 (N_4229,N_701,N_1538);
and U4230 (N_4230,N_2235,N_7);
nand U4231 (N_4231,N_2076,N_2348);
or U4232 (N_4232,N_1926,N_2168);
xnor U4233 (N_4233,N_1791,N_199);
xnor U4234 (N_4234,N_2080,N_288);
nor U4235 (N_4235,N_1687,N_75);
xnor U4236 (N_4236,N_2005,N_2845);
xnor U4237 (N_4237,N_1312,N_1973);
xnor U4238 (N_4238,N_998,N_2156);
or U4239 (N_4239,N_138,N_1629);
and U4240 (N_4240,N_2447,N_2664);
and U4241 (N_4241,N_1001,N_787);
and U4242 (N_4242,N_1902,N_784);
and U4243 (N_4243,N_879,N_2449);
nand U4244 (N_4244,N_2264,N_2716);
xor U4245 (N_4245,N_1618,N_1058);
nand U4246 (N_4246,N_1215,N_2613);
xnor U4247 (N_4247,N_1644,N_2668);
or U4248 (N_4248,N_2713,N_514);
nand U4249 (N_4249,N_1780,N_2646);
or U4250 (N_4250,N_1135,N_1891);
and U4251 (N_4251,N_917,N_2479);
xnor U4252 (N_4252,N_2489,N_1824);
or U4253 (N_4253,N_1282,N_675);
nand U4254 (N_4254,N_2157,N_92);
or U4255 (N_4255,N_968,N_2243);
and U4256 (N_4256,N_486,N_1857);
or U4257 (N_4257,N_1064,N_2717);
or U4258 (N_4258,N_461,N_1729);
nand U4259 (N_4259,N_2739,N_1259);
xor U4260 (N_4260,N_2966,N_2501);
nor U4261 (N_4261,N_1540,N_1414);
nor U4262 (N_4262,N_843,N_1719);
and U4263 (N_4263,N_458,N_1056);
nand U4264 (N_4264,N_88,N_1222);
xnor U4265 (N_4265,N_115,N_2286);
nor U4266 (N_4266,N_1921,N_1090);
and U4267 (N_4267,N_60,N_291);
xnor U4268 (N_4268,N_1779,N_1479);
xor U4269 (N_4269,N_1983,N_2325);
nand U4270 (N_4270,N_1342,N_1724);
xnor U4271 (N_4271,N_86,N_2831);
and U4272 (N_4272,N_1231,N_2906);
or U4273 (N_4273,N_931,N_1711);
and U4274 (N_4274,N_1075,N_350);
nand U4275 (N_4275,N_148,N_2088);
or U4276 (N_4276,N_209,N_867);
and U4277 (N_4277,N_1674,N_1195);
xnor U4278 (N_4278,N_135,N_2866);
nand U4279 (N_4279,N_2128,N_2540);
nor U4280 (N_4280,N_1727,N_1111);
nor U4281 (N_4281,N_617,N_2662);
xor U4282 (N_4282,N_2224,N_2418);
nor U4283 (N_4283,N_668,N_1109);
or U4284 (N_4284,N_2316,N_1100);
or U4285 (N_4285,N_2733,N_2374);
and U4286 (N_4286,N_805,N_937);
nand U4287 (N_4287,N_106,N_2705);
or U4288 (N_4288,N_2877,N_2789);
xnor U4289 (N_4289,N_1380,N_51);
xnor U4290 (N_4290,N_455,N_117);
xor U4291 (N_4291,N_2940,N_803);
or U4292 (N_4292,N_2251,N_2775);
and U4293 (N_4293,N_323,N_1270);
xnor U4294 (N_4294,N_553,N_1221);
nand U4295 (N_4295,N_300,N_591);
xnor U4296 (N_4296,N_1201,N_1839);
nand U4297 (N_4297,N_1994,N_253);
or U4298 (N_4298,N_1766,N_2203);
or U4299 (N_4299,N_2179,N_1858);
and U4300 (N_4300,N_901,N_2307);
nor U4301 (N_4301,N_1650,N_2089);
or U4302 (N_4302,N_1143,N_2331);
nor U4303 (N_4303,N_1428,N_607);
or U4304 (N_4304,N_2834,N_1965);
and U4305 (N_4305,N_764,N_17);
xnor U4306 (N_4306,N_570,N_2567);
or U4307 (N_4307,N_175,N_2651);
nor U4308 (N_4308,N_2465,N_1969);
nand U4309 (N_4309,N_1475,N_2698);
nand U4310 (N_4310,N_2974,N_262);
and U4311 (N_4311,N_2336,N_1569);
nand U4312 (N_4312,N_976,N_1392);
and U4313 (N_4313,N_1966,N_1377);
or U4314 (N_4314,N_384,N_2410);
nor U4315 (N_4315,N_211,N_2546);
nand U4316 (N_4316,N_2676,N_1287);
xor U4317 (N_4317,N_1786,N_2396);
or U4318 (N_4318,N_1230,N_2768);
or U4319 (N_4319,N_11,N_900);
nor U4320 (N_4320,N_1903,N_2144);
nor U4321 (N_4321,N_1991,N_1299);
nand U4322 (N_4322,N_1340,N_965);
nor U4323 (N_4323,N_1588,N_2558);
nor U4324 (N_4324,N_171,N_939);
xnor U4325 (N_4325,N_320,N_534);
nor U4326 (N_4326,N_102,N_2944);
and U4327 (N_4327,N_1390,N_283);
nor U4328 (N_4328,N_2252,N_2622);
and U4329 (N_4329,N_2829,N_1633);
and U4330 (N_4330,N_2015,N_2743);
and U4331 (N_4331,N_2329,N_429);
xnor U4332 (N_4332,N_2009,N_941);
nor U4333 (N_4333,N_443,N_710);
and U4334 (N_4334,N_1205,N_1930);
xnor U4335 (N_4335,N_2027,N_1407);
xnor U4336 (N_4336,N_1036,N_2643);
nor U4337 (N_4337,N_1934,N_993);
and U4338 (N_4338,N_793,N_658);
or U4339 (N_4339,N_1593,N_1685);
or U4340 (N_4340,N_952,N_2008);
or U4341 (N_4341,N_1292,N_1910);
nor U4342 (N_4342,N_671,N_2942);
xnor U4343 (N_4343,N_2100,N_2706);
or U4344 (N_4344,N_2025,N_1573);
and U4345 (N_4345,N_294,N_2816);
nand U4346 (N_4346,N_1089,N_841);
nand U4347 (N_4347,N_1800,N_1503);
and U4348 (N_4348,N_2139,N_111);
nand U4349 (N_4349,N_2345,N_2436);
nand U4350 (N_4350,N_2909,N_1389);
nor U4351 (N_4351,N_681,N_644);
nand U4352 (N_4352,N_815,N_963);
nor U4353 (N_4353,N_1558,N_956);
and U4354 (N_4354,N_1562,N_2982);
and U4355 (N_4355,N_1133,N_2910);
and U4356 (N_4356,N_2450,N_685);
nand U4357 (N_4357,N_1188,N_2738);
or U4358 (N_4358,N_1813,N_2837);
nand U4359 (N_4359,N_1611,N_648);
xor U4360 (N_4360,N_1598,N_2530);
and U4361 (N_4361,N_162,N_2873);
and U4362 (N_4362,N_646,N_898);
nand U4363 (N_4363,N_1713,N_2300);
nand U4364 (N_4364,N_603,N_494);
and U4365 (N_4365,N_1841,N_796);
or U4366 (N_4366,N_990,N_2488);
or U4367 (N_4367,N_2824,N_2811);
or U4368 (N_4368,N_2801,N_1284);
nor U4369 (N_4369,N_694,N_2112);
or U4370 (N_4370,N_2417,N_2355);
or U4371 (N_4371,N_2147,N_2323);
nor U4372 (N_4372,N_2278,N_1733);
nor U4373 (N_4373,N_792,N_52);
nand U4374 (N_4374,N_890,N_355);
or U4375 (N_4375,N_2671,N_2952);
and U4376 (N_4376,N_1985,N_1241);
nand U4377 (N_4377,N_2381,N_765);
or U4378 (N_4378,N_1809,N_2696);
nor U4379 (N_4379,N_2197,N_83);
or U4380 (N_4380,N_604,N_1533);
xnor U4381 (N_4381,N_1760,N_744);
and U4382 (N_4382,N_1716,N_1225);
xor U4383 (N_4383,N_1238,N_506);
nand U4384 (N_4384,N_1907,N_2694);
xor U4385 (N_4385,N_2095,N_312);
or U4386 (N_4386,N_414,N_1037);
xnor U4387 (N_4387,N_1656,N_535);
xnor U4388 (N_4388,N_2819,N_2922);
or U4389 (N_4389,N_1909,N_1161);
or U4390 (N_4390,N_1219,N_1638);
nand U4391 (N_4391,N_2182,N_1782);
nand U4392 (N_4392,N_985,N_537);
or U4393 (N_4393,N_2626,N_2607);
nand U4394 (N_4394,N_298,N_87);
or U4395 (N_4395,N_858,N_2850);
nor U4396 (N_4396,N_1944,N_1024);
nand U4397 (N_4397,N_181,N_2119);
nor U4398 (N_4398,N_1516,N_1812);
nor U4399 (N_4399,N_633,N_1054);
nor U4400 (N_4400,N_1924,N_1875);
and U4401 (N_4401,N_1466,N_723);
nor U4402 (N_4402,N_2269,N_2642);
xnor U4403 (N_4403,N_1136,N_2454);
nor U4404 (N_4404,N_2306,N_2281);
nand U4405 (N_4405,N_42,N_678);
or U4406 (N_4406,N_1798,N_2822);
or U4407 (N_4407,N_2474,N_2241);
nand U4408 (N_4408,N_246,N_2334);
xor U4409 (N_4409,N_934,N_448);
and U4410 (N_4410,N_1680,N_2349);
nand U4411 (N_4411,N_2466,N_1764);
or U4412 (N_4412,N_1335,N_1750);
and U4413 (N_4413,N_2083,N_225);
nand U4414 (N_4414,N_2021,N_2923);
xnor U4415 (N_4415,N_2260,N_1191);
and U4416 (N_4416,N_818,N_807);
or U4417 (N_4417,N_2263,N_2134);
xnor U4418 (N_4418,N_1124,N_2032);
and U4419 (N_4419,N_1690,N_1084);
or U4420 (N_4420,N_1156,N_82);
nand U4421 (N_4421,N_2859,N_57);
nand U4422 (N_4422,N_1016,N_2839);
or U4423 (N_4423,N_873,N_1057);
or U4424 (N_4424,N_1748,N_2991);
xor U4425 (N_4425,N_358,N_1989);
nor U4426 (N_4426,N_1264,N_645);
and U4427 (N_4427,N_1999,N_1248);
xnor U4428 (N_4428,N_808,N_1334);
or U4429 (N_4429,N_930,N_862);
or U4430 (N_4430,N_2688,N_2996);
and U4431 (N_4431,N_451,N_1744);
nand U4432 (N_4432,N_423,N_1313);
xnor U4433 (N_4433,N_104,N_2631);
or U4434 (N_4434,N_1982,N_1505);
nand U4435 (N_4435,N_2172,N_1553);
nand U4436 (N_4436,N_2129,N_1861);
or U4437 (N_4437,N_2585,N_1311);
xnor U4438 (N_4438,N_2700,N_242);
nor U4439 (N_4439,N_338,N_883);
or U4440 (N_4440,N_244,N_1620);
xor U4441 (N_4441,N_2377,N_238);
xnor U4442 (N_4442,N_855,N_640);
xnor U4443 (N_4443,N_248,N_154);
or U4444 (N_4444,N_391,N_2061);
xnor U4445 (N_4445,N_2684,N_2547);
nand U4446 (N_4446,N_201,N_1863);
or U4447 (N_4447,N_2326,N_1773);
or U4448 (N_4448,N_372,N_698);
or U4449 (N_4449,N_656,N_1029);
xnor U4450 (N_4450,N_2602,N_2344);
nor U4451 (N_4451,N_405,N_2335);
or U4452 (N_4452,N_2936,N_1296);
nor U4453 (N_4453,N_557,N_2977);
xnor U4454 (N_4454,N_421,N_1673);
or U4455 (N_4455,N_2527,N_2226);
or U4456 (N_4456,N_647,N_36);
xor U4457 (N_4457,N_679,N_1913);
or U4458 (N_4458,N_1403,N_234);
nand U4459 (N_4459,N_2303,N_1005);
or U4460 (N_4460,N_1158,N_1866);
nor U4461 (N_4461,N_2081,N_2430);
or U4462 (N_4462,N_400,N_1847);
or U4463 (N_4463,N_180,N_2439);
nand U4464 (N_4464,N_868,N_1548);
and U4465 (N_4465,N_549,N_2650);
xnor U4466 (N_4466,N_390,N_2999);
nand U4467 (N_4467,N_1295,N_396);
nand U4468 (N_4468,N_226,N_882);
nand U4469 (N_4469,N_398,N_2087);
or U4470 (N_4470,N_1872,N_463);
nand U4471 (N_4471,N_2398,N_1070);
nand U4472 (N_4472,N_2340,N_821);
xor U4473 (N_4473,N_871,N_56);
nand U4474 (N_4474,N_1978,N_688);
nand U4475 (N_4475,N_947,N_457);
nor U4476 (N_4476,N_975,N_676);
nor U4477 (N_4477,N_1608,N_2879);
xnor U4478 (N_4478,N_1268,N_436);
and U4479 (N_4479,N_2882,N_2481);
nor U4480 (N_4480,N_2641,N_334);
xor U4481 (N_4481,N_2889,N_2082);
and U4482 (N_4482,N_2085,N_1220);
and U4483 (N_4483,N_1369,N_1795);
nor U4484 (N_4484,N_2939,N_1708);
nand U4485 (N_4485,N_2708,N_612);
or U4486 (N_4486,N_2000,N_1574);
xor U4487 (N_4487,N_2216,N_147);
xor U4488 (N_4488,N_627,N_18);
xor U4489 (N_4489,N_1382,N_2972);
and U4490 (N_4490,N_1561,N_2672);
xor U4491 (N_4491,N_2587,N_131);
nand U4492 (N_4492,N_2572,N_1712);
nor U4493 (N_4493,N_704,N_611);
nand U4494 (N_4494,N_2557,N_1895);
or U4495 (N_4495,N_1300,N_708);
and U4496 (N_4496,N_970,N_558);
and U4497 (N_4497,N_1481,N_1884);
or U4498 (N_4498,N_153,N_526);
or U4499 (N_4499,N_816,N_2538);
xnor U4500 (N_4500,N_2938,N_1786);
nand U4501 (N_4501,N_721,N_2114);
nand U4502 (N_4502,N_312,N_1683);
or U4503 (N_4503,N_2791,N_1605);
or U4504 (N_4504,N_701,N_48);
xor U4505 (N_4505,N_750,N_2216);
nor U4506 (N_4506,N_599,N_820);
xor U4507 (N_4507,N_579,N_1977);
nand U4508 (N_4508,N_1841,N_2800);
nand U4509 (N_4509,N_534,N_1617);
nor U4510 (N_4510,N_2768,N_2246);
or U4511 (N_4511,N_224,N_2137);
nand U4512 (N_4512,N_354,N_2442);
nor U4513 (N_4513,N_2723,N_277);
nand U4514 (N_4514,N_1552,N_2188);
nor U4515 (N_4515,N_544,N_1216);
or U4516 (N_4516,N_1609,N_2702);
xnor U4517 (N_4517,N_165,N_329);
xnor U4518 (N_4518,N_2354,N_323);
nor U4519 (N_4519,N_2096,N_2017);
nor U4520 (N_4520,N_1840,N_1145);
xnor U4521 (N_4521,N_1955,N_290);
xnor U4522 (N_4522,N_1713,N_2934);
or U4523 (N_4523,N_2372,N_1830);
nand U4524 (N_4524,N_2126,N_2722);
nor U4525 (N_4525,N_102,N_1865);
nor U4526 (N_4526,N_2595,N_437);
or U4527 (N_4527,N_2511,N_347);
xnor U4528 (N_4528,N_901,N_2773);
xnor U4529 (N_4529,N_1135,N_1182);
nor U4530 (N_4530,N_963,N_1792);
nand U4531 (N_4531,N_894,N_342);
nand U4532 (N_4532,N_1698,N_2228);
xnor U4533 (N_4533,N_485,N_1353);
xnor U4534 (N_4534,N_13,N_2476);
nor U4535 (N_4535,N_1768,N_216);
and U4536 (N_4536,N_2383,N_1944);
nor U4537 (N_4537,N_1787,N_521);
and U4538 (N_4538,N_1729,N_2275);
nor U4539 (N_4539,N_1689,N_2021);
nand U4540 (N_4540,N_964,N_1365);
nand U4541 (N_4541,N_348,N_11);
nand U4542 (N_4542,N_1288,N_2090);
and U4543 (N_4543,N_334,N_2472);
nor U4544 (N_4544,N_1436,N_2704);
xor U4545 (N_4545,N_1721,N_564);
xor U4546 (N_4546,N_3,N_2771);
and U4547 (N_4547,N_2455,N_2184);
nor U4548 (N_4548,N_615,N_2461);
and U4549 (N_4549,N_1329,N_2999);
and U4550 (N_4550,N_53,N_2836);
or U4551 (N_4551,N_135,N_1946);
or U4552 (N_4552,N_1113,N_2678);
and U4553 (N_4553,N_1186,N_363);
or U4554 (N_4554,N_872,N_1557);
or U4555 (N_4555,N_421,N_2237);
xnor U4556 (N_4556,N_1198,N_481);
or U4557 (N_4557,N_2517,N_1060);
or U4558 (N_4558,N_2677,N_1330);
or U4559 (N_4559,N_429,N_2707);
and U4560 (N_4560,N_1664,N_251);
nand U4561 (N_4561,N_996,N_2011);
nand U4562 (N_4562,N_726,N_285);
or U4563 (N_4563,N_1577,N_2098);
nor U4564 (N_4564,N_2989,N_2168);
and U4565 (N_4565,N_2811,N_2063);
nand U4566 (N_4566,N_2661,N_2125);
and U4567 (N_4567,N_2364,N_355);
and U4568 (N_4568,N_583,N_1029);
xnor U4569 (N_4569,N_117,N_2057);
nand U4570 (N_4570,N_80,N_1500);
xor U4571 (N_4571,N_938,N_39);
and U4572 (N_4572,N_2568,N_2205);
and U4573 (N_4573,N_794,N_389);
or U4574 (N_4574,N_2619,N_78);
and U4575 (N_4575,N_2614,N_1059);
xor U4576 (N_4576,N_2273,N_2596);
and U4577 (N_4577,N_535,N_250);
or U4578 (N_4578,N_2474,N_2935);
and U4579 (N_4579,N_902,N_2382);
nor U4580 (N_4580,N_893,N_563);
or U4581 (N_4581,N_2964,N_2471);
or U4582 (N_4582,N_1415,N_937);
nand U4583 (N_4583,N_2348,N_1534);
or U4584 (N_4584,N_623,N_588);
nand U4585 (N_4585,N_645,N_2779);
or U4586 (N_4586,N_1418,N_168);
or U4587 (N_4587,N_149,N_2741);
or U4588 (N_4588,N_89,N_643);
nand U4589 (N_4589,N_884,N_2134);
and U4590 (N_4590,N_294,N_1840);
nor U4591 (N_4591,N_300,N_2426);
nand U4592 (N_4592,N_684,N_483);
nand U4593 (N_4593,N_799,N_2026);
and U4594 (N_4594,N_2272,N_990);
and U4595 (N_4595,N_2250,N_1539);
nor U4596 (N_4596,N_2026,N_1583);
xor U4597 (N_4597,N_1951,N_2695);
and U4598 (N_4598,N_2898,N_2159);
nand U4599 (N_4599,N_147,N_2667);
nand U4600 (N_4600,N_2594,N_1212);
or U4601 (N_4601,N_2900,N_229);
or U4602 (N_4602,N_1493,N_1680);
xnor U4603 (N_4603,N_698,N_2828);
or U4604 (N_4604,N_410,N_544);
or U4605 (N_4605,N_261,N_1561);
nand U4606 (N_4606,N_1693,N_1715);
and U4607 (N_4607,N_2532,N_123);
nor U4608 (N_4608,N_1600,N_1088);
or U4609 (N_4609,N_2854,N_2029);
and U4610 (N_4610,N_1756,N_2585);
and U4611 (N_4611,N_2051,N_1675);
xor U4612 (N_4612,N_1122,N_999);
or U4613 (N_4613,N_958,N_2926);
and U4614 (N_4614,N_2410,N_2450);
xor U4615 (N_4615,N_503,N_351);
or U4616 (N_4616,N_2196,N_743);
or U4617 (N_4617,N_801,N_503);
or U4618 (N_4618,N_1224,N_2165);
xor U4619 (N_4619,N_455,N_1967);
and U4620 (N_4620,N_2230,N_454);
and U4621 (N_4621,N_2928,N_1409);
nand U4622 (N_4622,N_2374,N_1644);
or U4623 (N_4623,N_1703,N_1939);
or U4624 (N_4624,N_2470,N_1972);
nand U4625 (N_4625,N_2819,N_590);
xnor U4626 (N_4626,N_1959,N_710);
nor U4627 (N_4627,N_1834,N_1256);
xnor U4628 (N_4628,N_1463,N_265);
and U4629 (N_4629,N_2400,N_2257);
and U4630 (N_4630,N_1068,N_1272);
nor U4631 (N_4631,N_700,N_2893);
xnor U4632 (N_4632,N_443,N_331);
and U4633 (N_4633,N_2085,N_2288);
xor U4634 (N_4634,N_144,N_268);
nand U4635 (N_4635,N_2377,N_1639);
nand U4636 (N_4636,N_2667,N_2545);
xnor U4637 (N_4637,N_772,N_2475);
and U4638 (N_4638,N_1659,N_1921);
and U4639 (N_4639,N_2584,N_2841);
nor U4640 (N_4640,N_918,N_1294);
nor U4641 (N_4641,N_4,N_219);
nand U4642 (N_4642,N_2084,N_1047);
nor U4643 (N_4643,N_1257,N_1754);
or U4644 (N_4644,N_1329,N_1879);
xor U4645 (N_4645,N_586,N_1690);
xnor U4646 (N_4646,N_1355,N_1079);
and U4647 (N_4647,N_442,N_176);
xnor U4648 (N_4648,N_623,N_1536);
nor U4649 (N_4649,N_1089,N_2547);
or U4650 (N_4650,N_508,N_2435);
nand U4651 (N_4651,N_2665,N_1775);
nor U4652 (N_4652,N_1742,N_1869);
nand U4653 (N_4653,N_2900,N_718);
nor U4654 (N_4654,N_2897,N_1397);
nand U4655 (N_4655,N_1415,N_1199);
and U4656 (N_4656,N_2788,N_111);
or U4657 (N_4657,N_447,N_2566);
xnor U4658 (N_4658,N_102,N_979);
or U4659 (N_4659,N_1509,N_489);
xnor U4660 (N_4660,N_1308,N_0);
and U4661 (N_4661,N_2573,N_1381);
and U4662 (N_4662,N_154,N_448);
nor U4663 (N_4663,N_321,N_2998);
nand U4664 (N_4664,N_2430,N_2422);
or U4665 (N_4665,N_1067,N_2131);
nor U4666 (N_4666,N_2030,N_1831);
xor U4667 (N_4667,N_1728,N_2192);
nand U4668 (N_4668,N_704,N_2236);
xnor U4669 (N_4669,N_1535,N_335);
or U4670 (N_4670,N_142,N_684);
or U4671 (N_4671,N_1880,N_2299);
nand U4672 (N_4672,N_607,N_1638);
and U4673 (N_4673,N_357,N_762);
xor U4674 (N_4674,N_1976,N_1349);
nor U4675 (N_4675,N_1227,N_569);
nand U4676 (N_4676,N_2545,N_174);
or U4677 (N_4677,N_377,N_2943);
nand U4678 (N_4678,N_2821,N_2175);
or U4679 (N_4679,N_1931,N_312);
nand U4680 (N_4680,N_822,N_2628);
nand U4681 (N_4681,N_1798,N_2727);
xor U4682 (N_4682,N_2585,N_1319);
and U4683 (N_4683,N_627,N_2023);
xor U4684 (N_4684,N_922,N_253);
or U4685 (N_4685,N_1315,N_1567);
nor U4686 (N_4686,N_487,N_1131);
nor U4687 (N_4687,N_2901,N_1986);
nand U4688 (N_4688,N_2958,N_1630);
nor U4689 (N_4689,N_2539,N_2945);
nand U4690 (N_4690,N_955,N_2344);
and U4691 (N_4691,N_1429,N_2613);
or U4692 (N_4692,N_2348,N_1674);
and U4693 (N_4693,N_2199,N_2047);
nor U4694 (N_4694,N_890,N_262);
nand U4695 (N_4695,N_1147,N_236);
and U4696 (N_4696,N_2582,N_1838);
or U4697 (N_4697,N_2916,N_112);
xnor U4698 (N_4698,N_2510,N_2160);
or U4699 (N_4699,N_632,N_1681);
or U4700 (N_4700,N_1658,N_2546);
xnor U4701 (N_4701,N_1117,N_1240);
and U4702 (N_4702,N_1406,N_1962);
nor U4703 (N_4703,N_605,N_143);
and U4704 (N_4704,N_1989,N_2731);
xnor U4705 (N_4705,N_2684,N_2746);
nand U4706 (N_4706,N_85,N_1231);
nand U4707 (N_4707,N_962,N_1242);
or U4708 (N_4708,N_2704,N_228);
nor U4709 (N_4709,N_740,N_1767);
and U4710 (N_4710,N_1596,N_277);
nor U4711 (N_4711,N_2952,N_1815);
and U4712 (N_4712,N_554,N_2114);
nor U4713 (N_4713,N_2656,N_567);
nor U4714 (N_4714,N_1938,N_1323);
nand U4715 (N_4715,N_1446,N_2626);
nand U4716 (N_4716,N_2789,N_220);
nor U4717 (N_4717,N_1349,N_1129);
xnor U4718 (N_4718,N_1790,N_1617);
and U4719 (N_4719,N_2033,N_133);
nor U4720 (N_4720,N_1827,N_436);
or U4721 (N_4721,N_870,N_1113);
or U4722 (N_4722,N_175,N_1629);
or U4723 (N_4723,N_2159,N_678);
and U4724 (N_4724,N_2119,N_576);
nor U4725 (N_4725,N_324,N_1878);
or U4726 (N_4726,N_2355,N_1560);
nor U4727 (N_4727,N_399,N_1838);
xnor U4728 (N_4728,N_2124,N_635);
or U4729 (N_4729,N_1842,N_1556);
or U4730 (N_4730,N_2226,N_277);
nor U4731 (N_4731,N_1475,N_2680);
and U4732 (N_4732,N_2229,N_822);
xnor U4733 (N_4733,N_2066,N_2421);
or U4734 (N_4734,N_522,N_2774);
nand U4735 (N_4735,N_2704,N_808);
xnor U4736 (N_4736,N_573,N_2037);
or U4737 (N_4737,N_1818,N_563);
xnor U4738 (N_4738,N_2873,N_2468);
and U4739 (N_4739,N_565,N_1270);
xnor U4740 (N_4740,N_33,N_2539);
or U4741 (N_4741,N_338,N_1448);
nor U4742 (N_4742,N_2462,N_1234);
nand U4743 (N_4743,N_1053,N_328);
or U4744 (N_4744,N_91,N_447);
nor U4745 (N_4745,N_380,N_1806);
or U4746 (N_4746,N_1882,N_841);
nand U4747 (N_4747,N_2062,N_2004);
xor U4748 (N_4748,N_2749,N_787);
nor U4749 (N_4749,N_2991,N_267);
xor U4750 (N_4750,N_940,N_397);
nor U4751 (N_4751,N_1046,N_1648);
nand U4752 (N_4752,N_1940,N_898);
xnor U4753 (N_4753,N_2515,N_2259);
xnor U4754 (N_4754,N_2079,N_454);
or U4755 (N_4755,N_1405,N_1382);
and U4756 (N_4756,N_400,N_2488);
or U4757 (N_4757,N_2946,N_1503);
nand U4758 (N_4758,N_2581,N_2949);
and U4759 (N_4759,N_1333,N_1471);
nand U4760 (N_4760,N_1953,N_1851);
or U4761 (N_4761,N_414,N_191);
xnor U4762 (N_4762,N_1631,N_1476);
and U4763 (N_4763,N_1523,N_2995);
or U4764 (N_4764,N_2909,N_425);
nand U4765 (N_4765,N_766,N_242);
nor U4766 (N_4766,N_83,N_1427);
xor U4767 (N_4767,N_71,N_1209);
and U4768 (N_4768,N_2265,N_1102);
and U4769 (N_4769,N_1520,N_891);
nor U4770 (N_4770,N_784,N_2285);
xnor U4771 (N_4771,N_2523,N_1162);
nand U4772 (N_4772,N_7,N_546);
nor U4773 (N_4773,N_1513,N_116);
xnor U4774 (N_4774,N_363,N_1815);
xnor U4775 (N_4775,N_962,N_631);
or U4776 (N_4776,N_1493,N_2181);
xnor U4777 (N_4777,N_153,N_46);
nand U4778 (N_4778,N_1965,N_2306);
nand U4779 (N_4779,N_546,N_1632);
xnor U4780 (N_4780,N_872,N_1228);
or U4781 (N_4781,N_505,N_495);
nand U4782 (N_4782,N_2405,N_1772);
nor U4783 (N_4783,N_2687,N_111);
nor U4784 (N_4784,N_2532,N_1801);
xnor U4785 (N_4785,N_1664,N_2438);
or U4786 (N_4786,N_2960,N_2777);
nand U4787 (N_4787,N_1863,N_1418);
and U4788 (N_4788,N_399,N_2929);
nor U4789 (N_4789,N_596,N_1886);
xor U4790 (N_4790,N_1781,N_69);
and U4791 (N_4791,N_882,N_34);
and U4792 (N_4792,N_1894,N_1533);
and U4793 (N_4793,N_1291,N_1232);
or U4794 (N_4794,N_2934,N_2285);
nor U4795 (N_4795,N_831,N_1149);
or U4796 (N_4796,N_819,N_1599);
and U4797 (N_4797,N_2196,N_2134);
and U4798 (N_4798,N_805,N_2658);
or U4799 (N_4799,N_1385,N_2783);
and U4800 (N_4800,N_251,N_1959);
xor U4801 (N_4801,N_1655,N_1332);
xnor U4802 (N_4802,N_1155,N_862);
nand U4803 (N_4803,N_872,N_1079);
nor U4804 (N_4804,N_2452,N_1200);
nand U4805 (N_4805,N_1473,N_2394);
or U4806 (N_4806,N_2252,N_1633);
nand U4807 (N_4807,N_766,N_1688);
and U4808 (N_4808,N_1591,N_1127);
nor U4809 (N_4809,N_1873,N_987);
nor U4810 (N_4810,N_1424,N_2443);
nand U4811 (N_4811,N_553,N_529);
or U4812 (N_4812,N_1263,N_2284);
nor U4813 (N_4813,N_2594,N_1344);
or U4814 (N_4814,N_1964,N_1119);
nand U4815 (N_4815,N_877,N_1609);
nand U4816 (N_4816,N_1176,N_1563);
and U4817 (N_4817,N_966,N_2883);
or U4818 (N_4818,N_2251,N_710);
or U4819 (N_4819,N_2871,N_1394);
and U4820 (N_4820,N_2072,N_2314);
xnor U4821 (N_4821,N_1786,N_706);
nor U4822 (N_4822,N_1066,N_1);
or U4823 (N_4823,N_323,N_1386);
and U4824 (N_4824,N_204,N_1604);
or U4825 (N_4825,N_1123,N_2353);
or U4826 (N_4826,N_58,N_225);
nor U4827 (N_4827,N_81,N_2673);
nor U4828 (N_4828,N_2986,N_1981);
and U4829 (N_4829,N_1590,N_1763);
xnor U4830 (N_4830,N_157,N_761);
or U4831 (N_4831,N_1277,N_1144);
nor U4832 (N_4832,N_1305,N_2959);
and U4833 (N_4833,N_2888,N_707);
nand U4834 (N_4834,N_1071,N_1949);
and U4835 (N_4835,N_2108,N_2094);
nand U4836 (N_4836,N_702,N_408);
and U4837 (N_4837,N_1258,N_475);
nor U4838 (N_4838,N_548,N_2952);
nand U4839 (N_4839,N_2001,N_1450);
or U4840 (N_4840,N_765,N_2778);
nand U4841 (N_4841,N_2028,N_611);
and U4842 (N_4842,N_260,N_1178);
and U4843 (N_4843,N_1210,N_1930);
nor U4844 (N_4844,N_677,N_2815);
xor U4845 (N_4845,N_78,N_2659);
and U4846 (N_4846,N_1770,N_1956);
and U4847 (N_4847,N_556,N_2019);
xnor U4848 (N_4848,N_2241,N_1098);
xor U4849 (N_4849,N_176,N_1153);
xnor U4850 (N_4850,N_521,N_1906);
nor U4851 (N_4851,N_2326,N_2842);
nand U4852 (N_4852,N_2370,N_1150);
or U4853 (N_4853,N_284,N_2166);
or U4854 (N_4854,N_1084,N_66);
nor U4855 (N_4855,N_312,N_252);
nor U4856 (N_4856,N_1180,N_529);
or U4857 (N_4857,N_2878,N_2091);
nand U4858 (N_4858,N_2376,N_1640);
xnor U4859 (N_4859,N_927,N_385);
or U4860 (N_4860,N_788,N_2721);
nand U4861 (N_4861,N_2325,N_2266);
and U4862 (N_4862,N_2104,N_627);
and U4863 (N_4863,N_838,N_2020);
and U4864 (N_4864,N_542,N_392);
xnor U4865 (N_4865,N_1929,N_2620);
and U4866 (N_4866,N_1373,N_1686);
or U4867 (N_4867,N_1432,N_2935);
nor U4868 (N_4868,N_1504,N_1858);
nor U4869 (N_4869,N_1051,N_2058);
xnor U4870 (N_4870,N_1483,N_2911);
and U4871 (N_4871,N_841,N_1324);
nor U4872 (N_4872,N_1603,N_338);
nor U4873 (N_4873,N_2262,N_2416);
xnor U4874 (N_4874,N_2075,N_1863);
nand U4875 (N_4875,N_54,N_2716);
or U4876 (N_4876,N_506,N_843);
or U4877 (N_4877,N_193,N_839);
nand U4878 (N_4878,N_277,N_2578);
nor U4879 (N_4879,N_2543,N_1564);
nor U4880 (N_4880,N_162,N_1795);
or U4881 (N_4881,N_2602,N_167);
or U4882 (N_4882,N_2923,N_893);
xor U4883 (N_4883,N_2187,N_2930);
nor U4884 (N_4884,N_1771,N_82);
xor U4885 (N_4885,N_1639,N_2660);
or U4886 (N_4886,N_1637,N_1297);
nand U4887 (N_4887,N_141,N_174);
nand U4888 (N_4888,N_288,N_805);
nor U4889 (N_4889,N_2057,N_1281);
or U4890 (N_4890,N_2758,N_1350);
nand U4891 (N_4891,N_1401,N_718);
nand U4892 (N_4892,N_1845,N_400);
and U4893 (N_4893,N_228,N_210);
nor U4894 (N_4894,N_580,N_778);
nand U4895 (N_4895,N_2753,N_1310);
xnor U4896 (N_4896,N_242,N_2218);
or U4897 (N_4897,N_1814,N_1003);
nor U4898 (N_4898,N_2711,N_594);
nor U4899 (N_4899,N_2939,N_667);
nor U4900 (N_4900,N_550,N_1499);
nand U4901 (N_4901,N_1885,N_2713);
or U4902 (N_4902,N_938,N_2697);
xnor U4903 (N_4903,N_1186,N_2043);
and U4904 (N_4904,N_1878,N_2259);
and U4905 (N_4905,N_885,N_749);
xnor U4906 (N_4906,N_1350,N_557);
or U4907 (N_4907,N_2093,N_352);
nand U4908 (N_4908,N_172,N_2368);
nor U4909 (N_4909,N_553,N_168);
nor U4910 (N_4910,N_787,N_2752);
and U4911 (N_4911,N_2789,N_1971);
or U4912 (N_4912,N_2520,N_921);
and U4913 (N_4913,N_717,N_790);
nor U4914 (N_4914,N_2486,N_2754);
xnor U4915 (N_4915,N_2284,N_2281);
and U4916 (N_4916,N_2155,N_1795);
nand U4917 (N_4917,N_1400,N_186);
nor U4918 (N_4918,N_250,N_1327);
nand U4919 (N_4919,N_2552,N_1195);
nor U4920 (N_4920,N_203,N_1057);
nand U4921 (N_4921,N_2134,N_1826);
or U4922 (N_4922,N_2598,N_2538);
xnor U4923 (N_4923,N_2904,N_926);
xor U4924 (N_4924,N_1014,N_192);
xnor U4925 (N_4925,N_2215,N_1027);
nor U4926 (N_4926,N_2590,N_2965);
xor U4927 (N_4927,N_2668,N_2520);
and U4928 (N_4928,N_2782,N_2499);
nand U4929 (N_4929,N_1146,N_2702);
xor U4930 (N_4930,N_1494,N_1634);
nand U4931 (N_4931,N_1229,N_2862);
nand U4932 (N_4932,N_1934,N_983);
xnor U4933 (N_4933,N_1034,N_1893);
xor U4934 (N_4934,N_2468,N_1697);
nor U4935 (N_4935,N_381,N_2099);
and U4936 (N_4936,N_1485,N_2103);
nor U4937 (N_4937,N_2860,N_1224);
and U4938 (N_4938,N_2038,N_1747);
xnor U4939 (N_4939,N_1306,N_2202);
xnor U4940 (N_4940,N_2176,N_2814);
nor U4941 (N_4941,N_1475,N_2313);
or U4942 (N_4942,N_177,N_1611);
xnor U4943 (N_4943,N_50,N_1682);
nand U4944 (N_4944,N_1633,N_113);
nand U4945 (N_4945,N_1636,N_920);
nand U4946 (N_4946,N_580,N_1433);
nand U4947 (N_4947,N_2705,N_2580);
or U4948 (N_4948,N_1756,N_2498);
xnor U4949 (N_4949,N_751,N_2831);
xor U4950 (N_4950,N_289,N_941);
and U4951 (N_4951,N_289,N_2124);
nand U4952 (N_4952,N_1368,N_2711);
or U4953 (N_4953,N_1838,N_1371);
xnor U4954 (N_4954,N_19,N_1530);
and U4955 (N_4955,N_1641,N_552);
or U4956 (N_4956,N_2597,N_1137);
xor U4957 (N_4957,N_1382,N_2676);
nand U4958 (N_4958,N_1241,N_2770);
xnor U4959 (N_4959,N_1210,N_2862);
or U4960 (N_4960,N_710,N_722);
xor U4961 (N_4961,N_288,N_506);
and U4962 (N_4962,N_2694,N_850);
xnor U4963 (N_4963,N_2993,N_2201);
xnor U4964 (N_4964,N_1239,N_1917);
nand U4965 (N_4965,N_80,N_1718);
and U4966 (N_4966,N_2605,N_1131);
and U4967 (N_4967,N_794,N_835);
nor U4968 (N_4968,N_1690,N_279);
xor U4969 (N_4969,N_2704,N_1731);
or U4970 (N_4970,N_656,N_1822);
nor U4971 (N_4971,N_1232,N_2039);
and U4972 (N_4972,N_2333,N_62);
or U4973 (N_4973,N_736,N_2604);
nand U4974 (N_4974,N_2339,N_1790);
nor U4975 (N_4975,N_2082,N_2539);
nor U4976 (N_4976,N_1515,N_608);
nand U4977 (N_4977,N_672,N_1397);
and U4978 (N_4978,N_1244,N_1650);
xor U4979 (N_4979,N_1419,N_2870);
nor U4980 (N_4980,N_2278,N_1024);
or U4981 (N_4981,N_1985,N_2296);
nand U4982 (N_4982,N_2067,N_924);
nand U4983 (N_4983,N_370,N_377);
and U4984 (N_4984,N_1769,N_2495);
nor U4985 (N_4985,N_1766,N_2321);
nor U4986 (N_4986,N_262,N_812);
xnor U4987 (N_4987,N_1562,N_2001);
and U4988 (N_4988,N_107,N_1036);
nor U4989 (N_4989,N_1056,N_2978);
nand U4990 (N_4990,N_742,N_2908);
nand U4991 (N_4991,N_1914,N_2524);
nand U4992 (N_4992,N_1115,N_2884);
xor U4993 (N_4993,N_2353,N_2506);
nand U4994 (N_4994,N_276,N_61);
nor U4995 (N_4995,N_1298,N_863);
xnor U4996 (N_4996,N_235,N_2782);
or U4997 (N_4997,N_2670,N_2605);
xor U4998 (N_4998,N_2593,N_2413);
xor U4999 (N_4999,N_2562,N_2977);
xnor U5000 (N_5000,N_1046,N_445);
nand U5001 (N_5001,N_544,N_2508);
and U5002 (N_5002,N_2973,N_2021);
nand U5003 (N_5003,N_348,N_1171);
nor U5004 (N_5004,N_1707,N_2143);
and U5005 (N_5005,N_1602,N_1351);
and U5006 (N_5006,N_817,N_1805);
or U5007 (N_5007,N_2640,N_1072);
and U5008 (N_5008,N_1550,N_736);
xnor U5009 (N_5009,N_1529,N_2184);
and U5010 (N_5010,N_2822,N_2646);
or U5011 (N_5011,N_2755,N_2478);
or U5012 (N_5012,N_786,N_2911);
nand U5013 (N_5013,N_1501,N_2982);
xnor U5014 (N_5014,N_2764,N_1976);
nand U5015 (N_5015,N_2603,N_2755);
nor U5016 (N_5016,N_151,N_165);
nor U5017 (N_5017,N_2968,N_1217);
nand U5018 (N_5018,N_669,N_708);
or U5019 (N_5019,N_1463,N_466);
nand U5020 (N_5020,N_2720,N_906);
xor U5021 (N_5021,N_1427,N_1223);
nor U5022 (N_5022,N_1560,N_357);
and U5023 (N_5023,N_1321,N_253);
or U5024 (N_5024,N_1294,N_2599);
or U5025 (N_5025,N_419,N_1060);
or U5026 (N_5026,N_103,N_739);
nand U5027 (N_5027,N_2649,N_2825);
nor U5028 (N_5028,N_646,N_2701);
or U5029 (N_5029,N_2365,N_372);
nand U5030 (N_5030,N_1711,N_2074);
nor U5031 (N_5031,N_2761,N_2311);
nand U5032 (N_5032,N_208,N_504);
nor U5033 (N_5033,N_669,N_2851);
nor U5034 (N_5034,N_1219,N_2915);
nor U5035 (N_5035,N_527,N_1479);
xnor U5036 (N_5036,N_2525,N_2011);
nor U5037 (N_5037,N_1849,N_354);
xnor U5038 (N_5038,N_2101,N_662);
or U5039 (N_5039,N_1205,N_1953);
nor U5040 (N_5040,N_1276,N_1970);
and U5041 (N_5041,N_490,N_1801);
nand U5042 (N_5042,N_1111,N_1476);
nand U5043 (N_5043,N_807,N_839);
nor U5044 (N_5044,N_2086,N_2359);
nand U5045 (N_5045,N_188,N_1554);
and U5046 (N_5046,N_570,N_2011);
and U5047 (N_5047,N_1506,N_1539);
and U5048 (N_5048,N_2240,N_2031);
or U5049 (N_5049,N_476,N_254);
xor U5050 (N_5050,N_1911,N_2107);
or U5051 (N_5051,N_705,N_1958);
or U5052 (N_5052,N_1947,N_2255);
nor U5053 (N_5053,N_1219,N_1718);
xor U5054 (N_5054,N_737,N_277);
or U5055 (N_5055,N_2993,N_1817);
nand U5056 (N_5056,N_1696,N_824);
nand U5057 (N_5057,N_1394,N_327);
or U5058 (N_5058,N_2597,N_991);
or U5059 (N_5059,N_110,N_2696);
or U5060 (N_5060,N_2933,N_1263);
xor U5061 (N_5061,N_1900,N_1824);
nand U5062 (N_5062,N_1852,N_1911);
and U5063 (N_5063,N_1183,N_1973);
and U5064 (N_5064,N_1493,N_2458);
nor U5065 (N_5065,N_1721,N_841);
or U5066 (N_5066,N_1871,N_971);
nand U5067 (N_5067,N_2174,N_1700);
and U5068 (N_5068,N_2315,N_1087);
xnor U5069 (N_5069,N_1678,N_1139);
and U5070 (N_5070,N_2623,N_1393);
xor U5071 (N_5071,N_2725,N_2778);
or U5072 (N_5072,N_1427,N_1064);
nand U5073 (N_5073,N_536,N_2925);
and U5074 (N_5074,N_1755,N_1451);
and U5075 (N_5075,N_542,N_1381);
xor U5076 (N_5076,N_2899,N_796);
nor U5077 (N_5077,N_1173,N_555);
xor U5078 (N_5078,N_1215,N_2168);
nor U5079 (N_5079,N_1821,N_1373);
or U5080 (N_5080,N_2084,N_1387);
xor U5081 (N_5081,N_1824,N_466);
nor U5082 (N_5082,N_1418,N_2128);
nand U5083 (N_5083,N_715,N_1301);
nand U5084 (N_5084,N_374,N_762);
and U5085 (N_5085,N_1055,N_2694);
xnor U5086 (N_5086,N_497,N_929);
xor U5087 (N_5087,N_1152,N_2448);
nor U5088 (N_5088,N_2922,N_2581);
or U5089 (N_5089,N_31,N_58);
nand U5090 (N_5090,N_1417,N_541);
or U5091 (N_5091,N_416,N_1492);
nor U5092 (N_5092,N_2569,N_817);
and U5093 (N_5093,N_2982,N_1288);
or U5094 (N_5094,N_907,N_148);
and U5095 (N_5095,N_1170,N_273);
nand U5096 (N_5096,N_2808,N_1701);
and U5097 (N_5097,N_1060,N_1050);
nor U5098 (N_5098,N_804,N_2631);
nand U5099 (N_5099,N_10,N_2393);
xor U5100 (N_5100,N_1417,N_582);
nor U5101 (N_5101,N_2070,N_392);
nand U5102 (N_5102,N_376,N_2792);
and U5103 (N_5103,N_1666,N_2796);
or U5104 (N_5104,N_626,N_2146);
or U5105 (N_5105,N_260,N_235);
and U5106 (N_5106,N_932,N_2934);
xnor U5107 (N_5107,N_1227,N_1469);
nand U5108 (N_5108,N_1825,N_2726);
nor U5109 (N_5109,N_770,N_2041);
and U5110 (N_5110,N_1655,N_225);
nor U5111 (N_5111,N_1884,N_275);
nand U5112 (N_5112,N_1174,N_1797);
xor U5113 (N_5113,N_1247,N_1334);
or U5114 (N_5114,N_749,N_2821);
or U5115 (N_5115,N_2622,N_2009);
xor U5116 (N_5116,N_2157,N_1525);
or U5117 (N_5117,N_731,N_321);
xor U5118 (N_5118,N_142,N_512);
or U5119 (N_5119,N_623,N_1020);
nor U5120 (N_5120,N_357,N_100);
xnor U5121 (N_5121,N_215,N_2603);
nand U5122 (N_5122,N_2880,N_1657);
xor U5123 (N_5123,N_968,N_1920);
or U5124 (N_5124,N_1003,N_1319);
nand U5125 (N_5125,N_1240,N_1665);
and U5126 (N_5126,N_99,N_1690);
nand U5127 (N_5127,N_852,N_72);
and U5128 (N_5128,N_976,N_614);
and U5129 (N_5129,N_2117,N_1356);
nand U5130 (N_5130,N_2142,N_2841);
nand U5131 (N_5131,N_1843,N_199);
nand U5132 (N_5132,N_2428,N_1477);
xnor U5133 (N_5133,N_2904,N_1095);
and U5134 (N_5134,N_1762,N_2708);
or U5135 (N_5135,N_250,N_481);
and U5136 (N_5136,N_185,N_1977);
nand U5137 (N_5137,N_2483,N_2266);
xor U5138 (N_5138,N_751,N_1873);
xor U5139 (N_5139,N_844,N_172);
nor U5140 (N_5140,N_212,N_1553);
and U5141 (N_5141,N_1425,N_650);
xnor U5142 (N_5142,N_1796,N_1086);
nand U5143 (N_5143,N_600,N_2885);
xnor U5144 (N_5144,N_1612,N_2571);
and U5145 (N_5145,N_2921,N_1012);
nand U5146 (N_5146,N_1575,N_1521);
nand U5147 (N_5147,N_1689,N_1703);
nor U5148 (N_5148,N_1755,N_734);
and U5149 (N_5149,N_2959,N_809);
and U5150 (N_5150,N_2214,N_1181);
xnor U5151 (N_5151,N_862,N_2582);
and U5152 (N_5152,N_2726,N_388);
and U5153 (N_5153,N_2998,N_1727);
nand U5154 (N_5154,N_2032,N_271);
nand U5155 (N_5155,N_2949,N_915);
nor U5156 (N_5156,N_468,N_1427);
nor U5157 (N_5157,N_2094,N_2089);
or U5158 (N_5158,N_637,N_1089);
nor U5159 (N_5159,N_1843,N_2879);
xnor U5160 (N_5160,N_2086,N_1897);
nand U5161 (N_5161,N_2755,N_2677);
nor U5162 (N_5162,N_1019,N_376);
or U5163 (N_5163,N_2635,N_2506);
or U5164 (N_5164,N_498,N_146);
nand U5165 (N_5165,N_2087,N_1815);
xnor U5166 (N_5166,N_1313,N_2202);
and U5167 (N_5167,N_96,N_393);
and U5168 (N_5168,N_315,N_1664);
and U5169 (N_5169,N_1483,N_1642);
nor U5170 (N_5170,N_2566,N_64);
nor U5171 (N_5171,N_40,N_1230);
nand U5172 (N_5172,N_1021,N_1791);
and U5173 (N_5173,N_706,N_2841);
nor U5174 (N_5174,N_1476,N_275);
nand U5175 (N_5175,N_622,N_1569);
nand U5176 (N_5176,N_59,N_1373);
nand U5177 (N_5177,N_2884,N_490);
nand U5178 (N_5178,N_406,N_1943);
xnor U5179 (N_5179,N_2356,N_1085);
or U5180 (N_5180,N_699,N_1091);
nor U5181 (N_5181,N_2442,N_1842);
xor U5182 (N_5182,N_2233,N_206);
and U5183 (N_5183,N_583,N_2710);
and U5184 (N_5184,N_25,N_909);
xor U5185 (N_5185,N_2644,N_934);
or U5186 (N_5186,N_885,N_1119);
nor U5187 (N_5187,N_144,N_2183);
nor U5188 (N_5188,N_2562,N_2556);
and U5189 (N_5189,N_96,N_2533);
or U5190 (N_5190,N_814,N_2861);
and U5191 (N_5191,N_502,N_1128);
and U5192 (N_5192,N_1741,N_2350);
xor U5193 (N_5193,N_2156,N_2809);
xor U5194 (N_5194,N_1981,N_1419);
and U5195 (N_5195,N_2705,N_2999);
nand U5196 (N_5196,N_2641,N_629);
and U5197 (N_5197,N_154,N_2918);
nor U5198 (N_5198,N_1917,N_1189);
xnor U5199 (N_5199,N_1196,N_211);
and U5200 (N_5200,N_793,N_1588);
nor U5201 (N_5201,N_518,N_890);
and U5202 (N_5202,N_1888,N_2214);
or U5203 (N_5203,N_1982,N_1525);
nand U5204 (N_5204,N_132,N_1355);
and U5205 (N_5205,N_1375,N_10);
or U5206 (N_5206,N_1036,N_1100);
xor U5207 (N_5207,N_2889,N_1512);
xor U5208 (N_5208,N_1743,N_2302);
xor U5209 (N_5209,N_2079,N_257);
nand U5210 (N_5210,N_1758,N_854);
nor U5211 (N_5211,N_1213,N_934);
and U5212 (N_5212,N_229,N_2993);
and U5213 (N_5213,N_2028,N_2025);
xnor U5214 (N_5214,N_387,N_473);
nor U5215 (N_5215,N_274,N_2097);
and U5216 (N_5216,N_2195,N_217);
nand U5217 (N_5217,N_736,N_790);
xnor U5218 (N_5218,N_2791,N_721);
nand U5219 (N_5219,N_2766,N_2878);
or U5220 (N_5220,N_2453,N_308);
and U5221 (N_5221,N_883,N_2171);
nor U5222 (N_5222,N_1522,N_1314);
or U5223 (N_5223,N_190,N_2747);
nand U5224 (N_5224,N_2533,N_1995);
or U5225 (N_5225,N_2325,N_1728);
xor U5226 (N_5226,N_1034,N_1232);
and U5227 (N_5227,N_891,N_1993);
xnor U5228 (N_5228,N_2137,N_2729);
xor U5229 (N_5229,N_59,N_2450);
xnor U5230 (N_5230,N_394,N_818);
nor U5231 (N_5231,N_1597,N_696);
or U5232 (N_5232,N_2121,N_1924);
or U5233 (N_5233,N_1732,N_527);
xnor U5234 (N_5234,N_2864,N_1684);
nand U5235 (N_5235,N_263,N_1978);
or U5236 (N_5236,N_1087,N_1356);
and U5237 (N_5237,N_760,N_1256);
nor U5238 (N_5238,N_2056,N_2020);
nor U5239 (N_5239,N_362,N_2302);
nand U5240 (N_5240,N_1081,N_2433);
or U5241 (N_5241,N_2961,N_2693);
or U5242 (N_5242,N_2128,N_1014);
or U5243 (N_5243,N_2930,N_2775);
xor U5244 (N_5244,N_2124,N_1320);
nor U5245 (N_5245,N_67,N_538);
or U5246 (N_5246,N_1400,N_2281);
xor U5247 (N_5247,N_93,N_152);
or U5248 (N_5248,N_1427,N_1447);
nor U5249 (N_5249,N_2065,N_682);
nand U5250 (N_5250,N_2133,N_1575);
nand U5251 (N_5251,N_1261,N_583);
or U5252 (N_5252,N_712,N_1432);
xnor U5253 (N_5253,N_1840,N_2248);
or U5254 (N_5254,N_669,N_214);
xor U5255 (N_5255,N_1064,N_949);
nor U5256 (N_5256,N_2772,N_1459);
xnor U5257 (N_5257,N_1365,N_2166);
xor U5258 (N_5258,N_700,N_592);
and U5259 (N_5259,N_1033,N_405);
or U5260 (N_5260,N_2278,N_1166);
and U5261 (N_5261,N_1152,N_1885);
or U5262 (N_5262,N_1687,N_1104);
nor U5263 (N_5263,N_2037,N_1973);
nand U5264 (N_5264,N_2407,N_1083);
and U5265 (N_5265,N_858,N_2417);
and U5266 (N_5266,N_1383,N_2657);
nand U5267 (N_5267,N_226,N_940);
or U5268 (N_5268,N_540,N_1461);
or U5269 (N_5269,N_2916,N_378);
nor U5270 (N_5270,N_657,N_207);
xnor U5271 (N_5271,N_1157,N_1701);
or U5272 (N_5272,N_1880,N_2553);
nor U5273 (N_5273,N_1640,N_2353);
nor U5274 (N_5274,N_1286,N_358);
nor U5275 (N_5275,N_2797,N_2037);
nand U5276 (N_5276,N_1318,N_654);
xnor U5277 (N_5277,N_241,N_2750);
xor U5278 (N_5278,N_2628,N_1357);
or U5279 (N_5279,N_1692,N_2910);
and U5280 (N_5280,N_1507,N_889);
nand U5281 (N_5281,N_1091,N_1935);
nor U5282 (N_5282,N_2281,N_1215);
nor U5283 (N_5283,N_2503,N_2154);
nand U5284 (N_5284,N_1901,N_484);
nand U5285 (N_5285,N_688,N_330);
xor U5286 (N_5286,N_715,N_1507);
xnor U5287 (N_5287,N_1197,N_1384);
and U5288 (N_5288,N_603,N_1091);
or U5289 (N_5289,N_1274,N_1127);
and U5290 (N_5290,N_1798,N_2135);
or U5291 (N_5291,N_1486,N_109);
xor U5292 (N_5292,N_1480,N_2361);
or U5293 (N_5293,N_1781,N_2415);
nor U5294 (N_5294,N_2176,N_698);
and U5295 (N_5295,N_2369,N_1957);
nor U5296 (N_5296,N_2714,N_1975);
nand U5297 (N_5297,N_2798,N_2744);
and U5298 (N_5298,N_1026,N_1890);
or U5299 (N_5299,N_1503,N_1858);
xor U5300 (N_5300,N_1690,N_264);
or U5301 (N_5301,N_553,N_1773);
nor U5302 (N_5302,N_1393,N_613);
nand U5303 (N_5303,N_1570,N_2920);
or U5304 (N_5304,N_1159,N_2602);
nand U5305 (N_5305,N_212,N_496);
xnor U5306 (N_5306,N_1798,N_1092);
and U5307 (N_5307,N_1518,N_402);
and U5308 (N_5308,N_541,N_1256);
or U5309 (N_5309,N_186,N_653);
nor U5310 (N_5310,N_333,N_22);
xor U5311 (N_5311,N_420,N_765);
nor U5312 (N_5312,N_2517,N_1860);
and U5313 (N_5313,N_2463,N_1277);
or U5314 (N_5314,N_900,N_1762);
and U5315 (N_5315,N_1425,N_1727);
nor U5316 (N_5316,N_1643,N_1823);
or U5317 (N_5317,N_2420,N_125);
nand U5318 (N_5318,N_462,N_981);
nor U5319 (N_5319,N_565,N_807);
nor U5320 (N_5320,N_1510,N_2841);
nand U5321 (N_5321,N_981,N_2663);
or U5322 (N_5322,N_1690,N_1456);
and U5323 (N_5323,N_1283,N_1867);
and U5324 (N_5324,N_267,N_949);
nor U5325 (N_5325,N_2710,N_935);
nand U5326 (N_5326,N_562,N_2177);
xnor U5327 (N_5327,N_2681,N_267);
or U5328 (N_5328,N_1150,N_2565);
and U5329 (N_5329,N_1,N_1065);
or U5330 (N_5330,N_825,N_2046);
nand U5331 (N_5331,N_1777,N_2517);
nand U5332 (N_5332,N_46,N_1404);
and U5333 (N_5333,N_1772,N_2269);
xor U5334 (N_5334,N_2785,N_2864);
nand U5335 (N_5335,N_898,N_2726);
and U5336 (N_5336,N_372,N_1648);
nor U5337 (N_5337,N_797,N_1484);
nand U5338 (N_5338,N_2557,N_418);
or U5339 (N_5339,N_1372,N_2156);
and U5340 (N_5340,N_458,N_1773);
xor U5341 (N_5341,N_2546,N_1138);
or U5342 (N_5342,N_2603,N_1102);
or U5343 (N_5343,N_2584,N_2147);
and U5344 (N_5344,N_680,N_2848);
nand U5345 (N_5345,N_495,N_2393);
and U5346 (N_5346,N_748,N_177);
nor U5347 (N_5347,N_860,N_2388);
or U5348 (N_5348,N_520,N_483);
nand U5349 (N_5349,N_1762,N_1456);
nor U5350 (N_5350,N_2953,N_2513);
xnor U5351 (N_5351,N_1621,N_279);
xor U5352 (N_5352,N_2696,N_1897);
xnor U5353 (N_5353,N_555,N_557);
xnor U5354 (N_5354,N_2908,N_299);
nand U5355 (N_5355,N_2060,N_645);
or U5356 (N_5356,N_1740,N_1367);
nand U5357 (N_5357,N_746,N_701);
xor U5358 (N_5358,N_1708,N_1652);
xnor U5359 (N_5359,N_2840,N_308);
xnor U5360 (N_5360,N_995,N_577);
and U5361 (N_5361,N_1263,N_712);
nand U5362 (N_5362,N_2949,N_2988);
xnor U5363 (N_5363,N_2126,N_875);
or U5364 (N_5364,N_2613,N_1199);
or U5365 (N_5365,N_1073,N_534);
nand U5366 (N_5366,N_1724,N_2352);
and U5367 (N_5367,N_377,N_62);
nor U5368 (N_5368,N_2007,N_466);
nor U5369 (N_5369,N_323,N_939);
nand U5370 (N_5370,N_1947,N_1984);
or U5371 (N_5371,N_1035,N_613);
or U5372 (N_5372,N_846,N_396);
nand U5373 (N_5373,N_2813,N_115);
nand U5374 (N_5374,N_638,N_2095);
and U5375 (N_5375,N_2370,N_2389);
nand U5376 (N_5376,N_84,N_930);
nand U5377 (N_5377,N_470,N_2120);
and U5378 (N_5378,N_2417,N_733);
xnor U5379 (N_5379,N_1385,N_1074);
xor U5380 (N_5380,N_471,N_1791);
nor U5381 (N_5381,N_1115,N_415);
nand U5382 (N_5382,N_824,N_981);
and U5383 (N_5383,N_662,N_209);
nor U5384 (N_5384,N_1154,N_1653);
xnor U5385 (N_5385,N_1013,N_1527);
nor U5386 (N_5386,N_2393,N_2960);
or U5387 (N_5387,N_2784,N_19);
xnor U5388 (N_5388,N_740,N_1193);
and U5389 (N_5389,N_456,N_369);
and U5390 (N_5390,N_2390,N_954);
nand U5391 (N_5391,N_1931,N_2336);
and U5392 (N_5392,N_2406,N_876);
and U5393 (N_5393,N_1429,N_2944);
nand U5394 (N_5394,N_287,N_1498);
and U5395 (N_5395,N_2338,N_1389);
nor U5396 (N_5396,N_1572,N_2937);
and U5397 (N_5397,N_1868,N_1307);
nor U5398 (N_5398,N_347,N_501);
nand U5399 (N_5399,N_85,N_685);
nand U5400 (N_5400,N_935,N_371);
nor U5401 (N_5401,N_179,N_1574);
nand U5402 (N_5402,N_2771,N_1396);
nand U5403 (N_5403,N_846,N_2086);
xor U5404 (N_5404,N_2571,N_804);
or U5405 (N_5405,N_926,N_398);
nor U5406 (N_5406,N_1037,N_415);
or U5407 (N_5407,N_1495,N_1558);
and U5408 (N_5408,N_2928,N_2915);
and U5409 (N_5409,N_2637,N_600);
nor U5410 (N_5410,N_485,N_1916);
nor U5411 (N_5411,N_1758,N_1144);
nor U5412 (N_5412,N_2380,N_1376);
nand U5413 (N_5413,N_2537,N_2473);
and U5414 (N_5414,N_1658,N_2822);
nand U5415 (N_5415,N_2201,N_2228);
and U5416 (N_5416,N_1731,N_1923);
or U5417 (N_5417,N_2962,N_1766);
nor U5418 (N_5418,N_2359,N_793);
nor U5419 (N_5419,N_1078,N_2457);
nor U5420 (N_5420,N_893,N_2474);
nand U5421 (N_5421,N_685,N_1446);
nand U5422 (N_5422,N_2859,N_1540);
nand U5423 (N_5423,N_442,N_1085);
and U5424 (N_5424,N_289,N_1595);
xor U5425 (N_5425,N_1673,N_2349);
or U5426 (N_5426,N_2567,N_1695);
xnor U5427 (N_5427,N_591,N_1533);
and U5428 (N_5428,N_404,N_12);
or U5429 (N_5429,N_2901,N_141);
nor U5430 (N_5430,N_2377,N_313);
nand U5431 (N_5431,N_917,N_2682);
nor U5432 (N_5432,N_2560,N_2974);
nand U5433 (N_5433,N_1183,N_2929);
xnor U5434 (N_5434,N_2398,N_907);
and U5435 (N_5435,N_2856,N_1332);
xnor U5436 (N_5436,N_2670,N_64);
and U5437 (N_5437,N_1912,N_2618);
nand U5438 (N_5438,N_1604,N_2255);
nand U5439 (N_5439,N_1383,N_550);
nand U5440 (N_5440,N_2264,N_227);
or U5441 (N_5441,N_1179,N_38);
nand U5442 (N_5442,N_1075,N_2784);
or U5443 (N_5443,N_1906,N_1087);
nand U5444 (N_5444,N_1520,N_2118);
nor U5445 (N_5445,N_818,N_985);
and U5446 (N_5446,N_2128,N_1781);
or U5447 (N_5447,N_918,N_553);
or U5448 (N_5448,N_436,N_1541);
xor U5449 (N_5449,N_84,N_1507);
xnor U5450 (N_5450,N_552,N_1509);
or U5451 (N_5451,N_828,N_1797);
xor U5452 (N_5452,N_2190,N_694);
nand U5453 (N_5453,N_2625,N_604);
and U5454 (N_5454,N_2972,N_2607);
or U5455 (N_5455,N_1196,N_2760);
nand U5456 (N_5456,N_19,N_1739);
nor U5457 (N_5457,N_1829,N_2734);
and U5458 (N_5458,N_1061,N_2351);
xnor U5459 (N_5459,N_1285,N_1117);
nand U5460 (N_5460,N_424,N_1072);
or U5461 (N_5461,N_837,N_1838);
or U5462 (N_5462,N_1145,N_1887);
nor U5463 (N_5463,N_1180,N_2075);
nor U5464 (N_5464,N_1976,N_2459);
or U5465 (N_5465,N_863,N_570);
xor U5466 (N_5466,N_588,N_73);
xnor U5467 (N_5467,N_362,N_613);
nor U5468 (N_5468,N_723,N_2776);
nor U5469 (N_5469,N_2027,N_2334);
and U5470 (N_5470,N_1969,N_2010);
xnor U5471 (N_5471,N_1416,N_1021);
or U5472 (N_5472,N_1733,N_2092);
nand U5473 (N_5473,N_1409,N_1004);
and U5474 (N_5474,N_816,N_215);
and U5475 (N_5475,N_1851,N_2156);
xnor U5476 (N_5476,N_1651,N_333);
or U5477 (N_5477,N_169,N_92);
nor U5478 (N_5478,N_2101,N_2217);
xnor U5479 (N_5479,N_537,N_2469);
xor U5480 (N_5480,N_863,N_329);
or U5481 (N_5481,N_1921,N_1418);
and U5482 (N_5482,N_1874,N_453);
nand U5483 (N_5483,N_478,N_19);
nand U5484 (N_5484,N_2891,N_1572);
and U5485 (N_5485,N_403,N_677);
xnor U5486 (N_5486,N_94,N_2070);
and U5487 (N_5487,N_1286,N_2721);
nand U5488 (N_5488,N_1265,N_318);
and U5489 (N_5489,N_1554,N_946);
nand U5490 (N_5490,N_1648,N_2360);
or U5491 (N_5491,N_893,N_926);
nand U5492 (N_5492,N_591,N_724);
or U5493 (N_5493,N_279,N_520);
and U5494 (N_5494,N_1325,N_2230);
nor U5495 (N_5495,N_2362,N_309);
xor U5496 (N_5496,N_744,N_2971);
nand U5497 (N_5497,N_2375,N_109);
and U5498 (N_5498,N_2838,N_1518);
nor U5499 (N_5499,N_85,N_2589);
xor U5500 (N_5500,N_1536,N_1253);
or U5501 (N_5501,N_1396,N_2973);
and U5502 (N_5502,N_2029,N_2958);
nand U5503 (N_5503,N_2861,N_2798);
xor U5504 (N_5504,N_533,N_52);
nor U5505 (N_5505,N_2998,N_2001);
nand U5506 (N_5506,N_1288,N_2111);
xnor U5507 (N_5507,N_840,N_2304);
xor U5508 (N_5508,N_1580,N_244);
nand U5509 (N_5509,N_769,N_385);
nor U5510 (N_5510,N_2795,N_2385);
nand U5511 (N_5511,N_2811,N_2085);
nor U5512 (N_5512,N_2294,N_1227);
xor U5513 (N_5513,N_2718,N_2885);
nor U5514 (N_5514,N_259,N_126);
nand U5515 (N_5515,N_2922,N_2373);
nand U5516 (N_5516,N_1346,N_1288);
nand U5517 (N_5517,N_1244,N_1871);
and U5518 (N_5518,N_1122,N_2600);
nor U5519 (N_5519,N_2977,N_1001);
nand U5520 (N_5520,N_2723,N_1879);
or U5521 (N_5521,N_2580,N_583);
nand U5522 (N_5522,N_1942,N_312);
nor U5523 (N_5523,N_2866,N_1485);
nand U5524 (N_5524,N_573,N_2274);
or U5525 (N_5525,N_765,N_277);
or U5526 (N_5526,N_1639,N_142);
xor U5527 (N_5527,N_436,N_917);
or U5528 (N_5528,N_2026,N_896);
xor U5529 (N_5529,N_735,N_68);
xor U5530 (N_5530,N_921,N_100);
xnor U5531 (N_5531,N_2443,N_195);
nand U5532 (N_5532,N_1159,N_2670);
xor U5533 (N_5533,N_2962,N_24);
nor U5534 (N_5534,N_814,N_2260);
nor U5535 (N_5535,N_1,N_500);
xnor U5536 (N_5536,N_654,N_2625);
xor U5537 (N_5537,N_992,N_2844);
or U5538 (N_5538,N_2266,N_1406);
nor U5539 (N_5539,N_8,N_822);
nand U5540 (N_5540,N_460,N_2967);
xnor U5541 (N_5541,N_318,N_2622);
xnor U5542 (N_5542,N_1695,N_2501);
nor U5543 (N_5543,N_761,N_290);
nand U5544 (N_5544,N_1707,N_1459);
nand U5545 (N_5545,N_1605,N_1999);
or U5546 (N_5546,N_1482,N_1148);
and U5547 (N_5547,N_1233,N_2931);
and U5548 (N_5548,N_71,N_333);
xnor U5549 (N_5549,N_1426,N_358);
and U5550 (N_5550,N_2315,N_2704);
xnor U5551 (N_5551,N_559,N_719);
nor U5552 (N_5552,N_488,N_2780);
nand U5553 (N_5553,N_1778,N_1920);
and U5554 (N_5554,N_2984,N_1863);
nand U5555 (N_5555,N_1347,N_831);
or U5556 (N_5556,N_2166,N_1346);
nand U5557 (N_5557,N_778,N_1834);
nand U5558 (N_5558,N_1523,N_1354);
nand U5559 (N_5559,N_913,N_436);
nor U5560 (N_5560,N_1875,N_326);
nor U5561 (N_5561,N_2154,N_1029);
xnor U5562 (N_5562,N_878,N_2637);
and U5563 (N_5563,N_174,N_588);
and U5564 (N_5564,N_1611,N_2237);
and U5565 (N_5565,N_1708,N_96);
xnor U5566 (N_5566,N_1542,N_1903);
nor U5567 (N_5567,N_697,N_1885);
and U5568 (N_5568,N_2076,N_373);
nor U5569 (N_5569,N_451,N_1202);
or U5570 (N_5570,N_2059,N_108);
or U5571 (N_5571,N_2510,N_1181);
nand U5572 (N_5572,N_1539,N_2374);
nor U5573 (N_5573,N_1904,N_29);
and U5574 (N_5574,N_575,N_88);
nand U5575 (N_5575,N_2018,N_212);
xor U5576 (N_5576,N_1532,N_2837);
nand U5577 (N_5577,N_1993,N_1298);
nor U5578 (N_5578,N_19,N_682);
nand U5579 (N_5579,N_1538,N_1121);
nor U5580 (N_5580,N_2887,N_2874);
and U5581 (N_5581,N_1780,N_1242);
nand U5582 (N_5582,N_2489,N_1869);
xor U5583 (N_5583,N_1598,N_965);
nor U5584 (N_5584,N_328,N_2002);
nor U5585 (N_5585,N_1157,N_1398);
nand U5586 (N_5586,N_402,N_897);
nor U5587 (N_5587,N_233,N_832);
and U5588 (N_5588,N_100,N_881);
and U5589 (N_5589,N_2768,N_30);
nor U5590 (N_5590,N_2380,N_1151);
nor U5591 (N_5591,N_1483,N_2);
and U5592 (N_5592,N_2597,N_1018);
nand U5593 (N_5593,N_1115,N_1744);
nand U5594 (N_5594,N_1853,N_1871);
and U5595 (N_5595,N_1989,N_515);
nand U5596 (N_5596,N_1936,N_667);
or U5597 (N_5597,N_1759,N_2706);
nand U5598 (N_5598,N_1589,N_2026);
xnor U5599 (N_5599,N_327,N_1619);
or U5600 (N_5600,N_647,N_1324);
nor U5601 (N_5601,N_1723,N_1837);
or U5602 (N_5602,N_145,N_1502);
nand U5603 (N_5603,N_2625,N_1179);
nor U5604 (N_5604,N_174,N_1822);
nand U5605 (N_5605,N_2459,N_2411);
nor U5606 (N_5606,N_996,N_2661);
or U5607 (N_5607,N_2270,N_199);
nand U5608 (N_5608,N_2850,N_506);
or U5609 (N_5609,N_902,N_210);
xor U5610 (N_5610,N_2175,N_2058);
nand U5611 (N_5611,N_2665,N_1256);
nor U5612 (N_5612,N_1043,N_1968);
and U5613 (N_5613,N_404,N_1394);
and U5614 (N_5614,N_1561,N_371);
nor U5615 (N_5615,N_1901,N_2594);
xor U5616 (N_5616,N_1178,N_2983);
nand U5617 (N_5617,N_308,N_1340);
nor U5618 (N_5618,N_2560,N_1517);
or U5619 (N_5619,N_1564,N_650);
and U5620 (N_5620,N_1525,N_43);
and U5621 (N_5621,N_157,N_2948);
nand U5622 (N_5622,N_2006,N_1590);
nand U5623 (N_5623,N_2410,N_1712);
nand U5624 (N_5624,N_693,N_2190);
xnor U5625 (N_5625,N_1465,N_2911);
and U5626 (N_5626,N_1190,N_551);
xnor U5627 (N_5627,N_2618,N_2402);
nor U5628 (N_5628,N_675,N_797);
nand U5629 (N_5629,N_2671,N_2130);
xor U5630 (N_5630,N_281,N_2031);
xnor U5631 (N_5631,N_1039,N_2362);
xnor U5632 (N_5632,N_2594,N_93);
xnor U5633 (N_5633,N_227,N_442);
nand U5634 (N_5634,N_807,N_1598);
nor U5635 (N_5635,N_482,N_1982);
nor U5636 (N_5636,N_737,N_1733);
xnor U5637 (N_5637,N_1446,N_1979);
or U5638 (N_5638,N_924,N_1111);
or U5639 (N_5639,N_886,N_5);
or U5640 (N_5640,N_1923,N_55);
nor U5641 (N_5641,N_2124,N_2100);
nor U5642 (N_5642,N_420,N_1363);
nor U5643 (N_5643,N_2291,N_1339);
xnor U5644 (N_5644,N_2372,N_740);
nand U5645 (N_5645,N_2623,N_1909);
and U5646 (N_5646,N_2798,N_1511);
xor U5647 (N_5647,N_791,N_1987);
or U5648 (N_5648,N_2375,N_2744);
nand U5649 (N_5649,N_61,N_2440);
and U5650 (N_5650,N_858,N_1504);
and U5651 (N_5651,N_1313,N_2025);
or U5652 (N_5652,N_2537,N_2251);
xor U5653 (N_5653,N_2301,N_2440);
nand U5654 (N_5654,N_197,N_2751);
xnor U5655 (N_5655,N_326,N_1091);
or U5656 (N_5656,N_2045,N_2976);
and U5657 (N_5657,N_98,N_1049);
and U5658 (N_5658,N_1561,N_1520);
xor U5659 (N_5659,N_1710,N_2683);
or U5660 (N_5660,N_2191,N_1031);
xor U5661 (N_5661,N_2121,N_597);
nand U5662 (N_5662,N_1978,N_1806);
and U5663 (N_5663,N_1958,N_135);
nor U5664 (N_5664,N_104,N_2128);
and U5665 (N_5665,N_828,N_2046);
and U5666 (N_5666,N_118,N_1056);
nand U5667 (N_5667,N_2553,N_573);
nand U5668 (N_5668,N_2303,N_1830);
nand U5669 (N_5669,N_2090,N_318);
nor U5670 (N_5670,N_2796,N_122);
nand U5671 (N_5671,N_1084,N_380);
nor U5672 (N_5672,N_2745,N_215);
nand U5673 (N_5673,N_50,N_2529);
and U5674 (N_5674,N_2306,N_1310);
nor U5675 (N_5675,N_2505,N_1060);
xnor U5676 (N_5676,N_2854,N_2526);
and U5677 (N_5677,N_120,N_714);
xor U5678 (N_5678,N_2651,N_443);
or U5679 (N_5679,N_1364,N_1294);
and U5680 (N_5680,N_2934,N_72);
or U5681 (N_5681,N_2675,N_1381);
or U5682 (N_5682,N_1100,N_744);
xor U5683 (N_5683,N_2177,N_2652);
nor U5684 (N_5684,N_164,N_1245);
nand U5685 (N_5685,N_1083,N_1593);
nor U5686 (N_5686,N_986,N_555);
and U5687 (N_5687,N_1376,N_2503);
nand U5688 (N_5688,N_2026,N_2331);
nor U5689 (N_5689,N_2049,N_859);
and U5690 (N_5690,N_568,N_2856);
or U5691 (N_5691,N_2864,N_828);
nor U5692 (N_5692,N_489,N_1619);
nand U5693 (N_5693,N_2993,N_1308);
and U5694 (N_5694,N_1069,N_1282);
or U5695 (N_5695,N_2251,N_2534);
or U5696 (N_5696,N_306,N_907);
xnor U5697 (N_5697,N_208,N_55);
nor U5698 (N_5698,N_1690,N_1275);
and U5699 (N_5699,N_402,N_1668);
nand U5700 (N_5700,N_1794,N_619);
nor U5701 (N_5701,N_1444,N_980);
xor U5702 (N_5702,N_1771,N_2616);
nor U5703 (N_5703,N_2898,N_2738);
or U5704 (N_5704,N_1169,N_38);
or U5705 (N_5705,N_557,N_2255);
and U5706 (N_5706,N_2719,N_1251);
xnor U5707 (N_5707,N_2935,N_2225);
xor U5708 (N_5708,N_2097,N_67);
nand U5709 (N_5709,N_617,N_2182);
nand U5710 (N_5710,N_441,N_2163);
nand U5711 (N_5711,N_977,N_223);
and U5712 (N_5712,N_1578,N_824);
or U5713 (N_5713,N_2543,N_523);
and U5714 (N_5714,N_791,N_2977);
or U5715 (N_5715,N_667,N_1947);
nor U5716 (N_5716,N_845,N_184);
nor U5717 (N_5717,N_1022,N_945);
and U5718 (N_5718,N_768,N_909);
nor U5719 (N_5719,N_2573,N_140);
xnor U5720 (N_5720,N_523,N_1363);
xnor U5721 (N_5721,N_1126,N_1875);
xnor U5722 (N_5722,N_2465,N_41);
or U5723 (N_5723,N_181,N_431);
or U5724 (N_5724,N_2957,N_2232);
nand U5725 (N_5725,N_2810,N_2523);
nor U5726 (N_5726,N_2148,N_1234);
nand U5727 (N_5727,N_1147,N_2261);
and U5728 (N_5728,N_2690,N_943);
xor U5729 (N_5729,N_2976,N_921);
nand U5730 (N_5730,N_2190,N_1018);
nand U5731 (N_5731,N_608,N_1173);
nor U5732 (N_5732,N_1039,N_2468);
nor U5733 (N_5733,N_2006,N_2154);
xor U5734 (N_5734,N_2072,N_1102);
nand U5735 (N_5735,N_1847,N_490);
xnor U5736 (N_5736,N_146,N_194);
or U5737 (N_5737,N_1171,N_2520);
or U5738 (N_5738,N_2300,N_2481);
xnor U5739 (N_5739,N_58,N_2450);
nand U5740 (N_5740,N_2629,N_2221);
and U5741 (N_5741,N_335,N_543);
xnor U5742 (N_5742,N_872,N_451);
nor U5743 (N_5743,N_1341,N_887);
or U5744 (N_5744,N_351,N_172);
nor U5745 (N_5745,N_1332,N_812);
nand U5746 (N_5746,N_122,N_1746);
nor U5747 (N_5747,N_2011,N_1643);
nand U5748 (N_5748,N_1371,N_1674);
nand U5749 (N_5749,N_203,N_554);
xor U5750 (N_5750,N_7,N_362);
or U5751 (N_5751,N_2932,N_2807);
and U5752 (N_5752,N_310,N_2759);
and U5753 (N_5753,N_2274,N_2640);
nor U5754 (N_5754,N_1948,N_1326);
xnor U5755 (N_5755,N_699,N_1878);
nor U5756 (N_5756,N_2246,N_1120);
nor U5757 (N_5757,N_2590,N_462);
nor U5758 (N_5758,N_200,N_553);
nand U5759 (N_5759,N_155,N_2696);
nor U5760 (N_5760,N_2729,N_425);
or U5761 (N_5761,N_1641,N_2930);
or U5762 (N_5762,N_620,N_1759);
and U5763 (N_5763,N_2811,N_462);
or U5764 (N_5764,N_1899,N_2670);
nand U5765 (N_5765,N_2149,N_1349);
xor U5766 (N_5766,N_1407,N_2870);
xor U5767 (N_5767,N_2247,N_1846);
nand U5768 (N_5768,N_1549,N_1182);
xnor U5769 (N_5769,N_1650,N_1901);
or U5770 (N_5770,N_2152,N_2735);
or U5771 (N_5771,N_1694,N_37);
nand U5772 (N_5772,N_2661,N_217);
and U5773 (N_5773,N_2744,N_850);
or U5774 (N_5774,N_1309,N_2789);
nor U5775 (N_5775,N_1468,N_1052);
nor U5776 (N_5776,N_376,N_820);
nand U5777 (N_5777,N_1419,N_1077);
nand U5778 (N_5778,N_1493,N_1489);
nand U5779 (N_5779,N_2204,N_1231);
and U5780 (N_5780,N_1113,N_2053);
xor U5781 (N_5781,N_469,N_2642);
nor U5782 (N_5782,N_1883,N_504);
xor U5783 (N_5783,N_425,N_1813);
xnor U5784 (N_5784,N_817,N_2108);
xor U5785 (N_5785,N_292,N_2621);
nor U5786 (N_5786,N_2399,N_1475);
and U5787 (N_5787,N_1126,N_330);
and U5788 (N_5788,N_1729,N_27);
nor U5789 (N_5789,N_1865,N_1716);
nand U5790 (N_5790,N_774,N_2503);
nor U5791 (N_5791,N_2007,N_2517);
xor U5792 (N_5792,N_28,N_1461);
nor U5793 (N_5793,N_590,N_1871);
nand U5794 (N_5794,N_1061,N_415);
nand U5795 (N_5795,N_1718,N_2171);
xor U5796 (N_5796,N_1655,N_1812);
and U5797 (N_5797,N_2740,N_2988);
and U5798 (N_5798,N_2089,N_2997);
or U5799 (N_5799,N_2014,N_2492);
xor U5800 (N_5800,N_2117,N_2742);
xor U5801 (N_5801,N_1275,N_832);
nor U5802 (N_5802,N_994,N_93);
nor U5803 (N_5803,N_1058,N_523);
xnor U5804 (N_5804,N_2404,N_2975);
nor U5805 (N_5805,N_1712,N_1772);
nor U5806 (N_5806,N_1056,N_389);
or U5807 (N_5807,N_1764,N_2);
xnor U5808 (N_5808,N_875,N_1356);
nor U5809 (N_5809,N_149,N_1984);
nand U5810 (N_5810,N_2745,N_447);
and U5811 (N_5811,N_583,N_2756);
or U5812 (N_5812,N_1440,N_1519);
or U5813 (N_5813,N_2234,N_2952);
nor U5814 (N_5814,N_838,N_17);
nor U5815 (N_5815,N_1024,N_2848);
or U5816 (N_5816,N_80,N_2151);
nand U5817 (N_5817,N_2437,N_1257);
and U5818 (N_5818,N_418,N_297);
or U5819 (N_5819,N_2528,N_1343);
nand U5820 (N_5820,N_1746,N_189);
and U5821 (N_5821,N_2348,N_1834);
xnor U5822 (N_5822,N_874,N_165);
xnor U5823 (N_5823,N_1209,N_1793);
nor U5824 (N_5824,N_1140,N_1717);
nand U5825 (N_5825,N_695,N_859);
or U5826 (N_5826,N_1888,N_997);
xnor U5827 (N_5827,N_2925,N_682);
nand U5828 (N_5828,N_1780,N_659);
nand U5829 (N_5829,N_1662,N_2505);
or U5830 (N_5830,N_2800,N_1087);
xnor U5831 (N_5831,N_735,N_1905);
nand U5832 (N_5832,N_1399,N_654);
nand U5833 (N_5833,N_1820,N_2631);
nand U5834 (N_5834,N_1755,N_201);
nor U5835 (N_5835,N_2321,N_2203);
and U5836 (N_5836,N_775,N_67);
nor U5837 (N_5837,N_1389,N_2655);
xnor U5838 (N_5838,N_842,N_1084);
nor U5839 (N_5839,N_327,N_136);
and U5840 (N_5840,N_2549,N_2152);
nand U5841 (N_5841,N_298,N_1649);
nand U5842 (N_5842,N_557,N_907);
or U5843 (N_5843,N_237,N_2004);
nor U5844 (N_5844,N_2696,N_1132);
nor U5845 (N_5845,N_46,N_850);
nor U5846 (N_5846,N_697,N_2836);
nor U5847 (N_5847,N_974,N_673);
nand U5848 (N_5848,N_809,N_1488);
xor U5849 (N_5849,N_2032,N_762);
and U5850 (N_5850,N_247,N_915);
xor U5851 (N_5851,N_1153,N_2009);
and U5852 (N_5852,N_1884,N_588);
or U5853 (N_5853,N_2506,N_2110);
xor U5854 (N_5854,N_1764,N_458);
xnor U5855 (N_5855,N_2877,N_2498);
and U5856 (N_5856,N_1364,N_223);
xor U5857 (N_5857,N_1594,N_2705);
or U5858 (N_5858,N_490,N_647);
xnor U5859 (N_5859,N_793,N_2940);
xnor U5860 (N_5860,N_92,N_1578);
or U5861 (N_5861,N_2794,N_253);
or U5862 (N_5862,N_1007,N_1061);
nand U5863 (N_5863,N_282,N_2372);
and U5864 (N_5864,N_873,N_492);
nand U5865 (N_5865,N_2863,N_1825);
nand U5866 (N_5866,N_865,N_801);
or U5867 (N_5867,N_1006,N_1838);
nand U5868 (N_5868,N_2170,N_2949);
nor U5869 (N_5869,N_2986,N_987);
nand U5870 (N_5870,N_1832,N_2392);
xnor U5871 (N_5871,N_2605,N_901);
xor U5872 (N_5872,N_2981,N_30);
nor U5873 (N_5873,N_2131,N_674);
nor U5874 (N_5874,N_2178,N_2585);
xnor U5875 (N_5875,N_1448,N_1990);
and U5876 (N_5876,N_2362,N_1215);
and U5877 (N_5877,N_2397,N_1673);
nand U5878 (N_5878,N_632,N_1255);
nor U5879 (N_5879,N_904,N_683);
xnor U5880 (N_5880,N_1716,N_2399);
or U5881 (N_5881,N_1457,N_1194);
xnor U5882 (N_5882,N_1096,N_1842);
nand U5883 (N_5883,N_640,N_710);
xor U5884 (N_5884,N_192,N_1886);
nor U5885 (N_5885,N_2586,N_1870);
and U5886 (N_5886,N_1413,N_2661);
nor U5887 (N_5887,N_2607,N_798);
nor U5888 (N_5888,N_1312,N_1132);
nand U5889 (N_5889,N_2807,N_1230);
or U5890 (N_5890,N_2602,N_942);
nor U5891 (N_5891,N_1241,N_207);
nand U5892 (N_5892,N_659,N_2753);
and U5893 (N_5893,N_975,N_2604);
xor U5894 (N_5894,N_1824,N_2817);
or U5895 (N_5895,N_1964,N_524);
nor U5896 (N_5896,N_1111,N_41);
and U5897 (N_5897,N_1971,N_2740);
nor U5898 (N_5898,N_1714,N_466);
nor U5899 (N_5899,N_243,N_1106);
xnor U5900 (N_5900,N_2173,N_2662);
xnor U5901 (N_5901,N_2915,N_2726);
xor U5902 (N_5902,N_129,N_1084);
and U5903 (N_5903,N_1724,N_993);
nor U5904 (N_5904,N_2201,N_899);
and U5905 (N_5905,N_1412,N_1454);
and U5906 (N_5906,N_1123,N_580);
or U5907 (N_5907,N_1365,N_1496);
xor U5908 (N_5908,N_2100,N_759);
or U5909 (N_5909,N_2612,N_1411);
nor U5910 (N_5910,N_2024,N_937);
nor U5911 (N_5911,N_977,N_1588);
xor U5912 (N_5912,N_526,N_793);
and U5913 (N_5913,N_2792,N_1730);
xor U5914 (N_5914,N_1109,N_173);
nand U5915 (N_5915,N_1544,N_1867);
nor U5916 (N_5916,N_1710,N_2629);
nand U5917 (N_5917,N_1435,N_682);
nand U5918 (N_5918,N_32,N_774);
nor U5919 (N_5919,N_293,N_1374);
and U5920 (N_5920,N_2129,N_2426);
or U5921 (N_5921,N_255,N_674);
or U5922 (N_5922,N_2516,N_483);
and U5923 (N_5923,N_2451,N_1893);
xor U5924 (N_5924,N_631,N_1209);
nand U5925 (N_5925,N_1773,N_308);
nor U5926 (N_5926,N_1270,N_420);
and U5927 (N_5927,N_1751,N_2793);
nor U5928 (N_5928,N_2851,N_395);
xnor U5929 (N_5929,N_2806,N_2471);
xor U5930 (N_5930,N_86,N_1725);
xnor U5931 (N_5931,N_840,N_1623);
nand U5932 (N_5932,N_1251,N_2683);
nor U5933 (N_5933,N_2088,N_2449);
and U5934 (N_5934,N_613,N_93);
nand U5935 (N_5935,N_2436,N_2551);
and U5936 (N_5936,N_846,N_1076);
nand U5937 (N_5937,N_590,N_1592);
or U5938 (N_5938,N_1320,N_2988);
nor U5939 (N_5939,N_941,N_1639);
nor U5940 (N_5940,N_377,N_1200);
xnor U5941 (N_5941,N_1990,N_2771);
or U5942 (N_5942,N_824,N_984);
nand U5943 (N_5943,N_908,N_1565);
nor U5944 (N_5944,N_2939,N_1863);
or U5945 (N_5945,N_2341,N_2509);
or U5946 (N_5946,N_2751,N_336);
nor U5947 (N_5947,N_2201,N_1907);
or U5948 (N_5948,N_44,N_2116);
nor U5949 (N_5949,N_1416,N_561);
xnor U5950 (N_5950,N_2264,N_2187);
or U5951 (N_5951,N_907,N_162);
nor U5952 (N_5952,N_1960,N_1961);
nand U5953 (N_5953,N_2749,N_1039);
nor U5954 (N_5954,N_1000,N_1228);
or U5955 (N_5955,N_309,N_143);
nor U5956 (N_5956,N_755,N_1124);
nand U5957 (N_5957,N_2954,N_1805);
nand U5958 (N_5958,N_2921,N_1703);
nor U5959 (N_5959,N_1235,N_2746);
and U5960 (N_5960,N_995,N_2162);
and U5961 (N_5961,N_132,N_2906);
nand U5962 (N_5962,N_234,N_1781);
or U5963 (N_5963,N_697,N_1568);
or U5964 (N_5964,N_2213,N_838);
or U5965 (N_5965,N_2284,N_1093);
nor U5966 (N_5966,N_2169,N_765);
xnor U5967 (N_5967,N_334,N_2486);
or U5968 (N_5968,N_1845,N_663);
or U5969 (N_5969,N_1676,N_2113);
and U5970 (N_5970,N_450,N_1255);
or U5971 (N_5971,N_435,N_2322);
nor U5972 (N_5972,N_2235,N_776);
and U5973 (N_5973,N_1669,N_2506);
nand U5974 (N_5974,N_2182,N_1234);
nor U5975 (N_5975,N_995,N_1202);
nand U5976 (N_5976,N_2682,N_1926);
nand U5977 (N_5977,N_2896,N_2168);
nor U5978 (N_5978,N_1894,N_2959);
xnor U5979 (N_5979,N_2413,N_510);
xnor U5980 (N_5980,N_1512,N_953);
or U5981 (N_5981,N_1574,N_1645);
nor U5982 (N_5982,N_1770,N_1191);
and U5983 (N_5983,N_725,N_2107);
nor U5984 (N_5984,N_1233,N_526);
nor U5985 (N_5985,N_372,N_2073);
xnor U5986 (N_5986,N_2600,N_2013);
and U5987 (N_5987,N_562,N_1769);
and U5988 (N_5988,N_607,N_1174);
or U5989 (N_5989,N_2692,N_358);
nor U5990 (N_5990,N_1333,N_2306);
or U5991 (N_5991,N_1316,N_1419);
or U5992 (N_5992,N_1190,N_234);
or U5993 (N_5993,N_1544,N_1217);
nor U5994 (N_5994,N_1661,N_436);
or U5995 (N_5995,N_2993,N_1082);
nor U5996 (N_5996,N_535,N_846);
and U5997 (N_5997,N_660,N_128);
nand U5998 (N_5998,N_919,N_93);
xor U5999 (N_5999,N_2716,N_302);
and U6000 (N_6000,N_3104,N_3393);
or U6001 (N_6001,N_4614,N_4338);
nor U6002 (N_6002,N_3671,N_3714);
nand U6003 (N_6003,N_4644,N_4224);
nand U6004 (N_6004,N_5401,N_3401);
nor U6005 (N_6005,N_3913,N_4785);
or U6006 (N_6006,N_3835,N_3061);
nor U6007 (N_6007,N_4109,N_4052);
or U6008 (N_6008,N_5131,N_4937);
or U6009 (N_6009,N_3911,N_4226);
or U6010 (N_6010,N_4555,N_4736);
or U6011 (N_6011,N_5929,N_3287);
and U6012 (N_6012,N_4911,N_4135);
or U6013 (N_6013,N_4046,N_4894);
xnor U6014 (N_6014,N_4769,N_3846);
or U6015 (N_6015,N_3149,N_4364);
and U6016 (N_6016,N_3323,N_4340);
nor U6017 (N_6017,N_5258,N_5964);
nand U6018 (N_6018,N_5578,N_5265);
nand U6019 (N_6019,N_4814,N_3662);
nand U6020 (N_6020,N_5823,N_3222);
nor U6021 (N_6021,N_4186,N_5686);
nand U6022 (N_6022,N_4506,N_4815);
nand U6023 (N_6023,N_4885,N_5482);
nor U6024 (N_6024,N_4801,N_3438);
or U6025 (N_6025,N_3439,N_3672);
or U6026 (N_6026,N_5911,N_3436);
nor U6027 (N_6027,N_4328,N_4978);
and U6028 (N_6028,N_4846,N_3334);
nor U6029 (N_6029,N_4444,N_4917);
and U6030 (N_6030,N_5314,N_4180);
nor U6031 (N_6031,N_4366,N_3923);
and U6032 (N_6032,N_4987,N_5642);
nor U6033 (N_6033,N_5245,N_5452);
xor U6034 (N_6034,N_5462,N_3018);
nor U6035 (N_6035,N_5613,N_4933);
nand U6036 (N_6036,N_5368,N_3216);
or U6037 (N_6037,N_3043,N_3109);
xnor U6038 (N_6038,N_5094,N_5114);
nor U6039 (N_6039,N_4733,N_4021);
nor U6040 (N_6040,N_3999,N_5286);
or U6041 (N_6041,N_5869,N_5287);
nor U6042 (N_6042,N_5212,N_3342);
xnor U6043 (N_6043,N_3268,N_3794);
or U6044 (N_6044,N_4268,N_3494);
nor U6045 (N_6045,N_3108,N_4476);
nor U6046 (N_6046,N_3632,N_3220);
and U6047 (N_6047,N_5325,N_5788);
nand U6048 (N_6048,N_5386,N_4207);
or U6049 (N_6049,N_3152,N_3724);
or U6050 (N_6050,N_4966,N_4193);
nand U6051 (N_6051,N_4155,N_5475);
nor U6052 (N_6052,N_3450,N_5033);
nand U6053 (N_6053,N_4333,N_4800);
and U6054 (N_6054,N_5139,N_4386);
and U6055 (N_6055,N_4915,N_4004);
nor U6056 (N_6056,N_4102,N_4250);
and U6057 (N_6057,N_3941,N_4093);
nor U6058 (N_6058,N_4127,N_3987);
nor U6059 (N_6059,N_3803,N_4922);
xnor U6060 (N_6060,N_5144,N_3037);
nor U6061 (N_6061,N_5825,N_3434);
xor U6062 (N_6062,N_3060,N_5075);
and U6063 (N_6063,N_5841,N_3965);
xnor U6064 (N_6064,N_5285,N_5444);
and U6065 (N_6065,N_4148,N_4737);
nor U6066 (N_6066,N_4635,N_3300);
xnor U6067 (N_6067,N_4128,N_5279);
or U6068 (N_6068,N_3716,N_4803);
or U6069 (N_6069,N_4070,N_3319);
xor U6070 (N_6070,N_5012,N_3900);
nand U6071 (N_6071,N_4205,N_4199);
nor U6072 (N_6072,N_3951,N_5090);
or U6073 (N_6073,N_4361,N_4271);
or U6074 (N_6074,N_4988,N_5594);
xor U6075 (N_6075,N_3212,N_4797);
and U6076 (N_6076,N_5775,N_4907);
nand U6077 (N_6077,N_3729,N_4437);
or U6078 (N_6078,N_5554,N_3458);
xor U6079 (N_6079,N_3136,N_5392);
nor U6080 (N_6080,N_4906,N_5540);
or U6081 (N_6081,N_3129,N_3521);
and U6082 (N_6082,N_4173,N_4400);
nor U6083 (N_6083,N_3648,N_4596);
nand U6084 (N_6084,N_4661,N_4358);
nor U6085 (N_6085,N_5189,N_5367);
nand U6086 (N_6086,N_3483,N_3255);
nor U6087 (N_6087,N_3224,N_5629);
nand U6088 (N_6088,N_4347,N_3002);
nand U6089 (N_6089,N_5785,N_5014);
nor U6090 (N_6090,N_4065,N_5845);
nand U6091 (N_6091,N_5416,N_5543);
and U6092 (N_6092,N_4081,N_4951);
nor U6093 (N_6093,N_5732,N_5988);
or U6094 (N_6094,N_3480,N_3301);
nand U6095 (N_6095,N_5501,N_4225);
and U6096 (N_6096,N_4934,N_5373);
xnor U6097 (N_6097,N_4645,N_4646);
nand U6098 (N_6098,N_5087,N_3190);
or U6099 (N_6099,N_4072,N_5609);
or U6100 (N_6100,N_4985,N_4952);
nor U6101 (N_6101,N_4221,N_5125);
or U6102 (N_6102,N_4238,N_5990);
nand U6103 (N_6103,N_4036,N_3554);
or U6104 (N_6104,N_5074,N_3415);
nor U6105 (N_6105,N_5941,N_4055);
or U6106 (N_6106,N_4330,N_5073);
or U6107 (N_6107,N_5730,N_4379);
xnor U6108 (N_6108,N_5611,N_4493);
xor U6109 (N_6109,N_3559,N_5659);
xor U6110 (N_6110,N_4680,N_4022);
or U6111 (N_6111,N_5067,N_5993);
xnor U6112 (N_6112,N_5630,N_5332);
nand U6113 (N_6113,N_3707,N_4816);
nand U6114 (N_6114,N_3605,N_5377);
nand U6115 (N_6115,N_3799,N_3995);
nand U6116 (N_6116,N_3782,N_3591);
or U6117 (N_6117,N_4377,N_4222);
nor U6118 (N_6118,N_3541,N_5565);
nor U6119 (N_6119,N_5644,N_5355);
and U6120 (N_6120,N_3423,N_4606);
and U6121 (N_6121,N_5342,N_4169);
and U6122 (N_6122,N_4416,N_5875);
and U6123 (N_6123,N_3012,N_3683);
nor U6124 (N_6124,N_5602,N_4099);
xnor U6125 (N_6125,N_3501,N_4683);
nand U6126 (N_6126,N_3141,N_4561);
and U6127 (N_6127,N_5161,N_4295);
nor U6128 (N_6128,N_3115,N_5826);
nand U6129 (N_6129,N_3736,N_5983);
xor U6130 (N_6130,N_5351,N_4090);
or U6131 (N_6131,N_3633,N_4182);
xor U6132 (N_6132,N_4475,N_4176);
and U6133 (N_6133,N_4983,N_3909);
nor U6134 (N_6134,N_3918,N_4343);
nand U6135 (N_6135,N_5747,N_4533);
xnor U6136 (N_6136,N_4172,N_3956);
or U6137 (N_6137,N_4527,N_3854);
nor U6138 (N_6138,N_5953,N_3738);
and U6139 (N_6139,N_3041,N_5300);
or U6140 (N_6140,N_5885,N_3841);
xor U6141 (N_6141,N_5054,N_4722);
or U6142 (N_6142,N_4054,N_4075);
xnor U6143 (N_6143,N_5782,N_4768);
nor U6144 (N_6144,N_4033,N_5404);
nand U6145 (N_6145,N_3471,N_4612);
or U6146 (N_6146,N_5205,N_5049);
nor U6147 (N_6147,N_5688,N_5595);
and U6148 (N_6148,N_3540,N_3154);
or U6149 (N_6149,N_3155,N_4152);
xnor U6150 (N_6150,N_3561,N_5772);
xnor U6151 (N_6151,N_5414,N_3784);
and U6152 (N_6152,N_5866,N_3394);
nor U6153 (N_6153,N_5761,N_4433);
or U6154 (N_6154,N_4097,N_4919);
and U6155 (N_6155,N_5844,N_3719);
nand U6156 (N_6156,N_4354,N_4970);
nand U6157 (N_6157,N_5650,N_3908);
nor U6158 (N_6158,N_3964,N_5917);
xnor U6159 (N_6159,N_5066,N_5079);
nor U6160 (N_6160,N_5445,N_4144);
xor U6161 (N_6161,N_5442,N_4427);
or U6162 (N_6162,N_3276,N_3311);
and U6163 (N_6163,N_4827,N_3443);
or U6164 (N_6164,N_4677,N_3919);
nand U6165 (N_6165,N_3040,N_4890);
xor U6166 (N_6166,N_5248,N_5238);
xor U6167 (N_6167,N_5798,N_4590);
nand U6168 (N_6168,N_3055,N_3512);
nor U6169 (N_6169,N_3747,N_4299);
or U6170 (N_6170,N_5320,N_4360);
xor U6171 (N_6171,N_4015,N_4842);
and U6172 (N_6172,N_5583,N_5899);
or U6173 (N_6173,N_5982,N_4651);
or U6174 (N_6174,N_3292,N_5227);
xnor U6175 (N_6175,N_3107,N_3499);
and U6176 (N_6176,N_5330,N_5810);
and U6177 (N_6177,N_4556,N_3444);
or U6178 (N_6178,N_4594,N_3601);
nor U6179 (N_6179,N_4626,N_3432);
xor U6180 (N_6180,N_4957,N_4844);
nand U6181 (N_6181,N_4467,N_4724);
and U6182 (N_6182,N_5834,N_3120);
nand U6183 (N_6183,N_3739,N_4939);
xnor U6184 (N_6184,N_3460,N_4168);
and U6185 (N_6185,N_3976,N_5878);
or U6186 (N_6186,N_3417,N_4552);
nand U6187 (N_6187,N_4613,N_5575);
nor U6188 (N_6188,N_5213,N_5310);
or U6189 (N_6189,N_3031,N_5068);
or U6190 (N_6190,N_5581,N_3510);
nand U6191 (N_6191,N_4992,N_5236);
nand U6192 (N_6192,N_5346,N_4779);
xor U6193 (N_6193,N_4454,N_4248);
or U6194 (N_6194,N_3333,N_5499);
or U6195 (N_6195,N_3685,N_4874);
xor U6196 (N_6196,N_5746,N_4368);
nor U6197 (N_6197,N_5391,N_5786);
xor U6198 (N_6198,N_5179,N_5040);
xor U6199 (N_6199,N_4794,N_5152);
nand U6200 (N_6200,N_3879,N_3217);
and U6201 (N_6201,N_5136,N_5909);
nand U6202 (N_6202,N_3160,N_5518);
xnor U6203 (N_6203,N_4270,N_3800);
and U6204 (N_6204,N_5784,N_4470);
or U6205 (N_6205,N_3164,N_4705);
xor U6206 (N_6206,N_5948,N_4279);
nand U6207 (N_6207,N_3505,N_5369);
nand U6208 (N_6208,N_4175,N_3409);
nand U6209 (N_6209,N_3889,N_4462);
nor U6210 (N_6210,N_5436,N_3240);
nor U6211 (N_6211,N_5928,N_3073);
or U6212 (N_6212,N_3111,N_4771);
xnor U6213 (N_6213,N_4287,N_4600);
nand U6214 (N_6214,N_4472,N_4851);
or U6215 (N_6215,N_5297,N_4411);
xnor U6216 (N_6216,N_5851,N_4905);
nand U6217 (N_6217,N_4947,N_4599);
xor U6218 (N_6218,N_3468,N_3326);
or U6219 (N_6219,N_4997,N_4068);
nand U6220 (N_6220,N_5544,N_3456);
or U6221 (N_6221,N_4137,N_3171);
and U6222 (N_6222,N_3649,N_4671);
nand U6223 (N_6223,N_5209,N_3962);
nor U6224 (N_6224,N_4272,N_5217);
or U6225 (N_6225,N_5316,N_5961);
and U6226 (N_6226,N_5133,N_4441);
nand U6227 (N_6227,N_4630,N_3230);
or U6228 (N_6228,N_4289,N_5753);
xnor U6229 (N_6229,N_5107,N_3762);
or U6230 (N_6230,N_4039,N_3388);
or U6231 (N_6231,N_5221,N_4979);
nor U6232 (N_6232,N_5076,N_3796);
xor U6233 (N_6233,N_5410,N_5042);
nand U6234 (N_6234,N_3653,N_4616);
nor U6235 (N_6235,N_3416,N_5237);
and U6236 (N_6236,N_5468,N_5713);
nor U6237 (N_6237,N_3270,N_4791);
nand U6238 (N_6238,N_4805,N_5038);
or U6239 (N_6239,N_5521,N_5047);
and U6240 (N_6240,N_3264,N_3448);
or U6241 (N_6241,N_5776,N_4447);
nand U6242 (N_6242,N_3143,N_3545);
xnor U6243 (N_6243,N_3691,N_3187);
and U6244 (N_6244,N_4048,N_3074);
xor U6245 (N_6245,N_5759,N_5787);
xnor U6246 (N_6246,N_5486,N_3677);
nor U6247 (N_6247,N_5662,N_3589);
xor U6248 (N_6248,N_4335,N_4514);
or U6249 (N_6249,N_3891,N_4264);
nor U6250 (N_6250,N_5466,N_5963);
or U6251 (N_6251,N_5743,N_4557);
or U6252 (N_6252,N_4657,N_4539);
nand U6253 (N_6253,N_3452,N_5494);
and U6254 (N_6254,N_5537,N_4926);
or U6255 (N_6255,N_5289,N_3244);
and U6256 (N_6256,N_3954,N_5335);
xnor U6257 (N_6257,N_4230,N_4134);
and U6258 (N_6258,N_4689,N_5526);
and U6259 (N_6259,N_4660,N_5914);
nor U6260 (N_6260,N_4445,N_4740);
and U6261 (N_6261,N_4956,N_5797);
and U6262 (N_6262,N_5958,N_3330);
and U6263 (N_6263,N_4359,N_4126);
and U6264 (N_6264,N_3528,N_5843);
xor U6265 (N_6265,N_5077,N_4776);
and U6266 (N_6266,N_3543,N_4942);
or U6267 (N_6267,N_5327,N_5848);
or U6268 (N_6268,N_3945,N_3937);
xnor U6269 (N_6269,N_3994,N_5569);
or U6270 (N_6270,N_3341,N_5740);
nand U6271 (N_6271,N_5925,N_3975);
or U6272 (N_6272,N_3433,N_5429);
nand U6273 (N_6273,N_3549,N_3502);
xor U6274 (N_6274,N_5546,N_5022);
xor U6275 (N_6275,N_5463,N_3294);
xor U6276 (N_6276,N_5803,N_5365);
nor U6277 (N_6277,N_5143,N_5374);
nand U6278 (N_6278,N_3419,N_5045);
or U6279 (N_6279,N_4973,N_4921);
and U6280 (N_6280,N_3898,N_4167);
nand U6281 (N_6281,N_5794,N_3743);
and U6282 (N_6282,N_5440,N_4893);
or U6283 (N_6283,N_3903,N_4969);
xor U6284 (N_6284,N_4331,N_3179);
xor U6285 (N_6285,N_4888,N_5005);
nand U6286 (N_6286,N_3117,N_4442);
xnor U6287 (N_6287,N_4005,N_3869);
nand U6288 (N_6288,N_5088,N_4076);
xor U6289 (N_6289,N_4242,N_3787);
or U6290 (N_6290,N_5908,N_5458);
nor U6291 (N_6291,N_3500,N_5789);
or U6292 (N_6292,N_5036,N_5201);
or U6293 (N_6293,N_5216,N_4253);
xor U6294 (N_6294,N_3305,N_5078);
or U6295 (N_6295,N_3820,N_5513);
xor U6296 (N_6296,N_4317,N_3877);
nand U6297 (N_6297,N_3777,N_3944);
xor U6298 (N_6298,N_4422,N_3135);
xor U6299 (N_6299,N_5294,N_5719);
nand U6300 (N_6300,N_4348,N_5835);
nor U6301 (N_6301,N_4310,N_3694);
xnor U6302 (N_6302,N_5415,N_5596);
and U6303 (N_6303,N_4061,N_3248);
xor U6304 (N_6304,N_4625,N_4391);
or U6305 (N_6305,N_3306,N_5766);
or U6306 (N_6306,N_3807,N_5109);
and U6307 (N_6307,N_4770,N_4321);
or U6308 (N_6308,N_3457,N_3094);
or U6309 (N_6309,N_5311,N_4266);
xnor U6310 (N_6310,N_5046,N_5915);
nand U6311 (N_6311,N_3385,N_3542);
or U6312 (N_6312,N_5449,N_5011);
or U6313 (N_6313,N_5396,N_3798);
or U6314 (N_6314,N_3201,N_3613);
and U6315 (N_6315,N_5100,N_4261);
xor U6316 (N_6316,N_4731,N_3378);
and U6317 (N_6317,N_3469,N_4355);
xnor U6318 (N_6318,N_5157,N_5485);
nor U6319 (N_6319,N_4875,N_4284);
xnor U6320 (N_6320,N_3358,N_5970);
nand U6321 (N_6321,N_4150,N_3093);
nand U6322 (N_6322,N_3013,N_5469);
nor U6323 (N_6323,N_3832,N_4838);
nand U6324 (N_6324,N_4357,N_4091);
and U6325 (N_6325,N_4799,N_4419);
and U6326 (N_6326,N_5456,N_4174);
xor U6327 (N_6327,N_4772,N_5210);
nand U6328 (N_6328,N_5943,N_4158);
xnor U6329 (N_6329,N_5095,N_3098);
nand U6330 (N_6330,N_5340,N_4967);
and U6331 (N_6331,N_5863,N_3726);
nand U6332 (N_6332,N_5994,N_4410);
nor U6333 (N_6333,N_5837,N_5657);
nor U6334 (N_6334,N_4667,N_3958);
nor U6335 (N_6335,N_5428,N_5293);
or U6336 (N_6336,N_5447,N_3427);
nor U6337 (N_6337,N_4859,N_4653);
xor U6338 (N_6338,N_3272,N_3884);
nand U6339 (N_6339,N_3916,N_4088);
and U6340 (N_6340,N_5271,N_5288);
xnor U6341 (N_6341,N_4315,N_4212);
nor U6342 (N_6342,N_4306,N_4456);
xor U6343 (N_6343,N_4504,N_3070);
nor U6344 (N_6344,N_5541,N_3095);
or U6345 (N_6345,N_3196,N_4214);
and U6346 (N_6346,N_4351,N_4981);
xor U6347 (N_6347,N_5813,N_5817);
nor U6348 (N_6348,N_5652,N_3467);
nor U6349 (N_6349,N_5225,N_4953);
nor U6350 (N_6350,N_5711,N_5039);
xor U6351 (N_6351,N_5187,N_3203);
and U6352 (N_6352,N_3934,N_4320);
nand U6353 (N_6353,N_5268,N_4045);
xor U6354 (N_6354,N_4488,N_3174);
nand U6355 (N_6355,N_3122,N_4711);
nand U6356 (N_6356,N_5651,N_3119);
xnor U6357 (N_6357,N_3485,N_3000);
and U6358 (N_6358,N_3278,N_3621);
nand U6359 (N_6359,N_3007,N_4718);
or U6360 (N_6360,N_3183,N_5099);
and U6361 (N_6361,N_4153,N_3147);
nand U6362 (N_6362,N_3076,N_3626);
xnor U6363 (N_6363,N_3004,N_5579);
nand U6364 (N_6364,N_3643,N_3451);
nand U6365 (N_6365,N_4398,N_3727);
and U6366 (N_6366,N_4750,N_5790);
or U6367 (N_6367,N_4636,N_4129);
and U6368 (N_6368,N_3860,N_3974);
nand U6369 (N_6369,N_5808,N_4699);
and U6370 (N_6370,N_5354,N_3562);
nor U6371 (N_6371,N_5868,N_3406);
and U6372 (N_6372,N_4177,N_3939);
and U6373 (N_6373,N_4949,N_4896);
and U6374 (N_6374,N_3144,N_4307);
or U6375 (N_6375,N_5646,N_3430);
or U6376 (N_6376,N_3986,N_3477);
xnor U6377 (N_6377,N_4766,N_3989);
and U6378 (N_6378,N_5163,N_5473);
nand U6379 (N_6379,N_4067,N_3068);
xor U6380 (N_6380,N_4030,N_3267);
and U6381 (N_6381,N_5206,N_4584);
xnor U6382 (N_6382,N_3705,N_4231);
xor U6383 (N_6383,N_5693,N_4654);
nor U6384 (N_6384,N_4693,N_3668);
nand U6385 (N_6385,N_5658,N_4611);
or U6386 (N_6386,N_4156,N_5018);
xnor U6387 (N_6387,N_4998,N_5944);
or U6388 (N_6388,N_5126,N_3809);
nand U6389 (N_6389,N_4512,N_3327);
and U6390 (N_6390,N_5742,N_5228);
nand U6391 (N_6391,N_4752,N_3524);
nor U6392 (N_6392,N_4929,N_5954);
nor U6393 (N_6393,N_4517,N_5336);
or U6394 (N_6394,N_3193,N_4466);
xnor U6395 (N_6395,N_3586,N_3130);
or U6396 (N_6396,N_5137,N_3382);
xor U6397 (N_6397,N_5815,N_3883);
xnor U6398 (N_6398,N_5906,N_3996);
xnor U6399 (N_6399,N_5274,N_4179);
and U6400 (N_6400,N_4515,N_3766);
nor U6401 (N_6401,N_3262,N_5203);
nor U6402 (N_6402,N_3089,N_5032);
nor U6403 (N_6403,N_3598,N_5767);
nor U6404 (N_6404,N_5549,N_4440);
xnor U6405 (N_6405,N_3779,N_3243);
nor U6406 (N_6406,N_4159,N_4764);
or U6407 (N_6407,N_5115,N_4424);
nand U6408 (N_6408,N_5381,N_4622);
nand U6409 (N_6409,N_3273,N_3157);
nand U6410 (N_6410,N_3855,N_3785);
nand U6411 (N_6411,N_3819,N_4297);
xor U6412 (N_6412,N_5256,N_5781);
xor U6413 (N_6413,N_3831,N_4765);
and U6414 (N_6414,N_4203,N_4418);
nand U6415 (N_6415,N_4847,N_5418);
nand U6416 (N_6416,N_3538,N_5106);
and U6417 (N_6417,N_4963,N_3511);
nand U6418 (N_6418,N_4944,N_5202);
or U6419 (N_6419,N_4619,N_3768);
or U6420 (N_6420,N_5348,N_5153);
nor U6421 (N_6421,N_4415,N_5120);
nand U6422 (N_6422,N_4735,N_5084);
or U6423 (N_6423,N_5031,N_5417);
nand U6424 (N_6424,N_3774,N_4523);
nand U6425 (N_6425,N_4236,N_3044);
and U6426 (N_6426,N_5995,N_4362);
and U6427 (N_6427,N_5771,N_4565);
or U6428 (N_6428,N_4868,N_4260);
or U6429 (N_6429,N_5586,N_4160);
nor U6430 (N_6430,N_4629,N_3379);
nand U6431 (N_6431,N_4218,N_3642);
nand U6432 (N_6432,N_5559,N_4849);
or U6433 (N_6433,N_4020,N_5111);
nor U6434 (N_6434,N_3609,N_3453);
and U6435 (N_6435,N_5496,N_5006);
xnor U6436 (N_6436,N_4530,N_5198);
xnor U6437 (N_6437,N_5122,N_3259);
nand U6438 (N_6438,N_4716,N_3717);
nor U6439 (N_6439,N_4319,N_4404);
nor U6440 (N_6440,N_4288,N_5799);
xnor U6441 (N_6441,N_3617,N_5757);
nor U6442 (N_6442,N_4959,N_4002);
xnor U6443 (N_6443,N_4522,N_4481);
xnor U6444 (N_6444,N_3328,N_5043);
and U6445 (N_6445,N_3213,N_5861);
nand U6446 (N_6446,N_3788,N_5034);
nand U6447 (N_6447,N_3517,N_5451);
or U6448 (N_6448,N_3952,N_5108);
nand U6449 (N_6449,N_3239,N_4780);
nor U6450 (N_6450,N_5857,N_4350);
and U6451 (N_6451,N_4687,N_5498);
nand U6452 (N_6452,N_5838,N_4100);
and U6453 (N_6453,N_5007,N_3343);
nor U6454 (N_6454,N_4531,N_3594);
xnor U6455 (N_6455,N_4833,N_3047);
nor U6456 (N_6456,N_4696,N_5896);
or U6457 (N_6457,N_5694,N_5756);
xor U6458 (N_6458,N_4825,N_5968);
nand U6459 (N_6459,N_4782,N_4637);
or U6460 (N_6460,N_4254,N_4303);
nand U6461 (N_6461,N_3737,N_3102);
xor U6462 (N_6462,N_3844,N_5426);
and U6463 (N_6463,N_3045,N_4808);
xor U6464 (N_6464,N_3261,N_3624);
xnor U6465 (N_6465,N_4031,N_5675);
and U6466 (N_6466,N_4935,N_3885);
xnor U6467 (N_6467,N_4247,N_4385);
and U6468 (N_6468,N_4080,N_5252);
xnor U6469 (N_6469,N_5898,N_5497);
or U6470 (N_6470,N_5082,N_4712);
nor U6471 (N_6471,N_3926,N_3254);
nor U6472 (N_6472,N_3162,N_3030);
nor U6473 (N_6473,N_3353,N_4142);
nor U6474 (N_6474,N_4941,N_3924);
or U6475 (N_6475,N_4603,N_5457);
nor U6476 (N_6476,N_3897,N_3861);
nand U6477 (N_6477,N_3126,N_5375);
nor U6478 (N_6478,N_3572,N_4285);
or U6479 (N_6479,N_4269,N_3697);
nor U6480 (N_6480,N_5183,N_4162);
or U6481 (N_6481,N_4146,N_3797);
nand U6482 (N_6482,N_5155,N_3314);
and U6483 (N_6483,N_3630,N_4314);
nor U6484 (N_6484,N_4495,N_4282);
nor U6485 (N_6485,N_5802,N_5347);
nor U6486 (N_6486,N_5962,N_4040);
and U6487 (N_6487,N_5975,N_5124);
nand U6488 (N_6488,N_4912,N_3232);
nor U6489 (N_6489,N_3548,N_3935);
or U6490 (N_6490,N_3063,N_4524);
or U6491 (N_6491,N_4678,N_3490);
or U6492 (N_6492,N_5910,N_4602);
nand U6493 (N_6493,N_4406,N_5762);
or U6494 (N_6494,N_4071,N_5146);
xor U6495 (N_6495,N_3863,N_4738);
nor U6496 (N_6496,N_4585,N_3946);
or U6497 (N_6497,N_4787,N_4188);
xor U6498 (N_6498,N_4564,N_5671);
nor U6499 (N_6499,N_5600,N_3969);
xnor U6500 (N_6500,N_5247,N_4058);
and U6501 (N_6501,N_5903,N_5338);
nor U6502 (N_6502,N_3318,N_5979);
xnor U6503 (N_6503,N_5992,N_4672);
xor U6504 (N_6504,N_4393,N_3057);
or U6505 (N_6505,N_5620,N_5180);
nand U6506 (N_6506,N_4401,N_3016);
nand U6507 (N_6507,N_5411,N_5678);
xnor U6508 (N_6508,N_3484,N_3687);
nand U6509 (N_6509,N_3810,N_5831);
and U6510 (N_6510,N_5550,N_5476);
nor U6511 (N_6511,N_3290,N_5263);
or U6512 (N_6512,N_3848,N_5741);
or U6513 (N_6513,N_5972,N_4049);
nor U6514 (N_6514,N_3873,N_4647);
and U6515 (N_6515,N_5687,N_5384);
or U6516 (N_6516,N_3634,N_3972);
nor U6517 (N_6517,N_5382,N_5627);
nor U6518 (N_6518,N_3425,N_4692);
or U6519 (N_6519,N_4044,N_4329);
nand U6520 (N_6520,N_4783,N_5178);
nand U6521 (N_6521,N_4448,N_4439);
xor U6522 (N_6522,N_3298,N_4528);
nor U6523 (N_6523,N_4777,N_3791);
nor U6524 (N_6524,N_3116,N_5495);
and U6525 (N_6525,N_3069,N_5621);
and U6526 (N_6526,N_5892,N_5884);
nand U6527 (N_6527,N_3478,N_4760);
nand U6528 (N_6528,N_4560,N_3646);
nand U6529 (N_6529,N_4628,N_5669);
and U6530 (N_6530,N_3019,N_4345);
nand U6531 (N_6531,N_4308,N_4706);
nor U6532 (N_6532,N_5946,N_4850);
xnor U6533 (N_6533,N_5349,N_5628);
xnor U6534 (N_6534,N_3197,N_5121);
xnor U6535 (N_6535,N_4500,N_4161);
xnor U6536 (N_6536,N_5441,N_5778);
xor U6537 (N_6537,N_3410,N_5306);
or U6538 (N_6538,N_3282,N_4325);
or U6539 (N_6539,N_5129,N_4111);
xnor U6540 (N_6540,N_5918,N_5359);
xor U6541 (N_6541,N_4709,N_5937);
and U6542 (N_6542,N_5166,N_4698);
or U6543 (N_6543,N_4417,N_3555);
or U6544 (N_6544,N_4316,N_5260);
nor U6545 (N_6545,N_5660,N_3930);
or U6546 (N_6546,N_3142,N_5233);
xor U6547 (N_6547,N_5530,N_5542);
xor U6548 (N_6548,N_5984,N_3288);
nand U6549 (N_6549,N_4388,N_4964);
nor U6550 (N_6550,N_3192,N_3256);
nor U6551 (N_6551,N_5319,N_3445);
xor U6552 (N_6552,N_3475,N_5733);
xor U6553 (N_6553,N_4136,N_5876);
xor U6554 (N_6554,N_3097,N_5438);
nor U6555 (N_6555,N_4496,N_3664);
xnor U6556 (N_6556,N_5357,N_3675);
nor U6557 (N_6557,N_3277,N_3868);
and U6558 (N_6558,N_3793,N_5147);
or U6559 (N_6559,N_3830,N_4220);
nand U6560 (N_6560,N_3583,N_5309);
nand U6561 (N_6561,N_3967,N_5717);
and U6562 (N_6562,N_4729,N_4183);
or U6563 (N_6563,N_3943,N_3571);
or U6564 (N_6564,N_3146,N_4553);
and U6565 (N_6565,N_4798,N_5655);
xor U6566 (N_6566,N_5872,N_4761);
or U6567 (N_6567,N_5966,N_3003);
xor U6568 (N_6568,N_5363,N_3048);
nand U6569 (N_6569,N_4121,N_3285);
nand U6570 (N_6570,N_3618,N_4394);
and U6571 (N_6571,N_5399,N_3058);
or U6572 (N_6572,N_5894,N_5930);
nand U6573 (N_6573,N_5241,N_5949);
nor U6574 (N_6574,N_3914,N_3289);
nand U6575 (N_6575,N_5886,N_4395);
nor U6576 (N_6576,N_4244,N_3495);
nor U6577 (N_6577,N_4449,N_5037);
and U6578 (N_6578,N_3728,N_4239);
xor U6579 (N_6579,N_4305,N_4758);
xor U6580 (N_6580,N_3706,N_4618);
and U6581 (N_6581,N_4025,N_5197);
and U6582 (N_6582,N_3764,N_5478);
nor U6583 (N_6583,N_4743,N_5159);
and U6584 (N_6584,N_5527,N_3920);
and U6585 (N_6585,N_3020,N_3823);
and U6586 (N_6586,N_3284,N_3059);
xnor U6587 (N_6587,N_4047,N_4721);
and U6588 (N_6588,N_3647,N_4508);
nand U6589 (N_6589,N_5315,N_5313);
nor U6590 (N_6590,N_5705,N_3291);
or U6591 (N_6591,N_4811,N_3322);
nor U6592 (N_6592,N_3681,N_3050);
nand U6593 (N_6593,N_3509,N_3564);
or U6594 (N_6594,N_5123,N_5637);
xnor U6595 (N_6595,N_3838,N_4570);
xor U6596 (N_6596,N_3595,N_4513);
xor U6597 (N_6597,N_5004,N_4918);
and U6598 (N_6598,N_5303,N_4559);
nand U6599 (N_6599,N_3488,N_4621);
nand U6600 (N_6600,N_3600,N_3532);
nand U6601 (N_6601,N_3250,N_3199);
and U6602 (N_6602,N_5862,N_3721);
nand U6603 (N_6603,N_5989,N_3340);
nor U6604 (N_6604,N_3408,N_4029);
xnor U6605 (N_6605,N_5667,N_4290);
nor U6606 (N_6606,N_4538,N_3274);
or U6607 (N_6607,N_5219,N_3874);
xnor U6608 (N_6608,N_4593,N_3857);
and U6609 (N_6609,N_5394,N_5768);
nor U6610 (N_6610,N_5534,N_3713);
xor U6611 (N_6611,N_3576,N_5361);
or U6612 (N_6612,N_5539,N_4273);
and U6613 (N_6613,N_3627,N_5517);
nor U6614 (N_6614,N_3578,N_3816);
and U6615 (N_6615,N_4324,N_3703);
xnor U6616 (N_6616,N_4286,N_5257);
xnor U6617 (N_6617,N_3363,N_3008);
and U6618 (N_6618,N_5551,N_3980);
or U6619 (N_6619,N_3389,N_3993);
xnor U6620 (N_6620,N_4477,N_3354);
nand U6621 (N_6621,N_3397,N_4105);
and U6622 (N_6622,N_3901,N_4124);
xnor U6623 (N_6623,N_3133,N_3915);
nand U6624 (N_6624,N_5001,N_5901);
and U6625 (N_6625,N_4624,N_4834);
and U6626 (N_6626,N_4640,N_3921);
nand U6627 (N_6627,N_5985,N_3113);
nor U6628 (N_6628,N_5976,N_5278);
xor U6629 (N_6629,N_4008,N_3066);
nor U6630 (N_6630,N_4018,N_3892);
xor U6631 (N_6631,N_5230,N_3862);
or U6632 (N_6632,N_5402,N_5443);
nand U6633 (N_6633,N_4154,N_4259);
or U6634 (N_6634,N_4277,N_3176);
xnor U6635 (N_6635,N_4390,N_5640);
xnor U6636 (N_6636,N_4063,N_3252);
nand U6637 (N_6637,N_5969,N_3597);
nor U6638 (N_6638,N_5322,N_5017);
nand U6639 (N_6639,N_3329,N_5877);
xor U6640 (N_6640,N_3704,N_3474);
nor U6641 (N_6641,N_3170,N_5455);
and U6642 (N_6642,N_3933,N_4389);
nor U6643 (N_6643,N_5779,N_3027);
xnor U6644 (N_6644,N_3833,N_4060);
nand U6645 (N_6645,N_3374,N_3983);
xor U6646 (N_6646,N_5830,N_4106);
or U6647 (N_6647,N_4923,N_5081);
xor U6648 (N_6648,N_4763,N_3657);
or U6649 (N_6649,N_4656,N_4053);
or U6650 (N_6650,N_5253,N_3673);
or U6651 (N_6651,N_4860,N_5453);
nor U6652 (N_6652,N_3712,N_4009);
nand U6653 (N_6653,N_4938,N_5158);
xor U6654 (N_6654,N_4715,N_4605);
xor U6655 (N_6655,N_3034,N_4634);
nor U6656 (N_6656,N_5025,N_5145);
xor U6657 (N_6657,N_4563,N_5679);
nand U6658 (N_6658,N_4820,N_4369);
nor U6659 (N_6659,N_5587,N_3182);
nand U6660 (N_6660,N_5085,N_3569);
nor U6661 (N_6661,N_5607,N_3880);
nand U6662 (N_6662,N_4708,N_5450);
and U6663 (N_6663,N_4019,N_4326);
nor U6664 (N_6664,N_3309,N_5804);
nand U6665 (N_6665,N_5570,N_5702);
and U6666 (N_6666,N_5722,N_4853);
nor U6667 (N_6667,N_4762,N_5128);
xnor U6668 (N_6668,N_3181,N_4006);
xor U6669 (N_6669,N_3313,N_5996);
or U6670 (N_6670,N_3867,N_4828);
and U6671 (N_6671,N_3959,N_3337);
xor U6672 (N_6672,N_3669,N_3645);
or U6673 (N_6673,N_3709,N_4810);
xnor U6674 (N_6674,N_3992,N_3604);
and U6675 (N_6675,N_4198,N_3208);
and U6676 (N_6676,N_3812,N_4208);
xnor U6677 (N_6677,N_4638,N_4592);
xnor U6678 (N_6678,N_5254,N_5821);
or U6679 (N_6679,N_5487,N_5665);
nor U6680 (N_6680,N_4191,N_3932);
and U6681 (N_6681,N_4732,N_5061);
or U6682 (N_6682,N_5140,N_4458);
nand U6683 (N_6683,N_3811,N_5755);
or U6684 (N_6684,N_5854,N_3553);
and U6685 (N_6685,N_5847,N_4405);
and U6686 (N_6686,N_4567,N_3888);
or U6687 (N_6687,N_4876,N_5950);
and U6688 (N_6688,N_5947,N_3850);
nand U6689 (N_6689,N_5057,N_4871);
nor U6690 (N_6690,N_5446,N_4034);
or U6691 (N_6691,N_3922,N_5113);
xnor U6692 (N_6692,N_4631,N_3128);
and U6693 (N_6693,N_5506,N_5239);
nor U6694 (N_6694,N_4858,N_4746);
and U6695 (N_6695,N_4240,N_4210);
nand U6696 (N_6696,N_3753,N_5721);
nor U6697 (N_6697,N_3821,N_5697);
nand U6698 (N_6698,N_4914,N_3953);
or U6699 (N_6699,N_3758,N_4710);
nand U6700 (N_6700,N_3025,N_3344);
and U6701 (N_6701,N_3949,N_5220);
xnor U6702 (N_6702,N_4510,N_5101);
xnor U6703 (N_6703,N_4407,N_4863);
and U6704 (N_6704,N_4756,N_4726);
nand U6705 (N_6705,N_5514,N_5093);
nor U6706 (N_6706,N_4571,N_4627);
nor U6707 (N_6707,N_3661,N_5063);
and U6708 (N_6708,N_4714,N_3825);
and U6709 (N_6709,N_5284,N_5477);
and U6710 (N_6710,N_5337,N_5933);
nor U6711 (N_6711,N_4902,N_3619);
and U6712 (N_6712,N_3757,N_3042);
or U6713 (N_6713,N_4955,N_4669);
xor U6714 (N_6714,N_5181,N_5523);
nand U6715 (N_6715,N_3817,N_3558);
nand U6716 (N_6716,N_4296,N_5070);
and U6717 (N_6717,N_3688,N_3824);
and U6718 (N_6718,N_4685,N_3229);
nand U6719 (N_6719,N_4381,N_3387);
or U6720 (N_6720,N_5154,N_5028);
xor U6721 (N_6721,N_5398,N_3899);
and U6722 (N_6722,N_3464,N_5117);
and U6723 (N_6723,N_5528,N_3984);
nor U6724 (N_6724,N_3590,N_3338);
nor U6725 (N_6725,N_4219,N_3498);
nor U6726 (N_6726,N_5421,N_5516);
and U6727 (N_6727,N_5188,N_5352);
or U6728 (N_6728,N_5921,N_4925);
xor U6729 (N_6729,N_4877,N_4910);
nand U6730 (N_6730,N_5645,N_4139);
nor U6731 (N_6731,N_4353,N_5172);
or U6732 (N_6732,N_5118,N_3188);
or U6733 (N_6733,N_4886,N_3279);
xor U6734 (N_6734,N_5971,N_4754);
xnor U6735 (N_6735,N_3925,N_4845);
xor U6736 (N_6736,N_5437,N_5616);
and U6737 (N_6737,N_5706,N_4471);
nand U6738 (N_6738,N_3878,N_5704);
or U6739 (N_6739,N_4681,N_3711);
or U6740 (N_6740,N_4235,N_3971);
xor U6741 (N_6741,N_3265,N_4831);
nor U6742 (N_6742,N_5223,N_5916);
or U6743 (N_6743,N_5643,N_4104);
xor U6744 (N_6744,N_4083,N_5390);
and U6745 (N_6745,N_5714,N_3763);
nor U6746 (N_6746,N_3271,N_3973);
xor U6747 (N_6747,N_5590,N_4753);
or U6748 (N_6748,N_5683,N_3837);
and U6749 (N_6749,N_3263,N_4066);
nand U6750 (N_6750,N_5328,N_3302);
or U6751 (N_6751,N_3442,N_5718);
and U6752 (N_6752,N_3177,N_4864);
and U6753 (N_6753,N_5408,N_4812);
nand U6754 (N_6754,N_3346,N_4541);
or U6755 (N_6755,N_4633,N_5888);
and U6756 (N_6756,N_4255,N_4879);
nor U6757 (N_6757,N_4554,N_4639);
xor U6758 (N_6758,N_4267,N_5572);
xnor U6759 (N_6759,N_5840,N_5016);
xor U6760 (N_6760,N_4586,N_4806);
or U6761 (N_6761,N_4376,N_5879);
or U6762 (N_6762,N_3398,N_4840);
nor U6763 (N_6763,N_4378,N_4932);
xnor U6764 (N_6764,N_4012,N_5556);
nand U6765 (N_6765,N_4149,N_3251);
nor U6766 (N_6766,N_5653,N_5677);
and U6767 (N_6767,N_5819,N_4217);
and U6768 (N_6768,N_4569,N_5934);
xor U6769 (N_6769,N_4759,N_3312);
and U6770 (N_6770,N_5601,N_5827);
xor U6771 (N_6771,N_3420,N_4841);
nand U6772 (N_6772,N_3235,N_4972);
or U6773 (N_6773,N_4492,N_5432);
xnor U6774 (N_6774,N_3350,N_5668);
xnor U6775 (N_6775,N_3981,N_3081);
or U6776 (N_6776,N_4598,N_5870);
nand U6777 (N_6777,N_3599,N_3231);
nand U6778 (N_6778,N_5281,N_4201);
xnor U6779 (N_6779,N_3539,N_3242);
and U6780 (N_6780,N_4256,N_4857);
nor U6781 (N_6781,N_3806,N_3391);
xor U6782 (N_6782,N_5612,N_4796);
nor U6783 (N_6783,N_5849,N_4995);
nand U6784 (N_6784,N_5750,N_4228);
xnor U6785 (N_6785,N_5685,N_5839);
and U6786 (N_6786,N_4120,N_3011);
or U6787 (N_6787,N_5207,N_4110);
xnor U6788 (N_6788,N_4502,N_3580);
nor U6789 (N_6789,N_3895,N_4178);
nor U6790 (N_6790,N_4744,N_5795);
nor U6791 (N_6791,N_4346,N_3101);
nand U6792 (N_6792,N_5832,N_4059);
nand U6793 (N_6793,N_5058,N_3169);
xor U6794 (N_6794,N_5923,N_3257);
and U6795 (N_6795,N_5186,N_4356);
or U6796 (N_6796,N_5508,N_5619);
nor U6797 (N_6797,N_5792,N_5341);
or U6798 (N_6798,N_4336,N_4813);
or U6799 (N_6799,N_4986,N_5246);
or U6800 (N_6800,N_4717,N_5545);
nand U6801 (N_6801,N_4945,N_4609);
nor U6802 (N_6802,N_4024,N_3942);
or U6803 (N_6803,N_4026,N_3293);
xnor U6804 (N_6804,N_4133,N_4251);
xnor U6805 (N_6805,N_4984,N_5385);
nand U6806 (N_6806,N_5053,N_3009);
and U6807 (N_6807,N_3096,N_3557);
nand U6808 (N_6808,N_5864,N_3091);
or U6809 (N_6809,N_5531,N_5796);
nand U6810 (N_6810,N_4587,N_3603);
nor U6811 (N_6811,N_4869,N_3461);
nor U6812 (N_6812,N_4119,N_4115);
or U6813 (N_6813,N_4518,N_3132);
or U6814 (N_6814,N_3361,N_4383);
nor U6815 (N_6815,N_3321,N_5977);
and U6816 (N_6816,N_5148,N_4659);
xnor U6817 (N_6817,N_5634,N_4582);
or U6818 (N_6818,N_4184,N_3403);
or U6819 (N_6819,N_5304,N_5691);
nand U6820 (N_6820,N_4028,N_5666);
nand U6821 (N_6821,N_4473,N_3492);
or U6822 (N_6822,N_5820,N_3670);
and U6823 (N_6823,N_3760,N_5261);
nor U6824 (N_6824,N_3616,N_4960);
or U6825 (N_6825,N_3733,N_4931);
and U6826 (N_6826,N_3886,N_3929);
nand U6827 (N_6827,N_5532,N_5940);
xor U6828 (N_6828,N_5698,N_5200);
xor U6829 (N_6829,N_4138,N_3606);
and U6830 (N_6830,N_3202,N_4425);
nor U6831 (N_6831,N_3307,N_3150);
nor U6832 (N_6832,N_3198,N_3504);
xor U6833 (N_6833,N_5728,N_5350);
or U6834 (N_6834,N_3826,N_5695);
nor U6835 (N_6835,N_4122,N_4085);
and U6836 (N_6836,N_5512,N_3376);
nor U6837 (N_6837,N_5484,N_5955);
and U6838 (N_6838,N_5712,N_4202);
and U6839 (N_6839,N_3676,N_3245);
xnor U6840 (N_6840,N_5760,N_4042);
xnor U6841 (N_6841,N_3735,N_4165);
nor U6842 (N_6842,N_5370,N_5670);
nand U6843 (N_6843,N_4503,N_3552);
or U6844 (N_6844,N_3221,N_4223);
xnor U6845 (N_6845,N_5599,N_5490);
xor U6846 (N_6846,N_3786,N_3625);
nor U6847 (N_6847,N_4434,N_3507);
nor U6848 (N_6848,N_3412,N_3701);
nor U6849 (N_6849,N_4691,N_4035);
or U6850 (N_6850,N_3767,N_4843);
nand U6851 (N_6851,N_5262,N_4595);
nor U6852 (N_6852,N_3525,N_3596);
and U6853 (N_6853,N_4195,N_4339);
xnor U6854 (N_6854,N_4293,N_4525);
or U6855 (N_6855,N_5959,N_4928);
and U6856 (N_6856,N_4568,N_4899);
nand U6857 (N_6857,N_3579,N_5564);
xnor U6858 (N_6858,N_3991,N_5266);
xor U6859 (N_6859,N_3927,N_4968);
or U6860 (N_6860,N_5822,N_4373);
xor U6861 (N_6861,N_3955,N_5480);
or U6862 (N_6862,N_5334,N_5676);
and U6863 (N_6863,N_4688,N_3623);
nand U6864 (N_6864,N_4344,N_3266);
or U6865 (N_6865,N_3140,N_5344);
xnor U6866 (N_6866,N_4884,N_5112);
xnor U6867 (N_6867,N_3778,N_3489);
nor U6868 (N_6868,N_4908,N_5769);
nand U6869 (N_6869,N_4982,N_4302);
or U6870 (N_6870,N_5734,N_4372);
or U6871 (N_6871,N_5852,N_4457);
xnor U6872 (N_6872,N_5904,N_5842);
nand U6873 (N_6873,N_4817,N_5502);
nand U6874 (N_6874,N_3801,N_4623);
nor U6875 (N_6875,N_5059,N_3575);
and U6876 (N_6876,N_4751,N_5089);
nor U6877 (N_6877,N_5503,N_3369);
nand U6878 (N_6878,N_3872,N_4719);
and U6879 (N_6879,N_4818,N_5701);
nand U6880 (N_6880,N_5273,N_5454);
and U6881 (N_6881,N_3390,N_4819);
and U6882 (N_6882,N_4241,N_3131);
nor U6883 (N_6883,N_4014,N_5744);
nor U6884 (N_6884,N_4209,N_3383);
nor U6885 (N_6885,N_4976,N_3902);
nor U6886 (N_6886,N_5568,N_4954);
or U6887 (N_6887,N_5836,N_4615);
xnor U6888 (N_6888,N_4257,N_5991);
nor U6889 (N_6889,N_4300,N_4641);
nand U6890 (N_6890,N_5500,N_3696);
nor U6891 (N_6891,N_5561,N_5891);
and U6892 (N_6892,N_5967,N_4607);
xor U6893 (N_6893,N_5282,N_3740);
or U6894 (N_6894,N_3638,N_3454);
or U6895 (N_6895,N_4507,N_3486);
or U6896 (N_6896,N_4384,N_5816);
nor U6897 (N_6897,N_4920,N_4123);
nand U6898 (N_6898,N_4069,N_5290);
and U6899 (N_6899,N_5887,N_5533);
nand U6900 (N_6900,N_4062,N_5211);
nor U6901 (N_6901,N_5105,N_4823);
nor U6902 (N_6902,N_3497,N_3702);
nor U6903 (N_6903,N_4511,N_3948);
nor U6904 (N_6904,N_3218,N_5242);
nor U6905 (N_6905,N_5801,N_4460);
nand U6906 (N_6906,N_4943,N_5618);
or U6907 (N_6907,N_5639,N_5598);
nand U6908 (N_6908,N_4087,N_5555);
or U6909 (N_6909,N_5935,N_5091);
xnor U6910 (N_6910,N_3310,N_3372);
nor U6911 (N_6911,N_4589,N_4830);
nor U6912 (N_6912,N_5773,N_5636);
nand U6913 (N_6913,N_3125,N_5013);
and U6914 (N_6914,N_4962,N_3637);
xor U6915 (N_6915,N_5150,N_5900);
xnor U6916 (N_6916,N_3936,N_3121);
or U6917 (N_6917,N_3365,N_3652);
nor U6918 (N_6918,N_4101,N_5871);
nor U6919 (N_6919,N_5874,N_5855);
or U6920 (N_6920,N_5096,N_5229);
nor U6921 (N_6921,N_4501,N_3866);
xor U6922 (N_6922,N_4889,N_3723);
nor U6923 (N_6923,N_3689,N_5614);
nor U6924 (N_6924,N_3839,N_5942);
nand U6925 (N_6925,N_4107,N_3400);
xnor U6926 (N_6926,N_5434,N_5459);
nor U6927 (N_6927,N_4632,N_4204);
nand U6928 (N_6928,N_5809,N_4003);
nand U6929 (N_6929,N_5739,N_5448);
and U6930 (N_6930,N_4233,N_5173);
nor U6931 (N_6931,N_5425,N_5828);
nor U6932 (N_6932,N_4130,N_5405);
and U6933 (N_6933,N_5175,N_5881);
or U6934 (N_6934,N_4578,N_3679);
nand U6935 (N_6935,N_3665,N_3184);
nand U6936 (N_6936,N_3871,N_5723);
xor U6937 (N_6937,N_5467,N_5552);
or U6938 (N_6938,N_3658,N_5044);
or U6939 (N_6939,N_4304,N_5604);
xor U6940 (N_6940,N_5292,N_3629);
xnor U6941 (N_6941,N_3405,N_5811);
nand U6942 (N_6942,N_3790,N_3772);
nand U6943 (N_6943,N_3537,N_3732);
xor U6944 (N_6944,N_3882,N_3209);
and U6945 (N_6945,N_4258,N_3033);
and U6946 (N_6946,N_5226,N_5932);
and U6947 (N_6947,N_5160,N_4084);
and U6948 (N_6948,N_5919,N_4428);
nand U6949 (N_6949,N_5264,N_4807);
nand U6950 (N_6950,N_3957,N_5474);
nand U6951 (N_6951,N_3666,N_5403);
nor U6952 (N_6952,N_4141,N_3424);
nor U6953 (N_6953,N_3628,N_4459);
or U6954 (N_6954,N_5275,N_5890);
and U6955 (N_6955,N_5372,N_4720);
nand U6956 (N_6956,N_4757,N_3366);
nand U6957 (N_6957,N_3692,N_3200);
nor U6958 (N_6958,N_5465,N_4309);
and U6959 (N_6959,N_4490,N_3684);
xnor U6960 (N_6960,N_4370,N_5214);
nand U6961 (N_6961,N_4784,N_3565);
xor U6962 (N_6962,N_5692,N_4670);
and U6963 (N_6963,N_4663,N_4903);
or U6964 (N_6964,N_4057,N_5507);
nand U6965 (N_6965,N_4227,N_5865);
nor U6966 (N_6966,N_3755,N_4294);
nand U6967 (N_6967,N_3465,N_5806);
nand U6968 (N_6968,N_3088,N_3299);
xor U6969 (N_6969,N_3026,N_3769);
nand U6970 (N_6970,N_4206,N_4064);
nor U6971 (N_6971,N_5680,N_3722);
xor U6972 (N_6972,N_5433,N_4465);
and U6973 (N_6973,N_3295,N_3631);
and U6974 (N_6974,N_4237,N_3015);
nand U6975 (N_6975,N_3636,N_4591);
nand U6976 (N_6976,N_3449,N_4793);
xor U6977 (N_6977,N_5102,N_3049);
xor U6978 (N_6978,N_4577,N_3345);
nor U6979 (N_6979,N_4778,N_5295);
and U6980 (N_6980,N_3966,N_5562);
or U6981 (N_6981,N_4363,N_4802);
nand U6982 (N_6982,N_4098,N_3893);
nor U6983 (N_6983,N_4679,N_4883);
nor U6984 (N_6984,N_4521,N_3180);
xnor U6985 (N_6985,N_5800,N_5737);
nor U6986 (N_6986,N_5707,N_3746);
xnor U6987 (N_6987,N_5807,N_3749);
xor U6988 (N_6988,N_3145,N_3395);
xnor U6989 (N_6989,N_5764,N_3896);
and U6990 (N_6990,N_4113,N_4147);
and U6991 (N_6991,N_5169,N_3017);
and U6992 (N_6992,N_3396,N_4392);
nor U6993 (N_6993,N_5312,N_5489);
xor U6994 (N_6994,N_3961,N_3418);
and U6995 (N_6995,N_5519,N_5255);
and U6996 (N_6996,N_3371,N_4664);
and U6997 (N_6997,N_3054,N_5973);
or U6998 (N_6998,N_5071,N_4604);
nand U6999 (N_6999,N_5104,N_5716);
or U7000 (N_7000,N_4723,N_4574);
and U7001 (N_7001,N_4870,N_3818);
or U7002 (N_7002,N_4588,N_5606);
and U7003 (N_7003,N_5170,N_3260);
or U7004 (N_7004,N_5765,N_5622);
nand U7005 (N_7005,N_4375,N_3570);
xor U7006 (N_7006,N_3380,N_4792);
nor U7007 (N_7007,N_4550,N_5931);
xor U7008 (N_7008,N_4610,N_3014);
nand U7009 (N_7009,N_5654,N_4051);
or U7010 (N_7010,N_5132,N_3756);
nor U7011 (N_7011,N_5727,N_5920);
xnor U7012 (N_7012,N_3970,N_3650);
or U7013 (N_7013,N_3038,N_3982);
nor U7014 (N_7014,N_5424,N_3592);
nor U7015 (N_7015,N_5987,N_4742);
nor U7016 (N_7016,N_3308,N_3022);
nand U7017 (N_7017,N_5060,N_5912);
and U7018 (N_7018,N_4200,N_4700);
nand U7019 (N_7019,N_3138,N_5196);
nor U7020 (N_7020,N_4461,N_4143);
xnor U7021 (N_7021,N_5051,N_4192);
nand U7022 (N_7022,N_5470,N_4662);
or U7023 (N_7023,N_5883,N_4262);
nand U7024 (N_7024,N_4478,N_3280);
nor U7025 (N_7025,N_3032,N_4668);
nor U7026 (N_7026,N_3533,N_4548);
nor U7027 (N_7027,N_5407,N_3336);
and U7028 (N_7028,N_3124,N_5538);
nand U7029 (N_7029,N_4413,N_3978);
nor U7030 (N_7030,N_3905,N_3977);
xor U7031 (N_7031,N_5805,N_3587);
nand U7032 (N_7032,N_5362,N_5610);
or U7033 (N_7033,N_3226,N_3950);
or U7034 (N_7034,N_3185,N_4892);
nor U7035 (N_7035,N_3751,N_3331);
xnor U7036 (N_7036,N_4516,N_3834);
and U7037 (N_7037,N_3582,N_3853);
or U7038 (N_7038,N_4725,N_3997);
and U7039 (N_7039,N_3963,N_4027);
xor U7040 (N_7040,N_4187,N_3466);
xor U7041 (N_7041,N_4648,N_4436);
nand U7042 (N_7042,N_3514,N_5780);
nand U7043 (N_7043,N_3563,N_5302);
xor U7044 (N_7044,N_4455,N_5190);
xnor U7045 (N_7045,N_4974,N_5873);
and U7046 (N_7046,N_4701,N_4332);
and U7047 (N_7047,N_5749,N_5626);
nand U7048 (N_7048,N_5623,N_3917);
nand U7049 (N_7049,N_5673,N_3827);
xnor U7050 (N_7050,N_3386,N_5774);
nand U7051 (N_7051,N_3215,N_4371);
or U7052 (N_7052,N_3377,N_4649);
or U7053 (N_7053,N_3335,N_3651);
or U7054 (N_7054,N_5656,N_5735);
nor U7055 (N_7055,N_4420,N_4573);
and U7056 (N_7056,N_5326,N_3087);
or U7057 (N_7057,N_3968,N_5305);
and U7058 (N_7058,N_4895,N_3053);
or U7059 (N_7059,N_5567,N_3316);
and U7060 (N_7060,N_5464,N_3072);
nor U7061 (N_7061,N_5002,N_3210);
xnor U7062 (N_7062,N_3660,N_5625);
nor U7063 (N_7063,N_4112,N_5234);
nand U7064 (N_7064,N_3402,N_5251);
nor U7065 (N_7065,N_5243,N_4397);
nor U7066 (N_7066,N_5030,N_3530);
or U7067 (N_7067,N_4786,N_3075);
nor U7068 (N_7068,N_5086,N_5731);
and U7069 (N_7069,N_3482,N_5945);
nor U7070 (N_7070,N_4873,N_5584);
nand U7071 (N_7071,N_3134,N_5566);
nand U7072 (N_7072,N_5576,N_3079);
or U7073 (N_7073,N_5395,N_5167);
xor U7074 (N_7074,N_4975,N_5648);
xor U7075 (N_7075,N_5481,N_4990);
or U7076 (N_7076,N_3588,N_3656);
or U7077 (N_7077,N_5383,N_3822);
and U7078 (N_7078,N_4092,N_5208);
nand U7079 (N_7079,N_5232,N_3988);
xnor U7080 (N_7080,N_5520,N_5525);
xor U7081 (N_7081,N_5259,N_4650);
nand U7082 (N_7082,N_4505,N_5317);
nor U7083 (N_7083,N_5431,N_4292);
and U7084 (N_7084,N_5406,N_3493);
nor U7085 (N_7085,N_3725,N_5184);
and U7086 (N_7086,N_5364,N_3035);
nand U7087 (N_7087,N_4412,N_4435);
nand U7088 (N_7088,N_5269,N_3759);
nand U7089 (N_7089,N_4832,N_5833);
and U7090 (N_7090,N_5343,N_3655);
and U7091 (N_7091,N_3547,N_3700);
or U7092 (N_7092,N_3165,N_5069);
and U7093 (N_7093,N_5419,N_3317);
nand U7094 (N_7094,N_3472,N_4774);
xor U7095 (N_7095,N_4900,N_4196);
and U7096 (N_7096,N_4323,N_5192);
and U7097 (N_7097,N_4166,N_5889);
and U7098 (N_7098,N_4498,N_3506);
nand U7099 (N_7099,N_3046,N_4583);
nor U7100 (N_7100,N_3607,N_3481);
nor U7101 (N_7101,N_4674,N_4023);
xor U7102 (N_7102,N_5818,N_4016);
or U7103 (N_7103,N_3906,N_3431);
nor U7104 (N_7104,N_5700,N_4773);
nor U7105 (N_7105,N_3219,N_3351);
nand U7106 (N_7106,N_5661,N_3487);
or U7107 (N_7107,N_3067,N_3859);
xor U7108 (N_7108,N_4734,N_5573);
nor U7109 (N_7109,N_3640,N_3912);
and U7110 (N_7110,N_5853,N_3515);
xor U7111 (N_7111,N_5003,N_3870);
xnor U7112 (N_7112,N_3865,N_4694);
and U7113 (N_7113,N_3447,N_3356);
and U7114 (N_7114,N_3612,N_3770);
nand U7115 (N_7115,N_5195,N_4013);
nand U7116 (N_7116,N_4767,N_3802);
or U7117 (N_7117,N_4283,N_3455);
nand U7118 (N_7118,N_4327,N_5064);
or U7119 (N_7119,N_5393,N_5751);
or U7120 (N_7120,N_5000,N_3858);
and U7121 (N_7121,N_3168,N_4826);
nor U7122 (N_7122,N_4275,N_3808);
and U7123 (N_7123,N_5699,N_3083);
nand U7124 (N_7124,N_3156,N_4374);
nand U7125 (N_7125,N_5353,N_4157);
and U7126 (N_7126,N_4809,N_5471);
nand U7127 (N_7127,N_4280,N_5738);
or U7128 (N_7128,N_4163,N_3568);
xor U7129 (N_7129,N_4898,N_4399);
xor U7130 (N_7130,N_5647,N_5020);
nor U7131 (N_7131,N_5856,N_5980);
nand U7132 (N_7132,N_5859,N_3435);
and U7133 (N_7133,N_5591,N_4697);
nor U7134 (N_7134,N_5023,N_4861);
nand U7135 (N_7135,N_5240,N_4909);
and U7136 (N_7136,N_4520,N_3370);
nand U7137 (N_7137,N_5435,N_3281);
nor U7138 (N_7138,N_3851,N_3105);
xor U7139 (N_7139,N_4489,N_4482);
nor U7140 (N_7140,N_3001,N_4409);
nand U7141 (N_7141,N_4652,N_5729);
xnor U7142 (N_7142,N_4468,N_5329);
and U7143 (N_7143,N_3663,N_4540);
and U7144 (N_7144,N_5829,N_3979);
xnor U7145 (N_7145,N_5400,N_3178);
xnor U7146 (N_7146,N_4077,N_3842);
xor U7147 (N_7147,N_4094,N_3325);
nand U7148 (N_7148,N_5199,N_3167);
xor U7149 (N_7149,N_5592,N_3503);
nor U7150 (N_7150,N_5703,N_5420);
or U7151 (N_7151,N_4140,N_3804);
or U7152 (N_7152,N_3360,N_3695);
nand U7153 (N_7153,N_4011,N_5547);
and U7154 (N_7154,N_3843,N_5323);
nor U7155 (N_7155,N_3106,N_3644);
nor U7156 (N_7156,N_4252,N_4038);
nor U7157 (N_7157,N_3375,N_5770);
xnor U7158 (N_7158,N_4103,N_4534);
and U7159 (N_7159,N_4483,N_3614);
xor U7160 (N_7160,N_3161,N_3421);
or U7161 (N_7161,N_3362,N_3078);
and U7162 (N_7162,N_3508,N_3720);
xor U7163 (N_7163,N_5880,N_3407);
xnor U7164 (N_7164,N_5560,N_4558);
or U7165 (N_7165,N_5488,N_5726);
or U7166 (N_7166,N_3875,N_3710);
nand U7167 (N_7167,N_5193,N_3163);
xnor U7168 (N_7168,N_5015,N_5812);
nand U7169 (N_7169,N_3931,N_3513);
or U7170 (N_7170,N_4839,N_5754);
nand U7171 (N_7171,N_3414,N_5585);
nand U7172 (N_7172,N_5907,N_4916);
xor U7173 (N_7173,N_3744,N_3446);
nand U7174 (N_7174,N_5127,N_5633);
or U7175 (N_7175,N_5593,N_5141);
nor U7176 (N_7176,N_5893,N_5684);
nor U7177 (N_7177,N_5283,N_4913);
and U7178 (N_7178,N_4499,N_5603);
nand U7179 (N_7179,N_4403,N_5672);
xor U7180 (N_7180,N_5185,N_3429);
nor U7181 (N_7181,N_5720,N_5615);
nand U7182 (N_7182,N_4856,N_5558);
xnor U7183 (N_7183,N_5577,N_4185);
and U7184 (N_7184,N_5149,N_5092);
nor U7185 (N_7185,N_3699,N_4666);
xnor U7186 (N_7186,N_4509,N_4263);
nand U7187 (N_7187,N_5663,N_4086);
or U7188 (N_7188,N_4655,N_4822);
nand U7189 (N_7189,N_5321,N_5624);
xnor U7190 (N_7190,N_5758,N_4690);
xnor U7191 (N_7191,N_4197,N_3223);
xnor U7192 (N_7192,N_3667,N_5009);
or U7193 (N_7193,N_4897,N_3357);
nand U7194 (N_7194,N_5905,N_3752);
and U7195 (N_7195,N_3275,N_4352);
or U7196 (N_7196,N_4872,N_5745);
or U7197 (N_7197,N_5174,N_3754);
and U7198 (N_7198,N_3320,N_3522);
and U7199 (N_7199,N_4181,N_3349);
and U7200 (N_7200,N_5224,N_4365);
nor U7201 (N_7201,N_5072,N_3186);
xnor U7202 (N_7202,N_3641,N_3241);
nand U7203 (N_7203,N_5641,N_5936);
nand U7204 (N_7204,N_5632,N_5065);
and U7205 (N_7205,N_5483,N_4010);
nand U7206 (N_7206,N_3815,N_5339);
and U7207 (N_7207,N_4862,N_4867);
nor U7208 (N_7208,N_5244,N_4789);
or U7209 (N_7209,N_5814,N_3550);
nor U7210 (N_7210,N_3531,N_3615);
nand U7211 (N_7211,N_4620,N_3339);
nor U7212 (N_7212,N_3092,N_3690);
nor U7213 (N_7213,N_4446,N_5504);
nand U7214 (N_7214,N_5460,N_4438);
or U7215 (N_7215,N_5846,N_4852);
xor U7216 (N_7216,N_3148,N_3894);
nor U7217 (N_7217,N_4882,N_4464);
xor U7218 (N_7218,N_3602,N_4151);
nand U7219 (N_7219,N_4380,N_5535);
xnor U7220 (N_7220,N_3114,N_4032);
nor U7221 (N_7221,N_3286,N_4904);
and U7222 (N_7222,N_4318,N_3056);
nor U7223 (N_7223,N_4056,N_4494);
or U7224 (N_7224,N_5397,N_4396);
or U7225 (N_7225,N_3813,N_5387);
or U7226 (N_7226,N_4479,N_5307);
or U7227 (N_7227,N_5324,N_4430);
xnor U7228 (N_7228,N_5165,N_4730);
nor U7229 (N_7229,N_4580,N_5098);
nand U7230 (N_7230,N_3173,N_5997);
nand U7231 (N_7231,N_4132,N_3139);
xor U7232 (N_7232,N_3610,N_5998);
or U7233 (N_7233,N_5681,N_4537);
and U7234 (N_7234,N_5710,N_4367);
nor U7235 (N_7235,N_5021,N_5218);
xnor U7236 (N_7236,N_4642,N_5029);
nor U7237 (N_7237,N_3577,N_3520);
and U7238 (N_7238,N_3593,N_5301);
nor U7239 (N_7239,N_4189,N_4739);
or U7240 (N_7240,N_5965,N_3151);
nand U7241 (N_7241,N_4545,N_5296);
or U7242 (N_7242,N_3084,N_5736);
and U7243 (N_7243,N_3536,N_5331);
nand U7244 (N_7244,N_5168,N_4675);
nor U7245 (N_7245,N_4866,N_4526);
xor U7246 (N_7246,N_4950,N_3783);
nand U7247 (N_7247,N_4337,N_4043);
nand U7248 (N_7248,N_3367,N_4643);
xor U7249 (N_7249,N_5492,N_4116);
and U7250 (N_7250,N_5388,N_3283);
and U7251 (N_7251,N_4432,N_3938);
nor U7252 (N_7252,N_5204,N_3085);
xnor U7253 (N_7253,N_4421,N_3741);
xor U7254 (N_7254,N_5055,N_5974);
and U7255 (N_7255,N_4017,N_4243);
nor U7256 (N_7256,N_3191,N_5412);
xor U7257 (N_7257,N_3373,N_4991);
or U7258 (N_7258,N_3100,N_4519);
or U7259 (N_7259,N_4948,N_4164);
nand U7260 (N_7260,N_5333,N_4727);
and U7261 (N_7261,N_3516,N_5708);
and U7262 (N_7262,N_3734,N_5215);
and U7263 (N_7263,N_4451,N_3771);
xnor U7264 (N_7264,N_5588,N_4835);
xnor U7265 (N_7265,N_3998,N_5194);
xnor U7266 (N_7266,N_5318,N_3153);
nor U7267 (N_7267,N_3023,N_3228);
nor U7268 (N_7268,N_3437,N_4431);
or U7269 (N_7269,N_5413,N_3158);
and U7270 (N_7270,N_5389,N_3246);
nor U7271 (N_7271,N_3518,N_3194);
xnor U7272 (N_7272,N_5674,N_4108);
nand U7273 (N_7273,N_5422,N_5119);
or U7274 (N_7274,N_3127,N_5580);
or U7275 (N_7275,N_4989,N_4001);
xor U7276 (N_7276,N_4443,N_5231);
and U7277 (N_7277,N_5510,N_3904);
nor U7278 (N_7278,N_3459,N_4145);
and U7279 (N_7279,N_3581,N_3534);
or U7280 (N_7280,N_5272,N_5222);
or U7281 (N_7281,N_5138,N_3776);
nand U7282 (N_7282,N_3175,N_4572);
nand U7283 (N_7283,N_5358,N_4713);
and U7284 (N_7284,N_3036,N_3708);
and U7285 (N_7285,N_5777,N_4311);
or U7286 (N_7286,N_5725,N_3368);
or U7287 (N_7287,N_5957,N_3422);
nand U7288 (N_7288,N_3440,N_3864);
nand U7289 (N_7289,N_5783,N_5423);
or U7290 (N_7290,N_3479,N_5709);
or U7291 (N_7291,N_3693,N_3123);
or U7292 (N_7292,N_4487,N_4414);
and U7293 (N_7293,N_4265,N_5427);
nand U7294 (N_7294,N_4118,N_3473);
nand U7295 (N_7295,N_4546,N_3852);
nand U7296 (N_7296,N_3428,N_5371);
xor U7297 (N_7297,N_4781,N_4617);
or U7298 (N_7298,N_3560,N_3635);
nor U7299 (N_7299,N_5035,N_5491);
or U7300 (N_7300,N_3526,N_3303);
or U7301 (N_7301,N_4695,N_4463);
xor U7302 (N_7302,N_4579,N_5461);
or U7303 (N_7303,N_4547,N_5752);
nor U7304 (N_7304,N_3359,N_3491);
or U7305 (N_7305,N_3381,N_4958);
or U7306 (N_7306,N_4930,N_3236);
xor U7307 (N_7307,N_3064,N_5608);
xor U7308 (N_7308,N_4450,N_3332);
xnor U7309 (N_7309,N_5597,N_5505);
xnor U7310 (N_7310,N_5270,N_4755);
and U7311 (N_7311,N_5360,N_4194);
or U7312 (N_7312,N_4749,N_5689);
and U7313 (N_7313,N_4423,N_4429);
nor U7314 (N_7314,N_3829,N_5378);
nor U7315 (N_7315,N_5010,N_5939);
and U7316 (N_7316,N_4936,N_5515);
nor U7317 (N_7317,N_4996,N_3206);
nand U7318 (N_7318,N_4836,N_4961);
nor U7319 (N_7319,N_5110,N_4880);
xor U7320 (N_7320,N_4665,N_5724);
or U7321 (N_7321,N_5981,N_5479);
and U7322 (N_7322,N_5529,N_3080);
and U7323 (N_7323,N_3795,N_3413);
xor U7324 (N_7324,N_5019,N_5472);
and U7325 (N_7325,N_5345,N_4041);
and U7326 (N_7326,N_4562,N_5649);
or U7327 (N_7327,N_5582,N_3052);
or U7328 (N_7328,N_4007,N_4865);
nor U7329 (N_7329,N_3910,N_3789);
nand U7330 (N_7330,N_3551,N_4274);
or U7331 (N_7331,N_5176,N_4878);
or U7332 (N_7332,N_3836,N_3698);
or U7333 (N_7333,N_4050,N_4543);
nor U7334 (N_7334,N_4532,N_4349);
nand U7335 (N_7335,N_4125,N_5250);
nand U7336 (N_7336,N_3674,N_3947);
xor U7337 (N_7337,N_4190,N_5922);
nor U7338 (N_7338,N_4073,N_4402);
xnor U7339 (N_7339,N_3269,N_3297);
or U7340 (N_7340,N_3567,N_3928);
xnor U7341 (N_7341,N_3476,N_5083);
or U7342 (N_7342,N_4312,N_5999);
nor U7343 (N_7343,N_4855,N_3773);
and U7344 (N_7344,N_3748,N_3584);
nand U7345 (N_7345,N_5103,N_3715);
xor U7346 (N_7346,N_5249,N_4536);
nand U7347 (N_7347,N_4965,N_4601);
and U7348 (N_7348,N_4682,N_5277);
nor U7349 (N_7349,N_4281,N_4117);
and U7350 (N_7350,N_4249,N_4575);
nand U7351 (N_7351,N_3845,N_3118);
nor U7352 (N_7352,N_3065,N_4703);
xor U7353 (N_7353,N_4608,N_5951);
xnor U7354 (N_7354,N_5379,N_3718);
xnor U7355 (N_7355,N_3233,N_3234);
or U7356 (N_7356,N_4676,N_3750);
and U7357 (N_7357,N_3775,N_3225);
nand U7358 (N_7358,N_5280,N_4213);
xor U7359 (N_7359,N_4686,N_3364);
or U7360 (N_7360,N_3110,N_3828);
xor U7361 (N_7361,N_3608,N_4474);
nor U7362 (N_7362,N_4453,N_3404);
nand U7363 (N_7363,N_3535,N_3519);
nand U7364 (N_7364,N_3680,N_5151);
and U7365 (N_7365,N_3411,N_3205);
nand U7366 (N_7366,N_4993,N_3805);
and U7367 (N_7367,N_3907,N_3021);
or U7368 (N_7368,N_3010,N_3620);
nor U7369 (N_7369,N_4245,N_4170);
nand U7370 (N_7370,N_5048,N_4977);
or U7371 (N_7371,N_3214,N_5308);
and U7372 (N_7372,N_5299,N_4824);
nand U7373 (N_7373,N_3985,N_5978);
xor U7374 (N_7374,N_5080,N_3573);
or U7375 (N_7375,N_4322,N_4469);
and U7376 (N_7376,N_5553,N_3082);
and U7377 (N_7377,N_4999,N_5791);
or U7378 (N_7378,N_3159,N_5276);
or U7379 (N_7379,N_5938,N_3227);
or U7380 (N_7380,N_4278,N_3249);
and U7381 (N_7381,N_3384,N_4114);
and U7382 (N_7382,N_3077,N_3006);
and U7383 (N_7383,N_4704,N_5366);
nand U7384 (N_7384,N_3441,N_3990);
nor U7385 (N_7385,N_3686,N_3556);
and U7386 (N_7386,N_4566,N_4485);
nand U7387 (N_7387,N_3856,N_3347);
or U7388 (N_7388,N_4497,N_5860);
xor U7389 (N_7389,N_5927,N_4387);
nor U7390 (N_7390,N_3574,N_3028);
xnor U7391 (N_7391,N_3024,N_3189);
nor U7392 (N_7392,N_3876,N_5134);
xnor U7393 (N_7393,N_3546,N_3730);
xnor U7394 (N_7394,N_5142,N_3544);
and U7395 (N_7395,N_4891,N_5409);
or U7396 (N_7396,N_5924,N_5571);
or U7397 (N_7397,N_3742,N_5171);
nor U7398 (N_7398,N_3887,N_4581);
or U7399 (N_7399,N_5960,N_3780);
nor U7400 (N_7400,N_3622,N_4234);
nor U7401 (N_7401,N_4171,N_5605);
xnor U7402 (N_7402,N_4748,N_3099);
nand U7403 (N_7403,N_5715,N_5631);
or U7404 (N_7404,N_4549,N_3529);
nor U7405 (N_7405,N_3237,N_3847);
nor U7406 (N_7406,N_5041,N_4728);
or U7407 (N_7407,N_4980,N_4747);
nor U7408 (N_7408,N_3324,N_4887);
nand U7409 (N_7409,N_4707,N_3355);
or U7410 (N_7410,N_5574,N_3960);
nand U7411 (N_7411,N_5056,N_3258);
or U7412 (N_7412,N_4079,N_5563);
xnor U7413 (N_7413,N_4037,N_4795);
and U7414 (N_7414,N_3195,N_5913);
nand U7415 (N_7415,N_5182,N_4788);
nor U7416 (N_7416,N_5696,N_5824);
or U7417 (N_7417,N_4096,N_3112);
xor U7418 (N_7418,N_4790,N_4291);
nand U7419 (N_7419,N_3071,N_4486);
xor U7420 (N_7420,N_3051,N_3659);
nand U7421 (N_7421,N_4741,N_5356);
nor U7422 (N_7422,N_5548,N_3462);
nand U7423 (N_7423,N_4408,N_5291);
xnor U7424 (N_7424,N_3348,N_5164);
nor U7425 (N_7425,N_4597,N_3745);
nand U7426 (N_7426,N_3890,N_3940);
xnor U7427 (N_7427,N_4535,N_4544);
nor U7428 (N_7428,N_3247,N_5867);
nand U7429 (N_7429,N_4074,N_3654);
nor U7430 (N_7430,N_5027,N_5050);
or U7431 (N_7431,N_5952,N_5376);
nand U7432 (N_7432,N_4673,N_4480);
nand U7433 (N_7433,N_5267,N_3296);
and U7434 (N_7434,N_5511,N_3204);
nand U7435 (N_7435,N_5986,N_5664);
and U7436 (N_7436,N_3352,N_3103);
xnor U7437 (N_7437,N_5682,N_3566);
xnor U7438 (N_7438,N_4576,N_3678);
or U7439 (N_7439,N_3005,N_3172);
nor U7440 (N_7440,N_5008,N_4342);
or U7441 (N_7441,N_5430,N_3585);
or U7442 (N_7442,N_3523,N_4095);
xor U7443 (N_7443,N_5850,N_4901);
nand U7444 (N_7444,N_5062,N_5882);
nand U7445 (N_7445,N_3765,N_4542);
xor U7446 (N_7446,N_4848,N_4301);
or U7447 (N_7447,N_4804,N_5522);
nor U7448 (N_7448,N_3253,N_3238);
or U7449 (N_7449,N_4452,N_4426);
xnor U7450 (N_7450,N_3496,N_4341);
nor U7451 (N_7451,N_5135,N_5895);
nor U7452 (N_7452,N_3814,N_4211);
nand U7453 (N_7453,N_3426,N_5635);
or U7454 (N_7454,N_4745,N_4702);
xor U7455 (N_7455,N_5097,N_4821);
nor U7456 (N_7456,N_5638,N_5380);
nor U7457 (N_7457,N_3463,N_5956);
nand U7458 (N_7458,N_5524,N_5024);
nor U7459 (N_7459,N_4971,N_5858);
or U7460 (N_7460,N_5130,N_3781);
or U7461 (N_7461,N_4082,N_5926);
xnor U7462 (N_7462,N_4216,N_4775);
xor U7463 (N_7463,N_5493,N_3881);
nand U7464 (N_7464,N_4927,N_4000);
nor U7465 (N_7465,N_3137,N_5617);
or U7466 (N_7466,N_4658,N_4215);
xnor U7467 (N_7467,N_4229,N_3090);
nand U7468 (N_7468,N_4881,N_4946);
xor U7469 (N_7469,N_5536,N_4684);
nor U7470 (N_7470,N_3315,N_3840);
nor U7471 (N_7471,N_3062,N_5298);
nor U7472 (N_7472,N_5191,N_3304);
and U7473 (N_7473,N_4994,N_3682);
and U7474 (N_7474,N_4491,N_5177);
nand U7475 (N_7475,N_5763,N_3792);
nand U7476 (N_7476,N_3731,N_5156);
xor U7477 (N_7477,N_3527,N_4837);
or U7478 (N_7478,N_4924,N_4529);
and U7479 (N_7479,N_3849,N_3029);
xnor U7480 (N_7480,N_3761,N_3211);
nor U7481 (N_7481,N_4089,N_4484);
nand U7482 (N_7482,N_4276,N_4382);
nor U7483 (N_7483,N_3611,N_5509);
or U7484 (N_7484,N_4298,N_4313);
xor U7485 (N_7485,N_4854,N_3639);
xnor U7486 (N_7486,N_5557,N_5052);
or U7487 (N_7487,N_3470,N_4078);
and U7488 (N_7488,N_4940,N_5026);
or U7489 (N_7489,N_5748,N_4551);
nand U7490 (N_7490,N_5235,N_3399);
and U7491 (N_7491,N_5162,N_5902);
xnor U7492 (N_7492,N_3392,N_5439);
xnor U7493 (N_7493,N_5589,N_3039);
and U7494 (N_7494,N_5116,N_4131);
xor U7495 (N_7495,N_4334,N_5793);
or U7496 (N_7496,N_4829,N_3207);
xor U7497 (N_7497,N_4246,N_5897);
and U7498 (N_7498,N_4232,N_5690);
and U7499 (N_7499,N_3086,N_3166);
and U7500 (N_7500,N_3447,N_5872);
and U7501 (N_7501,N_5749,N_3862);
xnor U7502 (N_7502,N_4075,N_5393);
nand U7503 (N_7503,N_3693,N_5698);
and U7504 (N_7504,N_3634,N_5028);
or U7505 (N_7505,N_3328,N_4137);
and U7506 (N_7506,N_3996,N_4052);
nand U7507 (N_7507,N_5966,N_4732);
nand U7508 (N_7508,N_4007,N_5247);
nor U7509 (N_7509,N_4234,N_3629);
or U7510 (N_7510,N_3404,N_5676);
nand U7511 (N_7511,N_5722,N_3685);
or U7512 (N_7512,N_5903,N_3871);
xnor U7513 (N_7513,N_5696,N_4938);
xor U7514 (N_7514,N_3681,N_4128);
nor U7515 (N_7515,N_3523,N_4447);
nand U7516 (N_7516,N_3288,N_3462);
nor U7517 (N_7517,N_4798,N_3322);
nor U7518 (N_7518,N_3041,N_4094);
or U7519 (N_7519,N_3473,N_4165);
nor U7520 (N_7520,N_4363,N_5441);
nor U7521 (N_7521,N_3761,N_4590);
nand U7522 (N_7522,N_3222,N_5925);
or U7523 (N_7523,N_3701,N_5886);
nor U7524 (N_7524,N_4832,N_4415);
or U7525 (N_7525,N_3818,N_4582);
nor U7526 (N_7526,N_5525,N_3483);
and U7527 (N_7527,N_5975,N_4475);
xor U7528 (N_7528,N_5631,N_3897);
and U7529 (N_7529,N_3789,N_3333);
nand U7530 (N_7530,N_4117,N_4857);
and U7531 (N_7531,N_5840,N_4153);
or U7532 (N_7532,N_5800,N_5424);
nor U7533 (N_7533,N_5494,N_4620);
or U7534 (N_7534,N_4397,N_3264);
nor U7535 (N_7535,N_5649,N_4076);
and U7536 (N_7536,N_4999,N_3895);
nand U7537 (N_7537,N_5108,N_4977);
nand U7538 (N_7538,N_3276,N_5187);
or U7539 (N_7539,N_5035,N_5885);
nor U7540 (N_7540,N_3555,N_5146);
or U7541 (N_7541,N_3708,N_5124);
nor U7542 (N_7542,N_5312,N_5765);
xnor U7543 (N_7543,N_4033,N_5738);
nand U7544 (N_7544,N_3937,N_4712);
nand U7545 (N_7545,N_4390,N_5103);
nand U7546 (N_7546,N_3545,N_5637);
nor U7547 (N_7547,N_3003,N_5690);
nand U7548 (N_7548,N_5757,N_4561);
and U7549 (N_7549,N_3250,N_4648);
or U7550 (N_7550,N_3495,N_3546);
nor U7551 (N_7551,N_5294,N_3017);
nor U7552 (N_7552,N_4594,N_3084);
or U7553 (N_7553,N_3645,N_5202);
nand U7554 (N_7554,N_4278,N_3742);
xor U7555 (N_7555,N_4744,N_5062);
nor U7556 (N_7556,N_4935,N_4906);
xor U7557 (N_7557,N_3799,N_3065);
nor U7558 (N_7558,N_4895,N_4603);
nand U7559 (N_7559,N_3718,N_3262);
nand U7560 (N_7560,N_5006,N_3766);
nand U7561 (N_7561,N_5731,N_3241);
and U7562 (N_7562,N_4476,N_4099);
nor U7563 (N_7563,N_3456,N_3338);
and U7564 (N_7564,N_5720,N_4882);
xor U7565 (N_7565,N_3344,N_3014);
nand U7566 (N_7566,N_4671,N_4013);
nor U7567 (N_7567,N_5954,N_5248);
nor U7568 (N_7568,N_4544,N_3620);
xor U7569 (N_7569,N_3701,N_4681);
and U7570 (N_7570,N_4634,N_3413);
nand U7571 (N_7571,N_5865,N_3508);
and U7572 (N_7572,N_5937,N_3461);
and U7573 (N_7573,N_4217,N_3381);
xnor U7574 (N_7574,N_5944,N_4442);
xnor U7575 (N_7575,N_4465,N_3763);
and U7576 (N_7576,N_3826,N_4068);
and U7577 (N_7577,N_4862,N_4641);
or U7578 (N_7578,N_4718,N_4094);
xnor U7579 (N_7579,N_3963,N_4059);
nand U7580 (N_7580,N_4526,N_3790);
or U7581 (N_7581,N_5802,N_3141);
nor U7582 (N_7582,N_5656,N_4585);
or U7583 (N_7583,N_5527,N_4117);
xnor U7584 (N_7584,N_3242,N_3640);
or U7585 (N_7585,N_3579,N_4709);
or U7586 (N_7586,N_4178,N_5760);
nand U7587 (N_7587,N_5861,N_5834);
or U7588 (N_7588,N_5153,N_4766);
nor U7589 (N_7589,N_4745,N_5424);
or U7590 (N_7590,N_3639,N_4041);
nor U7591 (N_7591,N_3351,N_4834);
or U7592 (N_7592,N_4554,N_3024);
xnor U7593 (N_7593,N_4518,N_4419);
or U7594 (N_7594,N_4442,N_3350);
nand U7595 (N_7595,N_3436,N_4964);
or U7596 (N_7596,N_4087,N_3955);
nor U7597 (N_7597,N_4387,N_4426);
xnor U7598 (N_7598,N_4055,N_5324);
nand U7599 (N_7599,N_3155,N_5380);
nor U7600 (N_7600,N_5528,N_4465);
or U7601 (N_7601,N_4725,N_5186);
nand U7602 (N_7602,N_5665,N_4097);
nand U7603 (N_7603,N_4243,N_5929);
nor U7604 (N_7604,N_4570,N_3691);
nand U7605 (N_7605,N_4912,N_3700);
xor U7606 (N_7606,N_5621,N_5829);
nand U7607 (N_7607,N_3891,N_3450);
nand U7608 (N_7608,N_5239,N_3243);
or U7609 (N_7609,N_3040,N_5334);
and U7610 (N_7610,N_4975,N_4131);
nand U7611 (N_7611,N_3453,N_4656);
xor U7612 (N_7612,N_3465,N_4801);
and U7613 (N_7613,N_4352,N_3654);
or U7614 (N_7614,N_3571,N_3756);
and U7615 (N_7615,N_5221,N_4039);
nand U7616 (N_7616,N_4440,N_5072);
and U7617 (N_7617,N_3036,N_3225);
and U7618 (N_7618,N_3199,N_5897);
xnor U7619 (N_7619,N_3342,N_5252);
or U7620 (N_7620,N_3766,N_5376);
and U7621 (N_7621,N_4349,N_5400);
nor U7622 (N_7622,N_4237,N_5216);
and U7623 (N_7623,N_4570,N_5377);
xnor U7624 (N_7624,N_3437,N_5616);
nor U7625 (N_7625,N_3255,N_5934);
nand U7626 (N_7626,N_5809,N_3162);
nand U7627 (N_7627,N_5065,N_3817);
and U7628 (N_7628,N_5936,N_5456);
nand U7629 (N_7629,N_5916,N_3290);
and U7630 (N_7630,N_4577,N_4829);
or U7631 (N_7631,N_4572,N_5343);
or U7632 (N_7632,N_5318,N_5254);
xnor U7633 (N_7633,N_4745,N_4256);
nor U7634 (N_7634,N_5672,N_5298);
or U7635 (N_7635,N_3306,N_3663);
nand U7636 (N_7636,N_5463,N_4465);
nor U7637 (N_7637,N_5080,N_5604);
xor U7638 (N_7638,N_4357,N_4136);
and U7639 (N_7639,N_4093,N_3221);
or U7640 (N_7640,N_3467,N_5831);
xnor U7641 (N_7641,N_3951,N_3489);
or U7642 (N_7642,N_5396,N_5732);
xor U7643 (N_7643,N_4793,N_3721);
nor U7644 (N_7644,N_4332,N_5910);
nor U7645 (N_7645,N_4472,N_5440);
nor U7646 (N_7646,N_4491,N_5306);
and U7647 (N_7647,N_5653,N_5994);
and U7648 (N_7648,N_4309,N_5384);
nor U7649 (N_7649,N_4295,N_5532);
and U7650 (N_7650,N_3466,N_5572);
or U7651 (N_7651,N_5337,N_4101);
nand U7652 (N_7652,N_3703,N_4331);
or U7653 (N_7653,N_4439,N_5142);
and U7654 (N_7654,N_4874,N_5015);
or U7655 (N_7655,N_3960,N_3009);
or U7656 (N_7656,N_5219,N_3824);
or U7657 (N_7657,N_5878,N_5651);
and U7658 (N_7658,N_3935,N_5814);
nand U7659 (N_7659,N_5395,N_3649);
nand U7660 (N_7660,N_4090,N_5041);
and U7661 (N_7661,N_4954,N_5073);
xor U7662 (N_7662,N_4986,N_5143);
and U7663 (N_7663,N_4795,N_4376);
or U7664 (N_7664,N_4011,N_5273);
nor U7665 (N_7665,N_3014,N_3518);
xnor U7666 (N_7666,N_4344,N_4649);
and U7667 (N_7667,N_3349,N_5884);
or U7668 (N_7668,N_3350,N_4045);
or U7669 (N_7669,N_4308,N_5617);
and U7670 (N_7670,N_4216,N_5772);
or U7671 (N_7671,N_4842,N_3894);
nand U7672 (N_7672,N_4723,N_5724);
and U7673 (N_7673,N_3794,N_4756);
or U7674 (N_7674,N_5807,N_3192);
and U7675 (N_7675,N_3359,N_3611);
or U7676 (N_7676,N_5592,N_4240);
nand U7677 (N_7677,N_5237,N_5840);
xor U7678 (N_7678,N_4955,N_5069);
and U7679 (N_7679,N_5946,N_3890);
nand U7680 (N_7680,N_4395,N_4428);
nor U7681 (N_7681,N_4968,N_5685);
nor U7682 (N_7682,N_3762,N_4854);
xnor U7683 (N_7683,N_3977,N_4090);
nor U7684 (N_7684,N_5338,N_3778);
and U7685 (N_7685,N_3339,N_3962);
nand U7686 (N_7686,N_4675,N_3427);
nand U7687 (N_7687,N_3010,N_3983);
or U7688 (N_7688,N_3673,N_5334);
nand U7689 (N_7689,N_3730,N_3560);
nor U7690 (N_7690,N_4779,N_5464);
and U7691 (N_7691,N_3525,N_3724);
and U7692 (N_7692,N_3957,N_4293);
or U7693 (N_7693,N_3197,N_4297);
nor U7694 (N_7694,N_4754,N_5449);
and U7695 (N_7695,N_4221,N_5472);
nand U7696 (N_7696,N_4723,N_3740);
and U7697 (N_7697,N_4434,N_5009);
and U7698 (N_7698,N_4048,N_4213);
xnor U7699 (N_7699,N_5500,N_3743);
xor U7700 (N_7700,N_4140,N_5618);
and U7701 (N_7701,N_5109,N_4469);
nand U7702 (N_7702,N_5878,N_4425);
nor U7703 (N_7703,N_3930,N_4395);
nor U7704 (N_7704,N_5724,N_3944);
nand U7705 (N_7705,N_5333,N_5951);
nor U7706 (N_7706,N_3715,N_5536);
xnor U7707 (N_7707,N_4431,N_5435);
or U7708 (N_7708,N_5148,N_5404);
or U7709 (N_7709,N_5090,N_3372);
nand U7710 (N_7710,N_4509,N_4401);
xor U7711 (N_7711,N_3458,N_5479);
or U7712 (N_7712,N_4787,N_3604);
or U7713 (N_7713,N_5535,N_4319);
or U7714 (N_7714,N_4624,N_3482);
and U7715 (N_7715,N_4981,N_4821);
xnor U7716 (N_7716,N_3608,N_5020);
or U7717 (N_7717,N_5902,N_4598);
and U7718 (N_7718,N_5667,N_3966);
xor U7719 (N_7719,N_5298,N_3100);
nand U7720 (N_7720,N_4165,N_4633);
nor U7721 (N_7721,N_3361,N_5274);
and U7722 (N_7722,N_4795,N_5055);
nor U7723 (N_7723,N_3832,N_5268);
nor U7724 (N_7724,N_5092,N_4048);
nand U7725 (N_7725,N_4569,N_5804);
and U7726 (N_7726,N_5960,N_4925);
and U7727 (N_7727,N_3398,N_4109);
nor U7728 (N_7728,N_3124,N_3932);
and U7729 (N_7729,N_4672,N_5024);
and U7730 (N_7730,N_5877,N_3486);
and U7731 (N_7731,N_4335,N_5878);
nor U7732 (N_7732,N_5019,N_4564);
nor U7733 (N_7733,N_4947,N_3460);
xor U7734 (N_7734,N_4352,N_3827);
xnor U7735 (N_7735,N_3922,N_3056);
nand U7736 (N_7736,N_5557,N_4652);
and U7737 (N_7737,N_3560,N_5962);
nand U7738 (N_7738,N_5705,N_4808);
xor U7739 (N_7739,N_3888,N_3341);
and U7740 (N_7740,N_3092,N_3438);
or U7741 (N_7741,N_4865,N_4878);
nor U7742 (N_7742,N_4400,N_5562);
and U7743 (N_7743,N_5543,N_4157);
and U7744 (N_7744,N_5417,N_3148);
or U7745 (N_7745,N_5751,N_4186);
xor U7746 (N_7746,N_4344,N_4571);
and U7747 (N_7747,N_5815,N_5051);
xor U7748 (N_7748,N_4948,N_4912);
nor U7749 (N_7749,N_5904,N_4904);
nor U7750 (N_7750,N_5642,N_3275);
or U7751 (N_7751,N_5843,N_4697);
and U7752 (N_7752,N_5446,N_4938);
xnor U7753 (N_7753,N_5987,N_3968);
and U7754 (N_7754,N_5353,N_3497);
nor U7755 (N_7755,N_3357,N_3969);
nor U7756 (N_7756,N_4399,N_5103);
nand U7757 (N_7757,N_5182,N_5102);
nor U7758 (N_7758,N_5820,N_5666);
and U7759 (N_7759,N_5004,N_3112);
nor U7760 (N_7760,N_4815,N_5859);
or U7761 (N_7761,N_5863,N_3314);
nor U7762 (N_7762,N_5740,N_5106);
nand U7763 (N_7763,N_5601,N_5319);
or U7764 (N_7764,N_3644,N_3255);
nor U7765 (N_7765,N_5313,N_4902);
nor U7766 (N_7766,N_3462,N_4473);
nor U7767 (N_7767,N_5961,N_3534);
xnor U7768 (N_7768,N_3605,N_4901);
nor U7769 (N_7769,N_3496,N_5893);
nand U7770 (N_7770,N_3890,N_4331);
nand U7771 (N_7771,N_5327,N_4979);
and U7772 (N_7772,N_5806,N_5564);
nor U7773 (N_7773,N_5159,N_3035);
or U7774 (N_7774,N_5817,N_3580);
xor U7775 (N_7775,N_3119,N_3390);
xnor U7776 (N_7776,N_5946,N_4038);
or U7777 (N_7777,N_3821,N_3769);
xnor U7778 (N_7778,N_5131,N_4870);
and U7779 (N_7779,N_5215,N_5289);
xor U7780 (N_7780,N_3960,N_5299);
or U7781 (N_7781,N_4631,N_4398);
and U7782 (N_7782,N_3395,N_5674);
and U7783 (N_7783,N_3850,N_5710);
nand U7784 (N_7784,N_3761,N_4453);
nor U7785 (N_7785,N_3350,N_3047);
or U7786 (N_7786,N_4256,N_5372);
and U7787 (N_7787,N_4707,N_3412);
or U7788 (N_7788,N_3241,N_4934);
nor U7789 (N_7789,N_3459,N_4478);
nor U7790 (N_7790,N_5914,N_5181);
or U7791 (N_7791,N_3360,N_5422);
nor U7792 (N_7792,N_5799,N_4261);
nor U7793 (N_7793,N_4673,N_3932);
nand U7794 (N_7794,N_5608,N_4435);
nor U7795 (N_7795,N_3756,N_3633);
or U7796 (N_7796,N_4150,N_4854);
xnor U7797 (N_7797,N_3979,N_4978);
nor U7798 (N_7798,N_5328,N_3733);
nand U7799 (N_7799,N_5310,N_3396);
xor U7800 (N_7800,N_3668,N_5250);
and U7801 (N_7801,N_5489,N_5575);
or U7802 (N_7802,N_4068,N_5205);
nand U7803 (N_7803,N_3444,N_3301);
and U7804 (N_7804,N_5246,N_5955);
xor U7805 (N_7805,N_4152,N_4272);
or U7806 (N_7806,N_4270,N_3689);
nor U7807 (N_7807,N_5528,N_5565);
nand U7808 (N_7808,N_4443,N_3889);
or U7809 (N_7809,N_3088,N_5346);
nand U7810 (N_7810,N_3169,N_3443);
nand U7811 (N_7811,N_3275,N_5887);
and U7812 (N_7812,N_5017,N_3765);
nor U7813 (N_7813,N_3578,N_3984);
xnor U7814 (N_7814,N_5401,N_3385);
xnor U7815 (N_7815,N_3316,N_3423);
or U7816 (N_7816,N_5998,N_5668);
nor U7817 (N_7817,N_3538,N_4397);
nand U7818 (N_7818,N_4627,N_4282);
xnor U7819 (N_7819,N_4947,N_5964);
and U7820 (N_7820,N_5323,N_3578);
and U7821 (N_7821,N_4066,N_4888);
xnor U7822 (N_7822,N_3282,N_5943);
or U7823 (N_7823,N_3593,N_5628);
and U7824 (N_7824,N_4734,N_4097);
nand U7825 (N_7825,N_4845,N_4182);
nor U7826 (N_7826,N_5360,N_5418);
and U7827 (N_7827,N_4454,N_4328);
or U7828 (N_7828,N_3638,N_3208);
or U7829 (N_7829,N_5012,N_3530);
nand U7830 (N_7830,N_4810,N_4456);
nor U7831 (N_7831,N_5147,N_5730);
xor U7832 (N_7832,N_4072,N_4465);
or U7833 (N_7833,N_4950,N_3047);
and U7834 (N_7834,N_4397,N_4753);
xor U7835 (N_7835,N_4377,N_5471);
nor U7836 (N_7836,N_4294,N_4926);
nor U7837 (N_7837,N_5698,N_5101);
nor U7838 (N_7838,N_3008,N_4009);
or U7839 (N_7839,N_4376,N_4462);
xor U7840 (N_7840,N_4200,N_5471);
xor U7841 (N_7841,N_4642,N_5480);
and U7842 (N_7842,N_5600,N_3051);
or U7843 (N_7843,N_4530,N_5589);
or U7844 (N_7844,N_4671,N_5737);
nand U7845 (N_7845,N_4336,N_5323);
and U7846 (N_7846,N_3358,N_4744);
nor U7847 (N_7847,N_4440,N_4493);
nor U7848 (N_7848,N_4110,N_5617);
xnor U7849 (N_7849,N_4180,N_3432);
nand U7850 (N_7850,N_3409,N_5484);
nor U7851 (N_7851,N_4258,N_4298);
nand U7852 (N_7852,N_5946,N_5943);
nor U7853 (N_7853,N_5567,N_5315);
or U7854 (N_7854,N_4070,N_5642);
and U7855 (N_7855,N_5355,N_3855);
or U7856 (N_7856,N_4082,N_4222);
xor U7857 (N_7857,N_5431,N_5149);
or U7858 (N_7858,N_5108,N_4716);
nor U7859 (N_7859,N_4735,N_5152);
nand U7860 (N_7860,N_4250,N_5088);
nor U7861 (N_7861,N_4904,N_3514);
xnor U7862 (N_7862,N_5767,N_3406);
nor U7863 (N_7863,N_3435,N_5458);
nor U7864 (N_7864,N_5220,N_4567);
nor U7865 (N_7865,N_5095,N_4441);
and U7866 (N_7866,N_5743,N_3913);
and U7867 (N_7867,N_5779,N_3623);
nor U7868 (N_7868,N_5285,N_4714);
or U7869 (N_7869,N_3043,N_4527);
xor U7870 (N_7870,N_4018,N_4646);
xnor U7871 (N_7871,N_5479,N_4115);
and U7872 (N_7872,N_5513,N_3844);
nor U7873 (N_7873,N_5241,N_3450);
nand U7874 (N_7874,N_3055,N_5247);
nor U7875 (N_7875,N_3270,N_5734);
and U7876 (N_7876,N_4558,N_5224);
or U7877 (N_7877,N_5616,N_4140);
and U7878 (N_7878,N_5548,N_3918);
nand U7879 (N_7879,N_4224,N_3865);
nor U7880 (N_7880,N_3806,N_5015);
nand U7881 (N_7881,N_5924,N_5128);
nor U7882 (N_7882,N_5318,N_3504);
xnor U7883 (N_7883,N_5113,N_5566);
nor U7884 (N_7884,N_4153,N_4280);
and U7885 (N_7885,N_3103,N_3441);
nand U7886 (N_7886,N_5094,N_3797);
nor U7887 (N_7887,N_4671,N_3029);
xor U7888 (N_7888,N_3048,N_5862);
nand U7889 (N_7889,N_4516,N_5463);
nand U7890 (N_7890,N_5982,N_5593);
or U7891 (N_7891,N_3552,N_5920);
xnor U7892 (N_7892,N_5415,N_5744);
nand U7893 (N_7893,N_4358,N_4008);
nor U7894 (N_7894,N_5951,N_3392);
nand U7895 (N_7895,N_4385,N_3644);
nand U7896 (N_7896,N_3887,N_4170);
or U7897 (N_7897,N_3624,N_5041);
xnor U7898 (N_7898,N_4050,N_5547);
xor U7899 (N_7899,N_5875,N_4829);
or U7900 (N_7900,N_5338,N_5931);
nand U7901 (N_7901,N_3186,N_5906);
xnor U7902 (N_7902,N_3051,N_3283);
and U7903 (N_7903,N_4136,N_3295);
nand U7904 (N_7904,N_4031,N_3886);
and U7905 (N_7905,N_5905,N_3733);
or U7906 (N_7906,N_4476,N_3502);
or U7907 (N_7907,N_5735,N_3125);
nand U7908 (N_7908,N_5232,N_5812);
or U7909 (N_7909,N_5863,N_3873);
nand U7910 (N_7910,N_4302,N_3601);
nand U7911 (N_7911,N_4865,N_5495);
nor U7912 (N_7912,N_5298,N_4135);
nand U7913 (N_7913,N_4058,N_5095);
xnor U7914 (N_7914,N_5649,N_4212);
or U7915 (N_7915,N_4536,N_5568);
or U7916 (N_7916,N_5571,N_4998);
or U7917 (N_7917,N_5614,N_5033);
nor U7918 (N_7918,N_3494,N_5116);
or U7919 (N_7919,N_3857,N_3407);
nor U7920 (N_7920,N_5158,N_4605);
nand U7921 (N_7921,N_3482,N_5098);
and U7922 (N_7922,N_5911,N_3800);
xnor U7923 (N_7923,N_3156,N_5967);
nand U7924 (N_7924,N_3020,N_5645);
nor U7925 (N_7925,N_4331,N_3317);
xnor U7926 (N_7926,N_4816,N_5979);
and U7927 (N_7927,N_3094,N_5466);
xor U7928 (N_7928,N_4038,N_5458);
nand U7929 (N_7929,N_4357,N_4699);
xor U7930 (N_7930,N_5396,N_4398);
nand U7931 (N_7931,N_3171,N_3706);
and U7932 (N_7932,N_4485,N_4479);
nor U7933 (N_7933,N_3961,N_3521);
or U7934 (N_7934,N_4219,N_3759);
xnor U7935 (N_7935,N_5350,N_5057);
nor U7936 (N_7936,N_5343,N_5401);
or U7937 (N_7937,N_3478,N_4614);
or U7938 (N_7938,N_5138,N_4341);
xnor U7939 (N_7939,N_4185,N_4369);
and U7940 (N_7940,N_4719,N_3914);
nand U7941 (N_7941,N_5117,N_5693);
nand U7942 (N_7942,N_4356,N_5566);
or U7943 (N_7943,N_3257,N_3816);
and U7944 (N_7944,N_5270,N_5087);
nor U7945 (N_7945,N_3014,N_5214);
nor U7946 (N_7946,N_3700,N_4471);
nor U7947 (N_7947,N_3056,N_3674);
and U7948 (N_7948,N_5936,N_4220);
or U7949 (N_7949,N_5139,N_3948);
nand U7950 (N_7950,N_4303,N_4515);
nor U7951 (N_7951,N_5360,N_5557);
xnor U7952 (N_7952,N_4252,N_3754);
nand U7953 (N_7953,N_5747,N_5899);
nand U7954 (N_7954,N_4628,N_3225);
nor U7955 (N_7955,N_5974,N_3101);
or U7956 (N_7956,N_5612,N_3222);
or U7957 (N_7957,N_3426,N_3903);
nor U7958 (N_7958,N_5035,N_4803);
and U7959 (N_7959,N_5727,N_3780);
and U7960 (N_7960,N_5015,N_5768);
or U7961 (N_7961,N_5976,N_3965);
or U7962 (N_7962,N_5542,N_5996);
nand U7963 (N_7963,N_3846,N_3180);
and U7964 (N_7964,N_5170,N_4343);
and U7965 (N_7965,N_3391,N_4934);
nand U7966 (N_7966,N_5673,N_4420);
xnor U7967 (N_7967,N_5542,N_3486);
or U7968 (N_7968,N_4716,N_4433);
or U7969 (N_7969,N_5494,N_5287);
and U7970 (N_7970,N_5075,N_4955);
nor U7971 (N_7971,N_3935,N_5522);
nor U7972 (N_7972,N_4698,N_4576);
nor U7973 (N_7973,N_4431,N_3502);
nor U7974 (N_7974,N_5679,N_5846);
xnor U7975 (N_7975,N_4512,N_4919);
and U7976 (N_7976,N_3811,N_3550);
xnor U7977 (N_7977,N_5679,N_5933);
nand U7978 (N_7978,N_5701,N_3581);
nand U7979 (N_7979,N_5410,N_3607);
nor U7980 (N_7980,N_5344,N_3724);
xor U7981 (N_7981,N_4278,N_4143);
nor U7982 (N_7982,N_5339,N_3796);
and U7983 (N_7983,N_4612,N_5781);
and U7984 (N_7984,N_4855,N_4647);
xor U7985 (N_7985,N_4735,N_3634);
or U7986 (N_7986,N_5548,N_5376);
and U7987 (N_7987,N_5606,N_3936);
or U7988 (N_7988,N_3065,N_5432);
nand U7989 (N_7989,N_3039,N_4265);
nor U7990 (N_7990,N_3012,N_5362);
xor U7991 (N_7991,N_3843,N_4414);
xor U7992 (N_7992,N_4698,N_5003);
xor U7993 (N_7993,N_4597,N_5275);
xor U7994 (N_7994,N_3775,N_5335);
nand U7995 (N_7995,N_5302,N_3433);
xor U7996 (N_7996,N_3651,N_4955);
nand U7997 (N_7997,N_5210,N_5024);
nand U7998 (N_7998,N_3347,N_3092);
or U7999 (N_7999,N_4418,N_5892);
nor U8000 (N_8000,N_5009,N_4078);
nand U8001 (N_8001,N_5636,N_4604);
or U8002 (N_8002,N_3352,N_5998);
and U8003 (N_8003,N_5239,N_3048);
xnor U8004 (N_8004,N_4229,N_5222);
nand U8005 (N_8005,N_5770,N_5356);
nand U8006 (N_8006,N_5161,N_4772);
nand U8007 (N_8007,N_4768,N_5437);
and U8008 (N_8008,N_4669,N_5612);
or U8009 (N_8009,N_4889,N_4649);
nand U8010 (N_8010,N_3306,N_3760);
nand U8011 (N_8011,N_5254,N_4921);
and U8012 (N_8012,N_5569,N_3027);
and U8013 (N_8013,N_3252,N_4731);
nor U8014 (N_8014,N_3060,N_5585);
nor U8015 (N_8015,N_5346,N_3445);
xnor U8016 (N_8016,N_5627,N_3796);
or U8017 (N_8017,N_4928,N_3003);
or U8018 (N_8018,N_4624,N_4943);
nor U8019 (N_8019,N_5048,N_5641);
xnor U8020 (N_8020,N_4486,N_5673);
nor U8021 (N_8021,N_5093,N_5881);
nor U8022 (N_8022,N_3462,N_5549);
nand U8023 (N_8023,N_3469,N_5204);
and U8024 (N_8024,N_3197,N_3747);
or U8025 (N_8025,N_3274,N_5092);
nor U8026 (N_8026,N_5520,N_5858);
nand U8027 (N_8027,N_3658,N_4608);
xor U8028 (N_8028,N_3865,N_3396);
xnor U8029 (N_8029,N_5477,N_5720);
and U8030 (N_8030,N_4520,N_3515);
nor U8031 (N_8031,N_3911,N_4969);
xnor U8032 (N_8032,N_4736,N_3224);
and U8033 (N_8033,N_3512,N_4660);
or U8034 (N_8034,N_3465,N_4790);
nand U8035 (N_8035,N_5075,N_3821);
and U8036 (N_8036,N_3693,N_3740);
or U8037 (N_8037,N_3024,N_3904);
or U8038 (N_8038,N_5448,N_3043);
xor U8039 (N_8039,N_4853,N_5394);
or U8040 (N_8040,N_5892,N_5352);
nor U8041 (N_8041,N_4315,N_3573);
xor U8042 (N_8042,N_3076,N_5760);
and U8043 (N_8043,N_5341,N_4466);
nor U8044 (N_8044,N_4356,N_4903);
or U8045 (N_8045,N_3072,N_5182);
xor U8046 (N_8046,N_5138,N_4007);
nand U8047 (N_8047,N_4576,N_4407);
nor U8048 (N_8048,N_5019,N_3205);
and U8049 (N_8049,N_3628,N_3361);
nand U8050 (N_8050,N_5359,N_3630);
nor U8051 (N_8051,N_5511,N_3061);
xor U8052 (N_8052,N_3899,N_4670);
or U8053 (N_8053,N_4870,N_4909);
nand U8054 (N_8054,N_5534,N_5252);
and U8055 (N_8055,N_3257,N_5559);
xnor U8056 (N_8056,N_5822,N_3035);
or U8057 (N_8057,N_5118,N_5032);
or U8058 (N_8058,N_5365,N_4808);
and U8059 (N_8059,N_5305,N_3756);
nand U8060 (N_8060,N_4712,N_3757);
nand U8061 (N_8061,N_4081,N_5492);
nor U8062 (N_8062,N_4620,N_3039);
nand U8063 (N_8063,N_5951,N_5287);
nor U8064 (N_8064,N_5001,N_5403);
nand U8065 (N_8065,N_3998,N_5966);
nor U8066 (N_8066,N_5750,N_3605);
and U8067 (N_8067,N_4974,N_3136);
and U8068 (N_8068,N_5945,N_3423);
and U8069 (N_8069,N_5267,N_3224);
xnor U8070 (N_8070,N_4836,N_5998);
xnor U8071 (N_8071,N_3416,N_4897);
xnor U8072 (N_8072,N_3649,N_5414);
nand U8073 (N_8073,N_5729,N_5687);
and U8074 (N_8074,N_5584,N_3519);
nand U8075 (N_8075,N_3714,N_3798);
xnor U8076 (N_8076,N_5919,N_3614);
and U8077 (N_8077,N_5192,N_5597);
xnor U8078 (N_8078,N_5614,N_4018);
or U8079 (N_8079,N_4435,N_4509);
nand U8080 (N_8080,N_4209,N_5818);
and U8081 (N_8081,N_5350,N_4147);
xor U8082 (N_8082,N_5093,N_5446);
nor U8083 (N_8083,N_4387,N_3878);
and U8084 (N_8084,N_4376,N_3045);
nor U8085 (N_8085,N_4926,N_4681);
nor U8086 (N_8086,N_5856,N_3279);
and U8087 (N_8087,N_3614,N_3135);
and U8088 (N_8088,N_4378,N_3985);
or U8089 (N_8089,N_3933,N_4480);
nand U8090 (N_8090,N_4634,N_5978);
or U8091 (N_8091,N_5277,N_4175);
nor U8092 (N_8092,N_4590,N_4169);
and U8093 (N_8093,N_4296,N_5390);
or U8094 (N_8094,N_4733,N_3210);
nand U8095 (N_8095,N_4367,N_5199);
and U8096 (N_8096,N_5909,N_3248);
xor U8097 (N_8097,N_4905,N_4511);
or U8098 (N_8098,N_4444,N_4406);
or U8099 (N_8099,N_4833,N_5566);
xnor U8100 (N_8100,N_4482,N_5263);
or U8101 (N_8101,N_4446,N_5222);
or U8102 (N_8102,N_4725,N_5134);
nand U8103 (N_8103,N_5495,N_4883);
or U8104 (N_8104,N_5201,N_4335);
nor U8105 (N_8105,N_5940,N_5611);
and U8106 (N_8106,N_3167,N_4043);
and U8107 (N_8107,N_4202,N_4992);
nor U8108 (N_8108,N_4634,N_3320);
nand U8109 (N_8109,N_5743,N_3858);
nand U8110 (N_8110,N_5434,N_5415);
nand U8111 (N_8111,N_4325,N_4879);
nor U8112 (N_8112,N_5323,N_5334);
nand U8113 (N_8113,N_3797,N_4806);
or U8114 (N_8114,N_4840,N_4414);
nor U8115 (N_8115,N_4175,N_3476);
and U8116 (N_8116,N_5200,N_3600);
nand U8117 (N_8117,N_4609,N_3661);
xor U8118 (N_8118,N_4656,N_5739);
nor U8119 (N_8119,N_3892,N_3216);
xnor U8120 (N_8120,N_3759,N_4390);
and U8121 (N_8121,N_5911,N_3391);
nor U8122 (N_8122,N_4514,N_4150);
or U8123 (N_8123,N_4984,N_4492);
nor U8124 (N_8124,N_4600,N_3969);
nand U8125 (N_8125,N_4213,N_3529);
nor U8126 (N_8126,N_5517,N_4810);
or U8127 (N_8127,N_5069,N_4361);
nand U8128 (N_8128,N_4124,N_3727);
nor U8129 (N_8129,N_5844,N_3872);
xor U8130 (N_8130,N_4987,N_5375);
xor U8131 (N_8131,N_3356,N_5160);
or U8132 (N_8132,N_4808,N_3184);
or U8133 (N_8133,N_3410,N_5150);
nor U8134 (N_8134,N_5412,N_5959);
and U8135 (N_8135,N_3273,N_3840);
or U8136 (N_8136,N_5765,N_5453);
nor U8137 (N_8137,N_5788,N_4309);
nor U8138 (N_8138,N_5763,N_4412);
nand U8139 (N_8139,N_3746,N_4602);
and U8140 (N_8140,N_4435,N_5172);
or U8141 (N_8141,N_5232,N_5768);
or U8142 (N_8142,N_3265,N_3299);
or U8143 (N_8143,N_4145,N_5430);
or U8144 (N_8144,N_3083,N_3618);
xor U8145 (N_8145,N_5969,N_4740);
nand U8146 (N_8146,N_4171,N_4206);
nor U8147 (N_8147,N_3929,N_5071);
nand U8148 (N_8148,N_5734,N_5390);
and U8149 (N_8149,N_5461,N_4843);
or U8150 (N_8150,N_4514,N_4467);
xnor U8151 (N_8151,N_5455,N_4150);
nand U8152 (N_8152,N_5417,N_5729);
nor U8153 (N_8153,N_4439,N_5792);
and U8154 (N_8154,N_4823,N_5299);
nor U8155 (N_8155,N_3272,N_4125);
and U8156 (N_8156,N_3959,N_3949);
nor U8157 (N_8157,N_4025,N_5070);
xor U8158 (N_8158,N_5687,N_3101);
xnor U8159 (N_8159,N_5979,N_3463);
nand U8160 (N_8160,N_3920,N_5835);
xnor U8161 (N_8161,N_5011,N_3231);
nor U8162 (N_8162,N_3649,N_3169);
nand U8163 (N_8163,N_4667,N_4356);
or U8164 (N_8164,N_4324,N_3318);
xnor U8165 (N_8165,N_4257,N_4848);
xnor U8166 (N_8166,N_3864,N_4357);
xor U8167 (N_8167,N_5134,N_5882);
nor U8168 (N_8168,N_3900,N_3574);
and U8169 (N_8169,N_5892,N_4941);
and U8170 (N_8170,N_3797,N_4640);
and U8171 (N_8171,N_5832,N_4582);
xnor U8172 (N_8172,N_3550,N_3202);
nand U8173 (N_8173,N_4610,N_3099);
or U8174 (N_8174,N_4013,N_5096);
and U8175 (N_8175,N_3930,N_4935);
nor U8176 (N_8176,N_3373,N_5338);
or U8177 (N_8177,N_5836,N_3125);
nor U8178 (N_8178,N_4698,N_5671);
nand U8179 (N_8179,N_5566,N_5774);
or U8180 (N_8180,N_3912,N_4965);
nor U8181 (N_8181,N_5748,N_5326);
or U8182 (N_8182,N_4644,N_5558);
nand U8183 (N_8183,N_5970,N_4643);
nand U8184 (N_8184,N_4245,N_5427);
nor U8185 (N_8185,N_3722,N_4565);
xnor U8186 (N_8186,N_3150,N_5289);
and U8187 (N_8187,N_4561,N_4338);
xnor U8188 (N_8188,N_4705,N_3720);
nand U8189 (N_8189,N_5903,N_5369);
and U8190 (N_8190,N_4826,N_4116);
nand U8191 (N_8191,N_4785,N_3053);
nor U8192 (N_8192,N_5510,N_5493);
or U8193 (N_8193,N_3198,N_3117);
and U8194 (N_8194,N_5589,N_4617);
nand U8195 (N_8195,N_3735,N_5387);
xnor U8196 (N_8196,N_3396,N_5389);
xnor U8197 (N_8197,N_3895,N_5342);
nor U8198 (N_8198,N_3234,N_5799);
xnor U8199 (N_8199,N_4215,N_4797);
and U8200 (N_8200,N_5483,N_5778);
and U8201 (N_8201,N_5693,N_5384);
nand U8202 (N_8202,N_3547,N_5196);
and U8203 (N_8203,N_3130,N_5717);
nand U8204 (N_8204,N_4892,N_5057);
or U8205 (N_8205,N_3675,N_4587);
and U8206 (N_8206,N_4927,N_3379);
and U8207 (N_8207,N_3531,N_3769);
nor U8208 (N_8208,N_3853,N_4784);
xnor U8209 (N_8209,N_4838,N_5456);
nand U8210 (N_8210,N_4390,N_3287);
or U8211 (N_8211,N_5454,N_5933);
or U8212 (N_8212,N_3569,N_3298);
or U8213 (N_8213,N_5444,N_3892);
nor U8214 (N_8214,N_5671,N_5166);
or U8215 (N_8215,N_5130,N_5007);
xnor U8216 (N_8216,N_4002,N_4549);
and U8217 (N_8217,N_4969,N_5290);
or U8218 (N_8218,N_4799,N_4073);
nor U8219 (N_8219,N_4623,N_3501);
nor U8220 (N_8220,N_3512,N_5302);
nand U8221 (N_8221,N_5330,N_3192);
and U8222 (N_8222,N_5574,N_3892);
or U8223 (N_8223,N_3992,N_4225);
nand U8224 (N_8224,N_5926,N_3630);
nand U8225 (N_8225,N_5175,N_5523);
and U8226 (N_8226,N_3956,N_3326);
or U8227 (N_8227,N_4574,N_5137);
xor U8228 (N_8228,N_3651,N_3739);
nand U8229 (N_8229,N_5131,N_5066);
and U8230 (N_8230,N_5316,N_5429);
nor U8231 (N_8231,N_4599,N_3446);
or U8232 (N_8232,N_3537,N_3398);
and U8233 (N_8233,N_5660,N_3973);
and U8234 (N_8234,N_4542,N_4591);
and U8235 (N_8235,N_5151,N_5760);
nand U8236 (N_8236,N_3076,N_4415);
nand U8237 (N_8237,N_5474,N_3984);
nand U8238 (N_8238,N_4058,N_3949);
or U8239 (N_8239,N_3977,N_4210);
and U8240 (N_8240,N_4092,N_3466);
or U8241 (N_8241,N_5491,N_5831);
nand U8242 (N_8242,N_3497,N_3389);
nand U8243 (N_8243,N_3199,N_5199);
nand U8244 (N_8244,N_5214,N_3798);
and U8245 (N_8245,N_4939,N_3992);
nor U8246 (N_8246,N_5359,N_4046);
nand U8247 (N_8247,N_3869,N_5728);
and U8248 (N_8248,N_4745,N_4214);
nor U8249 (N_8249,N_5716,N_5401);
and U8250 (N_8250,N_5959,N_3954);
nor U8251 (N_8251,N_4196,N_4981);
xor U8252 (N_8252,N_3188,N_3201);
xor U8253 (N_8253,N_3778,N_3829);
nand U8254 (N_8254,N_4052,N_4933);
or U8255 (N_8255,N_3664,N_3989);
nand U8256 (N_8256,N_5189,N_3157);
and U8257 (N_8257,N_3531,N_5013);
and U8258 (N_8258,N_3632,N_5324);
or U8259 (N_8259,N_5302,N_4198);
nand U8260 (N_8260,N_4296,N_5086);
xor U8261 (N_8261,N_3883,N_4421);
or U8262 (N_8262,N_5883,N_5605);
or U8263 (N_8263,N_5074,N_4445);
nor U8264 (N_8264,N_5999,N_5466);
and U8265 (N_8265,N_5910,N_3556);
or U8266 (N_8266,N_5020,N_3890);
and U8267 (N_8267,N_4607,N_4470);
or U8268 (N_8268,N_3626,N_5014);
nand U8269 (N_8269,N_5935,N_5204);
and U8270 (N_8270,N_4834,N_5625);
nor U8271 (N_8271,N_3606,N_5567);
xnor U8272 (N_8272,N_3995,N_5330);
or U8273 (N_8273,N_3334,N_5966);
nor U8274 (N_8274,N_4754,N_5537);
or U8275 (N_8275,N_5996,N_3803);
or U8276 (N_8276,N_3155,N_4439);
and U8277 (N_8277,N_4103,N_3611);
xor U8278 (N_8278,N_5382,N_4661);
and U8279 (N_8279,N_4490,N_3450);
xor U8280 (N_8280,N_4790,N_4606);
and U8281 (N_8281,N_3447,N_3116);
or U8282 (N_8282,N_3555,N_4483);
and U8283 (N_8283,N_4698,N_4136);
and U8284 (N_8284,N_5429,N_5440);
xor U8285 (N_8285,N_5855,N_3272);
and U8286 (N_8286,N_4887,N_3228);
xnor U8287 (N_8287,N_4288,N_3539);
nand U8288 (N_8288,N_5990,N_5875);
nor U8289 (N_8289,N_4043,N_3931);
xnor U8290 (N_8290,N_3276,N_3358);
and U8291 (N_8291,N_4856,N_3326);
xor U8292 (N_8292,N_4291,N_4725);
xor U8293 (N_8293,N_3240,N_4397);
nand U8294 (N_8294,N_3467,N_3776);
or U8295 (N_8295,N_5196,N_4192);
or U8296 (N_8296,N_3995,N_5462);
nor U8297 (N_8297,N_4097,N_3276);
or U8298 (N_8298,N_5712,N_4184);
and U8299 (N_8299,N_5930,N_4117);
and U8300 (N_8300,N_3489,N_3816);
xnor U8301 (N_8301,N_4973,N_4746);
and U8302 (N_8302,N_5547,N_5392);
and U8303 (N_8303,N_3956,N_4938);
nand U8304 (N_8304,N_5713,N_4426);
or U8305 (N_8305,N_4605,N_4153);
xor U8306 (N_8306,N_5743,N_5595);
and U8307 (N_8307,N_5333,N_3838);
xnor U8308 (N_8308,N_5227,N_4196);
and U8309 (N_8309,N_3500,N_3174);
nor U8310 (N_8310,N_5140,N_3876);
nor U8311 (N_8311,N_4640,N_5660);
or U8312 (N_8312,N_4979,N_4429);
nand U8313 (N_8313,N_5674,N_3615);
nor U8314 (N_8314,N_4828,N_5771);
or U8315 (N_8315,N_5209,N_5825);
or U8316 (N_8316,N_5917,N_3431);
or U8317 (N_8317,N_4474,N_5059);
nand U8318 (N_8318,N_3731,N_5883);
or U8319 (N_8319,N_5863,N_5562);
xor U8320 (N_8320,N_5704,N_4837);
nor U8321 (N_8321,N_3633,N_4303);
xor U8322 (N_8322,N_5703,N_3597);
nor U8323 (N_8323,N_4773,N_5360);
nand U8324 (N_8324,N_5511,N_5045);
nor U8325 (N_8325,N_5408,N_4592);
nand U8326 (N_8326,N_5047,N_3059);
xnor U8327 (N_8327,N_4476,N_3389);
nor U8328 (N_8328,N_3579,N_5808);
xor U8329 (N_8329,N_5290,N_3088);
or U8330 (N_8330,N_3949,N_5523);
nand U8331 (N_8331,N_5865,N_5991);
nor U8332 (N_8332,N_4459,N_5981);
or U8333 (N_8333,N_5437,N_3854);
xor U8334 (N_8334,N_3159,N_3783);
xor U8335 (N_8335,N_5972,N_3892);
nor U8336 (N_8336,N_5928,N_5845);
and U8337 (N_8337,N_4893,N_5817);
xor U8338 (N_8338,N_3676,N_4889);
xor U8339 (N_8339,N_5498,N_3637);
and U8340 (N_8340,N_5859,N_4314);
and U8341 (N_8341,N_3441,N_5446);
nor U8342 (N_8342,N_3393,N_5920);
nor U8343 (N_8343,N_4477,N_3054);
nor U8344 (N_8344,N_5679,N_5973);
xnor U8345 (N_8345,N_3447,N_3437);
nor U8346 (N_8346,N_4578,N_3732);
xnor U8347 (N_8347,N_4464,N_5537);
nand U8348 (N_8348,N_5180,N_5832);
nor U8349 (N_8349,N_4229,N_3332);
or U8350 (N_8350,N_4090,N_3978);
nand U8351 (N_8351,N_3946,N_3970);
nor U8352 (N_8352,N_3649,N_3919);
or U8353 (N_8353,N_5316,N_4849);
and U8354 (N_8354,N_5108,N_4825);
xnor U8355 (N_8355,N_4443,N_5402);
xor U8356 (N_8356,N_4636,N_5012);
or U8357 (N_8357,N_5838,N_3091);
nor U8358 (N_8358,N_5322,N_4927);
xnor U8359 (N_8359,N_4079,N_3195);
nand U8360 (N_8360,N_4484,N_3415);
or U8361 (N_8361,N_4095,N_5126);
xnor U8362 (N_8362,N_5891,N_3813);
nor U8363 (N_8363,N_4648,N_3854);
nand U8364 (N_8364,N_5736,N_5772);
nor U8365 (N_8365,N_5478,N_5202);
xor U8366 (N_8366,N_4206,N_4245);
xnor U8367 (N_8367,N_3489,N_4847);
nand U8368 (N_8368,N_3631,N_4651);
and U8369 (N_8369,N_3977,N_3385);
and U8370 (N_8370,N_3442,N_4405);
nor U8371 (N_8371,N_3408,N_4169);
xnor U8372 (N_8372,N_5606,N_4968);
nand U8373 (N_8373,N_5196,N_3588);
or U8374 (N_8374,N_3492,N_5212);
nand U8375 (N_8375,N_4006,N_4271);
and U8376 (N_8376,N_5288,N_5737);
nand U8377 (N_8377,N_4640,N_5748);
or U8378 (N_8378,N_3940,N_5084);
xnor U8379 (N_8379,N_4518,N_5518);
xor U8380 (N_8380,N_4892,N_4809);
and U8381 (N_8381,N_5897,N_3464);
or U8382 (N_8382,N_4012,N_5614);
or U8383 (N_8383,N_3601,N_4802);
and U8384 (N_8384,N_5505,N_3563);
or U8385 (N_8385,N_4187,N_3708);
xor U8386 (N_8386,N_4264,N_3435);
and U8387 (N_8387,N_3157,N_5865);
xnor U8388 (N_8388,N_4699,N_4405);
nand U8389 (N_8389,N_3663,N_5718);
or U8390 (N_8390,N_5461,N_5436);
and U8391 (N_8391,N_3967,N_3318);
nand U8392 (N_8392,N_4380,N_3247);
or U8393 (N_8393,N_5217,N_4354);
and U8394 (N_8394,N_5965,N_3500);
and U8395 (N_8395,N_3659,N_4147);
and U8396 (N_8396,N_5894,N_3848);
and U8397 (N_8397,N_3866,N_4379);
nor U8398 (N_8398,N_3282,N_3805);
nand U8399 (N_8399,N_3108,N_4204);
or U8400 (N_8400,N_4146,N_3239);
nand U8401 (N_8401,N_4068,N_4007);
nor U8402 (N_8402,N_3340,N_5026);
and U8403 (N_8403,N_4293,N_5346);
nand U8404 (N_8404,N_4304,N_4795);
nand U8405 (N_8405,N_4260,N_3713);
xor U8406 (N_8406,N_3486,N_5357);
or U8407 (N_8407,N_4072,N_3170);
xor U8408 (N_8408,N_3654,N_5319);
xnor U8409 (N_8409,N_3114,N_3863);
or U8410 (N_8410,N_3898,N_5829);
nand U8411 (N_8411,N_3332,N_4176);
or U8412 (N_8412,N_4936,N_5318);
and U8413 (N_8413,N_4090,N_3991);
or U8414 (N_8414,N_4133,N_4686);
or U8415 (N_8415,N_5426,N_5610);
nor U8416 (N_8416,N_3364,N_3858);
nor U8417 (N_8417,N_5247,N_3780);
nor U8418 (N_8418,N_4353,N_5885);
nand U8419 (N_8419,N_3329,N_5365);
or U8420 (N_8420,N_4417,N_3922);
xnor U8421 (N_8421,N_4801,N_5076);
nor U8422 (N_8422,N_3432,N_5737);
nand U8423 (N_8423,N_3195,N_3718);
or U8424 (N_8424,N_5435,N_4146);
nand U8425 (N_8425,N_4878,N_3106);
nand U8426 (N_8426,N_3466,N_4816);
and U8427 (N_8427,N_3672,N_4196);
nor U8428 (N_8428,N_3468,N_4317);
and U8429 (N_8429,N_5161,N_5102);
or U8430 (N_8430,N_4842,N_5362);
and U8431 (N_8431,N_4105,N_3510);
nor U8432 (N_8432,N_5367,N_5077);
nand U8433 (N_8433,N_4582,N_4510);
and U8434 (N_8434,N_4674,N_4329);
or U8435 (N_8435,N_4508,N_3008);
xnor U8436 (N_8436,N_5171,N_5373);
or U8437 (N_8437,N_5410,N_4959);
nor U8438 (N_8438,N_3078,N_4051);
and U8439 (N_8439,N_5916,N_4174);
and U8440 (N_8440,N_3497,N_4361);
or U8441 (N_8441,N_4921,N_5454);
and U8442 (N_8442,N_5991,N_4664);
nor U8443 (N_8443,N_5760,N_5551);
nor U8444 (N_8444,N_3740,N_3668);
xnor U8445 (N_8445,N_4771,N_5798);
xnor U8446 (N_8446,N_5055,N_5833);
nand U8447 (N_8447,N_5385,N_4429);
or U8448 (N_8448,N_3726,N_5081);
and U8449 (N_8449,N_5955,N_5418);
or U8450 (N_8450,N_3835,N_5868);
and U8451 (N_8451,N_4611,N_3375);
or U8452 (N_8452,N_3517,N_5458);
nor U8453 (N_8453,N_4900,N_4895);
nor U8454 (N_8454,N_5170,N_3232);
xor U8455 (N_8455,N_3052,N_4084);
nor U8456 (N_8456,N_4068,N_5949);
and U8457 (N_8457,N_4284,N_4388);
or U8458 (N_8458,N_4295,N_4336);
nand U8459 (N_8459,N_5285,N_5599);
nand U8460 (N_8460,N_4949,N_4427);
xnor U8461 (N_8461,N_4146,N_5222);
nor U8462 (N_8462,N_4340,N_3049);
nand U8463 (N_8463,N_5972,N_3101);
or U8464 (N_8464,N_5660,N_5546);
or U8465 (N_8465,N_4970,N_5695);
nor U8466 (N_8466,N_5655,N_3161);
nor U8467 (N_8467,N_4162,N_3373);
or U8468 (N_8468,N_3968,N_4694);
nand U8469 (N_8469,N_4256,N_5749);
or U8470 (N_8470,N_5615,N_3468);
xnor U8471 (N_8471,N_4444,N_3891);
nor U8472 (N_8472,N_3199,N_4374);
nor U8473 (N_8473,N_4680,N_5286);
and U8474 (N_8474,N_3685,N_5412);
nor U8475 (N_8475,N_3246,N_4792);
or U8476 (N_8476,N_5139,N_3352);
or U8477 (N_8477,N_4936,N_3834);
xor U8478 (N_8478,N_4964,N_4321);
nand U8479 (N_8479,N_4862,N_4562);
and U8480 (N_8480,N_3953,N_5308);
nand U8481 (N_8481,N_4794,N_3564);
nor U8482 (N_8482,N_3045,N_3911);
and U8483 (N_8483,N_5575,N_3680);
nor U8484 (N_8484,N_4575,N_4176);
nor U8485 (N_8485,N_5473,N_5839);
nand U8486 (N_8486,N_5599,N_3178);
or U8487 (N_8487,N_4815,N_4722);
and U8488 (N_8488,N_4742,N_4876);
and U8489 (N_8489,N_3087,N_5948);
nor U8490 (N_8490,N_3210,N_4738);
nand U8491 (N_8491,N_3256,N_4174);
nor U8492 (N_8492,N_5946,N_4107);
nand U8493 (N_8493,N_3809,N_4478);
nor U8494 (N_8494,N_3135,N_4681);
and U8495 (N_8495,N_4734,N_3196);
nand U8496 (N_8496,N_3655,N_4664);
or U8497 (N_8497,N_5007,N_5403);
nand U8498 (N_8498,N_4105,N_5308);
and U8499 (N_8499,N_5315,N_5488);
nand U8500 (N_8500,N_5374,N_4504);
nand U8501 (N_8501,N_3525,N_5506);
xor U8502 (N_8502,N_4968,N_5509);
nand U8503 (N_8503,N_3942,N_5216);
or U8504 (N_8504,N_5343,N_3567);
and U8505 (N_8505,N_3997,N_3872);
nor U8506 (N_8506,N_4390,N_5723);
or U8507 (N_8507,N_3660,N_4598);
nand U8508 (N_8508,N_3351,N_5857);
xnor U8509 (N_8509,N_4175,N_5197);
xor U8510 (N_8510,N_3458,N_3515);
nand U8511 (N_8511,N_4808,N_5594);
and U8512 (N_8512,N_3407,N_4294);
and U8513 (N_8513,N_3408,N_3600);
and U8514 (N_8514,N_3081,N_5232);
and U8515 (N_8515,N_3783,N_5036);
and U8516 (N_8516,N_3587,N_5065);
nor U8517 (N_8517,N_3142,N_5957);
xor U8518 (N_8518,N_4458,N_5587);
nand U8519 (N_8519,N_3388,N_5529);
or U8520 (N_8520,N_5150,N_3663);
and U8521 (N_8521,N_3238,N_5483);
or U8522 (N_8522,N_3377,N_4190);
and U8523 (N_8523,N_3312,N_5309);
or U8524 (N_8524,N_5961,N_5247);
and U8525 (N_8525,N_3010,N_3757);
xor U8526 (N_8526,N_3785,N_4423);
nand U8527 (N_8527,N_3038,N_3665);
nor U8528 (N_8528,N_3712,N_3447);
or U8529 (N_8529,N_5782,N_3804);
nand U8530 (N_8530,N_5002,N_3918);
and U8531 (N_8531,N_5178,N_4694);
nor U8532 (N_8532,N_3029,N_5152);
and U8533 (N_8533,N_3705,N_3980);
nor U8534 (N_8534,N_5253,N_3488);
nor U8535 (N_8535,N_4462,N_3023);
and U8536 (N_8536,N_3502,N_4975);
nand U8537 (N_8537,N_3744,N_3600);
xnor U8538 (N_8538,N_4382,N_3107);
or U8539 (N_8539,N_5696,N_4291);
nand U8540 (N_8540,N_5771,N_4817);
nand U8541 (N_8541,N_4544,N_3859);
nand U8542 (N_8542,N_5283,N_3368);
nand U8543 (N_8543,N_5840,N_3988);
nor U8544 (N_8544,N_5293,N_5050);
and U8545 (N_8545,N_4729,N_3226);
xor U8546 (N_8546,N_4560,N_4450);
or U8547 (N_8547,N_4102,N_4923);
or U8548 (N_8548,N_3801,N_5258);
xor U8549 (N_8549,N_4354,N_4498);
or U8550 (N_8550,N_3508,N_5383);
xor U8551 (N_8551,N_4028,N_5153);
or U8552 (N_8552,N_4668,N_4436);
nand U8553 (N_8553,N_3075,N_5662);
xnor U8554 (N_8554,N_3299,N_4220);
or U8555 (N_8555,N_5286,N_3711);
or U8556 (N_8556,N_4987,N_3106);
nor U8557 (N_8557,N_5103,N_5943);
or U8558 (N_8558,N_4770,N_5637);
xor U8559 (N_8559,N_5222,N_4838);
and U8560 (N_8560,N_5962,N_3991);
and U8561 (N_8561,N_5251,N_3542);
xnor U8562 (N_8562,N_3372,N_3797);
xnor U8563 (N_8563,N_4196,N_3568);
and U8564 (N_8564,N_4407,N_3233);
xor U8565 (N_8565,N_4751,N_4564);
and U8566 (N_8566,N_5834,N_5314);
nand U8567 (N_8567,N_4850,N_3427);
nor U8568 (N_8568,N_5556,N_5077);
nor U8569 (N_8569,N_4659,N_4977);
and U8570 (N_8570,N_5749,N_4543);
and U8571 (N_8571,N_5382,N_5141);
and U8572 (N_8572,N_4659,N_5702);
nand U8573 (N_8573,N_3161,N_5050);
nand U8574 (N_8574,N_4464,N_3599);
and U8575 (N_8575,N_4951,N_3338);
nor U8576 (N_8576,N_5891,N_4712);
nor U8577 (N_8577,N_3745,N_3752);
and U8578 (N_8578,N_4699,N_4889);
nor U8579 (N_8579,N_4707,N_5662);
nand U8580 (N_8580,N_5809,N_4374);
and U8581 (N_8581,N_5207,N_5056);
nand U8582 (N_8582,N_5308,N_3315);
xnor U8583 (N_8583,N_5961,N_3016);
xnor U8584 (N_8584,N_3548,N_5786);
xor U8585 (N_8585,N_3637,N_5176);
nand U8586 (N_8586,N_4648,N_5595);
and U8587 (N_8587,N_5691,N_5631);
nor U8588 (N_8588,N_3759,N_5068);
xor U8589 (N_8589,N_5527,N_4165);
nand U8590 (N_8590,N_3435,N_4964);
nand U8591 (N_8591,N_3409,N_3769);
nor U8592 (N_8592,N_3859,N_3142);
and U8593 (N_8593,N_4851,N_3609);
or U8594 (N_8594,N_5034,N_3895);
and U8595 (N_8595,N_5120,N_5115);
xor U8596 (N_8596,N_4018,N_5715);
nor U8597 (N_8597,N_4284,N_4087);
or U8598 (N_8598,N_4436,N_4494);
nor U8599 (N_8599,N_5061,N_5659);
nor U8600 (N_8600,N_4516,N_4177);
nand U8601 (N_8601,N_5649,N_4096);
nand U8602 (N_8602,N_4134,N_4949);
nor U8603 (N_8603,N_3751,N_5862);
nand U8604 (N_8604,N_3189,N_5590);
nand U8605 (N_8605,N_5773,N_3629);
nor U8606 (N_8606,N_5742,N_3343);
or U8607 (N_8607,N_5911,N_3103);
nand U8608 (N_8608,N_4392,N_3182);
and U8609 (N_8609,N_4267,N_5198);
nand U8610 (N_8610,N_5779,N_4830);
nor U8611 (N_8611,N_3968,N_5407);
xor U8612 (N_8612,N_4751,N_4994);
nand U8613 (N_8613,N_3139,N_4976);
xnor U8614 (N_8614,N_3551,N_4792);
nand U8615 (N_8615,N_4350,N_5305);
nand U8616 (N_8616,N_4629,N_5927);
nand U8617 (N_8617,N_5994,N_5858);
or U8618 (N_8618,N_4693,N_3688);
nor U8619 (N_8619,N_5820,N_5406);
or U8620 (N_8620,N_4957,N_3202);
nand U8621 (N_8621,N_4854,N_3854);
xnor U8622 (N_8622,N_3462,N_3286);
nor U8623 (N_8623,N_5981,N_3347);
nand U8624 (N_8624,N_5955,N_3529);
nor U8625 (N_8625,N_3818,N_4704);
nand U8626 (N_8626,N_4083,N_3196);
or U8627 (N_8627,N_5627,N_4582);
xnor U8628 (N_8628,N_3024,N_4494);
xnor U8629 (N_8629,N_5164,N_4800);
and U8630 (N_8630,N_4223,N_4095);
xnor U8631 (N_8631,N_3383,N_4267);
and U8632 (N_8632,N_3221,N_5512);
nand U8633 (N_8633,N_3371,N_4462);
nand U8634 (N_8634,N_5059,N_3455);
nand U8635 (N_8635,N_5128,N_3525);
or U8636 (N_8636,N_4281,N_3296);
xor U8637 (N_8637,N_4038,N_3756);
nor U8638 (N_8638,N_3546,N_4521);
xor U8639 (N_8639,N_4244,N_5533);
nand U8640 (N_8640,N_3053,N_3790);
and U8641 (N_8641,N_3505,N_3910);
or U8642 (N_8642,N_5584,N_5242);
nor U8643 (N_8643,N_4124,N_4389);
nor U8644 (N_8644,N_4497,N_5270);
xnor U8645 (N_8645,N_5222,N_5274);
or U8646 (N_8646,N_3557,N_4798);
nor U8647 (N_8647,N_3269,N_5182);
nand U8648 (N_8648,N_3016,N_3326);
or U8649 (N_8649,N_5147,N_3041);
xor U8650 (N_8650,N_5996,N_4572);
nor U8651 (N_8651,N_4065,N_4089);
xor U8652 (N_8652,N_3964,N_3305);
xnor U8653 (N_8653,N_4767,N_4972);
nand U8654 (N_8654,N_4392,N_4332);
nand U8655 (N_8655,N_4626,N_5474);
nand U8656 (N_8656,N_3668,N_5616);
and U8657 (N_8657,N_3403,N_4128);
and U8658 (N_8658,N_3586,N_5008);
nand U8659 (N_8659,N_5936,N_3526);
xnor U8660 (N_8660,N_4108,N_3605);
xnor U8661 (N_8661,N_3909,N_3694);
and U8662 (N_8662,N_4275,N_4466);
nor U8663 (N_8663,N_4736,N_3719);
and U8664 (N_8664,N_5684,N_4190);
nand U8665 (N_8665,N_5194,N_5121);
xnor U8666 (N_8666,N_5591,N_4482);
xnor U8667 (N_8667,N_3437,N_5546);
or U8668 (N_8668,N_3935,N_5231);
and U8669 (N_8669,N_3223,N_5097);
and U8670 (N_8670,N_5667,N_3723);
xor U8671 (N_8671,N_3074,N_4519);
nor U8672 (N_8672,N_5205,N_5143);
or U8673 (N_8673,N_4900,N_4520);
nor U8674 (N_8674,N_5214,N_3309);
xor U8675 (N_8675,N_3939,N_5741);
nand U8676 (N_8676,N_5566,N_3632);
nand U8677 (N_8677,N_5086,N_5076);
nand U8678 (N_8678,N_3862,N_5691);
or U8679 (N_8679,N_3971,N_5135);
nor U8680 (N_8680,N_3850,N_5719);
and U8681 (N_8681,N_5021,N_3848);
and U8682 (N_8682,N_5549,N_4771);
nand U8683 (N_8683,N_5033,N_3304);
and U8684 (N_8684,N_4769,N_5592);
and U8685 (N_8685,N_4675,N_4586);
nand U8686 (N_8686,N_5705,N_5789);
nand U8687 (N_8687,N_5433,N_4016);
nor U8688 (N_8688,N_3317,N_3096);
or U8689 (N_8689,N_3332,N_5798);
nand U8690 (N_8690,N_5551,N_4474);
nor U8691 (N_8691,N_3389,N_4736);
nor U8692 (N_8692,N_3049,N_4291);
and U8693 (N_8693,N_4913,N_4199);
nand U8694 (N_8694,N_4444,N_4050);
and U8695 (N_8695,N_4666,N_4392);
nand U8696 (N_8696,N_5789,N_5561);
or U8697 (N_8697,N_5186,N_3306);
nand U8698 (N_8698,N_4555,N_3449);
nor U8699 (N_8699,N_3309,N_3168);
xor U8700 (N_8700,N_3444,N_4845);
nand U8701 (N_8701,N_4278,N_3350);
and U8702 (N_8702,N_4846,N_3371);
xor U8703 (N_8703,N_3438,N_3639);
xor U8704 (N_8704,N_4448,N_3452);
and U8705 (N_8705,N_5271,N_3649);
or U8706 (N_8706,N_3365,N_4945);
and U8707 (N_8707,N_3715,N_5001);
nand U8708 (N_8708,N_4118,N_3427);
nor U8709 (N_8709,N_4048,N_4842);
xor U8710 (N_8710,N_4841,N_3665);
and U8711 (N_8711,N_4296,N_5695);
nand U8712 (N_8712,N_5854,N_3726);
xor U8713 (N_8713,N_3407,N_5483);
nand U8714 (N_8714,N_3052,N_3782);
and U8715 (N_8715,N_4977,N_3648);
nor U8716 (N_8716,N_3445,N_3700);
xnor U8717 (N_8717,N_4820,N_5544);
nand U8718 (N_8718,N_5007,N_3938);
nand U8719 (N_8719,N_5385,N_5519);
xor U8720 (N_8720,N_5040,N_5886);
nand U8721 (N_8721,N_5537,N_4983);
or U8722 (N_8722,N_3888,N_3983);
or U8723 (N_8723,N_3833,N_3201);
or U8724 (N_8724,N_3298,N_3115);
nor U8725 (N_8725,N_4252,N_4435);
xor U8726 (N_8726,N_5680,N_5399);
or U8727 (N_8727,N_3138,N_4285);
and U8728 (N_8728,N_3969,N_5930);
or U8729 (N_8729,N_5486,N_4688);
xor U8730 (N_8730,N_5812,N_4249);
and U8731 (N_8731,N_3264,N_3909);
nor U8732 (N_8732,N_5924,N_5627);
xnor U8733 (N_8733,N_5595,N_3748);
xor U8734 (N_8734,N_4468,N_5351);
xor U8735 (N_8735,N_3362,N_3008);
nand U8736 (N_8736,N_4185,N_3607);
and U8737 (N_8737,N_3028,N_3972);
nor U8738 (N_8738,N_4980,N_4644);
nand U8739 (N_8739,N_5644,N_5481);
or U8740 (N_8740,N_4403,N_5222);
nor U8741 (N_8741,N_4084,N_3839);
nor U8742 (N_8742,N_4130,N_5427);
nor U8743 (N_8743,N_3327,N_4154);
nand U8744 (N_8744,N_4964,N_4382);
xor U8745 (N_8745,N_3472,N_5594);
nor U8746 (N_8746,N_3613,N_4166);
or U8747 (N_8747,N_5276,N_5778);
xor U8748 (N_8748,N_5473,N_3436);
nand U8749 (N_8749,N_5759,N_4026);
nor U8750 (N_8750,N_4123,N_5249);
nor U8751 (N_8751,N_3073,N_3846);
or U8752 (N_8752,N_5403,N_3942);
and U8753 (N_8753,N_5316,N_5112);
or U8754 (N_8754,N_3576,N_4976);
nor U8755 (N_8755,N_4286,N_3826);
and U8756 (N_8756,N_3779,N_3603);
xnor U8757 (N_8757,N_4289,N_5975);
and U8758 (N_8758,N_5453,N_3430);
and U8759 (N_8759,N_3339,N_4957);
nand U8760 (N_8760,N_3570,N_3959);
nand U8761 (N_8761,N_5746,N_5138);
and U8762 (N_8762,N_3670,N_4185);
or U8763 (N_8763,N_5889,N_4195);
nor U8764 (N_8764,N_4401,N_3224);
nand U8765 (N_8765,N_5407,N_3598);
or U8766 (N_8766,N_4069,N_5619);
and U8767 (N_8767,N_3025,N_3882);
or U8768 (N_8768,N_3075,N_5774);
xnor U8769 (N_8769,N_3623,N_4692);
and U8770 (N_8770,N_4999,N_4329);
or U8771 (N_8771,N_5354,N_5186);
nand U8772 (N_8772,N_4271,N_5175);
and U8773 (N_8773,N_3275,N_5324);
or U8774 (N_8774,N_5460,N_3224);
nand U8775 (N_8775,N_3489,N_3541);
nand U8776 (N_8776,N_5516,N_3123);
nor U8777 (N_8777,N_3231,N_5241);
xnor U8778 (N_8778,N_4009,N_3553);
or U8779 (N_8779,N_4894,N_3371);
xnor U8780 (N_8780,N_3412,N_5582);
nand U8781 (N_8781,N_5867,N_5664);
nand U8782 (N_8782,N_3076,N_5124);
nor U8783 (N_8783,N_3962,N_4619);
nand U8784 (N_8784,N_4653,N_4394);
and U8785 (N_8785,N_4387,N_5539);
and U8786 (N_8786,N_3223,N_5252);
or U8787 (N_8787,N_3271,N_5599);
nor U8788 (N_8788,N_5142,N_5170);
xnor U8789 (N_8789,N_4656,N_4392);
nor U8790 (N_8790,N_5658,N_4087);
nand U8791 (N_8791,N_5794,N_5289);
xnor U8792 (N_8792,N_3362,N_5795);
or U8793 (N_8793,N_4250,N_5483);
and U8794 (N_8794,N_4147,N_3847);
and U8795 (N_8795,N_3429,N_3175);
or U8796 (N_8796,N_4446,N_4650);
nand U8797 (N_8797,N_5178,N_5680);
or U8798 (N_8798,N_3667,N_5893);
or U8799 (N_8799,N_4810,N_5928);
and U8800 (N_8800,N_5667,N_4590);
xor U8801 (N_8801,N_3000,N_4669);
nor U8802 (N_8802,N_4160,N_5450);
and U8803 (N_8803,N_3964,N_4013);
nor U8804 (N_8804,N_4290,N_5550);
and U8805 (N_8805,N_3151,N_4171);
and U8806 (N_8806,N_5147,N_3563);
or U8807 (N_8807,N_5333,N_5831);
and U8808 (N_8808,N_4871,N_3342);
and U8809 (N_8809,N_4004,N_5452);
nor U8810 (N_8810,N_4291,N_3974);
nand U8811 (N_8811,N_4324,N_3244);
xnor U8812 (N_8812,N_3604,N_3488);
nor U8813 (N_8813,N_5249,N_4939);
nand U8814 (N_8814,N_3933,N_5249);
or U8815 (N_8815,N_4090,N_4902);
and U8816 (N_8816,N_3104,N_4930);
nand U8817 (N_8817,N_5191,N_5838);
xnor U8818 (N_8818,N_3480,N_5704);
xor U8819 (N_8819,N_5624,N_4940);
or U8820 (N_8820,N_4441,N_5686);
nor U8821 (N_8821,N_5326,N_5389);
xnor U8822 (N_8822,N_3980,N_5230);
or U8823 (N_8823,N_4786,N_3104);
xnor U8824 (N_8824,N_4281,N_5403);
or U8825 (N_8825,N_3479,N_4432);
xnor U8826 (N_8826,N_5917,N_3573);
xor U8827 (N_8827,N_4736,N_4172);
xnor U8828 (N_8828,N_5740,N_4351);
nor U8829 (N_8829,N_3490,N_3721);
xor U8830 (N_8830,N_5614,N_4837);
nand U8831 (N_8831,N_3326,N_4470);
and U8832 (N_8832,N_3809,N_3126);
nand U8833 (N_8833,N_5945,N_3921);
nor U8834 (N_8834,N_4927,N_3815);
and U8835 (N_8835,N_5097,N_4215);
and U8836 (N_8836,N_5701,N_4937);
nand U8837 (N_8837,N_3501,N_3338);
xor U8838 (N_8838,N_3421,N_5975);
and U8839 (N_8839,N_4098,N_4324);
nand U8840 (N_8840,N_4973,N_5849);
or U8841 (N_8841,N_4127,N_4655);
nor U8842 (N_8842,N_5586,N_3077);
or U8843 (N_8843,N_5558,N_5595);
xor U8844 (N_8844,N_3481,N_4847);
xnor U8845 (N_8845,N_4989,N_3489);
nor U8846 (N_8846,N_4860,N_4352);
and U8847 (N_8847,N_5168,N_3107);
nor U8848 (N_8848,N_4651,N_5899);
nor U8849 (N_8849,N_5991,N_3472);
or U8850 (N_8850,N_3206,N_3405);
or U8851 (N_8851,N_3076,N_3523);
nand U8852 (N_8852,N_4672,N_3305);
nor U8853 (N_8853,N_4424,N_5262);
and U8854 (N_8854,N_3916,N_4630);
or U8855 (N_8855,N_3306,N_4600);
and U8856 (N_8856,N_5321,N_5086);
nor U8857 (N_8857,N_3685,N_3618);
or U8858 (N_8858,N_5680,N_5298);
xor U8859 (N_8859,N_4199,N_3752);
nor U8860 (N_8860,N_4889,N_4228);
nor U8861 (N_8861,N_3847,N_4175);
xor U8862 (N_8862,N_5001,N_4957);
nand U8863 (N_8863,N_4383,N_4284);
nor U8864 (N_8864,N_5627,N_5219);
or U8865 (N_8865,N_4631,N_3061);
xor U8866 (N_8866,N_5368,N_3167);
xnor U8867 (N_8867,N_5264,N_3297);
and U8868 (N_8868,N_5935,N_3486);
and U8869 (N_8869,N_3070,N_5742);
xor U8870 (N_8870,N_5210,N_3932);
xnor U8871 (N_8871,N_4417,N_4225);
nor U8872 (N_8872,N_4105,N_5217);
nand U8873 (N_8873,N_5993,N_3431);
and U8874 (N_8874,N_5144,N_5836);
or U8875 (N_8875,N_4422,N_5139);
nand U8876 (N_8876,N_5750,N_5622);
xnor U8877 (N_8877,N_5009,N_4839);
or U8878 (N_8878,N_4163,N_4277);
xor U8879 (N_8879,N_5295,N_4129);
nand U8880 (N_8880,N_3057,N_5721);
nand U8881 (N_8881,N_5012,N_3008);
nor U8882 (N_8882,N_5952,N_4045);
xor U8883 (N_8883,N_3989,N_5355);
or U8884 (N_8884,N_5748,N_4495);
xnor U8885 (N_8885,N_4678,N_3414);
or U8886 (N_8886,N_4001,N_3416);
or U8887 (N_8887,N_5523,N_3751);
xor U8888 (N_8888,N_5292,N_4466);
nand U8889 (N_8889,N_4169,N_3807);
and U8890 (N_8890,N_3499,N_3418);
or U8891 (N_8891,N_5613,N_3308);
or U8892 (N_8892,N_5229,N_5026);
xor U8893 (N_8893,N_3336,N_4722);
xor U8894 (N_8894,N_5961,N_4138);
nor U8895 (N_8895,N_4279,N_4470);
xor U8896 (N_8896,N_4762,N_3754);
and U8897 (N_8897,N_4581,N_3738);
or U8898 (N_8898,N_5739,N_3554);
nor U8899 (N_8899,N_5885,N_4881);
or U8900 (N_8900,N_4928,N_5620);
or U8901 (N_8901,N_4161,N_5872);
nor U8902 (N_8902,N_5309,N_5229);
xnor U8903 (N_8903,N_5156,N_3287);
nor U8904 (N_8904,N_4192,N_5930);
nor U8905 (N_8905,N_5495,N_3365);
nor U8906 (N_8906,N_4714,N_3740);
nand U8907 (N_8907,N_3523,N_4627);
and U8908 (N_8908,N_3897,N_5439);
xnor U8909 (N_8909,N_5165,N_5778);
nand U8910 (N_8910,N_5338,N_5126);
or U8911 (N_8911,N_5653,N_3642);
nor U8912 (N_8912,N_3315,N_3866);
and U8913 (N_8913,N_4381,N_4039);
and U8914 (N_8914,N_3041,N_5889);
and U8915 (N_8915,N_5457,N_4501);
xnor U8916 (N_8916,N_3543,N_4466);
nor U8917 (N_8917,N_3147,N_3421);
xnor U8918 (N_8918,N_5188,N_3046);
or U8919 (N_8919,N_4400,N_3320);
or U8920 (N_8920,N_4806,N_4754);
nand U8921 (N_8921,N_4535,N_5833);
xor U8922 (N_8922,N_5864,N_5299);
xor U8923 (N_8923,N_5663,N_3513);
nor U8924 (N_8924,N_3470,N_5410);
nor U8925 (N_8925,N_4400,N_5400);
and U8926 (N_8926,N_4845,N_3754);
nor U8927 (N_8927,N_4162,N_4699);
and U8928 (N_8928,N_5137,N_5020);
nor U8929 (N_8929,N_3647,N_5996);
nor U8930 (N_8930,N_5491,N_3343);
or U8931 (N_8931,N_3390,N_4155);
or U8932 (N_8932,N_4722,N_3407);
nand U8933 (N_8933,N_3825,N_5356);
nand U8934 (N_8934,N_5263,N_4402);
nor U8935 (N_8935,N_4722,N_5848);
xnor U8936 (N_8936,N_3699,N_4729);
and U8937 (N_8937,N_4927,N_5219);
or U8938 (N_8938,N_4817,N_4450);
or U8939 (N_8939,N_3584,N_4072);
xnor U8940 (N_8940,N_3071,N_5551);
nor U8941 (N_8941,N_3291,N_4182);
or U8942 (N_8942,N_5947,N_4500);
nand U8943 (N_8943,N_5336,N_5954);
or U8944 (N_8944,N_4677,N_4138);
and U8945 (N_8945,N_5547,N_3155);
and U8946 (N_8946,N_4379,N_5318);
xnor U8947 (N_8947,N_4772,N_4263);
nand U8948 (N_8948,N_3326,N_4582);
or U8949 (N_8949,N_4309,N_3548);
and U8950 (N_8950,N_3552,N_5642);
nor U8951 (N_8951,N_3657,N_5564);
nor U8952 (N_8952,N_5973,N_4322);
and U8953 (N_8953,N_3536,N_3886);
or U8954 (N_8954,N_3757,N_3648);
and U8955 (N_8955,N_3020,N_4161);
nor U8956 (N_8956,N_3611,N_5101);
or U8957 (N_8957,N_3576,N_5317);
or U8958 (N_8958,N_5405,N_5458);
or U8959 (N_8959,N_4955,N_4950);
xnor U8960 (N_8960,N_4347,N_5470);
nor U8961 (N_8961,N_5236,N_5331);
nand U8962 (N_8962,N_5425,N_3283);
xor U8963 (N_8963,N_5605,N_5664);
nor U8964 (N_8964,N_3723,N_3122);
and U8965 (N_8965,N_3231,N_4892);
nand U8966 (N_8966,N_3581,N_5602);
xor U8967 (N_8967,N_3703,N_4814);
or U8968 (N_8968,N_4165,N_4456);
nor U8969 (N_8969,N_4056,N_5159);
xor U8970 (N_8970,N_4663,N_5505);
xnor U8971 (N_8971,N_4843,N_3015);
and U8972 (N_8972,N_5203,N_4380);
nand U8973 (N_8973,N_4773,N_5603);
and U8974 (N_8974,N_4530,N_5532);
xnor U8975 (N_8975,N_4923,N_3111);
nor U8976 (N_8976,N_4369,N_4944);
or U8977 (N_8977,N_4611,N_4914);
and U8978 (N_8978,N_4574,N_4098);
nand U8979 (N_8979,N_3284,N_5354);
nand U8980 (N_8980,N_4151,N_5528);
or U8981 (N_8981,N_3337,N_3547);
nor U8982 (N_8982,N_3161,N_3388);
nand U8983 (N_8983,N_5915,N_3868);
nand U8984 (N_8984,N_4819,N_5196);
xor U8985 (N_8985,N_3598,N_3541);
nand U8986 (N_8986,N_3664,N_5325);
and U8987 (N_8987,N_5304,N_4879);
and U8988 (N_8988,N_5742,N_5363);
and U8989 (N_8989,N_4605,N_4269);
nand U8990 (N_8990,N_4888,N_5067);
or U8991 (N_8991,N_5875,N_4305);
xnor U8992 (N_8992,N_5442,N_4165);
or U8993 (N_8993,N_5592,N_3010);
nor U8994 (N_8994,N_3613,N_4332);
and U8995 (N_8995,N_3882,N_4418);
xor U8996 (N_8996,N_3415,N_3515);
and U8997 (N_8997,N_4703,N_3876);
nor U8998 (N_8998,N_3773,N_5304);
xor U8999 (N_8999,N_3118,N_3876);
and U9000 (N_9000,N_7873,N_6788);
and U9001 (N_9001,N_6171,N_6334);
xnor U9002 (N_9002,N_8352,N_8067);
nand U9003 (N_9003,N_7028,N_6534);
xnor U9004 (N_9004,N_8619,N_6708);
or U9005 (N_9005,N_7853,N_6315);
or U9006 (N_9006,N_7516,N_6143);
xor U9007 (N_9007,N_6576,N_6741);
and U9008 (N_9008,N_6084,N_7317);
and U9009 (N_9009,N_8798,N_8127);
or U9010 (N_9010,N_6349,N_8108);
nor U9011 (N_9011,N_6116,N_6193);
or U9012 (N_9012,N_6773,N_6217);
xor U9013 (N_9013,N_7956,N_7274);
nand U9014 (N_9014,N_6156,N_7348);
xor U9015 (N_9015,N_8451,N_8935);
xnor U9016 (N_9016,N_7554,N_6920);
or U9017 (N_9017,N_8507,N_6965);
nor U9018 (N_9018,N_8808,N_7155);
xnor U9019 (N_9019,N_8233,N_8629);
or U9020 (N_9020,N_7588,N_6563);
nand U9021 (N_9021,N_8363,N_6794);
or U9022 (N_9022,N_7659,N_7964);
or U9023 (N_9023,N_8026,N_7574);
nand U9024 (N_9024,N_6991,N_6699);
nand U9025 (N_9025,N_6780,N_7523);
and U9026 (N_9026,N_6742,N_7197);
and U9027 (N_9027,N_6119,N_8684);
nand U9028 (N_9028,N_7909,N_7826);
or U9029 (N_9029,N_8584,N_7815);
nand U9030 (N_9030,N_8424,N_6416);
xnor U9031 (N_9031,N_8217,N_6070);
nor U9032 (N_9032,N_8779,N_7865);
xor U9033 (N_9033,N_8630,N_6019);
nor U9034 (N_9034,N_7113,N_7386);
xor U9035 (N_9035,N_6287,N_8859);
xor U9036 (N_9036,N_8458,N_8946);
and U9037 (N_9037,N_6168,N_6746);
nor U9038 (N_9038,N_6836,N_8764);
nor U9039 (N_9039,N_7968,N_7535);
and U9040 (N_9040,N_8877,N_7112);
xor U9041 (N_9041,N_7316,N_8029);
nand U9042 (N_9042,N_8522,N_7785);
nand U9043 (N_9043,N_6274,N_8490);
nor U9044 (N_9044,N_6461,N_8440);
and U9045 (N_9045,N_8649,N_6378);
nor U9046 (N_9046,N_6237,N_6801);
nand U9047 (N_9047,N_8933,N_8661);
and U9048 (N_9048,N_7140,N_7441);
nand U9049 (N_9049,N_7335,N_6832);
nand U9050 (N_9050,N_6122,N_6927);
nor U9051 (N_9051,N_7200,N_8854);
nand U9052 (N_9052,N_7726,N_8014);
and U9053 (N_9053,N_6248,N_7125);
or U9054 (N_9054,N_7528,N_6969);
nand U9055 (N_9055,N_6958,N_8614);
nor U9056 (N_9056,N_8456,N_8884);
and U9057 (N_9057,N_7463,N_7116);
or U9058 (N_9058,N_8470,N_8774);
nor U9059 (N_9059,N_6729,N_6399);
nand U9060 (N_9060,N_8423,N_8287);
nor U9061 (N_9061,N_6292,N_8050);
and U9062 (N_9062,N_7373,N_8431);
or U9063 (N_9063,N_8413,N_7294);
xor U9064 (N_9064,N_7939,N_6063);
nand U9065 (N_9065,N_8883,N_7009);
and U9066 (N_9066,N_7560,N_8647);
xor U9067 (N_9067,N_8625,N_7144);
nand U9068 (N_9068,N_6553,N_8826);
xnor U9069 (N_9069,N_7589,N_8070);
and U9070 (N_9070,N_6649,N_6629);
nor U9071 (N_9071,N_7745,N_7042);
nand U9072 (N_9072,N_8719,N_7069);
nand U9073 (N_9073,N_6157,N_7425);
nor U9074 (N_9074,N_8567,N_8138);
and U9075 (N_9075,N_7398,N_7118);
nor U9076 (N_9076,N_6716,N_6703);
nand U9077 (N_9077,N_8392,N_6270);
nor U9078 (N_9078,N_6719,N_8472);
nand U9079 (N_9079,N_6772,N_6721);
and U9080 (N_9080,N_6342,N_8527);
and U9081 (N_9081,N_7552,N_6061);
nor U9082 (N_9082,N_8271,N_8715);
or U9083 (N_9083,N_6144,N_7037);
nor U9084 (N_9084,N_8191,N_6659);
nor U9085 (N_9085,N_7891,N_6694);
and U9086 (N_9086,N_7298,N_7885);
nor U9087 (N_9087,N_7164,N_8852);
and U9088 (N_9088,N_7446,N_7637);
and U9089 (N_9089,N_6360,N_6486);
nor U9090 (N_9090,N_8742,N_8480);
or U9091 (N_9091,N_8811,N_6367);
or U9092 (N_9092,N_7011,N_8623);
nand U9093 (N_9093,N_6722,N_7334);
and U9094 (N_9094,N_7310,N_7708);
nand U9095 (N_9095,N_7558,N_7262);
nand U9096 (N_9096,N_6176,N_6604);
nor U9097 (N_9097,N_7951,N_7026);
xnor U9098 (N_9098,N_7471,N_8190);
and U9099 (N_9099,N_7150,N_8252);
xnor U9100 (N_9100,N_8949,N_6779);
and U9101 (N_9101,N_7555,N_7323);
xor U9102 (N_9102,N_8375,N_8083);
nor U9103 (N_9103,N_7814,N_6410);
xor U9104 (N_9104,N_8747,N_6885);
nor U9105 (N_9105,N_6219,N_8677);
or U9106 (N_9106,N_6357,N_7212);
xor U9107 (N_9107,N_8559,N_8314);
xor U9108 (N_9108,N_8275,N_7598);
nor U9109 (N_9109,N_8421,N_8658);
nor U9110 (N_9110,N_6615,N_6295);
or U9111 (N_9111,N_8604,N_8330);
nand U9112 (N_9112,N_7654,N_7712);
xor U9113 (N_9113,N_6484,N_8187);
and U9114 (N_9114,N_8598,N_8934);
nand U9115 (N_9115,N_8267,N_7821);
xnor U9116 (N_9116,N_7754,N_7606);
nand U9117 (N_9117,N_7299,N_7252);
nand U9118 (N_9118,N_8109,N_8114);
nand U9119 (N_9119,N_7942,N_8161);
or U9120 (N_9120,N_7867,N_7085);
and U9121 (N_9121,N_6766,N_6014);
xor U9122 (N_9122,N_8056,N_7549);
and U9123 (N_9123,N_8006,N_8711);
and U9124 (N_9124,N_8732,N_8398);
nand U9125 (N_9125,N_7641,N_8009);
xor U9126 (N_9126,N_7937,N_6189);
or U9127 (N_9127,N_8230,N_8201);
or U9128 (N_9128,N_7190,N_6242);
nand U9129 (N_9129,N_8538,N_6690);
nand U9130 (N_9130,N_6782,N_7084);
or U9131 (N_9131,N_6427,N_7825);
and U9132 (N_9132,N_7897,N_8754);
xor U9133 (N_9133,N_7621,N_7350);
nand U9134 (N_9134,N_7248,N_6134);
nand U9135 (N_9135,N_6457,N_6730);
and U9136 (N_9136,N_8515,N_7353);
or U9137 (N_9137,N_8246,N_8427);
nand U9138 (N_9138,N_7497,N_8845);
nor U9139 (N_9139,N_6020,N_7344);
and U9140 (N_9140,N_6940,N_7965);
or U9141 (N_9141,N_6582,N_7571);
or U9142 (N_9142,N_6145,N_8627);
xnor U9143 (N_9143,N_6464,N_7918);
nand U9144 (N_9144,N_6053,N_8857);
xor U9145 (N_9145,N_8467,N_6137);
and U9146 (N_9146,N_8107,N_8838);
and U9147 (N_9147,N_8439,N_6133);
nor U9148 (N_9148,N_7638,N_8149);
nor U9149 (N_9149,N_7502,N_7223);
nor U9150 (N_9150,N_8713,N_8956);
nor U9151 (N_9151,N_8842,N_7627);
nor U9152 (N_9152,N_7068,N_8690);
or U9153 (N_9153,N_8052,N_7245);
or U9154 (N_9154,N_8321,N_7632);
nand U9155 (N_9155,N_8040,N_7031);
nand U9156 (N_9156,N_6241,N_8958);
xnor U9157 (N_9157,N_7635,N_7001);
and U9158 (N_9158,N_7476,N_6344);
nand U9159 (N_9159,N_7765,N_6449);
nor U9160 (N_9160,N_6692,N_6000);
xor U9161 (N_9161,N_8815,N_6790);
and U9162 (N_9162,N_8790,N_6065);
or U9163 (N_9163,N_8982,N_6191);
and U9164 (N_9164,N_6727,N_8915);
and U9165 (N_9165,N_7566,N_7004);
xor U9166 (N_9166,N_8037,N_6099);
nand U9167 (N_9167,N_8680,N_6804);
nand U9168 (N_9168,N_8539,N_7579);
and U9169 (N_9169,N_6331,N_8167);
or U9170 (N_9170,N_8137,N_8175);
nor U9171 (N_9171,N_6279,N_7370);
or U9172 (N_9172,N_6016,N_6756);
and U9173 (N_9173,N_8139,N_7626);
or U9174 (N_9174,N_8174,N_7599);
and U9175 (N_9175,N_6810,N_7913);
or U9176 (N_9176,N_6547,N_8612);
xor U9177 (N_9177,N_6711,N_6124);
nand U9178 (N_9178,N_7280,N_7686);
nor U9179 (N_9179,N_7972,N_7008);
nand U9180 (N_9180,N_6786,N_7910);
nand U9181 (N_9181,N_8498,N_6872);
nor U9182 (N_9182,N_7027,N_8353);
xnor U9183 (N_9183,N_7952,N_8843);
nand U9184 (N_9184,N_8894,N_8382);
and U9185 (N_9185,N_8529,N_6904);
nor U9186 (N_9186,N_7395,N_8760);
xor U9187 (N_9187,N_6158,N_6866);
nand U9188 (N_9188,N_6761,N_6839);
xnor U9189 (N_9189,N_7360,N_7926);
nand U9190 (N_9190,N_6894,N_6379);
xnor U9191 (N_9191,N_7157,N_8227);
nand U9192 (N_9192,N_8442,N_8476);
nand U9193 (N_9193,N_7800,N_8533);
and U9194 (N_9194,N_8755,N_8298);
or U9195 (N_9195,N_8870,N_7301);
nor U9196 (N_9196,N_6459,N_8061);
and U9197 (N_9197,N_7408,N_7322);
nand U9198 (N_9198,N_7493,N_7034);
xor U9199 (N_9199,N_8750,N_6566);
nand U9200 (N_9200,N_7227,N_8666);
and U9201 (N_9201,N_8657,N_6935);
nand U9202 (N_9202,N_6470,N_8950);
xor U9203 (N_9203,N_6261,N_8501);
nor U9204 (N_9204,N_6106,N_6059);
nor U9205 (N_9205,N_8181,N_7548);
xor U9206 (N_9206,N_6684,N_7556);
or U9207 (N_9207,N_7234,N_6235);
xnor U9208 (N_9208,N_6887,N_7445);
nor U9209 (N_9209,N_8136,N_7273);
xor U9210 (N_9210,N_7817,N_7840);
xnor U9211 (N_9211,N_8587,N_8436);
and U9212 (N_9212,N_7283,N_8202);
nor U9213 (N_9213,N_7473,N_6285);
or U9214 (N_9214,N_8827,N_7567);
or U9215 (N_9215,N_6071,N_6043);
and U9216 (N_9216,N_7169,N_8477);
or U9217 (N_9217,N_6787,N_6549);
and U9218 (N_9218,N_6903,N_7410);
nor U9219 (N_9219,N_7644,N_6283);
nor U9220 (N_9220,N_6712,N_7994);
xor U9221 (N_9221,N_8162,N_7469);
nand U9222 (N_9222,N_7247,N_7624);
or U9223 (N_9223,N_6207,N_6173);
and U9224 (N_9224,N_8012,N_7576);
and U9225 (N_9225,N_7788,N_6616);
nand U9226 (N_9226,N_7828,N_6622);
or U9227 (N_9227,N_7750,N_7547);
xor U9228 (N_9228,N_8333,N_8340);
nor U9229 (N_9229,N_6401,N_6469);
nand U9230 (N_9230,N_8917,N_8411);
and U9231 (N_9231,N_7767,N_6265);
and U9232 (N_9232,N_6186,N_7766);
xor U9233 (N_9233,N_7985,N_6101);
and U9234 (N_9234,N_6160,N_8441);
nor U9235 (N_9235,N_7747,N_7830);
or U9236 (N_9236,N_6500,N_6982);
nand U9237 (N_9237,N_6946,N_6232);
nand U9238 (N_9238,N_7304,N_7531);
xor U9239 (N_9239,N_8445,N_6233);
xnor U9240 (N_9240,N_6519,N_6371);
xor U9241 (N_9241,N_6928,N_8296);
or U9242 (N_9242,N_7770,N_7415);
or U9243 (N_9243,N_7202,N_6952);
nand U9244 (N_9244,N_8046,N_8575);
nor U9245 (N_9245,N_8351,N_8736);
and U9246 (N_9246,N_8608,N_6368);
xnor U9247 (N_9247,N_7563,N_6933);
and U9248 (N_9248,N_6151,N_7670);
or U9249 (N_9249,N_7209,N_6830);
or U9250 (N_9250,N_8342,N_8005);
nand U9251 (N_9251,N_7318,N_8931);
or U9252 (N_9252,N_6948,N_6296);
and U9253 (N_9253,N_7120,N_7604);
or U9254 (N_9254,N_7270,N_7315);
nor U9255 (N_9255,N_8970,N_7844);
and U9256 (N_9256,N_8251,N_7114);
nand U9257 (N_9257,N_6681,N_6531);
nand U9258 (N_9258,N_7551,N_8452);
nor U9259 (N_9259,N_8409,N_7387);
and U9260 (N_9260,N_8971,N_8473);
nand U9261 (N_9261,N_7489,N_6816);
nand U9262 (N_9262,N_7515,N_6573);
xnor U9263 (N_9263,N_7927,N_8513);
xnor U9264 (N_9264,N_6587,N_8752);
xor U9265 (N_9265,N_8987,N_7426);
nor U9266 (N_9266,N_8102,N_7839);
or U9267 (N_9267,N_6949,N_8022);
nand U9268 (N_9268,N_8344,N_6454);
nand U9269 (N_9269,N_8549,N_6299);
nor U9270 (N_9270,N_7281,N_6055);
or U9271 (N_9271,N_7416,N_6931);
xor U9272 (N_9272,N_8100,N_8601);
and U9273 (N_9273,N_8320,N_6393);
nand U9274 (N_9274,N_6642,N_6825);
and U9275 (N_9275,N_8961,N_7459);
nor U9276 (N_9276,N_6275,N_8617);
xor U9277 (N_9277,N_6975,N_6793);
and U9278 (N_9278,N_6436,N_7883);
nand U9279 (N_9279,N_7109,N_6149);
nand U9280 (N_9280,N_6523,N_7030);
nor U9281 (N_9281,N_7279,N_7191);
nor U9282 (N_9282,N_7886,N_6610);
nor U9283 (N_9283,N_7080,N_8992);
nor U9284 (N_9284,N_7479,N_8702);
or U9285 (N_9285,N_6613,N_8903);
nor U9286 (N_9286,N_8322,N_8002);
or U9287 (N_9287,N_8855,N_8142);
xor U9288 (N_9288,N_6685,N_6228);
and U9289 (N_9289,N_8027,N_7220);
nor U9290 (N_9290,N_6923,N_8239);
or U9291 (N_9291,N_7719,N_6889);
and U9292 (N_9292,N_8393,N_6089);
nand U9293 (N_9293,N_8667,N_8724);
or U9294 (N_9294,N_8652,N_7971);
nor U9295 (N_9295,N_7590,N_7752);
nand U9296 (N_9296,N_7126,N_7553);
xor U9297 (N_9297,N_7354,N_8031);
nor U9298 (N_9298,N_8672,N_8210);
nand U9299 (N_9299,N_6601,N_7619);
and U9300 (N_9300,N_7219,N_7934);
nand U9301 (N_9301,N_6184,N_8745);
and U9302 (N_9302,N_7796,N_8509);
xnor U9303 (N_9303,N_7748,N_6535);
or U9304 (N_9304,N_8603,N_6326);
xnor U9305 (N_9305,N_8080,N_7751);
or U9306 (N_9306,N_7863,N_6899);
or U9307 (N_9307,N_8192,N_8407);
xor U9308 (N_9308,N_6980,N_7153);
nor U9309 (N_9309,N_7849,N_8345);
and U9310 (N_9310,N_6971,N_8801);
nand U9311 (N_9311,N_7950,N_7406);
and U9312 (N_9312,N_8150,N_7457);
and U9313 (N_9313,N_7411,N_7777);
or U9314 (N_9314,N_6740,N_7625);
or U9315 (N_9315,N_7110,N_8846);
xor U9316 (N_9316,N_7837,N_7723);
xnor U9317 (N_9317,N_7940,N_8967);
xor U9318 (N_9318,N_8048,N_8128);
or U9319 (N_9319,N_6323,N_8990);
nand U9320 (N_9320,N_6395,N_8795);
or U9321 (N_9321,N_8555,N_7780);
nand U9322 (N_9322,N_8851,N_6828);
and U9323 (N_9323,N_8318,N_7633);
or U9324 (N_9324,N_8374,N_8803);
xnor U9325 (N_9325,N_6339,N_8552);
nor U9326 (N_9326,N_6201,N_7341);
or U9327 (N_9327,N_6526,N_6476);
nand U9328 (N_9328,N_7607,N_8385);
nand U9329 (N_9329,N_7403,N_6674);
xnor U9330 (N_9330,N_8823,N_7456);
xnor U9331 (N_9331,N_8562,N_6387);
nor U9332 (N_9332,N_8646,N_6770);
nor U9333 (N_9333,N_6890,N_6429);
and U9334 (N_9334,N_6064,N_7899);
and U9335 (N_9335,N_7225,N_7240);
and U9336 (N_9336,N_6892,N_7687);
nand U9337 (N_9337,N_6917,N_6878);
nor U9338 (N_9338,N_8908,N_8400);
and U9339 (N_9339,N_8639,N_8292);
nor U9340 (N_9340,N_8304,N_7119);
or U9341 (N_9341,N_8969,N_7389);
nor U9342 (N_9342,N_7409,N_8648);
nor U9343 (N_9343,N_7911,N_6418);
and U9344 (N_9344,N_8316,N_8700);
nand U9345 (N_9345,N_8809,N_6148);
or U9346 (N_9346,N_6081,N_7546);
nor U9347 (N_9347,N_8051,N_8396);
nor U9348 (N_9348,N_7018,N_6864);
nand U9349 (N_9349,N_6440,N_7134);
or U9350 (N_9350,N_6518,N_6709);
xor U9351 (N_9351,N_6293,N_8898);
nor U9352 (N_9352,N_8454,N_6961);
or U9353 (N_9353,N_6004,N_8124);
or U9354 (N_9354,N_8196,N_8081);
nand U9355 (N_9355,N_8521,N_6281);
xnor U9356 (N_9356,N_8880,N_7661);
nor U9357 (N_9357,N_8028,N_8493);
nand U9358 (N_9358,N_7056,N_7525);
xor U9359 (N_9359,N_6224,N_7276);
and U9360 (N_9360,N_7526,N_7465);
and U9361 (N_9361,N_8060,N_7443);
or U9362 (N_9362,N_6052,N_6791);
or U9363 (N_9363,N_8208,N_6951);
nor U9364 (N_9364,N_6468,N_7608);
nand U9365 (N_9365,N_6365,N_6506);
xor U9366 (N_9366,N_7915,N_6691);
and U9367 (N_9367,N_7356,N_6648);
nand U9368 (N_9368,N_7731,N_8899);
nor U9369 (N_9369,N_6271,N_6715);
nor U9370 (N_9370,N_7432,N_6200);
and U9371 (N_9371,N_8420,N_7562);
nor U9372 (N_9372,N_6252,N_8740);
and U9373 (N_9373,N_6789,N_7629);
or U9374 (N_9374,N_8016,N_6294);
or U9375 (N_9375,N_8159,N_8737);
xnor U9376 (N_9376,N_8044,N_8544);
or U9377 (N_9377,N_7980,N_6146);
or U9378 (N_9378,N_7363,N_8998);
nand U9379 (N_9379,N_6682,N_7154);
or U9380 (N_9380,N_8399,N_7268);
or U9381 (N_9381,N_8259,N_6842);
or U9382 (N_9382,N_7700,N_6546);
nand U9383 (N_9383,N_6944,N_7764);
and U9384 (N_9384,N_7652,N_7115);
and U9385 (N_9385,N_7916,N_6250);
xor U9386 (N_9386,N_8064,N_6574);
nor U9387 (N_9387,N_7312,N_8278);
nand U9388 (N_9388,N_7397,N_8328);
nor U9389 (N_9389,N_8678,N_8453);
nor U9390 (N_9390,N_7474,N_6494);
nor U9391 (N_9391,N_7992,N_8834);
and U9392 (N_9392,N_8829,N_7953);
nand U9393 (N_9393,N_6407,N_7047);
or U9394 (N_9394,N_6213,N_8095);
nor U9395 (N_9395,N_6088,N_7585);
and U9396 (N_9396,N_6455,N_6042);
nor U9397 (N_9397,N_6067,N_6117);
nand U9398 (N_9398,N_8593,N_8929);
and U9399 (N_9399,N_7539,N_6888);
and U9400 (N_9400,N_8788,N_7834);
or U9401 (N_9401,N_7870,N_8078);
xnor U9402 (N_9402,N_8238,N_7789);
nor U9403 (N_9403,N_6495,N_6211);
xnor U9404 (N_9404,N_7505,N_8879);
or U9405 (N_9405,N_8624,N_7597);
or U9406 (N_9406,N_7722,N_7584);
and U9407 (N_9407,N_6175,N_7962);
nor U9408 (N_9408,N_8054,N_8386);
nor U9409 (N_9409,N_6047,N_7529);
and U9410 (N_9410,N_8189,N_7366);
nor U9411 (N_9411,N_7685,N_8727);
or U9412 (N_9412,N_8637,N_7216);
and U9413 (N_9413,N_8730,N_8849);
nand U9414 (N_9414,N_7753,N_6205);
nand U9415 (N_9415,N_7186,N_7668);
and U9416 (N_9416,N_8810,N_7400);
or U9417 (N_9417,N_7448,N_6317);
nor U9418 (N_9418,N_6995,N_7508);
nand U9419 (N_9419,N_8506,N_8185);
nor U9420 (N_9420,N_8751,N_7846);
or U9421 (N_9421,N_7842,N_6330);
nand U9422 (N_9422,N_7798,N_8258);
or U9423 (N_9423,N_7933,N_6707);
xor U9424 (N_9424,N_6777,N_7982);
nor U9425 (N_9425,N_7999,N_8011);
xnor U9426 (N_9426,N_7369,N_8117);
nor U9427 (N_9427,N_6919,N_7775);
nor U9428 (N_9428,N_7773,N_7250);
nand U9429 (N_9429,N_7530,N_8841);
nor U9430 (N_9430,N_8674,N_8777);
xnor U9431 (N_9431,N_7133,N_8176);
and U9432 (N_9432,N_7663,N_7928);
nand U9433 (N_9433,N_7527,N_6098);
nor U9434 (N_9434,N_7228,N_8283);
and U9435 (N_9435,N_6868,N_7464);
and U9436 (N_9436,N_7561,N_8395);
or U9437 (N_9437,N_7824,N_7462);
xor U9438 (N_9438,N_6640,N_8426);
nand U9439 (N_9439,N_8379,N_8797);
xor U9440 (N_9440,N_7930,N_7377);
and U9441 (N_9441,N_8045,N_8609);
nor U9442 (N_9442,N_6569,N_6443);
nor U9443 (N_9443,N_7963,N_7781);
or U9444 (N_9444,N_8525,N_6819);
nor U9445 (N_9445,N_8682,N_6388);
nor U9446 (N_9446,N_6280,N_7207);
nand U9447 (N_9447,N_6492,N_7509);
xnor U9448 (N_9448,N_7615,N_7198);
and U9449 (N_9449,N_7935,N_6874);
or U9450 (N_9450,N_8844,N_6181);
or U9451 (N_9451,N_6661,N_7438);
or U9452 (N_9452,N_8309,N_8524);
xnor U9453 (N_9453,N_6583,N_7437);
nor U9454 (N_9454,N_6432,N_7613);
or U9455 (N_9455,N_7036,N_8878);
or U9456 (N_9456,N_7282,N_6343);
and U9457 (N_9457,N_8074,N_8010);
nor U9458 (N_9458,N_6482,N_8173);
and U9459 (N_9459,N_8642,N_8756);
xor U9460 (N_9460,N_6415,N_7647);
nor U9461 (N_9461,N_6700,N_7917);
xor U9462 (N_9462,N_7494,N_7170);
and U9463 (N_9463,N_8853,N_7093);
nor U9464 (N_9464,N_8118,N_8186);
or U9465 (N_9465,N_8554,N_7970);
xor U9466 (N_9466,N_6208,N_6543);
or U9467 (N_9467,N_6049,N_7264);
nand U9468 (N_9468,N_8361,N_6291);
xor U9469 (N_9469,N_8957,N_6258);
nand U9470 (N_9470,N_7492,N_8636);
nor U9471 (N_9471,N_7161,N_8373);
xor U9472 (N_9472,N_6747,N_8530);
nor U9473 (N_9473,N_6167,N_6515);
nor U9474 (N_9474,N_7311,N_6739);
nor U9475 (N_9475,N_8282,N_6845);
xor U9476 (N_9476,N_8821,N_8812);
and U9477 (N_9477,N_7759,N_7359);
nand U9478 (N_9478,N_6598,N_7337);
or U9479 (N_9479,N_6086,N_6979);
and U9480 (N_9480,N_8735,N_7165);
nand U9481 (N_9481,N_6654,N_8698);
nand U9482 (N_9482,N_7466,N_6288);
and U9483 (N_9483,N_8266,N_8558);
or U9484 (N_9484,N_8261,N_6579);
nand U9485 (N_9485,N_7480,N_6223);
or U9486 (N_9486,N_8966,N_7684);
and U9487 (N_9487,N_6863,N_6045);
nand U9488 (N_9488,N_6512,N_6007);
nor U9489 (N_9489,N_8705,N_7450);
and U9490 (N_9490,N_6900,N_6302);
nand U9491 (N_9491,N_8025,N_6366);
nand U9492 (N_9492,N_6797,N_6704);
or U9493 (N_9493,N_6238,N_8368);
nand U9494 (N_9494,N_6257,N_8195);
and U9495 (N_9495,N_7797,N_6272);
nor U9496 (N_9496,N_7107,N_6590);
and U9497 (N_9497,N_7536,N_8550);
xor U9498 (N_9498,N_7858,N_6509);
xor U9499 (N_9499,N_6714,N_7871);
nor U9500 (N_9500,N_8704,N_6220);
and U9501 (N_9501,N_7351,N_8388);
nand U9502 (N_9502,N_6155,N_8867);
xor U9503 (N_9503,N_7984,N_6911);
nor U9504 (N_9504,N_7671,N_8055);
nor U9505 (N_9505,N_8122,N_7058);
and U9506 (N_9506,N_6231,N_6140);
or U9507 (N_9507,N_8902,N_8850);
nor U9508 (N_9508,N_7993,N_8583);
and U9509 (N_9509,N_8172,N_6808);
xnor U9510 (N_9510,N_7453,N_8547);
xor U9511 (N_9511,N_6667,N_7201);
nor U9512 (N_9512,N_8260,N_6570);
nand U9513 (N_9513,N_8911,N_6775);
or U9514 (N_9514,N_6544,N_6597);
nor U9515 (N_9515,N_6752,N_8104);
and U9516 (N_9516,N_7384,N_7564);
xnor U9517 (N_9517,N_7049,N_7330);
and U9518 (N_9518,N_6853,N_8569);
xor U9519 (N_9519,N_7728,N_7306);
nor U9520 (N_9520,N_8640,N_6411);
nand U9521 (N_9521,N_6138,N_8669);
nor U9522 (N_9522,N_6905,N_8376);
and U9523 (N_9523,N_7055,N_6218);
nor U9524 (N_9524,N_6227,N_8783);
xor U9525 (N_9525,N_7087,N_8989);
nor U9526 (N_9526,N_8053,N_7592);
nor U9527 (N_9527,N_6269,N_6303);
xnor U9528 (N_9528,N_7149,N_7468);
or U9529 (N_9529,N_6066,N_6734);
nor U9530 (N_9530,N_7986,N_8775);
nor U9531 (N_9531,N_6972,N_6311);
xnor U9532 (N_9532,N_8403,N_7361);
and U9533 (N_9533,N_8089,N_8572);
and U9534 (N_9534,N_6796,N_7451);
xor U9535 (N_9535,N_7959,N_6107);
and U9536 (N_9536,N_6545,N_6487);
nor U9537 (N_9537,N_8372,N_8813);
nand U9538 (N_9538,N_6198,N_8599);
or U9539 (N_9539,N_8032,N_8468);
and U9540 (N_9540,N_6021,N_8944);
nand U9541 (N_9541,N_8947,N_6754);
nor U9542 (N_9542,N_7677,N_6884);
nor U9543 (N_9543,N_8731,N_6424);
nand U9544 (N_9544,N_6164,N_6239);
or U9545 (N_9545,N_8954,N_8876);
and U9546 (N_9546,N_7481,N_6751);
or U9547 (N_9547,N_8325,N_8694);
nor U9548 (N_9548,N_6136,N_8773);
and U9549 (N_9549,N_8119,N_8020);
and U9550 (N_9550,N_8975,N_6859);
nor U9551 (N_9551,N_6035,N_7596);
and U9552 (N_9552,N_8977,N_8247);
xor U9553 (N_9553,N_6676,N_6439);
nor U9554 (N_9554,N_6724,N_6572);
and U9555 (N_9555,N_8964,N_8900);
nand U9556 (N_9556,N_6128,N_7427);
xnor U9557 (N_9557,N_7580,N_6683);
nor U9558 (N_9558,N_6538,N_6108);
nand U9559 (N_9559,N_8519,N_8145);
xnor U9560 (N_9560,N_8090,N_6152);
nor U9561 (N_9561,N_6705,N_8833);
xor U9562 (N_9562,N_8226,N_6460);
xor U9563 (N_9563,N_7086,N_8800);
xor U9564 (N_9564,N_7924,N_8256);
and U9565 (N_9565,N_6319,N_7218);
and U9566 (N_9566,N_7823,N_8651);
and U9567 (N_9567,N_6425,N_7484);
nor U9568 (N_9568,N_8337,N_6361);
and U9569 (N_9569,N_6332,N_8069);
and U9570 (N_9570,N_6162,N_8329);
or U9571 (N_9571,N_7098,N_6996);
nor U9572 (N_9572,N_8099,N_8786);
nor U9573 (N_9573,N_8995,N_7691);
nand U9574 (N_9574,N_7936,N_6750);
nor U9575 (N_9575,N_7648,N_8086);
xor U9576 (N_9576,N_6174,N_7099);
or U9577 (N_9577,N_7287,N_6688);
xor U9578 (N_9578,N_7171,N_7614);
and U9579 (N_9579,N_6854,N_7045);
nand U9580 (N_9580,N_6824,N_8140);
and U9581 (N_9581,N_8092,N_6118);
and U9582 (N_9582,N_8551,N_7845);
and U9583 (N_9583,N_8543,N_6527);
xor U9584 (N_9584,N_7771,N_7707);
nor U9585 (N_9585,N_7183,N_7594);
nor U9586 (N_9586,N_8459,N_6873);
nor U9587 (N_9587,N_7760,N_6009);
nand U9588 (N_9588,N_6984,N_8508);
xor U9589 (N_9589,N_7716,N_8112);
or U9590 (N_9590,N_7673,N_8941);
nand U9591 (N_9591,N_7996,N_8865);
or U9592 (N_9592,N_6453,N_7478);
or U9593 (N_9593,N_8907,N_8300);
nor U9594 (N_9594,N_6338,N_8837);
and U9595 (N_9595,N_7019,N_7932);
xor U9596 (N_9596,N_7328,N_6994);
nor U9597 (N_9597,N_7860,N_7383);
xor U9598 (N_9598,N_6426,N_6438);
and U9599 (N_9599,N_6530,N_7550);
or U9600 (N_9600,N_7711,N_7269);
nor U9601 (N_9601,N_8804,N_8716);
xnor U9602 (N_9602,N_7023,N_8717);
or U9603 (N_9603,N_6800,N_7532);
or U9604 (N_9604,N_6203,N_8744);
xnor U9605 (N_9605,N_8725,N_7593);
nand U9606 (N_9606,N_6195,N_6170);
nor U9607 (N_9607,N_8221,N_7990);
or U9608 (N_9608,N_8041,N_7213);
and U9609 (N_9609,N_6307,N_8769);
nor U9610 (N_9610,N_7239,N_6290);
and U9611 (N_9611,N_7241,N_8600);
or U9612 (N_9612,N_6732,N_8955);
xor U9613 (N_9613,N_8213,N_7472);
or U9614 (N_9614,N_8302,N_8607);
or U9615 (N_9615,N_6623,N_6953);
nor U9616 (N_9616,N_6305,N_8422);
or U9617 (N_9617,N_7070,N_8708);
nand U9618 (N_9618,N_6584,N_7364);
nor U9619 (N_9619,N_8590,N_7238);
nand U9620 (N_9620,N_6306,N_6717);
nand U9621 (N_9621,N_7025,N_8447);
nor U9622 (N_9622,N_6341,N_7108);
xnor U9623 (N_9623,N_7417,N_7966);
or U9624 (N_9624,N_8244,N_6973);
nor U9625 (N_9625,N_7504,N_6054);
nand U9626 (N_9626,N_6069,N_8289);
and U9627 (N_9627,N_7224,N_8574);
nor U9628 (N_9628,N_8362,N_8789);
xor U9629 (N_9629,N_8297,N_8378);
and U9630 (N_9630,N_6672,N_7645);
nor U9631 (N_9631,N_7715,N_7960);
xnor U9632 (N_9632,N_7215,N_6026);
nand U9633 (N_9633,N_7424,N_6891);
and U9634 (N_9634,N_7880,N_8729);
or U9635 (N_9635,N_6383,N_7185);
and U9636 (N_9636,N_6580,N_7501);
nand U9637 (N_9637,N_7568,N_6079);
nor U9638 (N_9638,N_6422,N_8203);
xor U9639 (N_9639,N_8759,N_7979);
nor U9640 (N_9640,N_8770,N_7703);
and U9641 (N_9641,N_6127,N_8502);
xnor U9642 (N_9642,N_6404,N_6802);
nand U9643 (N_9643,N_7265,N_7309);
and U9644 (N_9644,N_6636,N_8595);
xnor U9645 (N_9645,N_6599,N_7639);
and U9646 (N_9646,N_6112,N_6974);
or U9647 (N_9647,N_7272,N_6651);
or U9648 (N_9648,N_8746,N_7431);
or U9649 (N_9649,N_7156,N_7208);
and U9650 (N_9650,N_8763,N_8463);
nor U9651 (N_9651,N_6028,N_7783);
nand U9652 (N_9652,N_8495,N_6843);
xor U9653 (N_9653,N_8796,N_8354);
or U9654 (N_9654,N_8241,N_7794);
xor U9655 (N_9655,N_8784,N_6044);
nand U9656 (N_9656,N_7292,N_8404);
or U9657 (N_9657,N_8448,N_7898);
and U9658 (N_9658,N_6466,N_6406);
nand U9659 (N_9659,N_7130,N_7314);
and U9660 (N_9660,N_8726,N_7895);
xor U9661 (N_9661,N_6630,N_6606);
nor U9662 (N_9662,N_7083,N_8659);
or U9663 (N_9663,N_8695,N_7617);
nand U9664 (N_9664,N_8339,N_7958);
nand U9665 (N_9665,N_6354,N_8401);
and U9666 (N_9666,N_6192,N_7660);
and U9667 (N_9667,N_6657,N_6934);
or U9668 (N_9668,N_7433,N_6352);
or U9669 (N_9669,N_8628,N_8387);
xnor U9670 (N_9670,N_8184,N_7404);
or U9671 (N_9671,N_8814,N_8341);
or U9672 (N_9672,N_8816,N_8910);
nand U9673 (N_9673,N_8475,N_8868);
or U9674 (N_9674,N_7904,N_6370);
nor U9675 (N_9675,N_7906,N_6989);
xor U9676 (N_9676,N_6893,N_6627);
and U9677 (N_9677,N_8437,N_6032);
xor U9678 (N_9678,N_7062,N_8381);
nor U9679 (N_9679,N_8116,N_6006);
or U9680 (N_9680,N_6329,N_7166);
nand U9681 (N_9681,N_7394,N_8734);
xor U9682 (N_9682,N_6304,N_7135);
and U9683 (N_9683,N_6665,N_6612);
nor U9684 (N_9684,N_6632,N_7831);
nor U9685 (N_9685,N_6165,N_8194);
and U9686 (N_9686,N_8959,N_6322);
and U9687 (N_9687,N_8151,N_6998);
xor U9688 (N_9688,N_7925,N_8541);
xor U9689 (N_9689,N_6608,N_7046);
nor U9690 (N_9690,N_6221,N_8205);
or U9691 (N_9691,N_8577,N_7565);
nor U9692 (N_9692,N_7878,N_6902);
nand U9693 (N_9693,N_6932,N_7941);
and U9694 (N_9694,N_7051,N_6490);
or U9695 (N_9695,N_7843,N_7572);
nor U9696 (N_9696,N_7889,N_7040);
or U9697 (N_9697,N_6723,N_7656);
or U9698 (N_9698,N_7736,N_8709);
nand U9699 (N_9699,N_7355,N_8220);
nand U9700 (N_9700,N_6614,N_6609);
nor U9701 (N_9701,N_6444,N_8450);
nand U9702 (N_9702,N_8824,N_8156);
xor U9703 (N_9703,N_7173,N_6178);
nor U9704 (N_9704,N_8644,N_6462);
and U9705 (N_9705,N_6641,N_8520);
and U9706 (N_9706,N_8429,N_8311);
nand U9707 (N_9707,N_6625,N_7284);
xnor U9708 (N_9708,N_7005,N_6728);
and U9709 (N_9709,N_7653,N_8198);
nand U9710 (N_9710,N_7496,N_6477);
and U9711 (N_9711,N_7434,N_8738);
or U9712 (N_9712,N_7022,N_6883);
and U9713 (N_9713,N_8308,N_7100);
or U9714 (N_9714,N_7778,N_6666);
and U9715 (N_9715,N_8214,N_7340);
nor U9716 (N_9716,N_7053,N_6249);
nand U9717 (N_9717,N_7435,N_7813);
nor U9718 (N_9718,N_6125,N_8200);
and U9719 (N_9719,N_8301,N_6060);
nor U9720 (N_9720,N_8281,N_8347);
xnor U9721 (N_9721,N_6244,N_6744);
nor U9722 (N_9722,N_6456,N_8979);
nand U9723 (N_9723,N_7181,N_6402);
nand U9724 (N_9724,N_7675,N_8358);
and U9725 (N_9725,N_8864,N_8697);
nand U9726 (N_9726,N_7717,N_8034);
xnor U9727 (N_9727,N_7943,N_6446);
nand U9728 (N_9728,N_7961,N_8088);
xnor U9729 (N_9729,N_7570,N_7600);
xnor U9730 (N_9730,N_8653,N_7542);
and U9731 (N_9731,N_6142,N_8356);
nor U9732 (N_9732,N_7701,N_8464);
nor U9733 (N_9733,N_7577,N_6671);
or U9734 (N_9734,N_6840,N_7802);
and U9735 (N_9735,N_6448,N_7147);
nor U9736 (N_9736,N_8043,N_7444);
and U9737 (N_9737,N_7714,N_6646);
xor U9738 (N_9738,N_8579,N_7650);
xor U9739 (N_9739,N_6548,N_6421);
and U9740 (N_9740,N_8780,N_8634);
nor U9741 (N_9741,N_6745,N_7506);
xor U9742 (N_9742,N_7740,N_8597);
xor U9743 (N_9743,N_8023,N_8980);
nand U9744 (N_9744,N_7096,N_8207);
nand U9745 (N_9745,N_6826,N_7987);
and U9746 (N_9746,N_7000,N_6471);
nand U9747 (N_9747,N_6314,N_7162);
nand U9748 (N_9748,N_8696,N_8272);
or U9749 (N_9749,N_8071,N_8062);
or U9750 (N_9750,N_8474,N_7015);
and U9751 (N_9751,N_7612,N_6023);
and U9752 (N_9752,N_6236,N_8066);
nor U9753 (N_9753,N_6736,N_7981);
or U9754 (N_9754,N_8807,N_7111);
nor U9755 (N_9755,N_6803,N_7610);
nor U9756 (N_9756,N_7705,N_8240);
nor U9757 (N_9757,N_6398,N_8517);
nand U9758 (N_9758,N_7672,N_6190);
nand U9759 (N_9759,N_7179,N_7091);
and U9760 (N_9760,N_7290,N_6695);
and U9761 (N_9761,N_6619,N_8015);
nand U9762 (N_9762,N_7032,N_8154);
nand U9763 (N_9763,N_7407,N_6909);
xnor U9764 (N_9764,N_8255,N_6532);
or U9765 (N_9765,N_8416,N_6080);
nand U9766 (N_9766,N_8141,N_7832);
nand U9767 (N_9767,N_8225,N_7300);
or U9768 (N_9768,N_8417,N_6833);
xnor U9769 (N_9769,N_7922,N_6340);
or U9770 (N_9770,N_6503,N_8285);
or U9771 (N_9771,N_8588,N_8568);
nand U9772 (N_9772,N_6087,N_6478);
xor U9773 (N_9773,N_6129,N_6215);
or U9774 (N_9774,N_8496,N_8155);
or U9775 (N_9775,N_6806,N_8038);
and U9776 (N_9776,N_8075,N_7737);
and U9777 (N_9777,N_7017,N_6090);
and U9778 (N_9778,N_7324,N_8564);
nand U9779 (N_9779,N_7513,N_8094);
nor U9780 (N_9780,N_6769,N_8869);
nor U9781 (N_9781,N_6852,N_6748);
xnor U9782 (N_9782,N_8206,N_6511);
nand U9783 (N_9783,N_6130,N_7713);
or U9784 (N_9784,N_6713,N_6963);
xor U9785 (N_9785,N_7698,N_6660);
nand U9786 (N_9786,N_8994,N_8613);
nand U9787 (N_9787,N_8631,N_7420);
xor U9788 (N_9788,N_7847,N_6262);
xor U9789 (N_9789,N_7422,N_8818);
nand U9790 (N_9790,N_8197,N_6259);
nor U9791 (N_9791,N_8976,N_6757);
xor U9792 (N_9792,N_6015,N_7706);
xnor U9793 (N_9793,N_6103,N_6177);
nand U9794 (N_9794,N_6856,N_8242);
nand U9795 (N_9795,N_8557,N_8035);
nor U9796 (N_9796,N_7196,N_7893);
or U9797 (N_9797,N_6277,N_7066);
or U9798 (N_9798,N_7657,N_6551);
nor U9799 (N_9799,N_7852,N_8665);
and U9800 (N_9800,N_7946,N_8924);
or U9801 (N_9801,N_6555,N_8178);
xor U9802 (N_9802,N_6417,N_6652);
nand U9803 (N_9803,N_8866,N_8776);
nand U9804 (N_9804,N_7603,N_8212);
nor U9805 (N_9805,N_7947,N_8291);
xnor U9806 (N_9806,N_7776,N_7735);
nand U9807 (N_9807,N_8951,N_8348);
nor U9808 (N_9808,N_7044,N_8681);
or U9809 (N_9809,N_6072,N_8457);
nand U9810 (N_9810,N_8262,N_8632);
and U9811 (N_9811,N_6960,N_7217);
xnor U9812 (N_9812,N_8610,N_7718);
nand U9813 (N_9813,N_7452,N_6765);
or U9814 (N_9814,N_8805,N_8936);
xor U9815 (N_9815,N_8021,N_6624);
nand U9816 (N_9816,N_8953,N_7266);
xnor U9817 (N_9817,N_6082,N_6335);
and U9818 (N_9818,N_7195,N_6226);
nand U9819 (N_9819,N_6778,N_6644);
and U9820 (N_9820,N_6618,N_8991);
xor U9821 (N_9821,N_7578,N_7249);
nand U9822 (N_9822,N_8707,N_7095);
nand U9823 (N_9823,N_8317,N_8701);
nand U9824 (N_9824,N_7697,N_7907);
and U9825 (N_9825,N_7174,N_8825);
xnor U9826 (N_9826,N_6498,N_7167);
nand U9827 (N_9827,N_7063,N_8836);
nor U9828 (N_9828,N_6479,N_7286);
or U9829 (N_9829,N_6821,N_6327);
xnor U9830 (N_9830,N_8721,N_8765);
or U9831 (N_9831,N_6898,N_7455);
and U9832 (N_9832,N_7854,N_7033);
and U9833 (N_9833,N_6792,N_7475);
and U9834 (N_9834,N_6321,N_6316);
nor U9835 (N_9835,N_8013,N_8875);
or U9836 (N_9836,N_7559,N_8269);
nor U9837 (N_9837,N_7375,N_6048);
nor U9838 (N_9838,N_7729,N_7896);
or U9839 (N_9839,N_7586,N_7319);
xnor U9840 (N_9840,N_6886,N_6559);
nand U9841 (N_9841,N_8714,N_8042);
or U9842 (N_9842,N_6012,N_6650);
nor U9843 (N_9843,N_6434,N_7362);
nand U9844 (N_9844,N_8573,N_8279);
or U9845 (N_9845,N_8231,N_6245);
nand U9846 (N_9846,N_7418,N_8257);
nand U9847 (N_9847,N_7296,N_6110);
xor U9848 (N_9848,N_8586,N_7977);
xor U9849 (N_9849,N_8219,N_8858);
xor U9850 (N_9850,N_6550,N_7634);
or U9851 (N_9851,N_7724,N_7277);
xor U9852 (N_9852,N_7242,N_7921);
or U9853 (N_9853,N_8602,N_7050);
and U9854 (N_9854,N_7540,N_7757);
and U9855 (N_9855,N_8673,N_8433);
and U9856 (N_9856,N_7175,N_6983);
nand U9857 (N_9857,N_8611,N_6726);
nand U9858 (N_9858,N_6031,N_6631);
nand U9859 (N_9859,N_8945,N_8482);
nand U9860 (N_9860,N_7689,N_6731);
nor U9861 (N_9861,N_8772,N_8671);
and U9862 (N_9862,N_6876,N_7811);
and U9863 (N_9863,N_6993,N_7061);
xnor U9864 (N_9864,N_7957,N_7152);
nor U9865 (N_9865,N_6634,N_6420);
xnor U9866 (N_9866,N_8932,N_8718);
nand U9867 (N_9867,N_6795,N_8000);
or U9868 (N_9868,N_6647,N_7694);
nand U9869 (N_9869,N_7378,N_7543);
nor U9870 (N_9870,N_7667,N_8723);
and U9871 (N_9871,N_6959,N_6701);
nor U9872 (N_9872,N_6011,N_6941);
nor U9873 (N_9873,N_6120,N_6621);
xor U9874 (N_9874,N_7710,N_8848);
or U9875 (N_9875,N_7014,N_6126);
xor U9876 (N_9876,N_7226,N_8461);
and U9877 (N_9877,N_7954,N_6161);
or U9878 (N_9878,N_6337,N_7949);
nand U9879 (N_9879,N_8571,N_6182);
and U9880 (N_9880,N_6286,N_7288);
xor U9881 (N_9881,N_8794,N_8978);
nand U9882 (N_9882,N_7016,N_8893);
and U9883 (N_9883,N_6702,N_8147);
xnor U9884 (N_9884,N_8248,N_7630);
nand U9885 (N_9885,N_6463,N_6018);
nand U9886 (N_9886,N_8455,N_6687);
or U9887 (N_9887,N_8860,N_8489);
or U9888 (N_9888,N_7477,N_8578);
or U9889 (N_9889,N_7923,N_8891);
or U9890 (N_9890,N_7182,N_7861);
or U9891 (N_9891,N_6664,N_8606);
or U9892 (N_9892,N_6034,N_6005);
nor U9893 (N_9893,N_7256,N_8856);
xor U9894 (N_9894,N_6499,N_7285);
or U9895 (N_9895,N_8103,N_8589);
nor U9896 (N_9896,N_7210,N_8968);
and U9897 (N_9897,N_6297,N_6831);
and U9898 (N_9898,N_8591,N_6520);
nand U9899 (N_9899,N_8229,N_6858);
or U9900 (N_9900,N_6753,N_8839);
nor U9901 (N_9901,N_6204,N_6749);
nor U9902 (N_9902,N_8135,N_7793);
xnor U9903 (N_9903,N_7812,N_7744);
nand U9904 (N_9904,N_7163,N_7605);
and U9905 (N_9905,N_7510,N_7989);
nor U9906 (N_9906,N_7743,N_8146);
xor U9907 (N_9907,N_6617,N_7372);
nand U9908 (N_9908,N_7890,N_6062);
or U9909 (N_9909,N_6926,N_6225);
nor U9910 (N_9910,N_6172,N_7727);
xor U9911 (N_9911,N_6981,N_8930);
nand U9912 (N_9912,N_7206,N_6865);
and U9913 (N_9913,N_7428,N_7189);
and U9914 (N_9914,N_6345,N_8158);
nand U9915 (N_9915,N_6915,N_6373);
xnor U9916 (N_9916,N_7007,N_6620);
nand U9917 (N_9917,N_7988,N_8822);
or U9918 (N_9918,N_7901,N_7090);
nor U9919 (N_9919,N_8237,N_8592);
and U9920 (N_9920,N_6214,N_6799);
nand U9921 (N_9921,N_6966,N_8594);
xor U9922 (N_9922,N_8511,N_7774);
nand U9923 (N_9923,N_6419,N_8712);
nor U9924 (N_9924,N_6992,N_6536);
or U9925 (N_9925,N_8418,N_8434);
nor U9926 (N_9926,N_7168,N_7127);
nor U9927 (N_9927,N_8280,N_8922);
nand U9928 (N_9928,N_6771,N_6602);
or U9929 (N_9929,N_7818,N_8357);
or U9930 (N_9930,N_8887,N_7178);
and U9931 (N_9931,N_8871,N_6475);
nor U9932 (N_9932,N_7755,N_7020);
nand U9933 (N_9933,N_6093,N_8546);
or U9934 (N_9934,N_6844,N_8397);
nand U9935 (N_9935,N_7092,N_6811);
xor U9936 (N_9936,N_8276,N_7948);
and U9937 (N_9937,N_8249,N_8897);
xor U9938 (N_9938,N_6408,N_8115);
nand U9939 (N_9939,N_7882,N_8762);
nand U9940 (N_9940,N_8927,N_7117);
nand U9941 (N_9941,N_7486,N_8582);
nor U9942 (N_9942,N_7260,N_7973);
nor U9943 (N_9943,N_7742,N_8545);
nor U9944 (N_9944,N_6001,N_7595);
xor U9945 (N_9945,N_7931,N_8912);
xnor U9946 (N_9946,N_7903,N_8315);
and U9947 (N_9947,N_8097,N_8091);
nor U9948 (N_9948,N_7399,N_6929);
and U9949 (N_9949,N_6179,N_7518);
or U9950 (N_9950,N_6662,N_8443);
xnor U9951 (N_9951,N_6094,N_8872);
nand U9952 (N_9952,N_8366,N_8832);
or U9953 (N_9953,N_6588,N_7978);
nor U9954 (N_9954,N_7763,N_8307);
xor U9955 (N_9955,N_8873,N_8974);
nand U9956 (N_9956,N_6567,N_8962);
xnor U9957 (N_9957,N_6922,N_7035);
or U9958 (N_9958,N_7786,N_6102);
and U9959 (N_9959,N_8365,N_8130);
and U9960 (N_9960,N_6414,N_8585);
nor U9961 (N_9961,N_6027,N_8534);
nor U9962 (N_9962,N_7503,N_8004);
nand U9963 (N_9963,N_8049,N_6141);
xor U9964 (N_9964,N_6552,N_8886);
xnor U9965 (N_9965,N_8466,N_6474);
nor U9966 (N_9966,N_7674,N_6392);
nor U9967 (N_9967,N_8319,N_8494);
and U9968 (N_9968,N_6040,N_8633);
xor U9969 (N_9969,N_8928,N_7075);
or U9970 (N_9970,N_6921,N_8105);
nand U9971 (N_9971,N_7636,N_6491);
or U9972 (N_9972,N_7231,N_8312);
nor U9973 (N_9973,N_6637,N_6153);
or U9974 (N_9974,N_6010,N_7749);
and U9975 (N_9975,N_6374,N_7892);
nor U9976 (N_9976,N_8683,N_6967);
and U9977 (N_9977,N_6121,N_7974);
and U9978 (N_9978,N_8101,N_8679);
or U9979 (N_9979,N_7221,N_8536);
nand U9980 (N_9980,N_8164,N_7214);
nand U9981 (N_9981,N_7320,N_6488);
nand U9982 (N_9982,N_8303,N_6850);
xnor U9983 (N_9983,N_8743,N_7041);
xnor U9984 (N_9984,N_6955,N_7944);
or U9985 (N_9985,N_6300,N_6581);
or U9986 (N_9986,N_6829,N_7094);
nand U9987 (N_9987,N_8504,N_8047);
nor U9988 (N_9988,N_7688,N_6377);
xnor U9989 (N_9989,N_6668,N_7145);
and U9990 (N_9990,N_7365,N_6869);
nand U9991 (N_9991,N_7176,N_7345);
nand U9992 (N_9992,N_8093,N_8621);
and U9993 (N_9993,N_7308,N_6986);
and U9994 (N_9994,N_6350,N_6510);
xnor U9995 (N_9995,N_6939,N_6522);
xor U9996 (N_9996,N_8830,N_8384);
or U9997 (N_9997,N_7390,N_8126);
xor U9998 (N_9998,N_8749,N_8984);
nor U9999 (N_9999,N_7799,N_6918);
and U10000 (N_10000,N_7263,N_6785);
xor U10001 (N_10001,N_6362,N_8224);
nand U10002 (N_10002,N_6413,N_6336);
or U10003 (N_10003,N_6111,N_6568);
or U10004 (N_10004,N_8923,N_7702);
nand U10005 (N_10005,N_7591,N_8668);
nand U10006 (N_10006,N_8781,N_7902);
or U10007 (N_10007,N_8110,N_8254);
xnor U10008 (N_10008,N_6783,N_6809);
nand U10009 (N_10009,N_8626,N_7679);
or U10010 (N_10010,N_6458,N_6386);
xor U10011 (N_10011,N_6254,N_6240);
and U10012 (N_10012,N_8402,N_8685);
or U10013 (N_10013,N_6003,N_7756);
or U10014 (N_10014,N_8656,N_6528);
nor U10015 (N_10015,N_8410,N_8905);
or U10016 (N_10016,N_8334,N_8499);
or U10017 (N_10017,N_8881,N_6405);
nand U10018 (N_10018,N_8654,N_7888);
nand U10019 (N_10019,N_6480,N_6180);
or U10020 (N_10020,N_8369,N_8017);
and U10021 (N_10021,N_6123,N_8565);
and U10022 (N_10022,N_6954,N_6943);
and U10023 (N_10023,N_6058,N_8514);
xor U10024 (N_10024,N_6268,N_6533);
nand U10025 (N_10025,N_6369,N_8675);
nand U10026 (N_10026,N_8670,N_8478);
or U10027 (N_10027,N_6784,N_6057);
or U10028 (N_10028,N_6805,N_6759);
or U10029 (N_10029,N_7313,N_7367);
nand U10030 (N_10030,N_8408,N_8981);
nor U10031 (N_10031,N_8650,N_7524);
xnor U10032 (N_10032,N_7021,N_6502);
nand U10033 (N_10033,N_6942,N_6760);
or U10034 (N_10034,N_8232,N_7054);
or U10035 (N_10035,N_6838,N_6013);
xor U10036 (N_10036,N_7609,N_6656);
or U10037 (N_10037,N_8152,N_8072);
nand U10038 (N_10038,N_7631,N_8556);
nor U10039 (N_10039,N_7379,N_8566);
xor U10040 (N_10040,N_7052,N_8085);
xnor U10041 (N_10041,N_8819,N_6860);
or U10042 (N_10042,N_6855,N_7123);
or U10043 (N_10043,N_7623,N_7761);
xnor U10044 (N_10044,N_6447,N_6348);
and U10045 (N_10045,N_7346,N_6251);
nor U10046 (N_10046,N_8986,N_6394);
or U10047 (N_10047,N_8082,N_7271);
and U10048 (N_10048,N_6867,N_7082);
or U10049 (N_10049,N_8581,N_6132);
and U10050 (N_10050,N_8432,N_8618);
or U10051 (N_10051,N_7381,N_8125);
xnor U10052 (N_10052,N_7488,N_7779);
or U10053 (N_10053,N_8030,N_8563);
or U10054 (N_10054,N_8516,N_7148);
nand U10055 (N_10055,N_8323,N_8532);
nor U10056 (N_10056,N_6516,N_7419);
xnor U10057 (N_10057,N_8007,N_7467);
nor U10058 (N_10058,N_6763,N_6298);
nand U10059 (N_10059,N_8033,N_8890);
xnor U10060 (N_10060,N_7233,N_7368);
nor U10061 (N_10061,N_6812,N_6820);
nor U10062 (N_10062,N_6950,N_8018);
nand U10063 (N_10063,N_7159,N_8960);
nand U10064 (N_10064,N_8952,N_8921);
nor U10065 (N_10065,N_6234,N_7333);
xor U10066 (N_10066,N_7640,N_7856);
nand U10067 (N_10067,N_7232,N_7131);
xor U10068 (N_10068,N_6913,N_6645);
nor U10069 (N_10069,N_8084,N_8895);
nor U10070 (N_10070,N_7074,N_8540);
nor U10071 (N_10071,N_6897,N_6987);
or U10072 (N_10072,N_6104,N_8576);
nand U10073 (N_10073,N_6435,N_6473);
and U10074 (N_10074,N_7038,N_6355);
and U10075 (N_10075,N_7012,N_6194);
and U10076 (N_10076,N_6517,N_6758);
nor U10077 (N_10077,N_6767,N_7391);
nor U10078 (N_10078,N_8861,N_7393);
xor U10079 (N_10079,N_8336,N_8940);
or U10080 (N_10080,N_7841,N_7402);
nand U10081 (N_10081,N_8144,N_8123);
xnor U10082 (N_10082,N_6289,N_8645);
xnor U10083 (N_10083,N_6578,N_8024);
nor U10084 (N_10084,N_7658,N_7810);
and U10085 (N_10085,N_6698,N_8346);
xnor U10086 (N_10086,N_6737,N_8817);
nor U10087 (N_10087,N_8518,N_6163);
nand U10088 (N_10088,N_7141,N_7089);
or U10089 (N_10089,N_7680,N_6467);
and U10090 (N_10090,N_6679,N_6437);
xnor U10091 (N_10091,N_8703,N_7920);
nor U10092 (N_10092,N_8901,N_7205);
nand U10093 (N_10093,N_7097,N_8160);
and U10094 (N_10094,N_8706,N_8462);
nand U10095 (N_10095,N_6908,N_7997);
nand U10096 (N_10096,N_7490,N_7430);
nand U10097 (N_10097,N_8503,N_7622);
nor U10098 (N_10098,N_6029,N_6318);
nor U10099 (N_10099,N_6328,N_6397);
or U10100 (N_10100,N_7699,N_8165);
or U10101 (N_10101,N_6085,N_7079);
nand U10102 (N_10102,N_6968,N_8428);
nand U10103 (N_10103,N_8828,N_8722);
nor U10104 (N_10104,N_6391,N_7295);
nor U10105 (N_10105,N_6956,N_7187);
and U10106 (N_10106,N_6628,N_6041);
nor U10107 (N_10107,N_7326,N_6875);
or U10108 (N_10108,N_8121,N_7105);
nor U10109 (N_10109,N_8638,N_6938);
and U10110 (N_10110,N_8350,N_7121);
nand U10111 (N_10111,N_6670,N_8733);
or U10112 (N_10112,N_6978,N_8497);
and U10113 (N_10113,N_6022,N_8120);
nand U10114 (N_10114,N_6489,N_7253);
nand U10115 (N_10115,N_8500,N_7693);
xor U10116 (N_10116,N_7704,N_8691);
nor U10117 (N_10117,N_7442,N_6039);
or U10118 (N_10118,N_7385,N_7139);
xnor U10119 (N_10119,N_6030,N_6564);
or U10120 (N_10120,N_7628,N_8096);
or U10121 (N_10121,N_7077,N_6680);
xnor U10122 (N_10122,N_7881,N_7307);
xor U10123 (N_10123,N_7557,N_8250);
and U10124 (N_10124,N_8364,N_8264);
or U10125 (N_10125,N_6823,N_8215);
nand U10126 (N_10126,N_8414,N_7602);
nand U10127 (N_10127,N_8290,N_8937);
nor U10128 (N_10128,N_6870,N_7073);
xnor U10129 (N_10129,N_8526,N_8741);
or U10130 (N_10130,N_6781,N_8438);
nor U10131 (N_10131,N_7912,N_6267);
or U10132 (N_10132,N_7692,N_7851);
or U10133 (N_10133,N_6755,N_6255);
or U10134 (N_10134,N_8799,N_7519);
nand U10135 (N_10135,N_6901,N_7872);
nand U10136 (N_10136,N_6078,N_6400);
nand U10137 (N_10137,N_7520,N_7461);
nor U10138 (N_10138,N_7376,N_6849);
or U10139 (N_10139,N_7649,N_8888);
xor U10140 (N_10140,N_6036,N_6964);
nand U10141 (N_10141,N_7739,N_6655);
nand U10142 (N_10142,N_7655,N_6914);
or U10143 (N_10143,N_7734,N_6611);
xnor U10144 (N_10144,N_6539,N_8885);
or U10145 (N_10145,N_8390,N_8343);
and U10146 (N_10146,N_7396,N_7908);
nand U10147 (N_10147,N_6896,N_7827);
nand U10148 (N_10148,N_7809,N_7060);
nand U10149 (N_10149,N_8771,N_7507);
nor U10150 (N_10150,N_8655,N_8542);
and U10151 (N_10151,N_6504,N_7967);
or U10152 (N_10152,N_7331,N_6159);
and U10153 (N_10153,N_8492,N_8389);
nor U10154 (N_10154,N_8380,N_6382);
nand U10155 (N_10155,N_6846,N_6282);
and U10156 (N_10156,N_8909,N_6216);
xnor U10157 (N_10157,N_8277,N_6591);
and U10158 (N_10158,N_6596,N_7423);
nor U10159 (N_10159,N_8767,N_7255);
and U10160 (N_10160,N_6188,N_7720);
nor U10161 (N_10161,N_6076,N_7454);
nor U10162 (N_10162,N_8963,N_7804);
or U10163 (N_10163,N_6529,N_8003);
and U10164 (N_10164,N_6097,N_6485);
or U10165 (N_10165,N_6600,N_7709);
and U10166 (N_10166,N_7421,N_8355);
or U10167 (N_10167,N_7392,N_6356);
and U10168 (N_10168,N_7029,N_7618);
and U10169 (N_10169,N_6150,N_6135);
nand U10170 (N_10170,N_8331,N_6433);
or U10171 (N_10171,N_8265,N_7010);
or U10172 (N_10172,N_8616,N_6187);
nand U10173 (N_10173,N_7064,N_7855);
nand U10174 (N_10174,N_8710,N_7343);
or U10175 (N_10175,N_7142,N_7500);
and U10176 (N_10176,N_8486,N_7875);
xnor U10177 (N_10177,N_7512,N_6051);
or U10178 (N_10178,N_6229,N_6083);
xnor U10179 (N_10179,N_6540,N_7278);
or U10180 (N_10180,N_6310,N_8596);
xnor U10181 (N_10181,N_7732,N_8077);
xor U10182 (N_10182,N_8039,N_6183);
nand U10183 (N_10183,N_6450,N_6364);
nor U10184 (N_10184,N_7347,N_8766);
nand U10185 (N_10185,N_6924,N_7829);
xor U10186 (N_10186,N_7405,N_8997);
nor U10187 (N_10187,N_6513,N_6483);
nand U10188 (N_10188,N_6384,N_7769);
xor U10189 (N_10189,N_6068,N_6358);
nand U10190 (N_10190,N_7998,N_8131);
xnor U10191 (N_10191,N_7900,N_6109);
nand U10192 (N_10192,N_7929,N_7768);
nand U10193 (N_10193,N_8076,N_7388);
and U10194 (N_10194,N_6276,N_8999);
xor U10195 (N_10195,N_8157,N_6442);
nor U10196 (N_10196,N_8211,N_8662);
nand U10197 (N_10197,N_7795,N_7013);
or U10198 (N_10198,N_8510,N_6762);
nand U10199 (N_10199,N_7151,N_8643);
and U10200 (N_10200,N_8802,N_7868);
nor U10201 (N_10201,N_7730,N_8561);
nor U10202 (N_10202,N_6658,N_6910);
nor U10203 (N_10203,N_8793,N_7569);
xor U10204 (N_10204,N_6380,N_6537);
nand U10205 (N_10205,N_7894,N_7517);
nand U10206 (N_10206,N_6673,N_6871);
and U10207 (N_10207,N_7914,N_6024);
and U10208 (N_10208,N_8008,N_8892);
nor U10209 (N_10209,N_7138,N_8243);
and U10210 (N_10210,N_6718,N_7820);
and U10211 (N_10211,N_7695,N_8787);
nor U10212 (N_10212,N_8663,N_7762);
or U10213 (N_10213,N_6363,N_7836);
nor U10214 (N_10214,N_6333,N_7819);
or U10215 (N_10215,N_8973,N_7521);
or U10216 (N_10216,N_7884,N_6359);
or U10217 (N_10217,N_8193,N_7485);
nand U10218 (N_10218,N_7222,N_8491);
and U10219 (N_10219,N_8761,N_6273);
nand U10220 (N_10220,N_8111,N_8087);
or U10221 (N_10221,N_6693,N_7859);
xnor U10222 (N_10222,N_8235,N_7611);
nand U10223 (N_10223,N_7682,N_7976);
xor U10224 (N_10224,N_8531,N_7024);
nand U10225 (N_10225,N_6073,N_6593);
or U10226 (N_10226,N_7275,N_6375);
and U10227 (N_10227,N_8134,N_6264);
xor U10228 (N_10228,N_8863,N_8748);
nand U10229 (N_10229,N_8171,N_6677);
xor U10230 (N_10230,N_6710,N_8622);
nor U10231 (N_10231,N_7076,N_7575);
nor U10232 (N_10232,N_7541,N_6514);
nor U10233 (N_10233,N_8073,N_8169);
and U10234 (N_10234,N_7065,N_7081);
nor U10235 (N_10235,N_7143,N_6206);
or U10236 (N_10236,N_8460,N_6697);
nand U10237 (N_10237,N_6508,N_7866);
and U10238 (N_10238,N_7072,N_7129);
nand U10239 (N_10239,N_7136,N_7482);
and U10240 (N_10240,N_6554,N_6957);
xnor U10241 (N_10241,N_8939,N_7088);
nand U10242 (N_10242,N_7101,N_8615);
or U10243 (N_10243,N_6589,N_7106);
xnor U10244 (N_10244,N_6817,N_6209);
or U10245 (N_10245,N_8360,N_8228);
nand U10246 (N_10246,N_7188,N_7995);
nand U10247 (N_10247,N_7791,N_8785);
and U10248 (N_10248,N_6607,N_6114);
or U10249 (N_10249,N_6675,N_6879);
nand U10250 (N_10250,N_6837,N_7104);
nor U10251 (N_10251,N_7864,N_6347);
and U10252 (N_10252,N_6313,N_8113);
or U10253 (N_10253,N_6696,N_8367);
nor U10254 (N_10254,N_7243,N_7938);
or U10255 (N_10255,N_7772,N_6862);
xor U10256 (N_10256,N_8222,N_7371);
and U10257 (N_10257,N_8234,N_7544);
nand U10258 (N_10258,N_7349,N_7808);
xnor U10259 (N_10259,N_6561,N_7869);
xnor U10260 (N_10260,N_8693,N_6501);
and U10261 (N_10261,N_8306,N_8001);
xnor U10262 (N_10262,N_8688,N_7676);
xnor U10263 (N_10263,N_6263,N_7678);
and U10264 (N_10264,N_7230,N_7582);
nand U10265 (N_10265,N_8129,N_7192);
xnor U10266 (N_10266,N_6050,N_6585);
nor U10267 (N_10267,N_7401,N_7137);
xnor U10268 (N_10268,N_7806,N_6095);
nor U10269 (N_10269,N_7983,N_7662);
or U10270 (N_10270,N_7124,N_8479);
nand U10271 (N_10271,N_7681,N_8692);
xnor U10272 (N_10272,N_8079,N_7822);
nor U10273 (N_10273,N_7251,N_6507);
and U10274 (N_10274,N_7132,N_8183);
nor U10275 (N_10275,N_8163,N_8791);
nand U10276 (N_10276,N_6353,N_6266);
nor U10277 (N_10277,N_6312,N_7581);
or U10278 (N_10278,N_7325,N_7975);
xor U10279 (N_10279,N_6243,N_6977);
or U10280 (N_10280,N_7199,N_7733);
or U10281 (N_10281,N_7601,N_7784);
xor U10282 (N_10282,N_8686,N_7039);
nor U10283 (N_10283,N_8019,N_8177);
nor U10284 (N_10284,N_6505,N_8143);
and U10285 (N_10285,N_7332,N_8377);
nand U10286 (N_10286,N_7043,N_8925);
nand U10287 (N_10287,N_7002,N_7339);
and U10288 (N_10288,N_8179,N_7665);
and U10289 (N_10289,N_6807,N_6403);
xnor U10290 (N_10290,N_7721,N_6092);
xor U10291 (N_10291,N_8188,N_7534);
nor U10292 (N_10292,N_8535,N_6430);
nand U10293 (N_10293,N_6764,N_6916);
nor U10294 (N_10294,N_6376,N_8993);
or U10295 (N_10295,N_6768,N_6653);
or U10296 (N_10296,N_7057,N_7254);
xnor U10297 (N_10297,N_8324,N_7048);
nand U10298 (N_10298,N_8299,N_8236);
nor U10299 (N_10299,N_6947,N_6105);
xnor U10300 (N_10300,N_8996,N_8326);
and U10301 (N_10301,N_8620,N_8204);
nand U10302 (N_10302,N_7833,N_8349);
nand U10303 (N_10303,N_6409,N_8553);
nor U10304 (N_10304,N_8943,N_7338);
or U10305 (N_10305,N_7235,N_7850);
xnor U10306 (N_10306,N_6278,N_7838);
nor U10307 (N_10307,N_6706,N_8699);
and U10308 (N_10308,N_8199,N_6881);
xor U10309 (N_10309,N_8058,N_8168);
and U10310 (N_10310,N_7122,N_8449);
xor U10311 (N_10311,N_7193,N_6848);
xnor U10312 (N_10312,N_8313,N_7816);
and U10313 (N_10313,N_6678,N_7449);
xnor U10314 (N_10314,N_8295,N_7177);
nor U10315 (N_10315,N_6524,N_6912);
and U10316 (N_10316,N_7128,N_8965);
or U10317 (N_10317,N_8512,N_8862);
xor U10318 (N_10318,N_8245,N_7180);
nor U10319 (N_10319,N_7067,N_6185);
xnor U10320 (N_10320,N_6496,N_8488);
and U10321 (N_10321,N_6603,N_6557);
xor U10322 (N_10322,N_7969,N_6841);
or U10323 (N_10323,N_6525,N_7204);
and U10324 (N_10324,N_8170,N_7620);
nor U10325 (N_10325,N_8106,N_7573);
nand U10326 (N_10326,N_7805,N_6976);
or U10327 (N_10327,N_7336,N_8270);
nor U10328 (N_10328,N_6985,N_8753);
nand U10329 (N_10329,N_6025,N_7439);
nand U10330 (N_10330,N_6210,N_6389);
xnor U10331 (N_10331,N_8036,N_6197);
xnor U10332 (N_10332,N_6196,N_7991);
xnor U10333 (N_10333,N_6738,N_7160);
nor U10334 (N_10334,N_6936,N_8209);
and U10335 (N_10335,N_7293,N_7244);
xnor U10336 (N_10336,N_7495,N_6169);
nor U10337 (N_10337,N_7352,N_8263);
nor U10338 (N_10338,N_7412,N_8166);
nor U10339 (N_10339,N_8635,N_8926);
and U10340 (N_10340,N_7514,N_6733);
and U10341 (N_10341,N_7289,N_8938);
or U10342 (N_10342,N_8430,N_7103);
nand U10343 (N_10343,N_6222,N_7358);
nand U10344 (N_10344,N_6390,N_7071);
and U10345 (N_10345,N_7146,N_7246);
xor U10346 (N_10346,N_7382,N_8483);
and U10347 (N_10347,N_7236,N_6017);
and U10348 (N_10348,N_8942,N_6669);
and U10349 (N_10349,N_7414,N_6577);
and U10350 (N_10350,N_7848,N_6937);
and U10351 (N_10351,N_7538,N_8739);
nor U10352 (N_10352,N_7158,N_6075);
nand U10353 (N_10353,N_8889,N_8641);
nor U10354 (N_10354,N_6827,N_7887);
and U10355 (N_10355,N_6877,N_7374);
nor U10356 (N_10356,N_8948,N_6556);
nand U10357 (N_10357,N_6396,N_8676);
nor U10358 (N_10358,N_8057,N_8405);
xor U10359 (N_10359,N_6847,N_7738);
or U10360 (N_10360,N_6626,N_7683);
xnor U10361 (N_10361,N_7790,N_7646);
or U10362 (N_10362,N_6835,N_8605);
xor U10363 (N_10363,N_6558,N_7413);
nand U10364 (N_10364,N_7905,N_8806);
nand U10365 (N_10365,N_8469,N_6735);
and U10366 (N_10366,N_8758,N_8660);
or U10367 (N_10367,N_7690,N_6743);
and U10368 (N_10368,N_6497,N_6774);
xor U10369 (N_10369,N_6451,N_8148);
or U10370 (N_10370,N_8689,N_7807);
nand U10371 (N_10371,N_7725,N_8419);
xnor U10372 (N_10372,N_6851,N_7537);
or U10373 (N_10373,N_8904,N_8153);
nand U10374 (N_10374,N_7758,N_7746);
xnor U10375 (N_10375,N_6212,N_8485);
or U10376 (N_10376,N_7321,N_8882);
nor U10377 (N_10377,N_6100,N_7583);
nor U10378 (N_10378,N_8253,N_6988);
nand U10379 (N_10379,N_7511,N_6131);
and U10380 (N_10380,N_8528,N_7955);
xnor U10381 (N_10381,N_6046,N_8560);
xor U10382 (N_10382,N_6033,N_7078);
nor U10383 (N_10383,N_7229,N_7616);
and U10384 (N_10384,N_6147,N_7642);
nand U10385 (N_10385,N_6091,N_7877);
nor U10386 (N_10386,N_8757,N_8294);
nor U10387 (N_10387,N_7184,N_6056);
nand U10388 (N_10388,N_6635,N_7302);
nor U10389 (N_10389,N_8305,N_8435);
and U10390 (N_10390,N_8274,N_8896);
and U10391 (N_10391,N_8505,N_8835);
or U10392 (N_10392,N_7357,N_6906);
nor U10393 (N_10393,N_8916,N_6605);
nand U10394 (N_10394,N_8273,N_6472);
xor U10395 (N_10395,N_8792,N_6562);
xnor U10396 (N_10396,N_8728,N_6199);
nor U10397 (N_10397,N_6834,N_8370);
nor U10398 (N_10398,N_8286,N_6260);
and U10399 (N_10399,N_8383,N_6541);
and U10400 (N_10400,N_7003,N_6113);
xnor U10401 (N_10401,N_8985,N_7919);
nor U10402 (N_10402,N_7522,N_8284);
nand U10403 (N_10403,N_8920,N_7006);
and U10404 (N_10404,N_8327,N_8847);
nand U10405 (N_10405,N_6595,N_6037);
and U10406 (N_10406,N_6230,N_8983);
or U10407 (N_10407,N_8068,N_8720);
xor U10408 (N_10408,N_8098,N_7329);
xor U10409 (N_10409,N_7945,N_6633);
nand U10410 (N_10410,N_6346,N_6308);
nor U10411 (N_10411,N_7491,N_7194);
nand U10412 (N_10412,N_6154,N_6663);
and U10413 (N_10413,N_7879,N_6818);
or U10414 (N_10414,N_6096,N_6441);
nor U10415 (N_10415,N_6565,N_8918);
nand U10416 (N_10416,N_7261,N_7327);
nand U10417 (N_10417,N_8570,N_8906);
and U10418 (N_10418,N_6412,N_7470);
xor U10419 (N_10419,N_7447,N_7258);
xor U10420 (N_10420,N_8182,N_8782);
xor U10421 (N_10421,N_8218,N_6575);
and U10422 (N_10422,N_6930,N_6720);
or U10423 (N_10423,N_6493,N_8180);
xor U10424 (N_10424,N_7792,N_7782);
nand U10425 (N_10425,N_6431,N_7059);
xnor U10426 (N_10426,N_8288,N_8359);
and U10427 (N_10427,N_6465,N_7696);
xor U10428 (N_10428,N_6907,N_7643);
nand U10429 (N_10429,N_6686,N_7587);
nor U10430 (N_10430,N_8268,N_6643);
nand U10431 (N_10431,N_6372,N_7380);
xnor U10432 (N_10432,N_8874,N_8335);
and U10433 (N_10433,N_6638,N_8465);
or U10434 (N_10434,N_7801,N_7876);
or U10435 (N_10435,N_7533,N_6202);
nor U10436 (N_10436,N_7545,N_6882);
and U10437 (N_10437,N_6594,N_6813);
nand U10438 (N_10438,N_7259,N_8371);
nand U10439 (N_10439,N_8216,N_7669);
nand U10440 (N_10440,N_8913,N_6351);
and U10441 (N_10441,N_7664,N_6895);
xor U10442 (N_10442,N_7741,N_8394);
nand U10443 (N_10443,N_6689,N_7483);
nor U10444 (N_10444,N_6822,N_7303);
nor U10445 (N_10445,N_8425,N_6246);
xor U10446 (N_10446,N_8391,N_7874);
nand U10447 (N_10447,N_8523,N_7803);
nor U10448 (N_10448,N_7857,N_6038);
and U10449 (N_10449,N_6798,N_6639);
and U10450 (N_10450,N_6990,N_6284);
or U10451 (N_10451,N_6428,N_6560);
or U10452 (N_10452,N_8914,N_6325);
nand U10453 (N_10453,N_6481,N_6776);
and U10454 (N_10454,N_8293,N_6592);
or U10455 (N_10455,N_6997,N_8481);
or U10456 (N_10456,N_6115,N_8487);
xnor U10457 (N_10457,N_7487,N_6945);
and U10458 (N_10458,N_7666,N_7342);
nand U10459 (N_10459,N_6857,N_6445);
or U10460 (N_10460,N_6301,N_7498);
nor U10461 (N_10461,N_7267,N_6385);
xnor U10462 (N_10462,N_8664,N_7102);
nand U10463 (N_10463,N_6320,N_6925);
nand U10464 (N_10464,N_6324,N_6970);
and U10465 (N_10465,N_8580,N_8820);
or U10466 (N_10466,N_8132,N_7429);
or U10467 (N_10467,N_6256,N_6166);
nor U10468 (N_10468,N_8471,N_8988);
xnor U10469 (N_10469,N_7237,N_7499);
xor U10470 (N_10470,N_8548,N_6381);
nor U10471 (N_10471,N_8133,N_6725);
and U10472 (N_10472,N_8768,N_8831);
xor U10473 (N_10473,N_8310,N_7291);
and U10474 (N_10474,N_6521,N_6008);
or U10475 (N_10475,N_6309,N_6586);
xor U10476 (N_10476,N_6999,N_8484);
and U10477 (N_10477,N_7257,N_8415);
or U10478 (N_10478,N_8840,N_6571);
or U10479 (N_10479,N_7305,N_6542);
xor U10480 (N_10480,N_8778,N_8537);
nand U10481 (N_10481,N_8687,N_8446);
nor U10482 (N_10482,N_8919,N_8059);
nor U10483 (N_10483,N_6814,N_8332);
nand U10484 (N_10484,N_6253,N_6139);
or U10485 (N_10485,N_7172,N_7211);
nor U10486 (N_10486,N_8223,N_6002);
nand U10487 (N_10487,N_7203,N_7862);
and U10488 (N_10488,N_8444,N_8065);
xnor U10489 (N_10489,N_8063,N_8972);
and U10490 (N_10490,N_6452,N_6247);
nand U10491 (N_10491,N_8406,N_7460);
xnor U10492 (N_10492,N_6962,N_8338);
nor U10493 (N_10493,N_7297,N_6074);
xor U10494 (N_10494,N_7651,N_7458);
or U10495 (N_10495,N_6077,N_7787);
xnor U10496 (N_10496,N_6861,N_8412);
nand U10497 (N_10497,N_6880,N_7436);
or U10498 (N_10498,N_6815,N_7835);
and U10499 (N_10499,N_6423,N_7440);
and U10500 (N_10500,N_8770,N_7137);
xnor U10501 (N_10501,N_6216,N_6411);
or U10502 (N_10502,N_8552,N_7207);
nor U10503 (N_10503,N_6728,N_8074);
nand U10504 (N_10504,N_6771,N_6959);
nand U10505 (N_10505,N_6845,N_8769);
nand U10506 (N_10506,N_8472,N_6284);
and U10507 (N_10507,N_8391,N_8922);
and U10508 (N_10508,N_8204,N_7057);
nor U10509 (N_10509,N_8780,N_7567);
and U10510 (N_10510,N_8530,N_8639);
or U10511 (N_10511,N_7597,N_6618);
and U10512 (N_10512,N_8744,N_6154);
nor U10513 (N_10513,N_6057,N_7024);
nand U10514 (N_10514,N_7823,N_6547);
or U10515 (N_10515,N_7124,N_6532);
xnor U10516 (N_10516,N_6535,N_6602);
nor U10517 (N_10517,N_6633,N_6733);
xor U10518 (N_10518,N_7099,N_7426);
or U10519 (N_10519,N_7992,N_6256);
nor U10520 (N_10520,N_6061,N_8778);
nor U10521 (N_10521,N_6484,N_7135);
nand U10522 (N_10522,N_7783,N_8439);
nand U10523 (N_10523,N_8865,N_8138);
or U10524 (N_10524,N_8709,N_8481);
nand U10525 (N_10525,N_6062,N_6208);
xnor U10526 (N_10526,N_7188,N_7325);
and U10527 (N_10527,N_6654,N_8552);
and U10528 (N_10528,N_6118,N_8851);
or U10529 (N_10529,N_8594,N_7553);
and U10530 (N_10530,N_7263,N_7473);
nor U10531 (N_10531,N_8877,N_6917);
xnor U10532 (N_10532,N_7064,N_7200);
xnor U10533 (N_10533,N_7295,N_8518);
xnor U10534 (N_10534,N_8175,N_7855);
or U10535 (N_10535,N_6260,N_6635);
nand U10536 (N_10536,N_8440,N_8004);
xnor U10537 (N_10537,N_8340,N_6120);
xnor U10538 (N_10538,N_7506,N_8353);
xor U10539 (N_10539,N_6425,N_7115);
nor U10540 (N_10540,N_6611,N_6719);
or U10541 (N_10541,N_6001,N_8308);
nor U10542 (N_10542,N_8682,N_6592);
nand U10543 (N_10543,N_8522,N_6969);
xor U10544 (N_10544,N_6817,N_7149);
nand U10545 (N_10545,N_7172,N_8276);
and U10546 (N_10546,N_7629,N_7127);
xnor U10547 (N_10547,N_8122,N_6683);
and U10548 (N_10548,N_8731,N_6930);
nor U10549 (N_10549,N_6546,N_8777);
and U10550 (N_10550,N_6274,N_7774);
nor U10551 (N_10551,N_6599,N_8195);
nand U10552 (N_10552,N_8821,N_6513);
or U10553 (N_10553,N_7251,N_7473);
or U10554 (N_10554,N_6305,N_7527);
and U10555 (N_10555,N_6995,N_7568);
nor U10556 (N_10556,N_6612,N_7956);
nand U10557 (N_10557,N_8376,N_7534);
or U10558 (N_10558,N_6064,N_6524);
nand U10559 (N_10559,N_7522,N_7802);
and U10560 (N_10560,N_6991,N_6479);
and U10561 (N_10561,N_6118,N_8471);
xnor U10562 (N_10562,N_8273,N_8330);
or U10563 (N_10563,N_7820,N_8502);
or U10564 (N_10564,N_8327,N_7495);
and U10565 (N_10565,N_8659,N_7461);
nand U10566 (N_10566,N_6737,N_8038);
or U10567 (N_10567,N_7343,N_6969);
xor U10568 (N_10568,N_8222,N_8635);
or U10569 (N_10569,N_7901,N_6326);
nand U10570 (N_10570,N_8564,N_7866);
xnor U10571 (N_10571,N_6508,N_6729);
xnor U10572 (N_10572,N_7634,N_8565);
xor U10573 (N_10573,N_7666,N_6902);
xor U10574 (N_10574,N_6458,N_7303);
or U10575 (N_10575,N_7860,N_6040);
nand U10576 (N_10576,N_8355,N_6406);
nor U10577 (N_10577,N_8200,N_6579);
and U10578 (N_10578,N_7082,N_6030);
and U10579 (N_10579,N_8758,N_8072);
nor U10580 (N_10580,N_6905,N_7186);
or U10581 (N_10581,N_7572,N_8828);
or U10582 (N_10582,N_6512,N_8271);
xnor U10583 (N_10583,N_8916,N_6336);
or U10584 (N_10584,N_7146,N_7400);
nand U10585 (N_10585,N_6152,N_6635);
or U10586 (N_10586,N_6726,N_6848);
nand U10587 (N_10587,N_8591,N_7577);
or U10588 (N_10588,N_7725,N_7432);
nand U10589 (N_10589,N_8679,N_8825);
nor U10590 (N_10590,N_6156,N_8999);
nor U10591 (N_10591,N_8036,N_6591);
xnor U10592 (N_10592,N_6225,N_8748);
xor U10593 (N_10593,N_6178,N_7044);
xnor U10594 (N_10594,N_7525,N_7731);
xor U10595 (N_10595,N_7041,N_6215);
or U10596 (N_10596,N_6207,N_8892);
xor U10597 (N_10597,N_7714,N_8186);
or U10598 (N_10598,N_8643,N_7358);
xor U10599 (N_10599,N_7494,N_6038);
nor U10600 (N_10600,N_8741,N_8363);
nand U10601 (N_10601,N_7397,N_6160);
and U10602 (N_10602,N_7291,N_8100);
or U10603 (N_10603,N_6607,N_6882);
nor U10604 (N_10604,N_7448,N_6263);
or U10605 (N_10605,N_8669,N_6220);
and U10606 (N_10606,N_8267,N_8039);
nand U10607 (N_10607,N_6695,N_8165);
or U10608 (N_10608,N_8619,N_8902);
and U10609 (N_10609,N_6576,N_6892);
nor U10610 (N_10610,N_8802,N_8798);
and U10611 (N_10611,N_7111,N_7244);
and U10612 (N_10612,N_7246,N_8213);
nor U10613 (N_10613,N_8671,N_7997);
and U10614 (N_10614,N_6765,N_8800);
nand U10615 (N_10615,N_6553,N_6311);
xor U10616 (N_10616,N_8798,N_6066);
nand U10617 (N_10617,N_8943,N_7016);
nand U10618 (N_10618,N_7843,N_6980);
xnor U10619 (N_10619,N_8952,N_8741);
and U10620 (N_10620,N_7642,N_7087);
nor U10621 (N_10621,N_7055,N_8044);
nor U10622 (N_10622,N_8580,N_6494);
or U10623 (N_10623,N_8814,N_8886);
and U10624 (N_10624,N_7523,N_6828);
xnor U10625 (N_10625,N_8045,N_8150);
or U10626 (N_10626,N_6957,N_6229);
or U10627 (N_10627,N_6724,N_8816);
nand U10628 (N_10628,N_8452,N_7267);
or U10629 (N_10629,N_6923,N_7195);
or U10630 (N_10630,N_6524,N_6675);
nand U10631 (N_10631,N_6966,N_8772);
nand U10632 (N_10632,N_8030,N_6036);
or U10633 (N_10633,N_7210,N_6250);
or U10634 (N_10634,N_8641,N_6287);
nand U10635 (N_10635,N_8433,N_7077);
or U10636 (N_10636,N_6918,N_8682);
and U10637 (N_10637,N_8013,N_7896);
nor U10638 (N_10638,N_8699,N_7692);
and U10639 (N_10639,N_6773,N_8955);
or U10640 (N_10640,N_8160,N_6482);
nand U10641 (N_10641,N_7013,N_7702);
nand U10642 (N_10642,N_6028,N_7807);
xnor U10643 (N_10643,N_8342,N_6680);
nand U10644 (N_10644,N_7283,N_6576);
and U10645 (N_10645,N_6971,N_7763);
xor U10646 (N_10646,N_7043,N_7672);
and U10647 (N_10647,N_6803,N_7421);
or U10648 (N_10648,N_7767,N_7060);
xnor U10649 (N_10649,N_8049,N_6362);
or U10650 (N_10650,N_7288,N_7136);
or U10651 (N_10651,N_6709,N_6269);
nand U10652 (N_10652,N_6548,N_8083);
nand U10653 (N_10653,N_6129,N_6489);
nor U10654 (N_10654,N_8940,N_6198);
nand U10655 (N_10655,N_8789,N_7306);
nand U10656 (N_10656,N_6601,N_6308);
and U10657 (N_10657,N_7578,N_6684);
nor U10658 (N_10658,N_7840,N_7417);
nor U10659 (N_10659,N_6395,N_6887);
and U10660 (N_10660,N_7524,N_8565);
and U10661 (N_10661,N_7937,N_8544);
nor U10662 (N_10662,N_8796,N_7369);
xnor U10663 (N_10663,N_7321,N_8165);
xor U10664 (N_10664,N_7976,N_8848);
or U10665 (N_10665,N_8377,N_6526);
or U10666 (N_10666,N_8635,N_8993);
nor U10667 (N_10667,N_7632,N_8450);
xnor U10668 (N_10668,N_7949,N_7922);
nor U10669 (N_10669,N_8485,N_8843);
nor U10670 (N_10670,N_7323,N_6841);
nand U10671 (N_10671,N_7654,N_8193);
nand U10672 (N_10672,N_6926,N_7494);
or U10673 (N_10673,N_7963,N_7450);
nand U10674 (N_10674,N_8095,N_7432);
nand U10675 (N_10675,N_6852,N_7875);
or U10676 (N_10676,N_6887,N_6081);
nor U10677 (N_10677,N_7252,N_8370);
or U10678 (N_10678,N_8187,N_7003);
xnor U10679 (N_10679,N_7590,N_8413);
or U10680 (N_10680,N_8192,N_6836);
or U10681 (N_10681,N_6993,N_6422);
nor U10682 (N_10682,N_8417,N_6982);
nand U10683 (N_10683,N_6172,N_7289);
or U10684 (N_10684,N_8075,N_7107);
nor U10685 (N_10685,N_6685,N_6058);
nor U10686 (N_10686,N_8722,N_7012);
nand U10687 (N_10687,N_7110,N_6196);
xor U10688 (N_10688,N_6053,N_7172);
and U10689 (N_10689,N_7704,N_7304);
or U10690 (N_10690,N_6938,N_6135);
or U10691 (N_10691,N_6604,N_6670);
nand U10692 (N_10692,N_8355,N_7847);
and U10693 (N_10693,N_6067,N_6016);
or U10694 (N_10694,N_7922,N_6194);
xnor U10695 (N_10695,N_6596,N_7783);
nor U10696 (N_10696,N_7173,N_6269);
nor U10697 (N_10697,N_6564,N_8658);
nor U10698 (N_10698,N_8029,N_7787);
nor U10699 (N_10699,N_8562,N_8949);
xor U10700 (N_10700,N_7458,N_8625);
xnor U10701 (N_10701,N_7274,N_6738);
or U10702 (N_10702,N_7094,N_7084);
xnor U10703 (N_10703,N_7976,N_7480);
xnor U10704 (N_10704,N_6923,N_8036);
and U10705 (N_10705,N_7322,N_7709);
nor U10706 (N_10706,N_7143,N_6976);
or U10707 (N_10707,N_6263,N_6942);
nand U10708 (N_10708,N_7786,N_7881);
xnor U10709 (N_10709,N_8373,N_8239);
xor U10710 (N_10710,N_7328,N_7172);
or U10711 (N_10711,N_7768,N_6482);
and U10712 (N_10712,N_8679,N_7438);
xor U10713 (N_10713,N_6653,N_6072);
nand U10714 (N_10714,N_7785,N_7962);
and U10715 (N_10715,N_8341,N_7548);
xnor U10716 (N_10716,N_7789,N_7687);
or U10717 (N_10717,N_8370,N_8669);
or U10718 (N_10718,N_8760,N_6267);
xor U10719 (N_10719,N_6021,N_6869);
nor U10720 (N_10720,N_7072,N_7760);
nor U10721 (N_10721,N_8010,N_7380);
and U10722 (N_10722,N_7834,N_7673);
and U10723 (N_10723,N_7530,N_8226);
nor U10724 (N_10724,N_6876,N_8676);
nand U10725 (N_10725,N_6662,N_8323);
and U10726 (N_10726,N_6728,N_7750);
nor U10727 (N_10727,N_7765,N_6121);
nand U10728 (N_10728,N_6995,N_6817);
or U10729 (N_10729,N_6112,N_7806);
nand U10730 (N_10730,N_6252,N_7977);
xor U10731 (N_10731,N_6282,N_6818);
and U10732 (N_10732,N_8426,N_7136);
xor U10733 (N_10733,N_8019,N_8944);
xor U10734 (N_10734,N_8586,N_6958);
nand U10735 (N_10735,N_7334,N_6772);
nor U10736 (N_10736,N_7881,N_8311);
nor U10737 (N_10737,N_7061,N_8540);
nor U10738 (N_10738,N_8428,N_7198);
and U10739 (N_10739,N_8750,N_8000);
and U10740 (N_10740,N_8993,N_7552);
xnor U10741 (N_10741,N_8338,N_7393);
or U10742 (N_10742,N_6756,N_7358);
and U10743 (N_10743,N_7842,N_8530);
or U10744 (N_10744,N_6773,N_7205);
nand U10745 (N_10745,N_8639,N_7950);
nor U10746 (N_10746,N_6409,N_8498);
or U10747 (N_10747,N_8223,N_8074);
xor U10748 (N_10748,N_8410,N_6219);
or U10749 (N_10749,N_6776,N_7187);
and U10750 (N_10750,N_6453,N_6879);
or U10751 (N_10751,N_8767,N_7838);
xor U10752 (N_10752,N_6012,N_6202);
xnor U10753 (N_10753,N_8415,N_6969);
nor U10754 (N_10754,N_8635,N_8602);
xor U10755 (N_10755,N_6745,N_7056);
and U10756 (N_10756,N_7410,N_6553);
nor U10757 (N_10757,N_8281,N_7468);
xnor U10758 (N_10758,N_8664,N_7502);
or U10759 (N_10759,N_8089,N_8311);
or U10760 (N_10760,N_6608,N_7980);
or U10761 (N_10761,N_7300,N_7210);
xnor U10762 (N_10762,N_7766,N_8190);
or U10763 (N_10763,N_6730,N_7531);
nand U10764 (N_10764,N_7076,N_7478);
nand U10765 (N_10765,N_6246,N_8515);
nor U10766 (N_10766,N_6905,N_8320);
or U10767 (N_10767,N_8478,N_8016);
xnor U10768 (N_10768,N_7803,N_7643);
nand U10769 (N_10769,N_8853,N_6095);
or U10770 (N_10770,N_7376,N_7782);
nor U10771 (N_10771,N_6522,N_8887);
or U10772 (N_10772,N_7038,N_7001);
xor U10773 (N_10773,N_8696,N_8431);
xnor U10774 (N_10774,N_6092,N_6613);
nand U10775 (N_10775,N_7545,N_7503);
and U10776 (N_10776,N_6368,N_6720);
nor U10777 (N_10777,N_7970,N_8302);
nand U10778 (N_10778,N_8018,N_6291);
or U10779 (N_10779,N_6056,N_7143);
or U10780 (N_10780,N_8231,N_8548);
nand U10781 (N_10781,N_6297,N_7532);
nand U10782 (N_10782,N_7831,N_7687);
and U10783 (N_10783,N_6332,N_6362);
or U10784 (N_10784,N_8168,N_6468);
nand U10785 (N_10785,N_6536,N_8512);
xnor U10786 (N_10786,N_7212,N_8271);
or U10787 (N_10787,N_7283,N_7243);
xor U10788 (N_10788,N_8376,N_6674);
nor U10789 (N_10789,N_8494,N_6381);
xnor U10790 (N_10790,N_7891,N_8037);
or U10791 (N_10791,N_6542,N_6136);
and U10792 (N_10792,N_7344,N_8396);
nand U10793 (N_10793,N_8608,N_8654);
and U10794 (N_10794,N_7316,N_6618);
nand U10795 (N_10795,N_7741,N_8441);
and U10796 (N_10796,N_7915,N_6163);
xnor U10797 (N_10797,N_6647,N_8968);
xor U10798 (N_10798,N_8353,N_6935);
and U10799 (N_10799,N_7077,N_8004);
and U10800 (N_10800,N_7196,N_6112);
xor U10801 (N_10801,N_8240,N_8014);
and U10802 (N_10802,N_6380,N_7087);
nand U10803 (N_10803,N_6370,N_7409);
or U10804 (N_10804,N_7014,N_6524);
xnor U10805 (N_10805,N_8619,N_8863);
nand U10806 (N_10806,N_7286,N_8137);
and U10807 (N_10807,N_8357,N_7901);
or U10808 (N_10808,N_6633,N_6926);
nor U10809 (N_10809,N_8807,N_8426);
nand U10810 (N_10810,N_7628,N_8513);
or U10811 (N_10811,N_7559,N_6449);
and U10812 (N_10812,N_6361,N_7521);
and U10813 (N_10813,N_6017,N_7846);
or U10814 (N_10814,N_8343,N_7060);
xnor U10815 (N_10815,N_8906,N_7140);
nor U10816 (N_10816,N_7437,N_6546);
nand U10817 (N_10817,N_7698,N_8843);
and U10818 (N_10818,N_6741,N_6539);
nand U10819 (N_10819,N_8449,N_8555);
xor U10820 (N_10820,N_7230,N_6376);
nor U10821 (N_10821,N_6177,N_8136);
or U10822 (N_10822,N_7106,N_8053);
and U10823 (N_10823,N_8717,N_6581);
or U10824 (N_10824,N_8013,N_7544);
or U10825 (N_10825,N_6604,N_6656);
or U10826 (N_10826,N_8157,N_6108);
and U10827 (N_10827,N_6383,N_8126);
xor U10828 (N_10828,N_8844,N_7516);
xnor U10829 (N_10829,N_8225,N_7892);
or U10830 (N_10830,N_7568,N_7044);
and U10831 (N_10831,N_7887,N_8537);
nand U10832 (N_10832,N_8341,N_7711);
nor U10833 (N_10833,N_6046,N_6718);
nor U10834 (N_10834,N_7914,N_8095);
nor U10835 (N_10835,N_6259,N_8205);
and U10836 (N_10836,N_8006,N_7702);
or U10837 (N_10837,N_8987,N_8900);
and U10838 (N_10838,N_7986,N_6162);
xor U10839 (N_10839,N_8518,N_8411);
nor U10840 (N_10840,N_7697,N_6770);
or U10841 (N_10841,N_8859,N_7698);
xor U10842 (N_10842,N_7215,N_8579);
and U10843 (N_10843,N_8084,N_7842);
nand U10844 (N_10844,N_6680,N_7818);
xor U10845 (N_10845,N_6516,N_7863);
xnor U10846 (N_10846,N_6828,N_8239);
nand U10847 (N_10847,N_8134,N_7954);
xnor U10848 (N_10848,N_6260,N_7053);
and U10849 (N_10849,N_7709,N_6239);
xnor U10850 (N_10850,N_7108,N_7349);
or U10851 (N_10851,N_8713,N_7861);
or U10852 (N_10852,N_6831,N_6657);
nand U10853 (N_10853,N_8275,N_7058);
or U10854 (N_10854,N_6211,N_8905);
xor U10855 (N_10855,N_6009,N_6977);
nor U10856 (N_10856,N_7338,N_8401);
xnor U10857 (N_10857,N_6008,N_8663);
and U10858 (N_10858,N_6227,N_7989);
or U10859 (N_10859,N_7260,N_7169);
nor U10860 (N_10860,N_6495,N_8567);
nand U10861 (N_10861,N_8722,N_7927);
xor U10862 (N_10862,N_7067,N_6915);
xor U10863 (N_10863,N_6820,N_8205);
or U10864 (N_10864,N_6336,N_8307);
and U10865 (N_10865,N_8687,N_7890);
xor U10866 (N_10866,N_7935,N_7754);
nor U10867 (N_10867,N_8914,N_8494);
nor U10868 (N_10868,N_6572,N_6580);
and U10869 (N_10869,N_6369,N_8355);
xnor U10870 (N_10870,N_7648,N_8511);
and U10871 (N_10871,N_6201,N_8058);
or U10872 (N_10872,N_6324,N_6462);
and U10873 (N_10873,N_7983,N_7975);
nor U10874 (N_10874,N_7611,N_6039);
nand U10875 (N_10875,N_7167,N_6443);
xnor U10876 (N_10876,N_7324,N_7879);
and U10877 (N_10877,N_6266,N_8331);
nor U10878 (N_10878,N_7178,N_7434);
nand U10879 (N_10879,N_8341,N_8674);
or U10880 (N_10880,N_8080,N_7621);
xnor U10881 (N_10881,N_8071,N_7715);
nor U10882 (N_10882,N_6949,N_7183);
and U10883 (N_10883,N_8077,N_7427);
and U10884 (N_10884,N_7272,N_8059);
and U10885 (N_10885,N_6677,N_8000);
xnor U10886 (N_10886,N_8156,N_6261);
or U10887 (N_10887,N_6579,N_6178);
xnor U10888 (N_10888,N_6528,N_7515);
or U10889 (N_10889,N_8369,N_7562);
or U10890 (N_10890,N_7626,N_8932);
nor U10891 (N_10891,N_6110,N_7563);
xor U10892 (N_10892,N_8599,N_6180);
nor U10893 (N_10893,N_7231,N_8024);
and U10894 (N_10894,N_7221,N_8821);
and U10895 (N_10895,N_7114,N_7624);
and U10896 (N_10896,N_8268,N_6542);
and U10897 (N_10897,N_8794,N_6009);
nand U10898 (N_10898,N_7448,N_7079);
or U10899 (N_10899,N_8641,N_8859);
xor U10900 (N_10900,N_7098,N_8707);
nand U10901 (N_10901,N_8974,N_7912);
or U10902 (N_10902,N_6772,N_8643);
nand U10903 (N_10903,N_8820,N_7777);
nor U10904 (N_10904,N_8586,N_6425);
nor U10905 (N_10905,N_8119,N_8115);
nand U10906 (N_10906,N_7212,N_6732);
and U10907 (N_10907,N_6827,N_7077);
xnor U10908 (N_10908,N_6569,N_8235);
nor U10909 (N_10909,N_8747,N_7321);
nand U10910 (N_10910,N_7114,N_7799);
nand U10911 (N_10911,N_8737,N_8426);
xor U10912 (N_10912,N_8552,N_6150);
xnor U10913 (N_10913,N_6432,N_6698);
and U10914 (N_10914,N_7906,N_6280);
and U10915 (N_10915,N_6190,N_6129);
nand U10916 (N_10916,N_7449,N_7466);
nor U10917 (N_10917,N_7854,N_8444);
or U10918 (N_10918,N_6701,N_8141);
xnor U10919 (N_10919,N_8822,N_7856);
and U10920 (N_10920,N_7181,N_6331);
nor U10921 (N_10921,N_6110,N_8202);
nor U10922 (N_10922,N_8336,N_8820);
nand U10923 (N_10923,N_7458,N_8008);
nor U10924 (N_10924,N_8306,N_8712);
nor U10925 (N_10925,N_6119,N_7466);
and U10926 (N_10926,N_8158,N_6704);
or U10927 (N_10927,N_8011,N_7727);
nand U10928 (N_10928,N_6044,N_8335);
nor U10929 (N_10929,N_7401,N_6468);
nor U10930 (N_10930,N_8225,N_7270);
and U10931 (N_10931,N_6238,N_7896);
and U10932 (N_10932,N_6377,N_8595);
nor U10933 (N_10933,N_7647,N_8984);
xnor U10934 (N_10934,N_7537,N_7029);
nor U10935 (N_10935,N_8340,N_6163);
or U10936 (N_10936,N_7034,N_8836);
nor U10937 (N_10937,N_6009,N_8951);
nor U10938 (N_10938,N_8374,N_8529);
nand U10939 (N_10939,N_7006,N_8228);
and U10940 (N_10940,N_7521,N_8199);
nor U10941 (N_10941,N_8791,N_6715);
xor U10942 (N_10942,N_6325,N_8796);
nand U10943 (N_10943,N_6655,N_6841);
xor U10944 (N_10944,N_7798,N_7044);
nand U10945 (N_10945,N_8878,N_6021);
xnor U10946 (N_10946,N_7958,N_8904);
nor U10947 (N_10947,N_7039,N_7638);
nand U10948 (N_10948,N_7188,N_7031);
or U10949 (N_10949,N_6005,N_6841);
or U10950 (N_10950,N_7407,N_8960);
nand U10951 (N_10951,N_8400,N_6046);
or U10952 (N_10952,N_8689,N_8212);
nor U10953 (N_10953,N_6146,N_8852);
or U10954 (N_10954,N_8997,N_8300);
nor U10955 (N_10955,N_8197,N_6510);
or U10956 (N_10956,N_7731,N_6443);
and U10957 (N_10957,N_6336,N_7879);
nand U10958 (N_10958,N_7253,N_6858);
nor U10959 (N_10959,N_8025,N_6732);
and U10960 (N_10960,N_8445,N_8244);
nor U10961 (N_10961,N_6352,N_7663);
xor U10962 (N_10962,N_6728,N_6345);
and U10963 (N_10963,N_7592,N_8488);
xnor U10964 (N_10964,N_6519,N_6266);
nor U10965 (N_10965,N_7551,N_6652);
and U10966 (N_10966,N_7262,N_7309);
xor U10967 (N_10967,N_8990,N_7373);
xnor U10968 (N_10968,N_6955,N_6777);
xor U10969 (N_10969,N_7813,N_8193);
nand U10970 (N_10970,N_7965,N_8269);
xor U10971 (N_10971,N_7833,N_7428);
nor U10972 (N_10972,N_8134,N_6883);
and U10973 (N_10973,N_6472,N_8083);
or U10974 (N_10974,N_6240,N_6516);
and U10975 (N_10975,N_6748,N_7240);
and U10976 (N_10976,N_8260,N_7681);
nand U10977 (N_10977,N_6034,N_7190);
nand U10978 (N_10978,N_6533,N_8007);
or U10979 (N_10979,N_8457,N_8048);
and U10980 (N_10980,N_6160,N_8083);
or U10981 (N_10981,N_8320,N_8361);
xor U10982 (N_10982,N_8642,N_6021);
xnor U10983 (N_10983,N_7208,N_7930);
xnor U10984 (N_10984,N_6412,N_6673);
and U10985 (N_10985,N_7661,N_6273);
nor U10986 (N_10986,N_8382,N_8124);
nand U10987 (N_10987,N_6151,N_7677);
and U10988 (N_10988,N_6620,N_7952);
nor U10989 (N_10989,N_7794,N_6645);
xor U10990 (N_10990,N_8042,N_8819);
and U10991 (N_10991,N_8566,N_8719);
xnor U10992 (N_10992,N_7398,N_7906);
and U10993 (N_10993,N_6679,N_6375);
nor U10994 (N_10994,N_7343,N_8146);
or U10995 (N_10995,N_8318,N_7334);
xor U10996 (N_10996,N_6424,N_6667);
nand U10997 (N_10997,N_7470,N_8682);
nor U10998 (N_10998,N_6394,N_8950);
or U10999 (N_10999,N_8474,N_6433);
nor U11000 (N_11000,N_8772,N_7165);
nand U11001 (N_11001,N_7678,N_8310);
and U11002 (N_11002,N_7694,N_8928);
and U11003 (N_11003,N_6073,N_6981);
or U11004 (N_11004,N_7355,N_6661);
nor U11005 (N_11005,N_6276,N_8983);
and U11006 (N_11006,N_7023,N_8193);
nand U11007 (N_11007,N_8469,N_6716);
nor U11008 (N_11008,N_7896,N_6697);
or U11009 (N_11009,N_6447,N_8236);
nand U11010 (N_11010,N_6922,N_6545);
or U11011 (N_11011,N_7253,N_6668);
xnor U11012 (N_11012,N_8240,N_6004);
nor U11013 (N_11013,N_8040,N_6020);
xnor U11014 (N_11014,N_6215,N_7829);
xor U11015 (N_11015,N_6113,N_8041);
nand U11016 (N_11016,N_7682,N_8877);
nand U11017 (N_11017,N_6723,N_8810);
xor U11018 (N_11018,N_6236,N_6843);
or U11019 (N_11019,N_7899,N_8012);
nand U11020 (N_11020,N_6265,N_6405);
and U11021 (N_11021,N_8938,N_8125);
and U11022 (N_11022,N_6608,N_6204);
xnor U11023 (N_11023,N_8119,N_8076);
or U11024 (N_11024,N_6909,N_8130);
and U11025 (N_11025,N_7601,N_6045);
xor U11026 (N_11026,N_8865,N_8565);
nor U11027 (N_11027,N_7867,N_7999);
nor U11028 (N_11028,N_8505,N_7213);
and U11029 (N_11029,N_8879,N_7537);
nor U11030 (N_11030,N_6153,N_8505);
nand U11031 (N_11031,N_6951,N_7279);
nand U11032 (N_11032,N_7516,N_6906);
and U11033 (N_11033,N_6621,N_6233);
nor U11034 (N_11034,N_6632,N_8847);
and U11035 (N_11035,N_6711,N_7090);
nand U11036 (N_11036,N_6980,N_6725);
and U11037 (N_11037,N_6077,N_6013);
nor U11038 (N_11038,N_8331,N_8229);
and U11039 (N_11039,N_8686,N_7057);
nand U11040 (N_11040,N_6000,N_6457);
nor U11041 (N_11041,N_7382,N_7680);
nand U11042 (N_11042,N_8418,N_6941);
or U11043 (N_11043,N_8109,N_7905);
nor U11044 (N_11044,N_7905,N_7121);
nor U11045 (N_11045,N_6409,N_8339);
xnor U11046 (N_11046,N_7198,N_7317);
and U11047 (N_11047,N_8233,N_8315);
nand U11048 (N_11048,N_7538,N_6979);
nand U11049 (N_11049,N_8799,N_8544);
xnor U11050 (N_11050,N_6521,N_6042);
xor U11051 (N_11051,N_6686,N_8960);
nor U11052 (N_11052,N_8568,N_7954);
and U11053 (N_11053,N_7687,N_6966);
nand U11054 (N_11054,N_7282,N_7621);
nand U11055 (N_11055,N_7476,N_7811);
nor U11056 (N_11056,N_8443,N_6235);
xor U11057 (N_11057,N_7773,N_6299);
nand U11058 (N_11058,N_8220,N_6026);
xor U11059 (N_11059,N_7006,N_8930);
nand U11060 (N_11060,N_7257,N_6144);
nor U11061 (N_11061,N_6442,N_7959);
xnor U11062 (N_11062,N_8926,N_7023);
nand U11063 (N_11063,N_7128,N_7324);
nand U11064 (N_11064,N_8039,N_6934);
nand U11065 (N_11065,N_7521,N_6334);
and U11066 (N_11066,N_8739,N_8586);
and U11067 (N_11067,N_7871,N_7713);
xnor U11068 (N_11068,N_7501,N_6671);
and U11069 (N_11069,N_7347,N_7538);
nor U11070 (N_11070,N_8696,N_7650);
xor U11071 (N_11071,N_8439,N_8634);
nor U11072 (N_11072,N_8203,N_8248);
nand U11073 (N_11073,N_8276,N_6388);
or U11074 (N_11074,N_6119,N_6056);
xnor U11075 (N_11075,N_6409,N_7386);
nor U11076 (N_11076,N_7377,N_6675);
nor U11077 (N_11077,N_6143,N_8374);
or U11078 (N_11078,N_8519,N_7055);
or U11079 (N_11079,N_6333,N_6501);
nor U11080 (N_11080,N_7082,N_6390);
nor U11081 (N_11081,N_7711,N_6106);
and U11082 (N_11082,N_6471,N_8865);
xnor U11083 (N_11083,N_8224,N_8341);
xnor U11084 (N_11084,N_8602,N_6847);
and U11085 (N_11085,N_6097,N_8675);
or U11086 (N_11086,N_8013,N_6930);
and U11087 (N_11087,N_7376,N_7191);
nand U11088 (N_11088,N_6452,N_7088);
nand U11089 (N_11089,N_7170,N_8561);
xnor U11090 (N_11090,N_7454,N_6663);
nand U11091 (N_11091,N_8826,N_6956);
nor U11092 (N_11092,N_8904,N_7614);
nand U11093 (N_11093,N_8429,N_7470);
and U11094 (N_11094,N_7952,N_6910);
xor U11095 (N_11095,N_6843,N_8781);
and U11096 (N_11096,N_7729,N_7529);
nand U11097 (N_11097,N_8197,N_6726);
or U11098 (N_11098,N_6894,N_8977);
or U11099 (N_11099,N_7033,N_7921);
or U11100 (N_11100,N_7147,N_8662);
xnor U11101 (N_11101,N_6990,N_7684);
nor U11102 (N_11102,N_8509,N_6531);
xnor U11103 (N_11103,N_6068,N_8681);
xor U11104 (N_11104,N_8996,N_8489);
nand U11105 (N_11105,N_6545,N_8475);
xnor U11106 (N_11106,N_7447,N_7165);
or U11107 (N_11107,N_7314,N_6849);
xor U11108 (N_11108,N_7923,N_7032);
xor U11109 (N_11109,N_8804,N_7064);
nand U11110 (N_11110,N_6875,N_8962);
xnor U11111 (N_11111,N_8766,N_8507);
and U11112 (N_11112,N_8135,N_8387);
or U11113 (N_11113,N_6761,N_7453);
and U11114 (N_11114,N_7584,N_7417);
nand U11115 (N_11115,N_8254,N_8739);
and U11116 (N_11116,N_7179,N_7949);
nand U11117 (N_11117,N_7898,N_6984);
and U11118 (N_11118,N_8622,N_7627);
or U11119 (N_11119,N_6631,N_8514);
and U11120 (N_11120,N_6148,N_7927);
nand U11121 (N_11121,N_7359,N_8962);
and U11122 (N_11122,N_7623,N_8229);
and U11123 (N_11123,N_6533,N_7919);
xor U11124 (N_11124,N_6165,N_8071);
xor U11125 (N_11125,N_8350,N_7902);
and U11126 (N_11126,N_7522,N_6806);
xor U11127 (N_11127,N_7538,N_6133);
nand U11128 (N_11128,N_6359,N_6125);
nor U11129 (N_11129,N_8529,N_6309);
nand U11130 (N_11130,N_6653,N_6199);
nor U11131 (N_11131,N_7346,N_7303);
nand U11132 (N_11132,N_6478,N_6691);
and U11133 (N_11133,N_7656,N_8962);
or U11134 (N_11134,N_8740,N_8827);
or U11135 (N_11135,N_7369,N_8993);
nor U11136 (N_11136,N_6057,N_7592);
xnor U11137 (N_11137,N_8939,N_7867);
nor U11138 (N_11138,N_6774,N_7939);
nor U11139 (N_11139,N_6705,N_7291);
nor U11140 (N_11140,N_7219,N_7815);
nand U11141 (N_11141,N_6189,N_8190);
and U11142 (N_11142,N_6281,N_7424);
and U11143 (N_11143,N_6881,N_8419);
xor U11144 (N_11144,N_8372,N_6645);
and U11145 (N_11145,N_6649,N_6489);
and U11146 (N_11146,N_6087,N_8464);
xor U11147 (N_11147,N_6374,N_6832);
nand U11148 (N_11148,N_8421,N_7535);
nand U11149 (N_11149,N_6635,N_7976);
xor U11150 (N_11150,N_7000,N_6032);
xnor U11151 (N_11151,N_6382,N_7236);
or U11152 (N_11152,N_7271,N_6879);
or U11153 (N_11153,N_6944,N_6939);
xnor U11154 (N_11154,N_7422,N_8367);
xor U11155 (N_11155,N_6015,N_8393);
and U11156 (N_11156,N_8451,N_8450);
or U11157 (N_11157,N_6250,N_8020);
nor U11158 (N_11158,N_8960,N_7740);
and U11159 (N_11159,N_6110,N_7755);
or U11160 (N_11160,N_6417,N_7615);
nor U11161 (N_11161,N_6295,N_6611);
nor U11162 (N_11162,N_7826,N_6673);
nand U11163 (N_11163,N_6152,N_8012);
and U11164 (N_11164,N_7778,N_7586);
xor U11165 (N_11165,N_8547,N_8427);
xnor U11166 (N_11166,N_8671,N_8403);
or U11167 (N_11167,N_6745,N_6469);
nor U11168 (N_11168,N_7207,N_6528);
nor U11169 (N_11169,N_7512,N_8763);
xor U11170 (N_11170,N_8152,N_7282);
or U11171 (N_11171,N_8641,N_6783);
or U11172 (N_11172,N_8657,N_6602);
nand U11173 (N_11173,N_8027,N_7770);
xor U11174 (N_11174,N_6394,N_8163);
xnor U11175 (N_11175,N_6259,N_7997);
or U11176 (N_11176,N_8561,N_7264);
nor U11177 (N_11177,N_7924,N_6720);
nor U11178 (N_11178,N_6678,N_8448);
xnor U11179 (N_11179,N_6496,N_6118);
nor U11180 (N_11180,N_6195,N_6394);
and U11181 (N_11181,N_6653,N_8538);
nand U11182 (N_11182,N_8943,N_7178);
or U11183 (N_11183,N_7894,N_6108);
xor U11184 (N_11184,N_8239,N_6240);
and U11185 (N_11185,N_7999,N_8488);
nand U11186 (N_11186,N_7272,N_8246);
xor U11187 (N_11187,N_8606,N_7347);
nand U11188 (N_11188,N_8460,N_6201);
and U11189 (N_11189,N_7353,N_7311);
nor U11190 (N_11190,N_7919,N_6284);
xor U11191 (N_11191,N_6198,N_7256);
and U11192 (N_11192,N_6254,N_8977);
or U11193 (N_11193,N_7152,N_8377);
xnor U11194 (N_11194,N_6058,N_8387);
and U11195 (N_11195,N_8906,N_6145);
and U11196 (N_11196,N_6803,N_8128);
or U11197 (N_11197,N_7952,N_8305);
nor U11198 (N_11198,N_8106,N_7426);
nand U11199 (N_11199,N_8700,N_6805);
or U11200 (N_11200,N_7429,N_7860);
and U11201 (N_11201,N_6663,N_8385);
xnor U11202 (N_11202,N_7814,N_8578);
or U11203 (N_11203,N_6617,N_6842);
and U11204 (N_11204,N_6648,N_7345);
nor U11205 (N_11205,N_7302,N_8583);
xnor U11206 (N_11206,N_7365,N_8003);
or U11207 (N_11207,N_6220,N_6966);
nand U11208 (N_11208,N_8230,N_8332);
and U11209 (N_11209,N_7120,N_8569);
or U11210 (N_11210,N_7303,N_7921);
xnor U11211 (N_11211,N_8341,N_8406);
nor U11212 (N_11212,N_7988,N_8340);
nor U11213 (N_11213,N_6640,N_6450);
and U11214 (N_11214,N_8330,N_8500);
nand U11215 (N_11215,N_6680,N_7996);
or U11216 (N_11216,N_8950,N_6000);
xnor U11217 (N_11217,N_8091,N_7803);
nand U11218 (N_11218,N_8275,N_7603);
or U11219 (N_11219,N_7848,N_8412);
xor U11220 (N_11220,N_8395,N_6813);
xor U11221 (N_11221,N_8423,N_8477);
xor U11222 (N_11222,N_8449,N_6882);
or U11223 (N_11223,N_6806,N_7036);
nand U11224 (N_11224,N_8438,N_8205);
and U11225 (N_11225,N_6234,N_8116);
xnor U11226 (N_11226,N_8700,N_6196);
or U11227 (N_11227,N_7646,N_7749);
and U11228 (N_11228,N_7269,N_7718);
or U11229 (N_11229,N_7450,N_7889);
nor U11230 (N_11230,N_6225,N_7225);
nor U11231 (N_11231,N_8706,N_8606);
nand U11232 (N_11232,N_6309,N_6608);
nor U11233 (N_11233,N_6691,N_7658);
and U11234 (N_11234,N_7639,N_6811);
xor U11235 (N_11235,N_7073,N_7116);
nand U11236 (N_11236,N_7639,N_8601);
xor U11237 (N_11237,N_8064,N_6023);
xor U11238 (N_11238,N_8748,N_6455);
xor U11239 (N_11239,N_8458,N_8920);
and U11240 (N_11240,N_7450,N_7100);
or U11241 (N_11241,N_6557,N_7424);
nor U11242 (N_11242,N_6997,N_6311);
or U11243 (N_11243,N_6404,N_7616);
nand U11244 (N_11244,N_8973,N_7992);
xnor U11245 (N_11245,N_7341,N_6331);
nor U11246 (N_11246,N_8171,N_8385);
or U11247 (N_11247,N_6617,N_8464);
and U11248 (N_11248,N_8073,N_6940);
nor U11249 (N_11249,N_7576,N_8541);
nand U11250 (N_11250,N_6903,N_6934);
nor U11251 (N_11251,N_8539,N_6941);
and U11252 (N_11252,N_6672,N_6360);
and U11253 (N_11253,N_6493,N_6046);
nand U11254 (N_11254,N_7544,N_8601);
nor U11255 (N_11255,N_8992,N_6290);
and U11256 (N_11256,N_7402,N_7589);
or U11257 (N_11257,N_6966,N_6453);
nand U11258 (N_11258,N_8759,N_8672);
or U11259 (N_11259,N_7218,N_7485);
and U11260 (N_11260,N_6016,N_7136);
nand U11261 (N_11261,N_6450,N_6794);
nor U11262 (N_11262,N_8122,N_8612);
nand U11263 (N_11263,N_7919,N_6927);
nor U11264 (N_11264,N_7322,N_7083);
nor U11265 (N_11265,N_6593,N_8269);
or U11266 (N_11266,N_6874,N_8599);
nand U11267 (N_11267,N_6419,N_8829);
nand U11268 (N_11268,N_8915,N_7768);
or U11269 (N_11269,N_6215,N_8699);
nand U11270 (N_11270,N_6097,N_8527);
nor U11271 (N_11271,N_6730,N_8240);
or U11272 (N_11272,N_7449,N_6083);
or U11273 (N_11273,N_8747,N_6779);
nor U11274 (N_11274,N_6515,N_8324);
xnor U11275 (N_11275,N_6710,N_8340);
nor U11276 (N_11276,N_6335,N_6558);
nand U11277 (N_11277,N_6185,N_6794);
and U11278 (N_11278,N_8391,N_6614);
nor U11279 (N_11279,N_8567,N_8909);
and U11280 (N_11280,N_6457,N_6504);
xnor U11281 (N_11281,N_8523,N_8642);
nor U11282 (N_11282,N_8384,N_6242);
and U11283 (N_11283,N_7635,N_8171);
nor U11284 (N_11284,N_8134,N_6433);
or U11285 (N_11285,N_8787,N_8618);
xor U11286 (N_11286,N_6631,N_8848);
or U11287 (N_11287,N_7504,N_6707);
xor U11288 (N_11288,N_8332,N_8870);
nor U11289 (N_11289,N_6648,N_7145);
or U11290 (N_11290,N_6263,N_7381);
or U11291 (N_11291,N_6260,N_8768);
nor U11292 (N_11292,N_6006,N_8945);
and U11293 (N_11293,N_8341,N_7319);
or U11294 (N_11294,N_8031,N_7799);
or U11295 (N_11295,N_6727,N_8138);
xor U11296 (N_11296,N_8545,N_6817);
xor U11297 (N_11297,N_8002,N_8824);
nand U11298 (N_11298,N_6236,N_8164);
nand U11299 (N_11299,N_8400,N_6066);
nor U11300 (N_11300,N_7240,N_8284);
xor U11301 (N_11301,N_7609,N_7902);
xnor U11302 (N_11302,N_6160,N_8545);
nand U11303 (N_11303,N_6361,N_7974);
nor U11304 (N_11304,N_8251,N_6969);
or U11305 (N_11305,N_8485,N_8592);
xor U11306 (N_11306,N_6897,N_7211);
nor U11307 (N_11307,N_7627,N_6325);
and U11308 (N_11308,N_7826,N_6063);
nand U11309 (N_11309,N_6850,N_6605);
xnor U11310 (N_11310,N_7370,N_8490);
xor U11311 (N_11311,N_6783,N_8738);
nand U11312 (N_11312,N_6109,N_8033);
xnor U11313 (N_11313,N_7585,N_8267);
or U11314 (N_11314,N_7239,N_6730);
or U11315 (N_11315,N_6253,N_6303);
and U11316 (N_11316,N_6942,N_6430);
or U11317 (N_11317,N_7305,N_7565);
nand U11318 (N_11318,N_6862,N_8119);
and U11319 (N_11319,N_6806,N_7322);
or U11320 (N_11320,N_6769,N_6471);
or U11321 (N_11321,N_8607,N_7560);
nand U11322 (N_11322,N_6603,N_7799);
and U11323 (N_11323,N_8419,N_6597);
or U11324 (N_11324,N_7535,N_7238);
or U11325 (N_11325,N_8796,N_7535);
or U11326 (N_11326,N_8061,N_8807);
or U11327 (N_11327,N_7838,N_8152);
nand U11328 (N_11328,N_8516,N_7872);
nor U11329 (N_11329,N_8017,N_6966);
xnor U11330 (N_11330,N_7104,N_8672);
or U11331 (N_11331,N_6024,N_6045);
and U11332 (N_11332,N_6828,N_7748);
nand U11333 (N_11333,N_6458,N_6763);
nand U11334 (N_11334,N_8956,N_7568);
and U11335 (N_11335,N_7817,N_6476);
or U11336 (N_11336,N_6767,N_7544);
and U11337 (N_11337,N_6784,N_7176);
xor U11338 (N_11338,N_6333,N_7102);
nor U11339 (N_11339,N_8805,N_6748);
and U11340 (N_11340,N_6894,N_7271);
nand U11341 (N_11341,N_8992,N_7324);
nand U11342 (N_11342,N_6553,N_8923);
nor U11343 (N_11343,N_7261,N_8723);
xnor U11344 (N_11344,N_6387,N_6982);
or U11345 (N_11345,N_6800,N_6388);
or U11346 (N_11346,N_8389,N_8783);
nor U11347 (N_11347,N_8676,N_7892);
nand U11348 (N_11348,N_8018,N_6176);
nand U11349 (N_11349,N_7965,N_6104);
nand U11350 (N_11350,N_8653,N_7672);
and U11351 (N_11351,N_7617,N_8518);
nor U11352 (N_11352,N_6748,N_7367);
or U11353 (N_11353,N_7142,N_7534);
xor U11354 (N_11354,N_6099,N_7002);
xor U11355 (N_11355,N_8036,N_6661);
nand U11356 (N_11356,N_8162,N_7497);
nor U11357 (N_11357,N_8980,N_7697);
nor U11358 (N_11358,N_6647,N_6890);
and U11359 (N_11359,N_8749,N_8742);
or U11360 (N_11360,N_8691,N_7538);
nand U11361 (N_11361,N_7407,N_8624);
nand U11362 (N_11362,N_8813,N_7221);
and U11363 (N_11363,N_8641,N_7912);
nand U11364 (N_11364,N_8333,N_7759);
nand U11365 (N_11365,N_7110,N_8836);
nand U11366 (N_11366,N_6071,N_7286);
and U11367 (N_11367,N_6111,N_7857);
nor U11368 (N_11368,N_7608,N_7549);
nor U11369 (N_11369,N_7491,N_7939);
and U11370 (N_11370,N_6072,N_6256);
nand U11371 (N_11371,N_6248,N_8856);
xnor U11372 (N_11372,N_8452,N_6926);
nand U11373 (N_11373,N_6082,N_8729);
or U11374 (N_11374,N_8415,N_7297);
or U11375 (N_11375,N_7879,N_8387);
nor U11376 (N_11376,N_8730,N_6685);
or U11377 (N_11377,N_7441,N_7532);
or U11378 (N_11378,N_6735,N_6023);
xor U11379 (N_11379,N_7250,N_8629);
nand U11380 (N_11380,N_7865,N_8021);
nor U11381 (N_11381,N_8297,N_7491);
nand U11382 (N_11382,N_8458,N_6953);
nand U11383 (N_11383,N_6369,N_8811);
and U11384 (N_11384,N_6462,N_7349);
nand U11385 (N_11385,N_7662,N_8501);
xnor U11386 (N_11386,N_8492,N_7521);
xnor U11387 (N_11387,N_8328,N_6219);
xor U11388 (N_11388,N_7280,N_8789);
or U11389 (N_11389,N_7341,N_7954);
or U11390 (N_11390,N_6068,N_8319);
or U11391 (N_11391,N_7577,N_6179);
nor U11392 (N_11392,N_7285,N_8560);
nand U11393 (N_11393,N_6472,N_7524);
nand U11394 (N_11394,N_8873,N_7008);
or U11395 (N_11395,N_6808,N_6756);
and U11396 (N_11396,N_6665,N_7667);
xnor U11397 (N_11397,N_8832,N_8393);
nand U11398 (N_11398,N_8328,N_6438);
xnor U11399 (N_11399,N_6049,N_7248);
and U11400 (N_11400,N_6532,N_7005);
nand U11401 (N_11401,N_8382,N_8307);
xnor U11402 (N_11402,N_6062,N_7129);
xor U11403 (N_11403,N_6306,N_8035);
xor U11404 (N_11404,N_7844,N_6255);
nand U11405 (N_11405,N_7256,N_6974);
or U11406 (N_11406,N_8797,N_7286);
nor U11407 (N_11407,N_6443,N_8332);
nand U11408 (N_11408,N_7709,N_6878);
and U11409 (N_11409,N_8717,N_6624);
nand U11410 (N_11410,N_7732,N_8900);
and U11411 (N_11411,N_6138,N_7671);
nand U11412 (N_11412,N_8633,N_7059);
or U11413 (N_11413,N_8361,N_8615);
or U11414 (N_11414,N_8619,N_8118);
nand U11415 (N_11415,N_6502,N_8923);
xnor U11416 (N_11416,N_8569,N_8439);
and U11417 (N_11417,N_6174,N_6117);
xor U11418 (N_11418,N_8541,N_6456);
xor U11419 (N_11419,N_8533,N_8923);
nand U11420 (N_11420,N_8942,N_7399);
nor U11421 (N_11421,N_6764,N_6715);
xor U11422 (N_11422,N_7297,N_8831);
xor U11423 (N_11423,N_7294,N_8610);
xor U11424 (N_11424,N_7422,N_8285);
nor U11425 (N_11425,N_7430,N_7059);
nand U11426 (N_11426,N_7511,N_6652);
or U11427 (N_11427,N_8903,N_8390);
xor U11428 (N_11428,N_7690,N_8042);
and U11429 (N_11429,N_8732,N_7505);
and U11430 (N_11430,N_6284,N_6311);
or U11431 (N_11431,N_6709,N_8971);
nor U11432 (N_11432,N_8388,N_7985);
or U11433 (N_11433,N_6825,N_8693);
xor U11434 (N_11434,N_8694,N_6183);
and U11435 (N_11435,N_8165,N_6196);
xor U11436 (N_11436,N_7145,N_8536);
or U11437 (N_11437,N_8161,N_6358);
xnor U11438 (N_11438,N_7645,N_8016);
nor U11439 (N_11439,N_6946,N_8857);
or U11440 (N_11440,N_8966,N_7481);
or U11441 (N_11441,N_7201,N_6572);
nand U11442 (N_11442,N_7768,N_7181);
nand U11443 (N_11443,N_7410,N_6186);
xnor U11444 (N_11444,N_6856,N_8139);
xor U11445 (N_11445,N_6634,N_8236);
nor U11446 (N_11446,N_7006,N_7300);
xnor U11447 (N_11447,N_7348,N_8345);
and U11448 (N_11448,N_7695,N_7794);
and U11449 (N_11449,N_7709,N_6623);
nor U11450 (N_11450,N_6959,N_7822);
xnor U11451 (N_11451,N_6703,N_8061);
or U11452 (N_11452,N_7660,N_6513);
nor U11453 (N_11453,N_6199,N_6287);
and U11454 (N_11454,N_8154,N_8147);
or U11455 (N_11455,N_6089,N_7578);
xor U11456 (N_11456,N_7621,N_7477);
or U11457 (N_11457,N_7383,N_6168);
or U11458 (N_11458,N_7631,N_6371);
or U11459 (N_11459,N_7897,N_8510);
nor U11460 (N_11460,N_6465,N_7147);
nor U11461 (N_11461,N_6526,N_7639);
nand U11462 (N_11462,N_8251,N_8672);
nor U11463 (N_11463,N_7784,N_7743);
xnor U11464 (N_11464,N_7525,N_7538);
nand U11465 (N_11465,N_6322,N_8888);
nor U11466 (N_11466,N_6338,N_8932);
xor U11467 (N_11467,N_6953,N_7872);
or U11468 (N_11468,N_8283,N_8383);
and U11469 (N_11469,N_6206,N_7768);
or U11470 (N_11470,N_7052,N_8328);
xnor U11471 (N_11471,N_6017,N_6176);
xnor U11472 (N_11472,N_6728,N_8998);
nor U11473 (N_11473,N_6458,N_7231);
nand U11474 (N_11474,N_7633,N_8987);
nand U11475 (N_11475,N_8573,N_8123);
or U11476 (N_11476,N_6673,N_6793);
xor U11477 (N_11477,N_8874,N_7719);
nor U11478 (N_11478,N_7179,N_6200);
nand U11479 (N_11479,N_7409,N_7254);
and U11480 (N_11480,N_8722,N_7751);
nand U11481 (N_11481,N_7526,N_8431);
xor U11482 (N_11482,N_7971,N_7699);
or U11483 (N_11483,N_7683,N_6399);
nand U11484 (N_11484,N_6902,N_7259);
xnor U11485 (N_11485,N_8711,N_6062);
nand U11486 (N_11486,N_7735,N_7095);
nor U11487 (N_11487,N_7464,N_6788);
nand U11488 (N_11488,N_6874,N_8227);
or U11489 (N_11489,N_6319,N_7268);
nand U11490 (N_11490,N_7451,N_7231);
xor U11491 (N_11491,N_6301,N_7867);
or U11492 (N_11492,N_6376,N_8579);
nor U11493 (N_11493,N_7562,N_7689);
nor U11494 (N_11494,N_7312,N_8054);
nand U11495 (N_11495,N_7940,N_6422);
xor U11496 (N_11496,N_6080,N_6763);
nor U11497 (N_11497,N_7633,N_8830);
nand U11498 (N_11498,N_6455,N_7455);
nand U11499 (N_11499,N_8841,N_6546);
or U11500 (N_11500,N_7993,N_6250);
xor U11501 (N_11501,N_8072,N_7515);
or U11502 (N_11502,N_7514,N_6641);
nand U11503 (N_11503,N_6886,N_7532);
nor U11504 (N_11504,N_7831,N_7692);
and U11505 (N_11505,N_8659,N_8067);
and U11506 (N_11506,N_6140,N_8409);
or U11507 (N_11507,N_8030,N_6897);
and U11508 (N_11508,N_8867,N_6894);
nand U11509 (N_11509,N_7516,N_6678);
nor U11510 (N_11510,N_8862,N_6133);
and U11511 (N_11511,N_8337,N_7244);
or U11512 (N_11512,N_6548,N_7346);
nand U11513 (N_11513,N_7158,N_6530);
nor U11514 (N_11514,N_6161,N_6149);
xnor U11515 (N_11515,N_6295,N_7675);
nor U11516 (N_11516,N_8275,N_6900);
nand U11517 (N_11517,N_6246,N_8278);
or U11518 (N_11518,N_8709,N_8291);
and U11519 (N_11519,N_7276,N_8430);
xor U11520 (N_11520,N_7216,N_8583);
and U11521 (N_11521,N_7309,N_8286);
or U11522 (N_11522,N_8633,N_7766);
and U11523 (N_11523,N_6465,N_7323);
nor U11524 (N_11524,N_8722,N_8408);
xor U11525 (N_11525,N_8553,N_7731);
xor U11526 (N_11526,N_7624,N_6780);
nand U11527 (N_11527,N_7736,N_7790);
xnor U11528 (N_11528,N_7266,N_8492);
nor U11529 (N_11529,N_6741,N_7588);
xnor U11530 (N_11530,N_7928,N_7117);
and U11531 (N_11531,N_7304,N_7204);
nor U11532 (N_11532,N_8550,N_6783);
xor U11533 (N_11533,N_7675,N_7227);
or U11534 (N_11534,N_6248,N_8271);
xor U11535 (N_11535,N_6846,N_6806);
and U11536 (N_11536,N_8485,N_7519);
xnor U11537 (N_11537,N_6612,N_7059);
nand U11538 (N_11538,N_6525,N_7853);
nand U11539 (N_11539,N_6075,N_6893);
or U11540 (N_11540,N_8305,N_6050);
xnor U11541 (N_11541,N_7515,N_8578);
nor U11542 (N_11542,N_7711,N_6619);
nor U11543 (N_11543,N_6327,N_6709);
xor U11544 (N_11544,N_7149,N_6421);
nand U11545 (N_11545,N_6334,N_8263);
nand U11546 (N_11546,N_7616,N_6094);
or U11547 (N_11547,N_7077,N_6670);
and U11548 (N_11548,N_7150,N_6841);
or U11549 (N_11549,N_7225,N_8489);
nand U11550 (N_11550,N_8501,N_7408);
nand U11551 (N_11551,N_8753,N_6050);
or U11552 (N_11552,N_8078,N_7688);
nor U11553 (N_11553,N_7926,N_7471);
xor U11554 (N_11554,N_6370,N_8543);
nand U11555 (N_11555,N_8216,N_6088);
and U11556 (N_11556,N_8107,N_8132);
and U11557 (N_11557,N_6363,N_8837);
or U11558 (N_11558,N_6254,N_6759);
xor U11559 (N_11559,N_6209,N_8722);
nor U11560 (N_11560,N_8708,N_8102);
or U11561 (N_11561,N_6968,N_6309);
nand U11562 (N_11562,N_6343,N_7551);
nor U11563 (N_11563,N_8383,N_8598);
and U11564 (N_11564,N_6014,N_7098);
or U11565 (N_11565,N_8763,N_7727);
and U11566 (N_11566,N_8776,N_8570);
xnor U11567 (N_11567,N_8507,N_8555);
nor U11568 (N_11568,N_8294,N_7798);
xnor U11569 (N_11569,N_8394,N_8116);
nand U11570 (N_11570,N_7623,N_7041);
or U11571 (N_11571,N_8893,N_7682);
or U11572 (N_11572,N_6951,N_6539);
nand U11573 (N_11573,N_7125,N_8594);
and U11574 (N_11574,N_6463,N_8106);
or U11575 (N_11575,N_8571,N_8632);
xnor U11576 (N_11576,N_6556,N_6702);
nor U11577 (N_11577,N_7220,N_6494);
nand U11578 (N_11578,N_8055,N_6677);
or U11579 (N_11579,N_8149,N_7006);
or U11580 (N_11580,N_7748,N_8680);
and U11581 (N_11581,N_6303,N_6239);
nand U11582 (N_11582,N_7754,N_7006);
nand U11583 (N_11583,N_6521,N_8391);
or U11584 (N_11584,N_6201,N_7830);
xor U11585 (N_11585,N_8336,N_6636);
and U11586 (N_11586,N_6099,N_7106);
and U11587 (N_11587,N_8322,N_6985);
or U11588 (N_11588,N_7389,N_6373);
xnor U11589 (N_11589,N_6704,N_6830);
xor U11590 (N_11590,N_6721,N_8910);
nand U11591 (N_11591,N_7439,N_7773);
xnor U11592 (N_11592,N_8043,N_8885);
or U11593 (N_11593,N_8599,N_8762);
nand U11594 (N_11594,N_6516,N_7353);
and U11595 (N_11595,N_7531,N_6068);
or U11596 (N_11596,N_6609,N_8803);
and U11597 (N_11597,N_8818,N_6045);
nor U11598 (N_11598,N_7218,N_8760);
xnor U11599 (N_11599,N_7797,N_6214);
and U11600 (N_11600,N_7969,N_6677);
and U11601 (N_11601,N_7518,N_6270);
nand U11602 (N_11602,N_7973,N_6306);
xnor U11603 (N_11603,N_8674,N_7407);
nand U11604 (N_11604,N_8765,N_8471);
nor U11605 (N_11605,N_8453,N_6825);
or U11606 (N_11606,N_8391,N_6570);
nor U11607 (N_11607,N_8970,N_6196);
nor U11608 (N_11608,N_6032,N_6753);
nor U11609 (N_11609,N_7934,N_7973);
nor U11610 (N_11610,N_6244,N_6080);
and U11611 (N_11611,N_8894,N_8275);
nor U11612 (N_11612,N_6992,N_6936);
nor U11613 (N_11613,N_6579,N_7260);
or U11614 (N_11614,N_6409,N_6770);
or U11615 (N_11615,N_7107,N_8926);
nand U11616 (N_11616,N_7726,N_6273);
and U11617 (N_11617,N_7786,N_7367);
and U11618 (N_11618,N_7139,N_7739);
and U11619 (N_11619,N_7142,N_8163);
nand U11620 (N_11620,N_8700,N_8846);
or U11621 (N_11621,N_6155,N_8481);
or U11622 (N_11622,N_6888,N_7947);
and U11623 (N_11623,N_7945,N_8831);
or U11624 (N_11624,N_8021,N_8535);
nor U11625 (N_11625,N_7841,N_8945);
or U11626 (N_11626,N_8624,N_8703);
xor U11627 (N_11627,N_6185,N_7005);
or U11628 (N_11628,N_6244,N_7381);
or U11629 (N_11629,N_6680,N_6781);
or U11630 (N_11630,N_8727,N_6390);
nand U11631 (N_11631,N_7226,N_8122);
xor U11632 (N_11632,N_6866,N_6663);
nor U11633 (N_11633,N_7878,N_8209);
nand U11634 (N_11634,N_8674,N_6849);
nand U11635 (N_11635,N_7247,N_6725);
xor U11636 (N_11636,N_8155,N_6018);
or U11637 (N_11637,N_8042,N_7644);
nor U11638 (N_11638,N_8438,N_8796);
or U11639 (N_11639,N_8999,N_8100);
nor U11640 (N_11640,N_7630,N_6067);
nand U11641 (N_11641,N_6819,N_8469);
nand U11642 (N_11642,N_6782,N_8541);
nor U11643 (N_11643,N_6901,N_7491);
xnor U11644 (N_11644,N_8835,N_6313);
and U11645 (N_11645,N_7511,N_8847);
nor U11646 (N_11646,N_6474,N_6720);
nand U11647 (N_11647,N_8971,N_8009);
xor U11648 (N_11648,N_6177,N_7187);
nand U11649 (N_11649,N_8939,N_8253);
xnor U11650 (N_11650,N_7640,N_7880);
nor U11651 (N_11651,N_8869,N_7207);
nand U11652 (N_11652,N_8890,N_8802);
nor U11653 (N_11653,N_8378,N_8268);
or U11654 (N_11654,N_8446,N_7615);
and U11655 (N_11655,N_8044,N_7400);
or U11656 (N_11656,N_6730,N_8376);
xnor U11657 (N_11657,N_6154,N_6116);
nand U11658 (N_11658,N_7308,N_6204);
nand U11659 (N_11659,N_7255,N_8752);
or U11660 (N_11660,N_8697,N_8876);
nor U11661 (N_11661,N_6606,N_7098);
nor U11662 (N_11662,N_6735,N_6314);
nand U11663 (N_11663,N_7108,N_6078);
nand U11664 (N_11664,N_6443,N_8939);
nand U11665 (N_11665,N_6625,N_6442);
xor U11666 (N_11666,N_7779,N_7633);
xor U11667 (N_11667,N_6381,N_8786);
and U11668 (N_11668,N_6416,N_7312);
nor U11669 (N_11669,N_7390,N_8452);
nor U11670 (N_11670,N_7626,N_7776);
and U11671 (N_11671,N_6098,N_8621);
nor U11672 (N_11672,N_8248,N_7003);
or U11673 (N_11673,N_6962,N_6984);
and U11674 (N_11674,N_6208,N_7755);
xnor U11675 (N_11675,N_8210,N_8368);
xnor U11676 (N_11676,N_8561,N_6379);
or U11677 (N_11677,N_6867,N_8002);
xnor U11678 (N_11678,N_8895,N_8903);
xnor U11679 (N_11679,N_7241,N_7285);
xnor U11680 (N_11680,N_8081,N_6051);
nor U11681 (N_11681,N_8544,N_6785);
nor U11682 (N_11682,N_7329,N_7594);
and U11683 (N_11683,N_6794,N_7309);
nand U11684 (N_11684,N_6786,N_7228);
or U11685 (N_11685,N_6722,N_7807);
or U11686 (N_11686,N_6021,N_6208);
xnor U11687 (N_11687,N_6345,N_7745);
xor U11688 (N_11688,N_8283,N_7762);
xnor U11689 (N_11689,N_6140,N_8940);
xor U11690 (N_11690,N_6548,N_8695);
nand U11691 (N_11691,N_8231,N_8454);
and U11692 (N_11692,N_7591,N_7241);
and U11693 (N_11693,N_7432,N_8156);
and U11694 (N_11694,N_7036,N_6829);
nor U11695 (N_11695,N_7249,N_6208);
xor U11696 (N_11696,N_7140,N_8106);
nor U11697 (N_11697,N_8704,N_7770);
nand U11698 (N_11698,N_7028,N_6830);
nor U11699 (N_11699,N_7513,N_7137);
xnor U11700 (N_11700,N_8580,N_8799);
or U11701 (N_11701,N_8599,N_7307);
or U11702 (N_11702,N_7855,N_8341);
and U11703 (N_11703,N_8243,N_6570);
xor U11704 (N_11704,N_7689,N_7509);
or U11705 (N_11705,N_7584,N_7626);
nor U11706 (N_11706,N_7309,N_6008);
and U11707 (N_11707,N_7643,N_7372);
and U11708 (N_11708,N_7766,N_6409);
or U11709 (N_11709,N_7801,N_6622);
xor U11710 (N_11710,N_8129,N_6821);
xnor U11711 (N_11711,N_8952,N_6118);
xnor U11712 (N_11712,N_7923,N_6166);
nor U11713 (N_11713,N_7358,N_6479);
nor U11714 (N_11714,N_7782,N_8210);
and U11715 (N_11715,N_7732,N_7255);
nor U11716 (N_11716,N_7164,N_7806);
or U11717 (N_11717,N_7041,N_6769);
or U11718 (N_11718,N_8962,N_8310);
or U11719 (N_11719,N_7847,N_6541);
and U11720 (N_11720,N_8214,N_8736);
xor U11721 (N_11721,N_8802,N_8111);
or U11722 (N_11722,N_6046,N_7104);
and U11723 (N_11723,N_8889,N_6657);
nand U11724 (N_11724,N_6180,N_7766);
or U11725 (N_11725,N_7877,N_6900);
and U11726 (N_11726,N_7529,N_6379);
nor U11727 (N_11727,N_7699,N_8184);
or U11728 (N_11728,N_6679,N_8358);
xor U11729 (N_11729,N_6924,N_6377);
xor U11730 (N_11730,N_8887,N_7577);
nand U11731 (N_11731,N_6181,N_7200);
or U11732 (N_11732,N_6655,N_6734);
xnor U11733 (N_11733,N_8402,N_6105);
xnor U11734 (N_11734,N_8964,N_6996);
nor U11735 (N_11735,N_7322,N_6305);
nand U11736 (N_11736,N_8725,N_6567);
or U11737 (N_11737,N_6946,N_7783);
nand U11738 (N_11738,N_6778,N_6011);
nor U11739 (N_11739,N_8129,N_8888);
xor U11740 (N_11740,N_7420,N_6707);
and U11741 (N_11741,N_7263,N_8059);
nand U11742 (N_11742,N_7064,N_8456);
xnor U11743 (N_11743,N_6001,N_7157);
xnor U11744 (N_11744,N_8260,N_6845);
nand U11745 (N_11745,N_8011,N_6157);
nor U11746 (N_11746,N_7965,N_6513);
or U11747 (N_11747,N_8651,N_8236);
and U11748 (N_11748,N_7759,N_6696);
or U11749 (N_11749,N_7791,N_8465);
or U11750 (N_11750,N_7995,N_7807);
or U11751 (N_11751,N_8620,N_8576);
xnor U11752 (N_11752,N_8832,N_6235);
nand U11753 (N_11753,N_6061,N_7415);
or U11754 (N_11754,N_8429,N_8935);
nand U11755 (N_11755,N_7660,N_7446);
nor U11756 (N_11756,N_6566,N_7297);
and U11757 (N_11757,N_6199,N_7490);
and U11758 (N_11758,N_6472,N_8128);
and U11759 (N_11759,N_7991,N_6236);
nand U11760 (N_11760,N_7848,N_6756);
nand U11761 (N_11761,N_7505,N_6851);
nor U11762 (N_11762,N_8876,N_8705);
and U11763 (N_11763,N_7662,N_7402);
nor U11764 (N_11764,N_8522,N_6737);
nor U11765 (N_11765,N_6235,N_7320);
or U11766 (N_11766,N_7887,N_7016);
nor U11767 (N_11767,N_8598,N_8722);
xnor U11768 (N_11768,N_6596,N_7320);
and U11769 (N_11769,N_7978,N_6079);
and U11770 (N_11770,N_8116,N_6219);
or U11771 (N_11771,N_7362,N_8015);
nand U11772 (N_11772,N_8579,N_8092);
nor U11773 (N_11773,N_8080,N_7120);
or U11774 (N_11774,N_6224,N_8502);
or U11775 (N_11775,N_7952,N_7505);
nand U11776 (N_11776,N_8828,N_8275);
nand U11777 (N_11777,N_6532,N_8531);
nand U11778 (N_11778,N_8322,N_6432);
xor U11779 (N_11779,N_6386,N_7703);
nor U11780 (N_11780,N_8603,N_8528);
xor U11781 (N_11781,N_8601,N_8010);
and U11782 (N_11782,N_6349,N_6898);
or U11783 (N_11783,N_8973,N_7650);
nor U11784 (N_11784,N_7351,N_6174);
or U11785 (N_11785,N_6596,N_8433);
nor U11786 (N_11786,N_7244,N_7769);
nor U11787 (N_11787,N_6971,N_6513);
nor U11788 (N_11788,N_8759,N_6315);
nor U11789 (N_11789,N_8267,N_7098);
nor U11790 (N_11790,N_8495,N_8413);
nor U11791 (N_11791,N_7492,N_6490);
and U11792 (N_11792,N_8661,N_7040);
and U11793 (N_11793,N_6551,N_7585);
and U11794 (N_11794,N_6757,N_8994);
and U11795 (N_11795,N_8498,N_6077);
xnor U11796 (N_11796,N_6103,N_8633);
xor U11797 (N_11797,N_7870,N_8884);
or U11798 (N_11798,N_7877,N_7029);
xnor U11799 (N_11799,N_6707,N_8926);
and U11800 (N_11800,N_7882,N_7084);
or U11801 (N_11801,N_8962,N_6408);
or U11802 (N_11802,N_6461,N_6728);
and U11803 (N_11803,N_6843,N_7135);
nand U11804 (N_11804,N_6548,N_7745);
or U11805 (N_11805,N_6161,N_6233);
xor U11806 (N_11806,N_8617,N_6568);
nor U11807 (N_11807,N_7778,N_6879);
xor U11808 (N_11808,N_7771,N_7030);
nand U11809 (N_11809,N_6108,N_7585);
nand U11810 (N_11810,N_7681,N_8784);
nor U11811 (N_11811,N_6632,N_8482);
nor U11812 (N_11812,N_6582,N_7870);
nand U11813 (N_11813,N_6901,N_8196);
nand U11814 (N_11814,N_8035,N_8685);
and U11815 (N_11815,N_7708,N_8386);
or U11816 (N_11816,N_8991,N_7786);
or U11817 (N_11817,N_7019,N_6061);
or U11818 (N_11818,N_8228,N_6769);
xor U11819 (N_11819,N_7599,N_7462);
and U11820 (N_11820,N_7793,N_6791);
nor U11821 (N_11821,N_6164,N_7520);
and U11822 (N_11822,N_8407,N_8120);
and U11823 (N_11823,N_6105,N_7890);
nor U11824 (N_11824,N_6437,N_7970);
nand U11825 (N_11825,N_8793,N_6325);
nand U11826 (N_11826,N_6583,N_6031);
and U11827 (N_11827,N_6102,N_7276);
nor U11828 (N_11828,N_8480,N_6014);
nor U11829 (N_11829,N_7336,N_8815);
and U11830 (N_11830,N_6163,N_7536);
xor U11831 (N_11831,N_8998,N_7460);
or U11832 (N_11832,N_6291,N_7722);
nor U11833 (N_11833,N_7941,N_8587);
nand U11834 (N_11834,N_8412,N_6458);
xor U11835 (N_11835,N_7032,N_7450);
or U11836 (N_11836,N_7246,N_8954);
nand U11837 (N_11837,N_7216,N_8472);
nor U11838 (N_11838,N_7203,N_7573);
or U11839 (N_11839,N_7345,N_6383);
nand U11840 (N_11840,N_7754,N_8421);
and U11841 (N_11841,N_8947,N_6909);
or U11842 (N_11842,N_8164,N_6365);
and U11843 (N_11843,N_6269,N_6816);
nor U11844 (N_11844,N_8823,N_7517);
nor U11845 (N_11845,N_6890,N_6961);
or U11846 (N_11846,N_6399,N_8912);
or U11847 (N_11847,N_7010,N_7300);
and U11848 (N_11848,N_7380,N_8832);
xor U11849 (N_11849,N_8481,N_8523);
or U11850 (N_11850,N_7694,N_8137);
nand U11851 (N_11851,N_6082,N_6434);
nand U11852 (N_11852,N_7301,N_7037);
nand U11853 (N_11853,N_6632,N_8643);
xnor U11854 (N_11854,N_8632,N_8151);
or U11855 (N_11855,N_8218,N_6400);
and U11856 (N_11856,N_8353,N_7426);
nand U11857 (N_11857,N_6607,N_6182);
and U11858 (N_11858,N_7937,N_7856);
nand U11859 (N_11859,N_7481,N_7784);
xnor U11860 (N_11860,N_6631,N_6786);
nor U11861 (N_11861,N_8262,N_8413);
and U11862 (N_11862,N_7274,N_6065);
nand U11863 (N_11863,N_8852,N_7917);
or U11864 (N_11864,N_7352,N_8469);
xnor U11865 (N_11865,N_6157,N_8315);
nand U11866 (N_11866,N_8780,N_8473);
and U11867 (N_11867,N_8626,N_7301);
nor U11868 (N_11868,N_7541,N_6246);
and U11869 (N_11869,N_7338,N_6642);
xnor U11870 (N_11870,N_6971,N_6118);
and U11871 (N_11871,N_7684,N_8923);
or U11872 (N_11872,N_7872,N_8277);
xor U11873 (N_11873,N_6443,N_6448);
or U11874 (N_11874,N_7475,N_8488);
and U11875 (N_11875,N_6476,N_7005);
and U11876 (N_11876,N_7104,N_7761);
nand U11877 (N_11877,N_6447,N_8177);
or U11878 (N_11878,N_6001,N_7520);
and U11879 (N_11879,N_6577,N_7975);
or U11880 (N_11880,N_7054,N_8266);
nand U11881 (N_11881,N_6805,N_8170);
and U11882 (N_11882,N_6160,N_8864);
nor U11883 (N_11883,N_6394,N_8182);
or U11884 (N_11884,N_8840,N_8952);
nor U11885 (N_11885,N_6516,N_6260);
xor U11886 (N_11886,N_8239,N_6766);
and U11887 (N_11887,N_8707,N_8306);
and U11888 (N_11888,N_8981,N_8260);
and U11889 (N_11889,N_8744,N_6055);
and U11890 (N_11890,N_8850,N_6441);
and U11891 (N_11891,N_7392,N_6007);
or U11892 (N_11892,N_8144,N_7482);
nor U11893 (N_11893,N_8839,N_6908);
and U11894 (N_11894,N_6789,N_7270);
or U11895 (N_11895,N_8239,N_7643);
nand U11896 (N_11896,N_8582,N_6216);
nor U11897 (N_11897,N_7196,N_8696);
xnor U11898 (N_11898,N_7722,N_8248);
xor U11899 (N_11899,N_7371,N_7585);
or U11900 (N_11900,N_7568,N_8621);
xnor U11901 (N_11901,N_8933,N_7869);
or U11902 (N_11902,N_8982,N_7914);
xnor U11903 (N_11903,N_6338,N_7379);
or U11904 (N_11904,N_6197,N_7305);
and U11905 (N_11905,N_7075,N_6339);
xor U11906 (N_11906,N_8502,N_8442);
and U11907 (N_11907,N_8907,N_6651);
and U11908 (N_11908,N_8440,N_8426);
nand U11909 (N_11909,N_7262,N_6914);
nand U11910 (N_11910,N_8651,N_7064);
and U11911 (N_11911,N_7928,N_7846);
nand U11912 (N_11912,N_7175,N_7196);
nand U11913 (N_11913,N_7598,N_8986);
or U11914 (N_11914,N_8344,N_8026);
or U11915 (N_11915,N_6089,N_7060);
xor U11916 (N_11916,N_7419,N_7907);
or U11917 (N_11917,N_7316,N_8659);
and U11918 (N_11918,N_8461,N_8549);
or U11919 (N_11919,N_6387,N_6595);
and U11920 (N_11920,N_6425,N_6588);
nand U11921 (N_11921,N_7589,N_6927);
or U11922 (N_11922,N_8302,N_7296);
xnor U11923 (N_11923,N_7102,N_8449);
xnor U11924 (N_11924,N_8556,N_8350);
xnor U11925 (N_11925,N_7848,N_7586);
xor U11926 (N_11926,N_7421,N_6623);
xor U11927 (N_11927,N_7772,N_6110);
or U11928 (N_11928,N_6500,N_7325);
nand U11929 (N_11929,N_7239,N_8378);
or U11930 (N_11930,N_8381,N_8789);
or U11931 (N_11931,N_8626,N_8461);
and U11932 (N_11932,N_7052,N_7067);
or U11933 (N_11933,N_7416,N_7670);
and U11934 (N_11934,N_7970,N_8074);
and U11935 (N_11935,N_8921,N_6469);
and U11936 (N_11936,N_8008,N_8672);
and U11937 (N_11937,N_6726,N_6252);
xnor U11938 (N_11938,N_7918,N_7581);
or U11939 (N_11939,N_6711,N_8112);
nor U11940 (N_11940,N_7685,N_8259);
nor U11941 (N_11941,N_7738,N_6851);
xor U11942 (N_11942,N_6645,N_7396);
nand U11943 (N_11943,N_6984,N_8821);
nand U11944 (N_11944,N_6035,N_6815);
nand U11945 (N_11945,N_8099,N_8736);
nor U11946 (N_11946,N_8842,N_6002);
nand U11947 (N_11947,N_6705,N_7674);
or U11948 (N_11948,N_8654,N_6159);
xor U11949 (N_11949,N_6428,N_6426);
xnor U11950 (N_11950,N_6168,N_7671);
and U11951 (N_11951,N_8664,N_7524);
xnor U11952 (N_11952,N_6947,N_7526);
xor U11953 (N_11953,N_8807,N_7978);
xnor U11954 (N_11954,N_7071,N_8906);
nor U11955 (N_11955,N_6240,N_6874);
xnor U11956 (N_11956,N_8168,N_6628);
nor U11957 (N_11957,N_6930,N_8078);
nor U11958 (N_11958,N_6037,N_7640);
xnor U11959 (N_11959,N_7231,N_6384);
nor U11960 (N_11960,N_7604,N_7665);
xor U11961 (N_11961,N_6222,N_6533);
nand U11962 (N_11962,N_7867,N_7569);
or U11963 (N_11963,N_8725,N_6621);
xor U11964 (N_11964,N_6586,N_8977);
xor U11965 (N_11965,N_7030,N_6688);
nand U11966 (N_11966,N_7604,N_7486);
xor U11967 (N_11967,N_6784,N_7986);
xor U11968 (N_11968,N_6260,N_7318);
and U11969 (N_11969,N_8231,N_7390);
nand U11970 (N_11970,N_6803,N_7265);
or U11971 (N_11971,N_6887,N_6050);
and U11972 (N_11972,N_7506,N_7052);
and U11973 (N_11973,N_6806,N_6042);
nand U11974 (N_11974,N_6329,N_7026);
and U11975 (N_11975,N_6757,N_6840);
nor U11976 (N_11976,N_6569,N_6529);
xor U11977 (N_11977,N_6619,N_6073);
nand U11978 (N_11978,N_7375,N_6183);
nand U11979 (N_11979,N_6472,N_6197);
nor U11980 (N_11980,N_8404,N_7981);
and U11981 (N_11981,N_6493,N_6178);
nand U11982 (N_11982,N_8166,N_7833);
nor U11983 (N_11983,N_8737,N_6629);
nor U11984 (N_11984,N_7788,N_8496);
and U11985 (N_11985,N_7531,N_6022);
xnor U11986 (N_11986,N_7472,N_7863);
or U11987 (N_11987,N_6382,N_7992);
nor U11988 (N_11988,N_6335,N_8814);
or U11989 (N_11989,N_7272,N_8315);
nand U11990 (N_11990,N_6822,N_6305);
and U11991 (N_11991,N_7435,N_8524);
xnor U11992 (N_11992,N_6260,N_6584);
nor U11993 (N_11993,N_6341,N_6389);
nand U11994 (N_11994,N_7258,N_6537);
nand U11995 (N_11995,N_7820,N_8092);
nor U11996 (N_11996,N_8609,N_8399);
and U11997 (N_11997,N_6566,N_7737);
nand U11998 (N_11998,N_7170,N_6026);
xnor U11999 (N_11999,N_6099,N_6246);
or U12000 (N_12000,N_10079,N_10747);
or U12001 (N_12001,N_11455,N_10737);
and U12002 (N_12002,N_11653,N_11382);
nand U12003 (N_12003,N_10617,N_9976);
and U12004 (N_12004,N_11631,N_11358);
xor U12005 (N_12005,N_9490,N_11868);
nand U12006 (N_12006,N_11585,N_10812);
or U12007 (N_12007,N_10135,N_11884);
or U12008 (N_12008,N_11371,N_10141);
xnor U12009 (N_12009,N_11827,N_11370);
and U12010 (N_12010,N_10901,N_10526);
or U12011 (N_12011,N_9028,N_11399);
xnor U12012 (N_12012,N_9732,N_10438);
nor U12013 (N_12013,N_11964,N_9434);
nor U12014 (N_12014,N_9524,N_11240);
xor U12015 (N_12015,N_10582,N_11211);
xor U12016 (N_12016,N_10293,N_10204);
xnor U12017 (N_12017,N_10058,N_11608);
xor U12018 (N_12018,N_9377,N_10382);
or U12019 (N_12019,N_10757,N_11084);
nor U12020 (N_12020,N_10097,N_9542);
nor U12021 (N_12021,N_9279,N_10252);
nor U12022 (N_12022,N_11496,N_9849);
and U12023 (N_12023,N_9906,N_10859);
and U12024 (N_12024,N_11584,N_11269);
nand U12025 (N_12025,N_11525,N_10938);
and U12026 (N_12026,N_9128,N_11580);
or U12027 (N_12027,N_11736,N_10697);
or U12028 (N_12028,N_10815,N_9010);
xnor U12029 (N_12029,N_11010,N_9289);
nor U12030 (N_12030,N_9192,N_9201);
or U12031 (N_12031,N_9474,N_10499);
nand U12032 (N_12032,N_10249,N_9553);
nor U12033 (N_12033,N_9773,N_10299);
or U12034 (N_12034,N_11095,N_9485);
nor U12035 (N_12035,N_11014,N_10885);
nor U12036 (N_12036,N_10422,N_11122);
nor U12037 (N_12037,N_10715,N_10969);
nand U12038 (N_12038,N_9903,N_9642);
nand U12039 (N_12039,N_10955,N_11688);
or U12040 (N_12040,N_9470,N_10831);
or U12041 (N_12041,N_9125,N_11899);
and U12042 (N_12042,N_9369,N_10552);
nor U12043 (N_12043,N_11731,N_10056);
nor U12044 (N_12044,N_10026,N_9562);
nand U12045 (N_12045,N_9082,N_10709);
or U12046 (N_12046,N_10842,N_11949);
and U12047 (N_12047,N_10661,N_10770);
or U12048 (N_12048,N_9647,N_9902);
xnor U12049 (N_12049,N_11882,N_11217);
nand U12050 (N_12050,N_9971,N_10295);
and U12051 (N_12051,N_9735,N_9393);
nand U12052 (N_12052,N_9725,N_11924);
nand U12053 (N_12053,N_10763,N_10896);
nor U12054 (N_12054,N_10194,N_9857);
or U12055 (N_12055,N_9568,N_10279);
xnor U12056 (N_12056,N_10017,N_9448);
nor U12057 (N_12057,N_11792,N_9364);
nor U12058 (N_12058,N_9968,N_11001);
xor U12059 (N_12059,N_10558,N_9919);
nand U12060 (N_12060,N_10045,N_9339);
nor U12061 (N_12061,N_9106,N_10577);
nand U12062 (N_12062,N_9811,N_9365);
nand U12063 (N_12063,N_11681,N_10137);
or U12064 (N_12064,N_10553,N_11454);
and U12065 (N_12065,N_9038,N_10450);
or U12066 (N_12066,N_11694,N_10121);
nand U12067 (N_12067,N_9331,N_10443);
or U12068 (N_12068,N_9931,N_9037);
nand U12069 (N_12069,N_9698,N_10483);
xnor U12070 (N_12070,N_10472,N_9834);
nand U12071 (N_12071,N_10992,N_11194);
xnor U12072 (N_12072,N_10177,N_11288);
nand U12073 (N_12073,N_10865,N_11247);
nor U12074 (N_12074,N_9679,N_11163);
and U12075 (N_12075,N_11669,N_10309);
nand U12076 (N_12076,N_9382,N_10801);
xor U12077 (N_12077,N_10030,N_9414);
and U12078 (N_12078,N_11775,N_9572);
or U12079 (N_12079,N_11283,N_10639);
nor U12080 (N_12080,N_11146,N_9652);
nor U12081 (N_12081,N_11875,N_11168);
xnor U12082 (N_12082,N_11975,N_11630);
and U12083 (N_12083,N_9317,N_10853);
and U12084 (N_12084,N_10966,N_11767);
nor U12085 (N_12085,N_10819,N_10287);
and U12086 (N_12086,N_9676,N_11241);
nand U12087 (N_12087,N_11192,N_10620);
nand U12088 (N_12088,N_9205,N_11396);
or U12089 (N_12089,N_9162,N_10457);
nand U12090 (N_12090,N_9439,N_11696);
xor U12091 (N_12091,N_11139,N_11150);
nor U12092 (N_12092,N_10386,N_11453);
nand U12093 (N_12093,N_10234,N_11250);
and U12094 (N_12094,N_9027,N_11867);
xnor U12095 (N_12095,N_9326,N_10367);
and U12096 (N_12096,N_11013,N_9189);
or U12097 (N_12097,N_10425,N_10888);
or U12098 (N_12098,N_9661,N_9061);
and U12099 (N_12099,N_10485,N_9210);
nand U12100 (N_12100,N_10108,N_10767);
or U12101 (N_12101,N_9353,N_9251);
nor U12102 (N_12102,N_11404,N_11801);
xor U12103 (N_12103,N_9874,N_11213);
xnor U12104 (N_12104,N_10434,N_11027);
nor U12105 (N_12105,N_11215,N_10439);
and U12106 (N_12106,N_11278,N_9825);
or U12107 (N_12107,N_11711,N_9686);
or U12108 (N_12108,N_9323,N_10729);
and U12109 (N_12109,N_9965,N_10075);
nand U12110 (N_12110,N_10481,N_10968);
nand U12111 (N_12111,N_11935,N_11167);
xor U12112 (N_12112,N_10740,N_11155);
or U12113 (N_12113,N_11860,N_9085);
or U12114 (N_12114,N_10406,N_9993);
nor U12115 (N_12115,N_10585,N_11892);
xor U12116 (N_12116,N_9079,N_10758);
xor U12117 (N_12117,N_10925,N_9822);
or U12118 (N_12118,N_11305,N_9612);
and U12119 (N_12119,N_10324,N_9445);
and U12120 (N_12120,N_11545,N_9321);
and U12121 (N_12121,N_11502,N_10214);
and U12122 (N_12122,N_10847,N_11579);
nor U12123 (N_12123,N_10496,N_10197);
and U12124 (N_12124,N_9113,N_11761);
or U12125 (N_12125,N_11577,N_9454);
xor U12126 (N_12126,N_11109,N_10903);
nor U12127 (N_12127,N_9748,N_11210);
and U12128 (N_12128,N_10836,N_10002);
nor U12129 (N_12129,N_10733,N_10724);
or U12130 (N_12130,N_10142,N_10061);
or U12131 (N_12131,N_11733,N_10818);
nor U12132 (N_12132,N_9300,N_10402);
and U12133 (N_12133,N_11800,N_11770);
xor U12134 (N_12134,N_11652,N_11818);
xnor U12135 (N_12135,N_9643,N_9688);
nand U12136 (N_12136,N_11642,N_10011);
or U12137 (N_12137,N_10001,N_11644);
and U12138 (N_12138,N_9549,N_10314);
xor U12139 (N_12139,N_9550,N_9759);
and U12140 (N_12140,N_9831,N_11672);
xor U12141 (N_12141,N_9699,N_10304);
nand U12142 (N_12142,N_9307,N_9928);
nand U12143 (N_12143,N_10112,N_10176);
nor U12144 (N_12144,N_9237,N_10826);
xnor U12145 (N_12145,N_9244,N_10291);
or U12146 (N_12146,N_11456,N_9386);
nand U12147 (N_12147,N_9555,N_9761);
nand U12148 (N_12148,N_10870,N_9755);
or U12149 (N_12149,N_9119,N_11402);
xor U12150 (N_12150,N_10101,N_9721);
or U12151 (N_12151,N_10361,N_10746);
nand U12152 (N_12152,N_11962,N_9540);
nor U12153 (N_12153,N_10538,N_9936);
xnor U12154 (N_12154,N_9363,N_10348);
nand U12155 (N_12155,N_11841,N_11451);
xor U12156 (N_12156,N_10677,N_11565);
or U12157 (N_12157,N_9603,N_10811);
or U12158 (N_12158,N_11203,N_9048);
and U12159 (N_12159,N_10655,N_11401);
or U12160 (N_12160,N_10940,N_10220);
and U12161 (N_12161,N_11074,N_10389);
nand U12162 (N_12162,N_9468,N_10212);
or U12163 (N_12163,N_10404,N_11259);
nand U12164 (N_12164,N_10650,N_10397);
xnor U12165 (N_12165,N_11183,N_11817);
xnor U12166 (N_12166,N_11966,N_11816);
nand U12167 (N_12167,N_10440,N_9145);
nand U12168 (N_12168,N_11160,N_10867);
xor U12169 (N_12169,N_11538,N_10630);
or U12170 (N_12170,N_11675,N_9980);
nor U12171 (N_12171,N_9990,N_10235);
and U12172 (N_12172,N_11737,N_10646);
xor U12173 (N_12173,N_11476,N_10714);
nand U12174 (N_12174,N_9019,N_10830);
xor U12175 (N_12175,N_9071,N_9973);
nand U12176 (N_12176,N_11279,N_9932);
nor U12177 (N_12177,N_11024,N_9987);
xnor U12178 (N_12178,N_9121,N_9366);
and U12179 (N_12179,N_9332,N_10446);
or U12180 (N_12180,N_10525,N_10883);
and U12181 (N_12181,N_11547,N_10890);
or U12182 (N_12182,N_9590,N_11510);
or U12183 (N_12183,N_9378,N_11106);
nor U12184 (N_12184,N_11275,N_10308);
and U12185 (N_12185,N_11133,N_9375);
nor U12186 (N_12186,N_11151,N_11003);
nand U12187 (N_12187,N_10821,N_10720);
or U12188 (N_12188,N_11632,N_10816);
nor U12189 (N_12189,N_10358,N_11338);
nor U12190 (N_12190,N_9728,N_9328);
nand U12191 (N_12191,N_11651,N_10979);
nand U12192 (N_12192,N_11888,N_9272);
and U12193 (N_12193,N_10312,N_10580);
nor U12194 (N_12194,N_11773,N_9102);
and U12195 (N_12195,N_11023,N_11286);
xnor U12196 (N_12196,N_10833,N_11484);
nand U12197 (N_12197,N_9505,N_11740);
xor U12198 (N_12198,N_10302,N_9295);
nand U12199 (N_12199,N_11216,N_10051);
nand U12200 (N_12200,N_9673,N_9632);
and U12201 (N_12201,N_9765,N_10791);
and U12202 (N_12202,N_9538,N_10512);
nand U12203 (N_12203,N_9335,N_11497);
nor U12204 (N_12204,N_9194,N_11755);
nor U12205 (N_12205,N_11504,N_9527);
or U12206 (N_12206,N_10921,N_9742);
or U12207 (N_12207,N_9704,N_10834);
xnor U12208 (N_12208,N_10046,N_9062);
xor U12209 (N_12209,N_10572,N_11610);
or U12210 (N_12210,N_11065,N_11578);
nand U12211 (N_12211,N_9737,N_9978);
nand U12212 (N_12212,N_9690,N_11965);
xnor U12213 (N_12213,N_10511,N_10687);
nor U12214 (N_12214,N_11274,N_11529);
and U12215 (N_12215,N_11141,N_11833);
xor U12216 (N_12216,N_11355,N_10962);
nand U12217 (N_12217,N_10829,N_11039);
and U12218 (N_12218,N_11197,N_11482);
nor U12219 (N_12219,N_11698,N_9779);
or U12220 (N_12220,N_10689,N_10814);
nor U12221 (N_12221,N_9025,N_11308);
nor U12222 (N_12222,N_11602,N_9873);
and U12223 (N_12223,N_10574,N_11500);
nor U12224 (N_12224,N_11749,N_9496);
nand U12225 (N_12225,N_9012,N_9620);
or U12226 (N_12226,N_9870,N_10578);
nand U12227 (N_12227,N_11470,N_11931);
xor U12228 (N_12228,N_9922,N_11016);
xor U12229 (N_12229,N_9529,N_11524);
and U12230 (N_12230,N_11102,N_11462);
xnor U12231 (N_12231,N_10201,N_10806);
nor U12232 (N_12232,N_11598,N_10390);
nor U12233 (N_12233,N_10619,N_11325);
and U12234 (N_12234,N_9443,N_9504);
nand U12235 (N_12235,N_11947,N_9087);
nand U12236 (N_12236,N_9401,N_9286);
and U12237 (N_12237,N_11281,N_9926);
and U12238 (N_12238,N_10900,N_11070);
nor U12239 (N_12239,N_10090,N_9705);
nand U12240 (N_12240,N_9488,N_9818);
nand U12241 (N_12241,N_10868,N_11595);
nor U12242 (N_12242,N_9940,N_9887);
nand U12243 (N_12243,N_11763,N_10631);
and U12244 (N_12244,N_9738,N_11969);
or U12245 (N_12245,N_11189,N_10255);
and U12246 (N_12246,N_9687,N_9517);
and U12247 (N_12247,N_11764,N_11921);
nand U12248 (N_12248,N_11385,N_10892);
nor U12249 (N_12249,N_11159,N_9238);
and U12250 (N_12250,N_11843,N_9949);
nand U12251 (N_12251,N_10636,N_11793);
xnor U12252 (N_12252,N_9930,N_9741);
or U12253 (N_12253,N_9075,N_9599);
nor U12254 (N_12254,N_10664,N_11509);
or U12255 (N_12255,N_9956,N_10592);
xor U12256 (N_12256,N_11444,N_11289);
xor U12257 (N_12257,N_11480,N_9081);
nor U12258 (N_12258,N_9843,N_11922);
or U12259 (N_12259,N_10266,N_11685);
or U12260 (N_12260,N_9703,N_9092);
nor U12261 (N_12261,N_11823,N_9267);
xnor U12262 (N_12262,N_10106,N_10712);
and U12263 (N_12263,N_11748,N_11658);
nor U12264 (N_12264,N_11036,N_11287);
nand U12265 (N_12265,N_9224,N_11090);
and U12266 (N_12266,N_11144,N_9660);
xor U12267 (N_12267,N_10573,N_10880);
nand U12268 (N_12268,N_9724,N_11762);
and U12269 (N_12269,N_10115,N_9036);
and U12270 (N_12270,N_9168,N_11808);
xnor U12271 (N_12271,N_10024,N_10837);
or U12272 (N_12272,N_9938,N_11410);
xor U12273 (N_12273,N_11774,N_10170);
or U12274 (N_12274,N_9607,N_11848);
nor U12275 (N_12275,N_10456,N_10341);
nor U12276 (N_12276,N_9548,N_10004);
nand U12277 (N_12277,N_10663,N_9442);
or U12278 (N_12278,N_11505,N_9114);
or U12279 (N_12279,N_9784,N_10828);
or U12280 (N_12280,N_9258,N_9855);
nand U12281 (N_12281,N_9150,N_9868);
xor U12282 (N_12282,N_9016,N_9491);
nor U12283 (N_12283,N_10104,N_10854);
nand U12284 (N_12284,N_10145,N_9510);
xnor U12285 (N_12285,N_11108,N_11904);
nand U12286 (N_12286,N_9275,N_10789);
nand U12287 (N_12287,N_11557,N_9856);
xor U12288 (N_12288,N_10366,N_11824);
nand U12289 (N_12289,N_10363,N_9946);
and U12290 (N_12290,N_11449,N_11349);
xor U12291 (N_12291,N_10612,N_10957);
or U12292 (N_12292,N_11125,N_11846);
nor U12293 (N_12293,N_10629,N_10705);
or U12294 (N_12294,N_10429,N_10823);
xor U12295 (N_12295,N_10419,N_9994);
xor U12296 (N_12296,N_10083,N_11649);
xor U12297 (N_12297,N_9122,N_11815);
and U12298 (N_12298,N_9381,N_10786);
nor U12299 (N_12299,N_11788,N_11026);
and U12300 (N_12300,N_11925,N_10445);
and U12301 (N_12301,N_10596,N_9702);
xor U12302 (N_12302,N_10565,N_10163);
and U12303 (N_12303,N_11959,N_9828);
xor U12304 (N_12304,N_11639,N_9935);
or U12305 (N_12305,N_11347,N_11621);
and U12306 (N_12306,N_11004,N_9750);
and U12307 (N_12307,N_11501,N_11235);
nor U12308 (N_12308,N_11376,N_10325);
nor U12309 (N_12309,N_10423,N_9158);
nand U12310 (N_12310,N_11663,N_11723);
xnor U12311 (N_12311,N_11854,N_9712);
nand U12312 (N_12312,N_9991,N_10171);
nand U12313 (N_12313,N_10994,N_9296);
nor U12314 (N_12314,N_9597,N_9533);
and U12315 (N_12315,N_10178,N_10515);
and U12316 (N_12316,N_11517,N_10020);
and U12317 (N_12317,N_10800,N_11754);
nand U12318 (N_12318,N_9086,N_9302);
xor U12319 (N_12319,N_11392,N_10760);
nand U12320 (N_12320,N_11628,N_10618);
and U12321 (N_12321,N_10217,N_9112);
nor U12322 (N_12322,N_11897,N_9511);
or U12323 (N_12323,N_11326,N_9766);
or U12324 (N_12324,N_11670,N_10123);
and U12325 (N_12325,N_10649,N_9910);
and U12326 (N_12326,N_9641,N_11709);
xor U12327 (N_12327,N_9869,N_11156);
or U12328 (N_12328,N_9436,N_10062);
or U12329 (N_12329,N_10586,N_9437);
nand U12330 (N_12330,N_9556,N_9090);
or U12331 (N_12331,N_9428,N_11814);
or U12332 (N_12332,N_9625,N_9039);
and U12333 (N_12333,N_9240,N_11536);
or U12334 (N_12334,N_10069,N_11342);
nor U12335 (N_12335,N_10084,N_9056);
nor U12336 (N_12336,N_9986,N_11486);
nand U12337 (N_12337,N_11311,N_11734);
or U12338 (N_12338,N_11543,N_11043);
and U12339 (N_12339,N_10224,N_10678);
or U12340 (N_12340,N_11292,N_10052);
and U12341 (N_12341,N_11072,N_9024);
or U12342 (N_12342,N_9480,N_10448);
or U12343 (N_12343,N_11604,N_11758);
or U12344 (N_12344,N_11080,N_9638);
nand U12345 (N_12345,N_10192,N_11873);
and U12346 (N_12346,N_11790,N_9290);
nand U12347 (N_12347,N_10587,N_11022);
or U12348 (N_12348,N_9723,N_9124);
or U12349 (N_12349,N_11691,N_10857);
xnor U12350 (N_12350,N_11330,N_11850);
nand U12351 (N_12351,N_9777,N_10949);
nor U12352 (N_12352,N_10977,N_9392);
xnor U12353 (N_12353,N_9604,N_10343);
xor U12354 (N_12354,N_11228,N_9404);
nor U12355 (N_12355,N_9084,N_11469);
and U12356 (N_12356,N_9355,N_9816);
xor U12357 (N_12357,N_9219,N_11950);
nor U12358 (N_12358,N_9337,N_10717);
nand U12359 (N_12359,N_10337,N_11320);
nand U12360 (N_12360,N_9927,N_10148);
nand U12361 (N_12361,N_11667,N_11555);
and U12362 (N_12362,N_9004,N_10305);
nor U12363 (N_12363,N_11968,N_9216);
xnor U12364 (N_12364,N_11378,N_9984);
nand U12365 (N_12365,N_10010,N_9654);
and U12366 (N_12366,N_11909,N_9068);
and U12367 (N_12367,N_9570,N_9804);
or U12368 (N_12368,N_10395,N_11485);
or U12369 (N_12369,N_9034,N_10080);
xor U12370 (N_12370,N_9720,N_10641);
nand U12371 (N_12371,N_11994,N_9829);
and U12372 (N_12372,N_10939,N_11393);
and U12373 (N_12373,N_10424,N_11834);
and U12374 (N_12374,N_10036,N_9093);
xnor U12375 (N_12375,N_11066,N_11648);
nor U12376 (N_12376,N_10748,N_9554);
or U12377 (N_12377,N_11541,N_11783);
xor U12378 (N_12378,N_9546,N_11623);
xnor U12379 (N_12379,N_10879,N_10745);
or U12380 (N_12380,N_11059,N_9583);
and U12381 (N_12381,N_10408,N_11088);
nand U12382 (N_12382,N_11479,N_10614);
xor U12383 (N_12383,N_11148,N_9547);
and U12384 (N_12384,N_10909,N_11645);
or U12385 (N_12385,N_9154,N_10500);
xnor U12386 (N_12386,N_9076,N_10184);
nor U12387 (N_12387,N_11138,N_9565);
and U12388 (N_12388,N_11838,N_11406);
and U12389 (N_12389,N_11437,N_10936);
nand U12390 (N_12390,N_10560,N_10477);
nand U12391 (N_12391,N_11902,N_9501);
nor U12392 (N_12392,N_11563,N_10182);
nor U12393 (N_12393,N_11526,N_11991);
nand U12394 (N_12394,N_9650,N_9571);
and U12395 (N_12395,N_10346,N_9291);
nor U12396 (N_12396,N_11394,N_9444);
nor U12397 (N_12397,N_9227,N_10285);
nand U12398 (N_12398,N_10643,N_10489);
xor U12399 (N_12399,N_11341,N_11521);
nand U12400 (N_12400,N_11415,N_11040);
or U12401 (N_12401,N_9080,N_9116);
xnor U12402 (N_12402,N_10945,N_9234);
and U12403 (N_12403,N_9613,N_9462);
nand U12404 (N_12404,N_9193,N_11379);
and U12405 (N_12405,N_11130,N_9202);
nand U12406 (N_12406,N_9165,N_10405);
nor U12407 (N_12407,N_11243,N_11008);
nand U12408 (N_12408,N_11666,N_9103);
xor U12409 (N_12409,N_10469,N_10431);
and U12410 (N_12410,N_10535,N_10878);
nand U12411 (N_12411,N_9178,N_10864);
nor U12412 (N_12412,N_10453,N_10685);
and U12413 (N_12413,N_9110,N_10263);
or U12414 (N_12414,N_9775,N_9808);
or U12415 (N_12415,N_9611,N_11886);
or U12416 (N_12416,N_11452,N_10211);
xor U12417 (N_12417,N_9026,N_10917);
nand U12418 (N_12418,N_11887,N_9314);
nand U12419 (N_12419,N_10954,N_11735);
or U12420 (N_12420,N_11791,N_11369);
nor U12421 (N_12421,N_11938,N_10849);
nand U12422 (N_12422,N_11928,N_11242);
xor U12423 (N_12423,N_9431,N_9710);
nand U12424 (N_12424,N_11515,N_11007);
and U12425 (N_12425,N_10093,N_11837);
xnor U12426 (N_12426,N_11616,N_9615);
nor U12427 (N_12427,N_10282,N_10344);
xor U12428 (N_12428,N_9865,N_11153);
xor U12429 (N_12429,N_11117,N_10229);
or U12430 (N_12430,N_10764,N_10033);
xor U12431 (N_12431,N_9769,N_9478);
or U12432 (N_12432,N_10463,N_11166);
xor U12433 (N_12433,N_11953,N_9361);
nand U12434 (N_12434,N_11052,N_10841);
nor U12435 (N_12435,N_11597,N_11785);
nor U12436 (N_12436,N_11971,N_11588);
nor U12437 (N_12437,N_9281,N_10604);
or U12438 (N_12438,N_11826,N_10236);
xor U12439 (N_12439,N_10076,N_10625);
xor U12440 (N_12440,N_11746,N_10738);
nand U12441 (N_12441,N_10374,N_10151);
or U12442 (N_12442,N_10877,N_11528);
xnor U12443 (N_12443,N_9805,N_9327);
or U12444 (N_12444,N_9396,N_9883);
or U12445 (N_12445,N_10329,N_9268);
and U12446 (N_12446,N_9999,N_9495);
and U12447 (N_12447,N_11020,N_11316);
nor U12448 (N_12448,N_10623,N_9574);
nand U12449 (N_12449,N_9798,N_11372);
or U12450 (N_12450,N_11865,N_10651);
and U12451 (N_12451,N_9526,N_10003);
nand U12452 (N_12452,N_9049,N_9616);
xnor U12453 (N_12453,N_10822,N_11046);
nand U12454 (N_12454,N_9706,N_9096);
nand U12455 (N_12455,N_10752,N_11299);
nand U12456 (N_12456,N_11019,N_11425);
nor U12457 (N_12457,N_11992,N_11803);
nand U12458 (N_12458,N_10064,N_11487);
and U12459 (N_12459,N_9484,N_11481);
or U12460 (N_12460,N_11589,N_10207);
nand U12461 (N_12461,N_9692,N_10259);
nand U12462 (N_12462,N_9347,N_9191);
xor U12463 (N_12463,N_10681,N_10985);
or U12464 (N_12464,N_10703,N_10567);
nand U12465 (N_12465,N_10095,N_10555);
xnor U12466 (N_12466,N_10049,N_11946);
nor U12467 (N_12467,N_11728,N_10594);
xnor U12468 (N_12468,N_11490,N_11942);
and U12469 (N_12469,N_9508,N_11781);
xnor U12470 (N_12470,N_11306,N_9871);
or U12471 (N_12471,N_10858,N_10233);
and U12472 (N_12472,N_10920,N_10218);
or U12473 (N_12473,N_9260,N_9783);
and U12474 (N_12474,N_9146,N_11307);
nor U12475 (N_12475,N_10042,N_9297);
nor U12476 (N_12476,N_10813,N_11493);
nor U12477 (N_12477,N_11223,N_11813);
nor U12478 (N_12478,N_11352,N_10368);
and U12479 (N_12479,N_10726,N_9681);
nor U12480 (N_12480,N_10381,N_11572);
nor U12481 (N_12481,N_9731,N_9341);
or U12482 (N_12482,N_9422,N_11353);
nand U12483 (N_12483,N_9091,N_9410);
nand U12484 (N_12484,N_11309,N_11086);
nor U12485 (N_12485,N_11558,N_9312);
or U12486 (N_12486,N_9476,N_10127);
or U12487 (N_12487,N_9860,N_10622);
nand U12488 (N_12488,N_11494,N_11067);
or U12489 (N_12489,N_9666,N_9042);
and U12490 (N_12490,N_9918,N_9787);
and U12491 (N_12491,N_10970,N_11498);
or U12492 (N_12492,N_9498,N_10465);
nor U12493 (N_12493,N_9557,N_9005);
nor U12494 (N_12494,N_11799,N_9921);
or U12495 (N_12495,N_11979,N_9876);
or U12496 (N_12496,N_11657,N_10281);
xor U12497 (N_12497,N_10509,N_10125);
or U12498 (N_12498,N_10369,N_11018);
nand U12499 (N_12499,N_9159,N_11703);
or U12500 (N_12500,N_10895,N_11849);
nand U12501 (N_12501,N_11706,N_11560);
nor U12502 (N_12502,N_11996,N_9197);
and U12503 (N_12503,N_10768,N_11583);
nand U12504 (N_12504,N_9100,N_10723);
xnor U12505 (N_12505,N_11948,N_9864);
xor U12506 (N_12506,N_9867,N_11032);
or U12507 (N_12507,N_10569,N_10162);
and U12508 (N_12508,N_10128,N_10284);
nor U12509 (N_12509,N_11041,N_10244);
nand U12510 (N_12510,N_10584,N_11284);
nand U12511 (N_12511,N_11298,N_10334);
xnor U12512 (N_12512,N_9634,N_10150);
and U12513 (N_12513,N_11472,N_11105);
nor U12514 (N_12514,N_11154,N_11276);
or U12515 (N_12515,N_10863,N_9053);
and U12516 (N_12516,N_10149,N_11795);
or U12517 (N_12517,N_11017,N_10615);
nor U12518 (N_12518,N_9925,N_11419);
nor U12519 (N_12519,N_11403,N_11977);
xor U12520 (N_12520,N_10546,N_9576);
and U12521 (N_12521,N_11891,N_11704);
xnor U12522 (N_12522,N_10332,N_11389);
nor U12523 (N_12523,N_11794,N_10897);
xnor U12524 (N_12524,N_10749,N_10517);
xor U12525 (N_12525,N_10247,N_10021);
and U12526 (N_12526,N_9543,N_10120);
nor U12527 (N_12527,N_11056,N_11802);
nand U12528 (N_12528,N_11556,N_9559);
nor U12529 (N_12529,N_9521,N_11157);
or U12530 (N_12530,N_10338,N_11967);
xor U12531 (N_12531,N_10959,N_9806);
nand U12532 (N_12532,N_9104,N_10261);
nand U12533 (N_12533,N_10231,N_11391);
nor U12534 (N_12534,N_11441,N_10802);
nand U12535 (N_12535,N_9535,N_10547);
nor U12536 (N_12536,N_9896,N_9195);
nor U12537 (N_12537,N_10039,N_11054);
and U12538 (N_12538,N_9023,N_11042);
nor U12539 (N_12539,N_9943,N_9249);
or U12540 (N_12540,N_9653,N_9763);
xor U12541 (N_12541,N_11321,N_10327);
nand U12542 (N_12542,N_9215,N_10657);
and U12543 (N_12543,N_10794,N_11477);
nor U12544 (N_12544,N_10725,N_10695);
and U12545 (N_12545,N_10195,N_11917);
or U12546 (N_12546,N_11442,N_10873);
or U12547 (N_12547,N_11941,N_9420);
and U12548 (N_12548,N_10750,N_10536);
or U12549 (N_12549,N_9744,N_9751);
nand U12550 (N_12550,N_9539,N_11617);
nand U12551 (N_12551,N_10600,N_9239);
nor U12552 (N_12552,N_10874,N_9610);
xor U12553 (N_12553,N_11131,N_10524);
nand U12554 (N_12554,N_10172,N_11798);
or U12555 (N_12555,N_11809,N_11546);
xnor U12556 (N_12556,N_9265,N_9952);
or U12557 (N_12557,N_10809,N_11570);
or U12558 (N_12558,N_11057,N_11951);
xor U12559 (N_12559,N_9608,N_11751);
nor U12560 (N_12560,N_10693,N_10006);
or U12561 (N_12561,N_10117,N_11926);
xnor U12562 (N_12562,N_10413,N_11147);
or U12563 (N_12563,N_11377,N_10354);
xnor U12564 (N_12564,N_9780,N_9362);
or U12565 (N_12565,N_11128,N_10444);
and U12566 (N_12566,N_11789,N_9951);
nand U12567 (N_12567,N_10262,N_9376);
nor U12568 (N_12568,N_9408,N_11434);
or U12569 (N_12569,N_9329,N_10215);
and U12570 (N_12570,N_9183,N_9664);
nor U12571 (N_12571,N_11340,N_9252);
or U12572 (N_12572,N_10851,N_10188);
and U12573 (N_12573,N_9380,N_11635);
nand U12574 (N_12574,N_11601,N_11380);
nand U12575 (N_12575,N_9276,N_9909);
and U12576 (N_12576,N_10887,N_11423);
nor U12577 (N_12577,N_11359,N_10050);
nand U12578 (N_12578,N_11835,N_10189);
or U12579 (N_12579,N_11302,N_9575);
nand U12580 (N_12580,N_9003,N_11264);
or U12581 (N_12581,N_10501,N_10875);
or U12582 (N_12582,N_9455,N_10060);
and U12583 (N_12583,N_9134,N_10447);
or U12584 (N_12584,N_9044,N_11842);
nand U12585 (N_12585,N_11218,N_11337);
xor U12586 (N_12586,N_11464,N_11025);
nor U12587 (N_12587,N_10350,N_9827);
or U12588 (N_12588,N_11678,N_9701);
nand U12589 (N_12589,N_10267,N_10937);
nand U12590 (N_12590,N_9969,N_11676);
and U12591 (N_12591,N_9507,N_9482);
xnor U12592 (N_12592,N_11246,N_11876);
xnor U12593 (N_12593,N_11508,N_9229);
nand U12594 (N_12594,N_11107,N_10730);
nor U12595 (N_12595,N_9088,N_9519);
xor U12596 (N_12596,N_9960,N_11445);
nand U12597 (N_12597,N_10915,N_10777);
or U12598 (N_12598,N_11945,N_9992);
nor U12599 (N_12599,N_10180,N_10185);
xnor U12600 (N_12600,N_10562,N_10059);
nand U12601 (N_12601,N_9107,N_9579);
nand U12602 (N_12602,N_9851,N_10411);
nand U12603 (N_12603,N_11466,N_9481);
or U12604 (N_12604,N_9722,N_9133);
and U12605 (N_12605,N_9452,N_9532);
xor U12606 (N_12606,N_9820,N_10784);
nor U12607 (N_12607,N_10778,N_10544);
nand U12608 (N_12608,N_9493,N_9354);
xor U12609 (N_12609,N_9727,N_11855);
and U12610 (N_12610,N_10015,N_11222);
nor U12611 (N_12611,N_9126,N_10948);
or U12612 (N_12612,N_9261,N_9947);
or U12613 (N_12613,N_10545,N_9069);
xor U12614 (N_12614,N_9862,N_9578);
and U12615 (N_12615,N_9899,N_10113);
nor U12616 (N_12616,N_10884,N_11383);
xnor U12617 (N_12617,N_10306,N_10335);
or U12618 (N_12618,N_11861,N_10303);
nor U12619 (N_12619,N_9220,N_11332);
or U12620 (N_12620,N_10640,N_11741);
nor U12621 (N_12621,N_10362,N_9352);
xnor U12622 (N_12622,N_9523,N_9402);
or U12623 (N_12623,N_10602,N_11712);
nand U12624 (N_12624,N_11634,N_9944);
nor U12625 (N_12625,N_9509,N_11960);
nand U12626 (N_12626,N_9788,N_11995);
or U12627 (N_12627,N_10935,N_10109);
xor U12628 (N_12628,N_10057,N_11804);
and U12629 (N_12629,N_9879,N_10513);
and U12630 (N_12630,N_10645,N_10668);
or U12631 (N_12631,N_11878,N_9319);
nand U12632 (N_12632,N_11158,N_10838);
nand U12633 (N_12633,N_11126,N_9754);
nor U12634 (N_12634,N_11721,N_11447);
nand U12635 (N_12635,N_9923,N_11273);
xnor U12636 (N_12636,N_10982,N_9413);
and U12637 (N_12637,N_10451,N_11174);
and U12638 (N_12638,N_10037,N_10773);
and U12639 (N_12639,N_10143,N_9163);
xnor U12640 (N_12640,N_9933,N_9320);
or U12641 (N_12641,N_11852,N_11474);
or U12642 (N_12642,N_9662,N_11784);
nand U12643 (N_12643,N_11143,N_9283);
xor U12644 (N_12644,N_11932,N_10609);
xnor U12645 (N_12645,N_9015,N_11753);
and U12646 (N_12646,N_9440,N_11518);
or U12647 (N_12647,N_10910,N_11587);
nor U12648 (N_12648,N_9941,N_9348);
or U12649 (N_12649,N_11354,N_11491);
nor U12650 (N_12650,N_9156,N_9631);
and U12651 (N_12651,N_11511,N_11576);
or U12652 (N_12652,N_11478,N_10311);
nand U12653 (N_12653,N_10379,N_9322);
nand U12654 (N_12654,N_9236,N_11831);
and U12655 (N_12655,N_10091,N_10296);
or U12656 (N_12656,N_10349,N_11115);
or U12657 (N_12657,N_10564,N_11607);
nor U12658 (N_12658,N_9198,N_10250);
nand U12659 (N_12659,N_11458,N_11976);
and U12660 (N_12660,N_10089,N_11532);
or U12661 (N_12661,N_9190,N_9400);
or U12662 (N_12662,N_9045,N_11079);
nor U12663 (N_12663,N_10087,N_11329);
nor U12664 (N_12664,N_10914,N_10376);
and U12665 (N_12665,N_9222,N_10494);
xnor U12666 (N_12666,N_10532,N_9293);
nand U12667 (N_12667,N_9520,N_9633);
xnor U12668 (N_12668,N_11053,N_10265);
or U12669 (N_12669,N_9453,N_9471);
and U12670 (N_12670,N_11810,N_9911);
nor U12671 (N_12671,N_10464,N_11725);
nand U12672 (N_12672,N_10186,N_10805);
nor U12673 (N_12673,N_10426,N_11457);
xnor U12674 (N_12674,N_9915,N_9101);
xor U12675 (N_12675,N_9752,N_9274);
or U12676 (N_12676,N_9046,N_10633);
nand U12677 (N_12677,N_11000,N_9733);
xnor U12678 (N_12678,N_11611,N_10399);
and U12679 (N_12679,N_9914,N_11270);
nand U12680 (N_12680,N_10323,N_10028);
xor U12681 (N_12681,N_11609,N_10029);
nand U12682 (N_12682,N_11718,N_11999);
and U12683 (N_12683,N_10415,N_9530);
and U12684 (N_12684,N_9793,N_10230);
nand U12685 (N_12685,N_11729,N_10941);
xnor U12686 (N_12686,N_9665,N_10551);
nor U12687 (N_12687,N_9671,N_10659);
and U12688 (N_12688,N_11819,N_9050);
nor U12689 (N_12689,N_9438,N_11319);
nor U12690 (N_12690,N_9067,N_10710);
or U12691 (N_12691,N_9983,N_11937);
or U12692 (N_12692,N_10315,N_11534);
nor U12693 (N_12693,N_10035,N_10347);
nand U12694 (N_12694,N_10078,N_10943);
xnor U12695 (N_12695,N_11343,N_11836);
and U12696 (N_12696,N_11600,N_9587);
nor U12697 (N_12697,N_10321,N_9340);
xnor U12698 (N_12698,N_9284,N_11082);
and U12699 (N_12699,N_9995,N_9187);
or U12700 (N_12700,N_9257,N_10624);
nand U12701 (N_12701,N_10022,N_10412);
xnor U12702 (N_12702,N_9957,N_9889);
nor U12703 (N_12703,N_9230,N_9730);
or U12704 (N_12704,N_9672,N_9586);
xnor U12705 (N_12705,N_11450,N_10208);
and U12706 (N_12706,N_9866,N_10421);
and U12707 (N_12707,N_10055,N_11448);
xnor U12708 (N_12708,N_11012,N_11127);
and U12709 (N_12709,N_10528,N_9346);
nand U12710 (N_12710,N_9477,N_11654);
nor U12711 (N_12711,N_10721,N_10098);
or U12712 (N_12712,N_9683,N_9656);
and U12713 (N_12713,N_9809,N_9996);
and U12714 (N_12714,N_11756,N_9398);
and U12715 (N_12715,N_10804,N_10196);
xnor U12716 (N_12716,N_11339,N_11068);
xor U12717 (N_12717,N_11720,N_9430);
or U12718 (N_12718,N_10183,N_10508);
xor U12719 (N_12719,N_9552,N_11869);
nand U12720 (N_12720,N_10377,N_11596);
or U12721 (N_12721,N_11345,N_11282);
nand U12722 (N_12722,N_10396,N_11285);
nor U12723 (N_12723,N_11592,N_10482);
xnor U12724 (N_12724,N_9231,N_9786);
or U12725 (N_12725,N_10967,N_9164);
or U12726 (N_12726,N_10351,N_10073);
and U12727 (N_12727,N_11460,N_10918);
nand U12728 (N_12728,N_9309,N_10342);
and U12729 (N_12729,N_10040,N_11564);
nand U12730 (N_12730,N_9255,N_11252);
nor U12731 (N_12731,N_11662,N_11759);
nor U12732 (N_12732,N_9512,N_9256);
nand U12733 (N_12733,N_10041,N_9278);
or U12734 (N_12734,N_10092,N_9266);
and U12735 (N_12735,N_10237,N_9262);
and U12736 (N_12736,N_11188,N_10216);
nand U12737 (N_12737,N_9800,N_11334);
nand U12738 (N_12738,N_10203,N_11796);
or U12739 (N_12739,N_11256,N_10817);
or U12740 (N_12740,N_11028,N_11913);
nor U12741 (N_12741,N_9878,N_10736);
and U12742 (N_12742,N_9636,N_9768);
and U12743 (N_12743,N_11851,N_11280);
xnor U12744 (N_12744,N_11743,N_9131);
nor U12745 (N_12745,N_11619,N_10654);
and U12746 (N_12746,N_10070,N_10591);
xor U12747 (N_12747,N_11880,N_9663);
nor U12748 (N_12748,N_9417,N_9845);
or U12749 (N_12749,N_11050,N_11559);
nor U12750 (N_12750,N_9835,N_10922);
or U12751 (N_12751,N_10027,N_10766);
xor U12752 (N_12752,N_10254,N_11752);
nand U12753 (N_12753,N_10475,N_9399);
nand U12754 (N_12754,N_10480,N_10974);
and U12755 (N_12755,N_11360,N_10164);
xnor U12756 (N_12756,N_10088,N_11424);
nand U12757 (N_12757,N_11297,N_9799);
and U12758 (N_12758,N_9043,N_9059);
or U12759 (N_12759,N_9217,N_9253);
nor U12760 (N_12760,N_10507,N_9308);
nand U12761 (N_12761,N_9945,N_10848);
nor U12762 (N_12762,N_10110,N_11045);
nor U12763 (N_12763,N_11730,N_10316);
or U12764 (N_12764,N_9235,N_11908);
and U12765 (N_12765,N_9429,N_10638);
nand U12766 (N_12766,N_9064,N_10902);
and U12767 (N_12767,N_10755,N_9228);
xor U12768 (N_12768,N_9982,N_9670);
nand U12769 (N_12769,N_9588,N_10384);
or U12770 (N_12770,N_9288,N_11397);
nand U12771 (N_12771,N_10563,N_10598);
or U12772 (N_12772,N_9817,N_10238);
or U12773 (N_12773,N_9898,N_10995);
xor U12774 (N_12774,N_11318,N_11333);
and U12775 (N_12775,N_11119,N_10597);
nor U12776 (N_12776,N_11467,N_9221);
and U12777 (N_12777,N_9668,N_10012);
nand U12778 (N_12778,N_11641,N_11097);
or U12779 (N_12779,N_11627,N_9916);
nor U12780 (N_12780,N_11738,N_9859);
xor U12781 (N_12781,N_10468,N_10611);
nand U12782 (N_12782,N_9465,N_9247);
and U12783 (N_12783,N_9407,N_10781);
and U12784 (N_12784,N_9875,N_9830);
and U12785 (N_12785,N_9877,N_10543);
and U12786 (N_12786,N_10711,N_9179);
nand U12787 (N_12787,N_9387,N_11906);
or U12788 (N_12788,N_11367,N_9138);
nor U12789 (N_12789,N_9203,N_11268);
nand U12790 (N_12790,N_10242,N_10138);
or U12791 (N_12791,N_10418,N_10014);
xnor U12792 (N_12792,N_10253,N_10132);
xnor U12793 (N_12793,N_11900,N_11061);
nor U12794 (N_12794,N_11181,N_10385);
nand U12795 (N_12795,N_9035,N_9433);
nand U12796 (N_12796,N_9882,N_9963);
or U12797 (N_12797,N_9826,N_9833);
nand U12798 (N_12798,N_9589,N_9885);
or U12799 (N_12799,N_11121,N_11315);
xnor U12800 (N_12800,N_10699,N_10166);
nor U12801 (N_12801,N_10514,N_11520);
nor U12802 (N_12802,N_10688,N_10796);
xor U12803 (N_12803,N_10984,N_10860);
xor U12804 (N_12804,N_10713,N_11912);
or U12805 (N_12805,N_10360,N_9305);
or U12806 (N_12806,N_9280,N_10769);
nor U12807 (N_12807,N_11582,N_9772);
and U12808 (N_12808,N_9767,N_11120);
and U12809 (N_12809,N_9373,N_10280);
or U12810 (N_12810,N_10007,N_11573);
nor U12811 (N_12811,N_9758,N_10772);
nor U12812 (N_12812,N_10759,N_11845);
and U12813 (N_12813,N_11533,N_11911);
xnor U12814 (N_12814,N_11407,N_9207);
nand U12815 (N_12815,N_9310,N_9895);
xnor U12816 (N_12816,N_10023,N_11267);
and U12817 (N_12817,N_9263,N_10270);
and U12818 (N_12818,N_10276,N_11551);
and U12819 (N_12819,N_9472,N_9359);
and U12820 (N_12820,N_10529,N_10718);
and U12821 (N_12821,N_11684,N_11422);
nand U12822 (N_12822,N_11727,N_11331);
nor U12823 (N_12823,N_10548,N_9564);
and U12824 (N_12824,N_11440,N_9646);
nor U12825 (N_12825,N_10790,N_9591);
xnor U12826 (N_12826,N_11629,N_10130);
nor U12827 (N_12827,N_11212,N_10333);
or U12828 (N_12828,N_11633,N_10916);
nor U12829 (N_12829,N_9492,N_11140);
and U12830 (N_12830,N_9890,N_11650);
xnor U12831 (N_12831,N_10856,N_9961);
or U12832 (N_12832,N_10286,N_11214);
or U12833 (N_12833,N_10331,N_10951);
nor U12834 (N_12834,N_11443,N_9457);
xnor U12835 (N_12835,N_9913,N_11112);
nand U12836 (N_12836,N_10669,N_9432);
nor U12837 (N_12837,N_10258,N_10503);
nor U12838 (N_12838,N_11655,N_11821);
nand U12839 (N_12839,N_11361,N_10339);
nor U12840 (N_12840,N_11972,N_11982);
and U12841 (N_12841,N_9350,N_9785);
or U12842 (N_12842,N_11111,N_10973);
nor U12843 (N_12843,N_11686,N_9762);
nor U12844 (N_12844,N_10605,N_10199);
and U12845 (N_12845,N_10133,N_9051);
nand U12846 (N_12846,N_10797,N_10398);
nor U12847 (N_12847,N_9609,N_11071);
nand U12848 (N_12848,N_9749,N_11944);
or U12849 (N_12849,N_9796,N_10159);
and U12850 (N_12850,N_11744,N_10317);
and U12851 (N_12851,N_11073,N_11896);
nand U12852 (N_12852,N_10742,N_11918);
xor U12853 (N_12853,N_11839,N_11514);
or U12854 (N_12854,N_10788,N_11980);
and U12855 (N_12855,N_9259,N_9694);
and U12856 (N_12856,N_9967,N_9836);
and U12857 (N_12857,N_10330,N_9757);
or U12858 (N_12858,N_10679,N_11237);
nor U12859 (N_12859,N_9595,N_11145);
or U12860 (N_12860,N_11489,N_9939);
nand U12861 (N_12861,N_10047,N_9729);
and U12862 (N_12862,N_11697,N_11062);
or U12863 (N_12863,N_10993,N_10139);
nor U12864 (N_12864,N_10370,N_10239);
nand U12865 (N_12865,N_11660,N_9153);
nor U12866 (N_12866,N_9739,N_9892);
nor U12867 (N_12867,N_11395,N_11513);
or U12868 (N_12868,N_11335,N_11782);
or U12869 (N_12869,N_9270,N_9585);
and U12870 (N_12870,N_11411,N_10144);
nor U12871 (N_12871,N_10326,N_11231);
and U12872 (N_12872,N_11209,N_11668);
and U12873 (N_12873,N_11384,N_9989);
nor U12874 (N_12874,N_9166,N_11605);
and U12875 (N_12875,N_10313,N_11885);
and U12876 (N_12876,N_11428,N_10245);
nand U12877 (N_12877,N_9074,N_10100);
nand U12878 (N_12878,N_11984,N_11544);
nor U12879 (N_12879,N_11087,N_11303);
nand U12880 (N_12880,N_9171,N_9489);
nor U12881 (N_12881,N_9700,N_11625);
or U12882 (N_12882,N_11225,N_9132);
nor U12883 (N_12883,N_9287,N_9954);
and U12884 (N_12884,N_9774,N_10540);
nand U12885 (N_12885,N_10126,N_11135);
nor U12886 (N_12886,N_11747,N_9172);
nor U12887 (N_12887,N_9105,N_10599);
or U12888 (N_12888,N_9013,N_10032);
nor U12889 (N_12889,N_11998,N_10637);
and U12890 (N_12890,N_10205,N_9977);
nor U12891 (N_12891,N_11172,N_10289);
nor U12892 (N_12892,N_11988,N_10428);
xnor U12893 (N_12893,N_11881,N_10066);
nor U12894 (N_12894,N_10906,N_10810);
and U12895 (N_12895,N_11857,N_10223);
or U12896 (N_12896,N_11232,N_11562);
nor U12897 (N_12897,N_10048,N_11175);
xnor U12898 (N_12898,N_11049,N_9970);
and U12899 (N_12899,N_10470,N_11682);
nor U12900 (N_12900,N_9605,N_11832);
or U12901 (N_12901,N_10771,N_9151);
xnor U12902 (N_12902,N_10065,N_10735);
or U12903 (N_12903,N_10158,N_10527);
xor U12904 (N_12904,N_10248,N_10077);
xor U12905 (N_12905,N_11327,N_10844);
or U12906 (N_12906,N_10671,N_9567);
xor U12907 (N_12907,N_11060,N_11768);
or U12908 (N_12908,N_9130,N_9789);
or U12909 (N_12909,N_9953,N_10852);
nand U12910 (N_12910,N_11997,N_11671);
nand U12911 (N_12911,N_11417,N_10607);
nand U12912 (N_12912,N_11750,N_10593);
and U12913 (N_12913,N_9325,N_11568);
xor U12914 (N_12914,N_9412,N_9734);
nor U12915 (N_12915,N_9411,N_10492);
or U12916 (N_12916,N_9838,N_9063);
nor U12917 (N_12917,N_10134,N_11317);
xor U12918 (N_12918,N_10521,N_9691);
or U12919 (N_12919,N_10256,N_9379);
or U12920 (N_12920,N_10799,N_9169);
or U12921 (N_12921,N_10785,N_9306);
or U12922 (N_12922,N_10310,N_9174);
nand U12923 (N_12923,N_10274,N_9823);
or U12924 (N_12924,N_9186,N_9177);
xnor U12925 (N_12925,N_10926,N_11830);
nand U12926 (N_12926,N_9537,N_10461);
nor U12927 (N_12927,N_11031,N_10850);
or U12928 (N_12928,N_11940,N_11626);
nor U12929 (N_12929,N_10260,N_11152);
xor U12930 (N_12930,N_11910,N_10018);
xnor U12931 (N_12931,N_9667,N_10571);
and U12932 (N_12932,N_9601,N_9368);
nor U12933 (N_12933,N_10998,N_9726);
nand U12934 (N_12934,N_9695,N_9569);
nor U12935 (N_12935,N_11171,N_9743);
nand U12936 (N_12936,N_10232,N_9446);
or U12937 (N_12937,N_9041,N_11015);
and U12938 (N_12938,N_11757,N_9563);
xor U12939 (N_12939,N_9245,N_9697);
and U12940 (N_12940,N_11047,N_9459);
nor U12941 (N_12941,N_9137,N_9406);
nor U12942 (N_12942,N_9502,N_9030);
and U12943 (N_12943,N_9937,N_9600);
or U12944 (N_12944,N_9684,N_11943);
xor U12945 (N_12945,N_10886,N_11905);
nor U12946 (N_12946,N_10378,N_11807);
nand U12947 (N_12947,N_11301,N_11920);
and U12948 (N_12948,N_9167,N_10556);
and U12949 (N_12949,N_11859,N_11978);
xnor U12950 (N_12950,N_10840,N_11162);
or U12951 (N_12951,N_11190,N_9066);
nor U12952 (N_12952,N_9175,N_11901);
and U12953 (N_12953,N_9515,N_11574);
nor U12954 (N_12954,N_11898,N_9301);
and U12955 (N_12955,N_11571,N_9920);
or U12956 (N_12956,N_11400,N_9531);
or U12957 (N_12957,N_11436,N_11713);
xnor U12958 (N_12958,N_11471,N_11114);
nand U12959 (N_12959,N_11989,N_9541);
or U12960 (N_12960,N_9657,N_11257);
and U12961 (N_12961,N_10099,N_10958);
or U12962 (N_12962,N_10774,N_9842);
nand U12963 (N_12963,N_9707,N_11064);
or U12964 (N_12964,N_10881,N_11646);
and U12965 (N_12965,N_10808,N_11324);
nor U12966 (N_12966,N_11224,N_11266);
nor U12967 (N_12967,N_10670,N_11346);
or U12968 (N_12968,N_10783,N_10298);
nand U12969 (N_12969,N_10662,N_11503);
or U12970 (N_12970,N_10652,N_9072);
xnor U12971 (N_12971,N_11594,N_9832);
and U12972 (N_12972,N_9881,N_11304);
or U12973 (N_12973,N_11132,N_10459);
and U12974 (N_12974,N_9651,N_10336);
or U12975 (N_12975,N_10716,N_10557);
nand U12976 (N_12976,N_9077,N_9528);
and U12977 (N_12977,N_11055,N_10432);
xnor U12978 (N_12978,N_11693,N_10191);
and U12979 (N_12979,N_9313,N_10845);
nand U12980 (N_12980,N_9111,N_11461);
xnor U12981 (N_12981,N_11726,N_9997);
xor U12982 (N_12982,N_9581,N_11044);
and U12983 (N_12983,N_9002,N_10294);
nand U12984 (N_12984,N_10085,N_10666);
nand U12985 (N_12985,N_9900,N_10673);
nand U12986 (N_12986,N_11766,N_9776);
nand U12987 (N_12987,N_10987,N_11078);
nor U12988 (N_12988,N_11561,N_10744);
and U12989 (N_12989,N_10442,N_10680);
nand U12990 (N_12990,N_10187,N_9972);
nand U12991 (N_12991,N_11234,N_11170);
nor U12992 (N_12992,N_11553,N_11249);
xor U12993 (N_12993,N_10210,N_10096);
or U12994 (N_12994,N_10102,N_10357);
nand U12995 (N_12995,N_11512,N_11468);
xnor U12996 (N_12996,N_11779,N_11357);
nand U12997 (N_12997,N_9513,N_11692);
nor U12998 (N_12998,N_10946,N_11261);
xnor U12999 (N_12999,N_9136,N_9421);
nand U13000 (N_13000,N_9333,N_9000);
and U13001 (N_13001,N_9929,N_9185);
or U13002 (N_13002,N_9065,N_9419);
xor U13003 (N_13003,N_9680,N_10122);
or U13004 (N_13004,N_11603,N_10616);
and U13005 (N_13005,N_10644,N_10016);
nor U13006 (N_13006,N_9623,N_10054);
nand U13007 (N_13007,N_10934,N_11116);
nor U13008 (N_13008,N_9464,N_9397);
and U13009 (N_13009,N_11702,N_10388);
and U13010 (N_13010,N_11104,N_11983);
nand U13011 (N_13011,N_11204,N_9073);
nand U13012 (N_13012,N_9908,N_11862);
nor U13013 (N_13013,N_9682,N_9242);
nor U13014 (N_13014,N_11435,N_10190);
or U13015 (N_13015,N_10996,N_9184);
nand U13016 (N_13016,N_9206,N_10621);
xor U13017 (N_13017,N_11638,N_9149);
nor U13018 (N_13018,N_10433,N_11083);
xor U13019 (N_13019,N_10561,N_9467);
xor U13020 (N_13020,N_11206,N_11291);
nand U13021 (N_13021,N_9677,N_9577);
xor U13022 (N_13022,N_9626,N_11806);
and U13023 (N_13023,N_10476,N_10533);
and U13024 (N_13024,N_9208,N_10861);
xnor U13025 (N_13025,N_11636,N_11939);
or U13026 (N_13026,N_10320,N_9522);
nor U13027 (N_13027,N_11184,N_9316);
or U13028 (N_13028,N_9182,N_9218);
or U13029 (N_13029,N_10882,N_10613);
and U13030 (N_13030,N_11263,N_9998);
nand U13031 (N_13031,N_11923,N_9802);
nand U13032 (N_13032,N_9055,N_11099);
or U13033 (N_13033,N_9709,N_10862);
and U13034 (N_13034,N_9029,N_9098);
nand U13035 (N_13035,N_9017,N_9358);
nand U13036 (N_13036,N_10972,N_10103);
xnor U13037 (N_13037,N_11081,N_9047);
or U13038 (N_13038,N_11539,N_9389);
xor U13039 (N_13039,N_11314,N_9525);
nand U13040 (N_13040,N_9790,N_10739);
nor U13041 (N_13041,N_11787,N_11777);
or U13042 (N_13042,N_11390,N_11567);
nor U13043 (N_13043,N_11465,N_9196);
nand U13044 (N_13044,N_9344,N_10307);
and U13045 (N_13045,N_10153,N_10460);
nor U13046 (N_13046,N_10462,N_11687);
and U13047 (N_13047,N_9819,N_9756);
or U13048 (N_13048,N_11123,N_10403);
xnor U13049 (N_13049,N_10932,N_9416);
nand U13050 (N_13050,N_9959,N_11523);
nor U13051 (N_13051,N_9771,N_11161);
nand U13052 (N_13052,N_11954,N_10765);
or U13053 (N_13053,N_11103,N_9814);
nor U13054 (N_13054,N_10290,N_10173);
or U13055 (N_13055,N_11037,N_11196);
nand U13056 (N_13056,N_11262,N_9622);
xnor U13057 (N_13057,N_11182,N_11178);
nor U13058 (N_13058,N_10391,N_10991);
xor U13059 (N_13059,N_11179,N_9628);
and U13060 (N_13060,N_10583,N_10493);
nor U13061 (N_13061,N_10795,N_11193);
nand U13062 (N_13062,N_11164,N_9696);
and U13063 (N_13063,N_10179,N_10275);
nand U13064 (N_13064,N_11191,N_11011);
or U13065 (N_13065,N_9181,N_9886);
nor U13066 (N_13066,N_9872,N_9233);
and U13067 (N_13067,N_11272,N_11871);
xnor U13068 (N_13068,N_10889,N_9277);
nand U13069 (N_13069,N_9629,N_11879);
nand U13070 (N_13070,N_9962,N_11005);
nand U13071 (N_13071,N_10743,N_10504);
and U13072 (N_13072,N_9254,N_10497);
nor U13073 (N_13073,N_9617,N_11409);
nor U13074 (N_13074,N_10271,N_10116);
or U13075 (N_13075,N_10505,N_11554);
xor U13076 (N_13076,N_10981,N_10762);
or U13077 (N_13077,N_11507,N_10520);
xor U13078 (N_13078,N_9394,N_11412);
nor U13079 (N_13079,N_10140,N_9861);
xnor U13080 (N_13080,N_11771,N_9160);
nand U13081 (N_13081,N_11914,N_11840);
nor U13082 (N_13082,N_11405,N_11322);
and U13083 (N_13083,N_11336,N_11381);
xnor U13084 (N_13084,N_10776,N_9441);
or U13085 (N_13085,N_10839,N_11294);
or U13086 (N_13086,N_11714,N_11344);
nand U13087 (N_13087,N_9649,N_11872);
nand U13088 (N_13088,N_10340,N_10213);
and U13089 (N_13089,N_11021,N_10479);
and U13090 (N_13090,N_11430,N_9848);
nor U13091 (N_13091,N_9614,N_9147);
xnor U13092 (N_13092,N_9966,N_10754);
nand U13093 (N_13093,N_10157,N_11708);
or U13094 (N_13094,N_10372,N_9466);
nor U13095 (N_13095,N_9463,N_9264);
nand U13096 (N_13096,N_10869,N_10980);
nand U13097 (N_13097,N_9118,N_9596);
nand U13098 (N_13098,N_9536,N_9630);
nand U13099 (N_13099,N_10430,N_10025);
nor U13100 (N_13100,N_10719,N_11207);
and U13101 (N_13101,N_10300,N_9143);
nand U13102 (N_13102,N_9450,N_11990);
xnor U13103 (N_13103,N_10181,N_10647);
nor U13104 (N_13104,N_11673,N_10319);
xor U13105 (N_13105,N_10522,N_10975);
xnor U13106 (N_13106,N_11724,N_10843);
xnor U13107 (N_13107,N_11719,N_11981);
nand U13108 (N_13108,N_9674,N_10775);
nor U13109 (N_13109,N_9473,N_11856);
or U13110 (N_13110,N_10779,N_9449);
and U13111 (N_13111,N_11812,N_11705);
nor U13112 (N_13112,N_11745,N_11874);
xnor U13113 (N_13113,N_10971,N_10905);
or U13114 (N_13114,N_9592,N_9282);
nor U13115 (N_13115,N_9880,N_11475);
nor U13116 (N_13116,N_9094,N_11038);
or U13117 (N_13117,N_9678,N_10684);
nand U13118 (N_13118,N_10124,N_9716);
nand U13119 (N_13119,N_10495,N_9669);
nand U13120 (N_13120,N_9545,N_9573);
nand U13121 (N_13121,N_10452,N_9427);
or U13122 (N_13122,N_10686,N_11048);
or U13123 (N_13123,N_11987,N_11613);
nand U13124 (N_13124,N_9083,N_10541);
nand U13125 (N_13125,N_9142,N_11113);
nor U13126 (N_13126,N_10044,N_9057);
xnor U13127 (N_13127,N_10803,N_10603);
nor U13128 (N_13128,N_11373,N_9447);
and U13129 (N_13129,N_10240,N_11323);
xor U13130 (N_13130,N_9021,N_10632);
xor U13131 (N_13131,N_9514,N_9200);
and U13132 (N_13132,N_11647,N_9405);
nand U13133 (N_13133,N_11136,N_9020);
or U13134 (N_13134,N_10531,N_11348);
xor U13135 (N_13135,N_10356,N_9658);
or U13136 (N_13136,N_9764,N_9837);
xnor U13137 (N_13137,N_9241,N_9033);
nand U13138 (N_13138,N_9950,N_10904);
and U13139 (N_13139,N_10146,N_9209);
or U13140 (N_13140,N_9336,N_11665);
and U13141 (N_13141,N_9770,N_10566);
nand U13142 (N_13142,N_10965,N_10394);
nor U13143 (N_13143,N_11916,N_10537);
nor U13144 (N_13144,N_11180,N_10534);
or U13145 (N_13145,N_11368,N_11006);
and U13146 (N_13146,N_10458,N_10924);
or U13147 (N_13147,N_11251,N_11221);
xnor U13148 (N_13148,N_11238,N_11847);
xor U13149 (N_13149,N_9391,N_10579);
and U13150 (N_13150,N_9451,N_10913);
and U13151 (N_13151,N_9852,N_11701);
and U13152 (N_13152,N_9500,N_10928);
and U13153 (N_13153,N_9810,N_10793);
nand U13154 (N_13154,N_11227,N_10081);
nand U13155 (N_13155,N_10219,N_11614);
and U13156 (N_13156,N_10435,N_9675);
nor U13157 (N_13157,N_10352,N_10147);
xor U13158 (N_13158,N_10722,N_10692);
or U13159 (N_13159,N_10753,N_9942);
or U13160 (N_13160,N_9334,N_9360);
nand U13161 (N_13161,N_10581,N_10155);
xor U13162 (N_13162,N_10690,N_9645);
and U13163 (N_13163,N_10136,N_10008);
and U13164 (N_13164,N_9460,N_10449);
xor U13165 (N_13165,N_10626,N_10665);
nor U13166 (N_13166,N_9343,N_9089);
nor U13167 (N_13167,N_10682,N_10927);
and U13168 (N_13168,N_10165,N_9621);
or U13169 (N_13169,N_11974,N_9979);
or U13170 (N_13170,N_9180,N_11313);
nor U13171 (N_13171,N_9844,N_9715);
nand U13172 (N_13172,N_11312,N_9213);
and U13173 (N_13173,N_11952,N_10702);
xnor U13174 (N_13174,N_10691,N_10221);
and U13175 (N_13175,N_10855,N_11296);
nand U13176 (N_13176,N_9888,N_11093);
xnor U13177 (N_13177,N_10243,N_11591);
xor U13178 (N_13178,N_10082,N_9964);
and U13179 (N_13179,N_10251,N_9821);
nand U13180 (N_13180,N_11092,N_9011);
and U13181 (N_13181,N_11590,N_9246);
or U13182 (N_13182,N_10933,N_10588);
or U13183 (N_13183,N_9173,N_11934);
and U13184 (N_13184,N_9243,N_9115);
or U13185 (N_13185,N_10373,N_10732);
or U13186 (N_13186,N_10929,N_10277);
nor U13187 (N_13187,N_9506,N_10074);
and U13188 (N_13188,N_11640,N_10950);
and U13189 (N_13189,N_10409,N_9109);
and U13190 (N_13190,N_11255,N_9299);
nor U13191 (N_13191,N_10273,N_11993);
nor U13192 (N_13192,N_10911,N_9170);
or U13193 (N_13193,N_10490,N_9155);
and U13194 (N_13194,N_10960,N_10978);
and U13195 (N_13195,N_9374,N_10111);
nand U13196 (N_13196,N_11433,N_10707);
xnor U13197 (N_13197,N_10570,N_10908);
nor U13198 (N_13198,N_11581,N_11659);
xor U13199 (N_13199,N_9475,N_11776);
nand U13200 (N_13200,N_10206,N_10701);
or U13201 (N_13201,N_9403,N_10964);
nand U13202 (N_13202,N_11058,N_10660);
and U13203 (N_13203,N_11230,N_9580);
nand U13204 (N_13204,N_11973,N_9594);
and U13205 (N_13205,N_10380,N_9424);
xor U13206 (N_13206,N_11695,N_9813);
nor U13207 (N_13207,N_11895,N_10518);
xnor U13208 (N_13208,N_9975,N_9853);
nor U13209 (N_13209,N_9349,N_11414);
nor U13210 (N_13210,N_10807,N_10484);
or U13211 (N_13211,N_9648,N_11118);
nand U13212 (N_13212,N_9560,N_11173);
nor U13213 (N_13213,N_11258,N_11883);
and U13214 (N_13214,N_9303,N_10700);
xnor U13215 (N_13215,N_9022,N_9561);
nand U13216 (N_13216,N_10628,N_11519);
nand U13217 (N_13217,N_9060,N_10269);
xnor U13218 (N_13218,N_9070,N_11683);
and U13219 (N_13219,N_10407,N_9981);
nor U13220 (N_13220,N_11820,N_9693);
xor U13221 (N_13221,N_10292,N_9894);
xor U13222 (N_13222,N_11328,N_10510);
nand U13223 (N_13223,N_9423,N_10835);
or U13224 (N_13224,N_9781,N_11205);
nand U13225 (N_13225,N_11797,N_10169);
nand U13226 (N_13226,N_10371,N_11516);
or U13227 (N_13227,N_10454,N_9801);
nor U13228 (N_13228,N_10355,N_9338);
nor U13229 (N_13229,N_11710,N_9058);
or U13230 (N_13230,N_9371,N_9225);
nand U13231 (N_13231,N_11416,N_9315);
or U13232 (N_13232,N_11828,N_9497);
or U13233 (N_13233,N_11426,N_10634);
nor U13234 (N_13234,N_10466,N_10471);
nand U13235 (N_13235,N_11098,N_11986);
or U13236 (N_13236,N_9689,N_11009);
or U13237 (N_13237,N_9534,N_10416);
nand U13238 (N_13238,N_9904,N_10107);
and U13239 (N_13239,N_11427,N_11933);
or U13240 (N_13240,N_10907,N_11531);
nor U13241 (N_13241,N_10930,N_11124);
nor U13242 (N_13242,N_11077,N_9794);
xnor U13243 (N_13243,N_10944,N_11722);
nand U13244 (N_13244,N_10931,N_10780);
xor U13245 (N_13245,N_9324,N_9955);
xnor U13246 (N_13246,N_11219,N_10328);
nand U13247 (N_13247,N_11732,N_9007);
nand U13248 (N_13248,N_10674,N_10193);
xnor U13249 (N_13249,N_10268,N_10278);
or U13250 (N_13250,N_11780,N_11699);
and U13251 (N_13251,N_9214,N_11030);
nor U13252 (N_13252,N_10947,N_9456);
or U13253 (N_13253,N_9655,N_10365);
nand U13254 (N_13254,N_10118,N_10473);
xor U13255 (N_13255,N_11229,N_11622);
or U13256 (N_13256,N_9223,N_11772);
or U13257 (N_13257,N_10919,N_10264);
and U13258 (N_13258,N_10105,N_11677);
xor U13259 (N_13259,N_10642,N_9863);
and U13260 (N_13260,N_10694,N_11890);
nor U13261 (N_13261,N_9212,N_9161);
nand U13262 (N_13262,N_11356,N_9135);
nor U13263 (N_13263,N_11707,N_11689);
or U13264 (N_13264,N_10174,N_9014);
xor U13265 (N_13265,N_10131,N_11233);
xor U13266 (N_13266,N_10608,N_11363);
nand U13267 (N_13267,N_9847,N_10168);
xor U13268 (N_13268,N_11822,N_9318);
or U13269 (N_13269,N_11540,N_11185);
nor U13270 (N_13270,N_10031,N_10559);
nor U13271 (N_13271,N_11664,N_11537);
xor U13272 (N_13272,N_10550,N_9839);
xnor U13273 (N_13273,N_10912,N_10487);
and U13274 (N_13274,N_9040,N_9120);
and U13275 (N_13275,N_10072,N_11829);
or U13276 (N_13276,N_9099,N_9840);
and U13277 (N_13277,N_11398,N_9304);
or U13278 (N_13278,N_10241,N_9250);
or U13279 (N_13279,N_10554,N_11110);
nand U13280 (N_13280,N_10167,N_11637);
nor U13281 (N_13281,N_9140,N_9760);
or U13282 (N_13282,N_11089,N_11439);
nor U13283 (N_13283,N_9372,N_11293);
nor U13284 (N_13284,N_11459,N_11226);
or U13285 (N_13285,N_11858,N_10741);
or U13286 (N_13286,N_9884,N_9097);
or U13287 (N_13287,N_9469,N_9294);
nor U13288 (N_13288,N_11569,N_11778);
or U13289 (N_13289,N_9248,N_11985);
xnor U13290 (N_13290,N_9435,N_11295);
nor U13291 (N_13291,N_9176,N_10198);
and U13292 (N_13292,N_9753,N_10953);
xor U13293 (N_13293,N_11593,N_10983);
nand U13294 (N_13294,N_9815,N_10590);
xor U13295 (N_13295,N_9018,N_10119);
nor U13296 (N_13296,N_9740,N_10427);
nand U13297 (N_13297,N_10272,N_9685);
nand U13298 (N_13298,N_10417,N_9746);
nor U13299 (N_13299,N_9518,N_9095);
and U13300 (N_13300,N_9141,N_9627);
or U13301 (N_13301,N_11350,N_9858);
and U13302 (N_13302,N_11096,N_10872);
nand U13303 (N_13303,N_9503,N_11100);
nand U13304 (N_13304,N_10675,N_10283);
xnor U13305 (N_13305,N_9718,N_9791);
nor U13306 (N_13306,N_10387,N_10708);
nand U13307 (N_13307,N_10420,N_10601);
and U13308 (N_13308,N_10322,N_9483);
nand U13309 (N_13309,N_9897,N_11364);
xor U13310 (N_13310,N_10000,N_10393);
nand U13311 (N_13311,N_9635,N_11956);
nor U13312 (N_13312,N_11930,N_9584);
or U13313 (N_13313,N_11387,N_11700);
xor U13314 (N_13314,N_10297,N_11248);
nor U13315 (N_13315,N_11245,N_11530);
or U13316 (N_13316,N_11101,N_11365);
and U13317 (N_13317,N_11889,N_10891);
and U13318 (N_13318,N_10228,N_11853);
nand U13319 (N_13319,N_10129,N_9148);
nand U13320 (N_13320,N_10898,N_9144);
nand U13321 (N_13321,N_9127,N_11375);
nand U13322 (N_13322,N_10359,N_10063);
xor U13323 (N_13323,N_11805,N_9052);
and U13324 (N_13324,N_10530,N_9395);
and U13325 (N_13325,N_11765,N_10676);
xnor U13326 (N_13326,N_10648,N_9948);
and U13327 (N_13327,N_9795,N_10114);
nor U13328 (N_13328,N_10067,N_9803);
nor U13329 (N_13329,N_11386,N_10606);
nand U13330 (N_13330,N_11085,N_10202);
and U13331 (N_13331,N_9640,N_10610);
and U13332 (N_13332,N_10364,N_10756);
xnor U13333 (N_13333,N_10997,N_10005);
xor U13334 (N_13334,N_11413,N_9719);
or U13335 (N_13335,N_9714,N_11716);
nand U13336 (N_13336,N_11177,N_9958);
and U13337 (N_13337,N_9624,N_11388);
nor U13338 (N_13338,N_9285,N_10222);
nor U13339 (N_13339,N_10160,N_9232);
nand U13340 (N_13340,N_11811,N_11915);
nor U13341 (N_13341,N_11506,N_11351);
and U13342 (N_13342,N_11742,N_9458);
nor U13343 (N_13343,N_10832,N_9551);
nand U13344 (N_13344,N_10488,N_11680);
or U13345 (N_13345,N_10961,N_10455);
xnor U13346 (N_13346,N_10568,N_11421);
nor U13347 (N_13347,N_9792,N_9988);
and U13348 (N_13348,N_9269,N_10401);
and U13349 (N_13349,N_10683,N_10154);
nand U13350 (N_13350,N_10246,N_9850);
xnor U13351 (N_13351,N_11877,N_10787);
and U13352 (N_13352,N_10175,N_10383);
xnor U13353 (N_13353,N_9912,N_11612);
nor U13354 (N_13354,N_10301,N_10043);
and U13355 (N_13355,N_11142,N_9745);
or U13356 (N_13356,N_9409,N_10942);
or U13357 (N_13357,N_11220,N_11198);
or U13358 (N_13358,N_9602,N_11029);
nand U13359 (N_13359,N_11165,N_9566);
nor U13360 (N_13360,N_11063,N_11961);
and U13361 (N_13361,N_10706,N_10893);
and U13362 (N_13362,N_11310,N_10353);
nor U13363 (N_13363,N_9311,N_10728);
or U13364 (N_13364,N_9006,N_11201);
nand U13365 (N_13365,N_9157,N_9974);
and U13366 (N_13366,N_9893,N_11408);
and U13367 (N_13367,N_10866,N_10549);
or U13368 (N_13368,N_11033,N_11620);
or U13369 (N_13369,N_11864,N_11656);
or U13370 (N_13370,N_10761,N_9934);
xor U13371 (N_13371,N_11550,N_11575);
or U13372 (N_13372,N_9824,N_11492);
and U13373 (N_13373,N_10516,N_10846);
nand U13374 (N_13374,N_9717,N_10696);
and U13375 (N_13375,N_10019,N_10034);
xor U13376 (N_13376,N_9383,N_11548);
or U13377 (N_13377,N_9841,N_11970);
nor U13378 (N_13378,N_9486,N_9032);
nor U13379 (N_13379,N_9891,N_11535);
or U13380 (N_13380,N_11542,N_10152);
or U13381 (N_13381,N_9001,N_11903);
nor U13382 (N_13382,N_10094,N_10782);
xor U13383 (N_13383,N_10653,N_9797);
and U13384 (N_13384,N_9009,N_9117);
nor U13385 (N_13385,N_9711,N_11463);
xor U13386 (N_13386,N_9807,N_9659);
xor U13387 (N_13387,N_11473,N_10345);
nor U13388 (N_13388,N_10318,N_10672);
and U13389 (N_13389,N_11076,N_9367);
and U13390 (N_13390,N_10798,N_11075);
and U13391 (N_13391,N_10542,N_9415);
nand U13392 (N_13392,N_9292,N_11176);
xnor U13393 (N_13393,N_11265,N_11527);
nand U13394 (N_13394,N_9199,N_9271);
nand U13395 (N_13395,N_10071,N_9985);
nand U13396 (N_13396,N_9345,N_9370);
nor U13397 (N_13397,N_9606,N_11488);
nand U13398 (N_13398,N_10989,N_11690);
and U13399 (N_13399,N_11362,N_10824);
xor U13400 (N_13400,N_11870,N_11606);
and U13401 (N_13401,N_9494,N_9342);
nand U13402 (N_13402,N_11893,N_11134);
nand U13403 (N_13403,N_10486,N_10436);
or U13404 (N_13404,N_11035,N_11129);
xnor U13405 (N_13405,N_9782,N_11187);
xnor U13406 (N_13406,N_9204,N_9078);
nor U13407 (N_13407,N_11239,N_11624);
xnor U13408 (N_13408,N_10899,N_11760);
nand U13409 (N_13409,N_9593,N_11034);
and U13410 (N_13410,N_11863,N_11446);
xnor U13411 (N_13411,N_10400,N_11566);
and U13412 (N_13412,N_9123,N_10595);
nand U13413 (N_13413,N_11431,N_9558);
nor U13414 (N_13414,N_11271,N_11927);
or U13415 (N_13415,N_10999,N_9598);
or U13416 (N_13416,N_9907,N_9426);
xnor U13417 (N_13417,N_9544,N_10209);
nor U13418 (N_13418,N_10519,N_10467);
and U13419 (N_13419,N_10414,N_9499);
nand U13420 (N_13420,N_10876,N_10731);
nor U13421 (N_13421,N_10952,N_11260);
nand U13422 (N_13422,N_10038,N_10086);
xnor U13423 (N_13423,N_11199,N_10575);
or U13424 (N_13424,N_11715,N_11195);
and U13425 (N_13425,N_11549,N_10727);
nand U13426 (N_13426,N_9139,N_10410);
and U13427 (N_13427,N_11739,N_10161);
nand U13428 (N_13428,N_9273,N_9901);
or U13429 (N_13429,N_10523,N_9747);
or U13430 (N_13430,N_11374,N_11894);
or U13431 (N_13431,N_11586,N_10068);
xnor U13432 (N_13432,N_10441,N_10956);
nand U13433 (N_13433,N_9854,N_10627);
and U13434 (N_13434,N_10871,N_11963);
or U13435 (N_13435,N_11069,N_10988);
and U13436 (N_13436,N_11769,N_11599);
nor U13437 (N_13437,N_11186,N_9129);
and U13438 (N_13438,N_11254,N_10751);
xor U13439 (N_13439,N_9330,N_9188);
or U13440 (N_13440,N_10827,N_9516);
and U13441 (N_13441,N_11844,N_10658);
and U13442 (N_13442,N_9461,N_10375);
or U13443 (N_13443,N_10156,N_11679);
or U13444 (N_13444,N_9356,N_10225);
nor U13445 (N_13445,N_11499,N_10576);
or U13446 (N_13446,N_11432,N_10894);
or U13447 (N_13447,N_11002,N_9846);
xor U13448 (N_13448,N_10257,N_11290);
nand U13449 (N_13449,N_10923,N_11955);
xor U13450 (N_13450,N_11200,N_10635);
and U13451 (N_13451,N_11957,N_9708);
nand U13452 (N_13452,N_10053,N_11300);
and U13453 (N_13453,N_9418,N_11051);
xnor U13454 (N_13454,N_11366,N_11094);
nand U13455 (N_13455,N_9388,N_11149);
xnor U13456 (N_13456,N_11420,N_9917);
xnor U13457 (N_13457,N_9619,N_11253);
or U13458 (N_13458,N_11429,N_9713);
and U13459 (N_13459,N_10792,N_11674);
nor U13460 (N_13460,N_11929,N_9644);
nor U13461 (N_13461,N_9778,N_9637);
or U13462 (N_13462,N_9425,N_9351);
nor U13463 (N_13463,N_9924,N_10976);
nand U13464 (N_13464,N_11137,N_9639);
or U13465 (N_13465,N_10227,N_9812);
nor U13466 (N_13466,N_9298,N_11618);
and U13467 (N_13467,N_10226,N_11483);
xor U13468 (N_13468,N_9905,N_10437);
xor U13469 (N_13469,N_9031,N_9008);
nor U13470 (N_13470,N_10506,N_11438);
nor U13471 (N_13471,N_10491,N_11495);
nand U13472 (N_13472,N_10539,N_11244);
and U13473 (N_13473,N_11825,N_9479);
nor U13474 (N_13474,N_10704,N_9390);
nand U13475 (N_13475,N_11277,N_9582);
xor U13476 (N_13476,N_10698,N_10825);
nor U13477 (N_13477,N_10667,N_9054);
nor U13478 (N_13478,N_9226,N_10474);
nor U13479 (N_13479,N_9487,N_10963);
and U13480 (N_13480,N_11958,N_11936);
nand U13481 (N_13481,N_11522,N_9618);
nand U13482 (N_13482,N_9736,N_11615);
nor U13483 (N_13483,N_10478,N_10009);
nand U13484 (N_13484,N_11919,N_11907);
or U13485 (N_13485,N_9357,N_11866);
nor U13486 (N_13486,N_11552,N_11643);
or U13487 (N_13487,N_11236,N_10392);
or U13488 (N_13488,N_10498,N_10502);
xnor U13489 (N_13489,N_10656,N_11661);
nor U13490 (N_13490,N_9108,N_11202);
nand U13491 (N_13491,N_9211,N_10200);
xor U13492 (N_13492,N_10986,N_10288);
or U13493 (N_13493,N_10734,N_11208);
nand U13494 (N_13494,N_9384,N_11091);
xor U13495 (N_13495,N_10990,N_10013);
nor U13496 (N_13496,N_10589,N_9152);
xnor U13497 (N_13497,N_10820,N_11418);
nand U13498 (N_13498,N_11169,N_11786);
or U13499 (N_13499,N_11717,N_9385);
or U13500 (N_13500,N_11110,N_9262);
xnor U13501 (N_13501,N_10943,N_10536);
nand U13502 (N_13502,N_11992,N_10299);
or U13503 (N_13503,N_10591,N_9213);
xnor U13504 (N_13504,N_11123,N_9142);
xor U13505 (N_13505,N_11782,N_10368);
xor U13506 (N_13506,N_11559,N_10246);
or U13507 (N_13507,N_9189,N_11247);
nor U13508 (N_13508,N_11212,N_11312);
and U13509 (N_13509,N_9140,N_9990);
xnor U13510 (N_13510,N_10710,N_9856);
xor U13511 (N_13511,N_9535,N_9211);
xor U13512 (N_13512,N_11941,N_9608);
and U13513 (N_13513,N_9207,N_9045);
nand U13514 (N_13514,N_10615,N_10028);
xor U13515 (N_13515,N_11100,N_10364);
or U13516 (N_13516,N_10487,N_11463);
and U13517 (N_13517,N_11098,N_9679);
or U13518 (N_13518,N_11077,N_10981);
xor U13519 (N_13519,N_9643,N_9007);
and U13520 (N_13520,N_9328,N_10408);
xor U13521 (N_13521,N_11983,N_10564);
and U13522 (N_13522,N_10830,N_11255);
or U13523 (N_13523,N_11175,N_11553);
nand U13524 (N_13524,N_9684,N_10363);
xor U13525 (N_13525,N_9530,N_11328);
or U13526 (N_13526,N_11945,N_10315);
nor U13527 (N_13527,N_10872,N_9455);
nor U13528 (N_13528,N_10746,N_9962);
nand U13529 (N_13529,N_9120,N_11783);
and U13530 (N_13530,N_10649,N_9809);
or U13531 (N_13531,N_10880,N_9022);
and U13532 (N_13532,N_9933,N_9562);
xnor U13533 (N_13533,N_11745,N_9840);
or U13534 (N_13534,N_9461,N_9846);
and U13535 (N_13535,N_11827,N_11710);
or U13536 (N_13536,N_10646,N_10191);
nor U13537 (N_13537,N_10079,N_9322);
xnor U13538 (N_13538,N_9077,N_11789);
xnor U13539 (N_13539,N_11627,N_9413);
and U13540 (N_13540,N_10165,N_9901);
or U13541 (N_13541,N_9428,N_9429);
or U13542 (N_13542,N_10229,N_9105);
and U13543 (N_13543,N_9563,N_9919);
and U13544 (N_13544,N_11319,N_11988);
and U13545 (N_13545,N_9289,N_11705);
nor U13546 (N_13546,N_9859,N_9033);
and U13547 (N_13547,N_10641,N_11916);
or U13548 (N_13548,N_10409,N_11420);
xor U13549 (N_13549,N_10624,N_11538);
nor U13550 (N_13550,N_9285,N_9540);
or U13551 (N_13551,N_11054,N_9609);
and U13552 (N_13552,N_9004,N_10598);
nand U13553 (N_13553,N_10044,N_10217);
nand U13554 (N_13554,N_10660,N_10338);
nand U13555 (N_13555,N_11811,N_11637);
nor U13556 (N_13556,N_10340,N_11096);
nand U13557 (N_13557,N_9760,N_9594);
xnor U13558 (N_13558,N_10419,N_11574);
xor U13559 (N_13559,N_9038,N_10548);
nand U13560 (N_13560,N_9655,N_11984);
or U13561 (N_13561,N_10564,N_10695);
nor U13562 (N_13562,N_9813,N_9048);
and U13563 (N_13563,N_11828,N_9400);
nand U13564 (N_13564,N_10663,N_9666);
nand U13565 (N_13565,N_9336,N_9648);
xor U13566 (N_13566,N_11333,N_9181);
and U13567 (N_13567,N_11572,N_10927);
or U13568 (N_13568,N_11549,N_10141);
xor U13569 (N_13569,N_11981,N_11661);
nor U13570 (N_13570,N_10381,N_11802);
or U13571 (N_13571,N_10081,N_9962);
nor U13572 (N_13572,N_9199,N_11915);
nor U13573 (N_13573,N_9055,N_9988);
and U13574 (N_13574,N_9682,N_9589);
xnor U13575 (N_13575,N_9077,N_10125);
xnor U13576 (N_13576,N_10727,N_11189);
xor U13577 (N_13577,N_11427,N_10955);
nand U13578 (N_13578,N_9530,N_9309);
or U13579 (N_13579,N_11588,N_11151);
xnor U13580 (N_13580,N_9909,N_11628);
and U13581 (N_13581,N_9607,N_9168);
nand U13582 (N_13582,N_10468,N_11024);
or U13583 (N_13583,N_10810,N_9481);
nand U13584 (N_13584,N_11715,N_9384);
nor U13585 (N_13585,N_10316,N_9341);
nand U13586 (N_13586,N_10042,N_11432);
nand U13587 (N_13587,N_10511,N_9307);
xor U13588 (N_13588,N_9296,N_11271);
nor U13589 (N_13589,N_9778,N_11041);
xnor U13590 (N_13590,N_11902,N_11101);
or U13591 (N_13591,N_10784,N_10645);
or U13592 (N_13592,N_9801,N_11400);
nor U13593 (N_13593,N_10699,N_10409);
nand U13594 (N_13594,N_11146,N_11603);
xnor U13595 (N_13595,N_11000,N_11614);
xor U13596 (N_13596,N_10557,N_9264);
nand U13597 (N_13597,N_11513,N_10931);
nor U13598 (N_13598,N_10858,N_11279);
nand U13599 (N_13599,N_9202,N_11975);
and U13600 (N_13600,N_10894,N_9904);
or U13601 (N_13601,N_10645,N_11778);
nand U13602 (N_13602,N_11409,N_9777);
and U13603 (N_13603,N_11041,N_11613);
xor U13604 (N_13604,N_10599,N_11196);
xnor U13605 (N_13605,N_9021,N_9833);
or U13606 (N_13606,N_9246,N_11785);
xor U13607 (N_13607,N_11644,N_10439);
nand U13608 (N_13608,N_9873,N_11841);
or U13609 (N_13609,N_9517,N_11801);
nand U13610 (N_13610,N_10901,N_10562);
xor U13611 (N_13611,N_11914,N_11024);
and U13612 (N_13612,N_11161,N_11590);
nor U13613 (N_13613,N_10477,N_10245);
nor U13614 (N_13614,N_11822,N_9233);
or U13615 (N_13615,N_11934,N_9436);
nand U13616 (N_13616,N_10553,N_11760);
and U13617 (N_13617,N_10801,N_11786);
or U13618 (N_13618,N_11838,N_9711);
nor U13619 (N_13619,N_10619,N_9860);
nand U13620 (N_13620,N_11616,N_11045);
xor U13621 (N_13621,N_9816,N_10147);
nor U13622 (N_13622,N_9921,N_11318);
or U13623 (N_13623,N_11103,N_9208);
nand U13624 (N_13624,N_9575,N_11293);
nand U13625 (N_13625,N_9946,N_11098);
xnor U13626 (N_13626,N_10688,N_10514);
nor U13627 (N_13627,N_9927,N_9396);
or U13628 (N_13628,N_10850,N_9978);
nand U13629 (N_13629,N_11265,N_11199);
and U13630 (N_13630,N_10088,N_9573);
xnor U13631 (N_13631,N_9304,N_10038);
xnor U13632 (N_13632,N_11894,N_11053);
nand U13633 (N_13633,N_11697,N_9128);
xor U13634 (N_13634,N_11247,N_9491);
or U13635 (N_13635,N_9230,N_10330);
or U13636 (N_13636,N_9712,N_10024);
and U13637 (N_13637,N_10129,N_11631);
or U13638 (N_13638,N_10710,N_11480);
and U13639 (N_13639,N_9760,N_11339);
nand U13640 (N_13640,N_10398,N_10005);
nand U13641 (N_13641,N_9812,N_9902);
nand U13642 (N_13642,N_9413,N_10696);
and U13643 (N_13643,N_9549,N_11542);
nor U13644 (N_13644,N_9883,N_9360);
xor U13645 (N_13645,N_9119,N_11002);
nor U13646 (N_13646,N_9347,N_9899);
or U13647 (N_13647,N_10734,N_9889);
and U13648 (N_13648,N_9382,N_11508);
nand U13649 (N_13649,N_10879,N_10560);
nand U13650 (N_13650,N_9628,N_9013);
and U13651 (N_13651,N_10645,N_11242);
and U13652 (N_13652,N_10546,N_11163);
nor U13653 (N_13653,N_9915,N_11774);
nand U13654 (N_13654,N_11954,N_9657);
nand U13655 (N_13655,N_9341,N_10620);
xnor U13656 (N_13656,N_11576,N_10178);
and U13657 (N_13657,N_10619,N_9474);
nand U13658 (N_13658,N_9344,N_9104);
nand U13659 (N_13659,N_11174,N_11376);
nor U13660 (N_13660,N_10890,N_9177);
nand U13661 (N_13661,N_11483,N_9525);
and U13662 (N_13662,N_10188,N_11484);
nor U13663 (N_13663,N_11627,N_11474);
xnor U13664 (N_13664,N_11860,N_10962);
xnor U13665 (N_13665,N_9111,N_11408);
nand U13666 (N_13666,N_11779,N_9387);
or U13667 (N_13667,N_9452,N_9178);
xor U13668 (N_13668,N_9895,N_11602);
xnor U13669 (N_13669,N_9067,N_9157);
xor U13670 (N_13670,N_11033,N_10194);
nor U13671 (N_13671,N_9537,N_10548);
nor U13672 (N_13672,N_10847,N_10532);
and U13673 (N_13673,N_11757,N_11224);
xnor U13674 (N_13674,N_9782,N_11052);
and U13675 (N_13675,N_10513,N_9348);
and U13676 (N_13676,N_10536,N_11128);
nor U13677 (N_13677,N_10994,N_10023);
or U13678 (N_13678,N_9303,N_9082);
and U13679 (N_13679,N_10623,N_11559);
or U13680 (N_13680,N_9296,N_10692);
xnor U13681 (N_13681,N_11811,N_11310);
and U13682 (N_13682,N_9069,N_10162);
nor U13683 (N_13683,N_11090,N_9980);
or U13684 (N_13684,N_10282,N_11576);
or U13685 (N_13685,N_11640,N_11123);
or U13686 (N_13686,N_10816,N_10569);
xnor U13687 (N_13687,N_11327,N_9273);
and U13688 (N_13688,N_9074,N_9096);
or U13689 (N_13689,N_9536,N_10054);
and U13690 (N_13690,N_10193,N_9634);
nand U13691 (N_13691,N_11845,N_10521);
nor U13692 (N_13692,N_9565,N_11808);
xor U13693 (N_13693,N_10750,N_9553);
and U13694 (N_13694,N_11132,N_10145);
nand U13695 (N_13695,N_9446,N_10188);
xor U13696 (N_13696,N_10931,N_11069);
or U13697 (N_13697,N_10812,N_10072);
nand U13698 (N_13698,N_11266,N_11106);
and U13699 (N_13699,N_11571,N_9313);
and U13700 (N_13700,N_10265,N_9684);
and U13701 (N_13701,N_9123,N_10350);
and U13702 (N_13702,N_9243,N_11869);
and U13703 (N_13703,N_11434,N_9654);
and U13704 (N_13704,N_10307,N_9917);
nor U13705 (N_13705,N_9878,N_11638);
and U13706 (N_13706,N_11211,N_11667);
or U13707 (N_13707,N_10011,N_9666);
nor U13708 (N_13708,N_9255,N_10109);
nand U13709 (N_13709,N_11470,N_10685);
nor U13710 (N_13710,N_9915,N_11330);
xor U13711 (N_13711,N_10774,N_10267);
and U13712 (N_13712,N_10387,N_11460);
and U13713 (N_13713,N_11363,N_11477);
or U13714 (N_13714,N_11015,N_11378);
xor U13715 (N_13715,N_9444,N_11175);
nor U13716 (N_13716,N_10275,N_10186);
and U13717 (N_13717,N_9486,N_10145);
xnor U13718 (N_13718,N_9163,N_9222);
nor U13719 (N_13719,N_11795,N_9475);
or U13720 (N_13720,N_11049,N_11215);
nand U13721 (N_13721,N_9538,N_10736);
nor U13722 (N_13722,N_11367,N_11797);
nand U13723 (N_13723,N_11817,N_9510);
nor U13724 (N_13724,N_9944,N_11816);
and U13725 (N_13725,N_9964,N_10083);
nor U13726 (N_13726,N_9369,N_9376);
or U13727 (N_13727,N_11304,N_11679);
nor U13728 (N_13728,N_10395,N_11584);
xnor U13729 (N_13729,N_10101,N_10583);
xor U13730 (N_13730,N_10819,N_10401);
or U13731 (N_13731,N_11859,N_9423);
nor U13732 (N_13732,N_11276,N_9883);
nor U13733 (N_13733,N_11352,N_10801);
nand U13734 (N_13734,N_11724,N_9804);
and U13735 (N_13735,N_11347,N_9088);
nand U13736 (N_13736,N_11523,N_9383);
and U13737 (N_13737,N_11831,N_11618);
or U13738 (N_13738,N_11074,N_10795);
nand U13739 (N_13739,N_11946,N_11763);
xnor U13740 (N_13740,N_9505,N_10015);
or U13741 (N_13741,N_9586,N_9472);
nand U13742 (N_13742,N_11790,N_11622);
nand U13743 (N_13743,N_11918,N_10269);
nor U13744 (N_13744,N_9669,N_10156);
or U13745 (N_13745,N_9970,N_9537);
or U13746 (N_13746,N_10629,N_10811);
or U13747 (N_13747,N_9473,N_9638);
or U13748 (N_13748,N_10006,N_10709);
and U13749 (N_13749,N_11358,N_9256);
and U13750 (N_13750,N_11361,N_11207);
xnor U13751 (N_13751,N_9850,N_9698);
xnor U13752 (N_13752,N_9913,N_11464);
nor U13753 (N_13753,N_10429,N_10447);
nand U13754 (N_13754,N_10088,N_10055);
and U13755 (N_13755,N_9526,N_9456);
nor U13756 (N_13756,N_10451,N_9592);
nor U13757 (N_13757,N_10821,N_9169);
and U13758 (N_13758,N_11155,N_11281);
nor U13759 (N_13759,N_11635,N_9441);
or U13760 (N_13760,N_11988,N_9217);
or U13761 (N_13761,N_11485,N_11543);
or U13762 (N_13762,N_11676,N_9610);
nand U13763 (N_13763,N_10760,N_11663);
nand U13764 (N_13764,N_11275,N_11314);
xnor U13765 (N_13765,N_10267,N_10891);
or U13766 (N_13766,N_11610,N_10588);
xor U13767 (N_13767,N_10320,N_11212);
nor U13768 (N_13768,N_11759,N_11237);
xnor U13769 (N_13769,N_11234,N_9949);
xor U13770 (N_13770,N_11651,N_10678);
and U13771 (N_13771,N_11748,N_11200);
and U13772 (N_13772,N_9889,N_10090);
nor U13773 (N_13773,N_11197,N_9619);
nor U13774 (N_13774,N_10332,N_9802);
and U13775 (N_13775,N_9417,N_10133);
xor U13776 (N_13776,N_9524,N_10629);
or U13777 (N_13777,N_10850,N_11883);
xor U13778 (N_13778,N_10188,N_9159);
xor U13779 (N_13779,N_10626,N_10985);
nor U13780 (N_13780,N_9739,N_11788);
xnor U13781 (N_13781,N_9849,N_10152);
nor U13782 (N_13782,N_9940,N_9644);
nor U13783 (N_13783,N_10620,N_10226);
nand U13784 (N_13784,N_9903,N_10309);
xor U13785 (N_13785,N_10777,N_10582);
nor U13786 (N_13786,N_9019,N_9838);
or U13787 (N_13787,N_11535,N_9922);
xor U13788 (N_13788,N_11361,N_11437);
xor U13789 (N_13789,N_11206,N_9722);
nor U13790 (N_13790,N_9394,N_10366);
nor U13791 (N_13791,N_10917,N_10088);
and U13792 (N_13792,N_9005,N_10388);
and U13793 (N_13793,N_10500,N_10852);
nor U13794 (N_13794,N_9634,N_11123);
xnor U13795 (N_13795,N_10319,N_9987);
nor U13796 (N_13796,N_11534,N_11543);
xnor U13797 (N_13797,N_10636,N_11534);
nor U13798 (N_13798,N_9102,N_9446);
and U13799 (N_13799,N_10067,N_9896);
nand U13800 (N_13800,N_11797,N_10508);
and U13801 (N_13801,N_9996,N_10624);
nor U13802 (N_13802,N_10590,N_11236);
and U13803 (N_13803,N_11420,N_10307);
and U13804 (N_13804,N_10417,N_11014);
or U13805 (N_13805,N_9111,N_11040);
or U13806 (N_13806,N_10602,N_9288);
and U13807 (N_13807,N_10038,N_10212);
or U13808 (N_13808,N_9944,N_9433);
or U13809 (N_13809,N_10747,N_10899);
and U13810 (N_13810,N_10853,N_9198);
or U13811 (N_13811,N_11533,N_9463);
xnor U13812 (N_13812,N_9009,N_10821);
nand U13813 (N_13813,N_9171,N_10307);
xnor U13814 (N_13814,N_11744,N_10255);
and U13815 (N_13815,N_11091,N_9478);
nor U13816 (N_13816,N_9639,N_10841);
and U13817 (N_13817,N_11512,N_11030);
or U13818 (N_13818,N_10250,N_11531);
xnor U13819 (N_13819,N_10941,N_10427);
nor U13820 (N_13820,N_11510,N_9842);
xnor U13821 (N_13821,N_11137,N_9881);
xnor U13822 (N_13822,N_10755,N_9786);
and U13823 (N_13823,N_11759,N_11844);
nor U13824 (N_13824,N_9698,N_10789);
and U13825 (N_13825,N_9047,N_9355);
or U13826 (N_13826,N_11043,N_11064);
xor U13827 (N_13827,N_9274,N_9283);
nor U13828 (N_13828,N_10478,N_11140);
and U13829 (N_13829,N_9826,N_9062);
nor U13830 (N_13830,N_11784,N_10965);
nand U13831 (N_13831,N_10383,N_9612);
xnor U13832 (N_13832,N_9754,N_11955);
or U13833 (N_13833,N_11123,N_10044);
or U13834 (N_13834,N_10364,N_10903);
nand U13835 (N_13835,N_10630,N_9336);
and U13836 (N_13836,N_9633,N_9393);
nor U13837 (N_13837,N_9024,N_11015);
nand U13838 (N_13838,N_9047,N_11471);
nor U13839 (N_13839,N_10801,N_11030);
or U13840 (N_13840,N_9303,N_11111);
xor U13841 (N_13841,N_9943,N_9646);
nor U13842 (N_13842,N_10057,N_10880);
nor U13843 (N_13843,N_10779,N_11352);
nor U13844 (N_13844,N_10268,N_9306);
xor U13845 (N_13845,N_11983,N_9992);
nor U13846 (N_13846,N_10529,N_10870);
and U13847 (N_13847,N_10101,N_9179);
nor U13848 (N_13848,N_11804,N_10759);
or U13849 (N_13849,N_9892,N_10856);
nand U13850 (N_13850,N_10089,N_9051);
and U13851 (N_13851,N_9806,N_11756);
or U13852 (N_13852,N_11166,N_11665);
or U13853 (N_13853,N_11975,N_11711);
xnor U13854 (N_13854,N_11681,N_9219);
and U13855 (N_13855,N_10700,N_9850);
and U13856 (N_13856,N_9969,N_10647);
or U13857 (N_13857,N_11285,N_10878);
or U13858 (N_13858,N_11030,N_10212);
and U13859 (N_13859,N_11971,N_11188);
and U13860 (N_13860,N_9477,N_11822);
xor U13861 (N_13861,N_10891,N_9165);
and U13862 (N_13862,N_11818,N_10007);
nor U13863 (N_13863,N_10807,N_9476);
nand U13864 (N_13864,N_10098,N_10626);
nand U13865 (N_13865,N_10383,N_10489);
or U13866 (N_13866,N_10431,N_10603);
nand U13867 (N_13867,N_9332,N_9979);
nor U13868 (N_13868,N_11023,N_11562);
nand U13869 (N_13869,N_10919,N_11633);
nand U13870 (N_13870,N_10267,N_10650);
xor U13871 (N_13871,N_10776,N_11271);
xor U13872 (N_13872,N_11294,N_10497);
xnor U13873 (N_13873,N_10004,N_9350);
nor U13874 (N_13874,N_10793,N_10058);
nand U13875 (N_13875,N_9766,N_10929);
or U13876 (N_13876,N_9966,N_9149);
or U13877 (N_13877,N_10467,N_10734);
and U13878 (N_13878,N_9585,N_10019);
xnor U13879 (N_13879,N_9036,N_10614);
nor U13880 (N_13880,N_10530,N_11484);
or U13881 (N_13881,N_10423,N_9910);
or U13882 (N_13882,N_9865,N_11357);
and U13883 (N_13883,N_11711,N_11614);
and U13884 (N_13884,N_9855,N_11700);
and U13885 (N_13885,N_11723,N_11257);
or U13886 (N_13886,N_10194,N_11190);
or U13887 (N_13887,N_11294,N_10000);
and U13888 (N_13888,N_10805,N_11201);
or U13889 (N_13889,N_9404,N_9837);
nand U13890 (N_13890,N_9956,N_9885);
nor U13891 (N_13891,N_9211,N_11202);
or U13892 (N_13892,N_10886,N_11000);
or U13893 (N_13893,N_10296,N_11583);
or U13894 (N_13894,N_10521,N_11145);
nor U13895 (N_13895,N_10911,N_9713);
nor U13896 (N_13896,N_10418,N_9077);
nor U13897 (N_13897,N_10595,N_9839);
and U13898 (N_13898,N_10274,N_11483);
nand U13899 (N_13899,N_11023,N_10471);
and U13900 (N_13900,N_11025,N_10965);
nor U13901 (N_13901,N_9529,N_11241);
and U13902 (N_13902,N_9729,N_10850);
and U13903 (N_13903,N_9573,N_9224);
or U13904 (N_13904,N_10983,N_10536);
xor U13905 (N_13905,N_11404,N_11686);
and U13906 (N_13906,N_11844,N_10485);
xor U13907 (N_13907,N_11341,N_10883);
or U13908 (N_13908,N_11178,N_11211);
and U13909 (N_13909,N_9159,N_10468);
nor U13910 (N_13910,N_11224,N_10938);
or U13911 (N_13911,N_9076,N_9406);
nand U13912 (N_13912,N_11320,N_9617);
nor U13913 (N_13913,N_11574,N_10022);
nand U13914 (N_13914,N_9848,N_11703);
xor U13915 (N_13915,N_9014,N_9876);
or U13916 (N_13916,N_10845,N_11516);
and U13917 (N_13917,N_11144,N_10944);
nor U13918 (N_13918,N_10128,N_11553);
xnor U13919 (N_13919,N_10316,N_10847);
nor U13920 (N_13920,N_11074,N_9940);
nand U13921 (N_13921,N_11576,N_11756);
and U13922 (N_13922,N_9315,N_11704);
and U13923 (N_13923,N_10202,N_9635);
or U13924 (N_13924,N_11300,N_9466);
and U13925 (N_13925,N_9502,N_11067);
nand U13926 (N_13926,N_9778,N_11170);
and U13927 (N_13927,N_9156,N_9807);
xor U13928 (N_13928,N_9180,N_11612);
xnor U13929 (N_13929,N_11847,N_9170);
nand U13930 (N_13930,N_10396,N_11359);
and U13931 (N_13931,N_10066,N_11711);
xor U13932 (N_13932,N_9710,N_10813);
and U13933 (N_13933,N_10458,N_9538);
nor U13934 (N_13934,N_10170,N_9150);
nand U13935 (N_13935,N_11871,N_11822);
nand U13936 (N_13936,N_9254,N_11033);
nor U13937 (N_13937,N_10423,N_10264);
xnor U13938 (N_13938,N_11536,N_9703);
xor U13939 (N_13939,N_10915,N_9690);
nand U13940 (N_13940,N_9778,N_9274);
nand U13941 (N_13941,N_10349,N_10858);
nor U13942 (N_13942,N_9242,N_10864);
nor U13943 (N_13943,N_10455,N_10101);
nand U13944 (N_13944,N_9761,N_10476);
or U13945 (N_13945,N_11333,N_10774);
xor U13946 (N_13946,N_11268,N_9298);
xnor U13947 (N_13947,N_9904,N_10430);
nand U13948 (N_13948,N_11542,N_10084);
nand U13949 (N_13949,N_9717,N_10791);
and U13950 (N_13950,N_10472,N_10547);
and U13951 (N_13951,N_11647,N_11067);
nand U13952 (N_13952,N_10777,N_10913);
nor U13953 (N_13953,N_10730,N_11919);
nor U13954 (N_13954,N_10561,N_9273);
xor U13955 (N_13955,N_11928,N_9967);
and U13956 (N_13956,N_10473,N_9918);
nor U13957 (N_13957,N_9889,N_9682);
nand U13958 (N_13958,N_9364,N_9383);
or U13959 (N_13959,N_11637,N_9157);
xor U13960 (N_13960,N_11080,N_11802);
and U13961 (N_13961,N_11293,N_10060);
or U13962 (N_13962,N_10000,N_10295);
nor U13963 (N_13963,N_10639,N_11491);
xnor U13964 (N_13964,N_9761,N_11469);
and U13965 (N_13965,N_11694,N_10568);
nor U13966 (N_13966,N_10923,N_10677);
nor U13967 (N_13967,N_10796,N_11412);
and U13968 (N_13968,N_11890,N_9786);
and U13969 (N_13969,N_9318,N_11614);
and U13970 (N_13970,N_11355,N_11174);
nand U13971 (N_13971,N_10286,N_10766);
nand U13972 (N_13972,N_9908,N_9347);
nor U13973 (N_13973,N_10541,N_9772);
or U13974 (N_13974,N_10559,N_11965);
and U13975 (N_13975,N_9181,N_9535);
nand U13976 (N_13976,N_11150,N_9824);
xor U13977 (N_13977,N_9170,N_9757);
xnor U13978 (N_13978,N_11351,N_11902);
xnor U13979 (N_13979,N_9551,N_9096);
nor U13980 (N_13980,N_9589,N_9529);
or U13981 (N_13981,N_10062,N_9422);
or U13982 (N_13982,N_9154,N_11305);
nand U13983 (N_13983,N_9553,N_11772);
nor U13984 (N_13984,N_10909,N_11255);
nand U13985 (N_13985,N_10120,N_10570);
xnor U13986 (N_13986,N_10659,N_10314);
nand U13987 (N_13987,N_9859,N_9035);
nand U13988 (N_13988,N_11051,N_11521);
nand U13989 (N_13989,N_10499,N_9544);
and U13990 (N_13990,N_11162,N_9445);
nand U13991 (N_13991,N_10038,N_10599);
and U13992 (N_13992,N_10233,N_9208);
or U13993 (N_13993,N_10652,N_10227);
and U13994 (N_13994,N_11235,N_9319);
xor U13995 (N_13995,N_11493,N_10721);
xor U13996 (N_13996,N_9114,N_10825);
nor U13997 (N_13997,N_10238,N_10273);
and U13998 (N_13998,N_9956,N_9923);
nor U13999 (N_13999,N_11715,N_11353);
and U14000 (N_14000,N_9271,N_9028);
and U14001 (N_14001,N_11720,N_10322);
nand U14002 (N_14002,N_10429,N_10698);
and U14003 (N_14003,N_10405,N_11820);
nand U14004 (N_14004,N_10111,N_9825);
nor U14005 (N_14005,N_11575,N_9473);
xnor U14006 (N_14006,N_11593,N_10139);
or U14007 (N_14007,N_11851,N_9099);
nor U14008 (N_14008,N_10426,N_9079);
nor U14009 (N_14009,N_11828,N_11358);
nand U14010 (N_14010,N_11039,N_9348);
or U14011 (N_14011,N_10932,N_11832);
nand U14012 (N_14012,N_11675,N_11112);
xor U14013 (N_14013,N_10304,N_9760);
and U14014 (N_14014,N_9711,N_9720);
or U14015 (N_14015,N_9681,N_10064);
and U14016 (N_14016,N_9169,N_10652);
nand U14017 (N_14017,N_9317,N_10277);
or U14018 (N_14018,N_10095,N_11986);
or U14019 (N_14019,N_10160,N_9775);
nor U14020 (N_14020,N_11817,N_9007);
and U14021 (N_14021,N_9672,N_11975);
or U14022 (N_14022,N_11403,N_9065);
or U14023 (N_14023,N_11830,N_11775);
and U14024 (N_14024,N_11708,N_11506);
nor U14025 (N_14025,N_10906,N_10116);
and U14026 (N_14026,N_9770,N_10306);
xnor U14027 (N_14027,N_9012,N_11044);
xor U14028 (N_14028,N_10724,N_9548);
nor U14029 (N_14029,N_10140,N_11447);
xor U14030 (N_14030,N_11840,N_11566);
or U14031 (N_14031,N_10633,N_11665);
and U14032 (N_14032,N_11925,N_9772);
nor U14033 (N_14033,N_10188,N_9593);
or U14034 (N_14034,N_10705,N_9894);
nand U14035 (N_14035,N_9599,N_10318);
nand U14036 (N_14036,N_10332,N_10682);
nand U14037 (N_14037,N_9132,N_9515);
nor U14038 (N_14038,N_10616,N_9360);
and U14039 (N_14039,N_11540,N_9802);
nor U14040 (N_14040,N_11038,N_9202);
nand U14041 (N_14041,N_9258,N_11491);
nor U14042 (N_14042,N_10762,N_10551);
nor U14043 (N_14043,N_10221,N_9863);
nand U14044 (N_14044,N_11269,N_9606);
or U14045 (N_14045,N_11614,N_9509);
xor U14046 (N_14046,N_10775,N_9528);
xor U14047 (N_14047,N_9434,N_11634);
and U14048 (N_14048,N_9781,N_11956);
nor U14049 (N_14049,N_11296,N_11971);
or U14050 (N_14050,N_10091,N_9860);
nor U14051 (N_14051,N_9416,N_10770);
xnor U14052 (N_14052,N_10243,N_11552);
or U14053 (N_14053,N_10519,N_10042);
and U14054 (N_14054,N_9576,N_11463);
and U14055 (N_14055,N_11498,N_11732);
nor U14056 (N_14056,N_10431,N_9817);
and U14057 (N_14057,N_11936,N_10311);
nor U14058 (N_14058,N_9251,N_9788);
xor U14059 (N_14059,N_9864,N_10870);
nor U14060 (N_14060,N_11188,N_11997);
nand U14061 (N_14061,N_9170,N_10436);
xor U14062 (N_14062,N_10487,N_9081);
nor U14063 (N_14063,N_10734,N_9395);
nor U14064 (N_14064,N_9792,N_10387);
nand U14065 (N_14065,N_10899,N_9353);
and U14066 (N_14066,N_10413,N_11572);
nor U14067 (N_14067,N_9128,N_11299);
and U14068 (N_14068,N_10114,N_11292);
nand U14069 (N_14069,N_10273,N_10574);
and U14070 (N_14070,N_10995,N_11935);
xnor U14071 (N_14071,N_9868,N_10267);
and U14072 (N_14072,N_10628,N_10315);
nor U14073 (N_14073,N_10993,N_9967);
xnor U14074 (N_14074,N_9461,N_10952);
nand U14075 (N_14075,N_11616,N_9286);
nor U14076 (N_14076,N_11169,N_10257);
and U14077 (N_14077,N_10284,N_9706);
xnor U14078 (N_14078,N_10918,N_9275);
nor U14079 (N_14079,N_9931,N_9586);
xnor U14080 (N_14080,N_10107,N_9447);
or U14081 (N_14081,N_10461,N_10258);
and U14082 (N_14082,N_11956,N_9670);
nor U14083 (N_14083,N_10940,N_9652);
nand U14084 (N_14084,N_10680,N_11423);
or U14085 (N_14085,N_9149,N_10580);
xnor U14086 (N_14086,N_9176,N_10692);
or U14087 (N_14087,N_10920,N_10812);
nand U14088 (N_14088,N_11281,N_10253);
nor U14089 (N_14089,N_9297,N_11389);
nor U14090 (N_14090,N_9048,N_9921);
nand U14091 (N_14091,N_9523,N_9904);
nand U14092 (N_14092,N_10081,N_10441);
xor U14093 (N_14093,N_9598,N_10623);
and U14094 (N_14094,N_11481,N_11237);
or U14095 (N_14095,N_9906,N_9889);
or U14096 (N_14096,N_10162,N_9794);
and U14097 (N_14097,N_9309,N_10769);
and U14098 (N_14098,N_9925,N_9379);
nand U14099 (N_14099,N_11301,N_9699);
nand U14100 (N_14100,N_10006,N_10409);
and U14101 (N_14101,N_10745,N_10983);
xor U14102 (N_14102,N_11377,N_10112);
or U14103 (N_14103,N_10416,N_9584);
or U14104 (N_14104,N_11048,N_11747);
nand U14105 (N_14105,N_10302,N_11833);
and U14106 (N_14106,N_11948,N_11077);
or U14107 (N_14107,N_9671,N_10534);
nand U14108 (N_14108,N_11641,N_10062);
or U14109 (N_14109,N_9884,N_9684);
nor U14110 (N_14110,N_11806,N_11735);
nand U14111 (N_14111,N_11632,N_9934);
or U14112 (N_14112,N_9127,N_11770);
nor U14113 (N_14113,N_9398,N_11955);
and U14114 (N_14114,N_9698,N_9147);
nand U14115 (N_14115,N_9475,N_9260);
nor U14116 (N_14116,N_11773,N_11192);
xor U14117 (N_14117,N_11000,N_11065);
or U14118 (N_14118,N_9355,N_10011);
or U14119 (N_14119,N_9951,N_10497);
and U14120 (N_14120,N_11462,N_9978);
xnor U14121 (N_14121,N_10174,N_10213);
or U14122 (N_14122,N_9096,N_10181);
or U14123 (N_14123,N_11773,N_9649);
xnor U14124 (N_14124,N_10634,N_11393);
nor U14125 (N_14125,N_9949,N_9561);
nor U14126 (N_14126,N_10115,N_11432);
or U14127 (N_14127,N_10682,N_11372);
and U14128 (N_14128,N_10381,N_9931);
nor U14129 (N_14129,N_10235,N_10712);
xor U14130 (N_14130,N_9928,N_10039);
nor U14131 (N_14131,N_11696,N_10032);
nor U14132 (N_14132,N_10658,N_9602);
nor U14133 (N_14133,N_9819,N_9395);
nor U14134 (N_14134,N_10297,N_10983);
xor U14135 (N_14135,N_10210,N_9941);
and U14136 (N_14136,N_9937,N_11944);
and U14137 (N_14137,N_10211,N_10517);
and U14138 (N_14138,N_10568,N_11283);
nand U14139 (N_14139,N_11357,N_11904);
or U14140 (N_14140,N_10399,N_11950);
nand U14141 (N_14141,N_10043,N_9582);
nand U14142 (N_14142,N_9045,N_11696);
nand U14143 (N_14143,N_10204,N_10427);
nand U14144 (N_14144,N_11612,N_11448);
nand U14145 (N_14145,N_11519,N_11736);
nand U14146 (N_14146,N_11049,N_9731);
and U14147 (N_14147,N_10769,N_11198);
nand U14148 (N_14148,N_10502,N_10783);
and U14149 (N_14149,N_9398,N_11234);
xor U14150 (N_14150,N_11244,N_9598);
or U14151 (N_14151,N_9721,N_9360);
xnor U14152 (N_14152,N_9664,N_11299);
xor U14153 (N_14153,N_9916,N_11295);
xor U14154 (N_14154,N_9521,N_9378);
or U14155 (N_14155,N_9644,N_11343);
and U14156 (N_14156,N_11697,N_9588);
and U14157 (N_14157,N_9471,N_10459);
or U14158 (N_14158,N_11471,N_10690);
nor U14159 (N_14159,N_10330,N_10798);
nor U14160 (N_14160,N_10803,N_10439);
nor U14161 (N_14161,N_11352,N_9862);
and U14162 (N_14162,N_10233,N_11078);
nand U14163 (N_14163,N_9529,N_11500);
xnor U14164 (N_14164,N_9526,N_9132);
nor U14165 (N_14165,N_10311,N_11420);
nor U14166 (N_14166,N_11464,N_10919);
and U14167 (N_14167,N_10844,N_9989);
or U14168 (N_14168,N_11421,N_9784);
nand U14169 (N_14169,N_11109,N_11056);
or U14170 (N_14170,N_11564,N_11025);
or U14171 (N_14171,N_10898,N_10728);
nand U14172 (N_14172,N_11290,N_11267);
nor U14173 (N_14173,N_9493,N_10817);
xnor U14174 (N_14174,N_11480,N_9727);
or U14175 (N_14175,N_9391,N_9302);
or U14176 (N_14176,N_9959,N_9819);
or U14177 (N_14177,N_9348,N_9845);
xnor U14178 (N_14178,N_9980,N_10737);
nand U14179 (N_14179,N_10749,N_10175);
nor U14180 (N_14180,N_11956,N_9672);
nor U14181 (N_14181,N_9091,N_10920);
and U14182 (N_14182,N_10068,N_9987);
and U14183 (N_14183,N_10632,N_11412);
or U14184 (N_14184,N_9377,N_9530);
nand U14185 (N_14185,N_9873,N_9692);
xnor U14186 (N_14186,N_11354,N_9806);
nor U14187 (N_14187,N_9886,N_10750);
and U14188 (N_14188,N_9461,N_10191);
nand U14189 (N_14189,N_11551,N_9412);
xor U14190 (N_14190,N_9795,N_9867);
xnor U14191 (N_14191,N_10686,N_11142);
xnor U14192 (N_14192,N_10723,N_10698);
xor U14193 (N_14193,N_9563,N_11132);
and U14194 (N_14194,N_11772,N_11866);
nor U14195 (N_14195,N_10056,N_9406);
nand U14196 (N_14196,N_10988,N_11266);
and U14197 (N_14197,N_10412,N_9250);
and U14198 (N_14198,N_10093,N_11934);
xnor U14199 (N_14199,N_9616,N_11072);
nand U14200 (N_14200,N_11915,N_11188);
or U14201 (N_14201,N_11669,N_9143);
xor U14202 (N_14202,N_9923,N_11350);
or U14203 (N_14203,N_10871,N_9634);
and U14204 (N_14204,N_11221,N_11236);
xor U14205 (N_14205,N_9144,N_11936);
and U14206 (N_14206,N_9263,N_11222);
nor U14207 (N_14207,N_10135,N_11992);
or U14208 (N_14208,N_9073,N_9238);
or U14209 (N_14209,N_10098,N_11089);
xnor U14210 (N_14210,N_11227,N_10786);
nor U14211 (N_14211,N_10389,N_11321);
and U14212 (N_14212,N_9613,N_11746);
nand U14213 (N_14213,N_9983,N_11723);
or U14214 (N_14214,N_9001,N_11388);
nor U14215 (N_14215,N_10663,N_11238);
nand U14216 (N_14216,N_11894,N_10114);
xnor U14217 (N_14217,N_11477,N_9435);
and U14218 (N_14218,N_9684,N_10336);
or U14219 (N_14219,N_9613,N_11821);
nand U14220 (N_14220,N_9895,N_10985);
xor U14221 (N_14221,N_10346,N_9956);
or U14222 (N_14222,N_11077,N_11494);
or U14223 (N_14223,N_10851,N_9026);
nand U14224 (N_14224,N_11625,N_11331);
nor U14225 (N_14225,N_10200,N_11768);
xnor U14226 (N_14226,N_10364,N_9741);
nor U14227 (N_14227,N_9155,N_11558);
and U14228 (N_14228,N_9762,N_9319);
nor U14229 (N_14229,N_10673,N_9644);
and U14230 (N_14230,N_11941,N_9642);
or U14231 (N_14231,N_11157,N_10452);
and U14232 (N_14232,N_10546,N_10882);
or U14233 (N_14233,N_11672,N_11836);
or U14234 (N_14234,N_9223,N_11689);
nor U14235 (N_14235,N_11909,N_11223);
xor U14236 (N_14236,N_11109,N_11031);
nor U14237 (N_14237,N_9463,N_9917);
xor U14238 (N_14238,N_9112,N_9415);
and U14239 (N_14239,N_11355,N_10899);
nor U14240 (N_14240,N_11056,N_10337);
or U14241 (N_14241,N_10328,N_10006);
and U14242 (N_14242,N_9907,N_9065);
nand U14243 (N_14243,N_11186,N_10945);
nand U14244 (N_14244,N_9625,N_11020);
nor U14245 (N_14245,N_9267,N_9555);
nor U14246 (N_14246,N_9906,N_11025);
nor U14247 (N_14247,N_10058,N_11593);
and U14248 (N_14248,N_10507,N_11973);
nand U14249 (N_14249,N_10201,N_9866);
xor U14250 (N_14250,N_10066,N_11588);
or U14251 (N_14251,N_10880,N_10320);
or U14252 (N_14252,N_9300,N_10060);
xnor U14253 (N_14253,N_11988,N_10336);
xor U14254 (N_14254,N_11534,N_11994);
and U14255 (N_14255,N_10145,N_11009);
xor U14256 (N_14256,N_10127,N_11671);
xnor U14257 (N_14257,N_11333,N_11604);
nand U14258 (N_14258,N_10160,N_10633);
nor U14259 (N_14259,N_10577,N_10107);
and U14260 (N_14260,N_11436,N_11899);
or U14261 (N_14261,N_11138,N_10122);
nand U14262 (N_14262,N_10020,N_10273);
nor U14263 (N_14263,N_10883,N_9317);
nand U14264 (N_14264,N_9465,N_11180);
xnor U14265 (N_14265,N_9737,N_9871);
nand U14266 (N_14266,N_9314,N_11141);
and U14267 (N_14267,N_11955,N_10490);
and U14268 (N_14268,N_10240,N_10572);
nand U14269 (N_14269,N_11342,N_9816);
nor U14270 (N_14270,N_9956,N_9027);
nor U14271 (N_14271,N_11824,N_11097);
and U14272 (N_14272,N_11799,N_9080);
or U14273 (N_14273,N_10051,N_10871);
nor U14274 (N_14274,N_10220,N_9408);
or U14275 (N_14275,N_10499,N_11703);
or U14276 (N_14276,N_9946,N_10721);
xor U14277 (N_14277,N_11609,N_9604);
nor U14278 (N_14278,N_10724,N_11056);
nor U14279 (N_14279,N_10272,N_9350);
nand U14280 (N_14280,N_11357,N_9405);
xor U14281 (N_14281,N_9548,N_9885);
nand U14282 (N_14282,N_11728,N_11619);
or U14283 (N_14283,N_10188,N_11659);
or U14284 (N_14284,N_9537,N_10037);
nor U14285 (N_14285,N_11961,N_11793);
nor U14286 (N_14286,N_9779,N_10462);
xnor U14287 (N_14287,N_10692,N_10979);
and U14288 (N_14288,N_10027,N_9380);
xor U14289 (N_14289,N_10554,N_11766);
or U14290 (N_14290,N_10658,N_11044);
xnor U14291 (N_14291,N_9710,N_11961);
or U14292 (N_14292,N_9860,N_9725);
nand U14293 (N_14293,N_10405,N_11021);
and U14294 (N_14294,N_10779,N_9843);
or U14295 (N_14295,N_11390,N_9841);
nand U14296 (N_14296,N_11518,N_9642);
or U14297 (N_14297,N_11206,N_10428);
or U14298 (N_14298,N_10371,N_9652);
nor U14299 (N_14299,N_11631,N_10758);
xnor U14300 (N_14300,N_10289,N_9632);
nor U14301 (N_14301,N_9362,N_11264);
nand U14302 (N_14302,N_10239,N_10830);
xnor U14303 (N_14303,N_10009,N_9897);
or U14304 (N_14304,N_11270,N_9107);
and U14305 (N_14305,N_11486,N_10305);
nor U14306 (N_14306,N_9306,N_9030);
nor U14307 (N_14307,N_10628,N_10375);
xnor U14308 (N_14308,N_11885,N_10098);
nor U14309 (N_14309,N_11132,N_11003);
xnor U14310 (N_14310,N_10042,N_10617);
or U14311 (N_14311,N_10049,N_11688);
and U14312 (N_14312,N_10033,N_9458);
nand U14313 (N_14313,N_11087,N_11780);
nand U14314 (N_14314,N_11298,N_11381);
nor U14315 (N_14315,N_11833,N_11904);
xor U14316 (N_14316,N_10724,N_9075);
and U14317 (N_14317,N_9416,N_10015);
nor U14318 (N_14318,N_10397,N_11142);
nand U14319 (N_14319,N_10766,N_9929);
xnor U14320 (N_14320,N_9891,N_9623);
nor U14321 (N_14321,N_9134,N_10116);
nor U14322 (N_14322,N_11215,N_11613);
xor U14323 (N_14323,N_10845,N_11114);
or U14324 (N_14324,N_11865,N_10015);
nand U14325 (N_14325,N_9604,N_10954);
and U14326 (N_14326,N_10011,N_10446);
nor U14327 (N_14327,N_10716,N_11595);
xor U14328 (N_14328,N_10383,N_9834);
nand U14329 (N_14329,N_11351,N_11740);
nor U14330 (N_14330,N_9059,N_11028);
xor U14331 (N_14331,N_11291,N_9858);
or U14332 (N_14332,N_11074,N_9109);
xnor U14333 (N_14333,N_10593,N_9994);
nor U14334 (N_14334,N_10409,N_9273);
xor U14335 (N_14335,N_9311,N_9871);
or U14336 (N_14336,N_10332,N_10055);
or U14337 (N_14337,N_9082,N_10945);
and U14338 (N_14338,N_10301,N_10634);
and U14339 (N_14339,N_10487,N_11501);
nand U14340 (N_14340,N_11823,N_11921);
xor U14341 (N_14341,N_11251,N_9802);
and U14342 (N_14342,N_11150,N_9733);
and U14343 (N_14343,N_11251,N_10638);
nand U14344 (N_14344,N_9099,N_9854);
xor U14345 (N_14345,N_9677,N_9066);
xnor U14346 (N_14346,N_10160,N_11177);
nor U14347 (N_14347,N_11020,N_11969);
nand U14348 (N_14348,N_9701,N_9276);
xnor U14349 (N_14349,N_9162,N_9924);
or U14350 (N_14350,N_11377,N_9165);
xor U14351 (N_14351,N_11540,N_10933);
nor U14352 (N_14352,N_11266,N_11599);
xor U14353 (N_14353,N_9005,N_10622);
nand U14354 (N_14354,N_11774,N_10447);
or U14355 (N_14355,N_9243,N_9727);
nor U14356 (N_14356,N_10648,N_9597);
nand U14357 (N_14357,N_9539,N_11433);
or U14358 (N_14358,N_9757,N_11047);
nor U14359 (N_14359,N_11936,N_10170);
nand U14360 (N_14360,N_9379,N_9481);
xnor U14361 (N_14361,N_9715,N_10728);
or U14362 (N_14362,N_11226,N_9756);
or U14363 (N_14363,N_9494,N_11990);
nand U14364 (N_14364,N_11436,N_11807);
nor U14365 (N_14365,N_10189,N_11486);
nor U14366 (N_14366,N_10246,N_11001);
and U14367 (N_14367,N_10146,N_11028);
nor U14368 (N_14368,N_9863,N_11501);
nand U14369 (N_14369,N_9518,N_11649);
or U14370 (N_14370,N_11347,N_10116);
and U14371 (N_14371,N_10542,N_11102);
or U14372 (N_14372,N_9593,N_10977);
or U14373 (N_14373,N_11828,N_9509);
xnor U14374 (N_14374,N_9003,N_11874);
xnor U14375 (N_14375,N_11670,N_9431);
nand U14376 (N_14376,N_9897,N_9402);
nor U14377 (N_14377,N_10939,N_10928);
and U14378 (N_14378,N_10488,N_11369);
xnor U14379 (N_14379,N_10926,N_10895);
xnor U14380 (N_14380,N_11601,N_9990);
or U14381 (N_14381,N_10426,N_11088);
nor U14382 (N_14382,N_9840,N_11141);
nor U14383 (N_14383,N_10441,N_10930);
xor U14384 (N_14384,N_9147,N_11526);
and U14385 (N_14385,N_11517,N_10856);
xnor U14386 (N_14386,N_9794,N_11033);
or U14387 (N_14387,N_11264,N_9776);
and U14388 (N_14388,N_10190,N_10577);
xor U14389 (N_14389,N_11791,N_11824);
xor U14390 (N_14390,N_10926,N_9507);
nor U14391 (N_14391,N_11810,N_9883);
xor U14392 (N_14392,N_9751,N_9848);
and U14393 (N_14393,N_11392,N_10501);
and U14394 (N_14394,N_10653,N_10470);
nand U14395 (N_14395,N_10139,N_10483);
nand U14396 (N_14396,N_11494,N_9128);
nor U14397 (N_14397,N_11595,N_9159);
xnor U14398 (N_14398,N_9457,N_11918);
xnor U14399 (N_14399,N_9260,N_11536);
nand U14400 (N_14400,N_9509,N_9229);
or U14401 (N_14401,N_9918,N_10578);
or U14402 (N_14402,N_11615,N_11952);
or U14403 (N_14403,N_9490,N_11975);
or U14404 (N_14404,N_9667,N_10995);
xor U14405 (N_14405,N_9214,N_10815);
nor U14406 (N_14406,N_9810,N_11711);
nor U14407 (N_14407,N_9781,N_11828);
nand U14408 (N_14408,N_10701,N_9739);
nor U14409 (N_14409,N_9701,N_11008);
nand U14410 (N_14410,N_9769,N_10436);
nand U14411 (N_14411,N_9560,N_11515);
nor U14412 (N_14412,N_10174,N_9046);
and U14413 (N_14413,N_10044,N_10623);
or U14414 (N_14414,N_11593,N_10714);
nand U14415 (N_14415,N_11324,N_11123);
nor U14416 (N_14416,N_9325,N_10126);
nand U14417 (N_14417,N_11123,N_11161);
and U14418 (N_14418,N_11381,N_10667);
or U14419 (N_14419,N_11915,N_11456);
or U14420 (N_14420,N_9867,N_9919);
nor U14421 (N_14421,N_10443,N_11301);
and U14422 (N_14422,N_9408,N_10110);
nand U14423 (N_14423,N_11884,N_9519);
nand U14424 (N_14424,N_10890,N_10068);
nand U14425 (N_14425,N_11102,N_9307);
nor U14426 (N_14426,N_10692,N_11171);
nor U14427 (N_14427,N_11439,N_11274);
or U14428 (N_14428,N_10965,N_10628);
and U14429 (N_14429,N_9051,N_11394);
and U14430 (N_14430,N_11763,N_11442);
nand U14431 (N_14431,N_10927,N_9381);
and U14432 (N_14432,N_9213,N_9062);
nor U14433 (N_14433,N_11932,N_9386);
and U14434 (N_14434,N_10701,N_9201);
nor U14435 (N_14435,N_11855,N_11622);
nand U14436 (N_14436,N_10918,N_9234);
nand U14437 (N_14437,N_9307,N_11895);
or U14438 (N_14438,N_10001,N_10860);
nand U14439 (N_14439,N_11311,N_10884);
xor U14440 (N_14440,N_10872,N_9829);
nand U14441 (N_14441,N_11237,N_9344);
and U14442 (N_14442,N_9573,N_9792);
nor U14443 (N_14443,N_10097,N_10999);
nand U14444 (N_14444,N_11464,N_11153);
nor U14445 (N_14445,N_9558,N_9848);
nand U14446 (N_14446,N_11105,N_10104);
nor U14447 (N_14447,N_10380,N_11646);
or U14448 (N_14448,N_9131,N_9677);
or U14449 (N_14449,N_10371,N_9051);
or U14450 (N_14450,N_9632,N_9685);
nand U14451 (N_14451,N_11283,N_11352);
or U14452 (N_14452,N_9117,N_9884);
xnor U14453 (N_14453,N_9714,N_10616);
or U14454 (N_14454,N_10620,N_9370);
nor U14455 (N_14455,N_11667,N_9056);
nand U14456 (N_14456,N_10714,N_11838);
nor U14457 (N_14457,N_9191,N_10841);
nand U14458 (N_14458,N_10055,N_10761);
and U14459 (N_14459,N_9795,N_11170);
and U14460 (N_14460,N_11513,N_11595);
xnor U14461 (N_14461,N_11272,N_11349);
nor U14462 (N_14462,N_10394,N_10632);
or U14463 (N_14463,N_10389,N_11450);
nor U14464 (N_14464,N_10044,N_9829);
or U14465 (N_14465,N_9113,N_11829);
xnor U14466 (N_14466,N_11823,N_9137);
and U14467 (N_14467,N_10036,N_11170);
xor U14468 (N_14468,N_9541,N_11168);
and U14469 (N_14469,N_11686,N_11419);
nand U14470 (N_14470,N_10617,N_9198);
xor U14471 (N_14471,N_9532,N_9667);
and U14472 (N_14472,N_10374,N_10454);
nand U14473 (N_14473,N_10380,N_10692);
nand U14474 (N_14474,N_11956,N_10055);
xnor U14475 (N_14475,N_11253,N_10174);
nand U14476 (N_14476,N_11118,N_10770);
nor U14477 (N_14477,N_10997,N_10437);
xnor U14478 (N_14478,N_11333,N_9037);
nand U14479 (N_14479,N_11920,N_11160);
nand U14480 (N_14480,N_9557,N_10699);
xor U14481 (N_14481,N_10890,N_11328);
nand U14482 (N_14482,N_11380,N_9593);
or U14483 (N_14483,N_10353,N_9878);
xnor U14484 (N_14484,N_10887,N_10503);
nand U14485 (N_14485,N_9369,N_9825);
xor U14486 (N_14486,N_10851,N_10394);
xor U14487 (N_14487,N_10980,N_9664);
and U14488 (N_14488,N_10735,N_10021);
nand U14489 (N_14489,N_11822,N_10877);
nand U14490 (N_14490,N_10049,N_11292);
nand U14491 (N_14491,N_10873,N_11357);
and U14492 (N_14492,N_11293,N_9862);
nor U14493 (N_14493,N_11325,N_11750);
or U14494 (N_14494,N_10423,N_9305);
xor U14495 (N_14495,N_11622,N_9304);
nor U14496 (N_14496,N_10203,N_10616);
nor U14497 (N_14497,N_11519,N_10807);
xnor U14498 (N_14498,N_10210,N_9479);
or U14499 (N_14499,N_11259,N_9596);
nor U14500 (N_14500,N_9617,N_9400);
nand U14501 (N_14501,N_10692,N_9401);
nor U14502 (N_14502,N_9942,N_9204);
nand U14503 (N_14503,N_9896,N_9965);
xnor U14504 (N_14504,N_10192,N_10955);
or U14505 (N_14505,N_9200,N_11446);
nor U14506 (N_14506,N_9018,N_9469);
or U14507 (N_14507,N_11939,N_9777);
or U14508 (N_14508,N_11183,N_10619);
xor U14509 (N_14509,N_11183,N_11854);
nor U14510 (N_14510,N_9545,N_9254);
nand U14511 (N_14511,N_9360,N_9686);
xor U14512 (N_14512,N_9467,N_11331);
xnor U14513 (N_14513,N_10237,N_10558);
xnor U14514 (N_14514,N_10202,N_10883);
and U14515 (N_14515,N_10723,N_10000);
xnor U14516 (N_14516,N_10464,N_9618);
or U14517 (N_14517,N_9110,N_10541);
or U14518 (N_14518,N_9279,N_10246);
nor U14519 (N_14519,N_10944,N_9716);
nor U14520 (N_14520,N_11910,N_9621);
nand U14521 (N_14521,N_11247,N_9429);
and U14522 (N_14522,N_9949,N_9324);
xor U14523 (N_14523,N_9954,N_11374);
xor U14524 (N_14524,N_10659,N_11142);
and U14525 (N_14525,N_10252,N_9906);
xnor U14526 (N_14526,N_10479,N_10559);
nor U14527 (N_14527,N_10529,N_11844);
or U14528 (N_14528,N_10108,N_9439);
and U14529 (N_14529,N_9111,N_9457);
nand U14530 (N_14530,N_11124,N_10151);
xnor U14531 (N_14531,N_10237,N_11452);
nand U14532 (N_14532,N_10387,N_10752);
nor U14533 (N_14533,N_9949,N_10481);
nand U14534 (N_14534,N_10198,N_10840);
and U14535 (N_14535,N_10194,N_9913);
and U14536 (N_14536,N_9144,N_9480);
or U14537 (N_14537,N_9305,N_11374);
xnor U14538 (N_14538,N_11236,N_10174);
or U14539 (N_14539,N_9749,N_9374);
and U14540 (N_14540,N_9042,N_9500);
nand U14541 (N_14541,N_11764,N_10791);
or U14542 (N_14542,N_9906,N_10616);
or U14543 (N_14543,N_9142,N_11092);
and U14544 (N_14544,N_9177,N_10855);
xor U14545 (N_14545,N_10471,N_10816);
or U14546 (N_14546,N_11086,N_10493);
nor U14547 (N_14547,N_9779,N_11703);
nor U14548 (N_14548,N_11442,N_9586);
nor U14549 (N_14549,N_10318,N_11210);
or U14550 (N_14550,N_9140,N_9704);
nand U14551 (N_14551,N_10950,N_11550);
nor U14552 (N_14552,N_10588,N_11928);
xnor U14553 (N_14553,N_11478,N_11155);
and U14554 (N_14554,N_11388,N_9755);
xnor U14555 (N_14555,N_11232,N_10843);
nand U14556 (N_14556,N_9373,N_10745);
or U14557 (N_14557,N_11110,N_11881);
or U14558 (N_14558,N_9592,N_11655);
xor U14559 (N_14559,N_10862,N_9204);
nand U14560 (N_14560,N_11930,N_11952);
nor U14561 (N_14561,N_10351,N_10101);
nand U14562 (N_14562,N_9409,N_10778);
nor U14563 (N_14563,N_11080,N_10958);
nor U14564 (N_14564,N_10271,N_10085);
and U14565 (N_14565,N_11695,N_10791);
nor U14566 (N_14566,N_9588,N_10699);
nand U14567 (N_14567,N_10570,N_10321);
xor U14568 (N_14568,N_11189,N_10675);
and U14569 (N_14569,N_11095,N_10242);
or U14570 (N_14570,N_9799,N_11976);
and U14571 (N_14571,N_10321,N_9753);
xor U14572 (N_14572,N_11389,N_9428);
nor U14573 (N_14573,N_11873,N_11632);
nor U14574 (N_14574,N_10612,N_11667);
xnor U14575 (N_14575,N_9912,N_11084);
nand U14576 (N_14576,N_9826,N_10184);
or U14577 (N_14577,N_11416,N_11647);
or U14578 (N_14578,N_9695,N_10440);
and U14579 (N_14579,N_10144,N_9263);
or U14580 (N_14580,N_11381,N_9736);
and U14581 (N_14581,N_9937,N_11349);
nor U14582 (N_14582,N_10184,N_10576);
xnor U14583 (N_14583,N_11403,N_9389);
nor U14584 (N_14584,N_11421,N_10653);
xor U14585 (N_14585,N_9737,N_11160);
or U14586 (N_14586,N_11935,N_11258);
or U14587 (N_14587,N_11529,N_11646);
or U14588 (N_14588,N_11228,N_11479);
nor U14589 (N_14589,N_9306,N_10732);
nand U14590 (N_14590,N_11252,N_9473);
xnor U14591 (N_14591,N_9842,N_10543);
xor U14592 (N_14592,N_9867,N_9074);
nor U14593 (N_14593,N_9075,N_9345);
and U14594 (N_14594,N_10389,N_10597);
nor U14595 (N_14595,N_9323,N_11961);
xor U14596 (N_14596,N_10428,N_11333);
and U14597 (N_14597,N_11299,N_9707);
or U14598 (N_14598,N_10970,N_10115);
nor U14599 (N_14599,N_11820,N_10325);
nand U14600 (N_14600,N_10230,N_10502);
nand U14601 (N_14601,N_10999,N_11416);
nand U14602 (N_14602,N_11529,N_11086);
and U14603 (N_14603,N_9010,N_11027);
nand U14604 (N_14604,N_10921,N_9054);
nand U14605 (N_14605,N_10247,N_11895);
xor U14606 (N_14606,N_10592,N_9213);
and U14607 (N_14607,N_9112,N_11828);
xnor U14608 (N_14608,N_10039,N_11488);
nand U14609 (N_14609,N_10003,N_11449);
xor U14610 (N_14610,N_10062,N_9625);
xor U14611 (N_14611,N_9915,N_11561);
xnor U14612 (N_14612,N_11932,N_10039);
nand U14613 (N_14613,N_11242,N_10421);
and U14614 (N_14614,N_11602,N_10212);
xnor U14615 (N_14615,N_11858,N_10800);
or U14616 (N_14616,N_10420,N_11308);
xnor U14617 (N_14617,N_10716,N_11948);
or U14618 (N_14618,N_11954,N_11267);
xnor U14619 (N_14619,N_11034,N_10576);
xor U14620 (N_14620,N_10040,N_11179);
nor U14621 (N_14621,N_10485,N_9594);
and U14622 (N_14622,N_11277,N_10373);
nor U14623 (N_14623,N_9495,N_11578);
and U14624 (N_14624,N_9695,N_11365);
nand U14625 (N_14625,N_9979,N_10003);
nand U14626 (N_14626,N_11716,N_9006);
nor U14627 (N_14627,N_11887,N_9525);
and U14628 (N_14628,N_9402,N_9838);
and U14629 (N_14629,N_9451,N_9977);
and U14630 (N_14630,N_10658,N_9269);
or U14631 (N_14631,N_11662,N_9161);
nand U14632 (N_14632,N_10122,N_9209);
and U14633 (N_14633,N_10017,N_10289);
and U14634 (N_14634,N_11607,N_11702);
xor U14635 (N_14635,N_11236,N_11256);
or U14636 (N_14636,N_10139,N_10901);
xor U14637 (N_14637,N_11576,N_10789);
xor U14638 (N_14638,N_9895,N_9605);
xor U14639 (N_14639,N_9456,N_9047);
nor U14640 (N_14640,N_11806,N_9331);
or U14641 (N_14641,N_9251,N_10247);
nand U14642 (N_14642,N_11047,N_9521);
nand U14643 (N_14643,N_10815,N_11909);
nor U14644 (N_14644,N_9155,N_10924);
xnor U14645 (N_14645,N_9554,N_10639);
xnor U14646 (N_14646,N_10066,N_9674);
xnor U14647 (N_14647,N_10802,N_10506);
xnor U14648 (N_14648,N_11540,N_11753);
nand U14649 (N_14649,N_9588,N_10034);
and U14650 (N_14650,N_11164,N_10750);
nor U14651 (N_14651,N_10959,N_10024);
nand U14652 (N_14652,N_9151,N_9909);
xnor U14653 (N_14653,N_10373,N_9827);
xnor U14654 (N_14654,N_9065,N_9275);
xnor U14655 (N_14655,N_10352,N_10453);
xnor U14656 (N_14656,N_9145,N_11901);
xor U14657 (N_14657,N_10484,N_10820);
nand U14658 (N_14658,N_11754,N_10896);
nor U14659 (N_14659,N_11599,N_9825);
nor U14660 (N_14660,N_11713,N_11015);
nand U14661 (N_14661,N_10140,N_11197);
xnor U14662 (N_14662,N_11099,N_9073);
xor U14663 (N_14663,N_10716,N_11082);
nand U14664 (N_14664,N_10876,N_9545);
and U14665 (N_14665,N_9696,N_11568);
and U14666 (N_14666,N_10933,N_11708);
nand U14667 (N_14667,N_10525,N_10484);
and U14668 (N_14668,N_11896,N_10651);
nor U14669 (N_14669,N_9774,N_9752);
xor U14670 (N_14670,N_9278,N_10254);
xor U14671 (N_14671,N_9393,N_9589);
nor U14672 (N_14672,N_10514,N_11205);
nand U14673 (N_14673,N_11990,N_10356);
nor U14674 (N_14674,N_11036,N_9743);
nand U14675 (N_14675,N_9978,N_10481);
or U14676 (N_14676,N_9689,N_11144);
xnor U14677 (N_14677,N_10658,N_9617);
nand U14678 (N_14678,N_9579,N_11424);
or U14679 (N_14679,N_10371,N_10171);
or U14680 (N_14680,N_10286,N_11469);
or U14681 (N_14681,N_10302,N_10570);
nor U14682 (N_14682,N_9607,N_11713);
nor U14683 (N_14683,N_9394,N_10820);
or U14684 (N_14684,N_9929,N_9723);
and U14685 (N_14685,N_11690,N_11691);
or U14686 (N_14686,N_9476,N_9083);
and U14687 (N_14687,N_10643,N_10542);
nor U14688 (N_14688,N_9134,N_9398);
and U14689 (N_14689,N_11999,N_10958);
and U14690 (N_14690,N_10218,N_9286);
or U14691 (N_14691,N_10189,N_10710);
nand U14692 (N_14692,N_9222,N_11426);
nand U14693 (N_14693,N_9666,N_11470);
and U14694 (N_14694,N_10719,N_10386);
nor U14695 (N_14695,N_10921,N_11250);
and U14696 (N_14696,N_9466,N_9791);
and U14697 (N_14697,N_11042,N_11446);
and U14698 (N_14698,N_11851,N_11811);
nor U14699 (N_14699,N_11816,N_11236);
nand U14700 (N_14700,N_9630,N_11210);
nand U14701 (N_14701,N_11464,N_11594);
xor U14702 (N_14702,N_9555,N_10818);
and U14703 (N_14703,N_11864,N_9665);
or U14704 (N_14704,N_9225,N_10161);
nor U14705 (N_14705,N_9412,N_11927);
xnor U14706 (N_14706,N_10776,N_11253);
or U14707 (N_14707,N_9010,N_9420);
nand U14708 (N_14708,N_10988,N_9013);
nand U14709 (N_14709,N_9514,N_11213);
or U14710 (N_14710,N_9640,N_11001);
nand U14711 (N_14711,N_10655,N_10784);
nand U14712 (N_14712,N_10655,N_10063);
and U14713 (N_14713,N_11701,N_11196);
xor U14714 (N_14714,N_10683,N_10019);
and U14715 (N_14715,N_10077,N_11713);
xor U14716 (N_14716,N_10131,N_10816);
nor U14717 (N_14717,N_9171,N_11806);
nand U14718 (N_14718,N_11693,N_11877);
nor U14719 (N_14719,N_11558,N_10342);
xnor U14720 (N_14720,N_10466,N_11719);
or U14721 (N_14721,N_11738,N_11634);
nor U14722 (N_14722,N_10113,N_9721);
nor U14723 (N_14723,N_11910,N_9097);
and U14724 (N_14724,N_9708,N_10913);
nand U14725 (N_14725,N_9110,N_9173);
or U14726 (N_14726,N_11519,N_10904);
or U14727 (N_14727,N_9958,N_10169);
nor U14728 (N_14728,N_10703,N_9981);
xnor U14729 (N_14729,N_10280,N_11710);
xor U14730 (N_14730,N_9708,N_11400);
and U14731 (N_14731,N_10695,N_10217);
nor U14732 (N_14732,N_10749,N_11601);
xor U14733 (N_14733,N_9087,N_9472);
xor U14734 (N_14734,N_11883,N_10538);
or U14735 (N_14735,N_11991,N_11139);
or U14736 (N_14736,N_10771,N_10084);
xnor U14737 (N_14737,N_11073,N_9156);
nor U14738 (N_14738,N_10011,N_10873);
or U14739 (N_14739,N_9677,N_10986);
or U14740 (N_14740,N_11459,N_11252);
xor U14741 (N_14741,N_11679,N_9185);
and U14742 (N_14742,N_9922,N_10730);
nor U14743 (N_14743,N_11503,N_11957);
and U14744 (N_14744,N_9009,N_10010);
nor U14745 (N_14745,N_11483,N_10144);
and U14746 (N_14746,N_9914,N_11660);
nand U14747 (N_14747,N_11735,N_11384);
or U14748 (N_14748,N_9662,N_10335);
nor U14749 (N_14749,N_9429,N_11184);
nor U14750 (N_14750,N_10318,N_9781);
nand U14751 (N_14751,N_11252,N_9466);
nor U14752 (N_14752,N_9600,N_10367);
xor U14753 (N_14753,N_10971,N_10514);
xnor U14754 (N_14754,N_10271,N_11513);
nand U14755 (N_14755,N_10985,N_9566);
nor U14756 (N_14756,N_11592,N_9728);
nor U14757 (N_14757,N_11014,N_10889);
and U14758 (N_14758,N_10559,N_11575);
or U14759 (N_14759,N_9444,N_9198);
nor U14760 (N_14760,N_9786,N_9761);
or U14761 (N_14761,N_10527,N_9231);
or U14762 (N_14762,N_11377,N_10162);
nor U14763 (N_14763,N_9638,N_9336);
and U14764 (N_14764,N_10864,N_9682);
or U14765 (N_14765,N_10909,N_11979);
and U14766 (N_14766,N_11423,N_11597);
or U14767 (N_14767,N_11783,N_9987);
or U14768 (N_14768,N_10733,N_9170);
or U14769 (N_14769,N_10750,N_9489);
or U14770 (N_14770,N_10331,N_11748);
xnor U14771 (N_14771,N_11937,N_10276);
and U14772 (N_14772,N_9494,N_9407);
nand U14773 (N_14773,N_10329,N_10403);
nand U14774 (N_14774,N_11419,N_10839);
xnor U14775 (N_14775,N_9612,N_11722);
or U14776 (N_14776,N_10452,N_9428);
nand U14777 (N_14777,N_10020,N_11159);
nor U14778 (N_14778,N_9975,N_11085);
nor U14779 (N_14779,N_10814,N_11084);
nor U14780 (N_14780,N_10151,N_11114);
or U14781 (N_14781,N_10298,N_10817);
xnor U14782 (N_14782,N_11078,N_11460);
nor U14783 (N_14783,N_11025,N_11921);
and U14784 (N_14784,N_10759,N_11642);
nand U14785 (N_14785,N_10009,N_10133);
or U14786 (N_14786,N_11134,N_10227);
xnor U14787 (N_14787,N_9601,N_10685);
and U14788 (N_14788,N_9647,N_9192);
nor U14789 (N_14789,N_10148,N_11125);
nor U14790 (N_14790,N_9999,N_11794);
nand U14791 (N_14791,N_10526,N_11251);
and U14792 (N_14792,N_9459,N_11909);
or U14793 (N_14793,N_9258,N_10415);
or U14794 (N_14794,N_10307,N_10662);
xor U14795 (N_14795,N_11126,N_10418);
xnor U14796 (N_14796,N_9009,N_9947);
or U14797 (N_14797,N_9417,N_11026);
xor U14798 (N_14798,N_11391,N_11106);
or U14799 (N_14799,N_9217,N_10528);
xor U14800 (N_14800,N_10932,N_9759);
nand U14801 (N_14801,N_10786,N_9283);
nand U14802 (N_14802,N_10634,N_10801);
xnor U14803 (N_14803,N_11346,N_10778);
xnor U14804 (N_14804,N_9517,N_10055);
nor U14805 (N_14805,N_9842,N_9157);
or U14806 (N_14806,N_9941,N_9090);
or U14807 (N_14807,N_11488,N_10327);
nand U14808 (N_14808,N_11711,N_9204);
nand U14809 (N_14809,N_10039,N_11576);
nor U14810 (N_14810,N_10393,N_10461);
xnor U14811 (N_14811,N_10524,N_9852);
nor U14812 (N_14812,N_10243,N_11219);
and U14813 (N_14813,N_11032,N_11822);
or U14814 (N_14814,N_9092,N_9367);
nor U14815 (N_14815,N_10293,N_10158);
and U14816 (N_14816,N_9415,N_9622);
nand U14817 (N_14817,N_11177,N_10427);
xnor U14818 (N_14818,N_10476,N_9604);
xor U14819 (N_14819,N_10137,N_11907);
or U14820 (N_14820,N_11034,N_11820);
or U14821 (N_14821,N_9893,N_11825);
nand U14822 (N_14822,N_11202,N_9237);
or U14823 (N_14823,N_11610,N_9134);
or U14824 (N_14824,N_10465,N_9118);
xor U14825 (N_14825,N_11056,N_11424);
and U14826 (N_14826,N_9454,N_9391);
xnor U14827 (N_14827,N_11183,N_11167);
nor U14828 (N_14828,N_9180,N_10840);
xor U14829 (N_14829,N_11933,N_9561);
nand U14830 (N_14830,N_10283,N_9766);
nand U14831 (N_14831,N_10115,N_11470);
xor U14832 (N_14832,N_10760,N_10700);
or U14833 (N_14833,N_9305,N_11538);
xor U14834 (N_14834,N_10103,N_9062);
nor U14835 (N_14835,N_11440,N_9701);
xnor U14836 (N_14836,N_11150,N_9982);
and U14837 (N_14837,N_10593,N_9987);
and U14838 (N_14838,N_9084,N_10839);
and U14839 (N_14839,N_10449,N_10862);
xor U14840 (N_14840,N_10255,N_10793);
xor U14841 (N_14841,N_11209,N_11440);
xor U14842 (N_14842,N_11293,N_11879);
nor U14843 (N_14843,N_11973,N_9512);
nor U14844 (N_14844,N_11544,N_9019);
and U14845 (N_14845,N_9259,N_9738);
or U14846 (N_14846,N_11032,N_9679);
xor U14847 (N_14847,N_10167,N_10441);
xnor U14848 (N_14848,N_10675,N_10061);
or U14849 (N_14849,N_10591,N_10916);
nand U14850 (N_14850,N_11190,N_9173);
xnor U14851 (N_14851,N_11784,N_10623);
and U14852 (N_14852,N_9832,N_11513);
and U14853 (N_14853,N_10270,N_9186);
and U14854 (N_14854,N_11639,N_11023);
and U14855 (N_14855,N_9373,N_10986);
xor U14856 (N_14856,N_10224,N_9266);
xor U14857 (N_14857,N_11311,N_11336);
or U14858 (N_14858,N_10165,N_9523);
and U14859 (N_14859,N_10656,N_11228);
nand U14860 (N_14860,N_11790,N_11455);
nor U14861 (N_14861,N_10322,N_10598);
nand U14862 (N_14862,N_10654,N_10452);
or U14863 (N_14863,N_9114,N_10191);
nand U14864 (N_14864,N_9874,N_9848);
or U14865 (N_14865,N_9446,N_11331);
nor U14866 (N_14866,N_10329,N_10823);
or U14867 (N_14867,N_9677,N_9379);
xor U14868 (N_14868,N_9123,N_10708);
nor U14869 (N_14869,N_10217,N_10395);
nand U14870 (N_14870,N_11599,N_9306);
or U14871 (N_14871,N_9675,N_9205);
or U14872 (N_14872,N_11781,N_11249);
or U14873 (N_14873,N_11700,N_10699);
nand U14874 (N_14874,N_10822,N_10597);
or U14875 (N_14875,N_10781,N_11869);
nor U14876 (N_14876,N_11757,N_10824);
or U14877 (N_14877,N_10887,N_11588);
nand U14878 (N_14878,N_9891,N_10774);
or U14879 (N_14879,N_9217,N_11288);
nor U14880 (N_14880,N_10717,N_9947);
xnor U14881 (N_14881,N_11198,N_10491);
or U14882 (N_14882,N_11736,N_9596);
nor U14883 (N_14883,N_11336,N_10519);
xor U14884 (N_14884,N_9463,N_9156);
and U14885 (N_14885,N_9177,N_11244);
or U14886 (N_14886,N_10450,N_9621);
xor U14887 (N_14887,N_10384,N_11484);
and U14888 (N_14888,N_10511,N_11878);
or U14889 (N_14889,N_10630,N_9598);
and U14890 (N_14890,N_11718,N_9610);
nand U14891 (N_14891,N_9362,N_9403);
nor U14892 (N_14892,N_11525,N_9593);
nand U14893 (N_14893,N_10905,N_10190);
nand U14894 (N_14894,N_9216,N_9703);
nand U14895 (N_14895,N_11379,N_10206);
nand U14896 (N_14896,N_9367,N_11991);
nand U14897 (N_14897,N_11062,N_11809);
nand U14898 (N_14898,N_10733,N_10506);
xnor U14899 (N_14899,N_10186,N_11097);
nor U14900 (N_14900,N_11523,N_10913);
or U14901 (N_14901,N_11547,N_11564);
xnor U14902 (N_14902,N_10570,N_11542);
and U14903 (N_14903,N_11350,N_11370);
xnor U14904 (N_14904,N_11821,N_9939);
and U14905 (N_14905,N_11313,N_11831);
nand U14906 (N_14906,N_9601,N_11606);
nor U14907 (N_14907,N_11782,N_9464);
and U14908 (N_14908,N_10182,N_10077);
and U14909 (N_14909,N_11504,N_10821);
nor U14910 (N_14910,N_10204,N_11094);
xor U14911 (N_14911,N_9197,N_11963);
nor U14912 (N_14912,N_11235,N_10799);
xor U14913 (N_14913,N_11442,N_11853);
nand U14914 (N_14914,N_9351,N_11467);
or U14915 (N_14915,N_10950,N_10122);
or U14916 (N_14916,N_11188,N_10884);
xnor U14917 (N_14917,N_9612,N_10531);
xor U14918 (N_14918,N_9734,N_10379);
or U14919 (N_14919,N_9161,N_9336);
nand U14920 (N_14920,N_11800,N_10685);
and U14921 (N_14921,N_10027,N_9986);
nor U14922 (N_14922,N_11999,N_11389);
nor U14923 (N_14923,N_11761,N_9545);
nor U14924 (N_14924,N_9442,N_10006);
nand U14925 (N_14925,N_10645,N_9081);
nand U14926 (N_14926,N_10556,N_11535);
nand U14927 (N_14927,N_10066,N_11181);
nand U14928 (N_14928,N_11217,N_9679);
and U14929 (N_14929,N_11172,N_10650);
and U14930 (N_14930,N_9126,N_9925);
or U14931 (N_14931,N_9561,N_9800);
xor U14932 (N_14932,N_9998,N_11222);
nor U14933 (N_14933,N_9317,N_9475);
or U14934 (N_14934,N_11808,N_9021);
xor U14935 (N_14935,N_9656,N_9581);
nand U14936 (N_14936,N_11000,N_10582);
and U14937 (N_14937,N_9833,N_11091);
nor U14938 (N_14938,N_9928,N_9129);
nand U14939 (N_14939,N_11254,N_10781);
or U14940 (N_14940,N_11582,N_9447);
nor U14941 (N_14941,N_9078,N_11216);
nor U14942 (N_14942,N_9025,N_10789);
and U14943 (N_14943,N_10937,N_11557);
or U14944 (N_14944,N_11798,N_11021);
and U14945 (N_14945,N_11175,N_9957);
xor U14946 (N_14946,N_9265,N_10308);
nor U14947 (N_14947,N_9664,N_10316);
nand U14948 (N_14948,N_10666,N_10973);
or U14949 (N_14949,N_11897,N_9240);
or U14950 (N_14950,N_9602,N_9007);
xor U14951 (N_14951,N_11644,N_9574);
nand U14952 (N_14952,N_11787,N_9663);
nor U14953 (N_14953,N_10665,N_9576);
xnor U14954 (N_14954,N_10938,N_9392);
and U14955 (N_14955,N_11479,N_11825);
and U14956 (N_14956,N_9657,N_9507);
nor U14957 (N_14957,N_9752,N_9101);
xnor U14958 (N_14958,N_11272,N_9810);
xor U14959 (N_14959,N_11030,N_10955);
xor U14960 (N_14960,N_10859,N_9141);
and U14961 (N_14961,N_10366,N_10251);
and U14962 (N_14962,N_9771,N_11137);
nor U14963 (N_14963,N_10372,N_10554);
and U14964 (N_14964,N_9942,N_10872);
xnor U14965 (N_14965,N_11008,N_9624);
nor U14966 (N_14966,N_11505,N_9802);
nand U14967 (N_14967,N_9451,N_9559);
nor U14968 (N_14968,N_11782,N_9633);
and U14969 (N_14969,N_9343,N_9653);
or U14970 (N_14970,N_11410,N_9384);
xor U14971 (N_14971,N_11455,N_11290);
nor U14972 (N_14972,N_9006,N_9055);
or U14973 (N_14973,N_11784,N_10541);
nor U14974 (N_14974,N_11431,N_9341);
nor U14975 (N_14975,N_9042,N_11178);
nor U14976 (N_14976,N_10138,N_11300);
xnor U14977 (N_14977,N_10493,N_10262);
or U14978 (N_14978,N_9819,N_11930);
nand U14979 (N_14979,N_10769,N_10826);
xor U14980 (N_14980,N_10741,N_11291);
or U14981 (N_14981,N_10044,N_11021);
nand U14982 (N_14982,N_11058,N_11558);
xnor U14983 (N_14983,N_10653,N_9473);
nand U14984 (N_14984,N_11064,N_10132);
xnor U14985 (N_14985,N_9609,N_9400);
and U14986 (N_14986,N_10674,N_10916);
nor U14987 (N_14987,N_11048,N_11525);
or U14988 (N_14988,N_10640,N_9519);
nor U14989 (N_14989,N_10010,N_11164);
or U14990 (N_14990,N_9181,N_9545);
xor U14991 (N_14991,N_10890,N_11091);
nor U14992 (N_14992,N_9549,N_10900);
and U14993 (N_14993,N_11405,N_11660);
xnor U14994 (N_14994,N_10275,N_9596);
or U14995 (N_14995,N_11516,N_10100);
xor U14996 (N_14996,N_11302,N_10685);
nor U14997 (N_14997,N_11296,N_10939);
or U14998 (N_14998,N_10715,N_9298);
or U14999 (N_14999,N_11256,N_11210);
xnor UO_0 (O_0,N_13978,N_12790);
nor UO_1 (O_1,N_13635,N_14350);
xor UO_2 (O_2,N_12264,N_12077);
and UO_3 (O_3,N_12196,N_14899);
and UO_4 (O_4,N_13153,N_13433);
or UO_5 (O_5,N_13767,N_13864);
or UO_6 (O_6,N_13477,N_13743);
nand UO_7 (O_7,N_12369,N_14715);
xnor UO_8 (O_8,N_13562,N_12366);
xnor UO_9 (O_9,N_13649,N_13081);
and UO_10 (O_10,N_12182,N_14950);
or UO_11 (O_11,N_12611,N_13855);
nor UO_12 (O_12,N_12362,N_13791);
nor UO_13 (O_13,N_12856,N_14727);
and UO_14 (O_14,N_12199,N_13308);
or UO_15 (O_15,N_12844,N_12555);
or UO_16 (O_16,N_12758,N_12042);
nor UO_17 (O_17,N_12481,N_13391);
or UO_18 (O_18,N_14716,N_14709);
or UO_19 (O_19,N_14896,N_14074);
xnor UO_20 (O_20,N_14435,N_13319);
xor UO_21 (O_21,N_14490,N_14151);
nor UO_22 (O_22,N_13733,N_14517);
xor UO_23 (O_23,N_13259,N_14166);
nand UO_24 (O_24,N_13628,N_12851);
xor UO_25 (O_25,N_12859,N_13727);
xnor UO_26 (O_26,N_13837,N_12935);
xnor UO_27 (O_27,N_14681,N_12837);
xnor UO_28 (O_28,N_14158,N_14313);
and UO_29 (O_29,N_14433,N_12144);
and UO_30 (O_30,N_13088,N_12721);
nor UO_31 (O_31,N_12630,N_14340);
nand UO_32 (O_32,N_12177,N_12338);
nand UO_33 (O_33,N_14276,N_13313);
or UO_34 (O_34,N_12812,N_13728);
nand UO_35 (O_35,N_13892,N_13957);
xor UO_36 (O_36,N_12324,N_12412);
xnor UO_37 (O_37,N_13806,N_12915);
nand UO_38 (O_38,N_13414,N_12785);
or UO_39 (O_39,N_14851,N_14410);
xor UO_40 (O_40,N_13739,N_12502);
and UO_41 (O_41,N_13651,N_14335);
nand UO_42 (O_42,N_14383,N_14870);
nor UO_43 (O_43,N_14280,N_13054);
and UO_44 (O_44,N_14565,N_12883);
xor UO_45 (O_45,N_13971,N_13009);
nand UO_46 (O_46,N_14979,N_14016);
xnor UO_47 (O_47,N_14949,N_12834);
and UO_48 (O_48,N_13075,N_14978);
or UO_49 (O_49,N_13621,N_13227);
nand UO_50 (O_50,N_12120,N_14695);
and UO_51 (O_51,N_12293,N_13918);
xor UO_52 (O_52,N_14954,N_12334);
xnor UO_53 (O_53,N_13389,N_13900);
or UO_54 (O_54,N_13291,N_13766);
nor UO_55 (O_55,N_14411,N_12082);
xor UO_56 (O_56,N_12662,N_13329);
nand UO_57 (O_57,N_13147,N_12356);
or UO_58 (O_58,N_13201,N_13467);
and UO_59 (O_59,N_13662,N_13236);
and UO_60 (O_60,N_14301,N_12748);
xor UO_61 (O_61,N_14933,N_12404);
nor UO_62 (O_62,N_13976,N_12413);
nor UO_63 (O_63,N_14468,N_14580);
and UO_64 (O_64,N_12169,N_14687);
xor UO_65 (O_65,N_13744,N_13263);
or UO_66 (O_66,N_14853,N_13383);
xnor UO_67 (O_67,N_12842,N_13126);
nand UO_68 (O_68,N_13018,N_12926);
xnor UO_69 (O_69,N_13481,N_13004);
xnor UO_70 (O_70,N_13321,N_13287);
and UO_71 (O_71,N_12776,N_13560);
nand UO_72 (O_72,N_13065,N_12745);
and UO_73 (O_73,N_13652,N_14538);
nand UO_74 (O_74,N_13202,N_14389);
xnor UO_75 (O_75,N_13397,N_14033);
nor UO_76 (O_76,N_12695,N_12713);
nor UO_77 (O_77,N_12849,N_12129);
xor UO_78 (O_78,N_12532,N_12557);
and UO_79 (O_79,N_12156,N_13556);
nor UO_80 (O_80,N_14807,N_14426);
nand UO_81 (O_81,N_13582,N_13184);
or UO_82 (O_82,N_12895,N_14965);
and UO_83 (O_83,N_14866,N_13993);
nor UO_84 (O_84,N_13629,N_14234);
xor UO_85 (O_85,N_12238,N_12863);
xor UO_86 (O_86,N_13008,N_13509);
and UO_87 (O_87,N_14236,N_13352);
and UO_88 (O_88,N_13617,N_12016);
or UO_89 (O_89,N_14206,N_14099);
or UO_90 (O_90,N_12353,N_13669);
nor UO_91 (O_91,N_13545,N_13317);
nand UO_92 (O_92,N_13353,N_13949);
nand UO_93 (O_93,N_12694,N_13595);
or UO_94 (O_94,N_14698,N_13819);
or UO_95 (O_95,N_14321,N_13984);
or UO_96 (O_96,N_13226,N_12361);
or UO_97 (O_97,N_13257,N_13809);
nor UO_98 (O_98,N_12956,N_13130);
and UO_99 (O_99,N_14941,N_13922);
xnor UO_100 (O_100,N_12137,N_14876);
or UO_101 (O_101,N_14745,N_13625);
xnor UO_102 (O_102,N_14772,N_14789);
nand UO_103 (O_103,N_13941,N_13742);
or UO_104 (O_104,N_13813,N_13932);
nand UO_105 (O_105,N_14144,N_14367);
and UO_106 (O_106,N_14635,N_13547);
nand UO_107 (O_107,N_14943,N_14169);
xnor UO_108 (O_108,N_14752,N_14699);
nand UO_109 (O_109,N_12648,N_13684);
xor UO_110 (O_110,N_13262,N_12610);
xor UO_111 (O_111,N_12145,N_13139);
nor UO_112 (O_112,N_12749,N_13638);
nand UO_113 (O_113,N_13475,N_13448);
nand UO_114 (O_114,N_13511,N_14358);
xnor UO_115 (O_115,N_12917,N_12744);
or UO_116 (O_116,N_14129,N_14393);
or UO_117 (O_117,N_14838,N_14275);
nor UO_118 (O_118,N_14667,N_14156);
nand UO_119 (O_119,N_14423,N_13031);
and UO_120 (O_120,N_12435,N_13069);
nand UO_121 (O_121,N_14138,N_12551);
xnor UO_122 (O_122,N_12406,N_13023);
xor UO_123 (O_123,N_14233,N_14955);
or UO_124 (O_124,N_13268,N_14605);
xnor UO_125 (O_125,N_13415,N_12691);
or UO_126 (O_126,N_12494,N_12051);
nor UO_127 (O_127,N_13149,N_12885);
or UO_128 (O_128,N_14175,N_12706);
nor UO_129 (O_129,N_13732,N_13798);
nor UO_130 (O_130,N_13218,N_13412);
nor UO_131 (O_131,N_13936,N_12882);
nand UO_132 (O_132,N_12957,N_14946);
or UO_133 (O_133,N_13176,N_13293);
or UO_134 (O_134,N_13135,N_12805);
nand UO_135 (O_135,N_13636,N_12258);
or UO_136 (O_136,N_14534,N_13568);
nand UO_137 (O_137,N_13030,N_14572);
nand UO_138 (O_138,N_12275,N_12425);
nand UO_139 (O_139,N_12417,N_14273);
or UO_140 (O_140,N_13856,N_13722);
nand UO_141 (O_141,N_13839,N_14747);
nand UO_142 (O_142,N_14827,N_14296);
nand UO_143 (O_143,N_12954,N_12465);
nor UO_144 (O_144,N_13999,N_12910);
xor UO_145 (O_145,N_13529,N_12268);
and UO_146 (O_146,N_12821,N_14720);
or UO_147 (O_147,N_14629,N_14835);
or UO_148 (O_148,N_14343,N_13285);
and UO_149 (O_149,N_14184,N_14997);
or UO_150 (O_150,N_12677,N_12020);
or UO_151 (O_151,N_13336,N_14504);
nor UO_152 (O_152,N_13893,N_13036);
nand UO_153 (O_153,N_14120,N_13314);
or UO_154 (O_154,N_12898,N_13913);
xor UO_155 (O_155,N_12559,N_12483);
nor UO_156 (O_156,N_14109,N_13356);
nor UO_157 (O_157,N_12024,N_13827);
nand UO_158 (O_158,N_12506,N_13915);
xnor UO_159 (O_159,N_13899,N_13294);
or UO_160 (O_160,N_12942,N_13605);
and UO_161 (O_161,N_13540,N_14052);
and UO_162 (O_162,N_12535,N_13155);
nand UO_163 (O_163,N_14163,N_13843);
xnor UO_164 (O_164,N_13377,N_12030);
or UO_165 (O_165,N_14224,N_12871);
or UO_166 (O_166,N_14930,N_12605);
nand UO_167 (O_167,N_12467,N_12067);
xor UO_168 (O_168,N_12218,N_12233);
xnor UO_169 (O_169,N_12344,N_12421);
or UO_170 (O_170,N_14643,N_12322);
and UO_171 (O_171,N_13960,N_12830);
nand UO_172 (O_172,N_14799,N_13058);
or UO_173 (O_173,N_14977,N_14028);
xnor UO_174 (O_174,N_12692,N_14586);
nand UO_175 (O_175,N_12598,N_12711);
and UO_176 (O_176,N_14083,N_14985);
xor UO_177 (O_177,N_14604,N_14748);
or UO_178 (O_178,N_13192,N_12438);
and UO_179 (O_179,N_14051,N_13896);
nor UO_180 (O_180,N_12158,N_13310);
xnor UO_181 (O_181,N_14489,N_14768);
and UO_182 (O_182,N_13025,N_13944);
xor UO_183 (O_183,N_13362,N_14352);
nor UO_184 (O_184,N_13842,N_13773);
xnor UO_185 (O_185,N_13051,N_12415);
or UO_186 (O_186,N_12806,N_12866);
xnor UO_187 (O_187,N_13882,N_14778);
nand UO_188 (O_188,N_12147,N_12831);
xor UO_189 (O_189,N_14975,N_12111);
or UO_190 (O_190,N_14858,N_13076);
xor UO_191 (O_191,N_14320,N_14769);
and UO_192 (O_192,N_14781,N_14812);
or UO_193 (O_193,N_13254,N_12004);
xor UO_194 (O_194,N_13079,N_12731);
or UO_195 (O_195,N_14159,N_14563);
nor UO_196 (O_196,N_13221,N_13368);
xnor UO_197 (O_197,N_14019,N_12347);
or UO_198 (O_198,N_14111,N_13951);
or UO_199 (O_199,N_13926,N_13979);
and UO_200 (O_200,N_12088,N_12793);
and UO_201 (O_201,N_13679,N_13363);
xnor UO_202 (O_202,N_14735,N_14114);
and UO_203 (O_203,N_13462,N_13042);
and UO_204 (O_204,N_14971,N_13988);
nand UO_205 (O_205,N_14274,N_14334);
nand UO_206 (O_206,N_12444,N_14327);
nand UO_207 (O_207,N_13771,N_14270);
xor UO_208 (O_208,N_13003,N_12044);
xnor UO_209 (O_209,N_12623,N_13698);
or UO_210 (O_210,N_12634,N_14685);
nor UO_211 (O_211,N_12337,N_12877);
nand UO_212 (O_212,N_14663,N_14872);
xor UO_213 (O_213,N_14951,N_14628);
nor UO_214 (O_214,N_14484,N_12697);
or UO_215 (O_215,N_13749,N_14392);
xnor UO_216 (O_216,N_13376,N_13062);
xnor UO_217 (O_217,N_12643,N_12835);
nand UO_218 (O_218,N_12582,N_12174);
nor UO_219 (O_219,N_13863,N_14372);
nor UO_220 (O_220,N_13333,N_13360);
or UO_221 (O_221,N_12259,N_14124);
nand UO_222 (O_222,N_12981,N_13750);
nor UO_223 (O_223,N_12389,N_14329);
xnor UO_224 (O_224,N_14888,N_13063);
and UO_225 (O_225,N_14326,N_12450);
nand UO_226 (O_226,N_13323,N_12803);
xnor UO_227 (O_227,N_12724,N_14214);
and UO_228 (O_228,N_14211,N_13061);
or UO_229 (O_229,N_12606,N_13425);
and UO_230 (O_230,N_14505,N_13027);
and UO_231 (O_231,N_14762,N_14331);
xnor UO_232 (O_232,N_12489,N_13760);
xnor UO_233 (O_233,N_12862,N_13538);
nor UO_234 (O_234,N_12759,N_14450);
xnor UO_235 (O_235,N_12115,N_14438);
nand UO_236 (O_236,N_12755,N_12720);
and UO_237 (O_237,N_13965,N_14314);
xnor UO_238 (O_238,N_12968,N_14623);
nor UO_239 (O_239,N_13029,N_14365);
xor UO_240 (O_240,N_12187,N_13041);
nand UO_241 (O_241,N_13386,N_14228);
and UO_242 (O_242,N_12326,N_12358);
xor UO_243 (O_243,N_14652,N_12305);
xnor UO_244 (O_244,N_14839,N_12038);
xor UO_245 (O_245,N_12712,N_14680);
or UO_246 (O_246,N_14302,N_13205);
xor UO_247 (O_247,N_13850,N_12511);
or UO_248 (O_248,N_13644,N_14904);
and UO_249 (O_249,N_13172,N_14692);
nor UO_250 (O_250,N_12041,N_13945);
and UO_251 (O_251,N_12487,N_14377);
or UO_252 (O_252,N_14469,N_12280);
or UO_253 (O_253,N_14493,N_13495);
or UO_254 (O_254,N_13056,N_13518);
or UO_255 (O_255,N_12927,N_14487);
nor UO_256 (O_256,N_14829,N_14025);
nand UO_257 (O_257,N_14195,N_14265);
and UO_258 (O_258,N_14834,N_14688);
or UO_259 (O_259,N_13464,N_14104);
or UO_260 (O_260,N_12140,N_13459);
nand UO_261 (O_261,N_13458,N_14179);
or UO_262 (O_262,N_14064,N_14671);
nand UO_263 (O_263,N_12544,N_12271);
xnor UO_264 (O_264,N_13115,N_14137);
nand UO_265 (O_265,N_14561,N_14649);
nand UO_266 (O_266,N_13752,N_14323);
nor UO_267 (O_267,N_14048,N_13347);
nand UO_268 (O_268,N_13493,N_12249);
nor UO_269 (O_269,N_12734,N_12323);
and UO_270 (O_270,N_13532,N_12860);
nor UO_271 (O_271,N_12523,N_13453);
nor UO_272 (O_272,N_14055,N_12874);
nand UO_273 (O_273,N_13134,N_14402);
or UO_274 (O_274,N_14336,N_12315);
nor UO_275 (O_275,N_14470,N_14989);
nand UO_276 (O_276,N_13898,N_12384);
and UO_277 (O_277,N_14887,N_13515);
nand UO_278 (O_278,N_13755,N_12272);
xor UO_279 (O_279,N_14012,N_12383);
or UO_280 (O_280,N_13197,N_13935);
or UO_281 (O_281,N_12161,N_12900);
and UO_282 (O_282,N_12390,N_14272);
xor UO_283 (O_283,N_12951,N_13074);
xor UO_284 (O_284,N_14444,N_14738);
and UO_285 (O_285,N_13534,N_14601);
or UO_286 (O_286,N_14293,N_14987);
nor UO_287 (O_287,N_12060,N_13354);
nor UO_288 (O_288,N_12922,N_14893);
nor UO_289 (O_289,N_13653,N_12352);
nand UO_290 (O_290,N_13418,N_13038);
xor UO_291 (O_291,N_12112,N_13429);
xor UO_292 (O_292,N_14714,N_12746);
or UO_293 (O_293,N_12223,N_14240);
xnor UO_294 (O_294,N_12241,N_14093);
nand UO_295 (O_295,N_12179,N_13120);
nand UO_296 (O_296,N_14564,N_14934);
nand UO_297 (O_297,N_14066,N_13726);
and UO_298 (O_298,N_13174,N_12318);
xnor UO_299 (O_299,N_12011,N_13589);
nand UO_300 (O_300,N_14506,N_12094);
nor UO_301 (O_301,N_13001,N_14848);
and UO_302 (O_302,N_12048,N_12876);
nand UO_303 (O_303,N_13840,N_12451);
and UO_304 (O_304,N_14204,N_13339);
xnor UO_305 (O_305,N_12828,N_12902);
and UO_306 (O_306,N_12747,N_14759);
nor UO_307 (O_307,N_12609,N_12001);
or UO_308 (O_308,N_13388,N_14004);
nand UO_309 (O_309,N_12864,N_13588);
and UO_310 (O_310,N_12059,N_13512);
xor UO_311 (O_311,N_12717,N_14961);
or UO_312 (O_312,N_13758,N_14128);
and UO_313 (O_313,N_13478,N_13359);
nor UO_314 (O_314,N_14386,N_12649);
nor UO_315 (O_315,N_13133,N_13154);
xnor UO_316 (O_316,N_13832,N_13504);
nor UO_317 (O_317,N_12043,N_14528);
or UO_318 (O_318,N_12750,N_13994);
nand UO_319 (O_319,N_13483,N_12991);
and UO_320 (O_320,N_13626,N_12650);
xnor UO_321 (O_321,N_14146,N_13402);
nand UO_322 (O_322,N_13920,N_14106);
nand UO_323 (O_323,N_12032,N_12313);
and UO_324 (O_324,N_12301,N_13812);
or UO_325 (O_325,N_12901,N_12567);
or UO_326 (O_326,N_14518,N_12961);
nand UO_327 (O_327,N_14957,N_12046);
nor UO_328 (O_328,N_12367,N_12297);
nor UO_329 (O_329,N_14057,N_12693);
or UO_330 (O_330,N_13704,N_13769);
nand UO_331 (O_331,N_13972,N_13472);
xor UO_332 (O_332,N_13923,N_14614);
or UO_333 (O_333,N_14330,N_13925);
xor UO_334 (O_334,N_12289,N_14816);
or UO_335 (O_335,N_14777,N_13200);
nand UO_336 (O_336,N_14626,N_13252);
nand UO_337 (O_337,N_14886,N_14600);
nor UO_338 (O_338,N_12385,N_14341);
nand UO_339 (O_339,N_14262,N_13666);
nor UO_340 (O_340,N_13044,N_12023);
xor UO_341 (O_341,N_12047,N_14067);
and UO_342 (O_342,N_14193,N_12185);
nor UO_343 (O_343,N_14814,N_13593);
xnor UO_344 (O_344,N_12992,N_14303);
and UO_345 (O_345,N_13232,N_14573);
and UO_346 (O_346,N_13690,N_12778);
or UO_347 (O_347,N_14471,N_14203);
nand UO_348 (O_348,N_12537,N_14292);
or UO_349 (O_349,N_14122,N_13366);
nand UO_350 (O_350,N_12854,N_12946);
xor UO_351 (O_351,N_14920,N_14147);
nand UO_352 (O_352,N_12267,N_13709);
or UO_353 (O_353,N_12287,N_14325);
nor UO_354 (O_354,N_13423,N_14480);
or UO_355 (O_355,N_13536,N_13114);
or UO_356 (O_356,N_14637,N_13408);
and UO_357 (O_357,N_13267,N_12867);
and UO_358 (O_358,N_14967,N_12260);
xor UO_359 (O_359,N_14982,N_14399);
nor UO_360 (O_360,N_14578,N_12243);
or UO_361 (O_361,N_14006,N_13675);
nand UO_362 (O_362,N_13455,N_13665);
nor UO_363 (O_363,N_13078,N_12012);
nand UO_364 (O_364,N_12843,N_13590);
or UO_365 (O_365,N_13122,N_13530);
and UO_366 (O_366,N_12125,N_12525);
xnor UO_367 (O_367,N_14220,N_12540);
and UO_368 (O_368,N_12845,N_13325);
nor UO_369 (O_369,N_13503,N_12784);
nor UO_370 (O_370,N_12325,N_12807);
or UO_371 (O_371,N_12897,N_12302);
nand UO_372 (O_372,N_12832,N_12312);
xnor UO_373 (O_373,N_12800,N_12150);
nand UO_374 (O_374,N_12869,N_12022);
nor UO_375 (O_375,N_12064,N_13270);
nor UO_376 (O_376,N_14645,N_14463);
xnor UO_377 (O_377,N_13631,N_13370);
nor UO_378 (O_378,N_14247,N_14523);
nand UO_379 (O_379,N_13298,N_13245);
and UO_380 (O_380,N_14105,N_13601);
and UO_381 (O_381,N_12918,N_13528);
nor UO_382 (O_382,N_13373,N_14854);
nand UO_383 (O_383,N_12645,N_13702);
xnor UO_384 (O_384,N_13158,N_12118);
nand UO_385 (O_385,N_14269,N_12127);
and UO_386 (O_386,N_14909,N_13874);
and UO_387 (O_387,N_12841,N_12090);
nand UO_388 (O_388,N_12732,N_13486);
or UO_389 (O_389,N_12890,N_12079);
xnor UO_390 (O_390,N_12222,N_13656);
xor UO_391 (O_391,N_13161,N_12943);
xor UO_392 (O_392,N_14542,N_14865);
and UO_393 (O_393,N_12827,N_14912);
xnor UO_394 (O_394,N_12121,N_14010);
and UO_395 (O_395,N_13106,N_13318);
and UO_396 (O_396,N_12808,N_12458);
or UO_397 (O_397,N_14889,N_13144);
nand UO_398 (O_398,N_13094,N_14071);
and UO_399 (O_399,N_14624,N_14429);
nand UO_400 (O_400,N_14213,N_14696);
nor UO_401 (O_401,N_14574,N_12442);
nand UO_402 (O_402,N_13833,N_13189);
or UO_403 (O_403,N_13607,N_14097);
nor UO_404 (O_404,N_14113,N_13775);
xnor UO_405 (O_405,N_13165,N_12251);
nand UO_406 (O_406,N_12063,N_13187);
nand UO_407 (O_407,N_14801,N_12892);
nor UO_408 (O_408,N_14774,N_12853);
xor UO_409 (O_409,N_12240,N_13533);
and UO_410 (O_410,N_12328,N_14910);
nand UO_411 (O_411,N_14364,N_14053);
and UO_412 (O_412,N_14237,N_14069);
nor UO_413 (O_413,N_14821,N_13177);
or UO_414 (O_414,N_12086,N_12363);
or UO_415 (O_415,N_14371,N_13664);
and UO_416 (O_416,N_12663,N_13962);
nand UO_417 (O_417,N_13085,N_14973);
or UO_418 (O_418,N_14255,N_14116);
nor UO_419 (O_419,N_13346,N_13282);
nor UO_420 (O_420,N_13860,N_12524);
xor UO_421 (O_421,N_14485,N_12343);
or UO_422 (O_422,N_12128,N_12180);
or UO_423 (O_423,N_14627,N_13734);
xnor UO_424 (O_424,N_12230,N_14640);
xor UO_425 (O_425,N_12207,N_13524);
xnor UO_426 (O_426,N_14757,N_13351);
or UO_427 (O_427,N_12080,N_14880);
nand UO_428 (O_428,N_13513,N_12789);
nand UO_429 (O_429,N_13740,N_12742);
and UO_430 (O_430,N_13703,N_12545);
or UO_431 (O_431,N_12183,N_12549);
xnor UO_432 (O_432,N_14474,N_14874);
nand UO_433 (O_433,N_13977,N_13330);
or UO_434 (O_434,N_12163,N_14186);
and UO_435 (O_435,N_13692,N_13148);
or UO_436 (O_436,N_13517,N_12938);
nor UO_437 (O_437,N_14672,N_14664);
xor UO_438 (O_438,N_14775,N_14907);
nor UO_439 (O_439,N_12996,N_13516);
nand UO_440 (O_440,N_13810,N_13442);
or UO_441 (O_441,N_14728,N_14661);
nand UO_442 (O_442,N_14408,N_12463);
nand UO_443 (O_443,N_13747,N_12887);
nand UO_444 (O_444,N_14345,N_14976);
nor UO_445 (O_445,N_12409,N_12773);
or UO_446 (O_446,N_12948,N_14923);
and UO_447 (O_447,N_14232,N_12424);
or UO_448 (O_448,N_14322,N_12584);
nor UO_449 (O_449,N_13279,N_12055);
xor UO_450 (O_450,N_14431,N_12528);
and UO_451 (O_451,N_12533,N_12420);
or UO_452 (O_452,N_14266,N_13372);
and UO_453 (O_453,N_13985,N_12165);
nand UO_454 (O_454,N_13875,N_14621);
nor UO_455 (O_455,N_13676,N_12432);
nor UO_456 (O_456,N_13577,N_12242);
xnor UO_457 (O_457,N_13214,N_13320);
or UO_458 (O_458,N_13680,N_12518);
xor UO_459 (O_459,N_14964,N_14861);
nand UO_460 (O_460,N_13328,N_13620);
xnor UO_461 (O_461,N_12542,N_14890);
and UO_462 (O_462,N_13278,N_14915);
xnor UO_463 (O_463,N_14200,N_14729);
and UO_464 (O_464,N_14183,N_13506);
nor UO_465 (O_465,N_13841,N_13411);
nor UO_466 (O_466,N_13342,N_12941);
nand UO_467 (O_467,N_12775,N_13124);
and UO_468 (O_468,N_13399,N_14355);
nor UO_469 (O_469,N_12791,N_12014);
and UO_470 (O_470,N_14787,N_13491);
and UO_471 (O_471,N_13683,N_12469);
nand UO_472 (O_472,N_13204,N_14388);
and UO_473 (O_473,N_12382,N_12794);
nand UO_474 (O_474,N_14811,N_13379);
xnor UO_475 (O_475,N_14583,N_13422);
nor UO_476 (O_476,N_12612,N_13343);
xor UO_477 (O_477,N_13569,N_12427);
xor UO_478 (O_478,N_12381,N_13852);
and UO_479 (O_479,N_13142,N_14676);
and UO_480 (O_480,N_12680,N_14291);
xnor UO_481 (O_481,N_13557,N_12893);
or UO_482 (O_482,N_13431,N_12636);
or UO_483 (O_483,N_14342,N_14921);
nand UO_484 (O_484,N_14094,N_12217);
nand UO_485 (O_485,N_12653,N_13658);
and UO_486 (O_486,N_14842,N_13667);
nand UO_487 (O_487,N_13998,N_13384);
nor UO_488 (O_488,N_14143,N_14205);
xnor UO_489 (O_489,N_14589,N_14859);
xnor UO_490 (O_490,N_14346,N_12577);
xnor UO_491 (O_491,N_14013,N_14647);
or UO_492 (O_492,N_12049,N_13865);
nor UO_493 (O_493,N_12684,N_13717);
or UO_494 (O_494,N_13434,N_13931);
or UO_495 (O_495,N_12933,N_13910);
and UO_496 (O_496,N_13095,N_14936);
nand UO_497 (O_497,N_13781,N_14980);
and UO_498 (O_498,N_14825,N_14308);
xnor UO_499 (O_499,N_13242,N_14000);
or UO_500 (O_500,N_14488,N_13815);
nor UO_501 (O_501,N_13946,N_12686);
and UO_502 (O_502,N_13273,N_13693);
and UO_503 (O_503,N_12689,N_12262);
xor UO_504 (O_504,N_13141,N_13844);
or UO_505 (O_505,N_13203,N_14836);
nor UO_506 (O_506,N_14502,N_14536);
nand UO_507 (O_507,N_12408,N_14465);
and UO_508 (O_508,N_13016,N_14446);
or UO_509 (O_509,N_12767,N_12920);
nor UO_510 (O_510,N_14042,N_13987);
xor UO_511 (O_511,N_12194,N_13138);
nand UO_512 (O_512,N_13300,N_14994);
and UO_513 (O_513,N_13033,N_13659);
xor UO_514 (O_514,N_13792,N_12906);
or UO_515 (O_515,N_12644,N_14086);
nand UO_516 (O_516,N_12716,N_12164);
or UO_517 (O_517,N_14368,N_14723);
xor UO_518 (O_518,N_12423,N_12798);
nand UO_519 (O_519,N_13969,N_13697);
or UO_520 (O_520,N_12886,N_13641);
nand UO_521 (O_521,N_14883,N_12062);
and UO_522 (O_522,N_12912,N_13447);
and UO_523 (O_523,N_13274,N_14719);
and UO_524 (O_524,N_12726,N_12459);
xor UO_525 (O_525,N_13216,N_14295);
nor UO_526 (O_526,N_12846,N_12960);
nand UO_527 (O_527,N_14473,N_13770);
nand UO_528 (O_528,N_12959,N_14333);
xnor UO_529 (O_529,N_14478,N_13312);
nor UO_530 (O_530,N_14659,N_12817);
or UO_531 (O_531,N_13387,N_14472);
and UO_532 (O_532,N_14639,N_14673);
or UO_533 (O_533,N_14570,N_13052);
nor UO_534 (O_534,N_14611,N_13816);
nor UO_535 (O_535,N_14513,N_14282);
or UO_536 (O_536,N_12604,N_13022);
xor UO_537 (O_537,N_12526,N_12529);
or UO_538 (O_538,N_13365,N_13190);
nor UO_539 (O_539,N_14284,N_14417);
or UO_540 (O_540,N_12285,N_14569);
or UO_541 (O_541,N_12407,N_14996);
and UO_542 (O_542,N_14537,N_13083);
nand UO_543 (O_543,N_12092,N_13289);
nor UO_544 (O_544,N_13045,N_14032);
nand UO_545 (O_545,N_13143,N_12321);
xor UO_546 (O_546,N_12105,N_13763);
nor UO_547 (O_547,N_12578,N_13974);
or UO_548 (O_548,N_13225,N_13660);
nand UO_549 (O_549,N_14118,N_13059);
and UO_550 (O_550,N_14922,N_14458);
nor UO_551 (O_551,N_13239,N_14516);
and UO_552 (O_552,N_14145,N_12671);
nand UO_553 (O_553,N_12221,N_14588);
and UO_554 (O_554,N_13299,N_12641);
or UO_555 (O_555,N_13654,N_13811);
and UO_556 (O_556,N_13034,N_13606);
or UO_557 (O_557,N_13990,N_12660);
and UO_558 (O_558,N_12857,N_13017);
and UO_559 (O_559,N_14660,N_13884);
or UO_560 (O_560,N_12211,N_13829);
nor UO_561 (O_561,N_14268,N_12678);
and UO_562 (O_562,N_14185,N_12498);
nand UO_563 (O_563,N_14885,N_13657);
or UO_564 (O_564,N_12492,N_12355);
nand UO_565 (O_565,N_12548,N_14078);
or UO_566 (O_566,N_13021,N_12513);
xnor UO_567 (O_567,N_12547,N_13753);
and UO_568 (O_568,N_12116,N_14746);
or UO_569 (O_569,N_14167,N_13244);
and UO_570 (O_570,N_12654,N_12411);
nor UO_571 (O_571,N_12894,N_13420);
nand UO_572 (O_572,N_14020,N_14654);
and UO_573 (O_573,N_12146,N_13871);
or UO_574 (O_574,N_12261,N_14644);
and UO_575 (O_575,N_12591,N_14925);
nand UO_576 (O_576,N_14315,N_12034);
xnor UO_577 (O_577,N_12531,N_14191);
xnor UO_578 (O_578,N_13006,N_12760);
and UO_579 (O_579,N_13406,N_12566);
xnor UO_580 (O_580,N_12206,N_12357);
and UO_581 (O_581,N_14993,N_12814);
nand UO_582 (O_582,N_12391,N_12945);
nor UO_583 (O_583,N_14514,N_14963);
nand UO_584 (O_584,N_12665,N_12205);
or UO_585 (O_585,N_12795,N_14613);
xnor UO_586 (O_586,N_13380,N_14855);
nor UO_587 (O_587,N_12215,N_13927);
and UO_588 (O_588,N_12093,N_13335);
and UO_589 (O_589,N_13870,N_13255);
and UO_590 (O_590,N_14591,N_12980);
and UO_591 (O_591,N_14180,N_12319);
and UO_592 (O_592,N_13084,N_13451);
nor UO_593 (O_593,N_14174,N_13761);
or UO_594 (O_594,N_13762,N_14027);
and UO_595 (O_595,N_12452,N_13764);
and UO_596 (O_596,N_13212,N_14337);
and UO_597 (O_597,N_12517,N_14771);
xnor UO_598 (O_598,N_13170,N_14641);
nand UO_599 (O_599,N_12735,N_13419);
or UO_600 (O_600,N_14316,N_13228);
xnor UO_601 (O_601,N_14873,N_14869);
nor UO_602 (O_602,N_14724,N_14394);
xor UO_603 (O_603,N_14646,N_12433);
xor UO_604 (O_604,N_14054,N_14575);
nand UO_605 (O_605,N_12763,N_14238);
nor UO_606 (O_606,N_14631,N_12594);
and UO_607 (O_607,N_14535,N_14711);
or UO_608 (O_608,N_14310,N_12588);
or UO_609 (O_609,N_12482,N_12561);
nor UO_610 (O_610,N_14153,N_14462);
xnor UO_611 (O_611,N_14362,N_14045);
and UO_612 (O_612,N_12681,N_14115);
and UO_613 (O_613,N_12342,N_14384);
nor UO_614 (O_614,N_12117,N_14823);
nand UO_615 (O_615,N_12679,N_13950);
nand UO_616 (O_616,N_13956,N_14261);
and UO_617 (O_617,N_12858,N_13663);
nor UO_618 (O_618,N_12453,N_12377);
nand UO_619 (O_619,N_12766,N_13916);
xor UO_620 (O_620,N_14710,N_14387);
nor UO_621 (O_621,N_12534,N_14080);
nor UO_622 (O_622,N_13904,N_12227);
or UO_623 (O_623,N_14798,N_14697);
xor UO_624 (O_624,N_14059,N_14095);
or UO_625 (O_625,N_13100,N_13756);
or UO_626 (O_626,N_12015,N_14419);
nor UO_627 (O_627,N_13521,N_12829);
nand UO_628 (O_628,N_14062,N_13952);
nor UO_629 (O_629,N_13470,N_14353);
nor UO_630 (O_630,N_13527,N_14087);
xnor UO_631 (O_631,N_12971,N_13057);
and UO_632 (O_632,N_14089,N_14625);
xnor UO_633 (O_633,N_14712,N_14283);
and UO_634 (O_634,N_12197,N_14281);
nand UO_635 (O_635,N_14751,N_13673);
xor UO_636 (O_636,N_12836,N_13011);
or UO_637 (O_637,N_12855,N_14892);
xnor UO_638 (O_638,N_14400,N_13401);
nor UO_639 (O_639,N_14198,N_13596);
xnor UO_640 (O_640,N_13456,N_14991);
and UO_641 (O_641,N_13047,N_12003);
nand UO_642 (O_642,N_12515,N_12470);
and UO_643 (O_643,N_14150,N_12429);
nand UO_644 (O_644,N_13297,N_14562);
nor UO_645 (O_645,N_13902,N_13535);
xor UO_646 (O_646,N_14457,N_14721);
and UO_647 (O_647,N_14134,N_13253);
or UO_648 (O_648,N_14413,N_12558);
nand UO_649 (O_649,N_13938,N_12255);
xnor UO_650 (O_650,N_14294,N_13807);
and UO_651 (O_651,N_14103,N_13718);
nor UO_652 (O_652,N_13729,N_12765);
and UO_653 (O_653,N_12710,N_12571);
xnor UO_654 (O_654,N_12536,N_12277);
nor UO_655 (O_655,N_13436,N_14686);
or UO_656 (O_656,N_13686,N_13525);
and UO_657 (O_657,N_13162,N_13000);
or UO_658 (O_658,N_12656,N_14416);
xor UO_659 (O_659,N_12603,N_13575);
nand UO_660 (O_660,N_14477,N_14190);
nor UO_661 (O_661,N_12278,N_12516);
and UO_662 (O_662,N_13460,N_14567);
nor UO_663 (O_663,N_14250,N_12704);
xor UO_664 (O_664,N_13055,N_12476);
nand UO_665 (O_665,N_12076,N_12572);
or UO_666 (O_666,N_13624,N_14897);
and UO_667 (O_667,N_13633,N_12965);
or UO_668 (O_668,N_14615,N_14598);
nor UO_669 (O_669,N_14073,N_12950);
and UO_670 (O_670,N_13355,N_14938);
xor UO_671 (O_671,N_14924,N_14168);
nand UO_672 (O_672,N_12539,N_12617);
nand UO_673 (O_673,N_14475,N_14123);
or UO_674 (O_674,N_13613,N_13129);
and UO_675 (O_675,N_13921,N_12899);
nor UO_676 (O_676,N_12040,N_12714);
nand UO_677 (O_677,N_14770,N_14454);
xor UO_678 (O_678,N_14522,N_12930);
or UO_679 (O_679,N_13385,N_13465);
xnor UO_680 (O_680,N_14005,N_13866);
and UO_681 (O_681,N_14249,N_14125);
nor UO_682 (O_682,N_12426,N_14555);
nor UO_683 (O_683,N_12993,N_12700);
nor UO_684 (O_684,N_13616,N_12581);
nand UO_685 (O_685,N_12069,N_13492);
xnor UO_686 (O_686,N_14041,N_14986);
xor UO_687 (O_687,N_13322,N_14347);
nand UO_688 (O_688,N_14606,N_12550);
and UO_689 (O_689,N_14656,N_13146);
or UO_690 (O_690,N_12018,N_12543);
nor UO_691 (O_691,N_13037,N_12698);
and UO_692 (O_692,N_13597,N_13830);
or UO_693 (O_693,N_14779,N_12436);
nand UO_694 (O_694,N_12216,N_14015);
nor UO_695 (O_695,N_12982,N_14901);
and UO_696 (O_696,N_13132,N_12496);
or UO_697 (O_697,N_12316,N_13677);
or UO_698 (O_698,N_14917,N_12007);
or UO_699 (O_699,N_14974,N_12676);
xnor UO_700 (O_700,N_13010,N_12512);
or UO_701 (O_701,N_14913,N_13785);
nand UO_702 (O_702,N_13395,N_14031);
or UO_703 (O_703,N_13145,N_14593);
nand UO_704 (O_704,N_13375,N_13404);
xor UO_705 (O_705,N_13539,N_12266);
xor UO_706 (O_706,N_14075,N_13937);
or UO_707 (O_707,N_14260,N_13237);
xor UO_708 (O_708,N_12659,N_13275);
and UO_709 (O_709,N_12881,N_14217);
xnor UO_710 (O_710,N_13382,N_14263);
and UO_711 (O_711,N_14786,N_12607);
xnor UO_712 (O_712,N_12033,N_14532);
and UO_713 (O_713,N_13378,N_12212);
nor UO_714 (O_714,N_14304,N_13191);
and UO_715 (O_715,N_14678,N_12071);
xor UO_716 (O_716,N_12108,N_14152);
or UO_717 (O_717,N_14132,N_12878);
and UO_718 (O_718,N_14448,N_14451);
nand UO_719 (O_719,N_12985,N_14359);
or UO_720 (O_720,N_14773,N_12647);
or UO_721 (O_721,N_13955,N_12176);
nor UO_722 (O_722,N_12657,N_12977);
xnor UO_723 (O_723,N_14306,N_14741);
xor UO_724 (O_724,N_12107,N_12987);
nand UO_725 (O_725,N_12410,N_14905);
xnor UO_726 (O_726,N_13507,N_14852);
nor UO_727 (O_727,N_14999,N_14085);
and UO_728 (O_728,N_14783,N_14879);
and UO_729 (O_729,N_14436,N_14357);
xnor UO_730 (O_730,N_13867,N_14221);
or UO_731 (O_731,N_12824,N_13572);
nand UO_732 (O_732,N_14023,N_13446);
nand UO_733 (O_733,N_14882,N_12964);
xor UO_734 (O_734,N_13853,N_12270);
nand UO_735 (O_735,N_12010,N_12932);
and UO_736 (O_736,N_14795,N_13501);
xnor UO_737 (O_737,N_12769,N_13432);
nand UO_738 (O_738,N_13991,N_14305);
nor UO_739 (O_739,N_13005,N_14090);
and UO_740 (O_740,N_12655,N_12159);
nor UO_741 (O_741,N_12477,N_12388);
and UO_742 (O_742,N_13440,N_14792);
nand UO_743 (O_743,N_12908,N_14026);
xor UO_744 (O_744,N_14894,N_13441);
xnor UO_745 (O_745,N_13367,N_13166);
nor UO_746 (O_746,N_14529,N_14047);
and UO_747 (O_747,N_14088,N_12310);
nor UO_748 (O_748,N_13332,N_12909);
nor UO_749 (O_749,N_13123,N_12919);
nand UO_750 (O_750,N_14927,N_14797);
nor UO_751 (O_751,N_12967,N_14968);
and UO_752 (O_752,N_13393,N_14501);
and UO_753 (O_753,N_14929,N_12101);
nand UO_754 (O_754,N_12786,N_14966);
nand UO_755 (O_755,N_13426,N_13724);
xor UO_756 (O_756,N_13803,N_12336);
or UO_757 (O_757,N_13183,N_12296);
nor UO_758 (O_758,N_14319,N_14653);
or UO_759 (O_759,N_14092,N_12562);
or UO_760 (O_760,N_12729,N_14142);
xnor UO_761 (O_761,N_13789,N_13219);
and UO_762 (O_762,N_12576,N_12952);
xor UO_763 (O_763,N_12944,N_14655);
xnor UO_764 (O_764,N_12246,N_13646);
and UO_765 (O_765,N_12696,N_12300);
nor UO_766 (O_766,N_12292,N_12035);
nand UO_767 (O_767,N_13151,N_13510);
or UO_768 (O_768,N_13118,N_13928);
or UO_769 (O_769,N_13272,N_13053);
nor UO_770 (O_770,N_12339,N_14403);
nor UO_771 (O_771,N_12601,N_13235);
nand UO_772 (O_772,N_13901,N_12625);
nand UO_773 (O_773,N_13966,N_13661);
and UO_774 (O_774,N_14530,N_13164);
nand UO_775 (O_775,N_13514,N_13064);
or UO_776 (O_776,N_14928,N_13240);
nor UO_777 (O_777,N_14822,N_13642);
nand UO_778 (O_778,N_12674,N_13110);
nor UO_779 (O_779,N_14212,N_13602);
nand UO_780 (O_780,N_12039,N_14030);
nor UO_781 (O_781,N_14636,N_12078);
and UO_782 (O_782,N_14210,N_13251);
and UO_783 (O_783,N_12168,N_13580);
nand UO_784 (O_784,N_14441,N_13583);
and UO_785 (O_785,N_14508,N_12756);
nor UO_786 (O_786,N_14229,N_12787);
and UO_787 (O_787,N_14267,N_13357);
and UO_788 (O_788,N_12570,N_14553);
xnor UO_789 (O_789,N_13438,N_14556);
nand UO_790 (O_790,N_12274,N_13409);
nor UO_791 (O_791,N_12000,N_13958);
nor UO_792 (O_792,N_12028,N_14794);
and UO_793 (O_793,N_14940,N_13463);
or UO_794 (O_794,N_13248,N_14467);
nand UO_795 (O_795,N_14510,N_14800);
and UO_796 (O_796,N_14397,N_14962);
nand UO_797 (O_797,N_13163,N_14207);
and UO_798 (O_798,N_13159,N_13828);
nor UO_799 (O_799,N_12119,N_12519);
xnor UO_800 (O_800,N_12801,N_12936);
or UO_801 (O_801,N_13020,N_14524);
and UO_802 (O_802,N_14891,N_13048);
xnor UO_803 (O_803,N_14763,N_14900);
xor UO_804 (O_804,N_12818,N_12762);
xnor UO_805 (O_805,N_13101,N_13716);
and UO_806 (O_806,N_12669,N_12131);
or UO_807 (O_807,N_13340,N_13805);
nand UO_808 (O_808,N_12393,N_13039);
nand UO_809 (O_809,N_12368,N_13028);
and UO_810 (O_810,N_12934,N_14197);
xnor UO_811 (O_811,N_13348,N_13073);
nand UO_812 (O_812,N_14459,N_13092);
nand UO_813 (O_813,N_12234,N_14133);
nor UO_814 (O_814,N_14065,N_12484);
and UO_815 (O_815,N_12998,N_13326);
nand UO_816 (O_816,N_12538,N_13443);
nor UO_817 (O_817,N_14937,N_13233);
nand UO_818 (O_818,N_12149,N_12279);
nand UO_819 (O_819,N_14689,N_14931);
or UO_820 (O_820,N_14286,N_12166);
or UO_821 (O_821,N_12811,N_14227);
nand UO_822 (O_822,N_13774,N_14935);
nand UO_823 (O_823,N_13883,N_14549);
or UO_824 (O_824,N_12631,N_13919);
or UO_825 (O_825,N_13211,N_14405);
nor UO_826 (O_826,N_13522,N_14121);
nand UO_827 (O_827,N_13341,N_14189);
or UO_828 (O_828,N_12799,N_12802);
or UO_829 (O_829,N_12291,N_13046);
nor UO_830 (O_830,N_14527,N_12978);
xnor UO_831 (O_831,N_14511,N_14483);
nand UO_832 (O_832,N_13707,N_12618);
xnor UO_833 (O_833,N_13639,N_14500);
and UO_834 (O_834,N_12740,N_12153);
nand UO_835 (O_835,N_12514,N_12387);
xor UO_836 (O_836,N_14434,N_13157);
nand UO_837 (O_837,N_13905,N_12333);
nor UO_838 (O_838,N_12719,N_13217);
or UO_839 (O_839,N_13277,N_14521);
nor UO_840 (O_840,N_14871,N_13599);
or UO_841 (O_841,N_12148,N_12587);
or UO_842 (O_842,N_12690,N_13911);
xor UO_843 (O_843,N_14170,N_14918);
xnor UO_844 (O_844,N_13349,N_13848);
nand UO_845 (O_845,N_12096,N_12702);
or UO_846 (O_846,N_14908,N_12008);
xnor UO_847 (O_847,N_13600,N_14597);
or UO_848 (O_848,N_14808,N_13186);
nand UO_849 (O_849,N_13914,N_12414);
nand UO_850 (O_850,N_14136,N_12733);
nor UO_851 (O_851,N_13361,N_13437);
xnor UO_852 (O_852,N_14037,N_12556);
xnor UO_853 (O_853,N_12276,N_13119);
and UO_854 (O_854,N_13302,N_13208);
xnor UO_855 (O_855,N_14638,N_12850);
and UO_856 (O_856,N_13713,N_13854);
nor UO_857 (O_857,N_14868,N_13929);
nand UO_858 (O_858,N_13428,N_12204);
xnor UO_859 (O_859,N_13563,N_13531);
nor UO_860 (O_860,N_14607,N_14650);
nor UO_861 (O_861,N_13594,N_13930);
xnor UO_862 (O_862,N_13374,N_14378);
xnor UO_863 (O_863,N_12375,N_12709);
and UO_864 (O_864,N_13947,N_12134);
xor UO_865 (O_865,N_13706,N_14682);
xor UO_866 (O_866,N_14043,N_13350);
and UO_867 (O_867,N_14739,N_14850);
and UO_868 (O_868,N_12083,N_14780);
nand UO_869 (O_869,N_12621,N_12106);
or UO_870 (O_870,N_13681,N_13645);
xnor UO_871 (O_871,N_14944,N_13392);
or UO_872 (O_872,N_14713,N_14633);
nor UO_873 (O_873,N_12298,N_13080);
nor UO_874 (O_874,N_13765,N_12741);
or UO_875 (O_875,N_13751,N_14110);
nor UO_876 (O_876,N_13831,N_13396);
nor UO_877 (O_877,N_13869,N_13292);
nor UO_878 (O_878,N_12461,N_12924);
or UO_879 (O_879,N_13735,N_12248);
nand UO_880 (O_880,N_13150,N_13570);
and UO_881 (O_881,N_13592,N_12688);
xnor UO_882 (O_882,N_13820,N_12507);
nand UO_883 (O_883,N_14253,N_12466);
nor UO_884 (O_884,N_14034,N_14076);
and UO_885 (O_885,N_14674,N_12632);
nand UO_886 (O_886,N_13614,N_12768);
and UO_887 (O_887,N_12213,N_12286);
nor UO_888 (O_888,N_14491,N_12508);
xnor UO_889 (O_889,N_13737,N_12509);
and UO_890 (O_890,N_13776,N_12896);
nand UO_891 (O_891,N_14461,N_14420);
nor UO_892 (O_892,N_13371,N_14881);
nand UO_893 (O_893,N_13885,N_12569);
nand UO_894 (O_894,N_12188,N_12100);
or UO_895 (O_895,N_14722,N_13795);
and UO_896 (O_896,N_12673,N_12913);
xnor UO_897 (O_897,N_13283,N_13835);
xor UO_898 (O_898,N_14351,N_13846);
or UO_899 (O_899,N_14243,N_12888);
or UO_900 (O_900,N_14072,N_13430);
xnor UO_901 (O_901,N_13561,N_14009);
xor UO_902 (O_902,N_13246,N_12317);
nor UO_903 (O_903,N_14793,N_12983);
nand UO_904 (O_904,N_12396,N_14691);
nand UO_905 (O_905,N_12257,N_12497);
nand UO_906 (O_906,N_12236,N_13266);
nand UO_907 (O_907,N_14373,N_14867);
and UO_908 (O_908,N_13611,N_12635);
or UO_909 (O_909,N_13598,N_12552);
and UO_910 (O_910,N_13131,N_12171);
or UO_911 (O_911,N_13156,N_13066);
nor UO_912 (O_912,N_13316,N_12192);
nor UO_913 (O_913,N_13961,N_13691);
nand UO_914 (O_914,N_13544,N_12554);
or UO_915 (O_915,N_12081,N_13489);
xnor UO_916 (O_916,N_14810,N_13416);
nand UO_917 (O_917,N_14531,N_14750);
nor UO_918 (O_918,N_13077,N_13851);
nor UO_919 (O_919,N_13574,N_12072);
nor UO_920 (O_920,N_13578,N_13444);
and UO_921 (O_921,N_12225,N_13222);
and UO_922 (O_922,N_14804,N_14443);
nand UO_923 (O_923,N_12602,N_12771);
nand UO_924 (O_924,N_14289,N_13067);
xnor UO_925 (O_925,N_13694,N_12398);
and UO_926 (O_926,N_12418,N_12637);
and UO_927 (O_927,N_14970,N_12167);
or UO_928 (O_928,N_14718,N_14571);
and UO_929 (O_929,N_14790,N_13584);
or UO_930 (O_930,N_13194,N_14177);
or UO_931 (O_931,N_12220,N_12380);
and UO_932 (O_932,N_14551,N_12019);
or UO_933 (O_933,N_14919,N_14140);
nor UO_934 (O_934,N_12457,N_12428);
nand UO_935 (O_935,N_13736,N_12976);
nand UO_936 (O_936,N_14056,N_13171);
nand UO_937 (O_937,N_14833,N_14414);
nor UO_938 (O_938,N_14849,N_12314);
or UO_939 (O_939,N_14796,N_14318);
xnor UO_940 (O_940,N_13258,N_14815);
xor UO_941 (O_941,N_14385,N_13215);
nor UO_942 (O_942,N_13934,N_12664);
nor UO_943 (O_943,N_13696,N_14526);
nor UO_944 (O_944,N_13195,N_14044);
and UO_945 (O_945,N_12722,N_14540);
nand UO_946 (O_946,N_12642,N_14877);
nor UO_947 (O_947,N_12579,N_14348);
xor UO_948 (O_948,N_14135,N_13199);
nand UO_949 (O_949,N_12098,N_12308);
nand UO_950 (O_950,N_14050,N_14309);
xor UO_951 (O_951,N_13817,N_14070);
nand UO_952 (O_952,N_12214,N_12629);
and UO_953 (O_953,N_13721,N_14391);
and UO_954 (O_954,N_14736,N_14705);
and UO_955 (O_955,N_13672,N_14029);
xor UO_956 (O_956,N_13612,N_14554);
xor UO_957 (O_957,N_14363,N_14456);
nor UO_958 (O_958,N_14806,N_13700);
nor UO_959 (O_959,N_12273,N_13714);
nor UO_960 (O_960,N_14539,N_13992);
xor UO_961 (O_961,N_12468,N_13229);
and UO_962 (O_962,N_13271,N_14776);
xor UO_963 (O_963,N_13963,N_12929);
or UO_964 (O_964,N_13032,N_14612);
xor UO_965 (O_965,N_13741,N_13647);
nor UO_966 (O_966,N_14863,N_13049);
or UO_967 (O_967,N_12066,N_12122);
xnor UO_968 (O_968,N_14548,N_12879);
nand UO_969 (O_969,N_12087,N_12904);
xnor UO_970 (O_970,N_12751,N_13784);
xor UO_971 (O_971,N_12013,N_13128);
and UO_972 (O_972,N_12037,N_13304);
nand UO_973 (O_973,N_12972,N_12191);
nor UO_974 (O_974,N_14758,N_14791);
xor UO_975 (O_975,N_13897,N_13699);
and UO_976 (O_976,N_14481,N_14700);
nor UO_977 (O_977,N_14657,N_12099);
xnor UO_978 (O_978,N_14164,N_13818);
and UO_979 (O_979,N_13608,N_13127);
and UO_980 (O_980,N_14079,N_12839);
nand UO_981 (O_981,N_14112,N_12202);
nor UO_982 (O_982,N_14409,N_13480);
or UO_983 (O_983,N_14246,N_13196);
or UO_984 (O_984,N_12560,N_12256);
nand UO_985 (O_985,N_14543,N_13185);
and UO_986 (O_986,N_13779,N_14324);
and UO_987 (O_987,N_12873,N_13173);
nor UO_988 (O_988,N_13778,N_12703);
nand UO_989 (O_989,N_13500,N_13558);
nand UO_990 (O_990,N_14512,N_12848);
xnor UO_991 (O_991,N_12195,N_12365);
and UO_992 (O_992,N_13327,N_12110);
nand UO_993 (O_993,N_14670,N_13305);
nand UO_994 (O_994,N_14258,N_12652);
xnor UO_995 (O_995,N_13256,N_13609);
or UO_996 (O_996,N_12624,N_13682);
nor UO_997 (O_997,N_13381,N_14172);
nand UO_998 (O_998,N_12065,N_14108);
and UO_999 (O_999,N_12474,N_13553);
and UO_1000 (O_1000,N_12813,N_13140);
xnor UO_1001 (O_1001,N_12335,N_14708);
or UO_1002 (O_1002,N_13344,N_13708);
and UO_1003 (O_1003,N_12478,N_12592);
nor UO_1004 (O_1004,N_12448,N_14733);
nor UO_1005 (O_1005,N_14430,N_12133);
nor UO_1006 (O_1006,N_13872,N_12907);
or UO_1007 (O_1007,N_14239,N_12189);
nand UO_1008 (O_1008,N_12070,N_13405);
xor UO_1009 (O_1009,N_13296,N_14843);
nand UO_1010 (O_1010,N_12490,N_13358);
nor UO_1011 (O_1011,N_12589,N_13799);
nand UO_1012 (O_1012,N_13909,N_13104);
xnor UO_1013 (O_1013,N_13688,N_14818);
xnor UO_1014 (O_1014,N_14662,N_14196);
xor UO_1015 (O_1015,N_12102,N_13712);
or UO_1016 (O_1016,N_13103,N_12586);
nand UO_1017 (O_1017,N_13206,N_13182);
nand UO_1018 (O_1018,N_14610,N_12304);
and UO_1019 (O_1019,N_14693,N_14520);
xor UO_1020 (O_1020,N_14830,N_13650);
nand UO_1021 (O_1021,N_12889,N_12781);
xor UO_1022 (O_1022,N_13997,N_13485);
or UO_1023 (O_1023,N_13821,N_12142);
nand UO_1024 (O_1024,N_14995,N_13917);
or UO_1025 (O_1025,N_13417,N_12949);
or UO_1026 (O_1026,N_12330,N_12244);
xor UO_1027 (O_1027,N_12553,N_14407);
nand UO_1028 (O_1028,N_12990,N_12792);
nor UO_1029 (O_1029,N_13276,N_12770);
and UO_1030 (O_1030,N_14061,N_14297);
and UO_1031 (O_1031,N_14131,N_13967);
xnor UO_1032 (O_1032,N_14507,N_13117);
nor UO_1033 (O_1033,N_12958,N_14960);
nand UO_1034 (O_1034,N_13627,N_13541);
and UO_1035 (O_1035,N_14608,N_13585);
nor UO_1036 (O_1036,N_14018,N_13295);
nand UO_1037 (O_1037,N_14165,N_14618);
nand UO_1038 (O_1038,N_12891,N_13670);
nand UO_1039 (O_1039,N_13193,N_12715);
and UO_1040 (O_1040,N_12419,N_14875);
and UO_1041 (O_1041,N_14202,N_13102);
xor UO_1042 (O_1042,N_13797,N_12245);
nand UO_1043 (O_1043,N_12640,N_13243);
nor UO_1044 (O_1044,N_12056,N_13634);
nand UO_1045 (O_1045,N_13369,N_14544);
nor UO_1046 (O_1046,N_12228,N_14354);
nand UO_1047 (O_1047,N_14594,N_13324);
and UO_1048 (O_1048,N_12937,N_14956);
and UO_1049 (O_1049,N_13746,N_13107);
xnor UO_1050 (O_1050,N_14035,N_14349);
nor UO_1051 (O_1051,N_13879,N_12239);
or UO_1052 (O_1052,N_12493,N_14130);
nand UO_1053 (O_1053,N_12160,N_12661);
or UO_1054 (O_1054,N_14499,N_14817);
nand UO_1055 (O_1055,N_12809,N_12728);
and UO_1056 (O_1056,N_13886,N_14648);
or UO_1057 (O_1057,N_13924,N_13908);
nor UO_1058 (O_1058,N_13858,N_12143);
nor UO_1059 (O_1059,N_12970,N_14492);
nand UO_1060 (O_1060,N_13989,N_12203);
nor UO_1061 (O_1061,N_13043,N_13331);
and UO_1062 (O_1062,N_14906,N_14683);
nand UO_1063 (O_1063,N_14222,N_12126);
nor UO_1064 (O_1064,N_14703,N_13548);
nor UO_1065 (O_1065,N_12527,N_14187);
nor UO_1066 (O_1066,N_12178,N_12585);
and UO_1067 (O_1067,N_13224,N_13167);
nor UO_1068 (O_1068,N_12200,N_12346);
nor UO_1069 (O_1069,N_14100,N_13281);
or UO_1070 (O_1070,N_13887,N_12865);
nor UO_1071 (O_1071,N_13881,N_13982);
nand UO_1072 (O_1072,N_14215,N_13648);
or UO_1073 (O_1073,N_14452,N_13024);
and UO_1074 (O_1074,N_13550,N_13105);
or UO_1075 (O_1075,N_12685,N_14926);
and UO_1076 (O_1076,N_12777,N_12074);
xor UO_1077 (O_1077,N_13738,N_12283);
nand UO_1078 (O_1078,N_14482,N_13014);
xor UO_1079 (O_1079,N_13026,N_13618);
nand UO_1080 (O_1080,N_12462,N_14077);
xor UO_1081 (O_1081,N_14702,N_14831);
nand UO_1082 (O_1082,N_12084,N_14730);
nor UO_1083 (O_1083,N_14898,N_14749);
nor UO_1084 (O_1084,N_12109,N_14036);
nand UO_1085 (O_1085,N_12613,N_14424);
or UO_1086 (O_1086,N_12501,N_12495);
xor UO_1087 (O_1087,N_14126,N_13407);
and UO_1088 (O_1088,N_14856,N_13230);
and UO_1089 (O_1089,N_13603,N_13772);
or UO_1090 (O_1090,N_12232,N_14828);
nor UO_1091 (O_1091,N_13981,N_12757);
or UO_1092 (O_1092,N_14225,N_13804);
xnor UO_1093 (O_1093,N_14003,N_14437);
nor UO_1094 (O_1094,N_14290,N_14117);
xor UO_1095 (O_1095,N_13498,N_12638);
nor UO_1096 (O_1096,N_12779,N_14008);
nand UO_1097 (O_1097,N_13777,N_12772);
nand UO_1098 (O_1098,N_13476,N_12590);
or UO_1099 (O_1099,N_14704,N_14192);
and UO_1100 (O_1100,N_12184,N_14547);
or UO_1101 (O_1101,N_14932,N_13725);
nand UO_1102 (O_1102,N_14466,N_14725);
nor UO_1103 (O_1103,N_12597,N_14486);
or UO_1104 (O_1104,N_12651,N_13796);
and UO_1105 (O_1105,N_12568,N_13070);
nor UO_1106 (O_1106,N_14427,N_13260);
nor UO_1107 (O_1107,N_14668,N_12209);
or UO_1108 (O_1108,N_12026,N_14761);
xnor UO_1109 (O_1109,N_14248,N_13630);
and UO_1110 (O_1110,N_12646,N_12443);
xor UO_1111 (O_1111,N_12403,N_13787);
and UO_1112 (O_1112,N_12345,N_14021);
nand UO_1113 (O_1113,N_13488,N_13687);
and UO_1114 (O_1114,N_13715,N_13152);
xnor UO_1115 (O_1115,N_14666,N_13137);
xnor UO_1116 (O_1116,N_14568,N_14509);
nor UO_1117 (O_1117,N_13973,N_12480);
and UO_1118 (O_1118,N_14845,N_12633);
or UO_1119 (O_1119,N_12172,N_14634);
nor UO_1120 (O_1120,N_13435,N_14300);
xnor UO_1121 (O_1121,N_12139,N_14590);
nand UO_1122 (O_1122,N_12123,N_12500);
nand UO_1123 (O_1123,N_14679,N_12546);
and UO_1124 (O_1124,N_13040,N_14519);
xor UO_1125 (O_1125,N_14844,N_14840);
nor UO_1126 (O_1126,N_14878,N_12455);
nand UO_1127 (O_1127,N_12774,N_14422);
nor UO_1128 (O_1128,N_13087,N_14098);
nor UO_1129 (O_1129,N_12504,N_14298);
nor UO_1130 (O_1130,N_12379,N_14595);
and UO_1131 (O_1131,N_13701,N_12947);
and UO_1132 (O_1132,N_14914,N_13284);
nor UO_1133 (O_1133,N_13695,N_13834);
nand UO_1134 (O_1134,N_14566,N_14161);
or UO_1135 (O_1135,N_14173,N_14107);
nor UO_1136 (O_1136,N_12005,N_13802);
xnor UO_1137 (O_1137,N_13086,N_13450);
or UO_1138 (O_1138,N_13427,N_14582);
nand UO_1139 (O_1139,N_12284,N_12783);
xor UO_1140 (O_1140,N_12378,N_13604);
nor UO_1141 (O_1141,N_13554,N_14058);
nor UO_1142 (O_1142,N_13269,N_14396);
xnor UO_1143 (O_1143,N_13564,N_12437);
and UO_1144 (O_1144,N_14230,N_12386);
xnor UO_1145 (O_1145,N_14199,N_14418);
xor UO_1146 (O_1146,N_12615,N_12224);
nand UO_1147 (O_1147,N_12210,N_14737);
or UO_1148 (O_1148,N_12329,N_12838);
xor UO_1149 (O_1149,N_12485,N_12600);
or UO_1150 (O_1150,N_13637,N_13261);
nor UO_1151 (O_1151,N_13439,N_12009);
nor UO_1152 (O_1152,N_13502,N_13906);
and UO_1153 (O_1153,N_12999,N_12130);
and UO_1154 (O_1154,N_12441,N_14557);
or UO_1155 (O_1155,N_14742,N_14375);
nand UO_1156 (O_1156,N_13730,N_14706);
xnor UO_1157 (O_1157,N_13181,N_12237);
xnor UO_1158 (O_1158,N_13889,N_14847);
nor UO_1159 (O_1159,N_12464,N_13180);
and UO_1160 (O_1160,N_14256,N_14756);
nor UO_1161 (O_1161,N_14998,N_13678);
nand UO_1162 (O_1162,N_12973,N_13111);
nand UO_1163 (O_1163,N_14208,N_13050);
xnor UO_1164 (O_1164,N_14550,N_14149);
and UO_1165 (O_1165,N_14360,N_14425);
nand UO_1166 (O_1166,N_13109,N_12675);
and UO_1167 (O_1167,N_13471,N_12364);
nor UO_1168 (O_1168,N_13290,N_14809);
nand UO_1169 (O_1169,N_13303,N_14734);
nor UO_1170 (O_1170,N_12796,N_12351);
nor UO_1171 (O_1171,N_14017,N_13745);
nand UO_1172 (O_1172,N_13250,N_14439);
nand UO_1173 (O_1173,N_12564,N_14382);
nor UO_1174 (O_1174,N_13220,N_14162);
nor UO_1175 (O_1175,N_12628,N_12752);
nand UO_1176 (O_1176,N_13995,N_13980);
and UO_1177 (O_1177,N_12201,N_12294);
nor UO_1178 (O_1178,N_14694,N_13113);
or UO_1179 (O_1179,N_13576,N_12058);
nor UO_1180 (O_1180,N_12282,N_14824);
nand UO_1181 (O_1181,N_12446,N_12235);
nor UO_1182 (O_1182,N_13786,N_12331);
nor UO_1183 (O_1183,N_13160,N_13519);
nor UO_1184 (O_1184,N_12135,N_12510);
and UO_1185 (O_1185,N_13996,N_14455);
or UO_1186 (O_1186,N_14356,N_14139);
nor UO_1187 (O_1187,N_13238,N_14972);
or UO_1188 (O_1188,N_14178,N_12054);
and UO_1189 (O_1189,N_13873,N_14460);
or UO_1190 (O_1190,N_12392,N_14218);
xnor UO_1191 (O_1191,N_12622,N_14819);
or UO_1192 (O_1192,N_12928,N_12050);
nand UO_1193 (O_1193,N_12311,N_14182);
xnor UO_1194 (O_1194,N_12186,N_12701);
nor UO_1195 (O_1195,N_12486,N_14001);
or UO_1196 (O_1196,N_13954,N_13888);
or UO_1197 (O_1197,N_13826,N_14767);
and UO_1198 (O_1198,N_12422,N_13878);
and UO_1199 (O_1199,N_14102,N_13345);
nand UO_1200 (O_1200,N_13711,N_13012);
or UO_1201 (O_1201,N_13566,N_12045);
nand UO_1202 (O_1202,N_12921,N_14432);
or UO_1203 (O_1203,N_13542,N_13496);
xor UO_1204 (O_1204,N_12672,N_12574);
and UO_1205 (O_1205,N_12006,N_13794);
nor UO_1206 (O_1206,N_13705,N_13097);
nor UO_1207 (O_1207,N_14096,N_13632);
nand UO_1208 (O_1208,N_13610,N_12374);
xor UO_1209 (O_1209,N_13468,N_14603);
nand UO_1210 (O_1210,N_14515,N_13822);
nor UO_1211 (O_1211,N_14024,N_12320);
nand UO_1212 (O_1212,N_14002,N_12405);
and UO_1213 (O_1213,N_13398,N_13121);
nor UO_1214 (O_1214,N_14983,N_13571);
or UO_1215 (O_1215,N_14339,N_12181);
xor UO_1216 (O_1216,N_13552,N_12488);
or UO_1217 (O_1217,N_14312,N_12911);
nand UO_1218 (O_1218,N_12154,N_14194);
nor UO_1219 (O_1219,N_14760,N_12782);
and UO_1220 (O_1220,N_14038,N_14366);
nor UO_1221 (O_1221,N_14271,N_14984);
nor UO_1222 (O_1222,N_13782,N_12439);
xor UO_1223 (O_1223,N_12473,N_14404);
and UO_1224 (O_1224,N_13942,N_12327);
xor UO_1225 (O_1225,N_14546,N_12025);
nor UO_1226 (O_1226,N_13943,N_12966);
nor UO_1227 (O_1227,N_13002,N_12269);
and UO_1228 (O_1228,N_12226,N_12402);
and UO_1229 (O_1229,N_12373,N_13685);
nand UO_1230 (O_1230,N_14753,N_14084);
and UO_1231 (O_1231,N_13394,N_13780);
nor UO_1232 (O_1232,N_14498,N_14805);
nor UO_1233 (O_1233,N_14684,N_14254);
and UO_1234 (O_1234,N_13868,N_13783);
and UO_1235 (O_1235,N_12348,N_12017);
and UO_1236 (O_1236,N_13482,N_13894);
or UO_1237 (O_1237,N_13823,N_13523);
xnor UO_1238 (O_1238,N_14155,N_12916);
xor UO_1239 (O_1239,N_12666,N_12219);
xor UO_1240 (O_1240,N_13857,N_12263);
and UO_1241 (O_1241,N_14596,N_14609);
and UO_1242 (O_1242,N_12986,N_12295);
nor UO_1243 (O_1243,N_12061,N_13619);
nor UO_1244 (O_1244,N_14552,N_12940);
nor UO_1245 (O_1245,N_12903,N_14421);
or UO_1246 (O_1246,N_12193,N_13559);
nand UO_1247 (O_1247,N_13112,N_14587);
or UO_1248 (O_1248,N_13466,N_14616);
nor UO_1249 (O_1249,N_14428,N_13091);
nand UO_1250 (O_1250,N_14257,N_13788);
nor UO_1251 (O_1251,N_13800,N_12475);
xor UO_1252 (O_1252,N_13847,N_12847);
xor UO_1253 (O_1253,N_14577,N_12667);
and UO_1254 (O_1254,N_14497,N_14398);
nand UO_1255 (O_1255,N_14219,N_12229);
xor UO_1256 (O_1256,N_13334,N_13940);
nor UO_1257 (O_1257,N_12091,N_12596);
xnor UO_1258 (O_1258,N_13311,N_13089);
or UO_1259 (O_1259,N_12253,N_14525);
nand UO_1260 (O_1260,N_13013,N_14665);
or UO_1261 (O_1261,N_12608,N_14201);
and UO_1262 (O_1262,N_13175,N_14902);
or UO_1263 (O_1263,N_13068,N_13188);
and UO_1264 (O_1264,N_13748,N_12627);
and UO_1265 (O_1265,N_12073,N_13015);
nand UO_1266 (O_1266,N_14223,N_13288);
and UO_1267 (O_1267,N_13546,N_12162);
nor UO_1268 (O_1268,N_12816,N_13301);
xor UO_1269 (O_1269,N_14412,N_12988);
xnor UO_1270 (O_1270,N_12639,N_13551);
nand UO_1271 (O_1271,N_14630,N_14911);
nand UO_1272 (O_1272,N_12416,N_12593);
nand UO_1273 (O_1273,N_12399,N_14782);
and UO_1274 (O_1274,N_13490,N_14602);
and UO_1275 (O_1275,N_14476,N_14558);
and UO_1276 (O_1276,N_12725,N_12460);
nor UO_1277 (O_1277,N_13759,N_12103);
or UO_1278 (O_1278,N_13754,N_14862);
or UO_1279 (O_1279,N_13939,N_14895);
nand UO_1280 (O_1280,N_14381,N_12923);
or UO_1281 (O_1281,N_12170,N_13526);
xor UO_1282 (O_1282,N_13364,N_14245);
nand UO_1283 (O_1283,N_14376,N_13836);
and UO_1284 (O_1284,N_12963,N_13072);
or UO_1285 (O_1285,N_13573,N_13178);
nand UO_1286 (O_1286,N_13306,N_12445);
or UO_1287 (O_1287,N_13249,N_14903);
xor UO_1288 (O_1288,N_14311,N_12031);
and UO_1289 (O_1289,N_14447,N_13970);
nor UO_1290 (O_1290,N_14011,N_14395);
nand UO_1291 (O_1291,N_12198,N_13801);
nand UO_1292 (O_1292,N_14209,N_12002);
or UO_1293 (O_1293,N_12521,N_12815);
and UO_1294 (O_1294,N_12975,N_14119);
or UO_1295 (O_1295,N_13209,N_12136);
xor UO_1296 (O_1296,N_12580,N_12151);
nand UO_1297 (O_1297,N_14091,N_14374);
and UO_1298 (O_1298,N_12360,N_13877);
and UO_1299 (O_1299,N_12372,N_12953);
or UO_1300 (O_1300,N_14049,N_14945);
xor UO_1301 (O_1301,N_14252,N_12823);
nand UO_1302 (O_1302,N_14707,N_12822);
xor UO_1303 (O_1303,N_12872,N_13975);
and UO_1304 (O_1304,N_12350,N_13169);
or UO_1305 (O_1305,N_13907,N_14442);
nor UO_1306 (O_1306,N_14560,N_13264);
xor UO_1307 (O_1307,N_13859,N_14171);
nand UO_1308 (O_1308,N_13469,N_14765);
nor UO_1309 (O_1309,N_14658,N_12764);
nand UO_1310 (O_1310,N_13473,N_13445);
nand UO_1311 (O_1311,N_14288,N_12804);
nor UO_1312 (O_1312,N_13757,N_13710);
xor UO_1313 (O_1313,N_13891,N_12761);
or UO_1314 (O_1314,N_14740,N_13307);
or UO_1315 (O_1315,N_14576,N_13723);
and UO_1316 (O_1316,N_14328,N_14440);
xnor UO_1317 (O_1317,N_12884,N_14154);
nand UO_1318 (O_1318,N_13234,N_14813);
nor UO_1319 (O_1319,N_12682,N_14495);
nand UO_1320 (O_1320,N_12788,N_14390);
or UO_1321 (O_1321,N_14677,N_12810);
and UO_1322 (O_1322,N_14244,N_12499);
nand UO_1323 (O_1323,N_14226,N_14242);
or UO_1324 (O_1324,N_14864,N_12265);
nand UO_1325 (O_1325,N_13487,N_14584);
nand UO_1326 (O_1326,N_13862,N_14022);
nand UO_1327 (O_1327,N_14754,N_13719);
nand UO_1328 (O_1328,N_12739,N_14332);
xnor UO_1329 (O_1329,N_14157,N_12868);
or UO_1330 (O_1330,N_13964,N_12401);
and UO_1331 (O_1331,N_12288,N_12431);
and UO_1332 (O_1332,N_13241,N_14127);
nand UO_1333 (O_1333,N_13586,N_12614);
xor UO_1334 (O_1334,N_12995,N_12825);
or UO_1335 (O_1335,N_13497,N_14803);
nand UO_1336 (O_1336,N_14040,N_14592);
xor UO_1337 (O_1337,N_13090,N_13825);
and UO_1338 (O_1338,N_14743,N_12095);
nor UO_1339 (O_1339,N_14959,N_12997);
xnor UO_1340 (O_1340,N_12254,N_13198);
nor UO_1341 (O_1341,N_12833,N_14188);
and UO_1342 (O_1342,N_13136,N_12705);
or UO_1343 (O_1343,N_12036,N_13587);
xnor UO_1344 (O_1344,N_12826,N_14620);
nand UO_1345 (O_1345,N_13309,N_12434);
and UO_1346 (O_1346,N_14401,N_13280);
or UO_1347 (O_1347,N_14953,N_13410);
nor UO_1348 (O_1348,N_13071,N_13671);
xor UO_1349 (O_1349,N_14785,N_12021);
xnor UO_1350 (O_1350,N_12491,N_14479);
nor UO_1351 (O_1351,N_13895,N_14379);
xnor UO_1352 (O_1352,N_13953,N_12861);
nor UO_1353 (O_1353,N_14369,N_13454);
and UO_1354 (O_1354,N_14496,N_14181);
nand UO_1355 (O_1355,N_14299,N_14846);
and UO_1356 (O_1356,N_12736,N_13508);
xor UO_1357 (O_1357,N_13494,N_13007);
nor UO_1358 (O_1358,N_12730,N_12027);
and UO_1359 (O_1359,N_13876,N_14826);
xnor UO_1360 (O_1360,N_12053,N_13424);
and UO_1361 (O_1361,N_12619,N_14060);
or UO_1362 (O_1362,N_13179,N_14942);
and UO_1363 (O_1363,N_14039,N_12332);
or UO_1364 (O_1364,N_12989,N_13543);
nor UO_1365 (O_1365,N_12699,N_12340);
and UO_1366 (O_1366,N_12114,N_13655);
nor UO_1367 (O_1367,N_12303,N_14764);
and UO_1368 (O_1368,N_14731,N_13581);
nor UO_1369 (O_1369,N_14837,N_12395);
xnor UO_1370 (O_1370,N_13968,N_14264);
or UO_1371 (O_1371,N_14176,N_14449);
or UO_1372 (O_1372,N_12931,N_12299);
nand UO_1373 (O_1373,N_13231,N_12479);
nand UO_1374 (O_1374,N_12503,N_12349);
nand UO_1375 (O_1375,N_13912,N_13986);
xor UO_1376 (O_1376,N_13421,N_14259);
nor UO_1377 (O_1377,N_13933,N_14642);
or UO_1378 (O_1378,N_12400,N_12394);
nor UO_1379 (O_1379,N_14669,N_12250);
nor UO_1380 (O_1380,N_12819,N_13223);
or UO_1381 (O_1381,N_13537,N_12029);
and UO_1382 (O_1382,N_13567,N_12994);
and UO_1383 (O_1383,N_12737,N_14969);
nand UO_1384 (O_1384,N_14251,N_13623);
nand UO_1385 (O_1385,N_12727,N_13479);
and UO_1386 (O_1386,N_13948,N_12341);
xnor UO_1387 (O_1387,N_14081,N_13098);
and UO_1388 (O_1388,N_12376,N_12753);
nor UO_1389 (O_1389,N_12820,N_14585);
or UO_1390 (O_1390,N_14755,N_14717);
and UO_1391 (O_1391,N_13207,N_14533);
or UO_1392 (O_1392,N_13096,N_14860);
or UO_1393 (O_1393,N_12754,N_13449);
nand UO_1394 (O_1394,N_14464,N_12939);
and UO_1395 (O_1395,N_14046,N_12668);
and UO_1396 (O_1396,N_13903,N_14141);
xnor UO_1397 (O_1397,N_12430,N_14788);
nand UO_1398 (O_1398,N_14981,N_12925);
nand UO_1399 (O_1399,N_12723,N_12974);
and UO_1400 (O_1400,N_14559,N_14445);
xor UO_1401 (O_1401,N_12359,N_12707);
nand UO_1402 (O_1402,N_12190,N_14726);
nand UO_1403 (O_1403,N_12471,N_14820);
nor UO_1404 (O_1404,N_12052,N_13720);
nand UO_1405 (O_1405,N_12141,N_12658);
nor UO_1406 (O_1406,N_12565,N_13338);
xor UO_1407 (O_1407,N_13452,N_14632);
and UO_1408 (O_1408,N_13579,N_12447);
or UO_1409 (O_1409,N_13768,N_12173);
xnor UO_1410 (O_1410,N_14279,N_12530);
xor UO_1411 (O_1411,N_12914,N_13814);
or UO_1412 (O_1412,N_12880,N_14285);
nand UO_1413 (O_1413,N_12599,N_14231);
xor UO_1414 (O_1414,N_14651,N_13413);
and UO_1415 (O_1415,N_14380,N_14101);
and UO_1416 (O_1416,N_14947,N_14884);
nand UO_1417 (O_1417,N_12456,N_12290);
or UO_1418 (O_1418,N_12743,N_13210);
nand UO_1419 (O_1419,N_12969,N_12440);
and UO_1420 (O_1420,N_14361,N_12520);
and UO_1421 (O_1421,N_12089,N_13731);
or UO_1422 (O_1422,N_14617,N_14992);
xor UO_1423 (O_1423,N_13674,N_13484);
xnor UO_1424 (O_1424,N_14952,N_13125);
or UO_1425 (O_1425,N_14948,N_12670);
nand UO_1426 (O_1426,N_13689,N_12979);
nor UO_1427 (O_1427,N_12231,N_14832);
nand UO_1428 (O_1428,N_12124,N_14732);
and UO_1429 (O_1429,N_14277,N_12371);
nand UO_1430 (O_1430,N_13099,N_12616);
or UO_1431 (O_1431,N_14494,N_14063);
xnor UO_1432 (O_1432,N_14287,N_14802);
nand UO_1433 (O_1433,N_12626,N_14581);
nand UO_1434 (O_1434,N_13622,N_12075);
or UO_1435 (O_1435,N_14958,N_13808);
xnor UO_1436 (O_1436,N_14307,N_14007);
or UO_1437 (O_1437,N_14744,N_14453);
nor UO_1438 (O_1438,N_14278,N_14939);
nor UO_1439 (O_1439,N_14160,N_13505);
xnor UO_1440 (O_1440,N_12281,N_12797);
nor UO_1441 (O_1441,N_14317,N_14241);
nand UO_1442 (O_1442,N_12085,N_12780);
nor UO_1443 (O_1443,N_13035,N_14148);
xnor UO_1444 (O_1444,N_13983,N_14784);
or UO_1445 (O_1445,N_13093,N_12962);
nor UO_1446 (O_1446,N_12852,N_12252);
or UO_1447 (O_1447,N_13890,N_12138);
xor UO_1448 (O_1448,N_12595,N_13108);
xor UO_1449 (O_1449,N_13337,N_14370);
xnor UO_1450 (O_1450,N_13845,N_13591);
or UO_1451 (O_1451,N_14701,N_12309);
nor UO_1452 (O_1452,N_14338,N_13247);
nor UO_1453 (O_1453,N_12157,N_14014);
and UO_1454 (O_1454,N_13265,N_14406);
or UO_1455 (O_1455,N_12573,N_12097);
or UO_1456 (O_1456,N_13668,N_12583);
or UO_1457 (O_1457,N_13168,N_12505);
nor UO_1458 (O_1458,N_13400,N_14619);
nand UO_1459 (O_1459,N_12472,N_12575);
or UO_1460 (O_1460,N_13861,N_12522);
and UO_1461 (O_1461,N_14766,N_12152);
xnor UO_1462 (O_1462,N_14503,N_13643);
xnor UO_1463 (O_1463,N_13499,N_12307);
or UO_1464 (O_1464,N_13849,N_13640);
or UO_1465 (O_1465,N_13082,N_12397);
and UO_1466 (O_1466,N_12132,N_12068);
nor UO_1467 (O_1467,N_14841,N_14216);
and UO_1468 (O_1468,N_12208,N_14235);
or UO_1469 (O_1469,N_13457,N_12354);
xnor UO_1470 (O_1470,N_14675,N_13520);
or UO_1471 (O_1471,N_14990,N_13838);
xnor UO_1472 (O_1472,N_12155,N_12738);
and UO_1473 (O_1473,N_12905,N_12370);
nor UO_1474 (O_1474,N_14344,N_12875);
nor UO_1475 (O_1475,N_13549,N_12454);
nand UO_1476 (O_1476,N_12541,N_13474);
or UO_1477 (O_1477,N_12449,N_13286);
nand UO_1478 (O_1478,N_12840,N_12563);
or UO_1479 (O_1479,N_13615,N_12687);
nand UO_1480 (O_1480,N_12247,N_13390);
nand UO_1481 (O_1481,N_13116,N_13403);
nand UO_1482 (O_1482,N_13555,N_14579);
nor UO_1483 (O_1483,N_14082,N_13824);
nor UO_1484 (O_1484,N_12104,N_12306);
or UO_1485 (O_1485,N_14988,N_14857);
xor UO_1486 (O_1486,N_13880,N_14541);
nand UO_1487 (O_1487,N_12057,N_13565);
nor UO_1488 (O_1488,N_13213,N_12683);
nor UO_1489 (O_1489,N_13461,N_13060);
nand UO_1490 (O_1490,N_13019,N_13315);
xnor UO_1491 (O_1491,N_14068,N_14415);
and UO_1492 (O_1492,N_14690,N_13793);
nand UO_1493 (O_1493,N_12955,N_12708);
xor UO_1494 (O_1494,N_12175,N_12718);
nor UO_1495 (O_1495,N_12620,N_12870);
nor UO_1496 (O_1496,N_14622,N_14545);
xor UO_1497 (O_1497,N_14599,N_12113);
nand UO_1498 (O_1498,N_13790,N_13959);
xnor UO_1499 (O_1499,N_12984,N_14916);
nand UO_1500 (O_1500,N_14871,N_14145);
nor UO_1501 (O_1501,N_12487,N_13412);
xor UO_1502 (O_1502,N_13670,N_12205);
and UO_1503 (O_1503,N_14097,N_12150);
or UO_1504 (O_1504,N_13090,N_12073);
xor UO_1505 (O_1505,N_13359,N_12348);
xor UO_1506 (O_1506,N_12180,N_14204);
xor UO_1507 (O_1507,N_13209,N_14024);
nor UO_1508 (O_1508,N_13134,N_12472);
or UO_1509 (O_1509,N_13809,N_12629);
nor UO_1510 (O_1510,N_14956,N_12855);
and UO_1511 (O_1511,N_12463,N_12675);
or UO_1512 (O_1512,N_13291,N_12178);
nand UO_1513 (O_1513,N_14993,N_13224);
nand UO_1514 (O_1514,N_13616,N_12245);
nand UO_1515 (O_1515,N_13143,N_12277);
or UO_1516 (O_1516,N_12369,N_13804);
and UO_1517 (O_1517,N_12304,N_12624);
or UO_1518 (O_1518,N_12745,N_14271);
and UO_1519 (O_1519,N_13442,N_14845);
and UO_1520 (O_1520,N_14425,N_14539);
and UO_1521 (O_1521,N_12635,N_14699);
or UO_1522 (O_1522,N_14348,N_12787);
or UO_1523 (O_1523,N_12079,N_14220);
xor UO_1524 (O_1524,N_13934,N_13229);
or UO_1525 (O_1525,N_12929,N_14045);
nand UO_1526 (O_1526,N_12626,N_12318);
nor UO_1527 (O_1527,N_13643,N_14464);
xor UO_1528 (O_1528,N_14571,N_14271);
or UO_1529 (O_1529,N_13683,N_12687);
nor UO_1530 (O_1530,N_13150,N_12816);
xor UO_1531 (O_1531,N_14850,N_14011);
or UO_1532 (O_1532,N_14887,N_14712);
nor UO_1533 (O_1533,N_13149,N_14800);
or UO_1534 (O_1534,N_12819,N_14516);
nor UO_1535 (O_1535,N_13078,N_12448);
xnor UO_1536 (O_1536,N_14306,N_14101);
or UO_1537 (O_1537,N_13334,N_14580);
nor UO_1538 (O_1538,N_14045,N_12526);
or UO_1539 (O_1539,N_12925,N_14393);
xnor UO_1540 (O_1540,N_12118,N_14674);
nand UO_1541 (O_1541,N_12906,N_12983);
nand UO_1542 (O_1542,N_14962,N_13039);
nor UO_1543 (O_1543,N_13048,N_13460);
nand UO_1544 (O_1544,N_13462,N_14654);
nor UO_1545 (O_1545,N_13201,N_13788);
nand UO_1546 (O_1546,N_14636,N_13666);
and UO_1547 (O_1547,N_12239,N_12924);
and UO_1548 (O_1548,N_14681,N_13652);
nor UO_1549 (O_1549,N_13285,N_13242);
or UO_1550 (O_1550,N_14510,N_12345);
nor UO_1551 (O_1551,N_13145,N_14227);
or UO_1552 (O_1552,N_13659,N_12081);
xor UO_1553 (O_1553,N_12458,N_14929);
or UO_1554 (O_1554,N_14212,N_12232);
xor UO_1555 (O_1555,N_12701,N_13908);
or UO_1556 (O_1556,N_12586,N_14831);
xor UO_1557 (O_1557,N_14159,N_13082);
xnor UO_1558 (O_1558,N_14773,N_13610);
nand UO_1559 (O_1559,N_12990,N_14575);
and UO_1560 (O_1560,N_13307,N_12855);
or UO_1561 (O_1561,N_14598,N_12196);
or UO_1562 (O_1562,N_14580,N_14443);
nand UO_1563 (O_1563,N_12470,N_13063);
or UO_1564 (O_1564,N_12106,N_13269);
or UO_1565 (O_1565,N_14227,N_13850);
nand UO_1566 (O_1566,N_14835,N_13102);
nor UO_1567 (O_1567,N_12611,N_14239);
and UO_1568 (O_1568,N_12757,N_13457);
or UO_1569 (O_1569,N_14314,N_14792);
xor UO_1570 (O_1570,N_14509,N_14277);
xor UO_1571 (O_1571,N_12455,N_14845);
and UO_1572 (O_1572,N_13262,N_12837);
or UO_1573 (O_1573,N_14169,N_13603);
nor UO_1574 (O_1574,N_12199,N_12806);
and UO_1575 (O_1575,N_13375,N_12596);
and UO_1576 (O_1576,N_14294,N_13535);
and UO_1577 (O_1577,N_12849,N_13385);
or UO_1578 (O_1578,N_13297,N_13678);
or UO_1579 (O_1579,N_12541,N_12269);
or UO_1580 (O_1580,N_12601,N_13731);
and UO_1581 (O_1581,N_14253,N_12103);
xnor UO_1582 (O_1582,N_12316,N_12807);
nand UO_1583 (O_1583,N_13790,N_12647);
and UO_1584 (O_1584,N_14775,N_12812);
nor UO_1585 (O_1585,N_12576,N_12903);
and UO_1586 (O_1586,N_12403,N_13194);
and UO_1587 (O_1587,N_13099,N_12372);
nor UO_1588 (O_1588,N_14805,N_14303);
nor UO_1589 (O_1589,N_13760,N_13889);
nor UO_1590 (O_1590,N_12856,N_14048);
and UO_1591 (O_1591,N_14514,N_14807);
nor UO_1592 (O_1592,N_13228,N_13569);
nor UO_1593 (O_1593,N_13997,N_13483);
xnor UO_1594 (O_1594,N_13885,N_13056);
nor UO_1595 (O_1595,N_14884,N_13047);
or UO_1596 (O_1596,N_12263,N_13545);
and UO_1597 (O_1597,N_14643,N_12693);
or UO_1598 (O_1598,N_12352,N_12231);
and UO_1599 (O_1599,N_14323,N_12055);
or UO_1600 (O_1600,N_13607,N_12659);
xnor UO_1601 (O_1601,N_12979,N_14923);
xnor UO_1602 (O_1602,N_14236,N_13188);
nor UO_1603 (O_1603,N_12841,N_14732);
or UO_1604 (O_1604,N_14281,N_12111);
nor UO_1605 (O_1605,N_13068,N_12615);
nor UO_1606 (O_1606,N_12792,N_14856);
nor UO_1607 (O_1607,N_13423,N_12204);
nor UO_1608 (O_1608,N_14905,N_12207);
nor UO_1609 (O_1609,N_14082,N_12368);
xor UO_1610 (O_1610,N_14727,N_13219);
nor UO_1611 (O_1611,N_14116,N_12575);
xor UO_1612 (O_1612,N_12540,N_13165);
nand UO_1613 (O_1613,N_13618,N_12662);
and UO_1614 (O_1614,N_12153,N_14663);
and UO_1615 (O_1615,N_13653,N_14056);
nand UO_1616 (O_1616,N_14573,N_14517);
and UO_1617 (O_1617,N_12999,N_12696);
or UO_1618 (O_1618,N_14201,N_13796);
nand UO_1619 (O_1619,N_13705,N_13603);
xnor UO_1620 (O_1620,N_14934,N_12423);
xnor UO_1621 (O_1621,N_12498,N_12063);
or UO_1622 (O_1622,N_12665,N_14778);
nor UO_1623 (O_1623,N_14786,N_14084);
and UO_1624 (O_1624,N_14396,N_13600);
xor UO_1625 (O_1625,N_13568,N_14775);
xor UO_1626 (O_1626,N_12042,N_12455);
nor UO_1627 (O_1627,N_14182,N_12356);
or UO_1628 (O_1628,N_14289,N_14448);
or UO_1629 (O_1629,N_13870,N_12564);
nor UO_1630 (O_1630,N_14539,N_14668);
and UO_1631 (O_1631,N_13136,N_14762);
and UO_1632 (O_1632,N_14085,N_13567);
or UO_1633 (O_1633,N_12590,N_12328);
and UO_1634 (O_1634,N_13398,N_13109);
xnor UO_1635 (O_1635,N_13040,N_14488);
xor UO_1636 (O_1636,N_13033,N_12191);
and UO_1637 (O_1637,N_14946,N_12716);
or UO_1638 (O_1638,N_12518,N_13511);
nand UO_1639 (O_1639,N_14223,N_14156);
xor UO_1640 (O_1640,N_12586,N_14651);
nor UO_1641 (O_1641,N_12986,N_14349);
or UO_1642 (O_1642,N_12573,N_13451);
and UO_1643 (O_1643,N_12420,N_12163);
or UO_1644 (O_1644,N_12061,N_12550);
or UO_1645 (O_1645,N_12018,N_14008);
or UO_1646 (O_1646,N_14229,N_12752);
and UO_1647 (O_1647,N_13800,N_14817);
and UO_1648 (O_1648,N_14735,N_14767);
nand UO_1649 (O_1649,N_14364,N_12438);
and UO_1650 (O_1650,N_14628,N_12169);
xor UO_1651 (O_1651,N_13227,N_13929);
or UO_1652 (O_1652,N_13562,N_13179);
or UO_1653 (O_1653,N_13723,N_14187);
or UO_1654 (O_1654,N_13872,N_14132);
nand UO_1655 (O_1655,N_13286,N_12235);
nor UO_1656 (O_1656,N_14725,N_14765);
and UO_1657 (O_1657,N_13578,N_14205);
nand UO_1658 (O_1658,N_13828,N_12522);
nand UO_1659 (O_1659,N_12228,N_12850);
or UO_1660 (O_1660,N_12604,N_13961);
nand UO_1661 (O_1661,N_14972,N_13455);
nor UO_1662 (O_1662,N_12777,N_12350);
nand UO_1663 (O_1663,N_14934,N_14046);
xnor UO_1664 (O_1664,N_14906,N_13970);
and UO_1665 (O_1665,N_14764,N_14600);
nor UO_1666 (O_1666,N_13400,N_14166);
xor UO_1667 (O_1667,N_14157,N_12286);
and UO_1668 (O_1668,N_12331,N_12666);
nor UO_1669 (O_1669,N_13593,N_13779);
or UO_1670 (O_1670,N_12099,N_14204);
nand UO_1671 (O_1671,N_12489,N_13635);
nand UO_1672 (O_1672,N_13829,N_13219);
and UO_1673 (O_1673,N_14210,N_12675);
nor UO_1674 (O_1674,N_12460,N_12058);
xor UO_1675 (O_1675,N_13426,N_12211);
and UO_1676 (O_1676,N_13828,N_14513);
and UO_1677 (O_1677,N_13035,N_14134);
nor UO_1678 (O_1678,N_12775,N_13376);
nor UO_1679 (O_1679,N_13412,N_12712);
nand UO_1680 (O_1680,N_14021,N_14956);
xor UO_1681 (O_1681,N_14079,N_12997);
or UO_1682 (O_1682,N_14509,N_12412);
and UO_1683 (O_1683,N_12329,N_12898);
nand UO_1684 (O_1684,N_13030,N_13564);
xnor UO_1685 (O_1685,N_12442,N_14369);
or UO_1686 (O_1686,N_14412,N_12187);
or UO_1687 (O_1687,N_14745,N_12936);
and UO_1688 (O_1688,N_13045,N_14899);
or UO_1689 (O_1689,N_14720,N_12668);
and UO_1690 (O_1690,N_14670,N_13943);
xnor UO_1691 (O_1691,N_14408,N_12010);
nand UO_1692 (O_1692,N_12551,N_13197);
and UO_1693 (O_1693,N_12294,N_13574);
xor UO_1694 (O_1694,N_13750,N_13865);
xor UO_1695 (O_1695,N_14237,N_12940);
or UO_1696 (O_1696,N_13234,N_12156);
or UO_1697 (O_1697,N_12797,N_13725);
xor UO_1698 (O_1698,N_13434,N_13953);
or UO_1699 (O_1699,N_14589,N_13118);
and UO_1700 (O_1700,N_14677,N_12726);
nor UO_1701 (O_1701,N_13168,N_13558);
or UO_1702 (O_1702,N_13051,N_14509);
nor UO_1703 (O_1703,N_14568,N_14751);
and UO_1704 (O_1704,N_13092,N_12401);
or UO_1705 (O_1705,N_13630,N_12876);
nand UO_1706 (O_1706,N_14785,N_13844);
and UO_1707 (O_1707,N_12548,N_12436);
nor UO_1708 (O_1708,N_14124,N_13785);
or UO_1709 (O_1709,N_14382,N_13259);
nor UO_1710 (O_1710,N_14956,N_14063);
nand UO_1711 (O_1711,N_14190,N_14177);
and UO_1712 (O_1712,N_14831,N_12375);
and UO_1713 (O_1713,N_13554,N_13040);
and UO_1714 (O_1714,N_13939,N_14142);
nor UO_1715 (O_1715,N_13048,N_13386);
nand UO_1716 (O_1716,N_13030,N_14577);
or UO_1717 (O_1717,N_12528,N_14117);
and UO_1718 (O_1718,N_13925,N_14865);
or UO_1719 (O_1719,N_14919,N_13107);
and UO_1720 (O_1720,N_13135,N_14209);
nand UO_1721 (O_1721,N_12308,N_13413);
nor UO_1722 (O_1722,N_13010,N_13339);
xor UO_1723 (O_1723,N_12664,N_14280);
nand UO_1724 (O_1724,N_12182,N_12406);
xnor UO_1725 (O_1725,N_14968,N_12762);
nor UO_1726 (O_1726,N_14555,N_14121);
nor UO_1727 (O_1727,N_12705,N_13324);
nand UO_1728 (O_1728,N_14944,N_12348);
and UO_1729 (O_1729,N_13043,N_13816);
nor UO_1730 (O_1730,N_14226,N_13730);
and UO_1731 (O_1731,N_13705,N_13833);
nand UO_1732 (O_1732,N_14689,N_12921);
nand UO_1733 (O_1733,N_12390,N_13573);
xor UO_1734 (O_1734,N_12016,N_14004);
nand UO_1735 (O_1735,N_12647,N_14819);
nor UO_1736 (O_1736,N_12515,N_13513);
xnor UO_1737 (O_1737,N_13640,N_13176);
nor UO_1738 (O_1738,N_13848,N_13627);
or UO_1739 (O_1739,N_14571,N_12321);
or UO_1740 (O_1740,N_13602,N_13327);
xnor UO_1741 (O_1741,N_12657,N_13026);
nand UO_1742 (O_1742,N_14211,N_12323);
and UO_1743 (O_1743,N_14136,N_13648);
nor UO_1744 (O_1744,N_12152,N_12071);
xor UO_1745 (O_1745,N_14647,N_12670);
or UO_1746 (O_1746,N_13637,N_12142);
nand UO_1747 (O_1747,N_14356,N_13662);
nand UO_1748 (O_1748,N_12095,N_13060);
nand UO_1749 (O_1749,N_13537,N_14818);
nor UO_1750 (O_1750,N_12791,N_12567);
nor UO_1751 (O_1751,N_12879,N_14198);
nor UO_1752 (O_1752,N_13384,N_12932);
xor UO_1753 (O_1753,N_12352,N_12805);
nand UO_1754 (O_1754,N_13227,N_12121);
and UO_1755 (O_1755,N_12353,N_13366);
nor UO_1756 (O_1756,N_12907,N_14947);
nor UO_1757 (O_1757,N_14459,N_12656);
xnor UO_1758 (O_1758,N_13958,N_13002);
xnor UO_1759 (O_1759,N_13128,N_12966);
nand UO_1760 (O_1760,N_12456,N_13214);
or UO_1761 (O_1761,N_13604,N_12538);
and UO_1762 (O_1762,N_13424,N_14285);
and UO_1763 (O_1763,N_14393,N_14046);
or UO_1764 (O_1764,N_13180,N_13047);
nor UO_1765 (O_1765,N_13891,N_13020);
or UO_1766 (O_1766,N_14941,N_14484);
nand UO_1767 (O_1767,N_12332,N_14849);
or UO_1768 (O_1768,N_12474,N_13870);
nand UO_1769 (O_1769,N_14392,N_14831);
nand UO_1770 (O_1770,N_14589,N_12330);
or UO_1771 (O_1771,N_14359,N_14264);
and UO_1772 (O_1772,N_14535,N_13017);
and UO_1773 (O_1773,N_13607,N_14564);
nor UO_1774 (O_1774,N_14103,N_13737);
or UO_1775 (O_1775,N_12357,N_13408);
and UO_1776 (O_1776,N_14072,N_13100);
nand UO_1777 (O_1777,N_14776,N_13000);
nor UO_1778 (O_1778,N_13319,N_13787);
xor UO_1779 (O_1779,N_14180,N_14393);
xnor UO_1780 (O_1780,N_12558,N_14344);
and UO_1781 (O_1781,N_14225,N_13879);
xor UO_1782 (O_1782,N_12084,N_14640);
xnor UO_1783 (O_1783,N_13367,N_14343);
and UO_1784 (O_1784,N_13908,N_13528);
xnor UO_1785 (O_1785,N_13480,N_12362);
nand UO_1786 (O_1786,N_12643,N_14209);
nor UO_1787 (O_1787,N_12563,N_14509);
and UO_1788 (O_1788,N_12193,N_13632);
or UO_1789 (O_1789,N_14290,N_13470);
nor UO_1790 (O_1790,N_14580,N_14674);
or UO_1791 (O_1791,N_12950,N_14659);
nor UO_1792 (O_1792,N_14850,N_12833);
xnor UO_1793 (O_1793,N_14371,N_12437);
nor UO_1794 (O_1794,N_13228,N_12795);
or UO_1795 (O_1795,N_14371,N_13736);
nand UO_1796 (O_1796,N_13380,N_12915);
nor UO_1797 (O_1797,N_13408,N_14291);
or UO_1798 (O_1798,N_14823,N_13740);
and UO_1799 (O_1799,N_12901,N_14468);
nand UO_1800 (O_1800,N_12598,N_14561);
or UO_1801 (O_1801,N_13592,N_14741);
nor UO_1802 (O_1802,N_12355,N_13616);
nand UO_1803 (O_1803,N_13648,N_13888);
nand UO_1804 (O_1804,N_12684,N_14700);
nor UO_1805 (O_1805,N_13228,N_14058);
or UO_1806 (O_1806,N_14389,N_13244);
nand UO_1807 (O_1807,N_14661,N_14262);
and UO_1808 (O_1808,N_12678,N_13947);
or UO_1809 (O_1809,N_14797,N_13193);
nand UO_1810 (O_1810,N_12341,N_14946);
nor UO_1811 (O_1811,N_13127,N_14027);
xor UO_1812 (O_1812,N_14793,N_12463);
nand UO_1813 (O_1813,N_12531,N_12263);
nand UO_1814 (O_1814,N_14053,N_13462);
and UO_1815 (O_1815,N_13807,N_12846);
nand UO_1816 (O_1816,N_14120,N_13498);
and UO_1817 (O_1817,N_12864,N_14593);
xnor UO_1818 (O_1818,N_12115,N_13562);
and UO_1819 (O_1819,N_12055,N_14113);
nand UO_1820 (O_1820,N_13377,N_14354);
and UO_1821 (O_1821,N_14576,N_14458);
nor UO_1822 (O_1822,N_12917,N_12445);
nor UO_1823 (O_1823,N_12607,N_13235);
nor UO_1824 (O_1824,N_12237,N_14402);
nor UO_1825 (O_1825,N_12846,N_12745);
xor UO_1826 (O_1826,N_12407,N_12384);
xor UO_1827 (O_1827,N_14279,N_13923);
xor UO_1828 (O_1828,N_12061,N_14374);
xor UO_1829 (O_1829,N_12875,N_14906);
or UO_1830 (O_1830,N_14258,N_13405);
and UO_1831 (O_1831,N_13417,N_13103);
nor UO_1832 (O_1832,N_14908,N_12044);
and UO_1833 (O_1833,N_14567,N_12875);
nor UO_1834 (O_1834,N_14870,N_13253);
and UO_1835 (O_1835,N_13440,N_12420);
or UO_1836 (O_1836,N_14945,N_13783);
and UO_1837 (O_1837,N_13272,N_14457);
or UO_1838 (O_1838,N_13771,N_14442);
nand UO_1839 (O_1839,N_12190,N_13555);
and UO_1840 (O_1840,N_14127,N_13708);
or UO_1841 (O_1841,N_13876,N_12695);
and UO_1842 (O_1842,N_13694,N_14219);
and UO_1843 (O_1843,N_14981,N_14069);
or UO_1844 (O_1844,N_14858,N_14644);
or UO_1845 (O_1845,N_14069,N_14081);
nor UO_1846 (O_1846,N_13538,N_14683);
nand UO_1847 (O_1847,N_13063,N_12717);
nand UO_1848 (O_1848,N_12101,N_14719);
and UO_1849 (O_1849,N_12716,N_13447);
nand UO_1850 (O_1850,N_13301,N_13075);
xor UO_1851 (O_1851,N_12083,N_12105);
or UO_1852 (O_1852,N_14291,N_13548);
nand UO_1853 (O_1853,N_12717,N_14899);
and UO_1854 (O_1854,N_14217,N_13007);
and UO_1855 (O_1855,N_14782,N_14030);
nand UO_1856 (O_1856,N_12843,N_13130);
nand UO_1857 (O_1857,N_14732,N_14387);
or UO_1858 (O_1858,N_12053,N_13551);
nand UO_1859 (O_1859,N_14188,N_14579);
nand UO_1860 (O_1860,N_14831,N_12689);
nor UO_1861 (O_1861,N_13113,N_14541);
xor UO_1862 (O_1862,N_12366,N_14442);
nand UO_1863 (O_1863,N_14430,N_13532);
nor UO_1864 (O_1864,N_14979,N_13254);
nand UO_1865 (O_1865,N_14199,N_12640);
and UO_1866 (O_1866,N_13318,N_13087);
nand UO_1867 (O_1867,N_12797,N_13480);
nor UO_1868 (O_1868,N_14974,N_12201);
and UO_1869 (O_1869,N_13761,N_13139);
xnor UO_1870 (O_1870,N_12199,N_14890);
xor UO_1871 (O_1871,N_14249,N_12459);
or UO_1872 (O_1872,N_14100,N_13106);
xnor UO_1873 (O_1873,N_13059,N_12163);
xor UO_1874 (O_1874,N_14902,N_13852);
xor UO_1875 (O_1875,N_13102,N_13747);
xor UO_1876 (O_1876,N_14388,N_14018);
or UO_1877 (O_1877,N_14799,N_13314);
xnor UO_1878 (O_1878,N_13349,N_12219);
nor UO_1879 (O_1879,N_13067,N_12259);
nand UO_1880 (O_1880,N_14726,N_14621);
nand UO_1881 (O_1881,N_13081,N_14306);
or UO_1882 (O_1882,N_13920,N_14632);
or UO_1883 (O_1883,N_13420,N_13157);
and UO_1884 (O_1884,N_12063,N_14602);
and UO_1885 (O_1885,N_14168,N_12029);
nand UO_1886 (O_1886,N_13697,N_14119);
or UO_1887 (O_1887,N_13607,N_13427);
xnor UO_1888 (O_1888,N_12427,N_13594);
and UO_1889 (O_1889,N_12248,N_12274);
or UO_1890 (O_1890,N_14141,N_12855);
xor UO_1891 (O_1891,N_13412,N_12671);
nor UO_1892 (O_1892,N_14186,N_13156);
nor UO_1893 (O_1893,N_12264,N_14720);
nand UO_1894 (O_1894,N_14302,N_12631);
xnor UO_1895 (O_1895,N_12819,N_14095);
nor UO_1896 (O_1896,N_13358,N_12667);
and UO_1897 (O_1897,N_14569,N_13880);
xnor UO_1898 (O_1898,N_14478,N_13942);
or UO_1899 (O_1899,N_14844,N_14678);
nand UO_1900 (O_1900,N_12075,N_12319);
and UO_1901 (O_1901,N_13968,N_14314);
or UO_1902 (O_1902,N_12478,N_14318);
and UO_1903 (O_1903,N_14780,N_14678);
and UO_1904 (O_1904,N_14156,N_12404);
nand UO_1905 (O_1905,N_12612,N_13088);
nor UO_1906 (O_1906,N_14754,N_12336);
and UO_1907 (O_1907,N_13908,N_13321);
nor UO_1908 (O_1908,N_14573,N_14427);
xnor UO_1909 (O_1909,N_12563,N_14911);
xnor UO_1910 (O_1910,N_13943,N_14218);
or UO_1911 (O_1911,N_13430,N_14543);
or UO_1912 (O_1912,N_13610,N_13292);
xor UO_1913 (O_1913,N_12540,N_13770);
xnor UO_1914 (O_1914,N_12787,N_12448);
or UO_1915 (O_1915,N_12412,N_14211);
or UO_1916 (O_1916,N_12504,N_14933);
and UO_1917 (O_1917,N_12710,N_14058);
nor UO_1918 (O_1918,N_12013,N_14388);
or UO_1919 (O_1919,N_12439,N_14032);
nand UO_1920 (O_1920,N_14099,N_12171);
nor UO_1921 (O_1921,N_12080,N_13705);
nor UO_1922 (O_1922,N_13791,N_14030);
and UO_1923 (O_1923,N_13506,N_13363);
and UO_1924 (O_1924,N_12443,N_12190);
nand UO_1925 (O_1925,N_12281,N_14794);
xor UO_1926 (O_1926,N_12809,N_13305);
and UO_1927 (O_1927,N_13032,N_13645);
nand UO_1928 (O_1928,N_13564,N_14644);
xor UO_1929 (O_1929,N_13642,N_14936);
and UO_1930 (O_1930,N_14100,N_13944);
and UO_1931 (O_1931,N_12163,N_12414);
or UO_1932 (O_1932,N_12526,N_13970);
or UO_1933 (O_1933,N_14919,N_14543);
xnor UO_1934 (O_1934,N_12486,N_13753);
xnor UO_1935 (O_1935,N_13991,N_14577);
or UO_1936 (O_1936,N_14509,N_14881);
and UO_1937 (O_1937,N_12504,N_14878);
nand UO_1938 (O_1938,N_14179,N_14790);
nand UO_1939 (O_1939,N_12734,N_13064);
nand UO_1940 (O_1940,N_13596,N_14220);
nand UO_1941 (O_1941,N_12164,N_14593);
nor UO_1942 (O_1942,N_13427,N_14835);
xnor UO_1943 (O_1943,N_12567,N_13217);
nand UO_1944 (O_1944,N_12777,N_12322);
nor UO_1945 (O_1945,N_14528,N_13343);
nand UO_1946 (O_1946,N_12806,N_14248);
xnor UO_1947 (O_1947,N_13717,N_13578);
and UO_1948 (O_1948,N_12655,N_12832);
nand UO_1949 (O_1949,N_13431,N_13261);
xor UO_1950 (O_1950,N_14203,N_13019);
nand UO_1951 (O_1951,N_14614,N_14550);
nand UO_1952 (O_1952,N_14912,N_14719);
nor UO_1953 (O_1953,N_13381,N_14479);
nor UO_1954 (O_1954,N_12838,N_13391);
nor UO_1955 (O_1955,N_14507,N_12908);
or UO_1956 (O_1956,N_13392,N_13849);
xnor UO_1957 (O_1957,N_12032,N_12809);
and UO_1958 (O_1958,N_12767,N_13200);
nand UO_1959 (O_1959,N_13127,N_13907);
nor UO_1960 (O_1960,N_12012,N_14751);
nand UO_1961 (O_1961,N_14335,N_14106);
nor UO_1962 (O_1962,N_12688,N_12374);
nor UO_1963 (O_1963,N_12223,N_13688);
and UO_1964 (O_1964,N_13343,N_12224);
nand UO_1965 (O_1965,N_14662,N_14333);
nor UO_1966 (O_1966,N_12354,N_12521);
or UO_1967 (O_1967,N_12815,N_13937);
and UO_1968 (O_1968,N_14987,N_14976);
xor UO_1969 (O_1969,N_14633,N_14495);
nor UO_1970 (O_1970,N_13370,N_13169);
or UO_1971 (O_1971,N_14381,N_14743);
or UO_1972 (O_1972,N_13340,N_13556);
nand UO_1973 (O_1973,N_13328,N_12530);
nand UO_1974 (O_1974,N_13945,N_12932);
xor UO_1975 (O_1975,N_12602,N_12789);
nor UO_1976 (O_1976,N_12252,N_12733);
and UO_1977 (O_1977,N_12842,N_14068);
xnor UO_1978 (O_1978,N_14513,N_12306);
nand UO_1979 (O_1979,N_12280,N_13457);
xor UO_1980 (O_1980,N_12121,N_14238);
nor UO_1981 (O_1981,N_14467,N_13495);
nor UO_1982 (O_1982,N_14696,N_12997);
nor UO_1983 (O_1983,N_13504,N_13165);
xnor UO_1984 (O_1984,N_13425,N_13349);
xnor UO_1985 (O_1985,N_13450,N_12162);
nand UO_1986 (O_1986,N_14072,N_12577);
or UO_1987 (O_1987,N_13477,N_13619);
nand UO_1988 (O_1988,N_13416,N_13436);
or UO_1989 (O_1989,N_12164,N_13075);
nor UO_1990 (O_1990,N_12737,N_14791);
nand UO_1991 (O_1991,N_13081,N_13034);
and UO_1992 (O_1992,N_14217,N_12260);
xnor UO_1993 (O_1993,N_12254,N_14483);
or UO_1994 (O_1994,N_14940,N_13415);
or UO_1995 (O_1995,N_14213,N_14920);
nand UO_1996 (O_1996,N_12145,N_14333);
or UO_1997 (O_1997,N_12012,N_13542);
xnor UO_1998 (O_1998,N_12636,N_14373);
xnor UO_1999 (O_1999,N_13965,N_13338);
endmodule