module basic_2000_20000_2500_100_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1966,In_1725);
or U1 (N_1,In_866,In_1870);
nand U2 (N_2,In_552,In_833);
nand U3 (N_3,In_1104,In_1317);
nand U4 (N_4,In_1599,In_1435);
xor U5 (N_5,In_199,In_363);
and U6 (N_6,In_1334,In_1103);
nand U7 (N_7,In_1237,In_1469);
xnor U8 (N_8,In_220,In_1574);
or U9 (N_9,In_138,In_37);
and U10 (N_10,In_1576,In_913);
nand U11 (N_11,In_99,In_120);
and U12 (N_12,In_788,In_544);
nor U13 (N_13,In_1090,In_427);
nor U14 (N_14,In_1701,In_864);
xnor U15 (N_15,In_971,In_1368);
nor U16 (N_16,In_300,In_1667);
xor U17 (N_17,In_791,In_1457);
xnor U18 (N_18,In_1621,In_93);
and U19 (N_19,In_1038,In_1482);
nor U20 (N_20,In_648,In_1152);
or U21 (N_21,In_70,In_283);
nand U22 (N_22,In_360,In_1306);
xor U23 (N_23,In_1211,In_1816);
and U24 (N_24,In_1142,In_295);
or U25 (N_25,In_690,In_1984);
nand U26 (N_26,In_21,In_921);
xor U27 (N_27,In_485,In_261);
nor U28 (N_28,In_539,In_69);
xnor U29 (N_29,In_201,In_171);
and U30 (N_30,In_270,In_978);
and U31 (N_31,In_103,In_774);
nand U32 (N_32,In_1866,In_1473);
xor U33 (N_33,In_1380,In_742);
nor U34 (N_34,In_907,In_1463);
or U35 (N_35,In_1112,In_1891);
or U36 (N_36,In_719,In_1625);
xnor U37 (N_37,In_400,In_1627);
nor U38 (N_38,In_383,In_1034);
or U39 (N_39,In_706,In_1254);
or U40 (N_40,In_845,In_1941);
and U41 (N_41,In_1834,In_1326);
xor U42 (N_42,In_1937,In_711);
and U43 (N_43,In_1699,In_899);
and U44 (N_44,In_1978,In_1758);
nor U45 (N_45,In_320,In_1572);
xor U46 (N_46,In_1029,In_1195);
and U47 (N_47,In_1845,In_871);
nor U48 (N_48,In_477,In_747);
xor U49 (N_49,In_1987,In_175);
nand U50 (N_50,In_1147,In_1786);
nor U51 (N_51,In_661,In_1311);
or U52 (N_52,In_1521,In_1780);
nand U53 (N_53,In_150,In_1120);
nand U54 (N_54,In_1278,In_1140);
xor U55 (N_55,In_1575,In_1461);
or U56 (N_56,In_869,In_243);
and U57 (N_57,In_386,In_650);
xor U58 (N_58,In_1442,In_373);
or U59 (N_59,In_556,In_792);
nand U60 (N_60,In_281,In_30);
nand U61 (N_61,In_1033,In_269);
nor U62 (N_62,In_514,In_1502);
nor U63 (N_63,In_1082,In_1549);
and U64 (N_64,In_821,In_1851);
and U65 (N_65,In_96,In_749);
or U66 (N_66,In_966,In_1656);
nor U67 (N_67,In_436,In_1020);
nand U68 (N_68,In_351,In_1266);
nand U69 (N_69,In_693,In_1300);
or U70 (N_70,In_805,In_1507);
or U71 (N_71,In_1044,In_211);
nand U72 (N_72,In_632,In_1624);
nand U73 (N_73,In_1001,In_1737);
nand U74 (N_74,In_624,In_439);
xnor U75 (N_75,In_1377,In_940);
or U76 (N_76,In_413,In_1060);
or U77 (N_77,In_223,In_1399);
xnor U78 (N_78,In_1935,In_252);
or U79 (N_79,In_1894,In_1923);
xor U80 (N_80,In_678,In_1822);
xor U81 (N_81,In_1241,In_106);
nand U82 (N_82,In_893,In_1880);
or U83 (N_83,In_583,In_854);
or U84 (N_84,In_258,In_276);
xor U85 (N_85,In_1253,In_536);
and U86 (N_86,In_1930,In_1610);
nand U87 (N_87,In_1212,In_963);
or U88 (N_88,In_898,In_610);
nand U89 (N_89,In_1421,In_1528);
nand U90 (N_90,In_916,In_1196);
nand U91 (N_91,In_1852,In_853);
and U92 (N_92,In_415,In_1012);
nor U93 (N_93,In_849,In_1312);
xnor U94 (N_94,In_1418,In_1782);
nor U95 (N_95,In_1213,In_1145);
xnor U96 (N_96,In_1976,In_558);
or U97 (N_97,In_1696,In_1531);
xor U98 (N_98,In_1445,In_852);
or U99 (N_99,In_372,In_1516);
or U100 (N_100,In_542,In_524);
xnor U101 (N_101,In_1285,In_1495);
xor U102 (N_102,In_1597,In_744);
and U103 (N_103,In_973,In_680);
nor U104 (N_104,In_1890,In_538);
and U105 (N_105,In_256,In_1491);
or U106 (N_106,In_1168,In_1231);
and U107 (N_107,In_1357,In_926);
and U108 (N_108,In_1708,In_860);
or U109 (N_109,In_1857,In_808);
nand U110 (N_110,In_550,In_599);
or U111 (N_111,In_130,In_265);
nor U112 (N_112,In_229,In_1484);
or U113 (N_113,In_1573,In_1932);
nand U114 (N_114,In_954,In_910);
xor U115 (N_115,In_1524,In_914);
and U116 (N_116,In_1390,In_1587);
nand U117 (N_117,In_1129,In_1692);
or U118 (N_118,In_81,In_667);
nand U119 (N_119,In_98,In_398);
or U120 (N_120,In_1776,In_365);
nand U121 (N_121,In_346,In_294);
nand U122 (N_122,In_100,In_381);
xor U123 (N_123,In_1194,In_24);
nand U124 (N_124,In_955,In_308);
xnor U125 (N_125,In_1592,In_1065);
xor U126 (N_126,In_990,In_594);
nor U127 (N_127,In_414,In_1441);
nor U128 (N_128,In_993,In_1366);
and U129 (N_129,In_141,In_1661);
xor U130 (N_130,In_1022,In_1316);
xor U131 (N_131,In_1819,In_1301);
xor U132 (N_132,In_1769,In_487);
nand U133 (N_133,In_1164,In_262);
and U134 (N_134,In_1471,In_1028);
or U135 (N_135,In_1601,In_753);
or U136 (N_136,In_154,In_32);
or U137 (N_137,In_430,In_1740);
or U138 (N_138,In_1273,In_423);
and U139 (N_139,In_911,In_1024);
or U140 (N_140,In_615,In_1844);
nand U141 (N_141,In_1478,In_33);
and U142 (N_142,In_406,In_301);
xor U143 (N_143,In_694,In_904);
or U144 (N_144,In_649,In_1620);
xor U145 (N_145,In_39,In_483);
nand U146 (N_146,In_104,In_405);
and U147 (N_147,In_1988,In_1553);
or U148 (N_148,In_1055,In_209);
nor U149 (N_149,In_1340,In_1450);
or U150 (N_150,In_1243,In_9);
or U151 (N_151,In_111,In_1973);
and U152 (N_152,In_416,In_1546);
nor U153 (N_153,In_1008,In_1807);
nand U154 (N_154,In_292,In_85);
nor U155 (N_155,In_1041,In_128);
or U156 (N_156,In_870,In_1475);
xor U157 (N_157,In_1210,In_472);
nand U158 (N_158,In_1270,In_1209);
nor U159 (N_159,In_1739,In_516);
nor U160 (N_160,In_927,In_684);
nand U161 (N_161,In_27,In_537);
or U162 (N_162,In_1623,In_961);
nor U163 (N_163,In_432,In_1432);
or U164 (N_164,In_461,In_1729);
or U165 (N_165,In_1189,In_486);
nand U166 (N_166,In_1626,In_738);
nor U167 (N_167,In_331,In_1548);
nor U168 (N_168,In_887,In_1359);
nand U169 (N_169,In_554,In_1386);
nand U170 (N_170,In_314,In_1026);
nor U171 (N_171,In_1867,In_1505);
or U172 (N_172,In_829,In_529);
xnor U173 (N_173,In_463,In_1183);
nand U174 (N_174,In_801,In_1288);
nor U175 (N_175,In_1422,In_254);
or U176 (N_176,In_1251,In_653);
nand U177 (N_177,In_1600,In_1617);
nand U178 (N_178,In_751,In_562);
xnor U179 (N_179,In_1287,In_417);
and U180 (N_180,In_1,In_1375);
or U181 (N_181,In_614,In_376);
nor U182 (N_182,In_1829,In_287);
nand U183 (N_183,In_356,In_1000);
and U184 (N_184,In_124,In_238);
nand U185 (N_185,In_1931,In_1203);
nand U186 (N_186,In_312,In_1897);
or U187 (N_187,In_1410,In_991);
and U188 (N_188,In_953,In_1293);
and U189 (N_189,In_1951,In_210);
or U190 (N_190,In_974,In_1622);
nand U191 (N_191,In_1335,In_1618);
xnor U192 (N_192,In_834,In_1296);
and U193 (N_193,In_717,In_1016);
and U194 (N_194,In_620,In_1248);
xor U195 (N_195,In_1582,In_1438);
and U196 (N_196,In_958,In_205);
or U197 (N_197,In_1174,In_1607);
and U198 (N_198,In_453,In_603);
or U199 (N_199,In_1957,In_972);
and U200 (N_200,In_1281,In_601);
or U201 (N_201,In_402,In_988);
nand U202 (N_202,In_306,In_718);
nand U203 (N_203,N_95,In_1043);
or U204 (N_204,N_142,In_714);
nor U205 (N_205,In_1814,In_1226);
or U206 (N_206,In_585,In_569);
and U207 (N_207,In_1700,In_1710);
nand U208 (N_208,In_876,In_1723);
and U209 (N_209,In_880,N_157);
and U210 (N_210,N_48,In_1709);
xnor U211 (N_211,In_172,In_669);
nor U212 (N_212,In_928,In_1734);
nor U213 (N_213,In_663,In_811);
nor U214 (N_214,In_1961,In_628);
nand U215 (N_215,In_1666,In_859);
xnor U216 (N_216,In_1675,In_1629);
nand U217 (N_217,In_1796,In_345);
and U218 (N_218,In_1439,In_1773);
nand U219 (N_219,In_944,N_19);
nand U220 (N_220,In_1123,In_1052);
nor U221 (N_221,In_702,In_490);
nand U222 (N_222,In_1489,In_772);
and U223 (N_223,In_1855,In_1721);
nand U224 (N_224,N_88,N_154);
xor U225 (N_225,In_1417,In_1101);
nand U226 (N_226,In_802,In_901);
or U227 (N_227,In_1458,In_1821);
and U228 (N_228,In_987,In_1113);
nand U229 (N_229,In_148,In_1651);
and U230 (N_230,In_1173,In_1839);
nand U231 (N_231,N_46,N_57);
nand U232 (N_232,In_942,In_875);
xnor U233 (N_233,In_284,In_445);
or U234 (N_234,In_1798,In_994);
or U235 (N_235,In_1076,In_403);
nand U236 (N_236,In_844,N_105);
and U237 (N_237,In_1545,In_1504);
or U238 (N_238,In_16,In_1088);
xnor U239 (N_239,In_546,In_1283);
or U240 (N_240,In_1771,In_184);
xor U241 (N_241,In_1967,In_563);
and U242 (N_242,In_310,In_855);
nor U243 (N_243,In_1793,In_531);
nor U244 (N_244,In_895,In_1964);
nor U245 (N_245,In_291,In_1010);
and U246 (N_246,In_1274,In_934);
nor U247 (N_247,In_605,In_827);
or U248 (N_248,In_674,In_824);
nand U249 (N_249,In_61,In_822);
xnor U250 (N_250,In_1434,In_631);
xor U251 (N_251,In_1394,In_1983);
and U252 (N_252,In_231,In_88);
or U253 (N_253,In_1615,In_1370);
nor U254 (N_254,In_906,In_1221);
or U255 (N_255,In_1825,In_1079);
xnor U256 (N_256,In_1778,In_236);
or U257 (N_257,In_754,In_1051);
xnor U258 (N_258,In_324,In_1722);
and U259 (N_259,In_1290,In_691);
nor U260 (N_260,In_228,In_1191);
xor U261 (N_261,In_1499,In_1464);
and U262 (N_262,In_634,In_1363);
nor U263 (N_263,In_503,N_140);
nor U264 (N_264,In_968,In_1327);
or U265 (N_265,In_1094,In_1824);
or U266 (N_266,In_159,In_638);
or U267 (N_267,In_1108,In_1423);
and U268 (N_268,In_1862,In_851);
and U269 (N_269,In_133,In_97);
xnor U270 (N_270,In_1025,N_81);
xnor U271 (N_271,In_1401,In_187);
nand U272 (N_272,In_1960,In_336);
nor U273 (N_273,In_580,In_160);
or U274 (N_274,In_1789,In_1384);
nand U275 (N_275,In_481,In_1009);
nand U276 (N_276,In_1838,In_743);
or U277 (N_277,In_1100,In_2);
nor U278 (N_278,In_1813,In_1811);
nand U279 (N_279,In_1519,In_1906);
nand U280 (N_280,In_1718,In_1234);
nor U281 (N_281,In_495,In_447);
and U282 (N_282,N_135,In_377);
or U283 (N_283,In_1985,In_429);
or U284 (N_284,In_1752,In_521);
xnor U285 (N_285,In_1356,In_786);
and U286 (N_286,In_1990,N_179);
or U287 (N_287,In_1480,In_46);
and U288 (N_288,In_1318,In_1325);
or U289 (N_289,In_1331,N_8);
or U290 (N_290,In_272,In_1856);
xor U291 (N_291,In_1229,In_492);
and U292 (N_292,In_361,N_11);
nand U293 (N_293,In_533,In_196);
and U294 (N_294,In_1202,In_448);
xor U295 (N_295,In_1083,N_141);
and U296 (N_296,In_731,In_1550);
xor U297 (N_297,In_1465,In_1002);
or U298 (N_298,In_1118,N_43);
and U299 (N_299,In_724,In_1508);
and U300 (N_300,In_1217,In_703);
xor U301 (N_301,N_54,In_1827);
nand U302 (N_302,In_652,In_568);
or U303 (N_303,In_68,In_671);
and U304 (N_304,In_1797,In_1056);
nand U305 (N_305,In_1228,In_1005);
nor U306 (N_306,In_1351,In_1259);
or U307 (N_307,In_1244,In_1077);
nor U308 (N_308,In_1854,N_174);
nor U309 (N_309,In_996,In_1665);
or U310 (N_310,In_843,In_756);
nor U311 (N_311,In_1955,In_1003);
nor U312 (N_312,In_1383,In_298);
or U313 (N_313,N_158,In_1250);
xor U314 (N_314,In_1818,In_1842);
nor U315 (N_315,In_912,In_362);
xnor U316 (N_316,In_115,In_188);
nor U317 (N_317,In_1058,In_685);
and U318 (N_318,In_1095,In_248);
nand U319 (N_319,In_1433,In_1648);
and U320 (N_320,In_948,In_657);
and U321 (N_321,In_549,In_1276);
and U322 (N_322,In_1977,In_1912);
xor U323 (N_323,N_132,In_83);
nand U324 (N_324,In_1321,In_139);
xnor U325 (N_325,In_1883,In_94);
nand U326 (N_326,In_31,In_584);
nor U327 (N_327,In_86,In_290);
and U328 (N_328,In_1411,In_280);
or U329 (N_329,In_1069,In_178);
xor U330 (N_330,In_1732,In_804);
and U331 (N_331,In_80,In_1346);
or U332 (N_332,In_50,In_1135);
nand U333 (N_333,In_1946,In_1888);
nand U334 (N_334,In_264,In_1460);
xor U335 (N_335,In_479,In_1201);
nand U336 (N_336,In_263,In_517);
xnor U337 (N_337,In_437,In_1858);
nor U338 (N_338,In_697,In_1373);
xnor U339 (N_339,In_750,In_905);
nor U340 (N_340,In_1949,In_1560);
or U341 (N_341,In_1927,In_1064);
xor U342 (N_342,In_710,In_672);
nand U343 (N_343,In_1218,In_1899);
nand U344 (N_344,In_1179,In_1098);
and U345 (N_345,In_1419,In_1903);
nand U346 (N_346,In_1676,In_709);
xor U347 (N_347,In_840,In_1995);
nand U348 (N_348,In_739,In_1641);
nor U349 (N_349,In_1670,In_1671);
nor U350 (N_350,N_126,In_1116);
nand U351 (N_351,In_181,In_488);
or U352 (N_352,In_1282,In_1470);
and U353 (N_353,In_129,In_191);
or U354 (N_354,In_1928,N_188);
xor U355 (N_355,N_133,In_1605);
and U356 (N_356,In_1902,In_440);
nand U357 (N_357,In_1262,In_75);
xor U358 (N_358,In_555,In_806);
and U359 (N_359,In_1875,In_572);
nor U360 (N_360,In_1496,In_450);
and U361 (N_361,In_1569,In_1379);
nor U362 (N_362,In_1182,In_877);
and U363 (N_363,In_1230,In_900);
xnor U364 (N_364,In_1148,N_22);
and U365 (N_365,N_90,In_858);
nand U366 (N_366,In_1677,In_621);
nor U367 (N_367,In_1593,N_162);
xnor U368 (N_368,In_12,In_1893);
and U369 (N_369,In_333,In_1887);
xnor U370 (N_370,In_1063,In_1766);
nor U371 (N_371,In_1777,In_1613);
and U372 (N_372,N_67,In_1804);
and U373 (N_373,In_1877,N_104);
nor U374 (N_374,In_1440,In_1690);
and U375 (N_375,In_570,In_1071);
nor U376 (N_376,In_1768,In_1454);
nor U377 (N_377,In_136,In_1606);
xnor U378 (N_378,In_666,N_134);
nor U379 (N_379,N_59,In_1014);
or U380 (N_380,In_66,In_8);
or U381 (N_381,In_1298,In_989);
and U382 (N_382,In_165,In_609);
or U383 (N_383,In_1013,In_1981);
nor U384 (N_384,In_198,In_177);
nor U385 (N_385,In_1091,N_64);
nand U386 (N_386,In_1110,N_176);
and U387 (N_387,In_1812,In_1246);
and U388 (N_388,In_950,In_579);
xor U389 (N_389,In_1204,In_1257);
and U390 (N_390,In_1896,In_757);
nand U391 (N_391,In_1188,In_787);
or U392 (N_392,N_136,N_198);
nand U393 (N_393,In_997,In_1735);
xor U394 (N_394,In_1004,In_557);
and U395 (N_395,In_1640,N_115);
xnor U396 (N_396,In_1925,In_1653);
nand U397 (N_397,In_186,In_337);
or U398 (N_398,In_459,In_0);
nand U399 (N_399,In_1898,N_73);
xnor U400 (N_400,In_452,In_515);
nand U401 (N_401,In_322,In_1303);
nor U402 (N_402,In_923,In_1205);
nor U403 (N_403,In_780,In_1663);
xor U404 (N_404,In_1403,In_1018);
xor U405 (N_405,In_1871,N_268);
nand U406 (N_406,N_85,In_1706);
xor U407 (N_407,In_836,In_915);
or U408 (N_408,In_867,In_161);
or U409 (N_409,In_1498,In_1494);
nor U410 (N_410,In_1815,N_98);
and U411 (N_411,In_1790,In_1345);
nand U412 (N_412,In_1688,N_302);
nand U413 (N_413,N_25,N_17);
xor U414 (N_414,In_1637,In_341);
and U415 (N_415,In_146,In_156);
xnor U416 (N_416,N_120,N_55);
nand U417 (N_417,In_1920,In_1772);
or U418 (N_418,In_730,In_354);
or U419 (N_419,In_713,In_1309);
nand U420 (N_420,N_262,In_1952);
and U421 (N_421,In_1352,In_34);
nor U422 (N_422,In_783,N_108);
or U423 (N_423,In_1275,In_342);
or U424 (N_424,N_369,In_1668);
nor U425 (N_425,In_1233,In_73);
and U426 (N_426,In_1167,N_168);
xor U427 (N_427,In_909,N_127);
or U428 (N_428,N_214,In_712);
or U429 (N_429,In_1319,In_396);
xnor U430 (N_430,In_687,In_309);
nor U431 (N_431,In_1783,In_1939);
and U432 (N_432,In_1727,In_1794);
or U433 (N_433,In_850,In_1568);
xnor U434 (N_434,N_165,In_1596);
or U435 (N_435,In_140,In_1608);
and U436 (N_436,In_409,In_886);
nand U437 (N_437,N_371,In_1707);
xnor U438 (N_438,In_1297,In_1348);
and U439 (N_439,N_202,In_1933);
or U440 (N_440,N_241,In_534);
or U441 (N_441,N_384,N_167);
and U442 (N_442,In_560,In_1087);
or U443 (N_443,In_387,In_484);
xor U444 (N_444,In_1436,In_986);
or U445 (N_445,In_113,In_832);
xor U446 (N_446,N_124,N_367);
and U447 (N_447,In_602,N_166);
and U448 (N_448,In_1878,N_354);
and U449 (N_449,In_547,In_575);
xnor U450 (N_450,In_704,N_192);
xor U451 (N_451,N_381,In_1415);
nor U452 (N_452,In_1481,In_779);
and U453 (N_453,In_1437,N_109);
or U454 (N_454,In_1350,In_105);
or U455 (N_455,In_1712,N_212);
or U456 (N_456,In_506,In_1302);
nand U457 (N_457,N_189,In_957);
nand U458 (N_458,In_359,In_812);
xor U459 (N_459,In_271,In_1806);
and U460 (N_460,In_1991,In_208);
nor U461 (N_461,In_1389,In_1649);
xor U462 (N_462,In_1965,In_449);
xnor U463 (N_463,In_1595,N_1);
xor U464 (N_464,In_1537,In_1956);
xor U465 (N_465,In_1907,In_607);
nand U466 (N_466,N_234,In_1570);
nand U467 (N_467,In_1242,In_540);
xor U468 (N_468,N_304,In_1042);
and U469 (N_469,In_740,In_795);
xnor U470 (N_470,N_32,In_155);
xnor U471 (N_471,In_1754,N_99);
and U472 (N_472,In_378,In_519);
xnor U473 (N_473,In_1542,In_608);
nand U474 (N_474,In_316,In_1738);
nor U475 (N_475,In_635,In_7);
nand U476 (N_476,In_1632,In_1998);
nand U477 (N_477,In_675,N_143);
or U478 (N_478,N_232,In_1208);
or U479 (N_479,In_1840,In_173);
xnor U480 (N_480,In_1068,In_1443);
nor U481 (N_481,In_1307,In_71);
xor U482 (N_482,In_1176,In_212);
or U483 (N_483,In_1770,In_1015);
nand U484 (N_484,In_716,In_1510);
or U485 (N_485,In_720,In_526);
or U486 (N_486,In_274,In_1150);
xnor U487 (N_487,In_293,In_330);
nand U488 (N_488,In_1566,In_1580);
nor U489 (N_489,N_298,In_576);
nor U490 (N_490,In_606,In_797);
or U491 (N_491,In_659,In_1832);
nor U492 (N_492,In_1074,In_101);
nor U493 (N_493,In_1385,N_252);
or U494 (N_494,In_482,In_1315);
or U495 (N_495,In_1039,In_881);
or U496 (N_496,In_1886,In_1555);
nor U497 (N_497,In_183,In_1067);
and U498 (N_498,In_699,In_1338);
nor U499 (N_499,N_396,In_84);
and U500 (N_500,N_121,In_637);
nand U501 (N_501,In_224,N_201);
xnor U502 (N_502,In_1017,In_397);
and U503 (N_503,In_1579,In_646);
xnor U504 (N_504,In_655,In_673);
nor U505 (N_505,In_1561,N_368);
nor U506 (N_506,In_1809,N_261);
nor U507 (N_507,N_30,In_1944);
or U508 (N_508,N_77,In_582);
nand U509 (N_509,In_393,In_1467);
and U510 (N_510,N_208,N_333);
and U511 (N_511,In_1872,In_1901);
nor U512 (N_512,In_158,In_1396);
nor U513 (N_513,In_323,In_1922);
nand U514 (N_514,In_489,N_26);
nor U515 (N_515,In_1070,In_119);
xnor U516 (N_516,In_941,N_373);
xnor U517 (N_517,In_350,N_346);
or U518 (N_518,In_424,In_434);
nand U519 (N_519,In_1784,N_350);
nand U520 (N_520,In_1636,In_1689);
or U521 (N_521,In_1490,In_1781);
nor U522 (N_522,In_1333,In_525);
or U523 (N_523,In_1134,N_160);
nor U524 (N_524,In_945,N_151);
or U525 (N_525,In_1085,In_1847);
and U526 (N_526,In_1996,In_729);
nand U527 (N_527,N_315,In_1962);
or U528 (N_528,N_97,In_1163);
nand U529 (N_529,N_360,In_932);
nor U530 (N_530,N_207,In_174);
nand U531 (N_531,In_222,In_1765);
and U532 (N_532,In_892,In_763);
or U533 (N_533,In_930,In_1693);
and U534 (N_534,In_1744,In_1048);
or U535 (N_535,In_616,In_10);
xnor U536 (N_536,In_1511,In_1564);
and U537 (N_537,N_288,In_1959);
nor U538 (N_538,N_122,In_935);
or U539 (N_539,In_78,In_1534);
nand U540 (N_540,N_10,In_1388);
nor U541 (N_541,In_1518,In_6);
xor U542 (N_542,In_1371,N_336);
or U543 (N_543,N_362,In_1633);
nor U544 (N_544,In_1376,In_838);
nor U545 (N_545,In_1895,In_268);
nand U546 (N_546,N_335,In_1277);
nor U547 (N_547,In_1645,N_101);
nor U548 (N_548,In_769,In_203);
or U549 (N_549,In_1169,N_163);
and U550 (N_550,In_1820,In_1731);
nor U551 (N_551,In_793,In_286);
xnor U552 (N_552,In_1787,In_225);
nor U553 (N_553,In_1817,In_167);
xnor U554 (N_554,In_166,In_370);
nand U555 (N_555,In_1199,In_1868);
xor U556 (N_556,In_1364,In_58);
nor U557 (N_557,In_462,In_1691);
nand U558 (N_558,N_280,N_310);
nand U559 (N_559,In_11,In_1247);
and U560 (N_560,In_765,In_596);
nor U561 (N_561,In_1520,N_397);
and U562 (N_562,In_1683,In_682);
nor U563 (N_563,In_1089,In_467);
nor U564 (N_564,In_1571,In_1743);
nor U565 (N_565,N_236,N_195);
and U566 (N_566,In_433,In_412);
nand U567 (N_567,In_1971,N_295);
nor U568 (N_568,In_282,In_1180);
xor U569 (N_569,In_1007,In_1105);
xor U570 (N_570,In_4,In_1159);
nand U571 (N_571,N_322,In_250);
xnor U572 (N_572,N_228,In_407);
and U573 (N_573,In_1075,N_70);
or U574 (N_574,In_642,In_748);
nand U575 (N_575,In_782,In_815);
xor U576 (N_576,In_504,N_215);
nand U577 (N_577,In_1979,In_1753);
xnor U578 (N_578,N_203,In_1023);
or U579 (N_579,In_1759,In_1304);
and U580 (N_580,In_1889,In_499);
or U581 (N_581,In_1835,In_214);
or U582 (N_582,In_1848,In_530);
nor U583 (N_583,N_71,In_1448);
nand U584 (N_584,N_110,In_679);
nand U585 (N_585,N_177,N_4);
nor U586 (N_586,In_458,In_1031);
and U587 (N_587,N_199,In_796);
nand U588 (N_588,In_1466,N_156);
xor U589 (N_589,In_1642,In_1919);
xor U590 (N_590,In_1562,In_180);
and U591 (N_591,In_874,N_211);
or U592 (N_592,In_1513,N_393);
and U593 (N_593,In_1329,In_1057);
or U594 (N_594,In_1404,In_1139);
and U595 (N_595,In_574,In_369);
or U596 (N_596,N_386,N_14);
xor U597 (N_597,N_123,In_1800);
or U598 (N_598,In_1157,In_1178);
or U599 (N_599,N_170,In_185);
and U600 (N_600,In_1405,N_531);
nand U601 (N_601,In_230,In_117);
nand U602 (N_602,In_761,In_908);
nor U603 (N_603,In_108,N_497);
nor U604 (N_604,In_1940,N_356);
xor U605 (N_605,In_677,In_1638);
nand U606 (N_606,N_282,N_487);
and U607 (N_607,In_1267,In_375);
and U608 (N_608,In_48,N_130);
and U609 (N_609,In_194,N_153);
xnor U610 (N_610,N_496,N_300);
nor U611 (N_611,In_980,N_405);
nand U612 (N_612,N_559,N_594);
nor U613 (N_613,N_486,In_1970);
nand U614 (N_614,In_857,N_424);
nand U615 (N_615,N_444,N_427);
nor U616 (N_616,N_33,In_1803);
xnor U617 (N_617,In_1092,In_95);
nor U618 (N_618,In_597,In_1551);
xor U619 (N_619,N_137,N_338);
and U620 (N_620,In_809,In_60);
xnor U621 (N_621,N_183,In_460);
and U622 (N_622,In_1252,In_1831);
nor U623 (N_623,In_1914,N_556);
nand U624 (N_624,In_960,In_762);
or U625 (N_625,In_1413,In_1369);
nand U626 (N_626,In_1130,In_17);
nor U627 (N_627,In_888,N_325);
or U628 (N_628,In_1861,N_148);
or U629 (N_629,In_131,N_45);
nand U630 (N_630,In_532,In_1751);
or U631 (N_631,N_511,N_265);
and U632 (N_632,In_1330,In_1046);
nor U633 (N_633,In_1745,N_512);
and U634 (N_634,In_1628,In_1910);
xor U635 (N_635,In_419,N_578);
nor U636 (N_636,In_1631,In_217);
nor U637 (N_637,In_1830,In_1323);
or U638 (N_638,N_320,In_1885);
nor U639 (N_639,In_1374,In_1506);
nor U640 (N_640,N_538,In_588);
xor U641 (N_641,In_259,N_31);
nand U642 (N_642,N_469,In_62);
nand U643 (N_643,In_1165,In_818);
nand U644 (N_644,In_1805,In_338);
xnor U645 (N_645,In_493,In_480);
nor U646 (N_646,In_1911,N_190);
nor U647 (N_647,N_509,In_1050);
nor U648 (N_648,In_586,In_428);
nor U649 (N_649,In_1543,In_658);
and U650 (N_650,N_545,In_670);
nor U651 (N_651,In_938,In_1828);
nor U652 (N_652,N_599,N_216);
xnor U653 (N_653,In_1236,In_143);
nor U654 (N_654,In_1604,In_1310);
nand U655 (N_655,N_383,In_630);
nand U656 (N_656,N_391,In_457);
xor U657 (N_657,In_152,In_771);
nand U658 (N_658,In_466,In_577);
nor U659 (N_659,N_425,In_523);
xnor U660 (N_660,In_878,N_205);
nor U661 (N_661,In_1873,In_1774);
and U662 (N_662,In_112,In_444);
and U663 (N_663,In_169,In_1062);
xor U664 (N_664,N_449,In_326);
nor U665 (N_665,In_826,N_518);
or U666 (N_666,In_766,In_1724);
nor U667 (N_667,In_1767,N_351);
xor U668 (N_668,In_343,N_184);
and U669 (N_669,In_810,In_1036);
xor U670 (N_670,N_308,In_1255);
and U671 (N_671,N_510,N_474);
nand U672 (N_672,In_1539,In_1673);
xor U673 (N_673,In_469,N_331);
nor U674 (N_674,In_1156,In_701);
xor U675 (N_675,In_949,In_510);
nand U676 (N_676,N_13,N_592);
or U677 (N_677,In_1954,N_76);
xor U678 (N_678,In_303,N_225);
or U679 (N_679,In_1530,N_358);
or U680 (N_680,N_388,N_585);
xnor U681 (N_681,N_169,N_451);
nand U682 (N_682,In_511,N_507);
nand U683 (N_683,N_401,N_477);
or U684 (N_684,In_153,In_1681);
xnor U685 (N_685,In_626,In_999);
xnor U686 (N_686,N_567,In_1171);
nor U687 (N_687,In_1552,N_279);
nor U688 (N_688,In_57,N_442);
nor U689 (N_689,N_36,In_1472);
and U690 (N_690,In_1261,In_681);
or U691 (N_691,In_1072,N_570);
nor U692 (N_692,In_856,In_25);
nand U693 (N_693,In_456,In_1121);
and U694 (N_694,In_425,In_1249);
xnor U695 (N_695,In_1515,In_1341);
and U696 (N_696,In_1144,In_1177);
and U697 (N_697,N_223,N_492);
nor U698 (N_698,In_918,In_1133);
xnor U699 (N_699,N_299,In_380);
and U700 (N_700,N_506,In_3);
nand U701 (N_701,N_283,In_1214);
nand U702 (N_702,In_700,In_226);
xnor U703 (N_703,N_348,N_292);
and U704 (N_704,In_1646,In_1468);
xor U705 (N_705,In_1387,In_1741);
nand U706 (N_706,N_404,In_1791);
or U707 (N_707,N_555,In_1557);
and U708 (N_708,N_119,N_479);
and U709 (N_709,In_227,In_1313);
nor U710 (N_710,N_565,In_689);
xnor U711 (N_711,In_426,In_528);
nand U712 (N_712,In_1032,In_1760);
or U713 (N_713,In_758,In_401);
xnor U714 (N_714,In_1583,In_883);
or U715 (N_715,In_936,In_831);
xor U716 (N_716,N_439,In_72);
or U717 (N_717,In_625,In_1446);
and U718 (N_718,In_195,N_422);
nand U719 (N_719,In_773,In_497);
or U720 (N_720,N_125,In_149);
or U721 (N_721,In_1652,In_277);
or U722 (N_722,In_1337,In_395);
or U723 (N_723,N_220,In_1657);
xnor U724 (N_724,In_520,In_91);
or U725 (N_725,N_560,N_38);
xnor U726 (N_726,In_1219,N_540);
nand U727 (N_727,In_132,N_317);
xor U728 (N_728,In_889,N_436);
xor U729 (N_729,N_29,In_545);
nand U730 (N_730,In_1992,In_145);
xor U731 (N_731,In_399,In_1968);
and U732 (N_732,In_1053,In_647);
xor U733 (N_733,In_564,In_1837);
nor U734 (N_734,N_558,N_253);
nor U735 (N_735,N_218,In_221);
nand U736 (N_736,In_1453,In_278);
nand U737 (N_737,In_1455,In_862);
nand U738 (N_738,In_865,N_593);
xnor U739 (N_739,In_1097,In_501);
or U740 (N_740,In_922,N_353);
and U741 (N_741,N_480,N_159);
or U742 (N_742,In_1155,N_464);
and U743 (N_743,In_26,N_467);
or U744 (N_744,N_118,In_364);
nand U745 (N_745,In_593,In_1578);
xnor U746 (N_746,In_1541,In_1324);
xnor U747 (N_747,In_1349,N_562);
nand U748 (N_748,N_535,N_264);
xor U749 (N_749,In_1908,In_1634);
nor U750 (N_750,N_175,In_1892);
xor U751 (N_751,In_507,N_347);
nand U752 (N_752,In_1603,In_1594);
and U753 (N_753,N_15,In_1080);
or U754 (N_754,In_1884,N_92);
or U755 (N_755,In_1378,In_1882);
nor U756 (N_756,In_688,In_1096);
nand U757 (N_757,In_273,N_529);
nor U758 (N_758,In_734,In_589);
xnor U759 (N_759,N_266,N_235);
xnor U760 (N_760,N_68,N_344);
or U761 (N_761,In_1332,N_324);
nor U762 (N_762,N_355,In_839);
nor U763 (N_763,In_1591,N_62);
and U764 (N_764,In_1493,In_109);
and U765 (N_765,In_1149,In_527);
nor U766 (N_766,In_636,In_1424);
xor U767 (N_767,In_1459,N_548);
nor U768 (N_768,In_1486,N_82);
nor U769 (N_769,In_1958,In_1755);
xnor U770 (N_770,In_1292,In_814);
or U771 (N_771,In_65,In_266);
nand U772 (N_772,In_931,In_640);
nor U773 (N_773,N_554,In_651);
nor U774 (N_774,In_1850,In_1295);
nor U775 (N_775,In_1073,N_517);
nand U776 (N_776,N_80,In_89);
nand U777 (N_777,In_438,N_489);
or U778 (N_778,In_1132,In_1558);
and U779 (N_779,N_246,In_1567);
nor U780 (N_780,N_9,In_1355);
xor U781 (N_781,In_1258,N_495);
and U782 (N_782,In_1107,N_240);
nand U783 (N_783,N_65,N_277);
and U784 (N_784,In_1540,In_1563);
xor U785 (N_785,N_463,In_1409);
or U786 (N_786,In_1239,In_1299);
nand U787 (N_787,In_777,In_983);
or U788 (N_788,In_1697,In_1619);
nand U789 (N_789,In_1444,In_1864);
or U790 (N_790,N_458,N_420);
or U791 (N_791,In_789,N_521);
nand U792 (N_792,In_1286,In_1452);
and U793 (N_793,N_468,In_470);
nand U794 (N_794,In_1197,N_272);
xnor U795 (N_795,In_368,In_847);
nor U796 (N_796,In_374,In_19);
nand U797 (N_797,In_1533,In_1565);
and U798 (N_798,N_145,In_1853);
nand U799 (N_799,In_981,In_725);
nand U800 (N_800,In_1294,N_206);
nor U801 (N_801,In_1736,In_841);
nand U802 (N_802,N_102,In_47);
nand U803 (N_803,N_723,N_452);
xor U804 (N_804,In_56,N_100);
xor U805 (N_805,N_505,N_374);
nor U806 (N_806,In_245,In_1027);
and U807 (N_807,N_462,In_357);
nor U808 (N_808,N_129,In_1660);
xor U809 (N_809,In_662,N_611);
nor U810 (N_810,N_693,In_1059);
xor U811 (N_811,In_43,In_1172);
nand U812 (N_812,N_634,In_1588);
or U813 (N_813,In_946,N_297);
xnor U814 (N_814,N_116,In_1393);
xor U815 (N_815,N_568,N_605);
nand U816 (N_816,N_44,N_481);
xnor U817 (N_817,In_1265,In_468);
nor U818 (N_818,N_485,N_343);
nand U819 (N_819,In_52,In_872);
or U820 (N_820,In_454,In_1131);
nand U821 (N_821,N_385,N_484);
and U822 (N_822,N_466,In_1381);
nor U823 (N_823,N_654,N_595);
or U824 (N_824,In_1447,In_1905);
nor U825 (N_825,In_28,In_604);
and U826 (N_826,N_434,In_394);
and U827 (N_827,N_460,In_1756);
xor U828 (N_828,N_672,In_1187);
xnor U829 (N_829,N_490,In_1926);
nor U830 (N_830,In_253,N_527);
nand U831 (N_831,In_1529,In_51);
or U832 (N_832,N_651,N_60);
nand U833 (N_833,In_1503,N_644);
and U834 (N_834,In_1146,N_229);
nand U835 (N_835,In_344,N_582);
nor U836 (N_836,In_18,N_653);
nor U837 (N_837,N_683,In_705);
xnor U838 (N_838,N_665,In_976);
and U839 (N_839,In_741,In_1788);
and U840 (N_840,N_89,In_803);
xnor U841 (N_841,N_756,In_125);
and U842 (N_842,N_441,In_49);
nor U843 (N_843,N_12,N_366);
and U844 (N_844,N_243,In_873);
nand U845 (N_845,In_722,In_137);
nor U846 (N_846,N_783,N_616);
xor U847 (N_847,N_244,N_631);
and U848 (N_848,In_726,In_123);
or U849 (N_849,N_433,In_1836);
nor U850 (N_850,In_979,N_667);
or U851 (N_851,In_1614,In_1975);
and U852 (N_852,In_1392,N_412);
nor U853 (N_853,N_785,N_239);
nand U854 (N_854,N_774,In_746);
nor U855 (N_855,In_1590,N_289);
nor U856 (N_856,In_410,In_654);
and U857 (N_857,N_619,In_1102);
nand U858 (N_858,In_1081,N_482);
nand U859 (N_859,N_306,N_37);
nand U860 (N_860,In_289,N_523);
nor U861 (N_861,In_1268,N_2);
nand U862 (N_862,N_522,In_216);
and U863 (N_863,In_1414,In_1801);
xnor U864 (N_864,In_82,In_299);
nor U865 (N_865,In_1602,In_1989);
and U866 (N_866,N_94,N_620);
nor U867 (N_867,In_455,In_1216);
and U868 (N_868,N_617,In_1019);
nor U869 (N_869,N_370,N_668);
and U870 (N_870,N_483,In_1488);
or U871 (N_871,N_430,N_794);
xnor U872 (N_872,N_504,In_1485);
xor U873 (N_873,N_147,In_745);
nand U874 (N_874,N_685,N_589);
and U875 (N_875,In_464,N_472);
and U876 (N_876,In_189,N_498);
nor U877 (N_877,N_768,In_1554);
and U878 (N_878,In_641,N_669);
nand U879 (N_879,N_703,In_695);
xor U880 (N_880,In_1222,In_435);
nand U881 (N_881,N_602,In_45);
xnor U882 (N_882,In_335,N_547);
nand U883 (N_883,In_1154,N_686);
or U884 (N_884,N_7,N_69);
nand U885 (N_885,In_755,In_1943);
nor U886 (N_886,In_1716,In_1280);
and U887 (N_887,In_1138,N_630);
nand U888 (N_888,In_1662,In_1682);
xnor U889 (N_889,N_701,In_885);
xor U890 (N_890,In_1532,N_51);
or U891 (N_891,In_1577,N_673);
nand U892 (N_892,In_267,N_743);
nand U893 (N_893,N_682,N_571);
or U894 (N_894,In_698,In_392);
nor U895 (N_895,N_695,N_622);
xnor U896 (N_896,In_764,N_777);
and U897 (N_897,In_500,N_561);
or U898 (N_898,N_514,N_251);
nand U899 (N_899,In_411,In_421);
or U900 (N_900,In_192,N_689);
xnor U901 (N_901,In_77,N_704);
nor U902 (N_902,In_134,N_74);
xnor U903 (N_903,In_1184,In_759);
and U904 (N_904,In_1517,In_985);
nand U905 (N_905,In_952,In_1702);
or U906 (N_906,In_279,In_1650);
xor U907 (N_907,In_1406,N_491);
and U908 (N_908,N_376,N_66);
or U909 (N_909,In_1589,N_440);
nor U910 (N_910,In_1609,In_1336);
and U911 (N_911,N_569,In_1170);
nand U912 (N_912,In_471,In_349);
or U913 (N_913,N_493,N_674);
xor U914 (N_914,N_731,In_969);
or U915 (N_915,In_307,In_708);
and U916 (N_916,N_410,N_372);
nand U917 (N_917,N_742,In_559);
xor U918 (N_918,In_1207,In_1106);
xnor U919 (N_919,N_471,N_528);
nand U920 (N_920,N_270,In_1291);
and U921 (N_921,In_321,N_645);
nor U922 (N_922,In_443,In_897);
nor U923 (N_923,In_304,N_146);
xor U924 (N_924,N_93,In_204);
or U925 (N_925,N_649,N_294);
or U926 (N_926,N_23,In_1999);
nor U927 (N_927,In_1680,In_382);
nor U928 (N_928,In_1559,In_1361);
xnor U929 (N_929,N_574,In_1762);
nor U930 (N_930,In_241,In_1192);
or U931 (N_931,In_206,N_716);
nand U932 (N_932,In_182,N_769);
xor U933 (N_933,N_197,In_781);
nand U934 (N_934,In_352,In_1644);
xnor U935 (N_935,In_1779,N_637);
nand U936 (N_936,N_72,In_578);
and U937 (N_937,In_1969,In_1726);
and U938 (N_938,In_1994,In_1126);
xor U939 (N_939,In_1185,N_263);
nor U940 (N_940,N_546,In_1353);
nand U941 (N_941,N_473,In_894);
or U942 (N_942,N_332,In_598);
xor U943 (N_943,In_1186,N_470);
xor U944 (N_944,In_721,In_643);
and U945 (N_945,N_274,In_1430);
and U946 (N_946,In_347,In_1358);
nand U947 (N_947,In_122,N_799);
or U948 (N_948,In_1269,In_451);
or U949 (N_949,In_591,In_644);
xor U950 (N_950,N_664,In_1040);
and U951 (N_951,N_96,In_35);
nand U952 (N_952,In_623,N_387);
or U953 (N_953,N_722,In_38);
and U954 (N_954,In_1021,N_112);
nor U955 (N_955,N_789,N_713);
or U956 (N_956,N_760,In_1993);
nor U957 (N_957,N_155,In_157);
nor U958 (N_958,In_1161,In_1030);
and U959 (N_959,In_1099,N_213);
xnor U960 (N_960,N_564,N_50);
nand U961 (N_961,N_150,In_107);
and U962 (N_962,In_1746,N_708);
or U963 (N_963,N_286,N_580);
and U964 (N_964,N_579,N_660);
and U965 (N_965,N_382,In_1117);
and U966 (N_966,N_526,N_128);
or U967 (N_967,In_1826,N_583);
nor U968 (N_968,In_1544,N_200);
nand U969 (N_969,In_1225,In_939);
nor U970 (N_970,N_224,In_29);
nor U971 (N_971,In_1279,N_106);
xnor U972 (N_972,N_342,N_24);
xor U973 (N_973,In_1764,N_305);
nor U974 (N_974,In_509,N_721);
nor U975 (N_975,In_1799,N_407);
nor U976 (N_976,In_1924,In_1654);
and U977 (N_977,N_86,N_639);
and U978 (N_978,N_718,In_1704);
nor U979 (N_979,In_1581,In_15);
nor U980 (N_980,In_1500,In_1412);
nand U981 (N_981,N_341,N_87);
or U982 (N_982,N_550,In_573);
and U983 (N_983,In_1742,N_632);
xor U984 (N_984,In_785,In_297);
xnor U985 (N_985,N_640,In_1795);
and U986 (N_986,In_257,N_603);
nor U987 (N_987,N_27,In_334);
nor U988 (N_988,In_622,N_752);
nor U989 (N_989,In_1686,In_676);
xnor U990 (N_990,N_587,N_49);
or U991 (N_991,In_126,In_502);
or U992 (N_992,N_584,In_1425);
or U993 (N_993,N_719,In_1344);
or U994 (N_994,N_329,In_215);
nand U995 (N_995,In_179,N_519);
xor U996 (N_996,In_1235,In_275);
and U997 (N_997,In_1122,N_696);
xor U998 (N_998,In_1538,In_1775);
nand U999 (N_999,N_380,N_58);
nand U1000 (N_1000,N_678,N_276);
nand U1001 (N_1001,N_609,In_1078);
xnor U1002 (N_1002,In_1748,N_415);
or U1003 (N_1003,N_949,N_544);
nand U1004 (N_1004,In_600,In_442);
xor U1005 (N_1005,N_476,N_865);
xor U1006 (N_1006,N_702,N_895);
nor U1007 (N_1007,N_532,In_1109);
nand U1008 (N_1008,In_943,N_699);
nor U1009 (N_1009,N_557,In_1833);
xor U1010 (N_1010,N_993,N_323);
nand U1011 (N_1011,N_186,N_194);
or U1012 (N_1012,N_961,N_725);
nor U1013 (N_1013,N_807,In_1982);
and U1014 (N_1014,N_377,In_127);
nand U1015 (N_1015,N_754,In_1264);
or U1016 (N_1016,In_1674,In_1308);
xnor U1017 (N_1017,N_745,In_296);
nand U1018 (N_1018,N_798,N_242);
xor U1019 (N_1019,N_963,In_219);
nor U1020 (N_1020,In_247,In_982);
xnor U1021 (N_1021,N_824,In_1125);
xor U1022 (N_1022,In_233,N_671);
xor U1023 (N_1023,In_1492,N_800);
nand U1024 (N_1024,N_296,N_996);
nand U1025 (N_1025,N_307,N_676);
nand U1026 (N_1026,In_1227,N_284);
nor U1027 (N_1027,In_1049,N_915);
or U1028 (N_1028,N_931,N_684);
or U1029 (N_1029,N_608,N_437);
nor U1030 (N_1030,N_808,In_1728);
xnor U1031 (N_1031,N_862,N_278);
and U1032 (N_1032,N_648,In_665);
xor U1033 (N_1033,N_290,N_729);
nor U1034 (N_1034,In_890,In_590);
nand U1035 (N_1035,In_1711,N_138);
xor U1036 (N_1036,In_727,N_400);
nor U1037 (N_1037,In_863,In_776);
nand U1038 (N_1038,N_47,N_221);
or U1039 (N_1039,N_995,In_1382);
xor U1040 (N_1040,In_518,In_1947);
xor U1041 (N_1041,N_748,In_1938);
nor U1042 (N_1042,In_200,N_516);
and U1043 (N_1043,In_1224,N_494);
or U1044 (N_1044,In_329,N_948);
and U1045 (N_1045,N_455,In_929);
nor U1046 (N_1046,In_197,In_1879);
xnor U1047 (N_1047,In_422,In_1158);
or U1048 (N_1048,In_1909,N_853);
nor U1049 (N_1049,N_914,In_1011);
and U1050 (N_1050,N_149,N_870);
xnor U1051 (N_1051,N_917,In_1647);
or U1052 (N_1052,N_6,In_1175);
or U1053 (N_1053,In_956,In_696);
xnor U1054 (N_1054,N_258,N_952);
xnor U1055 (N_1055,In_237,N_293);
xor U1056 (N_1056,In_1869,In_431);
xor U1057 (N_1057,In_418,N_709);
xnor U1058 (N_1058,In_618,N_894);
or U1059 (N_1059,N_784,N_563);
nor U1060 (N_1060,N_423,In_1616);
nand U1061 (N_1061,N_817,In_984);
nand U1062 (N_1062,In_1972,In_1703);
or U1063 (N_1063,N_955,N_921);
xnor U1064 (N_1064,N_726,In_884);
xor U1065 (N_1065,N_937,N_641);
nor U1066 (N_1066,In_1997,N_775);
nor U1067 (N_1067,In_1420,N_834);
nand U1068 (N_1068,N_610,N_524);
nor U1069 (N_1069,In_1929,N_848);
nor U1070 (N_1070,N_982,In_1320);
nand U1071 (N_1071,In_371,N_267);
xor U1072 (N_1072,N_764,N_363);
xor U1073 (N_1073,N_312,N_872);
and U1074 (N_1074,In_244,In_246);
xnor U1075 (N_1075,In_234,In_1525);
nor U1076 (N_1076,In_318,N_394);
or U1077 (N_1077,In_44,N_780);
nand U1078 (N_1078,In_1477,N_275);
xnor U1079 (N_1079,N_746,N_41);
nor U1080 (N_1080,N_222,N_662);
or U1081 (N_1081,N_891,In_1913);
xnor U1082 (N_1082,N_542,N_365);
and U1083 (N_1083,N_475,N_913);
nand U1084 (N_1084,In_116,In_319);
and U1085 (N_1085,N_938,In_1160);
nand U1086 (N_1086,N_705,N_359);
and U1087 (N_1087,N_349,N_328);
and U1088 (N_1088,In_1220,N_78);
xor U1089 (N_1089,N_34,N_431);
or U1090 (N_1090,N_233,N_209);
nor U1091 (N_1091,N_285,In_384);
and U1092 (N_1092,N_943,In_732);
xor U1093 (N_1093,N_659,N_788);
nand U1094 (N_1094,N_835,In_1128);
xor U1095 (N_1095,N_314,In_63);
nand U1096 (N_1096,In_925,N_852);
xor U1097 (N_1097,In_404,N_828);
or U1098 (N_1098,N_334,N_409);
nor U1099 (N_1099,N_782,In_1679);
and U1100 (N_1100,In_1556,In_1006);
nand U1101 (N_1101,N_990,In_1672);
nor U1102 (N_1102,N_846,In_1980);
nand U1103 (N_1103,N_967,N_841);
xor U1104 (N_1104,N_75,In_478);
nand U1105 (N_1105,In_1658,In_1598);
xor U1106 (N_1106,In_828,N_707);
nand U1107 (N_1107,In_541,In_1119);
nand U1108 (N_1108,N_792,N_503);
nand U1109 (N_1109,In_553,N_152);
nand U1110 (N_1110,In_505,In_1843);
nor U1111 (N_1111,In_1476,N_759);
and U1112 (N_1112,In_735,N_465);
xor U1113 (N_1113,In_1398,In_76);
nand U1114 (N_1114,N_956,N_204);
xor U1115 (N_1115,N_903,N_530);
and U1116 (N_1116,N_882,In_819);
xor U1117 (N_1117,N_499,In_1181);
or U1118 (N_1118,N_944,N_478);
xor U1119 (N_1119,In_110,N_898);
and U1120 (N_1120,N_951,In_1407);
or U1121 (N_1121,In_1841,In_992);
or U1122 (N_1122,In_784,N_823);
or U1123 (N_1123,N_210,In_629);
nor U1124 (N_1124,In_1876,N_180);
or U1125 (N_1125,N_364,In_565);
or U1126 (N_1126,N_858,In_1715);
and U1127 (N_1127,N_879,In_1904);
nor U1128 (N_1128,In_420,In_613);
or U1129 (N_1129,In_408,In_581);
xnor U1130 (N_1130,In_775,N_591);
nand U1131 (N_1131,In_1719,N_691);
or U1132 (N_1132,N_453,N_428);
xor U1133 (N_1133,In_1630,N_670);
nor U1134 (N_1134,In_879,N_392);
xnor U1135 (N_1135,In_353,N_411);
nand U1136 (N_1136,N_953,N_604);
and U1137 (N_1137,N_749,In_379);
or U1138 (N_1138,N_985,N_977);
nand U1139 (N_1139,In_656,N_779);
xnor U1140 (N_1140,In_861,In_1066);
xnor U1141 (N_1141,In_1687,In_1035);
xor U1142 (N_1142,N_330,N_925);
nor U1143 (N_1143,N_987,In_1136);
nand U1144 (N_1144,N_839,In_1479);
and U1145 (N_1145,N_681,In_14);
xnor U1146 (N_1146,N_793,In_74);
and U1147 (N_1147,In_1874,In_686);
nor U1148 (N_1148,In_1260,N_859);
nor U1149 (N_1149,In_1497,In_633);
nand U1150 (N_1150,In_778,N_551);
nor U1151 (N_1151,In_23,N_677);
nand U1152 (N_1152,In_1865,N_28);
and U1153 (N_1153,N_395,N_249);
nand U1154 (N_1154,In_903,N_981);
nor U1155 (N_1155,N_337,N_607);
and U1156 (N_1156,In_90,In_446);
nor U1157 (N_1157,In_1190,N_408);
and U1158 (N_1158,N_978,N_533);
nor U1159 (N_1159,In_1400,N_908);
and U1160 (N_1160,In_249,N_904);
nor U1161 (N_1161,N_435,N_379);
xor U1162 (N_1162,N_79,In_1695);
nor U1163 (N_1163,N_248,In_1354);
or U1164 (N_1164,N_869,In_548);
nor U1165 (N_1165,In_1792,In_1193);
nand U1166 (N_1166,In_494,N_131);
or U1167 (N_1167,In_366,N_217);
xnor U1168 (N_1168,N_52,In_1698);
and U1169 (N_1169,N_313,N_918);
nand U1170 (N_1170,N_740,In_475);
nor U1171 (N_1171,N_791,N_445);
xor U1172 (N_1172,In_388,N_231);
nand U1173 (N_1173,N_643,N_697);
nor U1174 (N_1174,N_172,In_64);
and U1175 (N_1175,N_456,N_886);
xnor U1176 (N_1176,N_161,N_973);
or U1177 (N_1177,N_389,In_1428);
xor U1178 (N_1178,In_816,N_650);
nand U1179 (N_1179,N_260,In_118);
nor U1180 (N_1180,N_39,N_316);
or U1181 (N_1181,N_536,N_922);
nand U1182 (N_1182,N_950,In_611);
or U1183 (N_1183,N_761,N_694);
xor U1184 (N_1184,N_847,N_688);
nand U1185 (N_1185,In_251,In_1037);
or U1186 (N_1186,In_902,In_522);
and U1187 (N_1187,N_720,N_113);
nand U1188 (N_1188,In_367,N_912);
nand U1189 (N_1189,In_1921,N_924);
xor U1190 (N_1190,N_849,In_325);
xnor U1191 (N_1191,In_1483,In_813);
or U1192 (N_1192,In_1314,In_1730);
nand U1193 (N_1193,N_906,In_1859);
nand U1194 (N_1194,In_794,In_1124);
xor U1195 (N_1195,N_340,N_960);
nand U1196 (N_1196,N_586,In_882);
nor U1197 (N_1197,N_291,In_595);
nand U1198 (N_1198,N_638,In_891);
or U1199 (N_1199,N_797,N_107);
nor U1200 (N_1200,N_1148,N_1079);
xor U1201 (N_1201,N_770,N_1111);
or U1202 (N_1202,In_207,N_875);
or U1203 (N_1203,N_416,N_1033);
and U1204 (N_1204,In_232,In_1240);
nand U1205 (N_1205,N_1133,N_1147);
or U1206 (N_1206,N_621,In_566);
nor U1207 (N_1207,N_1027,In_1535);
nand U1208 (N_1208,In_1763,N_311);
xor U1209 (N_1209,N_930,N_899);
nand U1210 (N_1210,N_755,N_144);
xor U1211 (N_1211,N_259,In_1115);
nand U1212 (N_1212,In_441,N_345);
xor U1213 (N_1213,N_375,N_0);
nand U1214 (N_1214,In_242,N_878);
or U1215 (N_1215,N_1104,In_1860);
and U1216 (N_1216,N_945,In_951);
nor U1217 (N_1217,In_1151,In_1289);
nand U1218 (N_1218,In_496,N_766);
xnor U1219 (N_1219,N_1061,In_733);
xnor U1220 (N_1220,N_647,In_328);
nor U1221 (N_1221,N_1059,N_450);
nor U1222 (N_1222,In_933,N_821);
nor U1223 (N_1223,N_181,N_836);
nor U1224 (N_1224,N_1194,N_999);
or U1225 (N_1225,N_273,N_833);
or U1226 (N_1226,N_596,N_16);
or U1227 (N_1227,In_1986,N_646);
or U1228 (N_1228,In_1684,In_164);
xor U1229 (N_1229,In_770,In_723);
xor U1230 (N_1230,In_168,N_1016);
or U1231 (N_1231,N_860,N_1019);
nand U1232 (N_1232,In_728,In_1238);
and U1233 (N_1233,N_805,N_1178);
nor U1234 (N_1234,N_1131,In_975);
xor U1235 (N_1235,N_1040,In_1863);
nand U1236 (N_1236,In_1747,N_1105);
and U1237 (N_1237,N_975,N_1021);
or U1238 (N_1238,N_1182,In_498);
nand U1239 (N_1239,In_1523,N_790);
or U1240 (N_1240,N_831,In_358);
nand U1241 (N_1241,N_1167,In_627);
xor U1242 (N_1242,N_227,In_1272);
nand U1243 (N_1243,N_1042,N_700);
and U1244 (N_1244,N_281,N_1114);
and U1245 (N_1245,N_61,N_173);
xor U1246 (N_1246,N_352,N_1097);
or U1247 (N_1247,N_910,N_692);
xnor U1248 (N_1248,In_1757,N_946);
or U1249 (N_1249,N_737,In_1785);
xor U1250 (N_1250,N_812,N_1012);
xnor U1251 (N_1251,N_1190,N_861);
or U1252 (N_1252,N_1064,N_1084);
and U1253 (N_1253,N_1075,In_59);
or U1254 (N_1254,N_525,N_247);
and U1255 (N_1255,In_1137,N_679);
and U1256 (N_1256,N_863,N_398);
and U1257 (N_1257,In_1416,N_675);
or U1258 (N_1258,In_1093,In_1974);
xor U1259 (N_1259,N_818,N_1045);
and U1260 (N_1260,N_21,N_1112);
nor U1261 (N_1261,In_288,N_1010);
or U1262 (N_1262,In_1365,In_1339);
xnor U1263 (N_1263,N_626,In_41);
xor U1264 (N_1264,N_309,In_315);
and U1265 (N_1265,N_1185,In_1900);
nand U1266 (N_1266,N_842,In_937);
or U1267 (N_1267,N_816,N_42);
nor U1268 (N_1268,N_612,N_1055);
nand U1269 (N_1269,In_1849,In_1945);
nor U1270 (N_1270,N_655,N_1069);
nand U1271 (N_1271,N_966,In_571);
xnor U1272 (N_1272,In_1749,N_615);
nand U1273 (N_1273,In_473,N_1095);
nor U1274 (N_1274,In_799,N_1176);
or U1275 (N_1275,In_332,In_1720);
and U1276 (N_1276,N_1046,N_361);
xor U1277 (N_1277,N_753,N_815);
nor U1278 (N_1278,N_744,N_926);
nor U1279 (N_1279,N_1078,In_962);
or U1280 (N_1280,N_301,N_1103);
nor U1281 (N_1281,N_1158,In_54);
nor U1282 (N_1282,N_1070,In_995);
and U1283 (N_1283,N_40,In_617);
and U1284 (N_1284,In_5,In_807);
and U1285 (N_1285,N_786,N_1051);
and U1286 (N_1286,N_1109,N_1041);
nor U1287 (N_1287,N_1157,N_850);
nor U1288 (N_1288,In_1284,N_868);
or U1289 (N_1289,N_1119,N_989);
or U1290 (N_1290,N_873,In_13);
xor U1291 (N_1291,N_418,In_619);
nand U1292 (N_1292,N_888,N_772);
and U1293 (N_1293,In_1263,N_549);
and U1294 (N_1294,N_171,N_553);
nand U1295 (N_1295,N_936,In_235);
nor U1296 (N_1296,N_613,N_911);
xnor U1297 (N_1297,N_20,N_730);
and U1298 (N_1298,N_974,N_303);
and U1299 (N_1299,In_592,N_957);
nand U1300 (N_1300,In_924,N_881);
nand U1301 (N_1301,N_576,N_196);
nand U1302 (N_1302,N_1191,N_636);
nor U1303 (N_1303,In_1694,In_1047);
xor U1304 (N_1304,N_929,N_1197);
and U1305 (N_1305,N_390,N_827);
nand U1306 (N_1306,N_714,N_1065);
or U1307 (N_1307,N_1018,In_1934);
xor U1308 (N_1308,In_474,N_429);
and U1309 (N_1309,N_1031,N_319);
nor U1310 (N_1310,N_226,N_964);
or U1311 (N_1311,N_566,In_348);
nand U1312 (N_1312,N_597,N_778);
nand U1313 (N_1313,In_1659,N_1047);
xnor U1314 (N_1314,N_762,N_103);
and U1315 (N_1315,In_1408,N_633);
nor U1316 (N_1316,In_1917,N_1181);
or U1317 (N_1317,N_1135,N_1101);
nand U1318 (N_1318,N_581,In_87);
nor U1319 (N_1319,N_1094,N_940);
xor U1320 (N_1320,N_1071,N_855);
nor U1321 (N_1321,N_992,N_758);
nor U1322 (N_1322,N_1091,N_900);
xor U1323 (N_1323,N_500,N_1171);
or U1324 (N_1324,N_864,N_1146);
nand U1325 (N_1325,N_628,N_1132);
or U1326 (N_1326,N_976,In_1585);
or U1327 (N_1327,N_970,N_1008);
nand U1328 (N_1328,N_421,In_476);
nor U1329 (N_1329,N_614,N_598);
nor U1330 (N_1330,In_170,N_1048);
xnor U1331 (N_1331,N_935,N_1011);
xor U1332 (N_1332,In_919,N_1142);
nor U1333 (N_1333,In_1343,In_391);
or U1334 (N_1334,In_1456,In_317);
xnor U1335 (N_1335,In_1948,In_1362);
nand U1336 (N_1336,In_1487,N_820);
nor U1337 (N_1337,In_965,In_1215);
xor U1338 (N_1338,N_1060,In_508);
nor U1339 (N_1339,N_1003,In_1427);
or U1340 (N_1340,N_733,In_40);
or U1341 (N_1341,N_1049,N_326);
or U1342 (N_1342,N_1180,N_1087);
and U1343 (N_1343,N_1023,N_625);
or U1344 (N_1344,N_1038,N_1098);
or U1345 (N_1345,N_1122,In_1474);
or U1346 (N_1346,N_735,In_1810);
and U1347 (N_1347,N_1024,N_1153);
nor U1348 (N_1348,N_883,In_896);
nand U1349 (N_1349,N_916,N_890);
xnor U1350 (N_1350,In_1429,N_1096);
xor U1351 (N_1351,N_321,N_968);
and U1352 (N_1352,N_254,N_825);
or U1353 (N_1353,N_5,N_1149);
or U1354 (N_1354,N_901,N_811);
xnor U1355 (N_1355,N_1100,N_1088);
or U1356 (N_1356,In_390,N_1160);
and U1357 (N_1357,N_1000,N_269);
xnor U1358 (N_1358,In_707,N_448);
nor U1359 (N_1359,In_285,N_739);
nand U1360 (N_1360,N_520,N_806);
and U1361 (N_1361,In_1223,N_771);
or U1362 (N_1362,N_1058,N_1089);
nor U1363 (N_1363,N_889,N_552);
nor U1364 (N_1364,In_1808,N_629);
xor U1365 (N_1365,N_843,N_287);
and U1366 (N_1366,N_652,N_1107);
nand U1367 (N_1367,In_1963,N_1118);
or U1368 (N_1368,N_998,In_1685);
nor U1369 (N_1369,N_488,N_1076);
nor U1370 (N_1370,N_763,N_63);
or U1371 (N_1371,N_958,N_844);
nor U1372 (N_1372,N_257,N_1144);
nand U1373 (N_1373,N_1092,N_1113);
or U1374 (N_1374,In_1953,N_1172);
and U1375 (N_1375,N_1174,N_1162);
xor U1376 (N_1376,N_657,In_513);
or U1377 (N_1377,In_964,In_1942);
xor U1378 (N_1378,In_767,N_459);
xor U1379 (N_1379,In_1449,N_1121);
xor U1380 (N_1380,N_751,In_144);
nor U1381 (N_1381,N_893,In_1206);
xnor U1382 (N_1382,N_414,In_752);
and U1383 (N_1383,N_1050,N_962);
nor U1384 (N_1384,N_1163,In_959);
xor U1385 (N_1385,N_932,In_1451);
nand U1386 (N_1386,N_1151,N_111);
nand U1387 (N_1387,N_1128,N_1090);
and U1388 (N_1388,N_1036,N_417);
nor U1389 (N_1389,N_1145,N_1086);
nand U1390 (N_1390,N_1110,N_724);
nand U1391 (N_1391,In_339,N_871);
xnor U1392 (N_1392,In_1045,N_443);
nand U1393 (N_1393,N_250,N_738);
or U1394 (N_1394,In_817,In_1245);
xor U1395 (N_1395,N_819,N_1039);
nor U1396 (N_1396,N_856,N_802);
xnor U1397 (N_1397,N_539,In_639);
xor U1398 (N_1398,N_606,N_727);
and U1399 (N_1399,In_1127,N_1117);
and U1400 (N_1400,N_984,N_947);
nor U1401 (N_1401,In_820,N_1184);
or U1402 (N_1402,N_1334,N_1355);
xor U1403 (N_1403,In_163,N_1356);
xor U1404 (N_1404,N_1261,N_877);
xor U1405 (N_1405,N_1319,N_1277);
xnor U1406 (N_1406,In_327,N_1085);
and U1407 (N_1407,N_1120,N_378);
or U1408 (N_1408,In_42,N_1136);
nand U1409 (N_1409,N_1188,N_1006);
nor U1410 (N_1410,N_1307,In_1678);
nor U1411 (N_1411,N_1192,N_1073);
nand U1412 (N_1412,N_1295,N_971);
and U1413 (N_1413,N_1308,In_837);
xor U1414 (N_1414,N_1170,N_1328);
or U1415 (N_1415,N_814,N_1243);
nand U1416 (N_1416,In_1397,N_454);
nor U1417 (N_1417,N_590,N_1327);
xor U1418 (N_1418,N_1316,In_1802);
or U1419 (N_1419,N_829,In_389);
nand U1420 (N_1420,N_845,N_1125);
nand U1421 (N_1421,N_1017,N_1235);
xor U1422 (N_1422,In_1669,N_1231);
xnor U1423 (N_1423,N_1375,N_1124);
nor U1424 (N_1424,N_1239,N_1126);
and U1425 (N_1425,In_53,In_768);
or U1426 (N_1426,N_732,N_874);
and U1427 (N_1427,N_965,In_1714);
and U1428 (N_1428,N_1229,In_20);
nor U1429 (N_1429,N_1363,N_1266);
xnor U1430 (N_1430,N_1338,N_767);
xor U1431 (N_1431,N_318,In_760);
or U1432 (N_1432,N_1028,N_986);
and U1433 (N_1433,N_923,N_854);
or U1434 (N_1434,N_1020,N_1081);
nor U1435 (N_1435,N_1253,N_193);
nand U1436 (N_1436,N_1269,In_543);
or U1437 (N_1437,N_822,N_1270);
nand U1438 (N_1438,N_83,N_543);
nor U1439 (N_1439,N_91,N_438);
or U1440 (N_1440,N_1116,N_1284);
xor U1441 (N_1441,N_1044,N_245);
nand U1442 (N_1442,N_757,In_800);
xor U1443 (N_1443,N_1156,N_1189);
and U1444 (N_1444,N_830,In_1232);
nand U1445 (N_1445,In_790,N_1102);
and U1446 (N_1446,N_773,N_1298);
nor U1447 (N_1447,N_919,In_1522);
nor U1448 (N_1448,N_1264,N_810);
and U1449 (N_1449,N_1329,N_809);
and U1450 (N_1450,N_1115,N_1140);
and U1451 (N_1451,N_1354,N_402);
or U1452 (N_1452,N_1336,In_920);
xnor U1453 (N_1453,N_1337,N_1164);
nor U1454 (N_1454,N_1238,N_1379);
nor U1455 (N_1455,N_1265,N_1240);
or U1456 (N_1456,N_1005,N_1285);
and U1457 (N_1457,N_1159,In_868);
nand U1458 (N_1458,In_1664,N_1317);
and U1459 (N_1459,N_717,N_635);
nand U1460 (N_1460,N_1224,N_406);
nand U1461 (N_1461,N_1177,N_1395);
xnor U1462 (N_1462,N_339,N_1205);
nand U1463 (N_1463,N_795,In_67);
nand U1464 (N_1464,N_813,N_1358);
and U1465 (N_1465,N_1173,N_1077);
xor U1466 (N_1466,N_3,N_1272);
nor U1467 (N_1467,N_1349,N_934);
nand U1468 (N_1468,N_1370,N_1009);
nand U1469 (N_1469,N_1385,In_683);
xor U1470 (N_1470,In_1054,N_1310);
xor U1471 (N_1471,N_1399,N_1226);
and U1472 (N_1472,N_1263,N_1234);
nand U1473 (N_1473,In_587,N_419);
nand U1474 (N_1474,N_1343,N_1382);
and U1475 (N_1475,N_1383,In_947);
nand U1476 (N_1476,In_92,N_804);
xnor U1477 (N_1477,N_1255,N_1154);
xor U1478 (N_1478,N_1384,N_1052);
or U1479 (N_1479,N_972,In_1950);
or U1480 (N_1480,N_1396,N_413);
and U1481 (N_1481,N_1271,In_240);
and U1482 (N_1482,N_1216,In_1918);
or U1483 (N_1483,In_1431,N_1199);
nor U1484 (N_1484,N_1309,N_1134);
and U1485 (N_1485,In_736,N_508);
or U1486 (N_1486,N_1360,N_457);
xor U1487 (N_1487,N_572,N_1378);
nand U1488 (N_1488,N_892,N_959);
nand U1489 (N_1489,N_803,N_1002);
nand U1490 (N_1490,N_979,N_690);
xnor U1491 (N_1491,N_1381,In_1586);
nand U1492 (N_1492,In_260,In_193);
and U1493 (N_1493,N_656,N_747);
and U1494 (N_1494,In_355,N_1323);
xnor U1495 (N_1495,N_1305,N_1391);
nor U1496 (N_1496,N_1315,N_1074);
and U1497 (N_1497,N_577,N_837);
nor U1498 (N_1498,N_1221,N_178);
and U1499 (N_1499,N_851,N_942);
nand U1500 (N_1500,N_18,In_1426);
xnor U1501 (N_1501,N_1340,N_1368);
or U1502 (N_1502,In_1509,N_461);
and U1503 (N_1503,In_645,N_1209);
nor U1504 (N_1504,In_1705,N_1213);
and U1505 (N_1505,N_1179,N_1293);
and U1506 (N_1506,N_787,In_1328);
nor U1507 (N_1507,N_1279,N_1034);
nor U1508 (N_1508,N_1251,N_1237);
nor U1509 (N_1509,N_1286,N_880);
nand U1510 (N_1510,N_1004,In_22);
or U1511 (N_1511,In_1305,N_1204);
or U1512 (N_1512,N_1274,N_1371);
xnor U1513 (N_1513,In_1061,N_1093);
and U1514 (N_1514,N_1275,In_1936);
and U1515 (N_1515,N_1304,N_1201);
and U1516 (N_1516,In_1111,N_238);
or U1517 (N_1517,N_182,N_1301);
or U1518 (N_1518,In_176,N_35);
or U1519 (N_1519,N_1325,N_1311);
or U1520 (N_1520,N_1331,N_1127);
and U1521 (N_1521,N_1053,N_734);
nor U1522 (N_1522,N_1099,N_988);
nand U1523 (N_1523,In_848,N_706);
and U1524 (N_1524,N_1290,N_185);
and U1525 (N_1525,N_1222,N_1359);
xor U1526 (N_1526,In_255,N_1241);
nor U1527 (N_1527,In_1153,N_1393);
or U1528 (N_1528,In_202,N_1392);
or U1529 (N_1529,N_1186,N_1022);
nand U1530 (N_1530,N_191,N_1208);
and U1531 (N_1531,N_1394,In_830);
xor U1532 (N_1532,N_53,N_1026);
nor U1533 (N_1533,In_1846,N_1068);
nand U1534 (N_1534,N_781,In_846);
xor U1535 (N_1535,N_902,N_1106);
xnor U1536 (N_1536,N_114,In_551);
nor U1537 (N_1537,N_627,N_1357);
nand U1538 (N_1538,N_1248,In_102);
nand U1539 (N_1539,N_765,N_885);
nor U1540 (N_1540,N_1377,In_36);
nand U1541 (N_1541,N_573,N_1278);
and U1542 (N_1542,In_1086,N_1244);
nor U1543 (N_1543,In_114,N_1350);
xnor U1544 (N_1544,N_1380,N_896);
xnor U1545 (N_1545,N_164,N_1312);
or U1546 (N_1546,N_237,N_832);
xor U1547 (N_1547,In_79,In_1717);
xor U1548 (N_1548,N_1014,N_623);
nand U1549 (N_1549,N_801,In_142);
xnor U1550 (N_1550,N_928,N_1062);
nand U1551 (N_1551,N_1398,N_1219);
and U1552 (N_1552,N_991,N_1376);
nor U1553 (N_1553,N_575,In_823);
nor U1554 (N_1554,N_1138,N_1037);
and U1555 (N_1555,In_239,N_1236);
and U1556 (N_1556,In_213,N_1150);
xor U1557 (N_1557,N_1227,N_1223);
nand U1558 (N_1558,N_1297,N_1082);
nor U1559 (N_1559,In_1527,N_230);
and U1560 (N_1560,N_711,N_432);
nor U1561 (N_1561,In_1372,N_1339);
nand U1562 (N_1562,N_1303,N_1063);
and U1563 (N_1563,N_541,N_1152);
nor U1564 (N_1564,N_1193,In_151);
nor U1565 (N_1565,N_1035,In_1611);
nor U1566 (N_1566,N_1001,N_1372);
or U1567 (N_1567,N_1043,N_857);
or U1568 (N_1568,N_1299,N_1007);
or U1569 (N_1569,In_1612,N_256);
xor U1570 (N_1570,N_1198,In_1512);
or U1571 (N_1571,N_1233,In_668);
nand U1572 (N_1572,N_1361,N_1321);
or U1573 (N_1573,In_1114,In_535);
xor U1574 (N_1574,In_1915,N_534);
nor U1575 (N_1575,N_867,N_1175);
xor U1576 (N_1576,N_1256,N_447);
or U1577 (N_1577,N_1333,N_1281);
nand U1578 (N_1578,N_983,In_465);
nand U1579 (N_1579,In_1360,N_1030);
nor U1580 (N_1580,N_1314,N_1313);
or U1581 (N_1581,N_687,In_825);
nand U1582 (N_1582,N_219,N_741);
xor U1583 (N_1583,N_969,N_826);
nor U1584 (N_1584,N_1210,N_884);
nor U1585 (N_1585,In_835,N_994);
xnor U1586 (N_1586,In_692,N_618);
or U1587 (N_1587,N_866,N_1374);
and U1588 (N_1588,In_491,N_728);
or U1589 (N_1589,N_1306,N_1280);
nand U1590 (N_1590,N_1168,N_1212);
xnor U1591 (N_1591,N_1351,N_840);
or U1592 (N_1592,In_798,N_1230);
xnor U1593 (N_1593,N_1347,In_340);
and U1594 (N_1594,N_1254,N_1353);
nor U1595 (N_1595,N_1207,In_1639);
or U1596 (N_1596,N_905,N_1362);
xnor U1597 (N_1597,In_1143,N_1318);
and U1598 (N_1598,N_954,N_1397);
xnor U1599 (N_1599,N_1066,N_1366);
nor U1600 (N_1600,N_1345,N_1489);
nor U1601 (N_1601,N_941,N_1445);
nand U1602 (N_1602,N_1503,In_147);
or U1603 (N_1603,N_1400,N_1225);
nor U1604 (N_1604,N_1499,N_1324);
nor U1605 (N_1605,N_1326,N_1543);
nand U1606 (N_1606,In_1823,N_1516);
nand U1607 (N_1607,In_1402,N_1508);
xnor U1608 (N_1608,N_1527,N_1013);
nor U1609 (N_1609,N_399,N_1463);
and U1610 (N_1610,N_1407,N_1488);
xor U1611 (N_1611,N_1585,N_1518);
xor U1612 (N_1612,N_1481,In_967);
nor U1613 (N_1613,N_1515,N_1389);
nand U1614 (N_1614,In_1347,N_1509);
xor U1615 (N_1615,N_1129,N_1536);
nor U1616 (N_1616,N_1411,In_567);
nand U1617 (N_1617,N_1547,N_1459);
and U1618 (N_1618,N_1486,N_515);
xnor U1619 (N_1619,N_1572,N_1564);
and U1620 (N_1620,N_1032,N_1420);
and U1621 (N_1621,N_907,N_1206);
and U1622 (N_1622,N_1414,N_1418);
nor U1623 (N_1623,N_715,N_1438);
nand U1624 (N_1624,N_1139,In_1166);
and U1625 (N_1625,N_927,N_1545);
xnor U1626 (N_1626,N_1507,N_1511);
xnor U1627 (N_1627,N_1451,N_1405);
or U1628 (N_1628,In_305,N_1195);
nor U1629 (N_1629,N_1531,N_1322);
nor U1630 (N_1630,N_1458,N_1415);
xnor U1631 (N_1631,N_1341,In_1761);
nand U1632 (N_1632,N_1402,N_1571);
and U1633 (N_1633,In_612,N_1015);
nor U1634 (N_1634,In_512,In_1643);
nor U1635 (N_1635,N_736,N_1524);
and U1636 (N_1636,N_1534,N_1302);
xnor U1637 (N_1637,N_1080,N_1196);
xnor U1638 (N_1638,N_1523,N_1583);
or U1639 (N_1639,N_1567,N_1448);
nand U1640 (N_1640,N_1447,N_887);
nand U1641 (N_1641,N_712,N_1498);
or U1642 (N_1642,N_1166,N_1465);
nor U1643 (N_1643,N_1483,N_1273);
nor U1644 (N_1644,N_1570,N_1369);
nand U1645 (N_1645,N_446,N_1586);
xor U1646 (N_1646,N_776,N_698);
and U1647 (N_1647,N_1590,N_1067);
or U1648 (N_1648,N_1517,N_1470);
nor U1649 (N_1649,N_1412,N_1423);
nor U1650 (N_1650,N_1436,N_1582);
nand U1651 (N_1651,N_1473,N_1596);
nand U1652 (N_1652,N_1344,N_1373);
xnor U1653 (N_1653,N_1259,N_624);
nor U1654 (N_1654,N_1267,N_1442);
xor U1655 (N_1655,In_1713,N_1548);
nor U1656 (N_1656,In_1750,N_1565);
and U1657 (N_1657,N_1578,In_1526);
xnor U1658 (N_1658,In_162,N_117);
or U1659 (N_1659,N_1476,N_1584);
nor U1660 (N_1660,N_1550,N_1455);
or U1661 (N_1661,N_1480,N_1282);
or U1662 (N_1662,N_1202,N_1403);
and U1663 (N_1663,N_1533,In_1916);
nor U1664 (N_1664,N_1549,N_1539);
nor U1665 (N_1665,N_1577,N_1246);
nand U1666 (N_1666,N_1587,N_1413);
nand U1667 (N_1667,N_1514,N_1544);
nor U1668 (N_1668,N_1477,N_1563);
nand U1669 (N_1669,N_1388,N_1592);
xnor U1670 (N_1670,N_1519,N_1528);
nand U1671 (N_1671,N_1183,N_1594);
nor U1672 (N_1672,N_1367,N_1540);
and U1673 (N_1673,N_1453,N_1203);
nand U1674 (N_1674,N_1551,N_1579);
xnor U1675 (N_1675,N_1462,N_1072);
nor U1676 (N_1676,N_1490,N_513);
or U1677 (N_1677,N_1252,N_1581);
xnor U1678 (N_1678,N_1141,N_1187);
and U1679 (N_1679,N_1342,N_666);
nand U1680 (N_1680,N_537,N_588);
nor U1681 (N_1681,N_271,N_1482);
nor U1682 (N_1682,N_1214,N_1332);
xor U1683 (N_1683,N_1546,N_1364);
or U1684 (N_1684,N_187,N_1575);
xnor U1685 (N_1685,N_1218,N_1496);
nand U1686 (N_1686,N_680,In_135);
xnor U1687 (N_1687,N_710,N_1296);
or U1688 (N_1688,N_1541,In_1367);
nor U1689 (N_1689,N_1472,N_1439);
nand U1690 (N_1690,N_1365,N_1215);
xnor U1691 (N_1691,N_1487,N_1268);
xor U1692 (N_1692,N_1537,N_1446);
and U1693 (N_1693,N_1220,N_1484);
xnor U1694 (N_1694,N_1555,N_1424);
or U1695 (N_1695,N_939,N_1471);
and U1696 (N_1696,N_1468,N_84);
or U1697 (N_1697,In_311,N_1538);
nand U1698 (N_1698,In_1536,N_1466);
or U1699 (N_1699,N_1408,N_1475);
xor U1700 (N_1700,N_1123,N_601);
nor U1701 (N_1701,N_1434,In_1395);
or U1702 (N_1702,N_876,N_1291);
xnor U1703 (N_1703,N_997,In_1514);
nand U1704 (N_1704,In_1733,N_1283);
nand U1705 (N_1705,In_1256,N_1429);
nor U1706 (N_1706,N_1294,N_1491);
and U1707 (N_1707,N_327,N_1430);
or U1708 (N_1708,N_1200,N_1242);
nor U1709 (N_1709,In_1198,N_426);
xnor U1710 (N_1710,In_1501,N_357);
xnor U1711 (N_1711,N_1444,In_1342);
or U1712 (N_1712,N_1588,N_501);
or U1713 (N_1713,N_1330,N_1292);
or U1714 (N_1714,In_1391,N_1474);
nor U1715 (N_1715,N_502,N_1530);
nand U1716 (N_1716,N_1165,N_56);
nor U1717 (N_1717,N_1559,N_663);
and U1718 (N_1718,In_1200,N_1493);
nand U1719 (N_1719,N_1217,N_1469);
nand U1720 (N_1720,N_1452,In_998);
or U1721 (N_1721,In_1635,In_1462);
nor U1722 (N_1722,In_1584,N_1574);
xor U1723 (N_1723,N_1561,N_1566);
xor U1724 (N_1724,N_139,N_1300);
nand U1725 (N_1725,N_1335,N_1525);
xnor U1726 (N_1726,N_1464,N_1556);
nand U1727 (N_1727,N_1211,N_1130);
or U1728 (N_1728,N_1428,N_1409);
nor U1729 (N_1729,In_664,N_1591);
xnor U1730 (N_1730,N_1598,N_1522);
xor U1731 (N_1731,N_1542,In_1271);
nor U1732 (N_1732,N_1532,In_385);
and U1733 (N_1733,N_1456,N_920);
nor U1734 (N_1734,In_737,N_1416);
nor U1735 (N_1735,N_1348,N_1262);
xor U1736 (N_1736,N_1506,N_403);
or U1737 (N_1737,N_897,N_1479);
and U1738 (N_1738,N_1593,In_1881);
xnor U1739 (N_1739,In_1547,N_1386);
xnor U1740 (N_1740,N_1485,N_1497);
xnor U1741 (N_1741,N_1513,In_561);
nor U1742 (N_1742,In_977,N_1169);
nand U1743 (N_1743,N_1417,N_1521);
nor U1744 (N_1744,N_1320,N_1057);
xnor U1745 (N_1745,N_1558,N_1404);
or U1746 (N_1746,N_1426,N_1597);
nand U1747 (N_1747,In_121,N_1569);
and U1748 (N_1748,N_1501,N_1390);
and U1749 (N_1749,N_1449,N_1580);
xnor U1750 (N_1750,N_1520,In_1322);
xor U1751 (N_1751,N_796,N_642);
nor U1752 (N_1752,N_1589,N_1425);
xnor U1753 (N_1753,N_1554,N_933);
and U1754 (N_1754,N_1287,In_1655);
nor U1755 (N_1755,N_1557,In_1084);
and U1756 (N_1756,N_1510,N_1401);
xnor U1757 (N_1757,N_1056,In_970);
nor U1758 (N_1758,N_600,N_1553);
nor U1759 (N_1759,N_1289,N_1535);
and U1760 (N_1760,N_1245,N_1054);
xnor U1761 (N_1761,N_1562,In_1162);
nand U1762 (N_1762,N_1595,N_1155);
or U1763 (N_1763,N_1257,N_1568);
or U1764 (N_1764,N_1495,N_1478);
nor U1765 (N_1765,N_1346,N_1108);
xor U1766 (N_1766,N_1494,N_1492);
xnor U1767 (N_1767,N_1387,N_1467);
or U1768 (N_1768,In_842,N_1137);
nor U1769 (N_1769,N_1437,N_255);
xnor U1770 (N_1770,N_1352,N_1460);
and U1771 (N_1771,In_190,N_1276);
nand U1772 (N_1772,N_1573,N_1247);
or U1773 (N_1773,N_1526,N_1576);
or U1774 (N_1774,In_660,N_1432);
nand U1775 (N_1775,N_1250,N_1443);
and U1776 (N_1776,N_1500,N_1410);
nor U1777 (N_1777,N_1505,N_1260);
and U1778 (N_1778,N_1232,In_302);
nor U1779 (N_1779,N_1457,N_661);
xnor U1780 (N_1780,N_1512,N_1427);
nor U1781 (N_1781,N_1228,N_1440);
and U1782 (N_1782,N_1025,N_1161);
nor U1783 (N_1783,N_909,N_980);
xor U1784 (N_1784,In_218,N_1560);
xor U1785 (N_1785,N_1421,N_750);
xor U1786 (N_1786,N_1461,N_1419);
nor U1787 (N_1787,N_1249,N_1504);
or U1788 (N_1788,In_917,N_1422);
nor U1789 (N_1789,In_715,N_1431);
nand U1790 (N_1790,N_658,N_1502);
xnor U1791 (N_1791,N_1454,N_1433);
and U1792 (N_1792,N_1435,N_838);
and U1793 (N_1793,N_1599,N_1029);
or U1794 (N_1794,N_1288,N_1083);
xor U1795 (N_1795,In_313,N_1450);
nand U1796 (N_1796,N_1529,N_1258);
xor U1797 (N_1797,In_55,N_1441);
or U1798 (N_1798,N_1143,In_1141);
and U1799 (N_1799,N_1406,N_1552);
xnor U1800 (N_1800,N_1711,N_1708);
and U1801 (N_1801,N_1752,N_1778);
nand U1802 (N_1802,N_1625,N_1654);
xnor U1803 (N_1803,N_1783,N_1730);
nor U1804 (N_1804,N_1723,N_1615);
nand U1805 (N_1805,N_1734,N_1640);
nor U1806 (N_1806,N_1683,N_1685);
xor U1807 (N_1807,N_1728,N_1756);
nand U1808 (N_1808,N_1686,N_1620);
or U1809 (N_1809,N_1697,N_1714);
nand U1810 (N_1810,N_1797,N_1786);
nand U1811 (N_1811,N_1757,N_1603);
or U1812 (N_1812,N_1624,N_1762);
or U1813 (N_1813,N_1767,N_1609);
xor U1814 (N_1814,N_1789,N_1736);
nor U1815 (N_1815,N_1785,N_1675);
nor U1816 (N_1816,N_1680,N_1749);
nand U1817 (N_1817,N_1692,N_1623);
xnor U1818 (N_1818,N_1776,N_1769);
or U1819 (N_1819,N_1798,N_1629);
nor U1820 (N_1820,N_1606,N_1662);
nor U1821 (N_1821,N_1733,N_1722);
nand U1822 (N_1822,N_1780,N_1658);
nor U1823 (N_1823,N_1731,N_1691);
xnor U1824 (N_1824,N_1725,N_1715);
and U1825 (N_1825,N_1792,N_1755);
and U1826 (N_1826,N_1706,N_1735);
or U1827 (N_1827,N_1741,N_1684);
and U1828 (N_1828,N_1775,N_1677);
xor U1829 (N_1829,N_1648,N_1637);
nor U1830 (N_1830,N_1643,N_1652);
or U1831 (N_1831,N_1724,N_1764);
nand U1832 (N_1832,N_1740,N_1768);
or U1833 (N_1833,N_1721,N_1777);
nand U1834 (N_1834,N_1617,N_1698);
or U1835 (N_1835,N_1754,N_1613);
or U1836 (N_1836,N_1701,N_1653);
and U1837 (N_1837,N_1744,N_1667);
or U1838 (N_1838,N_1699,N_1634);
or U1839 (N_1839,N_1737,N_1717);
or U1840 (N_1840,N_1738,N_1642);
or U1841 (N_1841,N_1663,N_1716);
and U1842 (N_1842,N_1784,N_1753);
nor U1843 (N_1843,N_1751,N_1618);
nor U1844 (N_1844,N_1622,N_1670);
and U1845 (N_1845,N_1781,N_1612);
nand U1846 (N_1846,N_1782,N_1687);
nand U1847 (N_1847,N_1705,N_1668);
xor U1848 (N_1848,N_1664,N_1743);
or U1849 (N_1849,N_1682,N_1770);
nor U1850 (N_1850,N_1616,N_1674);
or U1851 (N_1851,N_1633,N_1679);
or U1852 (N_1852,N_1689,N_1600);
nor U1853 (N_1853,N_1626,N_1796);
nand U1854 (N_1854,N_1759,N_1621);
nor U1855 (N_1855,N_1638,N_1678);
or U1856 (N_1856,N_1619,N_1688);
nand U1857 (N_1857,N_1646,N_1660);
and U1858 (N_1858,N_1631,N_1773);
nand U1859 (N_1859,N_1774,N_1604);
and U1860 (N_1860,N_1729,N_1702);
nor U1861 (N_1861,N_1709,N_1611);
nand U1862 (N_1862,N_1742,N_1700);
or U1863 (N_1863,N_1694,N_1710);
nand U1864 (N_1864,N_1748,N_1665);
or U1865 (N_1865,N_1632,N_1788);
nand U1866 (N_1866,N_1681,N_1732);
or U1867 (N_1867,N_1791,N_1790);
nand U1868 (N_1868,N_1639,N_1645);
or U1869 (N_1869,N_1727,N_1760);
xnor U1870 (N_1870,N_1713,N_1628);
nor U1871 (N_1871,N_1779,N_1766);
xor U1872 (N_1872,N_1644,N_1795);
and U1873 (N_1873,N_1747,N_1671);
or U1874 (N_1874,N_1690,N_1794);
nand U1875 (N_1875,N_1647,N_1676);
nand U1876 (N_1876,N_1787,N_1650);
nand U1877 (N_1877,N_1669,N_1719);
and U1878 (N_1878,N_1630,N_1771);
or U1879 (N_1879,N_1793,N_1746);
nand U1880 (N_1880,N_1720,N_1695);
xnor U1881 (N_1881,N_1673,N_1696);
or U1882 (N_1882,N_1651,N_1739);
xor U1883 (N_1883,N_1758,N_1602);
and U1884 (N_1884,N_1635,N_1656);
xnor U1885 (N_1885,N_1707,N_1750);
xnor U1886 (N_1886,N_1627,N_1763);
or U1887 (N_1887,N_1718,N_1649);
and U1888 (N_1888,N_1657,N_1614);
and U1889 (N_1889,N_1772,N_1693);
or U1890 (N_1890,N_1745,N_1672);
nor U1891 (N_1891,N_1761,N_1799);
and U1892 (N_1892,N_1607,N_1610);
xor U1893 (N_1893,N_1726,N_1659);
xnor U1894 (N_1894,N_1703,N_1608);
and U1895 (N_1895,N_1661,N_1641);
nand U1896 (N_1896,N_1655,N_1765);
or U1897 (N_1897,N_1712,N_1636);
nor U1898 (N_1898,N_1666,N_1601);
xnor U1899 (N_1899,N_1704,N_1605);
nor U1900 (N_1900,N_1737,N_1611);
nand U1901 (N_1901,N_1742,N_1793);
xor U1902 (N_1902,N_1606,N_1659);
and U1903 (N_1903,N_1732,N_1604);
nor U1904 (N_1904,N_1744,N_1673);
or U1905 (N_1905,N_1625,N_1688);
nand U1906 (N_1906,N_1617,N_1648);
or U1907 (N_1907,N_1759,N_1735);
xnor U1908 (N_1908,N_1796,N_1607);
nand U1909 (N_1909,N_1697,N_1613);
xor U1910 (N_1910,N_1715,N_1632);
nor U1911 (N_1911,N_1707,N_1677);
xnor U1912 (N_1912,N_1656,N_1794);
or U1913 (N_1913,N_1794,N_1715);
nor U1914 (N_1914,N_1714,N_1648);
or U1915 (N_1915,N_1777,N_1699);
nor U1916 (N_1916,N_1759,N_1793);
xor U1917 (N_1917,N_1738,N_1796);
nor U1918 (N_1918,N_1742,N_1711);
nor U1919 (N_1919,N_1653,N_1792);
nand U1920 (N_1920,N_1639,N_1791);
and U1921 (N_1921,N_1626,N_1612);
xor U1922 (N_1922,N_1784,N_1694);
nand U1923 (N_1923,N_1684,N_1698);
nor U1924 (N_1924,N_1653,N_1615);
nand U1925 (N_1925,N_1759,N_1601);
or U1926 (N_1926,N_1601,N_1783);
and U1927 (N_1927,N_1675,N_1732);
or U1928 (N_1928,N_1761,N_1653);
xnor U1929 (N_1929,N_1680,N_1621);
nor U1930 (N_1930,N_1617,N_1692);
xor U1931 (N_1931,N_1764,N_1657);
or U1932 (N_1932,N_1644,N_1787);
nand U1933 (N_1933,N_1652,N_1737);
nor U1934 (N_1934,N_1670,N_1723);
nor U1935 (N_1935,N_1638,N_1748);
and U1936 (N_1936,N_1787,N_1657);
or U1937 (N_1937,N_1770,N_1686);
nor U1938 (N_1938,N_1608,N_1601);
nor U1939 (N_1939,N_1742,N_1632);
xnor U1940 (N_1940,N_1617,N_1788);
or U1941 (N_1941,N_1749,N_1733);
or U1942 (N_1942,N_1702,N_1768);
nor U1943 (N_1943,N_1706,N_1769);
xor U1944 (N_1944,N_1745,N_1737);
or U1945 (N_1945,N_1682,N_1780);
or U1946 (N_1946,N_1669,N_1632);
and U1947 (N_1947,N_1748,N_1611);
or U1948 (N_1948,N_1771,N_1643);
and U1949 (N_1949,N_1633,N_1632);
nor U1950 (N_1950,N_1634,N_1675);
nand U1951 (N_1951,N_1682,N_1659);
or U1952 (N_1952,N_1639,N_1615);
xor U1953 (N_1953,N_1608,N_1698);
nand U1954 (N_1954,N_1675,N_1658);
nand U1955 (N_1955,N_1792,N_1726);
nor U1956 (N_1956,N_1777,N_1746);
nor U1957 (N_1957,N_1769,N_1765);
or U1958 (N_1958,N_1703,N_1646);
xnor U1959 (N_1959,N_1656,N_1762);
nor U1960 (N_1960,N_1780,N_1751);
xnor U1961 (N_1961,N_1780,N_1640);
or U1962 (N_1962,N_1737,N_1697);
xor U1963 (N_1963,N_1693,N_1642);
nand U1964 (N_1964,N_1785,N_1672);
and U1965 (N_1965,N_1758,N_1789);
xor U1966 (N_1966,N_1643,N_1671);
xnor U1967 (N_1967,N_1725,N_1658);
or U1968 (N_1968,N_1768,N_1640);
and U1969 (N_1969,N_1631,N_1764);
xor U1970 (N_1970,N_1734,N_1641);
and U1971 (N_1971,N_1690,N_1723);
or U1972 (N_1972,N_1652,N_1719);
nand U1973 (N_1973,N_1721,N_1684);
or U1974 (N_1974,N_1630,N_1617);
xnor U1975 (N_1975,N_1785,N_1775);
or U1976 (N_1976,N_1738,N_1655);
nand U1977 (N_1977,N_1757,N_1758);
nor U1978 (N_1978,N_1641,N_1662);
xnor U1979 (N_1979,N_1605,N_1650);
and U1980 (N_1980,N_1653,N_1770);
nor U1981 (N_1981,N_1613,N_1619);
nor U1982 (N_1982,N_1697,N_1600);
nand U1983 (N_1983,N_1639,N_1759);
nand U1984 (N_1984,N_1696,N_1612);
nor U1985 (N_1985,N_1786,N_1606);
nand U1986 (N_1986,N_1701,N_1692);
xor U1987 (N_1987,N_1723,N_1724);
nand U1988 (N_1988,N_1720,N_1652);
xnor U1989 (N_1989,N_1732,N_1658);
or U1990 (N_1990,N_1696,N_1715);
nor U1991 (N_1991,N_1697,N_1705);
and U1992 (N_1992,N_1770,N_1626);
and U1993 (N_1993,N_1662,N_1795);
or U1994 (N_1994,N_1781,N_1631);
or U1995 (N_1995,N_1792,N_1710);
xnor U1996 (N_1996,N_1780,N_1790);
and U1997 (N_1997,N_1768,N_1767);
nor U1998 (N_1998,N_1613,N_1672);
and U1999 (N_1999,N_1776,N_1796);
xnor U2000 (N_2000,N_1924,N_1962);
or U2001 (N_2001,N_1919,N_1952);
nand U2002 (N_2002,N_1928,N_1845);
xnor U2003 (N_2003,N_1875,N_1906);
xnor U2004 (N_2004,N_1802,N_1892);
nor U2005 (N_2005,N_1968,N_1812);
nand U2006 (N_2006,N_1997,N_1852);
and U2007 (N_2007,N_1827,N_1933);
or U2008 (N_2008,N_1832,N_1823);
or U2009 (N_2009,N_1903,N_1816);
and U2010 (N_2010,N_1958,N_1927);
xor U2011 (N_2011,N_1993,N_1831);
or U2012 (N_2012,N_1841,N_1806);
and U2013 (N_2013,N_1972,N_1946);
nand U2014 (N_2014,N_1964,N_1822);
nor U2015 (N_2015,N_1929,N_1884);
nor U2016 (N_2016,N_1874,N_1922);
xnor U2017 (N_2017,N_1820,N_1811);
nand U2018 (N_2018,N_1911,N_1848);
xor U2019 (N_2019,N_1853,N_1926);
nor U2020 (N_2020,N_1861,N_1866);
or U2021 (N_2021,N_1970,N_1881);
nand U2022 (N_2022,N_1979,N_1982);
xnor U2023 (N_2023,N_1809,N_1818);
or U2024 (N_2024,N_1954,N_1967);
nand U2025 (N_2025,N_1838,N_1961);
xnor U2026 (N_2026,N_1830,N_1920);
nor U2027 (N_2027,N_1888,N_1857);
nor U2028 (N_2028,N_1963,N_1956);
nor U2029 (N_2029,N_1902,N_1896);
or U2030 (N_2030,N_1807,N_1869);
xnor U2031 (N_2031,N_1989,N_1978);
nor U2032 (N_2032,N_1883,N_1940);
xnor U2033 (N_2033,N_1873,N_1951);
nor U2034 (N_2034,N_1905,N_1817);
or U2035 (N_2035,N_1834,N_1897);
nor U2036 (N_2036,N_1935,N_1813);
xnor U2037 (N_2037,N_1959,N_1858);
and U2038 (N_2038,N_1991,N_1942);
xnor U2039 (N_2039,N_1829,N_1988);
or U2040 (N_2040,N_1870,N_1901);
or U2041 (N_2041,N_1990,N_1994);
and U2042 (N_2042,N_1850,N_1981);
xnor U2043 (N_2043,N_1871,N_1980);
or U2044 (N_2044,N_1899,N_1907);
and U2045 (N_2045,N_1863,N_1868);
xnor U2046 (N_2046,N_1984,N_1879);
nor U2047 (N_2047,N_1810,N_1908);
and U2048 (N_2048,N_1955,N_1937);
nand U2049 (N_2049,N_1893,N_1814);
and U2050 (N_2050,N_1965,N_1925);
and U2051 (N_2051,N_1859,N_1886);
nand U2052 (N_2052,N_1918,N_1969);
nor U2053 (N_2053,N_1999,N_1915);
xor U2054 (N_2054,N_1900,N_1880);
and U2055 (N_2055,N_1916,N_1801);
nand U2056 (N_2056,N_1949,N_1844);
or U2057 (N_2057,N_1843,N_1932);
nand U2058 (N_2058,N_1931,N_1953);
nor U2059 (N_2059,N_1890,N_1862);
xor U2060 (N_2060,N_1891,N_1912);
or U2061 (N_2061,N_1914,N_1808);
nand U2062 (N_2062,N_1995,N_1950);
or U2063 (N_2063,N_1977,N_1986);
nor U2064 (N_2064,N_1889,N_1957);
nor U2065 (N_2065,N_1960,N_1936);
nor U2066 (N_2066,N_1847,N_1998);
or U2067 (N_2067,N_1882,N_1872);
nor U2068 (N_2068,N_1887,N_1839);
nand U2069 (N_2069,N_1948,N_1815);
and U2070 (N_2070,N_1909,N_1944);
and U2071 (N_2071,N_1849,N_1835);
nor U2072 (N_2072,N_1885,N_1913);
xor U2073 (N_2073,N_1846,N_1828);
and U2074 (N_2074,N_1974,N_1939);
nand U2075 (N_2075,N_1864,N_1966);
nor U2076 (N_2076,N_1923,N_1855);
xor U2077 (N_2077,N_1865,N_1856);
xor U2078 (N_2078,N_1917,N_1973);
nor U2079 (N_2079,N_1910,N_1840);
and U2080 (N_2080,N_1983,N_1943);
or U2081 (N_2081,N_1992,N_1867);
nor U2082 (N_2082,N_1985,N_1826);
xnor U2083 (N_2083,N_1842,N_1800);
nand U2084 (N_2084,N_1860,N_1876);
nor U2085 (N_2085,N_1805,N_1976);
xnor U2086 (N_2086,N_1851,N_1930);
or U2087 (N_2087,N_1947,N_1904);
and U2088 (N_2088,N_1941,N_1996);
nand U2089 (N_2089,N_1878,N_1971);
or U2090 (N_2090,N_1824,N_1877);
and U2091 (N_2091,N_1821,N_1833);
nand U2092 (N_2092,N_1894,N_1934);
nor U2093 (N_2093,N_1836,N_1921);
or U2094 (N_2094,N_1819,N_1825);
nor U2095 (N_2095,N_1803,N_1898);
xor U2096 (N_2096,N_1837,N_1804);
or U2097 (N_2097,N_1987,N_1854);
nand U2098 (N_2098,N_1945,N_1895);
or U2099 (N_2099,N_1938,N_1975);
nor U2100 (N_2100,N_1946,N_1966);
nor U2101 (N_2101,N_1995,N_1962);
nand U2102 (N_2102,N_1955,N_1848);
nand U2103 (N_2103,N_1900,N_1951);
xnor U2104 (N_2104,N_1807,N_1912);
nor U2105 (N_2105,N_1850,N_1882);
or U2106 (N_2106,N_1906,N_1809);
nor U2107 (N_2107,N_1881,N_1924);
nand U2108 (N_2108,N_1850,N_1830);
xor U2109 (N_2109,N_1888,N_1900);
and U2110 (N_2110,N_1844,N_1953);
nand U2111 (N_2111,N_1820,N_1890);
nand U2112 (N_2112,N_1881,N_1853);
and U2113 (N_2113,N_1989,N_1998);
and U2114 (N_2114,N_1940,N_1870);
nor U2115 (N_2115,N_1978,N_1959);
nand U2116 (N_2116,N_1818,N_1896);
nand U2117 (N_2117,N_1865,N_1993);
nor U2118 (N_2118,N_1825,N_1893);
and U2119 (N_2119,N_1997,N_1845);
nand U2120 (N_2120,N_1967,N_1899);
nand U2121 (N_2121,N_1854,N_1884);
nor U2122 (N_2122,N_1824,N_1819);
and U2123 (N_2123,N_1971,N_1897);
nor U2124 (N_2124,N_1803,N_1891);
xor U2125 (N_2125,N_1929,N_1814);
nor U2126 (N_2126,N_1856,N_1904);
or U2127 (N_2127,N_1844,N_1836);
xor U2128 (N_2128,N_1972,N_1886);
and U2129 (N_2129,N_1926,N_1845);
or U2130 (N_2130,N_1908,N_1960);
nor U2131 (N_2131,N_1850,N_1859);
or U2132 (N_2132,N_1872,N_1887);
nor U2133 (N_2133,N_1949,N_1880);
nand U2134 (N_2134,N_1868,N_1915);
and U2135 (N_2135,N_1899,N_1885);
or U2136 (N_2136,N_1884,N_1958);
and U2137 (N_2137,N_1909,N_1837);
and U2138 (N_2138,N_1920,N_1867);
nor U2139 (N_2139,N_1961,N_1801);
xor U2140 (N_2140,N_1971,N_1927);
and U2141 (N_2141,N_1896,N_1873);
and U2142 (N_2142,N_1955,N_1869);
nand U2143 (N_2143,N_1813,N_1801);
xnor U2144 (N_2144,N_1840,N_1811);
nor U2145 (N_2145,N_1939,N_1899);
xnor U2146 (N_2146,N_1832,N_1822);
and U2147 (N_2147,N_1819,N_1992);
nand U2148 (N_2148,N_1901,N_1861);
xnor U2149 (N_2149,N_1849,N_1902);
xnor U2150 (N_2150,N_1890,N_1923);
and U2151 (N_2151,N_1956,N_1842);
or U2152 (N_2152,N_1956,N_1873);
nand U2153 (N_2153,N_1945,N_1866);
nor U2154 (N_2154,N_1994,N_1950);
xor U2155 (N_2155,N_1983,N_1847);
nor U2156 (N_2156,N_1974,N_1904);
or U2157 (N_2157,N_1803,N_1845);
nor U2158 (N_2158,N_1937,N_1888);
xor U2159 (N_2159,N_1876,N_1848);
and U2160 (N_2160,N_1843,N_1808);
or U2161 (N_2161,N_1966,N_1902);
nor U2162 (N_2162,N_1871,N_1998);
and U2163 (N_2163,N_1841,N_1884);
xor U2164 (N_2164,N_1829,N_1856);
nand U2165 (N_2165,N_1961,N_1822);
and U2166 (N_2166,N_1904,N_1954);
nand U2167 (N_2167,N_1843,N_1960);
nand U2168 (N_2168,N_1903,N_1951);
nor U2169 (N_2169,N_1997,N_1930);
xor U2170 (N_2170,N_1866,N_1823);
or U2171 (N_2171,N_1911,N_1806);
and U2172 (N_2172,N_1812,N_1945);
and U2173 (N_2173,N_1936,N_1812);
nor U2174 (N_2174,N_1846,N_1994);
or U2175 (N_2175,N_1892,N_1831);
nand U2176 (N_2176,N_1826,N_1969);
or U2177 (N_2177,N_1971,N_1826);
or U2178 (N_2178,N_1808,N_1883);
and U2179 (N_2179,N_1888,N_1833);
or U2180 (N_2180,N_1804,N_1855);
or U2181 (N_2181,N_1875,N_1879);
and U2182 (N_2182,N_1811,N_1960);
and U2183 (N_2183,N_1823,N_1824);
and U2184 (N_2184,N_1917,N_1876);
nor U2185 (N_2185,N_1867,N_1936);
nor U2186 (N_2186,N_1857,N_1953);
xnor U2187 (N_2187,N_1959,N_1900);
xor U2188 (N_2188,N_1977,N_1891);
and U2189 (N_2189,N_1898,N_1839);
or U2190 (N_2190,N_1963,N_1883);
nor U2191 (N_2191,N_1888,N_1847);
xnor U2192 (N_2192,N_1950,N_1845);
xnor U2193 (N_2193,N_1949,N_1859);
and U2194 (N_2194,N_1972,N_1986);
and U2195 (N_2195,N_1808,N_1849);
and U2196 (N_2196,N_1859,N_1848);
or U2197 (N_2197,N_1883,N_1952);
or U2198 (N_2198,N_1833,N_1927);
or U2199 (N_2199,N_1942,N_1924);
and U2200 (N_2200,N_2027,N_2055);
nor U2201 (N_2201,N_2000,N_2140);
or U2202 (N_2202,N_2021,N_2127);
and U2203 (N_2203,N_2115,N_2112);
and U2204 (N_2204,N_2187,N_2105);
and U2205 (N_2205,N_2142,N_2113);
or U2206 (N_2206,N_2195,N_2028);
or U2207 (N_2207,N_2098,N_2147);
nor U2208 (N_2208,N_2198,N_2010);
xnor U2209 (N_2209,N_2188,N_2137);
xnor U2210 (N_2210,N_2051,N_2011);
and U2211 (N_2211,N_2003,N_2166);
or U2212 (N_2212,N_2158,N_2160);
or U2213 (N_2213,N_2154,N_2064);
or U2214 (N_2214,N_2075,N_2190);
nor U2215 (N_2215,N_2136,N_2179);
xor U2216 (N_2216,N_2184,N_2120);
nand U2217 (N_2217,N_2175,N_2036);
nor U2218 (N_2218,N_2052,N_2025);
xnor U2219 (N_2219,N_2099,N_2104);
xor U2220 (N_2220,N_2095,N_2085);
and U2221 (N_2221,N_2086,N_2199);
xnor U2222 (N_2222,N_2012,N_2065);
nand U2223 (N_2223,N_2111,N_2139);
nor U2224 (N_2224,N_2171,N_2096);
nand U2225 (N_2225,N_2033,N_2081);
or U2226 (N_2226,N_2059,N_2002);
and U2227 (N_2227,N_2071,N_2155);
or U2228 (N_2228,N_2173,N_2157);
and U2229 (N_2229,N_2082,N_2102);
nand U2230 (N_2230,N_2063,N_2034);
or U2231 (N_2231,N_2101,N_2076);
nand U2232 (N_2232,N_2056,N_2030);
or U2233 (N_2233,N_2159,N_2193);
or U2234 (N_2234,N_2196,N_2134);
or U2235 (N_2235,N_2191,N_2014);
xnor U2236 (N_2236,N_2167,N_2129);
xor U2237 (N_2237,N_2180,N_2005);
xnor U2238 (N_2238,N_2018,N_2131);
xor U2239 (N_2239,N_2077,N_2066);
xnor U2240 (N_2240,N_2124,N_2149);
nor U2241 (N_2241,N_2169,N_2009);
nand U2242 (N_2242,N_2045,N_2133);
or U2243 (N_2243,N_2126,N_2138);
xor U2244 (N_2244,N_2121,N_2168);
and U2245 (N_2245,N_2119,N_2132);
nor U2246 (N_2246,N_2044,N_2007);
xnor U2247 (N_2247,N_2172,N_2069);
and U2248 (N_2248,N_2143,N_2092);
and U2249 (N_2249,N_2083,N_2162);
and U2250 (N_2250,N_2151,N_2165);
or U2251 (N_2251,N_2079,N_2091);
and U2252 (N_2252,N_2019,N_2023);
and U2253 (N_2253,N_2181,N_2084);
or U2254 (N_2254,N_2185,N_2114);
nand U2255 (N_2255,N_2177,N_2043);
nor U2256 (N_2256,N_2093,N_2148);
or U2257 (N_2257,N_2047,N_2183);
nor U2258 (N_2258,N_2067,N_2072);
or U2259 (N_2259,N_2016,N_2060);
nor U2260 (N_2260,N_2089,N_2110);
xor U2261 (N_2261,N_2130,N_2194);
nor U2262 (N_2262,N_2017,N_2117);
nor U2263 (N_2263,N_2039,N_2057);
nand U2264 (N_2264,N_2118,N_2038);
and U2265 (N_2265,N_2146,N_2073);
xnor U2266 (N_2266,N_2078,N_2058);
nor U2267 (N_2267,N_2061,N_2189);
nor U2268 (N_2268,N_2094,N_2026);
xor U2269 (N_2269,N_2108,N_2037);
or U2270 (N_2270,N_2145,N_2074);
nand U2271 (N_2271,N_2144,N_2049);
and U2272 (N_2272,N_2068,N_2125);
xor U2273 (N_2273,N_2103,N_2106);
and U2274 (N_2274,N_2020,N_2150);
and U2275 (N_2275,N_2176,N_2053);
nor U2276 (N_2276,N_2178,N_2186);
nand U2277 (N_2277,N_2024,N_2192);
nand U2278 (N_2278,N_2090,N_2153);
nand U2279 (N_2279,N_2050,N_2128);
or U2280 (N_2280,N_2161,N_2001);
or U2281 (N_2281,N_2042,N_2046);
xnor U2282 (N_2282,N_2029,N_2097);
or U2283 (N_2283,N_2197,N_2135);
and U2284 (N_2284,N_2032,N_2006);
nand U2285 (N_2285,N_2015,N_2070);
and U2286 (N_2286,N_2088,N_2170);
xor U2287 (N_2287,N_2087,N_2054);
and U2288 (N_2288,N_2163,N_2040);
or U2289 (N_2289,N_2013,N_2062);
and U2290 (N_2290,N_2100,N_2182);
or U2291 (N_2291,N_2109,N_2164);
xnor U2292 (N_2292,N_2048,N_2174);
xor U2293 (N_2293,N_2080,N_2031);
and U2294 (N_2294,N_2008,N_2035);
or U2295 (N_2295,N_2141,N_2004);
xor U2296 (N_2296,N_2116,N_2122);
or U2297 (N_2297,N_2156,N_2123);
nand U2298 (N_2298,N_2022,N_2107);
nor U2299 (N_2299,N_2152,N_2041);
xor U2300 (N_2300,N_2173,N_2011);
or U2301 (N_2301,N_2166,N_2179);
xor U2302 (N_2302,N_2112,N_2061);
nand U2303 (N_2303,N_2084,N_2086);
nand U2304 (N_2304,N_2119,N_2123);
xor U2305 (N_2305,N_2068,N_2001);
or U2306 (N_2306,N_2024,N_2065);
nor U2307 (N_2307,N_2189,N_2117);
and U2308 (N_2308,N_2011,N_2119);
and U2309 (N_2309,N_2188,N_2149);
xnor U2310 (N_2310,N_2019,N_2067);
or U2311 (N_2311,N_2079,N_2177);
or U2312 (N_2312,N_2044,N_2092);
nand U2313 (N_2313,N_2072,N_2087);
and U2314 (N_2314,N_2169,N_2067);
nand U2315 (N_2315,N_2043,N_2151);
xor U2316 (N_2316,N_2148,N_2054);
nor U2317 (N_2317,N_2183,N_2121);
and U2318 (N_2318,N_2109,N_2010);
and U2319 (N_2319,N_2082,N_2004);
or U2320 (N_2320,N_2022,N_2177);
nand U2321 (N_2321,N_2029,N_2135);
and U2322 (N_2322,N_2029,N_2132);
and U2323 (N_2323,N_2080,N_2131);
nand U2324 (N_2324,N_2178,N_2117);
and U2325 (N_2325,N_2023,N_2027);
or U2326 (N_2326,N_2057,N_2157);
and U2327 (N_2327,N_2073,N_2065);
nor U2328 (N_2328,N_2191,N_2083);
xor U2329 (N_2329,N_2161,N_2108);
and U2330 (N_2330,N_2191,N_2163);
and U2331 (N_2331,N_2018,N_2127);
or U2332 (N_2332,N_2149,N_2152);
nand U2333 (N_2333,N_2119,N_2118);
nor U2334 (N_2334,N_2016,N_2125);
xor U2335 (N_2335,N_2085,N_2013);
xor U2336 (N_2336,N_2127,N_2152);
xor U2337 (N_2337,N_2117,N_2095);
and U2338 (N_2338,N_2185,N_2155);
nand U2339 (N_2339,N_2149,N_2020);
xor U2340 (N_2340,N_2081,N_2075);
and U2341 (N_2341,N_2117,N_2074);
or U2342 (N_2342,N_2098,N_2165);
nand U2343 (N_2343,N_2018,N_2029);
nand U2344 (N_2344,N_2054,N_2097);
and U2345 (N_2345,N_2067,N_2111);
and U2346 (N_2346,N_2168,N_2154);
nor U2347 (N_2347,N_2132,N_2075);
or U2348 (N_2348,N_2150,N_2016);
nand U2349 (N_2349,N_2122,N_2081);
xor U2350 (N_2350,N_2118,N_2085);
or U2351 (N_2351,N_2193,N_2030);
nand U2352 (N_2352,N_2156,N_2112);
nand U2353 (N_2353,N_2038,N_2072);
or U2354 (N_2354,N_2116,N_2126);
xnor U2355 (N_2355,N_2013,N_2111);
nand U2356 (N_2356,N_2164,N_2175);
or U2357 (N_2357,N_2112,N_2084);
nand U2358 (N_2358,N_2055,N_2154);
nor U2359 (N_2359,N_2078,N_2101);
nor U2360 (N_2360,N_2126,N_2125);
nand U2361 (N_2361,N_2195,N_2071);
nor U2362 (N_2362,N_2100,N_2185);
or U2363 (N_2363,N_2069,N_2061);
nand U2364 (N_2364,N_2089,N_2159);
xnor U2365 (N_2365,N_2146,N_2055);
nor U2366 (N_2366,N_2146,N_2127);
nand U2367 (N_2367,N_2023,N_2152);
or U2368 (N_2368,N_2023,N_2051);
and U2369 (N_2369,N_2130,N_2090);
nand U2370 (N_2370,N_2154,N_2125);
nor U2371 (N_2371,N_2012,N_2092);
nor U2372 (N_2372,N_2124,N_2062);
and U2373 (N_2373,N_2155,N_2149);
nand U2374 (N_2374,N_2052,N_2079);
xor U2375 (N_2375,N_2141,N_2006);
xor U2376 (N_2376,N_2116,N_2090);
nor U2377 (N_2377,N_2183,N_2130);
or U2378 (N_2378,N_2098,N_2080);
nand U2379 (N_2379,N_2074,N_2154);
and U2380 (N_2380,N_2040,N_2119);
nor U2381 (N_2381,N_2005,N_2132);
nand U2382 (N_2382,N_2107,N_2064);
and U2383 (N_2383,N_2157,N_2011);
xnor U2384 (N_2384,N_2150,N_2132);
or U2385 (N_2385,N_2187,N_2031);
nor U2386 (N_2386,N_2159,N_2023);
nand U2387 (N_2387,N_2027,N_2159);
and U2388 (N_2388,N_2046,N_2060);
or U2389 (N_2389,N_2083,N_2044);
nand U2390 (N_2390,N_2168,N_2129);
xor U2391 (N_2391,N_2006,N_2162);
nor U2392 (N_2392,N_2158,N_2145);
xor U2393 (N_2393,N_2071,N_2187);
nand U2394 (N_2394,N_2038,N_2114);
or U2395 (N_2395,N_2080,N_2060);
nand U2396 (N_2396,N_2057,N_2069);
nand U2397 (N_2397,N_2148,N_2124);
and U2398 (N_2398,N_2080,N_2183);
nor U2399 (N_2399,N_2004,N_2118);
xnor U2400 (N_2400,N_2340,N_2301);
xor U2401 (N_2401,N_2366,N_2385);
nor U2402 (N_2402,N_2376,N_2259);
or U2403 (N_2403,N_2381,N_2369);
xnor U2404 (N_2404,N_2265,N_2322);
xor U2405 (N_2405,N_2383,N_2315);
nand U2406 (N_2406,N_2353,N_2375);
nor U2407 (N_2407,N_2320,N_2226);
nand U2408 (N_2408,N_2219,N_2289);
nand U2409 (N_2409,N_2218,N_2267);
nand U2410 (N_2410,N_2348,N_2329);
or U2411 (N_2411,N_2223,N_2386);
and U2412 (N_2412,N_2208,N_2336);
nor U2413 (N_2413,N_2235,N_2360);
or U2414 (N_2414,N_2324,N_2312);
nand U2415 (N_2415,N_2247,N_2316);
or U2416 (N_2416,N_2397,N_2242);
nor U2417 (N_2417,N_2260,N_2305);
and U2418 (N_2418,N_2206,N_2290);
nor U2419 (N_2419,N_2245,N_2297);
or U2420 (N_2420,N_2335,N_2257);
nor U2421 (N_2421,N_2291,N_2258);
and U2422 (N_2422,N_2362,N_2342);
xnor U2423 (N_2423,N_2238,N_2354);
xor U2424 (N_2424,N_2359,N_2307);
xor U2425 (N_2425,N_2255,N_2205);
nand U2426 (N_2426,N_2358,N_2299);
xor U2427 (N_2427,N_2344,N_2234);
or U2428 (N_2428,N_2326,N_2288);
xnor U2429 (N_2429,N_2328,N_2274);
and U2430 (N_2430,N_2200,N_2241);
or U2431 (N_2431,N_2364,N_2283);
nand U2432 (N_2432,N_2293,N_2311);
xor U2433 (N_2433,N_2231,N_2314);
nor U2434 (N_2434,N_2261,N_2269);
or U2435 (N_2435,N_2252,N_2268);
and U2436 (N_2436,N_2282,N_2204);
xnor U2437 (N_2437,N_2377,N_2285);
nor U2438 (N_2438,N_2248,N_2343);
and U2439 (N_2439,N_2228,N_2334);
or U2440 (N_2440,N_2243,N_2229);
nor U2441 (N_2441,N_2217,N_2306);
nand U2442 (N_2442,N_2286,N_2276);
or U2443 (N_2443,N_2388,N_2302);
nand U2444 (N_2444,N_2230,N_2310);
nand U2445 (N_2445,N_2389,N_2210);
and U2446 (N_2446,N_2263,N_2399);
and U2447 (N_2447,N_2391,N_2361);
nand U2448 (N_2448,N_2321,N_2319);
nor U2449 (N_2449,N_2341,N_2374);
xnor U2450 (N_2450,N_2212,N_2393);
or U2451 (N_2451,N_2330,N_2213);
nor U2452 (N_2452,N_2378,N_2295);
xor U2453 (N_2453,N_2323,N_2363);
nor U2454 (N_2454,N_2251,N_2214);
or U2455 (N_2455,N_2365,N_2201);
nand U2456 (N_2456,N_2250,N_2207);
and U2457 (N_2457,N_2325,N_2209);
nand U2458 (N_2458,N_2271,N_2224);
and U2459 (N_2459,N_2202,N_2294);
nor U2460 (N_2460,N_2318,N_2277);
or U2461 (N_2461,N_2232,N_2327);
or U2462 (N_2462,N_2249,N_2333);
and U2463 (N_2463,N_2313,N_2370);
nor U2464 (N_2464,N_2239,N_2350);
and U2465 (N_2465,N_2211,N_2337);
nor U2466 (N_2466,N_2379,N_2394);
nor U2467 (N_2467,N_2246,N_2253);
and U2468 (N_2468,N_2356,N_2398);
xor U2469 (N_2469,N_2300,N_2352);
nor U2470 (N_2470,N_2256,N_2244);
xor U2471 (N_2471,N_2390,N_2221);
nand U2472 (N_2472,N_2395,N_2220);
or U2473 (N_2473,N_2296,N_2287);
and U2474 (N_2474,N_2346,N_2347);
or U2475 (N_2475,N_2279,N_2372);
xor U2476 (N_2476,N_2236,N_2351);
nand U2477 (N_2477,N_2264,N_2308);
nand U2478 (N_2478,N_2371,N_2281);
nor U2479 (N_2479,N_2222,N_2357);
or U2480 (N_2480,N_2338,N_2225);
xor U2481 (N_2481,N_2396,N_2303);
nand U2482 (N_2482,N_2284,N_2273);
and U2483 (N_2483,N_2233,N_2292);
nand U2484 (N_2484,N_2331,N_2387);
and U2485 (N_2485,N_2237,N_2309);
nand U2486 (N_2486,N_2272,N_2215);
nand U2487 (N_2487,N_2368,N_2203);
nor U2488 (N_2488,N_2339,N_2384);
and U2489 (N_2489,N_2317,N_2240);
and U2490 (N_2490,N_2355,N_2304);
nor U2491 (N_2491,N_2227,N_2367);
or U2492 (N_2492,N_2382,N_2254);
and U2493 (N_2493,N_2216,N_2270);
nand U2494 (N_2494,N_2298,N_2262);
nand U2495 (N_2495,N_2392,N_2380);
nor U2496 (N_2496,N_2280,N_2345);
xor U2497 (N_2497,N_2278,N_2332);
or U2498 (N_2498,N_2373,N_2275);
or U2499 (N_2499,N_2266,N_2349);
and U2500 (N_2500,N_2222,N_2288);
and U2501 (N_2501,N_2351,N_2384);
xnor U2502 (N_2502,N_2277,N_2321);
xnor U2503 (N_2503,N_2301,N_2247);
xor U2504 (N_2504,N_2332,N_2240);
nand U2505 (N_2505,N_2302,N_2381);
nor U2506 (N_2506,N_2244,N_2232);
nor U2507 (N_2507,N_2280,N_2271);
and U2508 (N_2508,N_2338,N_2245);
or U2509 (N_2509,N_2231,N_2210);
or U2510 (N_2510,N_2201,N_2268);
or U2511 (N_2511,N_2385,N_2287);
or U2512 (N_2512,N_2292,N_2287);
or U2513 (N_2513,N_2262,N_2308);
xnor U2514 (N_2514,N_2222,N_2353);
and U2515 (N_2515,N_2348,N_2366);
or U2516 (N_2516,N_2291,N_2234);
nand U2517 (N_2517,N_2390,N_2264);
and U2518 (N_2518,N_2260,N_2258);
or U2519 (N_2519,N_2339,N_2228);
nor U2520 (N_2520,N_2399,N_2371);
nand U2521 (N_2521,N_2305,N_2281);
or U2522 (N_2522,N_2252,N_2278);
or U2523 (N_2523,N_2218,N_2291);
or U2524 (N_2524,N_2267,N_2370);
nand U2525 (N_2525,N_2339,N_2348);
and U2526 (N_2526,N_2343,N_2385);
nor U2527 (N_2527,N_2237,N_2331);
nand U2528 (N_2528,N_2346,N_2324);
nor U2529 (N_2529,N_2331,N_2262);
xnor U2530 (N_2530,N_2338,N_2312);
nand U2531 (N_2531,N_2394,N_2213);
nand U2532 (N_2532,N_2359,N_2383);
and U2533 (N_2533,N_2286,N_2265);
or U2534 (N_2534,N_2317,N_2336);
or U2535 (N_2535,N_2257,N_2238);
xnor U2536 (N_2536,N_2357,N_2359);
or U2537 (N_2537,N_2340,N_2286);
nand U2538 (N_2538,N_2251,N_2369);
or U2539 (N_2539,N_2301,N_2217);
nor U2540 (N_2540,N_2331,N_2240);
and U2541 (N_2541,N_2272,N_2267);
and U2542 (N_2542,N_2321,N_2256);
nand U2543 (N_2543,N_2206,N_2331);
nor U2544 (N_2544,N_2331,N_2261);
nor U2545 (N_2545,N_2250,N_2213);
xor U2546 (N_2546,N_2251,N_2348);
or U2547 (N_2547,N_2334,N_2380);
and U2548 (N_2548,N_2215,N_2228);
or U2549 (N_2549,N_2203,N_2399);
and U2550 (N_2550,N_2365,N_2217);
nor U2551 (N_2551,N_2294,N_2299);
or U2552 (N_2552,N_2371,N_2283);
and U2553 (N_2553,N_2335,N_2321);
nor U2554 (N_2554,N_2381,N_2334);
nand U2555 (N_2555,N_2392,N_2236);
or U2556 (N_2556,N_2331,N_2388);
xor U2557 (N_2557,N_2256,N_2249);
or U2558 (N_2558,N_2220,N_2240);
nor U2559 (N_2559,N_2268,N_2205);
xnor U2560 (N_2560,N_2292,N_2346);
xnor U2561 (N_2561,N_2265,N_2319);
nand U2562 (N_2562,N_2376,N_2202);
nand U2563 (N_2563,N_2297,N_2294);
nor U2564 (N_2564,N_2353,N_2384);
nor U2565 (N_2565,N_2297,N_2342);
and U2566 (N_2566,N_2329,N_2369);
or U2567 (N_2567,N_2256,N_2217);
or U2568 (N_2568,N_2375,N_2274);
or U2569 (N_2569,N_2287,N_2283);
nand U2570 (N_2570,N_2376,N_2393);
or U2571 (N_2571,N_2222,N_2243);
and U2572 (N_2572,N_2382,N_2256);
nand U2573 (N_2573,N_2352,N_2244);
and U2574 (N_2574,N_2261,N_2359);
or U2575 (N_2575,N_2341,N_2336);
nand U2576 (N_2576,N_2340,N_2245);
nor U2577 (N_2577,N_2304,N_2204);
xor U2578 (N_2578,N_2337,N_2238);
and U2579 (N_2579,N_2246,N_2206);
nor U2580 (N_2580,N_2218,N_2290);
or U2581 (N_2581,N_2236,N_2270);
xor U2582 (N_2582,N_2206,N_2330);
or U2583 (N_2583,N_2274,N_2213);
nand U2584 (N_2584,N_2342,N_2232);
and U2585 (N_2585,N_2242,N_2289);
nor U2586 (N_2586,N_2251,N_2309);
nor U2587 (N_2587,N_2303,N_2217);
nor U2588 (N_2588,N_2393,N_2322);
and U2589 (N_2589,N_2376,N_2232);
nor U2590 (N_2590,N_2241,N_2372);
or U2591 (N_2591,N_2326,N_2277);
nand U2592 (N_2592,N_2317,N_2269);
xnor U2593 (N_2593,N_2289,N_2350);
xnor U2594 (N_2594,N_2211,N_2296);
nor U2595 (N_2595,N_2399,N_2219);
xnor U2596 (N_2596,N_2372,N_2323);
nand U2597 (N_2597,N_2243,N_2207);
nor U2598 (N_2598,N_2234,N_2383);
nor U2599 (N_2599,N_2361,N_2375);
nand U2600 (N_2600,N_2407,N_2400);
xor U2601 (N_2601,N_2577,N_2571);
and U2602 (N_2602,N_2490,N_2528);
nand U2603 (N_2603,N_2547,N_2440);
xor U2604 (N_2604,N_2414,N_2521);
or U2605 (N_2605,N_2546,N_2574);
nand U2606 (N_2606,N_2413,N_2494);
or U2607 (N_2607,N_2420,N_2512);
and U2608 (N_2608,N_2444,N_2581);
nor U2609 (N_2609,N_2438,N_2520);
nand U2610 (N_2610,N_2415,N_2426);
nor U2611 (N_2611,N_2524,N_2543);
and U2612 (N_2612,N_2431,N_2466);
xor U2613 (N_2613,N_2507,N_2575);
or U2614 (N_2614,N_2578,N_2503);
nor U2615 (N_2615,N_2569,N_2510);
nand U2616 (N_2616,N_2452,N_2540);
or U2617 (N_2617,N_2573,N_2504);
nand U2618 (N_2618,N_2559,N_2437);
nor U2619 (N_2619,N_2454,N_2427);
xnor U2620 (N_2620,N_2481,N_2486);
xnor U2621 (N_2621,N_2410,N_2537);
and U2622 (N_2622,N_2594,N_2498);
and U2623 (N_2623,N_2457,N_2473);
nand U2624 (N_2624,N_2424,N_2471);
xor U2625 (N_2625,N_2565,N_2549);
and U2626 (N_2626,N_2472,N_2553);
and U2627 (N_2627,N_2517,N_2497);
xnor U2628 (N_2628,N_2552,N_2582);
xor U2629 (N_2629,N_2429,N_2448);
nor U2630 (N_2630,N_2408,N_2422);
nor U2631 (N_2631,N_2491,N_2511);
and U2632 (N_2632,N_2596,N_2580);
nand U2633 (N_2633,N_2576,N_2525);
nor U2634 (N_2634,N_2423,N_2434);
and U2635 (N_2635,N_2545,N_2566);
nand U2636 (N_2636,N_2502,N_2519);
and U2637 (N_2637,N_2514,N_2475);
xor U2638 (N_2638,N_2539,N_2458);
or U2639 (N_2639,N_2428,N_2450);
or U2640 (N_2640,N_2592,N_2522);
or U2641 (N_2641,N_2593,N_2595);
nand U2642 (N_2642,N_2402,N_2432);
and U2643 (N_2643,N_2585,N_2561);
nand U2644 (N_2644,N_2599,N_2579);
and U2645 (N_2645,N_2459,N_2401);
and U2646 (N_2646,N_2462,N_2598);
nor U2647 (N_2647,N_2456,N_2455);
or U2648 (N_2648,N_2554,N_2405);
or U2649 (N_2649,N_2416,N_2530);
or U2650 (N_2650,N_2412,N_2597);
and U2651 (N_2651,N_2474,N_2442);
or U2652 (N_2652,N_2584,N_2469);
nand U2653 (N_2653,N_2556,N_2590);
nand U2654 (N_2654,N_2463,N_2526);
nand U2655 (N_2655,N_2588,N_2446);
nor U2656 (N_2656,N_2451,N_2447);
and U2657 (N_2657,N_2435,N_2499);
nor U2658 (N_2658,N_2419,N_2403);
nand U2659 (N_2659,N_2433,N_2557);
or U2660 (N_2660,N_2587,N_2468);
and U2661 (N_2661,N_2548,N_2411);
or U2662 (N_2662,N_2449,N_2550);
nand U2663 (N_2663,N_2404,N_2476);
and U2664 (N_2664,N_2453,N_2441);
and U2665 (N_2665,N_2505,N_2445);
or U2666 (N_2666,N_2436,N_2562);
and U2667 (N_2667,N_2464,N_2478);
xnor U2668 (N_2668,N_2479,N_2538);
and U2669 (N_2669,N_2509,N_2583);
or U2670 (N_2670,N_2513,N_2586);
or U2671 (N_2671,N_2515,N_2564);
or U2672 (N_2672,N_2488,N_2443);
xnor U2673 (N_2673,N_2572,N_2558);
nor U2674 (N_2674,N_2551,N_2482);
or U2675 (N_2675,N_2532,N_2487);
or U2676 (N_2676,N_2496,N_2555);
nor U2677 (N_2677,N_2535,N_2567);
nand U2678 (N_2678,N_2500,N_2421);
nand U2679 (N_2679,N_2529,N_2493);
nor U2680 (N_2680,N_2568,N_2589);
nor U2681 (N_2681,N_2465,N_2508);
nand U2682 (N_2682,N_2495,N_2541);
nand U2683 (N_2683,N_2470,N_2536);
or U2684 (N_2684,N_2523,N_2544);
nor U2685 (N_2685,N_2489,N_2477);
and U2686 (N_2686,N_2461,N_2485);
or U2687 (N_2687,N_2430,N_2563);
and U2688 (N_2688,N_2516,N_2460);
nor U2689 (N_2689,N_2467,N_2501);
and U2690 (N_2690,N_2518,N_2533);
nor U2691 (N_2691,N_2591,N_2534);
and U2692 (N_2692,N_2480,N_2439);
nand U2693 (N_2693,N_2506,N_2570);
nand U2694 (N_2694,N_2409,N_2492);
nor U2695 (N_2695,N_2527,N_2483);
and U2696 (N_2696,N_2417,N_2531);
and U2697 (N_2697,N_2425,N_2560);
xor U2698 (N_2698,N_2418,N_2484);
and U2699 (N_2699,N_2406,N_2542);
xnor U2700 (N_2700,N_2587,N_2502);
or U2701 (N_2701,N_2525,N_2511);
or U2702 (N_2702,N_2485,N_2489);
xnor U2703 (N_2703,N_2463,N_2584);
or U2704 (N_2704,N_2428,N_2434);
nand U2705 (N_2705,N_2559,N_2497);
and U2706 (N_2706,N_2497,N_2594);
and U2707 (N_2707,N_2548,N_2466);
nand U2708 (N_2708,N_2517,N_2576);
nor U2709 (N_2709,N_2429,N_2414);
nor U2710 (N_2710,N_2453,N_2588);
and U2711 (N_2711,N_2412,N_2573);
and U2712 (N_2712,N_2426,N_2555);
nand U2713 (N_2713,N_2584,N_2458);
or U2714 (N_2714,N_2541,N_2589);
xor U2715 (N_2715,N_2521,N_2598);
and U2716 (N_2716,N_2522,N_2544);
xnor U2717 (N_2717,N_2566,N_2406);
or U2718 (N_2718,N_2466,N_2452);
or U2719 (N_2719,N_2424,N_2457);
nor U2720 (N_2720,N_2411,N_2434);
or U2721 (N_2721,N_2484,N_2470);
nand U2722 (N_2722,N_2476,N_2571);
xor U2723 (N_2723,N_2466,N_2520);
nand U2724 (N_2724,N_2550,N_2412);
or U2725 (N_2725,N_2539,N_2443);
nand U2726 (N_2726,N_2564,N_2474);
nand U2727 (N_2727,N_2460,N_2589);
nor U2728 (N_2728,N_2479,N_2559);
nor U2729 (N_2729,N_2454,N_2585);
nor U2730 (N_2730,N_2474,N_2596);
xnor U2731 (N_2731,N_2573,N_2424);
xor U2732 (N_2732,N_2567,N_2508);
xnor U2733 (N_2733,N_2491,N_2484);
or U2734 (N_2734,N_2420,N_2407);
nand U2735 (N_2735,N_2499,N_2427);
nor U2736 (N_2736,N_2585,N_2438);
and U2737 (N_2737,N_2565,N_2486);
nand U2738 (N_2738,N_2465,N_2469);
xnor U2739 (N_2739,N_2569,N_2492);
nand U2740 (N_2740,N_2431,N_2437);
xnor U2741 (N_2741,N_2474,N_2404);
nor U2742 (N_2742,N_2493,N_2426);
nand U2743 (N_2743,N_2480,N_2579);
xnor U2744 (N_2744,N_2493,N_2540);
nor U2745 (N_2745,N_2402,N_2487);
nand U2746 (N_2746,N_2415,N_2560);
nor U2747 (N_2747,N_2584,N_2512);
xor U2748 (N_2748,N_2588,N_2587);
nand U2749 (N_2749,N_2585,N_2555);
and U2750 (N_2750,N_2511,N_2485);
nand U2751 (N_2751,N_2425,N_2476);
nand U2752 (N_2752,N_2437,N_2408);
nand U2753 (N_2753,N_2417,N_2420);
nor U2754 (N_2754,N_2444,N_2519);
xor U2755 (N_2755,N_2465,N_2586);
and U2756 (N_2756,N_2582,N_2556);
nor U2757 (N_2757,N_2589,N_2432);
nor U2758 (N_2758,N_2432,N_2439);
and U2759 (N_2759,N_2519,N_2476);
xnor U2760 (N_2760,N_2588,N_2570);
nor U2761 (N_2761,N_2466,N_2459);
nand U2762 (N_2762,N_2443,N_2563);
nor U2763 (N_2763,N_2419,N_2451);
or U2764 (N_2764,N_2525,N_2474);
and U2765 (N_2765,N_2512,N_2553);
nor U2766 (N_2766,N_2477,N_2546);
nand U2767 (N_2767,N_2477,N_2418);
or U2768 (N_2768,N_2431,N_2485);
and U2769 (N_2769,N_2561,N_2472);
nor U2770 (N_2770,N_2430,N_2474);
and U2771 (N_2771,N_2498,N_2452);
nor U2772 (N_2772,N_2475,N_2463);
or U2773 (N_2773,N_2406,N_2568);
xnor U2774 (N_2774,N_2530,N_2492);
or U2775 (N_2775,N_2587,N_2583);
and U2776 (N_2776,N_2423,N_2522);
or U2777 (N_2777,N_2534,N_2410);
nor U2778 (N_2778,N_2446,N_2456);
or U2779 (N_2779,N_2574,N_2598);
nor U2780 (N_2780,N_2484,N_2415);
xnor U2781 (N_2781,N_2475,N_2562);
and U2782 (N_2782,N_2402,N_2598);
xnor U2783 (N_2783,N_2451,N_2506);
nor U2784 (N_2784,N_2595,N_2504);
xnor U2785 (N_2785,N_2525,N_2509);
xor U2786 (N_2786,N_2562,N_2437);
or U2787 (N_2787,N_2426,N_2432);
nor U2788 (N_2788,N_2502,N_2579);
nand U2789 (N_2789,N_2508,N_2495);
nor U2790 (N_2790,N_2433,N_2439);
and U2791 (N_2791,N_2509,N_2529);
nand U2792 (N_2792,N_2599,N_2418);
nand U2793 (N_2793,N_2574,N_2480);
nand U2794 (N_2794,N_2587,N_2530);
or U2795 (N_2795,N_2474,N_2457);
nand U2796 (N_2796,N_2461,N_2589);
and U2797 (N_2797,N_2409,N_2557);
and U2798 (N_2798,N_2487,N_2506);
nand U2799 (N_2799,N_2512,N_2543);
nor U2800 (N_2800,N_2781,N_2744);
or U2801 (N_2801,N_2759,N_2635);
xor U2802 (N_2802,N_2717,N_2785);
xnor U2803 (N_2803,N_2794,N_2733);
nand U2804 (N_2804,N_2692,N_2609);
nand U2805 (N_2805,N_2703,N_2767);
xnor U2806 (N_2806,N_2710,N_2667);
xnor U2807 (N_2807,N_2725,N_2658);
nand U2808 (N_2808,N_2693,N_2648);
or U2809 (N_2809,N_2684,N_2790);
nand U2810 (N_2810,N_2752,N_2685);
xnor U2811 (N_2811,N_2629,N_2657);
nor U2812 (N_2812,N_2656,N_2672);
nand U2813 (N_2813,N_2784,N_2668);
nand U2814 (N_2814,N_2610,N_2614);
nand U2815 (N_2815,N_2628,N_2756);
xnor U2816 (N_2816,N_2601,N_2603);
and U2817 (N_2817,N_2731,N_2772);
nor U2818 (N_2818,N_2771,N_2737);
xnor U2819 (N_2819,N_2793,N_2604);
or U2820 (N_2820,N_2741,N_2618);
xor U2821 (N_2821,N_2663,N_2686);
nor U2822 (N_2822,N_2779,N_2679);
nand U2823 (N_2823,N_2704,N_2702);
or U2824 (N_2824,N_2732,N_2798);
xnor U2825 (N_2825,N_2718,N_2766);
or U2826 (N_2826,N_2627,N_2722);
and U2827 (N_2827,N_2606,N_2762);
or U2828 (N_2828,N_2637,N_2757);
and U2829 (N_2829,N_2651,N_2632);
nand U2830 (N_2830,N_2743,N_2600);
nand U2831 (N_2831,N_2792,N_2626);
xnor U2832 (N_2832,N_2716,N_2749);
nand U2833 (N_2833,N_2676,N_2775);
and U2834 (N_2834,N_2763,N_2664);
and U2835 (N_2835,N_2713,N_2639);
xor U2836 (N_2836,N_2611,N_2705);
xnor U2837 (N_2837,N_2788,N_2768);
nand U2838 (N_2838,N_2797,N_2765);
xnor U2839 (N_2839,N_2642,N_2647);
and U2840 (N_2840,N_2706,N_2770);
nor U2841 (N_2841,N_2735,N_2782);
nand U2842 (N_2842,N_2612,N_2755);
or U2843 (N_2843,N_2753,N_2747);
nand U2844 (N_2844,N_2646,N_2750);
or U2845 (N_2845,N_2660,N_2689);
and U2846 (N_2846,N_2746,N_2727);
or U2847 (N_2847,N_2630,N_2720);
and U2848 (N_2848,N_2690,N_2758);
or U2849 (N_2849,N_2649,N_2724);
nand U2850 (N_2850,N_2673,N_2624);
nor U2851 (N_2851,N_2621,N_2777);
or U2852 (N_2852,N_2776,N_2728);
nor U2853 (N_2853,N_2683,N_2674);
nor U2854 (N_2854,N_2653,N_2745);
xor U2855 (N_2855,N_2677,N_2729);
and U2856 (N_2856,N_2734,N_2778);
nand U2857 (N_2857,N_2764,N_2751);
xor U2858 (N_2858,N_2760,N_2738);
nor U2859 (N_2859,N_2709,N_2670);
or U2860 (N_2860,N_2799,N_2698);
and U2861 (N_2861,N_2742,N_2625);
nand U2862 (N_2862,N_2633,N_2696);
and U2863 (N_2863,N_2721,N_2616);
and U2864 (N_2864,N_2620,N_2631);
xor U2865 (N_2865,N_2617,N_2643);
or U2866 (N_2866,N_2619,N_2796);
and U2867 (N_2867,N_2789,N_2708);
or U2868 (N_2868,N_2701,N_2655);
nand U2869 (N_2869,N_2680,N_2682);
nor U2870 (N_2870,N_2661,N_2636);
nand U2871 (N_2871,N_2613,N_2783);
nor U2872 (N_2872,N_2769,N_2666);
xnor U2873 (N_2873,N_2622,N_2650);
and U2874 (N_2874,N_2739,N_2786);
nor U2875 (N_2875,N_2687,N_2714);
nand U2876 (N_2876,N_2723,N_2795);
nand U2877 (N_2877,N_2754,N_2652);
nor U2878 (N_2878,N_2707,N_2699);
nand U2879 (N_2879,N_2736,N_2644);
xor U2880 (N_2880,N_2691,N_2659);
and U2881 (N_2881,N_2761,N_2602);
xor U2882 (N_2882,N_2740,N_2654);
nand U2883 (N_2883,N_2774,N_2748);
nand U2884 (N_2884,N_2662,N_2675);
nand U2885 (N_2885,N_2678,N_2634);
xnor U2886 (N_2886,N_2773,N_2608);
or U2887 (N_2887,N_2711,N_2671);
or U2888 (N_2888,N_2641,N_2780);
and U2889 (N_2889,N_2715,N_2681);
xnor U2890 (N_2890,N_2787,N_2638);
nor U2891 (N_2891,N_2726,N_2669);
xnor U2892 (N_2892,N_2623,N_2688);
and U2893 (N_2893,N_2697,N_2645);
and U2894 (N_2894,N_2730,N_2607);
nor U2895 (N_2895,N_2665,N_2791);
xor U2896 (N_2896,N_2719,N_2615);
nand U2897 (N_2897,N_2700,N_2695);
or U2898 (N_2898,N_2605,N_2640);
or U2899 (N_2899,N_2694,N_2712);
or U2900 (N_2900,N_2767,N_2726);
nand U2901 (N_2901,N_2750,N_2731);
and U2902 (N_2902,N_2612,N_2741);
and U2903 (N_2903,N_2664,N_2722);
nor U2904 (N_2904,N_2780,N_2618);
and U2905 (N_2905,N_2738,N_2661);
nand U2906 (N_2906,N_2734,N_2662);
nand U2907 (N_2907,N_2756,N_2787);
xor U2908 (N_2908,N_2701,N_2735);
and U2909 (N_2909,N_2744,N_2757);
and U2910 (N_2910,N_2757,N_2692);
or U2911 (N_2911,N_2764,N_2739);
and U2912 (N_2912,N_2632,N_2732);
nor U2913 (N_2913,N_2618,N_2610);
nor U2914 (N_2914,N_2772,N_2703);
xor U2915 (N_2915,N_2683,N_2776);
and U2916 (N_2916,N_2624,N_2793);
nor U2917 (N_2917,N_2755,N_2644);
xor U2918 (N_2918,N_2762,N_2798);
and U2919 (N_2919,N_2795,N_2642);
nand U2920 (N_2920,N_2643,N_2640);
nand U2921 (N_2921,N_2672,N_2648);
nand U2922 (N_2922,N_2681,N_2674);
xnor U2923 (N_2923,N_2660,N_2737);
xnor U2924 (N_2924,N_2609,N_2684);
or U2925 (N_2925,N_2661,N_2767);
nor U2926 (N_2926,N_2697,N_2729);
or U2927 (N_2927,N_2675,N_2623);
nand U2928 (N_2928,N_2653,N_2789);
or U2929 (N_2929,N_2656,N_2677);
nor U2930 (N_2930,N_2750,N_2682);
nor U2931 (N_2931,N_2718,N_2773);
nor U2932 (N_2932,N_2665,N_2762);
or U2933 (N_2933,N_2738,N_2755);
or U2934 (N_2934,N_2707,N_2690);
or U2935 (N_2935,N_2774,N_2612);
or U2936 (N_2936,N_2673,N_2797);
xor U2937 (N_2937,N_2795,N_2676);
nor U2938 (N_2938,N_2616,N_2635);
nor U2939 (N_2939,N_2647,N_2702);
nor U2940 (N_2940,N_2783,N_2751);
nand U2941 (N_2941,N_2627,N_2658);
nand U2942 (N_2942,N_2651,N_2679);
or U2943 (N_2943,N_2672,N_2738);
xnor U2944 (N_2944,N_2791,N_2654);
nand U2945 (N_2945,N_2788,N_2628);
and U2946 (N_2946,N_2604,N_2693);
or U2947 (N_2947,N_2690,N_2656);
nor U2948 (N_2948,N_2624,N_2759);
nand U2949 (N_2949,N_2626,N_2715);
xor U2950 (N_2950,N_2741,N_2608);
nor U2951 (N_2951,N_2643,N_2742);
or U2952 (N_2952,N_2718,N_2735);
and U2953 (N_2953,N_2692,N_2707);
nand U2954 (N_2954,N_2778,N_2671);
nand U2955 (N_2955,N_2686,N_2602);
and U2956 (N_2956,N_2677,N_2794);
or U2957 (N_2957,N_2726,N_2769);
xnor U2958 (N_2958,N_2747,N_2756);
and U2959 (N_2959,N_2626,N_2748);
nor U2960 (N_2960,N_2623,N_2691);
xnor U2961 (N_2961,N_2742,N_2603);
nand U2962 (N_2962,N_2626,N_2775);
or U2963 (N_2963,N_2701,N_2659);
xor U2964 (N_2964,N_2692,N_2773);
xor U2965 (N_2965,N_2736,N_2647);
and U2966 (N_2966,N_2694,N_2648);
xnor U2967 (N_2967,N_2761,N_2775);
xnor U2968 (N_2968,N_2605,N_2663);
xor U2969 (N_2969,N_2753,N_2645);
or U2970 (N_2970,N_2642,N_2702);
or U2971 (N_2971,N_2753,N_2705);
and U2972 (N_2972,N_2736,N_2789);
nor U2973 (N_2973,N_2673,N_2738);
nand U2974 (N_2974,N_2617,N_2713);
nand U2975 (N_2975,N_2692,N_2620);
xor U2976 (N_2976,N_2629,N_2745);
or U2977 (N_2977,N_2676,N_2778);
xnor U2978 (N_2978,N_2743,N_2721);
xnor U2979 (N_2979,N_2616,N_2626);
nor U2980 (N_2980,N_2679,N_2666);
or U2981 (N_2981,N_2787,N_2758);
xor U2982 (N_2982,N_2760,N_2741);
and U2983 (N_2983,N_2767,N_2722);
nand U2984 (N_2984,N_2653,N_2797);
or U2985 (N_2985,N_2682,N_2601);
nand U2986 (N_2986,N_2625,N_2728);
nand U2987 (N_2987,N_2729,N_2756);
nor U2988 (N_2988,N_2709,N_2639);
or U2989 (N_2989,N_2711,N_2762);
nand U2990 (N_2990,N_2715,N_2656);
and U2991 (N_2991,N_2687,N_2632);
or U2992 (N_2992,N_2779,N_2743);
or U2993 (N_2993,N_2762,N_2658);
nand U2994 (N_2994,N_2680,N_2743);
xnor U2995 (N_2995,N_2667,N_2726);
nand U2996 (N_2996,N_2761,N_2610);
and U2997 (N_2997,N_2688,N_2772);
xor U2998 (N_2998,N_2761,N_2675);
nor U2999 (N_2999,N_2737,N_2744);
xor U3000 (N_3000,N_2965,N_2992);
nand U3001 (N_3001,N_2912,N_2820);
xor U3002 (N_3002,N_2808,N_2875);
nor U3003 (N_3003,N_2938,N_2861);
nand U3004 (N_3004,N_2930,N_2852);
nor U3005 (N_3005,N_2903,N_2975);
or U3006 (N_3006,N_2893,N_2884);
or U3007 (N_3007,N_2879,N_2942);
nor U3008 (N_3008,N_2946,N_2896);
xnor U3009 (N_3009,N_2842,N_2918);
or U3010 (N_3010,N_2866,N_2881);
nand U3011 (N_3011,N_2859,N_2906);
or U3012 (N_3012,N_2983,N_2821);
and U3013 (N_3013,N_2892,N_2956);
xor U3014 (N_3014,N_2828,N_2978);
nor U3015 (N_3015,N_2940,N_2995);
or U3016 (N_3016,N_2891,N_2888);
nor U3017 (N_3017,N_2923,N_2972);
nor U3018 (N_3018,N_2890,N_2927);
nor U3019 (N_3019,N_2911,N_2813);
and U3020 (N_3020,N_2981,N_2921);
and U3021 (N_3021,N_2837,N_2849);
nor U3022 (N_3022,N_2967,N_2948);
and U3023 (N_3023,N_2908,N_2999);
xor U3024 (N_3024,N_2936,N_2864);
nand U3025 (N_3025,N_2984,N_2959);
or U3026 (N_3026,N_2939,N_2979);
or U3027 (N_3027,N_2865,N_2924);
nand U3028 (N_3028,N_2922,N_2913);
or U3029 (N_3029,N_2834,N_2819);
nor U3030 (N_3030,N_2832,N_2800);
nand U3031 (N_3031,N_2883,N_2878);
nor U3032 (N_3032,N_2846,N_2873);
nor U3033 (N_3033,N_2909,N_2931);
nand U3034 (N_3034,N_2805,N_2966);
xnor U3035 (N_3035,N_2961,N_2947);
nor U3036 (N_3036,N_2886,N_2987);
nand U3037 (N_3037,N_2860,N_2920);
or U3038 (N_3038,N_2841,N_2843);
nor U3039 (N_3039,N_2985,N_2885);
xor U3040 (N_3040,N_2815,N_2840);
nor U3041 (N_3041,N_2960,N_2933);
or U3042 (N_3042,N_2934,N_2835);
and U3043 (N_3043,N_2848,N_2863);
and U3044 (N_3044,N_2929,N_2900);
xor U3045 (N_3045,N_2845,N_2824);
or U3046 (N_3046,N_2818,N_2963);
and U3047 (N_3047,N_2889,N_2910);
or U3048 (N_3048,N_2833,N_2806);
xor U3049 (N_3049,N_2973,N_2952);
xnor U3050 (N_3050,N_2809,N_2974);
nand U3051 (N_3051,N_2954,N_2964);
xor U3052 (N_3052,N_2998,N_2919);
or U3053 (N_3053,N_2810,N_2976);
or U3054 (N_3054,N_2950,N_2914);
or U3055 (N_3055,N_2851,N_2994);
and U3056 (N_3056,N_2953,N_2988);
xnor U3057 (N_3057,N_2989,N_2844);
and U3058 (N_3058,N_2904,N_2867);
or U3059 (N_3059,N_2836,N_2801);
nor U3060 (N_3060,N_2907,N_2858);
nor U3061 (N_3061,N_2802,N_2944);
and U3062 (N_3062,N_2857,N_2894);
xor U3063 (N_3063,N_2982,N_2814);
nor U3064 (N_3064,N_2868,N_2968);
nor U3065 (N_3065,N_2869,N_2877);
or U3066 (N_3066,N_2986,N_2807);
xor U3067 (N_3067,N_2870,N_2977);
nor U3068 (N_3068,N_2917,N_2941);
and U3069 (N_3069,N_2997,N_2839);
or U3070 (N_3070,N_2943,N_2902);
or U3071 (N_3071,N_2958,N_2928);
nand U3072 (N_3072,N_2826,N_2897);
nand U3073 (N_3073,N_2895,N_2955);
nand U3074 (N_3074,N_2935,N_2816);
and U3075 (N_3075,N_2887,N_2949);
nor U3076 (N_3076,N_2853,N_2970);
and U3077 (N_3077,N_2830,N_2990);
nor U3078 (N_3078,N_2822,N_2825);
and U3079 (N_3079,N_2829,N_2969);
nor U3080 (N_3080,N_2937,N_2991);
and U3081 (N_3081,N_2957,N_2962);
and U3082 (N_3082,N_2862,N_2803);
or U3083 (N_3083,N_2827,N_2831);
xor U3084 (N_3084,N_2925,N_2838);
xnor U3085 (N_3085,N_2916,N_2898);
nand U3086 (N_3086,N_2915,N_2847);
nor U3087 (N_3087,N_2804,N_2817);
and U3088 (N_3088,N_2876,N_2872);
and U3089 (N_3089,N_2850,N_2971);
nand U3090 (N_3090,N_2812,N_2899);
and U3091 (N_3091,N_2811,N_2926);
and U3092 (N_3092,N_2880,N_2980);
or U3093 (N_3093,N_2855,N_2932);
nand U3094 (N_3094,N_2882,N_2905);
and U3095 (N_3095,N_2945,N_2871);
or U3096 (N_3096,N_2856,N_2854);
nand U3097 (N_3097,N_2951,N_2901);
nor U3098 (N_3098,N_2874,N_2993);
and U3099 (N_3099,N_2823,N_2996);
xor U3100 (N_3100,N_2856,N_2995);
and U3101 (N_3101,N_2863,N_2969);
xnor U3102 (N_3102,N_2990,N_2806);
nand U3103 (N_3103,N_2819,N_2802);
or U3104 (N_3104,N_2871,N_2902);
or U3105 (N_3105,N_2866,N_2890);
or U3106 (N_3106,N_2820,N_2879);
or U3107 (N_3107,N_2864,N_2813);
nor U3108 (N_3108,N_2996,N_2879);
or U3109 (N_3109,N_2826,N_2951);
and U3110 (N_3110,N_2871,N_2915);
xnor U3111 (N_3111,N_2988,N_2868);
nand U3112 (N_3112,N_2933,N_2864);
nand U3113 (N_3113,N_2989,N_2817);
nand U3114 (N_3114,N_2936,N_2932);
nand U3115 (N_3115,N_2854,N_2877);
and U3116 (N_3116,N_2975,N_2880);
xnor U3117 (N_3117,N_2820,N_2837);
xor U3118 (N_3118,N_2986,N_2825);
or U3119 (N_3119,N_2909,N_2955);
or U3120 (N_3120,N_2967,N_2849);
xnor U3121 (N_3121,N_2999,N_2951);
nor U3122 (N_3122,N_2918,N_2957);
and U3123 (N_3123,N_2926,N_2915);
or U3124 (N_3124,N_2949,N_2987);
nand U3125 (N_3125,N_2845,N_2833);
xnor U3126 (N_3126,N_2915,N_2909);
xnor U3127 (N_3127,N_2919,N_2934);
nor U3128 (N_3128,N_2820,N_2934);
nand U3129 (N_3129,N_2990,N_2941);
or U3130 (N_3130,N_2901,N_2859);
xnor U3131 (N_3131,N_2802,N_2865);
or U3132 (N_3132,N_2802,N_2982);
nand U3133 (N_3133,N_2828,N_2937);
nor U3134 (N_3134,N_2896,N_2900);
or U3135 (N_3135,N_2904,N_2921);
and U3136 (N_3136,N_2957,N_2806);
xnor U3137 (N_3137,N_2865,N_2912);
or U3138 (N_3138,N_2937,N_2806);
xor U3139 (N_3139,N_2841,N_2814);
nor U3140 (N_3140,N_2847,N_2906);
xor U3141 (N_3141,N_2969,N_2849);
and U3142 (N_3142,N_2859,N_2858);
and U3143 (N_3143,N_2905,N_2844);
or U3144 (N_3144,N_2925,N_2928);
or U3145 (N_3145,N_2801,N_2864);
or U3146 (N_3146,N_2909,N_2986);
and U3147 (N_3147,N_2846,N_2893);
nor U3148 (N_3148,N_2880,N_2985);
and U3149 (N_3149,N_2930,N_2990);
nand U3150 (N_3150,N_2858,N_2990);
nand U3151 (N_3151,N_2959,N_2906);
xor U3152 (N_3152,N_2951,N_2962);
or U3153 (N_3153,N_2899,N_2848);
xor U3154 (N_3154,N_2954,N_2820);
and U3155 (N_3155,N_2830,N_2836);
or U3156 (N_3156,N_2847,N_2800);
nor U3157 (N_3157,N_2832,N_2833);
and U3158 (N_3158,N_2879,N_2912);
nor U3159 (N_3159,N_2936,N_2912);
nor U3160 (N_3160,N_2823,N_2829);
and U3161 (N_3161,N_2829,N_2987);
xnor U3162 (N_3162,N_2900,N_2970);
and U3163 (N_3163,N_2848,N_2963);
or U3164 (N_3164,N_2845,N_2829);
and U3165 (N_3165,N_2861,N_2863);
nor U3166 (N_3166,N_2865,N_2900);
xor U3167 (N_3167,N_2901,N_2935);
and U3168 (N_3168,N_2954,N_2975);
xor U3169 (N_3169,N_2818,N_2995);
and U3170 (N_3170,N_2874,N_2933);
xnor U3171 (N_3171,N_2951,N_2875);
and U3172 (N_3172,N_2832,N_2825);
or U3173 (N_3173,N_2986,N_2927);
or U3174 (N_3174,N_2975,N_2864);
nand U3175 (N_3175,N_2875,N_2824);
or U3176 (N_3176,N_2942,N_2985);
or U3177 (N_3177,N_2950,N_2926);
and U3178 (N_3178,N_2947,N_2946);
and U3179 (N_3179,N_2918,N_2863);
nor U3180 (N_3180,N_2862,N_2910);
nand U3181 (N_3181,N_2949,N_2842);
or U3182 (N_3182,N_2940,N_2966);
or U3183 (N_3183,N_2958,N_2805);
nand U3184 (N_3184,N_2985,N_2939);
and U3185 (N_3185,N_2865,N_2962);
or U3186 (N_3186,N_2864,N_2850);
xor U3187 (N_3187,N_2988,N_2911);
nand U3188 (N_3188,N_2906,N_2948);
and U3189 (N_3189,N_2876,N_2847);
and U3190 (N_3190,N_2994,N_2990);
nor U3191 (N_3191,N_2861,N_2932);
xnor U3192 (N_3192,N_2903,N_2865);
nand U3193 (N_3193,N_2996,N_2915);
nor U3194 (N_3194,N_2896,N_2813);
or U3195 (N_3195,N_2858,N_2893);
nor U3196 (N_3196,N_2821,N_2851);
and U3197 (N_3197,N_2807,N_2853);
and U3198 (N_3198,N_2984,N_2830);
or U3199 (N_3199,N_2810,N_2892);
nor U3200 (N_3200,N_3107,N_3123);
and U3201 (N_3201,N_3140,N_3159);
nand U3202 (N_3202,N_3092,N_3065);
nor U3203 (N_3203,N_3091,N_3181);
nor U3204 (N_3204,N_3147,N_3194);
or U3205 (N_3205,N_3075,N_3099);
or U3206 (N_3206,N_3130,N_3030);
xor U3207 (N_3207,N_3115,N_3139);
xor U3208 (N_3208,N_3137,N_3150);
nor U3209 (N_3209,N_3010,N_3083);
nor U3210 (N_3210,N_3097,N_3000);
and U3211 (N_3211,N_3031,N_3160);
nand U3212 (N_3212,N_3105,N_3015);
or U3213 (N_3213,N_3164,N_3165);
or U3214 (N_3214,N_3157,N_3153);
or U3215 (N_3215,N_3032,N_3122);
xor U3216 (N_3216,N_3043,N_3119);
or U3217 (N_3217,N_3005,N_3182);
and U3218 (N_3218,N_3067,N_3021);
xnor U3219 (N_3219,N_3076,N_3135);
and U3220 (N_3220,N_3085,N_3132);
nand U3221 (N_3221,N_3176,N_3024);
xnor U3222 (N_3222,N_3114,N_3184);
or U3223 (N_3223,N_3109,N_3002);
xnor U3224 (N_3224,N_3025,N_3033);
nor U3225 (N_3225,N_3127,N_3061);
and U3226 (N_3226,N_3170,N_3174);
and U3227 (N_3227,N_3177,N_3156);
or U3228 (N_3228,N_3047,N_3138);
and U3229 (N_3229,N_3073,N_3198);
xor U3230 (N_3230,N_3003,N_3191);
or U3231 (N_3231,N_3103,N_3192);
or U3232 (N_3232,N_3056,N_3133);
nor U3233 (N_3233,N_3087,N_3069);
nor U3234 (N_3234,N_3155,N_3095);
nand U3235 (N_3235,N_3086,N_3016);
nand U3236 (N_3236,N_3058,N_3066);
nor U3237 (N_3237,N_3178,N_3173);
or U3238 (N_3238,N_3151,N_3028);
nand U3239 (N_3239,N_3042,N_3187);
or U3240 (N_3240,N_3126,N_3007);
or U3241 (N_3241,N_3046,N_3027);
nand U3242 (N_3242,N_3082,N_3175);
nand U3243 (N_3243,N_3131,N_3172);
nand U3244 (N_3244,N_3145,N_3041);
nor U3245 (N_3245,N_3018,N_3022);
xor U3246 (N_3246,N_3196,N_3072);
xnor U3247 (N_3247,N_3062,N_3179);
xnor U3248 (N_3248,N_3071,N_3106);
or U3249 (N_3249,N_3189,N_3185);
nand U3250 (N_3250,N_3129,N_3104);
and U3251 (N_3251,N_3112,N_3057);
and U3252 (N_3252,N_3149,N_3144);
nor U3253 (N_3253,N_3134,N_3146);
xnor U3254 (N_3254,N_3152,N_3120);
xor U3255 (N_3255,N_3166,N_3055);
and U3256 (N_3256,N_3044,N_3154);
xnor U3257 (N_3257,N_3118,N_3052);
xor U3258 (N_3258,N_3008,N_3195);
or U3259 (N_3259,N_3020,N_3001);
and U3260 (N_3260,N_3136,N_3169);
nand U3261 (N_3261,N_3110,N_3079);
xnor U3262 (N_3262,N_3078,N_3029);
nor U3263 (N_3263,N_3053,N_3186);
nand U3264 (N_3264,N_3193,N_3050);
nand U3265 (N_3265,N_3012,N_3142);
nor U3266 (N_3266,N_3163,N_3128);
and U3267 (N_3267,N_3006,N_3102);
nor U3268 (N_3268,N_3036,N_3148);
and U3269 (N_3269,N_3038,N_3048);
nor U3270 (N_3270,N_3035,N_3088);
nor U3271 (N_3271,N_3188,N_3100);
and U3272 (N_3272,N_3113,N_3108);
nand U3273 (N_3273,N_3125,N_3049);
nand U3274 (N_3274,N_3098,N_3117);
nand U3275 (N_3275,N_3045,N_3019);
nand U3276 (N_3276,N_3094,N_3060);
xnor U3277 (N_3277,N_3096,N_3011);
nand U3278 (N_3278,N_3059,N_3023);
nand U3279 (N_3279,N_3070,N_3171);
nor U3280 (N_3280,N_3180,N_3014);
or U3281 (N_3281,N_3101,N_3080);
nand U3282 (N_3282,N_3199,N_3013);
nor U3283 (N_3283,N_3081,N_3089);
or U3284 (N_3284,N_3074,N_3161);
nand U3285 (N_3285,N_3143,N_3068);
or U3286 (N_3286,N_3051,N_3063);
nand U3287 (N_3287,N_3039,N_3111);
or U3288 (N_3288,N_3026,N_3116);
xor U3289 (N_3289,N_3158,N_3197);
or U3290 (N_3290,N_3077,N_3090);
nand U3291 (N_3291,N_3162,N_3093);
xnor U3292 (N_3292,N_3183,N_3054);
nor U3293 (N_3293,N_3084,N_3017);
and U3294 (N_3294,N_3190,N_3037);
nor U3295 (N_3295,N_3168,N_3141);
xnor U3296 (N_3296,N_3004,N_3009);
xnor U3297 (N_3297,N_3124,N_3034);
xor U3298 (N_3298,N_3040,N_3167);
nand U3299 (N_3299,N_3064,N_3121);
xor U3300 (N_3300,N_3033,N_3000);
or U3301 (N_3301,N_3197,N_3116);
nor U3302 (N_3302,N_3111,N_3012);
and U3303 (N_3303,N_3090,N_3088);
nor U3304 (N_3304,N_3121,N_3089);
xor U3305 (N_3305,N_3043,N_3125);
or U3306 (N_3306,N_3003,N_3107);
and U3307 (N_3307,N_3041,N_3038);
nor U3308 (N_3308,N_3085,N_3009);
nand U3309 (N_3309,N_3107,N_3127);
or U3310 (N_3310,N_3137,N_3000);
nor U3311 (N_3311,N_3165,N_3143);
xnor U3312 (N_3312,N_3073,N_3182);
nor U3313 (N_3313,N_3189,N_3187);
nor U3314 (N_3314,N_3002,N_3145);
and U3315 (N_3315,N_3030,N_3027);
nand U3316 (N_3316,N_3006,N_3065);
xor U3317 (N_3317,N_3098,N_3088);
xor U3318 (N_3318,N_3008,N_3169);
and U3319 (N_3319,N_3104,N_3001);
and U3320 (N_3320,N_3119,N_3134);
nor U3321 (N_3321,N_3126,N_3085);
xor U3322 (N_3322,N_3169,N_3095);
xor U3323 (N_3323,N_3079,N_3131);
nor U3324 (N_3324,N_3178,N_3183);
and U3325 (N_3325,N_3105,N_3037);
nand U3326 (N_3326,N_3045,N_3126);
nand U3327 (N_3327,N_3176,N_3172);
nor U3328 (N_3328,N_3075,N_3089);
nand U3329 (N_3329,N_3019,N_3005);
xor U3330 (N_3330,N_3084,N_3101);
and U3331 (N_3331,N_3056,N_3188);
xor U3332 (N_3332,N_3174,N_3100);
nor U3333 (N_3333,N_3176,N_3182);
nand U3334 (N_3334,N_3088,N_3158);
nor U3335 (N_3335,N_3172,N_3024);
nor U3336 (N_3336,N_3192,N_3167);
xnor U3337 (N_3337,N_3180,N_3076);
nand U3338 (N_3338,N_3001,N_3058);
nor U3339 (N_3339,N_3150,N_3182);
nor U3340 (N_3340,N_3065,N_3186);
nand U3341 (N_3341,N_3119,N_3158);
and U3342 (N_3342,N_3179,N_3175);
or U3343 (N_3343,N_3072,N_3110);
and U3344 (N_3344,N_3171,N_3062);
xnor U3345 (N_3345,N_3055,N_3025);
nand U3346 (N_3346,N_3125,N_3005);
and U3347 (N_3347,N_3169,N_3051);
and U3348 (N_3348,N_3080,N_3017);
nand U3349 (N_3349,N_3137,N_3058);
nand U3350 (N_3350,N_3075,N_3178);
and U3351 (N_3351,N_3167,N_3034);
nand U3352 (N_3352,N_3082,N_3080);
nor U3353 (N_3353,N_3118,N_3139);
and U3354 (N_3354,N_3117,N_3061);
or U3355 (N_3355,N_3124,N_3138);
and U3356 (N_3356,N_3152,N_3112);
and U3357 (N_3357,N_3125,N_3027);
or U3358 (N_3358,N_3140,N_3094);
or U3359 (N_3359,N_3025,N_3000);
xnor U3360 (N_3360,N_3115,N_3088);
or U3361 (N_3361,N_3135,N_3174);
and U3362 (N_3362,N_3148,N_3143);
xor U3363 (N_3363,N_3007,N_3043);
xnor U3364 (N_3364,N_3064,N_3019);
nor U3365 (N_3365,N_3154,N_3059);
or U3366 (N_3366,N_3038,N_3060);
xor U3367 (N_3367,N_3157,N_3087);
xnor U3368 (N_3368,N_3008,N_3062);
or U3369 (N_3369,N_3192,N_3121);
nor U3370 (N_3370,N_3004,N_3021);
nand U3371 (N_3371,N_3079,N_3068);
or U3372 (N_3372,N_3164,N_3033);
nand U3373 (N_3373,N_3065,N_3098);
nand U3374 (N_3374,N_3105,N_3018);
or U3375 (N_3375,N_3045,N_3018);
xnor U3376 (N_3376,N_3009,N_3012);
or U3377 (N_3377,N_3062,N_3133);
or U3378 (N_3378,N_3146,N_3009);
and U3379 (N_3379,N_3031,N_3070);
or U3380 (N_3380,N_3072,N_3194);
xor U3381 (N_3381,N_3013,N_3190);
nor U3382 (N_3382,N_3032,N_3049);
nor U3383 (N_3383,N_3032,N_3113);
nand U3384 (N_3384,N_3048,N_3155);
xnor U3385 (N_3385,N_3017,N_3075);
and U3386 (N_3386,N_3098,N_3043);
nand U3387 (N_3387,N_3089,N_3021);
nor U3388 (N_3388,N_3149,N_3133);
and U3389 (N_3389,N_3167,N_3179);
or U3390 (N_3390,N_3154,N_3077);
xor U3391 (N_3391,N_3068,N_3185);
xor U3392 (N_3392,N_3130,N_3183);
nand U3393 (N_3393,N_3153,N_3083);
nor U3394 (N_3394,N_3070,N_3040);
or U3395 (N_3395,N_3103,N_3187);
nand U3396 (N_3396,N_3146,N_3086);
nor U3397 (N_3397,N_3082,N_3008);
and U3398 (N_3398,N_3000,N_3117);
xor U3399 (N_3399,N_3118,N_3120);
and U3400 (N_3400,N_3240,N_3299);
nand U3401 (N_3401,N_3265,N_3286);
or U3402 (N_3402,N_3315,N_3354);
nor U3403 (N_3403,N_3264,N_3276);
xor U3404 (N_3404,N_3340,N_3391);
or U3405 (N_3405,N_3289,N_3318);
and U3406 (N_3406,N_3233,N_3210);
and U3407 (N_3407,N_3230,N_3229);
or U3408 (N_3408,N_3360,N_3239);
nor U3409 (N_3409,N_3313,N_3358);
xor U3410 (N_3410,N_3320,N_3303);
xnor U3411 (N_3411,N_3282,N_3242);
xnor U3412 (N_3412,N_3349,N_3385);
or U3413 (N_3413,N_3347,N_3307);
xor U3414 (N_3414,N_3369,N_3367);
and U3415 (N_3415,N_3371,N_3259);
and U3416 (N_3416,N_3281,N_3243);
nor U3417 (N_3417,N_3396,N_3312);
xnor U3418 (N_3418,N_3308,N_3221);
xnor U3419 (N_3419,N_3317,N_3351);
nand U3420 (N_3420,N_3258,N_3208);
nand U3421 (N_3421,N_3332,N_3355);
or U3422 (N_3422,N_3368,N_3342);
xnor U3423 (N_3423,N_3205,N_3272);
nand U3424 (N_3424,N_3370,N_3363);
nand U3425 (N_3425,N_3231,N_3298);
nand U3426 (N_3426,N_3393,N_3302);
xnor U3427 (N_3427,N_3241,N_3321);
nand U3428 (N_3428,N_3237,N_3292);
and U3429 (N_3429,N_3295,N_3341);
xnor U3430 (N_3430,N_3333,N_3225);
xor U3431 (N_3431,N_3365,N_3350);
xor U3432 (N_3432,N_3395,N_3390);
or U3433 (N_3433,N_3375,N_3222);
nand U3434 (N_3434,N_3219,N_3334);
nand U3435 (N_3435,N_3343,N_3212);
nand U3436 (N_3436,N_3253,N_3206);
or U3437 (N_3437,N_3389,N_3274);
xnor U3438 (N_3438,N_3263,N_3373);
and U3439 (N_3439,N_3204,N_3293);
and U3440 (N_3440,N_3257,N_3279);
xnor U3441 (N_3441,N_3394,N_3338);
nand U3442 (N_3442,N_3344,N_3361);
and U3443 (N_3443,N_3203,N_3324);
xnor U3444 (N_3444,N_3245,N_3252);
nor U3445 (N_3445,N_3328,N_3228);
and U3446 (N_3446,N_3238,N_3304);
xnor U3447 (N_3447,N_3356,N_3201);
and U3448 (N_3448,N_3366,N_3346);
or U3449 (N_3449,N_3209,N_3277);
xnor U3450 (N_3450,N_3336,N_3378);
xnor U3451 (N_3451,N_3382,N_3235);
nand U3452 (N_3452,N_3376,N_3251);
nand U3453 (N_3453,N_3256,N_3300);
or U3454 (N_3454,N_3323,N_3284);
and U3455 (N_3455,N_3337,N_3329);
xor U3456 (N_3456,N_3398,N_3290);
xor U3457 (N_3457,N_3246,N_3268);
nand U3458 (N_3458,N_3339,N_3260);
or U3459 (N_3459,N_3244,N_3306);
xor U3460 (N_3460,N_3326,N_3215);
or U3461 (N_3461,N_3269,N_3377);
nor U3462 (N_3462,N_3202,N_3353);
xor U3463 (N_3463,N_3226,N_3275);
or U3464 (N_3464,N_3325,N_3291);
and U3465 (N_3465,N_3374,N_3310);
nor U3466 (N_3466,N_3362,N_3248);
nor U3467 (N_3467,N_3254,N_3359);
or U3468 (N_3468,N_3218,N_3379);
or U3469 (N_3469,N_3236,N_3234);
nor U3470 (N_3470,N_3255,N_3386);
and U3471 (N_3471,N_3262,N_3216);
and U3472 (N_3472,N_3288,N_3267);
nand U3473 (N_3473,N_3392,N_3380);
and U3474 (N_3474,N_3220,N_3348);
xor U3475 (N_3475,N_3283,N_3296);
or U3476 (N_3476,N_3322,N_3270);
nand U3477 (N_3477,N_3247,N_3266);
or U3478 (N_3478,N_3319,N_3227);
or U3479 (N_3479,N_3327,N_3335);
xnor U3480 (N_3480,N_3214,N_3381);
nor U3481 (N_3481,N_3285,N_3217);
nor U3482 (N_3482,N_3345,N_3287);
and U3483 (N_3483,N_3211,N_3357);
nor U3484 (N_3484,N_3261,N_3311);
xor U3485 (N_3485,N_3372,N_3399);
nand U3486 (N_3486,N_3309,N_3232);
nand U3487 (N_3487,N_3305,N_3314);
xor U3488 (N_3488,N_3388,N_3223);
and U3489 (N_3489,N_3280,N_3250);
nand U3490 (N_3490,N_3364,N_3200);
xnor U3491 (N_3491,N_3397,N_3331);
or U3492 (N_3492,N_3249,N_3301);
nor U3493 (N_3493,N_3316,N_3387);
or U3494 (N_3494,N_3273,N_3271);
nand U3495 (N_3495,N_3330,N_3278);
or U3496 (N_3496,N_3383,N_3207);
or U3497 (N_3497,N_3294,N_3352);
xor U3498 (N_3498,N_3384,N_3213);
nand U3499 (N_3499,N_3224,N_3297);
nand U3500 (N_3500,N_3267,N_3285);
and U3501 (N_3501,N_3232,N_3246);
nand U3502 (N_3502,N_3353,N_3374);
xnor U3503 (N_3503,N_3230,N_3220);
xnor U3504 (N_3504,N_3301,N_3291);
and U3505 (N_3505,N_3278,N_3266);
and U3506 (N_3506,N_3245,N_3282);
xnor U3507 (N_3507,N_3274,N_3342);
nor U3508 (N_3508,N_3218,N_3348);
nor U3509 (N_3509,N_3312,N_3286);
nand U3510 (N_3510,N_3272,N_3368);
or U3511 (N_3511,N_3330,N_3218);
nand U3512 (N_3512,N_3330,N_3348);
and U3513 (N_3513,N_3338,N_3254);
nor U3514 (N_3514,N_3304,N_3201);
and U3515 (N_3515,N_3233,N_3379);
and U3516 (N_3516,N_3267,N_3271);
and U3517 (N_3517,N_3330,N_3283);
nor U3518 (N_3518,N_3340,N_3310);
or U3519 (N_3519,N_3346,N_3308);
xnor U3520 (N_3520,N_3237,N_3248);
or U3521 (N_3521,N_3261,N_3371);
and U3522 (N_3522,N_3326,N_3221);
and U3523 (N_3523,N_3260,N_3383);
or U3524 (N_3524,N_3248,N_3340);
nand U3525 (N_3525,N_3346,N_3229);
and U3526 (N_3526,N_3388,N_3372);
xnor U3527 (N_3527,N_3243,N_3231);
nand U3528 (N_3528,N_3358,N_3253);
and U3529 (N_3529,N_3353,N_3287);
xor U3530 (N_3530,N_3263,N_3395);
nand U3531 (N_3531,N_3303,N_3332);
nor U3532 (N_3532,N_3244,N_3380);
and U3533 (N_3533,N_3364,N_3395);
or U3534 (N_3534,N_3336,N_3352);
nor U3535 (N_3535,N_3367,N_3307);
and U3536 (N_3536,N_3361,N_3268);
and U3537 (N_3537,N_3318,N_3309);
xnor U3538 (N_3538,N_3288,N_3380);
nand U3539 (N_3539,N_3368,N_3392);
nor U3540 (N_3540,N_3243,N_3258);
and U3541 (N_3541,N_3303,N_3233);
nor U3542 (N_3542,N_3346,N_3211);
nor U3543 (N_3543,N_3361,N_3234);
xor U3544 (N_3544,N_3312,N_3373);
nor U3545 (N_3545,N_3238,N_3374);
xnor U3546 (N_3546,N_3206,N_3348);
or U3547 (N_3547,N_3343,N_3353);
xnor U3548 (N_3548,N_3209,N_3257);
xor U3549 (N_3549,N_3266,N_3356);
nand U3550 (N_3550,N_3355,N_3255);
and U3551 (N_3551,N_3399,N_3256);
xnor U3552 (N_3552,N_3275,N_3287);
and U3553 (N_3553,N_3282,N_3338);
and U3554 (N_3554,N_3361,N_3273);
nor U3555 (N_3555,N_3337,N_3398);
nand U3556 (N_3556,N_3386,N_3393);
and U3557 (N_3557,N_3231,N_3301);
and U3558 (N_3558,N_3219,N_3398);
nor U3559 (N_3559,N_3277,N_3203);
nor U3560 (N_3560,N_3268,N_3286);
xor U3561 (N_3561,N_3338,N_3265);
nor U3562 (N_3562,N_3267,N_3348);
xor U3563 (N_3563,N_3233,N_3387);
xnor U3564 (N_3564,N_3374,N_3264);
nand U3565 (N_3565,N_3207,N_3288);
nand U3566 (N_3566,N_3320,N_3387);
nor U3567 (N_3567,N_3326,N_3367);
and U3568 (N_3568,N_3357,N_3273);
or U3569 (N_3569,N_3332,N_3260);
xnor U3570 (N_3570,N_3338,N_3356);
nand U3571 (N_3571,N_3268,N_3217);
xnor U3572 (N_3572,N_3208,N_3352);
nor U3573 (N_3573,N_3260,N_3326);
nand U3574 (N_3574,N_3399,N_3373);
nand U3575 (N_3575,N_3211,N_3354);
nor U3576 (N_3576,N_3339,N_3288);
and U3577 (N_3577,N_3306,N_3329);
or U3578 (N_3578,N_3311,N_3366);
xnor U3579 (N_3579,N_3260,N_3384);
or U3580 (N_3580,N_3352,N_3362);
nor U3581 (N_3581,N_3311,N_3221);
or U3582 (N_3582,N_3332,N_3238);
or U3583 (N_3583,N_3336,N_3304);
nor U3584 (N_3584,N_3389,N_3254);
and U3585 (N_3585,N_3241,N_3323);
xor U3586 (N_3586,N_3263,N_3392);
xnor U3587 (N_3587,N_3371,N_3300);
nor U3588 (N_3588,N_3369,N_3332);
xnor U3589 (N_3589,N_3317,N_3327);
or U3590 (N_3590,N_3387,N_3270);
xnor U3591 (N_3591,N_3394,N_3337);
nor U3592 (N_3592,N_3293,N_3327);
and U3593 (N_3593,N_3331,N_3245);
and U3594 (N_3594,N_3201,N_3299);
nand U3595 (N_3595,N_3259,N_3217);
and U3596 (N_3596,N_3206,N_3216);
nand U3597 (N_3597,N_3288,N_3397);
nand U3598 (N_3598,N_3347,N_3210);
or U3599 (N_3599,N_3330,N_3205);
xnor U3600 (N_3600,N_3549,N_3406);
nor U3601 (N_3601,N_3460,N_3495);
and U3602 (N_3602,N_3489,N_3517);
and U3603 (N_3603,N_3470,N_3492);
or U3604 (N_3604,N_3473,N_3426);
or U3605 (N_3605,N_3519,N_3497);
nor U3606 (N_3606,N_3518,N_3432);
and U3607 (N_3607,N_3547,N_3560);
nand U3608 (N_3608,N_3593,N_3417);
nor U3609 (N_3609,N_3450,N_3498);
nor U3610 (N_3610,N_3580,N_3506);
or U3611 (N_3611,N_3453,N_3563);
or U3612 (N_3612,N_3404,N_3456);
xnor U3613 (N_3613,N_3402,N_3494);
or U3614 (N_3614,N_3420,N_3505);
xnor U3615 (N_3615,N_3533,N_3477);
or U3616 (N_3616,N_3427,N_3469);
and U3617 (N_3617,N_3446,N_3541);
nor U3618 (N_3618,N_3493,N_3448);
nor U3619 (N_3619,N_3578,N_3485);
xor U3620 (N_3620,N_3561,N_3554);
or U3621 (N_3621,N_3586,N_3438);
nor U3622 (N_3622,N_3548,N_3525);
nand U3623 (N_3623,N_3418,N_3464);
nor U3624 (N_3624,N_3502,N_3577);
or U3625 (N_3625,N_3522,N_3556);
xnor U3626 (N_3626,N_3584,N_3598);
and U3627 (N_3627,N_3421,N_3551);
and U3628 (N_3628,N_3481,N_3490);
and U3629 (N_3629,N_3430,N_3457);
or U3630 (N_3630,N_3546,N_3466);
or U3631 (N_3631,N_3403,N_3447);
or U3632 (N_3632,N_3500,N_3527);
or U3633 (N_3633,N_3413,N_3487);
xor U3634 (N_3634,N_3491,N_3574);
or U3635 (N_3635,N_3520,N_3442);
nor U3636 (N_3636,N_3583,N_3542);
nand U3637 (N_3637,N_3504,N_3559);
and U3638 (N_3638,N_3434,N_3483);
xor U3639 (N_3639,N_3599,N_3445);
or U3640 (N_3640,N_3568,N_3524);
nand U3641 (N_3641,N_3458,N_3440);
nand U3642 (N_3642,N_3597,N_3443);
nand U3643 (N_3643,N_3496,N_3572);
nor U3644 (N_3644,N_3461,N_3422);
and U3645 (N_3645,N_3462,N_3590);
xnor U3646 (N_3646,N_3452,N_3408);
xnor U3647 (N_3647,N_3595,N_3455);
or U3648 (N_3648,N_3410,N_3569);
and U3649 (N_3649,N_3400,N_3585);
and U3650 (N_3650,N_3482,N_3409);
or U3651 (N_3651,N_3509,N_3565);
nor U3652 (N_3652,N_3564,N_3537);
nor U3653 (N_3653,N_3552,N_3571);
and U3654 (N_3654,N_3539,N_3530);
and U3655 (N_3655,N_3401,N_3511);
nand U3656 (N_3656,N_3463,N_3471);
nor U3657 (N_3657,N_3555,N_3573);
xnor U3658 (N_3658,N_3540,N_3449);
xnor U3659 (N_3659,N_3475,N_3562);
and U3660 (N_3660,N_3579,N_3407);
nor U3661 (N_3661,N_3405,N_3587);
nand U3662 (N_3662,N_3431,N_3435);
or U3663 (N_3663,N_3523,N_3451);
nand U3664 (N_3664,N_3553,N_3467);
xor U3665 (N_3665,N_3536,N_3508);
or U3666 (N_3666,N_3479,N_3575);
and U3667 (N_3667,N_3513,N_3544);
xor U3668 (N_3668,N_3570,N_3472);
xor U3669 (N_3669,N_3474,N_3557);
nand U3670 (N_3670,N_3528,N_3558);
nand U3671 (N_3671,N_3424,N_3596);
or U3672 (N_3672,N_3476,N_3567);
and U3673 (N_3673,N_3501,N_3588);
or U3674 (N_3674,N_3412,N_3459);
nor U3675 (N_3675,N_3484,N_3480);
nand U3676 (N_3676,N_3439,N_3419);
nor U3677 (N_3677,N_3550,N_3433);
nor U3678 (N_3678,N_3521,N_3425);
xor U3679 (N_3679,N_3488,N_3566);
nand U3680 (N_3680,N_3514,N_3423);
nand U3681 (N_3681,N_3526,N_3532);
or U3682 (N_3682,N_3592,N_3535);
or U3683 (N_3683,N_3529,N_3415);
nand U3684 (N_3684,N_3429,N_3531);
nand U3685 (N_3685,N_3499,N_3486);
or U3686 (N_3686,N_3576,N_3591);
and U3687 (N_3687,N_3510,N_3411);
xnor U3688 (N_3688,N_3468,N_3416);
nand U3689 (N_3689,N_3516,N_3437);
nor U3690 (N_3690,N_3582,N_3441);
nor U3691 (N_3691,N_3454,N_3538);
nor U3692 (N_3692,N_3589,N_3444);
xor U3693 (N_3693,N_3428,N_3478);
and U3694 (N_3694,N_3545,N_3594);
nand U3695 (N_3695,N_3503,N_3543);
nor U3696 (N_3696,N_3512,N_3436);
or U3697 (N_3697,N_3465,N_3581);
nor U3698 (N_3698,N_3414,N_3515);
or U3699 (N_3699,N_3507,N_3534);
nor U3700 (N_3700,N_3454,N_3509);
and U3701 (N_3701,N_3597,N_3494);
and U3702 (N_3702,N_3500,N_3409);
and U3703 (N_3703,N_3417,N_3569);
or U3704 (N_3704,N_3475,N_3588);
nor U3705 (N_3705,N_3571,N_3593);
nand U3706 (N_3706,N_3404,N_3487);
nor U3707 (N_3707,N_3402,N_3403);
nor U3708 (N_3708,N_3505,N_3597);
nor U3709 (N_3709,N_3589,N_3572);
xnor U3710 (N_3710,N_3460,N_3437);
or U3711 (N_3711,N_3559,N_3400);
or U3712 (N_3712,N_3513,N_3552);
nor U3713 (N_3713,N_3450,N_3495);
or U3714 (N_3714,N_3454,N_3511);
nor U3715 (N_3715,N_3432,N_3474);
xor U3716 (N_3716,N_3421,N_3567);
nor U3717 (N_3717,N_3558,N_3445);
xnor U3718 (N_3718,N_3545,N_3423);
or U3719 (N_3719,N_3553,N_3413);
nand U3720 (N_3720,N_3429,N_3564);
xor U3721 (N_3721,N_3444,N_3503);
and U3722 (N_3722,N_3575,N_3489);
and U3723 (N_3723,N_3492,N_3413);
xnor U3724 (N_3724,N_3472,N_3426);
and U3725 (N_3725,N_3579,N_3405);
or U3726 (N_3726,N_3536,N_3568);
xor U3727 (N_3727,N_3468,N_3558);
nand U3728 (N_3728,N_3522,N_3569);
or U3729 (N_3729,N_3409,N_3538);
xnor U3730 (N_3730,N_3469,N_3502);
nor U3731 (N_3731,N_3557,N_3589);
xnor U3732 (N_3732,N_3501,N_3463);
nor U3733 (N_3733,N_3418,N_3448);
and U3734 (N_3734,N_3413,N_3536);
or U3735 (N_3735,N_3518,N_3516);
or U3736 (N_3736,N_3435,N_3581);
or U3737 (N_3737,N_3494,N_3485);
nand U3738 (N_3738,N_3576,N_3414);
xor U3739 (N_3739,N_3426,N_3425);
xnor U3740 (N_3740,N_3532,N_3533);
or U3741 (N_3741,N_3455,N_3591);
or U3742 (N_3742,N_3484,N_3578);
nand U3743 (N_3743,N_3527,N_3495);
nand U3744 (N_3744,N_3401,N_3499);
xor U3745 (N_3745,N_3535,N_3505);
nor U3746 (N_3746,N_3565,N_3493);
nor U3747 (N_3747,N_3482,N_3577);
nand U3748 (N_3748,N_3482,N_3567);
xnor U3749 (N_3749,N_3434,N_3404);
and U3750 (N_3750,N_3409,N_3522);
and U3751 (N_3751,N_3515,N_3441);
xor U3752 (N_3752,N_3564,N_3464);
nor U3753 (N_3753,N_3500,N_3587);
and U3754 (N_3754,N_3467,N_3492);
xor U3755 (N_3755,N_3469,N_3598);
or U3756 (N_3756,N_3578,N_3410);
and U3757 (N_3757,N_3590,N_3496);
and U3758 (N_3758,N_3490,N_3515);
nand U3759 (N_3759,N_3593,N_3530);
nand U3760 (N_3760,N_3417,N_3410);
nand U3761 (N_3761,N_3492,N_3403);
and U3762 (N_3762,N_3534,N_3597);
nand U3763 (N_3763,N_3475,N_3542);
nand U3764 (N_3764,N_3541,N_3597);
nor U3765 (N_3765,N_3430,N_3411);
and U3766 (N_3766,N_3512,N_3591);
nor U3767 (N_3767,N_3568,N_3525);
or U3768 (N_3768,N_3432,N_3400);
and U3769 (N_3769,N_3468,N_3404);
and U3770 (N_3770,N_3430,N_3585);
nand U3771 (N_3771,N_3464,N_3546);
nand U3772 (N_3772,N_3462,N_3418);
xor U3773 (N_3773,N_3581,N_3445);
or U3774 (N_3774,N_3451,N_3516);
nor U3775 (N_3775,N_3591,N_3599);
nor U3776 (N_3776,N_3567,N_3555);
nor U3777 (N_3777,N_3518,N_3586);
and U3778 (N_3778,N_3409,N_3490);
and U3779 (N_3779,N_3540,N_3557);
and U3780 (N_3780,N_3584,N_3478);
and U3781 (N_3781,N_3516,N_3528);
nor U3782 (N_3782,N_3535,N_3548);
xnor U3783 (N_3783,N_3512,N_3497);
and U3784 (N_3784,N_3418,N_3408);
or U3785 (N_3785,N_3512,N_3571);
nand U3786 (N_3786,N_3550,N_3485);
and U3787 (N_3787,N_3505,N_3596);
nor U3788 (N_3788,N_3566,N_3477);
and U3789 (N_3789,N_3458,N_3566);
xor U3790 (N_3790,N_3524,N_3502);
nand U3791 (N_3791,N_3594,N_3528);
nor U3792 (N_3792,N_3449,N_3554);
or U3793 (N_3793,N_3481,N_3578);
and U3794 (N_3794,N_3416,N_3506);
nor U3795 (N_3795,N_3598,N_3537);
and U3796 (N_3796,N_3462,N_3416);
and U3797 (N_3797,N_3428,N_3545);
and U3798 (N_3798,N_3426,N_3565);
xor U3799 (N_3799,N_3581,N_3493);
or U3800 (N_3800,N_3650,N_3770);
xor U3801 (N_3801,N_3753,N_3761);
nor U3802 (N_3802,N_3752,N_3697);
nor U3803 (N_3803,N_3696,N_3744);
nor U3804 (N_3804,N_3667,N_3669);
and U3805 (N_3805,N_3642,N_3663);
or U3806 (N_3806,N_3647,N_3689);
nand U3807 (N_3807,N_3732,N_3799);
nand U3808 (N_3808,N_3639,N_3608);
or U3809 (N_3809,N_3680,N_3660);
nor U3810 (N_3810,N_3609,N_3622);
and U3811 (N_3811,N_3794,N_3740);
xnor U3812 (N_3812,N_3726,N_3727);
xnor U3813 (N_3813,N_3638,N_3754);
or U3814 (N_3814,N_3798,N_3618);
nor U3815 (N_3815,N_3699,N_3755);
xnor U3816 (N_3816,N_3735,N_3777);
nor U3817 (N_3817,N_3709,N_3614);
nor U3818 (N_3818,N_3653,N_3652);
and U3819 (N_3819,N_3664,N_3778);
nand U3820 (N_3820,N_3651,N_3640);
and U3821 (N_3821,N_3792,N_3678);
nor U3822 (N_3822,N_3665,N_3644);
nor U3823 (N_3823,N_3655,N_3722);
xnor U3824 (N_3824,N_3635,N_3739);
nor U3825 (N_3825,N_3780,N_3705);
or U3826 (N_3826,N_3704,N_3685);
and U3827 (N_3827,N_3672,N_3748);
and U3828 (N_3828,N_3751,N_3648);
nand U3829 (N_3829,N_3781,N_3769);
and U3830 (N_3830,N_3700,N_3782);
and U3831 (N_3831,N_3602,N_3677);
nor U3832 (N_3832,N_3624,N_3716);
xor U3833 (N_3833,N_3715,N_3750);
and U3834 (N_3834,N_3757,N_3646);
nor U3835 (N_3835,N_3641,N_3633);
and U3836 (N_3836,N_3707,N_3723);
and U3837 (N_3837,N_3675,N_3758);
nor U3838 (N_3838,N_3733,N_3785);
xnor U3839 (N_3839,N_3615,N_3725);
nand U3840 (N_3840,N_3773,N_3737);
xor U3841 (N_3841,N_3661,N_3788);
nand U3842 (N_3842,N_3712,N_3643);
xor U3843 (N_3843,N_3654,N_3631);
xnor U3844 (N_3844,N_3742,N_3759);
or U3845 (N_3845,N_3666,N_3698);
or U3846 (N_3846,N_3606,N_3747);
nand U3847 (N_3847,N_3714,N_3637);
or U3848 (N_3848,N_3687,N_3625);
and U3849 (N_3849,N_3718,N_3783);
and U3850 (N_3850,N_3779,N_3749);
nor U3851 (N_3851,N_3670,N_3766);
xnor U3852 (N_3852,N_3713,N_3605);
or U3853 (N_3853,N_3724,N_3676);
or U3854 (N_3854,N_3656,N_3765);
or U3855 (N_3855,N_3619,N_3600);
xnor U3856 (N_3856,N_3682,N_3623);
or U3857 (N_3857,N_3789,N_3786);
nor U3858 (N_3858,N_3763,N_3708);
xnor U3859 (N_3859,N_3774,N_3632);
nor U3860 (N_3860,N_3694,N_3610);
nor U3861 (N_3861,N_3673,N_3603);
or U3862 (N_3862,N_3719,N_3791);
xor U3863 (N_3863,N_3681,N_3775);
xor U3864 (N_3864,N_3691,N_3688);
nor U3865 (N_3865,N_3621,N_3686);
or U3866 (N_3866,N_3745,N_3706);
nand U3867 (N_3867,N_3702,N_3787);
and U3868 (N_3868,N_3649,N_3627);
nand U3869 (N_3869,N_3668,N_3604);
xor U3870 (N_3870,N_3795,N_3626);
or U3871 (N_3871,N_3693,N_3738);
and U3872 (N_3872,N_3692,N_3730);
nor U3873 (N_3873,N_3797,N_3729);
and U3874 (N_3874,N_3762,N_3690);
nor U3875 (N_3875,N_3746,N_3743);
nand U3876 (N_3876,N_3628,N_3645);
or U3877 (N_3877,N_3703,N_3616);
nand U3878 (N_3878,N_3784,N_3768);
xnor U3879 (N_3879,N_3728,N_3620);
xor U3880 (N_3880,N_3657,N_3695);
xor U3881 (N_3881,N_3710,N_3636);
or U3882 (N_3882,N_3607,N_3683);
nor U3883 (N_3883,N_3658,N_3629);
or U3884 (N_3884,N_3767,N_3796);
xnor U3885 (N_3885,N_3662,N_3630);
or U3886 (N_3886,N_3711,N_3793);
or U3887 (N_3887,N_3756,N_3772);
nor U3888 (N_3888,N_3659,N_3720);
nand U3889 (N_3889,N_3613,N_3736);
xor U3890 (N_3890,N_3717,N_3679);
and U3891 (N_3891,N_3617,N_3764);
nor U3892 (N_3892,N_3612,N_3731);
and U3893 (N_3893,N_3776,N_3734);
or U3894 (N_3894,N_3760,N_3674);
or U3895 (N_3895,N_3701,N_3741);
xnor U3896 (N_3896,N_3634,N_3684);
xnor U3897 (N_3897,N_3771,N_3601);
nand U3898 (N_3898,N_3611,N_3721);
nand U3899 (N_3899,N_3671,N_3790);
or U3900 (N_3900,N_3707,N_3749);
nor U3901 (N_3901,N_3738,N_3794);
xnor U3902 (N_3902,N_3729,N_3792);
nand U3903 (N_3903,N_3681,N_3702);
and U3904 (N_3904,N_3735,N_3609);
nand U3905 (N_3905,N_3731,N_3616);
nor U3906 (N_3906,N_3704,N_3749);
nor U3907 (N_3907,N_3766,N_3796);
and U3908 (N_3908,N_3790,N_3702);
xor U3909 (N_3909,N_3735,N_3645);
nor U3910 (N_3910,N_3730,N_3652);
and U3911 (N_3911,N_3767,N_3610);
xnor U3912 (N_3912,N_3796,N_3691);
xor U3913 (N_3913,N_3681,N_3755);
and U3914 (N_3914,N_3685,N_3708);
xnor U3915 (N_3915,N_3606,N_3615);
nor U3916 (N_3916,N_3616,N_3757);
or U3917 (N_3917,N_3600,N_3680);
and U3918 (N_3918,N_3760,N_3763);
nand U3919 (N_3919,N_3765,N_3688);
nand U3920 (N_3920,N_3702,N_3720);
xor U3921 (N_3921,N_3721,N_3746);
xnor U3922 (N_3922,N_3673,N_3687);
nor U3923 (N_3923,N_3771,N_3737);
and U3924 (N_3924,N_3671,N_3677);
nor U3925 (N_3925,N_3674,N_3692);
or U3926 (N_3926,N_3605,N_3704);
xor U3927 (N_3927,N_3696,N_3761);
nand U3928 (N_3928,N_3787,N_3713);
or U3929 (N_3929,N_3664,N_3633);
xor U3930 (N_3930,N_3793,N_3732);
nand U3931 (N_3931,N_3798,N_3690);
and U3932 (N_3932,N_3695,N_3615);
nor U3933 (N_3933,N_3604,N_3618);
nor U3934 (N_3934,N_3730,N_3731);
or U3935 (N_3935,N_3610,N_3777);
or U3936 (N_3936,N_3681,N_3669);
nor U3937 (N_3937,N_3690,N_3633);
and U3938 (N_3938,N_3640,N_3610);
xnor U3939 (N_3939,N_3789,N_3726);
or U3940 (N_3940,N_3767,N_3789);
or U3941 (N_3941,N_3781,N_3771);
nor U3942 (N_3942,N_3718,N_3772);
xnor U3943 (N_3943,N_3620,N_3793);
nand U3944 (N_3944,N_3727,N_3658);
and U3945 (N_3945,N_3772,N_3708);
nor U3946 (N_3946,N_3610,N_3772);
and U3947 (N_3947,N_3759,N_3736);
and U3948 (N_3948,N_3636,N_3783);
nor U3949 (N_3949,N_3706,N_3686);
nor U3950 (N_3950,N_3654,N_3614);
xor U3951 (N_3951,N_3669,N_3736);
and U3952 (N_3952,N_3755,N_3731);
nand U3953 (N_3953,N_3608,N_3642);
xor U3954 (N_3954,N_3669,N_3612);
nor U3955 (N_3955,N_3601,N_3744);
nor U3956 (N_3956,N_3657,N_3624);
and U3957 (N_3957,N_3799,N_3772);
nand U3958 (N_3958,N_3709,N_3651);
and U3959 (N_3959,N_3768,N_3741);
nor U3960 (N_3960,N_3746,N_3688);
or U3961 (N_3961,N_3610,N_3778);
or U3962 (N_3962,N_3623,N_3619);
xnor U3963 (N_3963,N_3675,N_3704);
or U3964 (N_3964,N_3686,N_3727);
nor U3965 (N_3965,N_3669,N_3677);
xor U3966 (N_3966,N_3791,N_3609);
and U3967 (N_3967,N_3656,N_3711);
and U3968 (N_3968,N_3721,N_3763);
and U3969 (N_3969,N_3626,N_3792);
nor U3970 (N_3970,N_3782,N_3651);
nand U3971 (N_3971,N_3724,N_3796);
xor U3972 (N_3972,N_3730,N_3691);
xor U3973 (N_3973,N_3720,N_3655);
xor U3974 (N_3974,N_3782,N_3703);
nand U3975 (N_3975,N_3699,N_3745);
xnor U3976 (N_3976,N_3743,N_3656);
and U3977 (N_3977,N_3602,N_3745);
nand U3978 (N_3978,N_3734,N_3727);
or U3979 (N_3979,N_3675,N_3732);
nor U3980 (N_3980,N_3642,N_3701);
nand U3981 (N_3981,N_3646,N_3676);
xnor U3982 (N_3982,N_3640,N_3738);
nor U3983 (N_3983,N_3697,N_3613);
and U3984 (N_3984,N_3693,N_3622);
nand U3985 (N_3985,N_3702,N_3783);
and U3986 (N_3986,N_3739,N_3753);
or U3987 (N_3987,N_3709,N_3797);
nand U3988 (N_3988,N_3799,N_3694);
nand U3989 (N_3989,N_3731,N_3772);
and U3990 (N_3990,N_3731,N_3685);
and U3991 (N_3991,N_3770,N_3627);
xnor U3992 (N_3992,N_3618,N_3795);
or U3993 (N_3993,N_3621,N_3794);
and U3994 (N_3994,N_3737,N_3780);
or U3995 (N_3995,N_3723,N_3688);
xnor U3996 (N_3996,N_3611,N_3747);
nand U3997 (N_3997,N_3690,N_3781);
nor U3998 (N_3998,N_3708,N_3780);
and U3999 (N_3999,N_3795,N_3758);
and U4000 (N_4000,N_3881,N_3910);
xnor U4001 (N_4001,N_3984,N_3823);
or U4002 (N_4002,N_3946,N_3845);
nor U4003 (N_4003,N_3816,N_3821);
nand U4004 (N_4004,N_3942,N_3998);
and U4005 (N_4005,N_3976,N_3980);
or U4006 (N_4006,N_3992,N_3920);
xor U4007 (N_4007,N_3907,N_3955);
and U4008 (N_4008,N_3892,N_3990);
and U4009 (N_4009,N_3827,N_3801);
or U4010 (N_4010,N_3915,N_3906);
or U4011 (N_4011,N_3864,N_3891);
xor U4012 (N_4012,N_3939,N_3988);
and U4013 (N_4013,N_3850,N_3838);
nand U4014 (N_4014,N_3909,N_3900);
xnor U4015 (N_4015,N_3828,N_3833);
or U4016 (N_4016,N_3888,N_3814);
or U4017 (N_4017,N_3812,N_3974);
and U4018 (N_4018,N_3804,N_3951);
and U4019 (N_4019,N_3839,N_3822);
and U4020 (N_4020,N_3897,N_3894);
nand U4021 (N_4021,N_3935,N_3825);
or U4022 (N_4022,N_3913,N_3918);
nor U4023 (N_4023,N_3805,N_3862);
nor U4024 (N_4024,N_3965,N_3912);
xor U4025 (N_4025,N_3882,N_3972);
nand U4026 (N_4026,N_3869,N_3978);
nand U4027 (N_4027,N_3880,N_3923);
and U4028 (N_4028,N_3847,N_3886);
xor U4029 (N_4029,N_3904,N_3849);
or U4030 (N_4030,N_3943,N_3962);
xnor U4031 (N_4031,N_3809,N_3859);
nand U4032 (N_4032,N_3985,N_3930);
and U4033 (N_4033,N_3963,N_3879);
nor U4034 (N_4034,N_3863,N_3875);
xnor U4035 (N_4035,N_3952,N_3934);
nor U4036 (N_4036,N_3947,N_3977);
nand U4037 (N_4037,N_3853,N_3959);
nand U4038 (N_4038,N_3903,N_3948);
nor U4039 (N_4039,N_3926,N_3840);
nor U4040 (N_4040,N_3818,N_3994);
nor U4041 (N_4041,N_3914,N_3928);
nor U4042 (N_4042,N_3803,N_3945);
or U4043 (N_4043,N_3929,N_3961);
nor U4044 (N_4044,N_3931,N_3884);
nor U4045 (N_4045,N_3848,N_3970);
or U4046 (N_4046,N_3867,N_3968);
or U4047 (N_4047,N_3933,N_3831);
nor U4048 (N_4048,N_3989,N_3979);
xnor U4049 (N_4049,N_3890,N_3973);
nor U4050 (N_4050,N_3983,N_3820);
xnor U4051 (N_4051,N_3878,N_3981);
or U4052 (N_4052,N_3834,N_3986);
nand U4053 (N_4053,N_3830,N_3922);
xor U4054 (N_4054,N_3868,N_3919);
and U4055 (N_4055,N_3877,N_3806);
and U4056 (N_4056,N_3911,N_3819);
nor U4057 (N_4057,N_3832,N_3960);
nor U4058 (N_4058,N_3873,N_3885);
nand U4059 (N_4059,N_3811,N_3921);
and U4060 (N_4060,N_3902,N_3995);
and U4061 (N_4061,N_3856,N_3971);
nor U4062 (N_4062,N_3872,N_3846);
xnor U4063 (N_4063,N_3861,N_3944);
and U4064 (N_4064,N_3997,N_3855);
and U4065 (N_4065,N_3829,N_3975);
and U4066 (N_4066,N_3844,N_3949);
and U4067 (N_4067,N_3987,N_3836);
and U4068 (N_4068,N_3813,N_3842);
xor U4069 (N_4069,N_3800,N_3993);
nand U4070 (N_4070,N_3843,N_3953);
nand U4071 (N_4071,N_3866,N_3893);
nand U4072 (N_4072,N_3815,N_3940);
or U4073 (N_4073,N_3883,N_3950);
and U4074 (N_4074,N_3901,N_3941);
and U4075 (N_4075,N_3924,N_3810);
or U4076 (N_4076,N_3932,N_3826);
and U4077 (N_4077,N_3982,N_3967);
or U4078 (N_4078,N_3996,N_3991);
xnor U4079 (N_4079,N_3837,N_3969);
and U4080 (N_4080,N_3876,N_3954);
nand U4081 (N_4081,N_3927,N_3937);
xnor U4082 (N_4082,N_3874,N_3899);
and U4083 (N_4083,N_3807,N_3824);
xnor U4084 (N_4084,N_3835,N_3857);
xnor U4085 (N_4085,N_3808,N_3852);
nand U4086 (N_4086,N_3817,N_3896);
or U4087 (N_4087,N_3860,N_3895);
or U4088 (N_4088,N_3958,N_3854);
or U4089 (N_4089,N_3851,N_3905);
nor U4090 (N_4090,N_3908,N_3925);
and U4091 (N_4091,N_3841,N_3870);
nand U4092 (N_4092,N_3938,N_3865);
or U4093 (N_4093,N_3964,N_3802);
and U4094 (N_4094,N_3887,N_3956);
nor U4095 (N_4095,N_3917,N_3936);
or U4096 (N_4096,N_3916,N_3966);
xnor U4097 (N_4097,N_3999,N_3889);
xor U4098 (N_4098,N_3898,N_3871);
and U4099 (N_4099,N_3858,N_3957);
nor U4100 (N_4100,N_3979,N_3905);
nor U4101 (N_4101,N_3874,N_3896);
xor U4102 (N_4102,N_3924,N_3891);
nand U4103 (N_4103,N_3864,N_3920);
xnor U4104 (N_4104,N_3880,N_3861);
and U4105 (N_4105,N_3923,N_3868);
xor U4106 (N_4106,N_3801,N_3931);
nor U4107 (N_4107,N_3864,N_3851);
nand U4108 (N_4108,N_3970,N_3950);
xnor U4109 (N_4109,N_3830,N_3817);
or U4110 (N_4110,N_3874,N_3892);
and U4111 (N_4111,N_3809,N_3929);
xnor U4112 (N_4112,N_3991,N_3902);
xnor U4113 (N_4113,N_3899,N_3915);
xnor U4114 (N_4114,N_3867,N_3846);
xnor U4115 (N_4115,N_3844,N_3887);
nand U4116 (N_4116,N_3854,N_3817);
or U4117 (N_4117,N_3852,N_3815);
xor U4118 (N_4118,N_3927,N_3955);
nor U4119 (N_4119,N_3933,N_3900);
and U4120 (N_4120,N_3986,N_3875);
or U4121 (N_4121,N_3950,N_3955);
nor U4122 (N_4122,N_3844,N_3816);
nor U4123 (N_4123,N_3856,N_3879);
nand U4124 (N_4124,N_3830,N_3933);
and U4125 (N_4125,N_3850,N_3969);
xor U4126 (N_4126,N_3981,N_3924);
and U4127 (N_4127,N_3918,N_3936);
or U4128 (N_4128,N_3863,N_3821);
nor U4129 (N_4129,N_3864,N_3925);
and U4130 (N_4130,N_3908,N_3883);
and U4131 (N_4131,N_3918,N_3999);
or U4132 (N_4132,N_3869,N_3861);
nand U4133 (N_4133,N_3840,N_3854);
or U4134 (N_4134,N_3947,N_3920);
xor U4135 (N_4135,N_3974,N_3971);
nor U4136 (N_4136,N_3815,N_3875);
nor U4137 (N_4137,N_3935,N_3888);
and U4138 (N_4138,N_3852,N_3935);
xor U4139 (N_4139,N_3971,N_3894);
and U4140 (N_4140,N_3988,N_3992);
nand U4141 (N_4141,N_3881,N_3951);
nand U4142 (N_4142,N_3873,N_3979);
nor U4143 (N_4143,N_3968,N_3979);
or U4144 (N_4144,N_3889,N_3895);
nor U4145 (N_4145,N_3960,N_3807);
and U4146 (N_4146,N_3865,N_3936);
nand U4147 (N_4147,N_3986,N_3852);
xor U4148 (N_4148,N_3956,N_3883);
or U4149 (N_4149,N_3929,N_3930);
and U4150 (N_4150,N_3884,N_3873);
or U4151 (N_4151,N_3945,N_3900);
xor U4152 (N_4152,N_3995,N_3884);
nor U4153 (N_4153,N_3877,N_3937);
and U4154 (N_4154,N_3946,N_3979);
nand U4155 (N_4155,N_3987,N_3975);
and U4156 (N_4156,N_3848,N_3908);
nand U4157 (N_4157,N_3900,N_3966);
nand U4158 (N_4158,N_3827,N_3963);
nand U4159 (N_4159,N_3854,N_3925);
xnor U4160 (N_4160,N_3977,N_3849);
and U4161 (N_4161,N_3979,N_3862);
and U4162 (N_4162,N_3876,N_3854);
xor U4163 (N_4163,N_3876,N_3971);
nor U4164 (N_4164,N_3946,N_3895);
and U4165 (N_4165,N_3902,N_3820);
nand U4166 (N_4166,N_3858,N_3864);
and U4167 (N_4167,N_3805,N_3860);
nand U4168 (N_4168,N_3853,N_3894);
nor U4169 (N_4169,N_3823,N_3832);
or U4170 (N_4170,N_3924,N_3986);
and U4171 (N_4171,N_3960,N_3984);
and U4172 (N_4172,N_3811,N_3841);
nand U4173 (N_4173,N_3940,N_3951);
xor U4174 (N_4174,N_3933,N_3921);
xor U4175 (N_4175,N_3819,N_3901);
and U4176 (N_4176,N_3810,N_3914);
nor U4177 (N_4177,N_3973,N_3875);
nor U4178 (N_4178,N_3854,N_3827);
nand U4179 (N_4179,N_3807,N_3922);
xnor U4180 (N_4180,N_3851,N_3937);
nand U4181 (N_4181,N_3912,N_3949);
nor U4182 (N_4182,N_3915,N_3892);
and U4183 (N_4183,N_3926,N_3879);
and U4184 (N_4184,N_3990,N_3949);
nand U4185 (N_4185,N_3920,N_3828);
and U4186 (N_4186,N_3940,N_3871);
xnor U4187 (N_4187,N_3841,N_3859);
nor U4188 (N_4188,N_3813,N_3975);
and U4189 (N_4189,N_3989,N_3924);
nand U4190 (N_4190,N_3821,N_3888);
xor U4191 (N_4191,N_3896,N_3867);
nand U4192 (N_4192,N_3807,N_3860);
nand U4193 (N_4193,N_3952,N_3933);
and U4194 (N_4194,N_3950,N_3935);
xnor U4195 (N_4195,N_3965,N_3933);
nand U4196 (N_4196,N_3855,N_3905);
and U4197 (N_4197,N_3864,N_3877);
nand U4198 (N_4198,N_3965,N_3907);
xnor U4199 (N_4199,N_3942,N_3982);
or U4200 (N_4200,N_4062,N_4162);
nand U4201 (N_4201,N_4040,N_4069);
nand U4202 (N_4202,N_4073,N_4108);
nand U4203 (N_4203,N_4014,N_4024);
nand U4204 (N_4204,N_4180,N_4083);
nor U4205 (N_4205,N_4025,N_4046);
or U4206 (N_4206,N_4159,N_4179);
nor U4207 (N_4207,N_4037,N_4116);
and U4208 (N_4208,N_4186,N_4063);
nor U4209 (N_4209,N_4154,N_4100);
nand U4210 (N_4210,N_4161,N_4006);
or U4211 (N_4211,N_4175,N_4156);
and U4212 (N_4212,N_4009,N_4044);
nor U4213 (N_4213,N_4047,N_4127);
and U4214 (N_4214,N_4051,N_4032);
and U4215 (N_4215,N_4131,N_4199);
nor U4216 (N_4216,N_4042,N_4057);
xnor U4217 (N_4217,N_4048,N_4089);
nor U4218 (N_4218,N_4023,N_4039);
or U4219 (N_4219,N_4145,N_4173);
nand U4220 (N_4220,N_4123,N_4115);
and U4221 (N_4221,N_4169,N_4004);
xor U4222 (N_4222,N_4177,N_4184);
nand U4223 (N_4223,N_4005,N_4084);
nor U4224 (N_4224,N_4003,N_4031);
xnor U4225 (N_4225,N_4026,N_4007);
nand U4226 (N_4226,N_4114,N_4150);
nand U4227 (N_4227,N_4020,N_4078);
nand U4228 (N_4228,N_4129,N_4136);
xor U4229 (N_4229,N_4105,N_4170);
xnor U4230 (N_4230,N_4076,N_4091);
nor U4231 (N_4231,N_4112,N_4163);
or U4232 (N_4232,N_4178,N_4144);
nand U4233 (N_4233,N_4135,N_4053);
nor U4234 (N_4234,N_4172,N_4030);
or U4235 (N_4235,N_4096,N_4194);
and U4236 (N_4236,N_4052,N_4142);
nand U4237 (N_4237,N_4121,N_4125);
and U4238 (N_4238,N_4110,N_4064);
xor U4239 (N_4239,N_4017,N_4176);
nor U4240 (N_4240,N_4068,N_4167);
xor U4241 (N_4241,N_4081,N_4043);
nor U4242 (N_4242,N_4058,N_4072);
nor U4243 (N_4243,N_4067,N_4138);
xor U4244 (N_4244,N_4124,N_4001);
or U4245 (N_4245,N_4097,N_4033);
xnor U4246 (N_4246,N_4034,N_4189);
nor U4247 (N_4247,N_4122,N_4029);
or U4248 (N_4248,N_4041,N_4158);
and U4249 (N_4249,N_4019,N_4092);
or U4250 (N_4250,N_4107,N_4012);
or U4251 (N_4251,N_4008,N_4140);
or U4252 (N_4252,N_4120,N_4147);
xnor U4253 (N_4253,N_4060,N_4056);
and U4254 (N_4254,N_4182,N_4198);
nand U4255 (N_4255,N_4071,N_4010);
xnor U4256 (N_4256,N_4049,N_4059);
nor U4257 (N_4257,N_4036,N_4011);
and U4258 (N_4258,N_4111,N_4197);
and U4259 (N_4259,N_4132,N_4185);
xor U4260 (N_4260,N_4168,N_4146);
nor U4261 (N_4261,N_4134,N_4151);
and U4262 (N_4262,N_4143,N_4035);
and U4263 (N_4263,N_4165,N_4174);
nor U4264 (N_4264,N_4113,N_4187);
nor U4265 (N_4265,N_4117,N_4079);
or U4266 (N_4266,N_4166,N_4149);
and U4267 (N_4267,N_4016,N_4139);
or U4268 (N_4268,N_4061,N_4088);
or U4269 (N_4269,N_4028,N_4104);
nand U4270 (N_4270,N_4045,N_4128);
and U4271 (N_4271,N_4119,N_4086);
and U4272 (N_4272,N_4103,N_4191);
nor U4273 (N_4273,N_4155,N_4022);
and U4274 (N_4274,N_4015,N_4018);
xnor U4275 (N_4275,N_4082,N_4080);
xnor U4276 (N_4276,N_4190,N_4183);
and U4277 (N_4277,N_4137,N_4098);
nor U4278 (N_4278,N_4070,N_4160);
and U4279 (N_4279,N_4153,N_4085);
xor U4280 (N_4280,N_4095,N_4181);
nor U4281 (N_4281,N_4133,N_4087);
nand U4282 (N_4282,N_4074,N_4118);
nor U4283 (N_4283,N_4193,N_4164);
or U4284 (N_4284,N_4075,N_4141);
or U4285 (N_4285,N_4090,N_4188);
xnor U4286 (N_4286,N_4055,N_4192);
nand U4287 (N_4287,N_4065,N_4027);
nor U4288 (N_4288,N_4099,N_4038);
xnor U4289 (N_4289,N_4130,N_4126);
nor U4290 (N_4290,N_4054,N_4157);
and U4291 (N_4291,N_4195,N_4171);
nor U4292 (N_4292,N_4102,N_4077);
xnor U4293 (N_4293,N_4021,N_4109);
and U4294 (N_4294,N_4094,N_4002);
nand U4295 (N_4295,N_4066,N_4106);
nand U4296 (N_4296,N_4148,N_4152);
nor U4297 (N_4297,N_4000,N_4101);
xnor U4298 (N_4298,N_4050,N_4013);
and U4299 (N_4299,N_4196,N_4093);
nor U4300 (N_4300,N_4150,N_4082);
nor U4301 (N_4301,N_4014,N_4194);
or U4302 (N_4302,N_4023,N_4073);
nor U4303 (N_4303,N_4016,N_4022);
and U4304 (N_4304,N_4157,N_4057);
nand U4305 (N_4305,N_4036,N_4170);
nand U4306 (N_4306,N_4009,N_4187);
and U4307 (N_4307,N_4068,N_4124);
nor U4308 (N_4308,N_4195,N_4070);
or U4309 (N_4309,N_4052,N_4175);
nor U4310 (N_4310,N_4151,N_4193);
and U4311 (N_4311,N_4118,N_4180);
xor U4312 (N_4312,N_4053,N_4030);
or U4313 (N_4313,N_4052,N_4025);
nor U4314 (N_4314,N_4022,N_4177);
nand U4315 (N_4315,N_4059,N_4102);
nand U4316 (N_4316,N_4058,N_4144);
and U4317 (N_4317,N_4169,N_4001);
or U4318 (N_4318,N_4022,N_4100);
xor U4319 (N_4319,N_4125,N_4164);
nand U4320 (N_4320,N_4060,N_4019);
or U4321 (N_4321,N_4183,N_4165);
or U4322 (N_4322,N_4106,N_4031);
or U4323 (N_4323,N_4022,N_4143);
nand U4324 (N_4324,N_4116,N_4191);
nor U4325 (N_4325,N_4073,N_4061);
and U4326 (N_4326,N_4081,N_4102);
or U4327 (N_4327,N_4041,N_4069);
xnor U4328 (N_4328,N_4150,N_4039);
or U4329 (N_4329,N_4058,N_4005);
nand U4330 (N_4330,N_4064,N_4067);
nand U4331 (N_4331,N_4141,N_4168);
xor U4332 (N_4332,N_4050,N_4146);
xor U4333 (N_4333,N_4165,N_4145);
nand U4334 (N_4334,N_4010,N_4149);
nand U4335 (N_4335,N_4198,N_4166);
nand U4336 (N_4336,N_4157,N_4052);
nor U4337 (N_4337,N_4170,N_4148);
nor U4338 (N_4338,N_4157,N_4096);
or U4339 (N_4339,N_4131,N_4041);
or U4340 (N_4340,N_4194,N_4139);
nor U4341 (N_4341,N_4092,N_4079);
and U4342 (N_4342,N_4190,N_4080);
xor U4343 (N_4343,N_4010,N_4015);
xnor U4344 (N_4344,N_4067,N_4075);
xnor U4345 (N_4345,N_4009,N_4182);
nand U4346 (N_4346,N_4165,N_4078);
nor U4347 (N_4347,N_4176,N_4095);
nand U4348 (N_4348,N_4098,N_4103);
nor U4349 (N_4349,N_4009,N_4047);
and U4350 (N_4350,N_4009,N_4137);
nor U4351 (N_4351,N_4110,N_4135);
xor U4352 (N_4352,N_4003,N_4107);
and U4353 (N_4353,N_4142,N_4101);
xor U4354 (N_4354,N_4199,N_4069);
xnor U4355 (N_4355,N_4046,N_4106);
or U4356 (N_4356,N_4142,N_4120);
nor U4357 (N_4357,N_4058,N_4149);
xnor U4358 (N_4358,N_4123,N_4182);
nor U4359 (N_4359,N_4143,N_4061);
xor U4360 (N_4360,N_4177,N_4024);
nand U4361 (N_4361,N_4091,N_4025);
and U4362 (N_4362,N_4119,N_4017);
and U4363 (N_4363,N_4145,N_4032);
nor U4364 (N_4364,N_4190,N_4061);
nand U4365 (N_4365,N_4179,N_4064);
nand U4366 (N_4366,N_4146,N_4086);
nor U4367 (N_4367,N_4062,N_4095);
and U4368 (N_4368,N_4195,N_4064);
xnor U4369 (N_4369,N_4118,N_4142);
or U4370 (N_4370,N_4095,N_4157);
or U4371 (N_4371,N_4055,N_4131);
xnor U4372 (N_4372,N_4196,N_4076);
nand U4373 (N_4373,N_4084,N_4081);
or U4374 (N_4374,N_4128,N_4046);
nor U4375 (N_4375,N_4158,N_4072);
or U4376 (N_4376,N_4085,N_4032);
nand U4377 (N_4377,N_4052,N_4140);
xnor U4378 (N_4378,N_4173,N_4070);
nor U4379 (N_4379,N_4111,N_4020);
nor U4380 (N_4380,N_4139,N_4006);
nor U4381 (N_4381,N_4066,N_4013);
or U4382 (N_4382,N_4161,N_4003);
or U4383 (N_4383,N_4068,N_4019);
xnor U4384 (N_4384,N_4024,N_4121);
and U4385 (N_4385,N_4077,N_4120);
xor U4386 (N_4386,N_4015,N_4178);
or U4387 (N_4387,N_4032,N_4101);
and U4388 (N_4388,N_4013,N_4041);
xnor U4389 (N_4389,N_4163,N_4169);
nor U4390 (N_4390,N_4076,N_4189);
nand U4391 (N_4391,N_4065,N_4028);
xor U4392 (N_4392,N_4189,N_4120);
nand U4393 (N_4393,N_4131,N_4085);
or U4394 (N_4394,N_4144,N_4071);
xnor U4395 (N_4395,N_4069,N_4034);
nor U4396 (N_4396,N_4026,N_4125);
or U4397 (N_4397,N_4191,N_4073);
or U4398 (N_4398,N_4024,N_4186);
xor U4399 (N_4399,N_4100,N_4043);
nor U4400 (N_4400,N_4244,N_4234);
or U4401 (N_4401,N_4247,N_4366);
or U4402 (N_4402,N_4384,N_4305);
nor U4403 (N_4403,N_4308,N_4232);
and U4404 (N_4404,N_4383,N_4381);
and U4405 (N_4405,N_4278,N_4386);
nor U4406 (N_4406,N_4289,N_4246);
and U4407 (N_4407,N_4358,N_4322);
nand U4408 (N_4408,N_4370,N_4367);
and U4409 (N_4409,N_4346,N_4375);
nand U4410 (N_4410,N_4251,N_4213);
and U4411 (N_4411,N_4240,N_4226);
nor U4412 (N_4412,N_4336,N_4345);
nor U4413 (N_4413,N_4365,N_4248);
or U4414 (N_4414,N_4307,N_4295);
or U4415 (N_4415,N_4235,N_4355);
or U4416 (N_4416,N_4343,N_4229);
nor U4417 (N_4417,N_4283,N_4364);
or U4418 (N_4418,N_4260,N_4220);
and U4419 (N_4419,N_4316,N_4395);
or U4420 (N_4420,N_4337,N_4396);
nand U4421 (N_4421,N_4362,N_4200);
nand U4422 (N_4422,N_4382,N_4211);
nand U4423 (N_4423,N_4369,N_4378);
and U4424 (N_4424,N_4368,N_4321);
and U4425 (N_4425,N_4205,N_4301);
nor U4426 (N_4426,N_4224,N_4217);
or U4427 (N_4427,N_4252,N_4284);
xnor U4428 (N_4428,N_4363,N_4311);
nor U4429 (N_4429,N_4238,N_4390);
or U4430 (N_4430,N_4243,N_4288);
nor U4431 (N_4431,N_4222,N_4285);
xor U4432 (N_4432,N_4318,N_4389);
and U4433 (N_4433,N_4331,N_4227);
xor U4434 (N_4434,N_4344,N_4256);
nor U4435 (N_4435,N_4253,N_4201);
nor U4436 (N_4436,N_4261,N_4372);
nand U4437 (N_4437,N_4236,N_4249);
nand U4438 (N_4438,N_4310,N_4399);
nand U4439 (N_4439,N_4280,N_4275);
nor U4440 (N_4440,N_4324,N_4350);
and U4441 (N_4441,N_4373,N_4304);
nor U4442 (N_4442,N_4287,N_4203);
and U4443 (N_4443,N_4279,N_4274);
or U4444 (N_4444,N_4290,N_4377);
nand U4445 (N_4445,N_4320,N_4385);
nand U4446 (N_4446,N_4323,N_4380);
nand U4447 (N_4447,N_4272,N_4263);
xnor U4448 (N_4448,N_4202,N_4347);
nand U4449 (N_4449,N_4300,N_4398);
nand U4450 (N_4450,N_4268,N_4333);
nand U4451 (N_4451,N_4326,N_4269);
xnor U4452 (N_4452,N_4335,N_4264);
nand U4453 (N_4453,N_4237,N_4233);
nand U4454 (N_4454,N_4221,N_4298);
and U4455 (N_4455,N_4352,N_4214);
xor U4456 (N_4456,N_4327,N_4204);
and U4457 (N_4457,N_4348,N_4277);
or U4458 (N_4458,N_4306,N_4293);
xnor U4459 (N_4459,N_4267,N_4239);
nand U4460 (N_4460,N_4357,N_4339);
and U4461 (N_4461,N_4297,N_4328);
nor U4462 (N_4462,N_4259,N_4262);
nor U4463 (N_4463,N_4241,N_4282);
nand U4464 (N_4464,N_4271,N_4265);
nand U4465 (N_4465,N_4250,N_4245);
xor U4466 (N_4466,N_4317,N_4266);
nand U4467 (N_4467,N_4309,N_4354);
xor U4468 (N_4468,N_4315,N_4360);
nand U4469 (N_4469,N_4356,N_4242);
xor U4470 (N_4470,N_4349,N_4257);
xor U4471 (N_4471,N_4294,N_4299);
xor U4472 (N_4472,N_4330,N_4314);
nand U4473 (N_4473,N_4292,N_4230);
nand U4474 (N_4474,N_4359,N_4281);
nand U4475 (N_4475,N_4388,N_4332);
xor U4476 (N_4476,N_4225,N_4329);
xnor U4477 (N_4477,N_4258,N_4270);
nand U4478 (N_4478,N_4371,N_4218);
nor U4479 (N_4479,N_4353,N_4231);
and U4480 (N_4480,N_4276,N_4391);
nor U4481 (N_4481,N_4273,N_4361);
and U4482 (N_4482,N_4342,N_4341);
or U4483 (N_4483,N_4215,N_4208);
and U4484 (N_4484,N_4209,N_4312);
nor U4485 (N_4485,N_4379,N_4219);
and U4486 (N_4486,N_4319,N_4374);
and U4487 (N_4487,N_4228,N_4325);
nand U4488 (N_4488,N_4376,N_4303);
or U4489 (N_4489,N_4334,N_4392);
nand U4490 (N_4490,N_4340,N_4313);
nor U4491 (N_4491,N_4207,N_4338);
xor U4492 (N_4492,N_4394,N_4351);
or U4493 (N_4493,N_4397,N_4206);
nand U4494 (N_4494,N_4255,N_4254);
and U4495 (N_4495,N_4286,N_4291);
xnor U4496 (N_4496,N_4216,N_4302);
xor U4497 (N_4497,N_4387,N_4393);
and U4498 (N_4498,N_4212,N_4296);
and U4499 (N_4499,N_4223,N_4210);
nand U4500 (N_4500,N_4301,N_4391);
xnor U4501 (N_4501,N_4340,N_4351);
nor U4502 (N_4502,N_4233,N_4372);
and U4503 (N_4503,N_4352,N_4232);
nor U4504 (N_4504,N_4200,N_4299);
and U4505 (N_4505,N_4263,N_4288);
nand U4506 (N_4506,N_4376,N_4273);
and U4507 (N_4507,N_4242,N_4248);
and U4508 (N_4508,N_4315,N_4304);
and U4509 (N_4509,N_4325,N_4252);
nor U4510 (N_4510,N_4263,N_4393);
and U4511 (N_4511,N_4219,N_4251);
and U4512 (N_4512,N_4346,N_4224);
nor U4513 (N_4513,N_4275,N_4277);
nand U4514 (N_4514,N_4257,N_4225);
and U4515 (N_4515,N_4315,N_4254);
and U4516 (N_4516,N_4307,N_4213);
xor U4517 (N_4517,N_4255,N_4323);
nand U4518 (N_4518,N_4343,N_4306);
nand U4519 (N_4519,N_4260,N_4253);
and U4520 (N_4520,N_4257,N_4363);
and U4521 (N_4521,N_4304,N_4290);
nor U4522 (N_4522,N_4217,N_4243);
xnor U4523 (N_4523,N_4327,N_4225);
nand U4524 (N_4524,N_4392,N_4238);
nand U4525 (N_4525,N_4378,N_4376);
nand U4526 (N_4526,N_4378,N_4314);
nor U4527 (N_4527,N_4258,N_4205);
and U4528 (N_4528,N_4214,N_4317);
xor U4529 (N_4529,N_4228,N_4345);
or U4530 (N_4530,N_4368,N_4266);
nor U4531 (N_4531,N_4205,N_4354);
xor U4532 (N_4532,N_4282,N_4221);
xnor U4533 (N_4533,N_4264,N_4337);
and U4534 (N_4534,N_4218,N_4317);
xor U4535 (N_4535,N_4351,N_4226);
and U4536 (N_4536,N_4355,N_4379);
nand U4537 (N_4537,N_4347,N_4252);
nand U4538 (N_4538,N_4293,N_4282);
nand U4539 (N_4539,N_4372,N_4362);
and U4540 (N_4540,N_4290,N_4369);
or U4541 (N_4541,N_4236,N_4291);
or U4542 (N_4542,N_4380,N_4304);
and U4543 (N_4543,N_4264,N_4298);
nand U4544 (N_4544,N_4330,N_4397);
nand U4545 (N_4545,N_4349,N_4358);
nor U4546 (N_4546,N_4379,N_4260);
and U4547 (N_4547,N_4256,N_4264);
and U4548 (N_4548,N_4311,N_4343);
or U4549 (N_4549,N_4251,N_4353);
and U4550 (N_4550,N_4217,N_4303);
nand U4551 (N_4551,N_4216,N_4363);
or U4552 (N_4552,N_4277,N_4296);
nand U4553 (N_4553,N_4375,N_4251);
xor U4554 (N_4554,N_4396,N_4390);
and U4555 (N_4555,N_4372,N_4399);
nor U4556 (N_4556,N_4299,N_4271);
and U4557 (N_4557,N_4313,N_4222);
nand U4558 (N_4558,N_4247,N_4219);
nand U4559 (N_4559,N_4219,N_4359);
nor U4560 (N_4560,N_4307,N_4267);
xnor U4561 (N_4561,N_4206,N_4221);
and U4562 (N_4562,N_4207,N_4231);
and U4563 (N_4563,N_4235,N_4366);
nor U4564 (N_4564,N_4301,N_4283);
nor U4565 (N_4565,N_4270,N_4301);
and U4566 (N_4566,N_4322,N_4252);
and U4567 (N_4567,N_4299,N_4318);
nand U4568 (N_4568,N_4325,N_4384);
nand U4569 (N_4569,N_4384,N_4212);
nor U4570 (N_4570,N_4241,N_4299);
or U4571 (N_4571,N_4231,N_4343);
or U4572 (N_4572,N_4241,N_4256);
nand U4573 (N_4573,N_4364,N_4331);
nor U4574 (N_4574,N_4345,N_4317);
and U4575 (N_4575,N_4375,N_4283);
nor U4576 (N_4576,N_4243,N_4245);
and U4577 (N_4577,N_4206,N_4300);
and U4578 (N_4578,N_4330,N_4213);
and U4579 (N_4579,N_4341,N_4214);
nor U4580 (N_4580,N_4330,N_4375);
nand U4581 (N_4581,N_4231,N_4314);
nor U4582 (N_4582,N_4253,N_4345);
xnor U4583 (N_4583,N_4308,N_4283);
nor U4584 (N_4584,N_4213,N_4211);
nand U4585 (N_4585,N_4393,N_4351);
or U4586 (N_4586,N_4339,N_4285);
and U4587 (N_4587,N_4296,N_4386);
or U4588 (N_4588,N_4388,N_4227);
or U4589 (N_4589,N_4263,N_4201);
nor U4590 (N_4590,N_4365,N_4383);
nor U4591 (N_4591,N_4338,N_4388);
xor U4592 (N_4592,N_4317,N_4249);
or U4593 (N_4593,N_4291,N_4388);
nor U4594 (N_4594,N_4293,N_4337);
and U4595 (N_4595,N_4238,N_4339);
nand U4596 (N_4596,N_4227,N_4298);
and U4597 (N_4597,N_4308,N_4355);
and U4598 (N_4598,N_4232,N_4201);
nor U4599 (N_4599,N_4224,N_4312);
and U4600 (N_4600,N_4470,N_4485);
xnor U4601 (N_4601,N_4477,N_4590);
or U4602 (N_4602,N_4592,N_4463);
xor U4603 (N_4603,N_4599,N_4448);
nand U4604 (N_4604,N_4566,N_4551);
nand U4605 (N_4605,N_4428,N_4583);
xnor U4606 (N_4606,N_4402,N_4472);
and U4607 (N_4607,N_4575,N_4579);
xor U4608 (N_4608,N_4567,N_4416);
nor U4609 (N_4609,N_4437,N_4562);
xnor U4610 (N_4610,N_4513,N_4527);
and U4611 (N_4611,N_4500,N_4464);
nor U4612 (N_4612,N_4552,N_4438);
xnor U4613 (N_4613,N_4507,N_4582);
xnor U4614 (N_4614,N_4439,N_4491);
nor U4615 (N_4615,N_4473,N_4496);
nand U4616 (N_4616,N_4517,N_4430);
nand U4617 (N_4617,N_4581,N_4518);
xnor U4618 (N_4618,N_4434,N_4556);
nand U4619 (N_4619,N_4492,N_4521);
or U4620 (N_4620,N_4523,N_4542);
nand U4621 (N_4621,N_4429,N_4431);
or U4622 (N_4622,N_4411,N_4539);
nand U4623 (N_4623,N_4432,N_4421);
nor U4624 (N_4624,N_4482,N_4455);
and U4625 (N_4625,N_4515,N_4487);
or U4626 (N_4626,N_4418,N_4405);
and U4627 (N_4627,N_4474,N_4536);
nor U4628 (N_4628,N_4449,N_4593);
or U4629 (N_4629,N_4506,N_4458);
and U4630 (N_4630,N_4445,N_4489);
and U4631 (N_4631,N_4502,N_4412);
and U4632 (N_4632,N_4471,N_4454);
nand U4633 (N_4633,N_4444,N_4565);
nor U4634 (N_4634,N_4525,N_4529);
nor U4635 (N_4635,N_4588,N_4465);
or U4636 (N_4636,N_4501,N_4570);
xnor U4637 (N_4637,N_4469,N_4443);
xor U4638 (N_4638,N_4435,N_4451);
and U4639 (N_4639,N_4541,N_4433);
and U4640 (N_4640,N_4450,N_4481);
and U4641 (N_4641,N_4544,N_4591);
and U4642 (N_4642,N_4425,N_4505);
and U4643 (N_4643,N_4484,N_4457);
xnor U4644 (N_4644,N_4598,N_4490);
nand U4645 (N_4645,N_4503,N_4400);
xnor U4646 (N_4646,N_4414,N_4440);
xor U4647 (N_4647,N_4597,N_4595);
nor U4648 (N_4648,N_4537,N_4554);
xnor U4649 (N_4649,N_4587,N_4528);
and U4650 (N_4650,N_4584,N_4569);
nand U4651 (N_4651,N_4585,N_4531);
xnor U4652 (N_4652,N_4514,N_4422);
nand U4653 (N_4653,N_4538,N_4409);
or U4654 (N_4654,N_4511,N_4512);
nor U4655 (N_4655,N_4532,N_4546);
and U4656 (N_4656,N_4488,N_4419);
or U4657 (N_4657,N_4533,N_4526);
nand U4658 (N_4658,N_4519,N_4480);
nor U4659 (N_4659,N_4547,N_4446);
or U4660 (N_4660,N_4540,N_4543);
and U4661 (N_4661,N_4589,N_4466);
xor U4662 (N_4662,N_4453,N_4545);
nor U4663 (N_4663,N_4550,N_4407);
nor U4664 (N_4664,N_4410,N_4548);
and U4665 (N_4665,N_4403,N_4459);
or U4666 (N_4666,N_4498,N_4564);
xor U4667 (N_4667,N_4460,N_4535);
nor U4668 (N_4668,N_4571,N_4559);
nand U4669 (N_4669,N_4555,N_4499);
or U4670 (N_4670,N_4596,N_4553);
or U4671 (N_4671,N_4549,N_4586);
nor U4672 (N_4672,N_4572,N_4494);
and U4673 (N_4673,N_4462,N_4504);
xor U4674 (N_4674,N_4479,N_4524);
or U4675 (N_4675,N_4478,N_4577);
or U4676 (N_4676,N_4476,N_4408);
and U4677 (N_4677,N_4520,N_4576);
nor U4678 (N_4678,N_4468,N_4497);
nand U4679 (N_4679,N_4420,N_4442);
and U4680 (N_4680,N_4413,N_4461);
xnor U4681 (N_4681,N_4594,N_4568);
nand U4682 (N_4682,N_4580,N_4534);
and U4683 (N_4683,N_4426,N_4558);
and U4684 (N_4684,N_4417,N_4493);
nor U4685 (N_4685,N_4401,N_4467);
and U4686 (N_4686,N_4509,N_4427);
nand U4687 (N_4687,N_4475,N_4486);
xor U4688 (N_4688,N_4424,N_4415);
nand U4689 (N_4689,N_4456,N_4530);
nor U4690 (N_4690,N_4423,N_4452);
nor U4691 (N_4691,N_4447,N_4557);
xor U4692 (N_4692,N_4560,N_4495);
xor U4693 (N_4693,N_4483,N_4441);
and U4694 (N_4694,N_4578,N_4406);
or U4695 (N_4695,N_4510,N_4516);
nor U4696 (N_4696,N_4573,N_4522);
nand U4697 (N_4697,N_4574,N_4436);
xor U4698 (N_4698,N_4404,N_4561);
or U4699 (N_4699,N_4508,N_4563);
and U4700 (N_4700,N_4457,N_4471);
xor U4701 (N_4701,N_4597,N_4416);
xor U4702 (N_4702,N_4594,N_4436);
nor U4703 (N_4703,N_4437,N_4556);
and U4704 (N_4704,N_4598,N_4485);
and U4705 (N_4705,N_4465,N_4596);
nand U4706 (N_4706,N_4578,N_4496);
nand U4707 (N_4707,N_4485,N_4484);
or U4708 (N_4708,N_4563,N_4510);
nand U4709 (N_4709,N_4470,N_4437);
nor U4710 (N_4710,N_4440,N_4462);
and U4711 (N_4711,N_4425,N_4503);
xnor U4712 (N_4712,N_4532,N_4483);
or U4713 (N_4713,N_4531,N_4465);
nand U4714 (N_4714,N_4447,N_4599);
nor U4715 (N_4715,N_4527,N_4521);
xnor U4716 (N_4716,N_4589,N_4501);
and U4717 (N_4717,N_4426,N_4488);
nand U4718 (N_4718,N_4539,N_4437);
nand U4719 (N_4719,N_4594,N_4427);
nor U4720 (N_4720,N_4510,N_4580);
or U4721 (N_4721,N_4521,N_4458);
nand U4722 (N_4722,N_4447,N_4590);
xnor U4723 (N_4723,N_4463,N_4589);
xnor U4724 (N_4724,N_4588,N_4564);
or U4725 (N_4725,N_4408,N_4456);
or U4726 (N_4726,N_4571,N_4411);
nor U4727 (N_4727,N_4587,N_4540);
nor U4728 (N_4728,N_4553,N_4523);
xnor U4729 (N_4729,N_4408,N_4416);
or U4730 (N_4730,N_4405,N_4542);
nand U4731 (N_4731,N_4540,N_4503);
or U4732 (N_4732,N_4405,N_4491);
xnor U4733 (N_4733,N_4573,N_4416);
and U4734 (N_4734,N_4462,N_4542);
or U4735 (N_4735,N_4498,N_4575);
nand U4736 (N_4736,N_4556,N_4429);
and U4737 (N_4737,N_4513,N_4536);
xor U4738 (N_4738,N_4486,N_4590);
or U4739 (N_4739,N_4474,N_4525);
nor U4740 (N_4740,N_4537,N_4498);
nor U4741 (N_4741,N_4471,N_4453);
xor U4742 (N_4742,N_4449,N_4482);
and U4743 (N_4743,N_4559,N_4449);
and U4744 (N_4744,N_4568,N_4565);
nor U4745 (N_4745,N_4441,N_4489);
nand U4746 (N_4746,N_4483,N_4433);
nand U4747 (N_4747,N_4490,N_4462);
nand U4748 (N_4748,N_4458,N_4520);
or U4749 (N_4749,N_4502,N_4474);
and U4750 (N_4750,N_4579,N_4441);
nor U4751 (N_4751,N_4416,N_4532);
xnor U4752 (N_4752,N_4466,N_4475);
and U4753 (N_4753,N_4587,N_4541);
and U4754 (N_4754,N_4452,N_4582);
nand U4755 (N_4755,N_4473,N_4560);
or U4756 (N_4756,N_4556,N_4499);
or U4757 (N_4757,N_4576,N_4552);
xor U4758 (N_4758,N_4438,N_4567);
or U4759 (N_4759,N_4473,N_4431);
nand U4760 (N_4760,N_4596,N_4541);
xnor U4761 (N_4761,N_4475,N_4498);
nand U4762 (N_4762,N_4514,N_4413);
nand U4763 (N_4763,N_4462,N_4446);
or U4764 (N_4764,N_4419,N_4424);
nand U4765 (N_4765,N_4567,N_4481);
or U4766 (N_4766,N_4473,N_4416);
and U4767 (N_4767,N_4461,N_4541);
xnor U4768 (N_4768,N_4465,N_4475);
nor U4769 (N_4769,N_4451,N_4578);
and U4770 (N_4770,N_4465,N_4421);
nor U4771 (N_4771,N_4450,N_4445);
or U4772 (N_4772,N_4469,N_4581);
nand U4773 (N_4773,N_4402,N_4460);
and U4774 (N_4774,N_4513,N_4530);
or U4775 (N_4775,N_4455,N_4554);
xnor U4776 (N_4776,N_4522,N_4566);
or U4777 (N_4777,N_4454,N_4591);
xnor U4778 (N_4778,N_4498,N_4468);
nor U4779 (N_4779,N_4573,N_4424);
nand U4780 (N_4780,N_4425,N_4538);
xor U4781 (N_4781,N_4425,N_4588);
or U4782 (N_4782,N_4545,N_4427);
nand U4783 (N_4783,N_4409,N_4433);
nor U4784 (N_4784,N_4446,N_4455);
and U4785 (N_4785,N_4479,N_4505);
xor U4786 (N_4786,N_4598,N_4496);
nand U4787 (N_4787,N_4419,N_4535);
or U4788 (N_4788,N_4425,N_4578);
nand U4789 (N_4789,N_4585,N_4565);
and U4790 (N_4790,N_4440,N_4499);
or U4791 (N_4791,N_4413,N_4489);
nor U4792 (N_4792,N_4579,N_4584);
nand U4793 (N_4793,N_4515,N_4570);
xnor U4794 (N_4794,N_4420,N_4545);
nor U4795 (N_4795,N_4479,N_4578);
and U4796 (N_4796,N_4467,N_4560);
nor U4797 (N_4797,N_4429,N_4441);
xnor U4798 (N_4798,N_4565,N_4548);
nor U4799 (N_4799,N_4480,N_4490);
nor U4800 (N_4800,N_4617,N_4624);
nor U4801 (N_4801,N_4757,N_4703);
xor U4802 (N_4802,N_4753,N_4727);
nand U4803 (N_4803,N_4786,N_4649);
and U4804 (N_4804,N_4738,N_4618);
nand U4805 (N_4805,N_4758,N_4730);
xnor U4806 (N_4806,N_4756,N_4683);
xnor U4807 (N_4807,N_4712,N_4791);
or U4808 (N_4808,N_4680,N_4611);
nor U4809 (N_4809,N_4735,N_4783);
nor U4810 (N_4810,N_4781,N_4760);
nand U4811 (N_4811,N_4769,N_4613);
nor U4812 (N_4812,N_4655,N_4685);
nor U4813 (N_4813,N_4736,N_4795);
and U4814 (N_4814,N_4720,N_4654);
nand U4815 (N_4815,N_4749,N_4750);
nand U4816 (N_4816,N_4622,N_4716);
nor U4817 (N_4817,N_4652,N_4722);
or U4818 (N_4818,N_4714,N_4774);
or U4819 (N_4819,N_4710,N_4635);
nand U4820 (N_4820,N_4693,N_4612);
nand U4821 (N_4821,N_4694,N_4733);
nand U4822 (N_4822,N_4796,N_4637);
nor U4823 (N_4823,N_4616,N_4775);
and U4824 (N_4824,N_4789,N_4793);
and U4825 (N_4825,N_4762,N_4662);
and U4826 (N_4826,N_4653,N_4681);
or U4827 (N_4827,N_4602,N_4747);
and U4828 (N_4828,N_4724,N_4755);
xnor U4829 (N_4829,N_4642,N_4670);
nand U4830 (N_4830,N_4661,N_4676);
nand U4831 (N_4831,N_4644,N_4682);
and U4832 (N_4832,N_4744,N_4764);
and U4833 (N_4833,N_4679,N_4748);
nor U4834 (N_4834,N_4631,N_4659);
nor U4835 (N_4835,N_4698,N_4706);
or U4836 (N_4836,N_4672,N_4606);
xor U4837 (N_4837,N_4713,N_4717);
nand U4838 (N_4838,N_4636,N_4677);
and U4839 (N_4839,N_4741,N_4700);
and U4840 (N_4840,N_4684,N_4785);
xor U4841 (N_4841,N_4797,N_4726);
nand U4842 (N_4842,N_4686,N_4643);
xor U4843 (N_4843,N_4790,N_4719);
nor U4844 (N_4844,N_4751,N_4620);
and U4845 (N_4845,N_4605,N_4792);
nand U4846 (N_4846,N_4725,N_4634);
nor U4847 (N_4847,N_4678,N_4615);
and U4848 (N_4848,N_4777,N_4664);
xnor U4849 (N_4849,N_4767,N_4692);
nand U4850 (N_4850,N_4699,N_4673);
xor U4851 (N_4851,N_4708,N_4711);
nand U4852 (N_4852,N_4763,N_4731);
nand U4853 (N_4853,N_4675,N_4721);
nand U4854 (N_4854,N_4743,N_4604);
nand U4855 (N_4855,N_4705,N_4665);
or U4856 (N_4856,N_4776,N_4632);
and U4857 (N_4857,N_4688,N_4794);
or U4858 (N_4858,N_4667,N_4697);
xnor U4859 (N_4859,N_4627,N_4666);
nor U4860 (N_4860,N_4729,N_4773);
xor U4861 (N_4861,N_4765,N_4650);
nand U4862 (N_4862,N_4734,N_4746);
nand U4863 (N_4863,N_4609,N_4778);
nor U4864 (N_4864,N_4732,N_4770);
xor U4865 (N_4865,N_4779,N_4646);
nand U4866 (N_4866,N_4651,N_4715);
nor U4867 (N_4867,N_4648,N_4660);
nand U4868 (N_4868,N_4621,N_4623);
nor U4869 (N_4869,N_4772,N_4740);
nor U4870 (N_4870,N_4671,N_4752);
nor U4871 (N_4871,N_4787,N_4614);
and U4872 (N_4872,N_4780,N_4641);
xnor U4873 (N_4873,N_4601,N_4647);
or U4874 (N_4874,N_4625,N_4603);
and U4875 (N_4875,N_4728,N_4695);
xor U4876 (N_4876,N_4669,N_4619);
and U4877 (N_4877,N_4626,N_4742);
nand U4878 (N_4878,N_4630,N_4739);
xnor U4879 (N_4879,N_4737,N_4663);
or U4880 (N_4880,N_4610,N_4798);
xnor U4881 (N_4881,N_4656,N_4718);
or U4882 (N_4882,N_4771,N_4782);
nand U4883 (N_4883,N_4628,N_4707);
or U4884 (N_4884,N_4701,N_4639);
nand U4885 (N_4885,N_4784,N_4689);
and U4886 (N_4886,N_4657,N_4600);
or U4887 (N_4887,N_4768,N_4629);
nor U4888 (N_4888,N_4608,N_4723);
nand U4889 (N_4889,N_4674,N_4754);
and U4890 (N_4890,N_4709,N_4607);
nor U4891 (N_4891,N_4691,N_4658);
nor U4892 (N_4892,N_4761,N_4745);
xor U4893 (N_4893,N_4759,N_4645);
xor U4894 (N_4894,N_4799,N_4687);
nor U4895 (N_4895,N_4690,N_4640);
nor U4896 (N_4896,N_4766,N_4696);
xnor U4897 (N_4897,N_4788,N_4633);
or U4898 (N_4898,N_4638,N_4704);
nor U4899 (N_4899,N_4702,N_4668);
nor U4900 (N_4900,N_4716,N_4610);
and U4901 (N_4901,N_4663,N_4724);
and U4902 (N_4902,N_4614,N_4641);
xor U4903 (N_4903,N_4720,N_4647);
or U4904 (N_4904,N_4729,N_4624);
nor U4905 (N_4905,N_4751,N_4614);
or U4906 (N_4906,N_4619,N_4708);
xor U4907 (N_4907,N_4734,N_4790);
nor U4908 (N_4908,N_4680,N_4652);
nand U4909 (N_4909,N_4776,N_4672);
or U4910 (N_4910,N_4718,N_4753);
xnor U4911 (N_4911,N_4676,N_4684);
or U4912 (N_4912,N_4764,N_4697);
nand U4913 (N_4913,N_4707,N_4634);
or U4914 (N_4914,N_4719,N_4721);
xor U4915 (N_4915,N_4664,N_4617);
and U4916 (N_4916,N_4772,N_4709);
or U4917 (N_4917,N_4717,N_4789);
xor U4918 (N_4918,N_4784,N_4670);
or U4919 (N_4919,N_4765,N_4726);
nor U4920 (N_4920,N_4601,N_4698);
nor U4921 (N_4921,N_4752,N_4767);
xnor U4922 (N_4922,N_4767,N_4693);
or U4923 (N_4923,N_4634,N_4619);
and U4924 (N_4924,N_4647,N_4734);
nand U4925 (N_4925,N_4650,N_4641);
and U4926 (N_4926,N_4773,N_4723);
nor U4927 (N_4927,N_4762,N_4660);
nor U4928 (N_4928,N_4760,N_4684);
or U4929 (N_4929,N_4648,N_4646);
nor U4930 (N_4930,N_4616,N_4657);
and U4931 (N_4931,N_4719,N_4739);
and U4932 (N_4932,N_4694,N_4708);
or U4933 (N_4933,N_4785,N_4675);
and U4934 (N_4934,N_4718,N_4678);
nor U4935 (N_4935,N_4623,N_4643);
and U4936 (N_4936,N_4665,N_4735);
and U4937 (N_4937,N_4658,N_4750);
or U4938 (N_4938,N_4612,N_4646);
nor U4939 (N_4939,N_4736,N_4707);
or U4940 (N_4940,N_4735,N_4697);
and U4941 (N_4941,N_4601,N_4699);
and U4942 (N_4942,N_4642,N_4710);
xor U4943 (N_4943,N_4766,N_4770);
and U4944 (N_4944,N_4776,N_4634);
xnor U4945 (N_4945,N_4610,N_4612);
and U4946 (N_4946,N_4789,N_4784);
nor U4947 (N_4947,N_4799,N_4647);
nand U4948 (N_4948,N_4775,N_4633);
nand U4949 (N_4949,N_4724,N_4617);
nand U4950 (N_4950,N_4650,N_4706);
nand U4951 (N_4951,N_4763,N_4777);
and U4952 (N_4952,N_4702,N_4688);
nor U4953 (N_4953,N_4796,N_4629);
and U4954 (N_4954,N_4735,N_4660);
xor U4955 (N_4955,N_4640,N_4771);
or U4956 (N_4956,N_4636,N_4717);
nand U4957 (N_4957,N_4618,N_4772);
nand U4958 (N_4958,N_4713,N_4770);
or U4959 (N_4959,N_4708,N_4635);
nor U4960 (N_4960,N_4771,N_4758);
and U4961 (N_4961,N_4785,N_4665);
nand U4962 (N_4962,N_4603,N_4708);
or U4963 (N_4963,N_4686,N_4733);
xnor U4964 (N_4964,N_4749,N_4607);
or U4965 (N_4965,N_4744,N_4753);
nor U4966 (N_4966,N_4718,N_4789);
xor U4967 (N_4967,N_4725,N_4721);
and U4968 (N_4968,N_4693,N_4684);
xnor U4969 (N_4969,N_4660,N_4668);
or U4970 (N_4970,N_4734,N_4777);
nand U4971 (N_4971,N_4733,N_4717);
nor U4972 (N_4972,N_4788,N_4698);
xnor U4973 (N_4973,N_4675,N_4705);
and U4974 (N_4974,N_4729,N_4746);
or U4975 (N_4975,N_4772,N_4686);
xnor U4976 (N_4976,N_4704,N_4667);
and U4977 (N_4977,N_4686,N_4607);
or U4978 (N_4978,N_4780,N_4773);
nor U4979 (N_4979,N_4677,N_4754);
and U4980 (N_4980,N_4694,N_4729);
or U4981 (N_4981,N_4753,N_4742);
or U4982 (N_4982,N_4657,N_4629);
and U4983 (N_4983,N_4622,N_4725);
xor U4984 (N_4984,N_4666,N_4735);
and U4985 (N_4985,N_4669,N_4760);
and U4986 (N_4986,N_4722,N_4720);
and U4987 (N_4987,N_4631,N_4675);
nand U4988 (N_4988,N_4689,N_4736);
nand U4989 (N_4989,N_4723,N_4795);
nand U4990 (N_4990,N_4769,N_4643);
nor U4991 (N_4991,N_4699,N_4650);
nand U4992 (N_4992,N_4706,N_4732);
and U4993 (N_4993,N_4739,N_4715);
or U4994 (N_4994,N_4681,N_4798);
or U4995 (N_4995,N_4636,N_4653);
or U4996 (N_4996,N_4710,N_4798);
or U4997 (N_4997,N_4745,N_4641);
or U4998 (N_4998,N_4707,N_4610);
nand U4999 (N_4999,N_4693,N_4668);
or U5000 (N_5000,N_4891,N_4856);
nand U5001 (N_5001,N_4930,N_4813);
nor U5002 (N_5002,N_4844,N_4977);
xor U5003 (N_5003,N_4944,N_4952);
or U5004 (N_5004,N_4826,N_4836);
or U5005 (N_5005,N_4913,N_4890);
or U5006 (N_5006,N_4854,N_4837);
xnor U5007 (N_5007,N_4804,N_4992);
xnor U5008 (N_5008,N_4858,N_4941);
nand U5009 (N_5009,N_4909,N_4898);
nor U5010 (N_5010,N_4865,N_4876);
nand U5011 (N_5011,N_4949,N_4871);
nand U5012 (N_5012,N_4892,N_4985);
and U5013 (N_5013,N_4907,N_4961);
and U5014 (N_5014,N_4827,N_4845);
and U5015 (N_5015,N_4995,N_4888);
or U5016 (N_5016,N_4882,N_4936);
nand U5017 (N_5017,N_4934,N_4868);
nand U5018 (N_5018,N_4808,N_4942);
and U5019 (N_5019,N_4911,N_4965);
xnor U5020 (N_5020,N_4846,N_4902);
xor U5021 (N_5021,N_4993,N_4805);
xor U5022 (N_5022,N_4801,N_4839);
and U5023 (N_5023,N_4991,N_4863);
nand U5024 (N_5024,N_4809,N_4974);
nor U5025 (N_5025,N_4953,N_4864);
nand U5026 (N_5026,N_4927,N_4853);
and U5027 (N_5027,N_4917,N_4842);
nand U5028 (N_5028,N_4883,N_4946);
xor U5029 (N_5029,N_4803,N_4861);
nor U5030 (N_5030,N_4960,N_4926);
nor U5031 (N_5031,N_4929,N_4816);
or U5032 (N_5032,N_4951,N_4957);
xor U5033 (N_5033,N_4981,N_4962);
or U5034 (N_5034,N_4894,N_4835);
or U5035 (N_5035,N_4959,N_4878);
nand U5036 (N_5036,N_4859,N_4824);
nand U5037 (N_5037,N_4935,N_4885);
nand U5038 (N_5038,N_4820,N_4975);
and U5039 (N_5039,N_4822,N_4806);
and U5040 (N_5040,N_4931,N_4982);
and U5041 (N_5041,N_4947,N_4921);
nor U5042 (N_5042,N_4880,N_4821);
xnor U5043 (N_5043,N_4850,N_4922);
and U5044 (N_5044,N_4976,N_4849);
nor U5045 (N_5045,N_4905,N_4904);
and U5046 (N_5046,N_4815,N_4938);
nand U5047 (N_5047,N_4989,N_4870);
nor U5048 (N_5048,N_4825,N_4954);
nand U5049 (N_5049,N_4834,N_4895);
nor U5050 (N_5050,N_4994,N_4940);
or U5051 (N_5051,N_4908,N_4851);
nor U5052 (N_5052,N_4969,N_4972);
xor U5053 (N_5053,N_4852,N_4967);
nand U5054 (N_5054,N_4830,N_4920);
nor U5055 (N_5055,N_4963,N_4984);
nor U5056 (N_5056,N_4862,N_4901);
or U5057 (N_5057,N_4906,N_4828);
nand U5058 (N_5058,N_4973,N_4923);
nand U5059 (N_5059,N_4915,N_4866);
and U5060 (N_5060,N_4914,N_4996);
nand U5061 (N_5061,N_4860,N_4843);
xnor U5062 (N_5062,N_4925,N_4829);
or U5063 (N_5063,N_4887,N_4833);
xor U5064 (N_5064,N_4848,N_4988);
or U5065 (N_5065,N_4968,N_4812);
xnor U5066 (N_5066,N_4910,N_4950);
xnor U5067 (N_5067,N_4875,N_4937);
or U5068 (N_5068,N_4838,N_4990);
nand U5069 (N_5069,N_4945,N_4867);
or U5070 (N_5070,N_4823,N_4872);
nor U5071 (N_5071,N_4884,N_4817);
and U5072 (N_5072,N_4847,N_4928);
nand U5073 (N_5073,N_4818,N_4998);
xnor U5074 (N_5074,N_4970,N_4855);
nand U5075 (N_5075,N_4958,N_4877);
and U5076 (N_5076,N_4983,N_4933);
or U5077 (N_5077,N_4948,N_4924);
and U5078 (N_5078,N_4819,N_4919);
nand U5079 (N_5079,N_4943,N_4873);
nand U5080 (N_5080,N_4997,N_4978);
nor U5081 (N_5081,N_4903,N_4840);
nand U5082 (N_5082,N_4896,N_4899);
xnor U5083 (N_5083,N_4966,N_4955);
nor U5084 (N_5084,N_4971,N_4918);
and U5085 (N_5085,N_4889,N_4987);
and U5086 (N_5086,N_4881,N_4879);
xnor U5087 (N_5087,N_4800,N_4897);
nor U5088 (N_5088,N_4810,N_4857);
xor U5089 (N_5089,N_4886,N_4916);
or U5090 (N_5090,N_4980,N_4999);
or U5091 (N_5091,N_4979,N_4811);
xnor U5092 (N_5092,N_4814,N_4956);
nor U5093 (N_5093,N_4807,N_4831);
nor U5094 (N_5094,N_4874,N_4986);
nor U5095 (N_5095,N_4869,N_4900);
or U5096 (N_5096,N_4932,N_4893);
xor U5097 (N_5097,N_4964,N_4841);
or U5098 (N_5098,N_4939,N_4802);
nand U5099 (N_5099,N_4832,N_4912);
nand U5100 (N_5100,N_4871,N_4937);
or U5101 (N_5101,N_4914,N_4865);
or U5102 (N_5102,N_4901,N_4918);
xnor U5103 (N_5103,N_4881,N_4977);
or U5104 (N_5104,N_4945,N_4846);
nand U5105 (N_5105,N_4966,N_4836);
nor U5106 (N_5106,N_4874,N_4925);
nand U5107 (N_5107,N_4932,N_4937);
and U5108 (N_5108,N_4804,N_4979);
nor U5109 (N_5109,N_4999,N_4944);
and U5110 (N_5110,N_4962,N_4902);
nor U5111 (N_5111,N_4902,N_4903);
nand U5112 (N_5112,N_4983,N_4850);
xor U5113 (N_5113,N_4892,N_4960);
nor U5114 (N_5114,N_4918,N_4995);
and U5115 (N_5115,N_4831,N_4927);
nor U5116 (N_5116,N_4839,N_4836);
xor U5117 (N_5117,N_4879,N_4938);
and U5118 (N_5118,N_4905,N_4946);
nand U5119 (N_5119,N_4927,N_4864);
or U5120 (N_5120,N_4838,N_4871);
nand U5121 (N_5121,N_4858,N_4933);
or U5122 (N_5122,N_4926,N_4987);
nand U5123 (N_5123,N_4932,N_4825);
or U5124 (N_5124,N_4970,N_4900);
nor U5125 (N_5125,N_4916,N_4913);
nor U5126 (N_5126,N_4870,N_4843);
xor U5127 (N_5127,N_4907,N_4830);
or U5128 (N_5128,N_4931,N_4995);
nor U5129 (N_5129,N_4995,N_4882);
xnor U5130 (N_5130,N_4994,N_4960);
or U5131 (N_5131,N_4904,N_4871);
and U5132 (N_5132,N_4928,N_4833);
xnor U5133 (N_5133,N_4888,N_4929);
nor U5134 (N_5134,N_4802,N_4853);
nand U5135 (N_5135,N_4885,N_4801);
and U5136 (N_5136,N_4932,N_4820);
xor U5137 (N_5137,N_4984,N_4952);
nand U5138 (N_5138,N_4864,N_4877);
and U5139 (N_5139,N_4905,N_4922);
xnor U5140 (N_5140,N_4999,N_4987);
xnor U5141 (N_5141,N_4849,N_4870);
nor U5142 (N_5142,N_4925,N_4823);
nand U5143 (N_5143,N_4911,N_4822);
nand U5144 (N_5144,N_4800,N_4802);
xnor U5145 (N_5145,N_4910,N_4904);
or U5146 (N_5146,N_4831,N_4983);
nor U5147 (N_5147,N_4944,N_4930);
xor U5148 (N_5148,N_4847,N_4920);
or U5149 (N_5149,N_4893,N_4908);
or U5150 (N_5150,N_4999,N_4898);
xor U5151 (N_5151,N_4983,N_4988);
or U5152 (N_5152,N_4931,N_4944);
xnor U5153 (N_5153,N_4861,N_4877);
nor U5154 (N_5154,N_4907,N_4833);
nand U5155 (N_5155,N_4885,N_4948);
xnor U5156 (N_5156,N_4996,N_4993);
or U5157 (N_5157,N_4922,N_4856);
nand U5158 (N_5158,N_4967,N_4804);
or U5159 (N_5159,N_4925,N_4899);
or U5160 (N_5160,N_4925,N_4883);
nor U5161 (N_5161,N_4922,N_4928);
xnor U5162 (N_5162,N_4895,N_4861);
nand U5163 (N_5163,N_4917,N_4900);
nand U5164 (N_5164,N_4937,N_4974);
nand U5165 (N_5165,N_4939,N_4973);
and U5166 (N_5166,N_4903,N_4969);
nor U5167 (N_5167,N_4912,N_4805);
nor U5168 (N_5168,N_4930,N_4828);
xor U5169 (N_5169,N_4886,N_4853);
xnor U5170 (N_5170,N_4918,N_4888);
nand U5171 (N_5171,N_4874,N_4886);
or U5172 (N_5172,N_4804,N_4870);
xnor U5173 (N_5173,N_4957,N_4882);
xor U5174 (N_5174,N_4844,N_4953);
nand U5175 (N_5175,N_4874,N_4843);
nor U5176 (N_5176,N_4889,N_4903);
nor U5177 (N_5177,N_4891,N_4841);
nand U5178 (N_5178,N_4802,N_4947);
nand U5179 (N_5179,N_4934,N_4820);
nand U5180 (N_5180,N_4965,N_4843);
nand U5181 (N_5181,N_4802,N_4999);
nor U5182 (N_5182,N_4941,N_4968);
nand U5183 (N_5183,N_4946,N_4897);
and U5184 (N_5184,N_4845,N_4969);
xnor U5185 (N_5185,N_4965,N_4852);
xor U5186 (N_5186,N_4967,N_4871);
nand U5187 (N_5187,N_4868,N_4833);
xor U5188 (N_5188,N_4802,N_4955);
nand U5189 (N_5189,N_4829,N_4850);
xnor U5190 (N_5190,N_4990,N_4932);
nand U5191 (N_5191,N_4960,N_4861);
xnor U5192 (N_5192,N_4865,N_4878);
xnor U5193 (N_5193,N_4888,N_4816);
and U5194 (N_5194,N_4902,N_4875);
nor U5195 (N_5195,N_4998,N_4816);
nor U5196 (N_5196,N_4966,N_4956);
or U5197 (N_5197,N_4897,N_4894);
or U5198 (N_5198,N_4870,N_4959);
and U5199 (N_5199,N_4874,N_4947);
and U5200 (N_5200,N_5041,N_5198);
or U5201 (N_5201,N_5106,N_5028);
nor U5202 (N_5202,N_5123,N_5159);
xnor U5203 (N_5203,N_5064,N_5182);
or U5204 (N_5204,N_5141,N_5070);
or U5205 (N_5205,N_5167,N_5194);
nand U5206 (N_5206,N_5017,N_5184);
nor U5207 (N_5207,N_5090,N_5134);
xnor U5208 (N_5208,N_5018,N_5131);
or U5209 (N_5209,N_5195,N_5132);
and U5210 (N_5210,N_5037,N_5163);
xnor U5211 (N_5211,N_5053,N_5170);
and U5212 (N_5212,N_5181,N_5061);
and U5213 (N_5213,N_5110,N_5162);
xor U5214 (N_5214,N_5035,N_5027);
or U5215 (N_5215,N_5021,N_5169);
nand U5216 (N_5216,N_5096,N_5179);
nand U5217 (N_5217,N_5055,N_5078);
nand U5218 (N_5218,N_5072,N_5192);
and U5219 (N_5219,N_5099,N_5080);
or U5220 (N_5220,N_5087,N_5083);
nand U5221 (N_5221,N_5124,N_5190);
nand U5222 (N_5222,N_5039,N_5178);
nor U5223 (N_5223,N_5048,N_5006);
nand U5224 (N_5224,N_5091,N_5156);
nor U5225 (N_5225,N_5020,N_5109);
xnor U5226 (N_5226,N_5177,N_5149);
and U5227 (N_5227,N_5172,N_5101);
or U5228 (N_5228,N_5043,N_5119);
and U5229 (N_5229,N_5145,N_5160);
and U5230 (N_5230,N_5098,N_5157);
nor U5231 (N_5231,N_5089,N_5081);
nor U5232 (N_5232,N_5050,N_5044);
nand U5233 (N_5233,N_5042,N_5153);
or U5234 (N_5234,N_5077,N_5007);
or U5235 (N_5235,N_5173,N_5186);
or U5236 (N_5236,N_5012,N_5082);
nor U5237 (N_5237,N_5144,N_5103);
and U5238 (N_5238,N_5092,N_5111);
xor U5239 (N_5239,N_5002,N_5175);
nor U5240 (N_5240,N_5067,N_5116);
nor U5241 (N_5241,N_5030,N_5117);
and U5242 (N_5242,N_5069,N_5105);
nand U5243 (N_5243,N_5095,N_5112);
and U5244 (N_5244,N_5128,N_5196);
or U5245 (N_5245,N_5088,N_5031);
and U5246 (N_5246,N_5024,N_5188);
or U5247 (N_5247,N_5146,N_5189);
nand U5248 (N_5248,N_5154,N_5097);
nor U5249 (N_5249,N_5122,N_5049);
or U5250 (N_5250,N_5045,N_5150);
and U5251 (N_5251,N_5147,N_5071);
nor U5252 (N_5252,N_5001,N_5022);
xnor U5253 (N_5253,N_5046,N_5056);
and U5254 (N_5254,N_5023,N_5136);
xor U5255 (N_5255,N_5032,N_5137);
and U5256 (N_5256,N_5015,N_5166);
or U5257 (N_5257,N_5010,N_5086);
and U5258 (N_5258,N_5073,N_5054);
nor U5259 (N_5259,N_5094,N_5040);
or U5260 (N_5260,N_5085,N_5065);
xnor U5261 (N_5261,N_5187,N_5129);
and U5262 (N_5262,N_5164,N_5193);
nand U5263 (N_5263,N_5075,N_5114);
or U5264 (N_5264,N_5051,N_5084);
and U5265 (N_5265,N_5093,N_5100);
or U5266 (N_5266,N_5142,N_5118);
or U5267 (N_5267,N_5108,N_5176);
nor U5268 (N_5268,N_5013,N_5019);
and U5269 (N_5269,N_5168,N_5197);
xnor U5270 (N_5270,N_5059,N_5115);
and U5271 (N_5271,N_5025,N_5014);
nor U5272 (N_5272,N_5034,N_5148);
xnor U5273 (N_5273,N_5058,N_5180);
xnor U5274 (N_5274,N_5029,N_5152);
and U5275 (N_5275,N_5135,N_5161);
nor U5276 (N_5276,N_5011,N_5009);
nand U5277 (N_5277,N_5151,N_5033);
xnor U5278 (N_5278,N_5155,N_5133);
xor U5279 (N_5279,N_5016,N_5004);
nand U5280 (N_5280,N_5143,N_5165);
xnor U5281 (N_5281,N_5130,N_5057);
and U5282 (N_5282,N_5066,N_5052);
nand U5283 (N_5283,N_5171,N_5102);
nor U5284 (N_5284,N_5008,N_5062);
and U5285 (N_5285,N_5121,N_5125);
and U5286 (N_5286,N_5063,N_5079);
nor U5287 (N_5287,N_5120,N_5076);
and U5288 (N_5288,N_5038,N_5140);
nand U5289 (N_5289,N_5199,N_5068);
nand U5290 (N_5290,N_5158,N_5113);
or U5291 (N_5291,N_5026,N_5127);
nor U5292 (N_5292,N_5139,N_5036);
or U5293 (N_5293,N_5174,N_5183);
and U5294 (N_5294,N_5104,N_5005);
nand U5295 (N_5295,N_5047,N_5185);
nand U5296 (N_5296,N_5003,N_5126);
nor U5297 (N_5297,N_5138,N_5074);
nand U5298 (N_5298,N_5060,N_5000);
and U5299 (N_5299,N_5107,N_5191);
xor U5300 (N_5300,N_5165,N_5169);
nand U5301 (N_5301,N_5180,N_5050);
or U5302 (N_5302,N_5097,N_5112);
or U5303 (N_5303,N_5123,N_5111);
or U5304 (N_5304,N_5089,N_5164);
or U5305 (N_5305,N_5017,N_5159);
nor U5306 (N_5306,N_5186,N_5184);
or U5307 (N_5307,N_5113,N_5050);
or U5308 (N_5308,N_5158,N_5127);
nand U5309 (N_5309,N_5020,N_5115);
nor U5310 (N_5310,N_5027,N_5038);
or U5311 (N_5311,N_5049,N_5180);
nand U5312 (N_5312,N_5158,N_5015);
or U5313 (N_5313,N_5064,N_5128);
or U5314 (N_5314,N_5143,N_5044);
and U5315 (N_5315,N_5139,N_5004);
nand U5316 (N_5316,N_5019,N_5008);
xor U5317 (N_5317,N_5167,N_5172);
xor U5318 (N_5318,N_5030,N_5088);
nand U5319 (N_5319,N_5008,N_5106);
xor U5320 (N_5320,N_5009,N_5021);
nand U5321 (N_5321,N_5103,N_5099);
nand U5322 (N_5322,N_5172,N_5150);
nor U5323 (N_5323,N_5077,N_5103);
or U5324 (N_5324,N_5135,N_5058);
nand U5325 (N_5325,N_5189,N_5119);
xor U5326 (N_5326,N_5096,N_5002);
or U5327 (N_5327,N_5124,N_5034);
nand U5328 (N_5328,N_5081,N_5182);
and U5329 (N_5329,N_5023,N_5144);
or U5330 (N_5330,N_5057,N_5073);
or U5331 (N_5331,N_5023,N_5068);
or U5332 (N_5332,N_5007,N_5088);
nor U5333 (N_5333,N_5008,N_5176);
nor U5334 (N_5334,N_5009,N_5132);
or U5335 (N_5335,N_5169,N_5188);
and U5336 (N_5336,N_5083,N_5160);
nand U5337 (N_5337,N_5098,N_5073);
xor U5338 (N_5338,N_5093,N_5005);
nand U5339 (N_5339,N_5006,N_5036);
xnor U5340 (N_5340,N_5045,N_5061);
and U5341 (N_5341,N_5026,N_5090);
or U5342 (N_5342,N_5051,N_5160);
or U5343 (N_5343,N_5056,N_5153);
or U5344 (N_5344,N_5177,N_5174);
xor U5345 (N_5345,N_5036,N_5174);
nand U5346 (N_5346,N_5035,N_5034);
and U5347 (N_5347,N_5162,N_5077);
nand U5348 (N_5348,N_5005,N_5125);
nor U5349 (N_5349,N_5086,N_5037);
or U5350 (N_5350,N_5035,N_5104);
nand U5351 (N_5351,N_5022,N_5174);
nand U5352 (N_5352,N_5125,N_5015);
xor U5353 (N_5353,N_5033,N_5065);
nand U5354 (N_5354,N_5159,N_5050);
xnor U5355 (N_5355,N_5073,N_5171);
xnor U5356 (N_5356,N_5089,N_5133);
nand U5357 (N_5357,N_5158,N_5016);
and U5358 (N_5358,N_5171,N_5021);
xor U5359 (N_5359,N_5098,N_5105);
nand U5360 (N_5360,N_5077,N_5172);
xor U5361 (N_5361,N_5012,N_5183);
nand U5362 (N_5362,N_5094,N_5130);
or U5363 (N_5363,N_5063,N_5081);
nand U5364 (N_5364,N_5171,N_5004);
nor U5365 (N_5365,N_5063,N_5132);
xnor U5366 (N_5366,N_5058,N_5063);
or U5367 (N_5367,N_5103,N_5008);
or U5368 (N_5368,N_5118,N_5193);
and U5369 (N_5369,N_5125,N_5163);
nand U5370 (N_5370,N_5144,N_5091);
and U5371 (N_5371,N_5122,N_5054);
and U5372 (N_5372,N_5169,N_5123);
and U5373 (N_5373,N_5190,N_5016);
nor U5374 (N_5374,N_5035,N_5161);
or U5375 (N_5375,N_5067,N_5032);
or U5376 (N_5376,N_5138,N_5191);
xnor U5377 (N_5377,N_5192,N_5146);
or U5378 (N_5378,N_5001,N_5096);
nand U5379 (N_5379,N_5062,N_5161);
nor U5380 (N_5380,N_5016,N_5159);
xor U5381 (N_5381,N_5115,N_5159);
xnor U5382 (N_5382,N_5019,N_5058);
nor U5383 (N_5383,N_5156,N_5093);
xor U5384 (N_5384,N_5045,N_5152);
and U5385 (N_5385,N_5073,N_5092);
and U5386 (N_5386,N_5190,N_5013);
and U5387 (N_5387,N_5050,N_5158);
and U5388 (N_5388,N_5061,N_5062);
nor U5389 (N_5389,N_5085,N_5077);
or U5390 (N_5390,N_5135,N_5075);
nor U5391 (N_5391,N_5047,N_5098);
nand U5392 (N_5392,N_5150,N_5179);
xor U5393 (N_5393,N_5199,N_5030);
nor U5394 (N_5394,N_5149,N_5044);
xor U5395 (N_5395,N_5059,N_5138);
and U5396 (N_5396,N_5087,N_5091);
xor U5397 (N_5397,N_5111,N_5147);
nor U5398 (N_5398,N_5137,N_5196);
or U5399 (N_5399,N_5127,N_5018);
and U5400 (N_5400,N_5308,N_5238);
xor U5401 (N_5401,N_5302,N_5307);
nand U5402 (N_5402,N_5243,N_5393);
xor U5403 (N_5403,N_5374,N_5306);
xor U5404 (N_5404,N_5279,N_5256);
nor U5405 (N_5405,N_5325,N_5204);
nor U5406 (N_5406,N_5331,N_5276);
nand U5407 (N_5407,N_5251,N_5270);
or U5408 (N_5408,N_5346,N_5313);
or U5409 (N_5409,N_5309,N_5336);
nor U5410 (N_5410,N_5376,N_5392);
and U5411 (N_5411,N_5362,N_5310);
nor U5412 (N_5412,N_5277,N_5350);
and U5413 (N_5413,N_5314,N_5343);
or U5414 (N_5414,N_5261,N_5284);
xnor U5415 (N_5415,N_5356,N_5345);
nand U5416 (N_5416,N_5354,N_5207);
or U5417 (N_5417,N_5280,N_5332);
or U5418 (N_5418,N_5287,N_5388);
nor U5419 (N_5419,N_5214,N_5372);
xnor U5420 (N_5420,N_5249,N_5230);
nor U5421 (N_5421,N_5379,N_5295);
nor U5422 (N_5422,N_5337,N_5344);
or U5423 (N_5423,N_5371,N_5361);
or U5424 (N_5424,N_5244,N_5395);
nand U5425 (N_5425,N_5380,N_5351);
xor U5426 (N_5426,N_5367,N_5315);
or U5427 (N_5427,N_5262,N_5268);
xor U5428 (N_5428,N_5381,N_5202);
and U5429 (N_5429,N_5398,N_5209);
nand U5430 (N_5430,N_5291,N_5324);
or U5431 (N_5431,N_5369,N_5352);
nand U5432 (N_5432,N_5228,N_5258);
xnor U5433 (N_5433,N_5382,N_5320);
nor U5434 (N_5434,N_5218,N_5300);
and U5435 (N_5435,N_5357,N_5215);
xor U5436 (N_5436,N_5223,N_5236);
xor U5437 (N_5437,N_5390,N_5281);
and U5438 (N_5438,N_5328,N_5237);
nor U5439 (N_5439,N_5389,N_5377);
xnor U5440 (N_5440,N_5232,N_5327);
xor U5441 (N_5441,N_5304,N_5267);
nand U5442 (N_5442,N_5274,N_5253);
nand U5443 (N_5443,N_5205,N_5342);
nor U5444 (N_5444,N_5335,N_5365);
and U5445 (N_5445,N_5363,N_5241);
nor U5446 (N_5446,N_5222,N_5316);
xor U5447 (N_5447,N_5293,N_5340);
xnor U5448 (N_5448,N_5255,N_5358);
or U5449 (N_5449,N_5233,N_5278);
or U5450 (N_5450,N_5397,N_5245);
or U5451 (N_5451,N_5264,N_5334);
xor U5452 (N_5452,N_5200,N_5387);
xor U5453 (N_5453,N_5323,N_5297);
nand U5454 (N_5454,N_5311,N_5257);
xor U5455 (N_5455,N_5269,N_5290);
or U5456 (N_5456,N_5385,N_5364);
nor U5457 (N_5457,N_5282,N_5373);
xnor U5458 (N_5458,N_5213,N_5286);
xor U5459 (N_5459,N_5247,N_5378);
nor U5460 (N_5460,N_5321,N_5203);
nor U5461 (N_5461,N_5242,N_5299);
nand U5462 (N_5462,N_5239,N_5386);
or U5463 (N_5463,N_5259,N_5329);
or U5464 (N_5464,N_5368,N_5330);
or U5465 (N_5465,N_5394,N_5229);
nand U5466 (N_5466,N_5210,N_5201);
xor U5467 (N_5467,N_5353,N_5355);
or U5468 (N_5468,N_5391,N_5235);
nand U5469 (N_5469,N_5319,N_5208);
and U5470 (N_5470,N_5231,N_5226);
nand U5471 (N_5471,N_5296,N_5217);
nor U5472 (N_5472,N_5219,N_5396);
and U5473 (N_5473,N_5303,N_5384);
and U5474 (N_5474,N_5234,N_5285);
nand U5475 (N_5475,N_5305,N_5375);
or U5476 (N_5476,N_5211,N_5318);
xor U5477 (N_5477,N_5266,N_5312);
nand U5478 (N_5478,N_5338,N_5220);
nor U5479 (N_5479,N_5216,N_5246);
or U5480 (N_5480,N_5360,N_5370);
and U5481 (N_5481,N_5339,N_5341);
xor U5482 (N_5482,N_5212,N_5347);
and U5483 (N_5483,N_5227,N_5289);
nand U5484 (N_5484,N_5322,N_5271);
nand U5485 (N_5485,N_5240,N_5399);
nand U5486 (N_5486,N_5224,N_5326);
nor U5487 (N_5487,N_5366,N_5221);
and U5488 (N_5488,N_5317,N_5298);
and U5489 (N_5489,N_5288,N_5283);
or U5490 (N_5490,N_5265,N_5333);
nand U5491 (N_5491,N_5383,N_5254);
xnor U5492 (N_5492,N_5250,N_5272);
and U5493 (N_5493,N_5273,N_5260);
or U5494 (N_5494,N_5275,N_5263);
nand U5495 (N_5495,N_5301,N_5206);
and U5496 (N_5496,N_5248,N_5225);
xnor U5497 (N_5497,N_5348,N_5294);
and U5498 (N_5498,N_5359,N_5349);
nor U5499 (N_5499,N_5292,N_5252);
nor U5500 (N_5500,N_5225,N_5239);
nand U5501 (N_5501,N_5375,N_5391);
or U5502 (N_5502,N_5362,N_5394);
or U5503 (N_5503,N_5278,N_5336);
nor U5504 (N_5504,N_5269,N_5286);
xor U5505 (N_5505,N_5231,N_5388);
and U5506 (N_5506,N_5210,N_5249);
and U5507 (N_5507,N_5341,N_5297);
xnor U5508 (N_5508,N_5393,N_5302);
nor U5509 (N_5509,N_5287,N_5273);
or U5510 (N_5510,N_5389,N_5375);
and U5511 (N_5511,N_5381,N_5358);
nor U5512 (N_5512,N_5321,N_5283);
xor U5513 (N_5513,N_5291,N_5206);
and U5514 (N_5514,N_5398,N_5333);
and U5515 (N_5515,N_5359,N_5345);
xor U5516 (N_5516,N_5351,N_5315);
nor U5517 (N_5517,N_5307,N_5290);
or U5518 (N_5518,N_5200,N_5278);
and U5519 (N_5519,N_5316,N_5277);
and U5520 (N_5520,N_5209,N_5258);
or U5521 (N_5521,N_5234,N_5287);
nand U5522 (N_5522,N_5358,N_5294);
and U5523 (N_5523,N_5337,N_5209);
or U5524 (N_5524,N_5345,N_5227);
nand U5525 (N_5525,N_5210,N_5264);
nand U5526 (N_5526,N_5256,N_5327);
or U5527 (N_5527,N_5282,N_5269);
xor U5528 (N_5528,N_5350,N_5272);
xnor U5529 (N_5529,N_5311,N_5293);
nand U5530 (N_5530,N_5387,N_5275);
xnor U5531 (N_5531,N_5389,N_5202);
nand U5532 (N_5532,N_5253,N_5222);
nand U5533 (N_5533,N_5280,N_5213);
xnor U5534 (N_5534,N_5372,N_5285);
nand U5535 (N_5535,N_5228,N_5380);
or U5536 (N_5536,N_5306,N_5242);
nand U5537 (N_5537,N_5216,N_5341);
nand U5538 (N_5538,N_5334,N_5277);
nor U5539 (N_5539,N_5341,N_5257);
and U5540 (N_5540,N_5336,N_5350);
nand U5541 (N_5541,N_5231,N_5301);
xnor U5542 (N_5542,N_5308,N_5363);
xor U5543 (N_5543,N_5332,N_5387);
nor U5544 (N_5544,N_5321,N_5327);
and U5545 (N_5545,N_5275,N_5308);
nand U5546 (N_5546,N_5287,N_5251);
and U5547 (N_5547,N_5333,N_5295);
nor U5548 (N_5548,N_5328,N_5228);
nor U5549 (N_5549,N_5202,N_5356);
or U5550 (N_5550,N_5219,N_5378);
or U5551 (N_5551,N_5323,N_5349);
or U5552 (N_5552,N_5219,N_5338);
and U5553 (N_5553,N_5209,N_5342);
or U5554 (N_5554,N_5243,N_5269);
and U5555 (N_5555,N_5224,N_5208);
xor U5556 (N_5556,N_5325,N_5253);
and U5557 (N_5557,N_5248,N_5299);
nor U5558 (N_5558,N_5216,N_5362);
or U5559 (N_5559,N_5328,N_5279);
and U5560 (N_5560,N_5353,N_5359);
nor U5561 (N_5561,N_5307,N_5314);
and U5562 (N_5562,N_5272,N_5261);
or U5563 (N_5563,N_5295,N_5297);
nor U5564 (N_5564,N_5228,N_5338);
or U5565 (N_5565,N_5343,N_5267);
or U5566 (N_5566,N_5271,N_5236);
and U5567 (N_5567,N_5324,N_5318);
nand U5568 (N_5568,N_5310,N_5375);
nor U5569 (N_5569,N_5217,N_5300);
nand U5570 (N_5570,N_5350,N_5329);
nor U5571 (N_5571,N_5234,N_5237);
or U5572 (N_5572,N_5231,N_5200);
nand U5573 (N_5573,N_5233,N_5225);
or U5574 (N_5574,N_5323,N_5253);
or U5575 (N_5575,N_5266,N_5236);
or U5576 (N_5576,N_5364,N_5378);
or U5577 (N_5577,N_5359,N_5283);
nor U5578 (N_5578,N_5300,N_5321);
and U5579 (N_5579,N_5382,N_5304);
or U5580 (N_5580,N_5368,N_5247);
and U5581 (N_5581,N_5318,N_5206);
or U5582 (N_5582,N_5341,N_5239);
or U5583 (N_5583,N_5350,N_5392);
nor U5584 (N_5584,N_5337,N_5262);
or U5585 (N_5585,N_5252,N_5324);
and U5586 (N_5586,N_5342,N_5301);
nand U5587 (N_5587,N_5383,N_5270);
xor U5588 (N_5588,N_5266,N_5290);
or U5589 (N_5589,N_5364,N_5240);
nor U5590 (N_5590,N_5346,N_5349);
or U5591 (N_5591,N_5367,N_5303);
or U5592 (N_5592,N_5341,N_5264);
nor U5593 (N_5593,N_5343,N_5268);
xor U5594 (N_5594,N_5227,N_5319);
nor U5595 (N_5595,N_5219,N_5252);
or U5596 (N_5596,N_5329,N_5304);
nor U5597 (N_5597,N_5307,N_5213);
or U5598 (N_5598,N_5252,N_5243);
xor U5599 (N_5599,N_5254,N_5358);
xnor U5600 (N_5600,N_5511,N_5409);
xnor U5601 (N_5601,N_5540,N_5522);
or U5602 (N_5602,N_5500,N_5421);
or U5603 (N_5603,N_5476,N_5578);
nand U5604 (N_5604,N_5486,N_5449);
xor U5605 (N_5605,N_5422,N_5458);
and U5606 (N_5606,N_5544,N_5460);
or U5607 (N_5607,N_5520,N_5574);
and U5608 (N_5608,N_5594,N_5597);
nand U5609 (N_5609,N_5580,N_5525);
nand U5610 (N_5610,N_5526,N_5494);
or U5611 (N_5611,N_5450,N_5535);
or U5612 (N_5612,N_5541,N_5568);
or U5613 (N_5613,N_5531,N_5402);
or U5614 (N_5614,N_5404,N_5466);
nand U5615 (N_5615,N_5475,N_5400);
or U5616 (N_5616,N_5472,N_5576);
nand U5617 (N_5617,N_5566,N_5595);
xnor U5618 (N_5618,N_5425,N_5585);
or U5619 (N_5619,N_5579,N_5413);
or U5620 (N_5620,N_5459,N_5545);
nand U5621 (N_5621,N_5473,N_5438);
nor U5622 (N_5622,N_5447,N_5408);
xor U5623 (N_5623,N_5468,N_5599);
xor U5624 (N_5624,N_5453,N_5452);
nor U5625 (N_5625,N_5560,N_5434);
and U5626 (N_5626,N_5565,N_5529);
nor U5627 (N_5627,N_5489,N_5417);
or U5628 (N_5628,N_5441,N_5477);
or U5629 (N_5629,N_5528,N_5495);
nand U5630 (N_5630,N_5502,N_5546);
nor U5631 (N_5631,N_5598,N_5499);
or U5632 (N_5632,N_5589,N_5462);
nand U5633 (N_5633,N_5534,N_5573);
xnor U5634 (N_5634,N_5485,N_5401);
xor U5635 (N_5635,N_5474,N_5515);
nor U5636 (N_5636,N_5406,N_5551);
xnor U5637 (N_5637,N_5439,N_5581);
nand U5638 (N_5638,N_5420,N_5550);
nor U5639 (N_5639,N_5547,N_5442);
and U5640 (N_5640,N_5443,N_5479);
xnor U5641 (N_5641,N_5465,N_5538);
and U5642 (N_5642,N_5505,N_5507);
nor U5643 (N_5643,N_5510,N_5567);
nor U5644 (N_5644,N_5457,N_5497);
or U5645 (N_5645,N_5569,N_5419);
nand U5646 (N_5646,N_5533,N_5501);
nor U5647 (N_5647,N_5558,N_5537);
xnor U5648 (N_5648,N_5521,N_5467);
or U5649 (N_5649,N_5509,N_5590);
nor U5650 (N_5650,N_5418,N_5432);
and U5651 (N_5651,N_5436,N_5410);
nor U5652 (N_5652,N_5414,N_5480);
or U5653 (N_5653,N_5423,N_5490);
nand U5654 (N_5654,N_5571,N_5557);
nand U5655 (N_5655,N_5559,N_5464);
and U5656 (N_5656,N_5548,N_5433);
or U5657 (N_5657,N_5487,N_5416);
nand U5658 (N_5658,N_5426,N_5491);
or U5659 (N_5659,N_5575,N_5517);
xor U5660 (N_5660,N_5539,N_5563);
or U5661 (N_5661,N_5481,N_5455);
and U5662 (N_5662,N_5508,N_5478);
or U5663 (N_5663,N_5556,N_5445);
nand U5664 (N_5664,N_5428,N_5483);
nor U5665 (N_5665,N_5593,N_5542);
nor U5666 (N_5666,N_5446,N_5424);
or U5667 (N_5667,N_5584,N_5572);
or U5668 (N_5668,N_5403,N_5412);
xnor U5669 (N_5669,N_5577,N_5407);
xnor U5670 (N_5670,N_5549,N_5555);
and U5671 (N_5671,N_5504,N_5519);
nor U5672 (N_5672,N_5586,N_5469);
nand U5673 (N_5673,N_5461,N_5543);
nor U5674 (N_5674,N_5503,N_5587);
nand U5675 (N_5675,N_5513,N_5553);
nor U5676 (N_5676,N_5518,N_5440);
nand U5677 (N_5677,N_5470,N_5411);
and U5678 (N_5678,N_5431,N_5583);
xnor U5679 (N_5679,N_5484,N_5454);
or U5680 (N_5680,N_5523,N_5493);
or U5681 (N_5681,N_5444,N_5592);
or U5682 (N_5682,N_5427,N_5536);
or U5683 (N_5683,N_5488,N_5512);
and U5684 (N_5684,N_5532,N_5562);
and U5685 (N_5685,N_5561,N_5514);
or U5686 (N_5686,N_5492,N_5471);
nand U5687 (N_5687,N_5430,N_5451);
nand U5688 (N_5688,N_5516,N_5448);
xor U5689 (N_5689,N_5588,N_5435);
nor U5690 (N_5690,N_5524,N_5554);
xnor U5691 (N_5691,N_5415,N_5463);
or U5692 (N_5692,N_5482,N_5429);
or U5693 (N_5693,N_5496,N_5498);
xor U5694 (N_5694,N_5564,N_5582);
nor U5695 (N_5695,N_5405,N_5456);
xor U5696 (N_5696,N_5437,N_5530);
nand U5697 (N_5697,N_5591,N_5552);
and U5698 (N_5698,N_5596,N_5506);
or U5699 (N_5699,N_5527,N_5570);
or U5700 (N_5700,N_5585,N_5482);
nand U5701 (N_5701,N_5435,N_5546);
xnor U5702 (N_5702,N_5596,N_5410);
nor U5703 (N_5703,N_5514,N_5460);
nor U5704 (N_5704,N_5592,N_5482);
or U5705 (N_5705,N_5480,N_5536);
nor U5706 (N_5706,N_5448,N_5472);
nor U5707 (N_5707,N_5431,N_5469);
or U5708 (N_5708,N_5483,N_5408);
xor U5709 (N_5709,N_5426,N_5434);
nand U5710 (N_5710,N_5461,N_5410);
or U5711 (N_5711,N_5491,N_5524);
nor U5712 (N_5712,N_5577,N_5557);
xor U5713 (N_5713,N_5533,N_5549);
and U5714 (N_5714,N_5497,N_5450);
nor U5715 (N_5715,N_5584,N_5503);
nor U5716 (N_5716,N_5541,N_5534);
nand U5717 (N_5717,N_5490,N_5591);
and U5718 (N_5718,N_5467,N_5581);
nor U5719 (N_5719,N_5526,N_5438);
nor U5720 (N_5720,N_5412,N_5491);
nor U5721 (N_5721,N_5569,N_5467);
nor U5722 (N_5722,N_5409,N_5517);
or U5723 (N_5723,N_5583,N_5476);
nand U5724 (N_5724,N_5550,N_5465);
xor U5725 (N_5725,N_5473,N_5508);
nor U5726 (N_5726,N_5549,N_5498);
or U5727 (N_5727,N_5420,N_5424);
and U5728 (N_5728,N_5454,N_5566);
and U5729 (N_5729,N_5481,N_5555);
nand U5730 (N_5730,N_5590,N_5558);
or U5731 (N_5731,N_5469,N_5549);
nand U5732 (N_5732,N_5514,N_5458);
nor U5733 (N_5733,N_5463,N_5529);
nand U5734 (N_5734,N_5524,N_5427);
or U5735 (N_5735,N_5468,N_5459);
or U5736 (N_5736,N_5468,N_5504);
nand U5737 (N_5737,N_5539,N_5568);
and U5738 (N_5738,N_5555,N_5514);
or U5739 (N_5739,N_5560,N_5557);
xnor U5740 (N_5740,N_5532,N_5513);
or U5741 (N_5741,N_5447,N_5455);
xnor U5742 (N_5742,N_5459,N_5500);
and U5743 (N_5743,N_5585,N_5481);
or U5744 (N_5744,N_5543,N_5439);
and U5745 (N_5745,N_5487,N_5523);
nand U5746 (N_5746,N_5495,N_5455);
nor U5747 (N_5747,N_5478,N_5459);
and U5748 (N_5748,N_5519,N_5527);
and U5749 (N_5749,N_5453,N_5414);
nor U5750 (N_5750,N_5500,N_5559);
xnor U5751 (N_5751,N_5598,N_5453);
or U5752 (N_5752,N_5573,N_5591);
nor U5753 (N_5753,N_5547,N_5556);
and U5754 (N_5754,N_5408,N_5471);
nor U5755 (N_5755,N_5511,N_5462);
and U5756 (N_5756,N_5504,N_5514);
nand U5757 (N_5757,N_5494,N_5556);
or U5758 (N_5758,N_5481,N_5432);
xor U5759 (N_5759,N_5565,N_5590);
nand U5760 (N_5760,N_5524,N_5590);
or U5761 (N_5761,N_5502,N_5570);
xor U5762 (N_5762,N_5409,N_5578);
and U5763 (N_5763,N_5563,N_5556);
xor U5764 (N_5764,N_5554,N_5505);
and U5765 (N_5765,N_5405,N_5487);
nand U5766 (N_5766,N_5470,N_5498);
or U5767 (N_5767,N_5483,N_5574);
xor U5768 (N_5768,N_5543,N_5421);
xor U5769 (N_5769,N_5450,N_5540);
or U5770 (N_5770,N_5537,N_5462);
xor U5771 (N_5771,N_5542,N_5487);
xnor U5772 (N_5772,N_5405,N_5426);
nand U5773 (N_5773,N_5597,N_5579);
xor U5774 (N_5774,N_5434,N_5470);
and U5775 (N_5775,N_5515,N_5527);
nand U5776 (N_5776,N_5555,N_5451);
or U5777 (N_5777,N_5488,N_5477);
nand U5778 (N_5778,N_5450,N_5445);
and U5779 (N_5779,N_5511,N_5432);
nand U5780 (N_5780,N_5425,N_5519);
or U5781 (N_5781,N_5513,N_5575);
nor U5782 (N_5782,N_5493,N_5542);
xor U5783 (N_5783,N_5538,N_5560);
or U5784 (N_5784,N_5579,N_5440);
xor U5785 (N_5785,N_5446,N_5581);
or U5786 (N_5786,N_5500,N_5430);
or U5787 (N_5787,N_5509,N_5550);
xnor U5788 (N_5788,N_5412,N_5557);
xor U5789 (N_5789,N_5542,N_5427);
or U5790 (N_5790,N_5505,N_5464);
or U5791 (N_5791,N_5510,N_5462);
or U5792 (N_5792,N_5572,N_5526);
xnor U5793 (N_5793,N_5494,N_5410);
or U5794 (N_5794,N_5437,N_5462);
nor U5795 (N_5795,N_5469,N_5485);
xnor U5796 (N_5796,N_5480,N_5404);
nor U5797 (N_5797,N_5575,N_5579);
and U5798 (N_5798,N_5471,N_5533);
nor U5799 (N_5799,N_5435,N_5570);
nand U5800 (N_5800,N_5660,N_5785);
and U5801 (N_5801,N_5606,N_5680);
and U5802 (N_5802,N_5604,N_5796);
nor U5803 (N_5803,N_5645,N_5757);
and U5804 (N_5804,N_5664,N_5745);
nor U5805 (N_5805,N_5706,N_5779);
xor U5806 (N_5806,N_5666,N_5612);
nor U5807 (N_5807,N_5759,N_5635);
and U5808 (N_5808,N_5696,N_5717);
and U5809 (N_5809,N_5633,N_5682);
or U5810 (N_5810,N_5691,N_5636);
xnor U5811 (N_5811,N_5624,N_5668);
nand U5812 (N_5812,N_5653,N_5637);
or U5813 (N_5813,N_5610,N_5767);
nand U5814 (N_5814,N_5685,N_5716);
nand U5815 (N_5815,N_5616,N_5721);
or U5816 (N_5816,N_5790,N_5791);
xnor U5817 (N_5817,N_5750,N_5792);
or U5818 (N_5818,N_5763,N_5688);
nor U5819 (N_5819,N_5741,N_5742);
nand U5820 (N_5820,N_5772,N_5657);
xnor U5821 (N_5821,N_5622,N_5619);
nor U5822 (N_5822,N_5708,N_5778);
nand U5823 (N_5823,N_5651,N_5683);
and U5824 (N_5824,N_5747,N_5630);
or U5825 (N_5825,N_5729,N_5638);
nor U5826 (N_5826,N_5611,N_5614);
xnor U5827 (N_5827,N_5697,N_5629);
and U5828 (N_5828,N_5758,N_5781);
nand U5829 (N_5829,N_5655,N_5711);
or U5830 (N_5830,N_5658,N_5665);
or U5831 (N_5831,N_5786,N_5615);
nand U5832 (N_5832,N_5783,N_5765);
or U5833 (N_5833,N_5602,N_5672);
and U5834 (N_5834,N_5601,N_5631);
nor U5835 (N_5835,N_5648,N_5733);
xor U5836 (N_5836,N_5746,N_5650);
and U5837 (N_5837,N_5709,N_5764);
xnor U5838 (N_5838,N_5752,N_5663);
xor U5839 (N_5839,N_5620,N_5656);
nor U5840 (N_5840,N_5674,N_5659);
or U5841 (N_5841,N_5724,N_5609);
nor U5842 (N_5842,N_5773,N_5710);
nor U5843 (N_5843,N_5699,N_5693);
nor U5844 (N_5844,N_5797,N_5727);
nand U5845 (N_5845,N_5705,N_5755);
xnor U5846 (N_5846,N_5760,N_5689);
nor U5847 (N_5847,N_5669,N_5723);
or U5848 (N_5848,N_5702,N_5725);
and U5849 (N_5849,N_5799,N_5769);
nand U5850 (N_5850,N_5780,N_5798);
or U5851 (N_5851,N_5632,N_5627);
nor U5852 (N_5852,N_5670,N_5738);
xnor U5853 (N_5853,N_5737,N_5644);
and U5854 (N_5854,N_5639,N_5618);
nand U5855 (N_5855,N_5684,N_5646);
xor U5856 (N_5856,N_5628,N_5679);
nand U5857 (N_5857,N_5613,N_5695);
and U5858 (N_5858,N_5740,N_5603);
and U5859 (N_5859,N_5777,N_5782);
or U5860 (N_5860,N_5720,N_5681);
xor U5861 (N_5861,N_5718,N_5643);
and U5862 (N_5862,N_5676,N_5704);
nand U5863 (N_5863,N_5735,N_5625);
or U5864 (N_5864,N_5748,N_5605);
and U5865 (N_5865,N_5623,N_5712);
nor U5866 (N_5866,N_5607,N_5686);
nand U5867 (N_5867,N_5774,N_5793);
nor U5868 (N_5868,N_5621,N_5701);
nor U5869 (N_5869,N_5756,N_5739);
nand U5870 (N_5870,N_5687,N_5776);
and U5871 (N_5871,N_5673,N_5743);
nor U5872 (N_5872,N_5654,N_5730);
nand U5873 (N_5873,N_5749,N_5707);
nand U5874 (N_5874,N_5634,N_5784);
nor U5875 (N_5875,N_5794,N_5649);
and U5876 (N_5876,N_5734,N_5694);
nand U5877 (N_5877,N_5652,N_5640);
nor U5878 (N_5878,N_5715,N_5736);
and U5879 (N_5879,N_5667,N_5642);
nand U5880 (N_5880,N_5771,N_5700);
and U5881 (N_5881,N_5671,N_5719);
and U5882 (N_5882,N_5795,N_5690);
or U5883 (N_5883,N_5766,N_5761);
nand U5884 (N_5884,N_5661,N_5641);
and U5885 (N_5885,N_5714,N_5626);
and U5886 (N_5886,N_5617,N_5726);
xor U5887 (N_5887,N_5703,N_5744);
xnor U5888 (N_5888,N_5722,N_5662);
or U5889 (N_5889,N_5787,N_5788);
xor U5890 (N_5890,N_5732,N_5675);
nor U5891 (N_5891,N_5762,N_5751);
or U5892 (N_5892,N_5775,N_5600);
and U5893 (N_5893,N_5728,N_5647);
nand U5894 (N_5894,N_5768,N_5754);
xnor U5895 (N_5895,N_5713,N_5608);
xnor U5896 (N_5896,N_5692,N_5789);
xnor U5897 (N_5897,N_5770,N_5677);
xnor U5898 (N_5898,N_5698,N_5731);
and U5899 (N_5899,N_5753,N_5678);
nor U5900 (N_5900,N_5705,N_5737);
nor U5901 (N_5901,N_5695,N_5793);
xor U5902 (N_5902,N_5709,N_5673);
nor U5903 (N_5903,N_5653,N_5649);
xor U5904 (N_5904,N_5617,N_5635);
and U5905 (N_5905,N_5769,N_5688);
nor U5906 (N_5906,N_5674,N_5797);
nor U5907 (N_5907,N_5773,N_5671);
xnor U5908 (N_5908,N_5709,N_5632);
xnor U5909 (N_5909,N_5686,N_5788);
nand U5910 (N_5910,N_5760,N_5604);
nor U5911 (N_5911,N_5732,N_5726);
nand U5912 (N_5912,N_5614,N_5773);
nand U5913 (N_5913,N_5657,N_5661);
nand U5914 (N_5914,N_5789,N_5761);
xnor U5915 (N_5915,N_5621,N_5770);
and U5916 (N_5916,N_5623,N_5653);
and U5917 (N_5917,N_5697,N_5777);
nor U5918 (N_5918,N_5643,N_5687);
nor U5919 (N_5919,N_5601,N_5753);
nand U5920 (N_5920,N_5738,N_5731);
or U5921 (N_5921,N_5796,N_5643);
nand U5922 (N_5922,N_5778,N_5799);
nand U5923 (N_5923,N_5770,N_5706);
nor U5924 (N_5924,N_5725,N_5790);
nor U5925 (N_5925,N_5693,N_5719);
xnor U5926 (N_5926,N_5621,N_5709);
nor U5927 (N_5927,N_5683,N_5616);
or U5928 (N_5928,N_5668,N_5777);
xor U5929 (N_5929,N_5700,N_5645);
xor U5930 (N_5930,N_5714,N_5615);
and U5931 (N_5931,N_5722,N_5690);
or U5932 (N_5932,N_5796,N_5779);
and U5933 (N_5933,N_5721,N_5712);
and U5934 (N_5934,N_5764,N_5797);
and U5935 (N_5935,N_5633,N_5731);
and U5936 (N_5936,N_5706,N_5701);
nand U5937 (N_5937,N_5696,N_5737);
or U5938 (N_5938,N_5784,N_5798);
nand U5939 (N_5939,N_5761,N_5606);
and U5940 (N_5940,N_5663,N_5703);
xnor U5941 (N_5941,N_5717,N_5799);
nand U5942 (N_5942,N_5678,N_5714);
nand U5943 (N_5943,N_5667,N_5665);
or U5944 (N_5944,N_5790,N_5792);
nor U5945 (N_5945,N_5732,N_5733);
and U5946 (N_5946,N_5684,N_5769);
and U5947 (N_5947,N_5689,N_5647);
nor U5948 (N_5948,N_5615,N_5664);
nand U5949 (N_5949,N_5739,N_5742);
xnor U5950 (N_5950,N_5655,N_5772);
xor U5951 (N_5951,N_5732,N_5697);
nand U5952 (N_5952,N_5655,N_5620);
xor U5953 (N_5953,N_5688,N_5706);
xor U5954 (N_5954,N_5675,N_5699);
xnor U5955 (N_5955,N_5724,N_5637);
and U5956 (N_5956,N_5785,N_5727);
nor U5957 (N_5957,N_5772,N_5716);
or U5958 (N_5958,N_5772,N_5753);
xnor U5959 (N_5959,N_5691,N_5649);
and U5960 (N_5960,N_5650,N_5778);
and U5961 (N_5961,N_5619,N_5627);
xnor U5962 (N_5962,N_5761,N_5738);
nand U5963 (N_5963,N_5703,N_5636);
xnor U5964 (N_5964,N_5652,N_5780);
nand U5965 (N_5965,N_5679,N_5688);
nand U5966 (N_5966,N_5769,N_5645);
nand U5967 (N_5967,N_5794,N_5712);
or U5968 (N_5968,N_5689,N_5612);
or U5969 (N_5969,N_5752,N_5657);
xnor U5970 (N_5970,N_5773,N_5652);
or U5971 (N_5971,N_5770,N_5740);
xnor U5972 (N_5972,N_5691,N_5743);
and U5973 (N_5973,N_5650,N_5769);
nand U5974 (N_5974,N_5704,N_5771);
nand U5975 (N_5975,N_5771,N_5604);
nor U5976 (N_5976,N_5764,N_5710);
nand U5977 (N_5977,N_5648,N_5693);
nor U5978 (N_5978,N_5766,N_5607);
or U5979 (N_5979,N_5741,N_5634);
nand U5980 (N_5980,N_5726,N_5779);
nand U5981 (N_5981,N_5792,N_5675);
nor U5982 (N_5982,N_5764,N_5796);
nor U5983 (N_5983,N_5632,N_5752);
or U5984 (N_5984,N_5723,N_5620);
or U5985 (N_5985,N_5633,N_5790);
and U5986 (N_5986,N_5631,N_5648);
xnor U5987 (N_5987,N_5639,N_5660);
and U5988 (N_5988,N_5727,N_5668);
nor U5989 (N_5989,N_5721,N_5620);
and U5990 (N_5990,N_5643,N_5764);
or U5991 (N_5991,N_5710,N_5787);
nand U5992 (N_5992,N_5609,N_5753);
xnor U5993 (N_5993,N_5605,N_5640);
and U5994 (N_5994,N_5654,N_5612);
nor U5995 (N_5995,N_5741,N_5684);
or U5996 (N_5996,N_5619,N_5693);
nand U5997 (N_5997,N_5636,N_5692);
nand U5998 (N_5998,N_5791,N_5641);
nor U5999 (N_5999,N_5640,N_5745);
and U6000 (N_6000,N_5866,N_5936);
nand U6001 (N_6001,N_5868,N_5885);
and U6002 (N_6002,N_5810,N_5935);
xnor U6003 (N_6003,N_5800,N_5846);
and U6004 (N_6004,N_5921,N_5830);
nor U6005 (N_6005,N_5979,N_5916);
nand U6006 (N_6006,N_5961,N_5833);
nor U6007 (N_6007,N_5822,N_5896);
nor U6008 (N_6008,N_5886,N_5985);
or U6009 (N_6009,N_5827,N_5906);
or U6010 (N_6010,N_5869,N_5857);
nor U6011 (N_6011,N_5843,N_5972);
and U6012 (N_6012,N_5995,N_5853);
or U6013 (N_6013,N_5953,N_5944);
and U6014 (N_6014,N_5820,N_5958);
or U6015 (N_6015,N_5839,N_5941);
xor U6016 (N_6016,N_5887,N_5975);
nand U6017 (N_6017,N_5879,N_5855);
and U6018 (N_6018,N_5931,N_5809);
and U6019 (N_6019,N_5912,N_5952);
and U6020 (N_6020,N_5997,N_5837);
nor U6021 (N_6021,N_5851,N_5890);
and U6022 (N_6022,N_5844,N_5957);
or U6023 (N_6023,N_5899,N_5905);
and U6024 (N_6024,N_5946,N_5978);
nand U6025 (N_6025,N_5963,N_5920);
or U6026 (N_6026,N_5836,N_5804);
xor U6027 (N_6027,N_5854,N_5956);
or U6028 (N_6028,N_5864,N_5924);
nand U6029 (N_6029,N_5955,N_5973);
nor U6030 (N_6030,N_5852,N_5909);
nand U6031 (N_6031,N_5917,N_5913);
and U6032 (N_6032,N_5976,N_5943);
nand U6033 (N_6033,N_5966,N_5823);
and U6034 (N_6034,N_5949,N_5863);
and U6035 (N_6035,N_5834,N_5938);
nor U6036 (N_6036,N_5841,N_5805);
nor U6037 (N_6037,N_5821,N_5932);
and U6038 (N_6038,N_5945,N_5968);
or U6039 (N_6039,N_5950,N_5872);
or U6040 (N_6040,N_5951,N_5914);
nand U6041 (N_6041,N_5962,N_5990);
xnor U6042 (N_6042,N_5933,N_5895);
and U6043 (N_6043,N_5897,N_5986);
or U6044 (N_6044,N_5954,N_5867);
or U6045 (N_6045,N_5981,N_5816);
and U6046 (N_6046,N_5988,N_5918);
nor U6047 (N_6047,N_5904,N_5992);
and U6048 (N_6048,N_5859,N_5898);
xor U6049 (N_6049,N_5892,N_5911);
and U6050 (N_6050,N_5835,N_5860);
nor U6051 (N_6051,N_5888,N_5807);
and U6052 (N_6052,N_5808,N_5960);
and U6053 (N_6053,N_5881,N_5965);
or U6054 (N_6054,N_5993,N_5891);
nor U6055 (N_6055,N_5883,N_5828);
nor U6056 (N_6056,N_5824,N_5934);
and U6057 (N_6057,N_5803,N_5873);
and U6058 (N_6058,N_5877,N_5937);
nand U6059 (N_6059,N_5858,N_5996);
xnor U6060 (N_6060,N_5959,N_5889);
nor U6061 (N_6061,N_5984,N_5999);
xor U6062 (N_6062,N_5806,N_5825);
nor U6063 (N_6063,N_5901,N_5910);
nand U6064 (N_6064,N_5818,N_5819);
nand U6065 (N_6065,N_5919,N_5940);
nand U6066 (N_6066,N_5974,N_5838);
xnor U6067 (N_6067,N_5967,N_5903);
nand U6068 (N_6068,N_5811,N_5876);
and U6069 (N_6069,N_5871,N_5849);
xor U6070 (N_6070,N_5894,N_5878);
or U6071 (N_6071,N_5964,N_5925);
nor U6072 (N_6072,N_5870,N_5862);
or U6073 (N_6073,N_5927,N_5942);
or U6074 (N_6074,N_5907,N_5845);
and U6075 (N_6075,N_5948,N_5882);
and U6076 (N_6076,N_5893,N_5832);
nand U6077 (N_6077,N_5982,N_5848);
nand U6078 (N_6078,N_5826,N_5801);
nor U6079 (N_6079,N_5861,N_5969);
nand U6080 (N_6080,N_5929,N_5875);
xnor U6081 (N_6081,N_5998,N_5850);
xnor U6082 (N_6082,N_5884,N_5829);
xnor U6083 (N_6083,N_5831,N_5814);
xor U6084 (N_6084,N_5812,N_5880);
and U6085 (N_6085,N_5926,N_5915);
xor U6086 (N_6086,N_5970,N_5922);
nand U6087 (N_6087,N_5815,N_5802);
or U6088 (N_6088,N_5840,N_5865);
and U6089 (N_6089,N_5856,N_5947);
nand U6090 (N_6090,N_5971,N_5939);
nor U6091 (N_6091,N_5923,N_5813);
nor U6092 (N_6092,N_5983,N_5874);
nand U6093 (N_6093,N_5842,N_5989);
and U6094 (N_6094,N_5930,N_5977);
nor U6095 (N_6095,N_5928,N_5817);
and U6096 (N_6096,N_5987,N_5902);
nor U6097 (N_6097,N_5908,N_5847);
nor U6098 (N_6098,N_5900,N_5994);
nor U6099 (N_6099,N_5980,N_5991);
or U6100 (N_6100,N_5894,N_5992);
or U6101 (N_6101,N_5856,N_5874);
xor U6102 (N_6102,N_5997,N_5926);
xnor U6103 (N_6103,N_5824,N_5974);
or U6104 (N_6104,N_5890,N_5926);
or U6105 (N_6105,N_5975,N_5889);
nor U6106 (N_6106,N_5867,N_5881);
nor U6107 (N_6107,N_5894,N_5952);
and U6108 (N_6108,N_5851,N_5887);
nor U6109 (N_6109,N_5889,N_5966);
and U6110 (N_6110,N_5846,N_5985);
nand U6111 (N_6111,N_5996,N_5997);
xnor U6112 (N_6112,N_5858,N_5816);
xor U6113 (N_6113,N_5939,N_5933);
or U6114 (N_6114,N_5868,N_5956);
nand U6115 (N_6115,N_5903,N_5973);
nor U6116 (N_6116,N_5981,N_5813);
or U6117 (N_6117,N_5926,N_5977);
or U6118 (N_6118,N_5801,N_5992);
nor U6119 (N_6119,N_5869,N_5999);
nand U6120 (N_6120,N_5966,N_5949);
xnor U6121 (N_6121,N_5921,N_5820);
nor U6122 (N_6122,N_5823,N_5890);
or U6123 (N_6123,N_5926,N_5858);
nor U6124 (N_6124,N_5961,N_5972);
or U6125 (N_6125,N_5961,N_5990);
and U6126 (N_6126,N_5804,N_5979);
nor U6127 (N_6127,N_5881,N_5895);
or U6128 (N_6128,N_5836,N_5841);
nor U6129 (N_6129,N_5858,N_5951);
and U6130 (N_6130,N_5983,N_5842);
nor U6131 (N_6131,N_5892,N_5870);
nor U6132 (N_6132,N_5875,N_5848);
nand U6133 (N_6133,N_5954,N_5840);
nand U6134 (N_6134,N_5811,N_5975);
nor U6135 (N_6135,N_5824,N_5995);
and U6136 (N_6136,N_5922,N_5866);
or U6137 (N_6137,N_5989,N_5984);
or U6138 (N_6138,N_5867,N_5828);
and U6139 (N_6139,N_5941,N_5922);
or U6140 (N_6140,N_5887,N_5870);
or U6141 (N_6141,N_5913,N_5841);
or U6142 (N_6142,N_5915,N_5930);
nand U6143 (N_6143,N_5811,N_5813);
and U6144 (N_6144,N_5923,N_5826);
or U6145 (N_6145,N_5935,N_5856);
and U6146 (N_6146,N_5833,N_5861);
nand U6147 (N_6147,N_5835,N_5842);
or U6148 (N_6148,N_5850,N_5986);
nand U6149 (N_6149,N_5810,N_5804);
and U6150 (N_6150,N_5982,N_5950);
or U6151 (N_6151,N_5976,N_5841);
nand U6152 (N_6152,N_5876,N_5960);
and U6153 (N_6153,N_5983,N_5860);
nor U6154 (N_6154,N_5817,N_5807);
or U6155 (N_6155,N_5842,N_5893);
nor U6156 (N_6156,N_5884,N_5874);
xor U6157 (N_6157,N_5883,N_5988);
or U6158 (N_6158,N_5910,N_5919);
xor U6159 (N_6159,N_5815,N_5829);
xor U6160 (N_6160,N_5961,N_5963);
nand U6161 (N_6161,N_5820,N_5818);
nand U6162 (N_6162,N_5925,N_5894);
nor U6163 (N_6163,N_5804,N_5988);
or U6164 (N_6164,N_5838,N_5836);
nor U6165 (N_6165,N_5838,N_5845);
and U6166 (N_6166,N_5945,N_5805);
and U6167 (N_6167,N_5839,N_5975);
nor U6168 (N_6168,N_5901,N_5900);
xor U6169 (N_6169,N_5848,N_5836);
xor U6170 (N_6170,N_5841,N_5940);
or U6171 (N_6171,N_5802,N_5866);
and U6172 (N_6172,N_5898,N_5808);
or U6173 (N_6173,N_5800,N_5826);
xor U6174 (N_6174,N_5871,N_5910);
and U6175 (N_6175,N_5862,N_5976);
xor U6176 (N_6176,N_5928,N_5978);
nor U6177 (N_6177,N_5926,N_5827);
nand U6178 (N_6178,N_5913,N_5991);
or U6179 (N_6179,N_5977,N_5830);
nand U6180 (N_6180,N_5969,N_5876);
nor U6181 (N_6181,N_5852,N_5928);
xor U6182 (N_6182,N_5945,N_5914);
nand U6183 (N_6183,N_5872,N_5916);
nand U6184 (N_6184,N_5944,N_5864);
nand U6185 (N_6185,N_5804,N_5954);
nor U6186 (N_6186,N_5834,N_5845);
nor U6187 (N_6187,N_5964,N_5911);
or U6188 (N_6188,N_5950,N_5887);
nand U6189 (N_6189,N_5888,N_5914);
nor U6190 (N_6190,N_5929,N_5855);
nor U6191 (N_6191,N_5857,N_5893);
and U6192 (N_6192,N_5931,N_5997);
xnor U6193 (N_6193,N_5838,N_5898);
and U6194 (N_6194,N_5867,N_5873);
nand U6195 (N_6195,N_5907,N_5838);
xnor U6196 (N_6196,N_5884,N_5894);
nor U6197 (N_6197,N_5981,N_5837);
nor U6198 (N_6198,N_5848,N_5890);
or U6199 (N_6199,N_5841,N_5804);
or U6200 (N_6200,N_6009,N_6148);
or U6201 (N_6201,N_6059,N_6118);
nand U6202 (N_6202,N_6157,N_6172);
and U6203 (N_6203,N_6089,N_6036);
nor U6204 (N_6204,N_6188,N_6198);
nand U6205 (N_6205,N_6095,N_6136);
nor U6206 (N_6206,N_6022,N_6049);
or U6207 (N_6207,N_6086,N_6011);
nor U6208 (N_6208,N_6031,N_6184);
nand U6209 (N_6209,N_6017,N_6038);
xor U6210 (N_6210,N_6150,N_6028);
or U6211 (N_6211,N_6080,N_6063);
xor U6212 (N_6212,N_6025,N_6064);
nor U6213 (N_6213,N_6012,N_6046);
or U6214 (N_6214,N_6173,N_6152);
and U6215 (N_6215,N_6085,N_6183);
and U6216 (N_6216,N_6195,N_6190);
xnor U6217 (N_6217,N_6193,N_6196);
nand U6218 (N_6218,N_6001,N_6083);
nor U6219 (N_6219,N_6032,N_6014);
nand U6220 (N_6220,N_6051,N_6103);
or U6221 (N_6221,N_6078,N_6033);
nand U6222 (N_6222,N_6174,N_6069);
nor U6223 (N_6223,N_6087,N_6181);
or U6224 (N_6224,N_6013,N_6048);
nor U6225 (N_6225,N_6029,N_6062);
nor U6226 (N_6226,N_6004,N_6113);
nand U6227 (N_6227,N_6115,N_6096);
or U6228 (N_6228,N_6018,N_6159);
or U6229 (N_6229,N_6101,N_6041);
and U6230 (N_6230,N_6000,N_6125);
nor U6231 (N_6231,N_6026,N_6002);
and U6232 (N_6232,N_6139,N_6177);
and U6233 (N_6233,N_6175,N_6132);
and U6234 (N_6234,N_6109,N_6197);
and U6235 (N_6235,N_6058,N_6108);
xnor U6236 (N_6236,N_6137,N_6146);
xor U6237 (N_6237,N_6072,N_6077);
and U6238 (N_6238,N_6194,N_6191);
xnor U6239 (N_6239,N_6044,N_6135);
xor U6240 (N_6240,N_6156,N_6007);
nand U6241 (N_6241,N_6057,N_6145);
nand U6242 (N_6242,N_6182,N_6006);
nand U6243 (N_6243,N_6093,N_6106);
and U6244 (N_6244,N_6088,N_6158);
or U6245 (N_6245,N_6043,N_6116);
nor U6246 (N_6246,N_6040,N_6008);
nand U6247 (N_6247,N_6039,N_6075);
xnor U6248 (N_6248,N_6161,N_6005);
and U6249 (N_6249,N_6126,N_6168);
nand U6250 (N_6250,N_6164,N_6024);
or U6251 (N_6251,N_6073,N_6171);
nor U6252 (N_6252,N_6037,N_6060);
and U6253 (N_6253,N_6144,N_6084);
or U6254 (N_6254,N_6104,N_6045);
or U6255 (N_6255,N_6147,N_6098);
nand U6256 (N_6256,N_6153,N_6052);
nor U6257 (N_6257,N_6128,N_6129);
nand U6258 (N_6258,N_6185,N_6023);
nor U6259 (N_6259,N_6133,N_6124);
or U6260 (N_6260,N_6030,N_6019);
xor U6261 (N_6261,N_6092,N_6079);
nor U6262 (N_6262,N_6163,N_6111);
and U6263 (N_6263,N_6169,N_6071);
xor U6264 (N_6264,N_6143,N_6070);
nor U6265 (N_6265,N_6138,N_6081);
and U6266 (N_6266,N_6020,N_6076);
and U6267 (N_6267,N_6107,N_6015);
nand U6268 (N_6268,N_6053,N_6054);
xor U6269 (N_6269,N_6091,N_6162);
xnor U6270 (N_6270,N_6149,N_6021);
nand U6271 (N_6271,N_6186,N_6056);
or U6272 (N_6272,N_6121,N_6068);
nand U6273 (N_6273,N_6141,N_6154);
nand U6274 (N_6274,N_6035,N_6155);
and U6275 (N_6275,N_6122,N_6114);
or U6276 (N_6276,N_6055,N_6074);
nand U6277 (N_6277,N_6027,N_6067);
or U6278 (N_6278,N_6166,N_6102);
or U6279 (N_6279,N_6120,N_6066);
nand U6280 (N_6280,N_6176,N_6189);
and U6281 (N_6281,N_6016,N_6105);
or U6282 (N_6282,N_6142,N_6127);
or U6283 (N_6283,N_6160,N_6010);
xnor U6284 (N_6284,N_6131,N_6140);
and U6285 (N_6285,N_6061,N_6034);
and U6286 (N_6286,N_6042,N_6099);
or U6287 (N_6287,N_6178,N_6165);
xor U6288 (N_6288,N_6170,N_6151);
and U6289 (N_6289,N_6090,N_6065);
and U6290 (N_6290,N_6082,N_6050);
nor U6291 (N_6291,N_6123,N_6199);
xnor U6292 (N_6292,N_6047,N_6119);
nand U6293 (N_6293,N_6130,N_6180);
and U6294 (N_6294,N_6094,N_6110);
nor U6295 (N_6295,N_6179,N_6100);
or U6296 (N_6296,N_6192,N_6117);
xor U6297 (N_6297,N_6187,N_6112);
and U6298 (N_6298,N_6134,N_6167);
xnor U6299 (N_6299,N_6003,N_6097);
and U6300 (N_6300,N_6188,N_6076);
nor U6301 (N_6301,N_6055,N_6195);
or U6302 (N_6302,N_6143,N_6153);
xnor U6303 (N_6303,N_6139,N_6071);
or U6304 (N_6304,N_6025,N_6081);
and U6305 (N_6305,N_6128,N_6018);
nand U6306 (N_6306,N_6112,N_6102);
xnor U6307 (N_6307,N_6004,N_6096);
nor U6308 (N_6308,N_6056,N_6184);
nor U6309 (N_6309,N_6130,N_6138);
and U6310 (N_6310,N_6138,N_6116);
nand U6311 (N_6311,N_6127,N_6147);
xor U6312 (N_6312,N_6075,N_6043);
nand U6313 (N_6313,N_6174,N_6112);
nor U6314 (N_6314,N_6075,N_6095);
nor U6315 (N_6315,N_6037,N_6058);
xor U6316 (N_6316,N_6192,N_6029);
nor U6317 (N_6317,N_6094,N_6025);
nor U6318 (N_6318,N_6127,N_6031);
and U6319 (N_6319,N_6052,N_6154);
nand U6320 (N_6320,N_6175,N_6057);
or U6321 (N_6321,N_6166,N_6165);
and U6322 (N_6322,N_6148,N_6188);
xor U6323 (N_6323,N_6048,N_6128);
nor U6324 (N_6324,N_6039,N_6062);
nand U6325 (N_6325,N_6013,N_6055);
xor U6326 (N_6326,N_6095,N_6073);
or U6327 (N_6327,N_6115,N_6085);
nand U6328 (N_6328,N_6171,N_6001);
nand U6329 (N_6329,N_6036,N_6092);
nand U6330 (N_6330,N_6022,N_6090);
and U6331 (N_6331,N_6009,N_6135);
nand U6332 (N_6332,N_6148,N_6143);
xor U6333 (N_6333,N_6033,N_6127);
xnor U6334 (N_6334,N_6144,N_6181);
and U6335 (N_6335,N_6122,N_6041);
nor U6336 (N_6336,N_6051,N_6152);
or U6337 (N_6337,N_6069,N_6128);
nand U6338 (N_6338,N_6053,N_6122);
nand U6339 (N_6339,N_6067,N_6182);
nand U6340 (N_6340,N_6144,N_6046);
and U6341 (N_6341,N_6067,N_6181);
and U6342 (N_6342,N_6177,N_6056);
xnor U6343 (N_6343,N_6138,N_6139);
and U6344 (N_6344,N_6107,N_6030);
nand U6345 (N_6345,N_6181,N_6062);
nand U6346 (N_6346,N_6019,N_6047);
nor U6347 (N_6347,N_6021,N_6031);
xnor U6348 (N_6348,N_6106,N_6105);
nand U6349 (N_6349,N_6118,N_6160);
and U6350 (N_6350,N_6029,N_6164);
xnor U6351 (N_6351,N_6117,N_6198);
or U6352 (N_6352,N_6069,N_6108);
or U6353 (N_6353,N_6152,N_6127);
nand U6354 (N_6354,N_6173,N_6027);
or U6355 (N_6355,N_6148,N_6076);
nor U6356 (N_6356,N_6047,N_6055);
xnor U6357 (N_6357,N_6189,N_6111);
or U6358 (N_6358,N_6155,N_6133);
xnor U6359 (N_6359,N_6028,N_6148);
nor U6360 (N_6360,N_6066,N_6168);
or U6361 (N_6361,N_6190,N_6044);
or U6362 (N_6362,N_6048,N_6181);
and U6363 (N_6363,N_6028,N_6091);
nand U6364 (N_6364,N_6017,N_6031);
and U6365 (N_6365,N_6141,N_6001);
nand U6366 (N_6366,N_6128,N_6103);
or U6367 (N_6367,N_6169,N_6134);
nor U6368 (N_6368,N_6188,N_6172);
nor U6369 (N_6369,N_6060,N_6099);
and U6370 (N_6370,N_6199,N_6130);
or U6371 (N_6371,N_6172,N_6183);
or U6372 (N_6372,N_6163,N_6190);
nand U6373 (N_6373,N_6111,N_6138);
nor U6374 (N_6374,N_6125,N_6108);
nand U6375 (N_6375,N_6018,N_6033);
nor U6376 (N_6376,N_6114,N_6108);
nor U6377 (N_6377,N_6081,N_6158);
or U6378 (N_6378,N_6022,N_6111);
and U6379 (N_6379,N_6084,N_6097);
and U6380 (N_6380,N_6018,N_6146);
or U6381 (N_6381,N_6098,N_6068);
or U6382 (N_6382,N_6116,N_6027);
xor U6383 (N_6383,N_6185,N_6118);
and U6384 (N_6384,N_6010,N_6059);
or U6385 (N_6385,N_6012,N_6065);
and U6386 (N_6386,N_6144,N_6193);
and U6387 (N_6387,N_6172,N_6061);
nand U6388 (N_6388,N_6062,N_6074);
nor U6389 (N_6389,N_6184,N_6132);
nor U6390 (N_6390,N_6160,N_6046);
or U6391 (N_6391,N_6130,N_6129);
xnor U6392 (N_6392,N_6128,N_6147);
xnor U6393 (N_6393,N_6042,N_6063);
nand U6394 (N_6394,N_6126,N_6095);
xor U6395 (N_6395,N_6168,N_6093);
or U6396 (N_6396,N_6137,N_6077);
xor U6397 (N_6397,N_6135,N_6159);
and U6398 (N_6398,N_6027,N_6077);
nor U6399 (N_6399,N_6128,N_6153);
xnor U6400 (N_6400,N_6307,N_6275);
xnor U6401 (N_6401,N_6205,N_6389);
and U6402 (N_6402,N_6255,N_6394);
and U6403 (N_6403,N_6238,N_6281);
and U6404 (N_6404,N_6237,N_6257);
nor U6405 (N_6405,N_6256,N_6339);
or U6406 (N_6406,N_6251,N_6223);
nand U6407 (N_6407,N_6336,N_6371);
nand U6408 (N_6408,N_6326,N_6213);
nor U6409 (N_6409,N_6364,N_6321);
or U6410 (N_6410,N_6274,N_6309);
nand U6411 (N_6411,N_6249,N_6385);
nand U6412 (N_6412,N_6342,N_6357);
nor U6413 (N_6413,N_6291,N_6219);
nand U6414 (N_6414,N_6324,N_6315);
and U6415 (N_6415,N_6368,N_6383);
and U6416 (N_6416,N_6360,N_6304);
and U6417 (N_6417,N_6397,N_6333);
and U6418 (N_6418,N_6280,N_6317);
or U6419 (N_6419,N_6367,N_6253);
and U6420 (N_6420,N_6395,N_6267);
or U6421 (N_6421,N_6334,N_6209);
xor U6422 (N_6422,N_6240,N_6374);
or U6423 (N_6423,N_6245,N_6378);
and U6424 (N_6424,N_6277,N_6252);
and U6425 (N_6425,N_6361,N_6391);
nor U6426 (N_6426,N_6396,N_6262);
nand U6427 (N_6427,N_6311,N_6289);
or U6428 (N_6428,N_6201,N_6313);
nand U6429 (N_6429,N_6387,N_6375);
or U6430 (N_6430,N_6355,N_6233);
or U6431 (N_6431,N_6384,N_6327);
or U6432 (N_6432,N_6300,N_6379);
nand U6433 (N_6433,N_6398,N_6325);
xnor U6434 (N_6434,N_6369,N_6386);
xnor U6435 (N_6435,N_6295,N_6218);
and U6436 (N_6436,N_6380,N_6376);
xor U6437 (N_6437,N_6299,N_6335);
nor U6438 (N_6438,N_6363,N_6263);
and U6439 (N_6439,N_6270,N_6346);
nand U6440 (N_6440,N_6235,N_6316);
and U6441 (N_6441,N_6344,N_6246);
nor U6442 (N_6442,N_6210,N_6328);
or U6443 (N_6443,N_6232,N_6258);
and U6444 (N_6444,N_6388,N_6259);
xnor U6445 (N_6445,N_6296,N_6207);
nor U6446 (N_6446,N_6260,N_6338);
nor U6447 (N_6447,N_6382,N_6276);
xnor U6448 (N_6448,N_6217,N_6293);
or U6449 (N_6449,N_6362,N_6393);
nor U6450 (N_6450,N_6312,N_6265);
nand U6451 (N_6451,N_6337,N_6211);
or U6452 (N_6452,N_6202,N_6297);
or U6453 (N_6453,N_6248,N_6279);
nor U6454 (N_6454,N_6266,N_6377);
or U6455 (N_6455,N_6352,N_6347);
or U6456 (N_6456,N_6332,N_6216);
nand U6457 (N_6457,N_6239,N_6323);
xnor U6458 (N_6458,N_6345,N_6206);
nand U6459 (N_6459,N_6225,N_6243);
xnor U6460 (N_6460,N_6200,N_6340);
nand U6461 (N_6461,N_6208,N_6349);
xor U6462 (N_6462,N_6322,N_6222);
and U6463 (N_6463,N_6372,N_6241);
nor U6464 (N_6464,N_6278,N_6306);
or U6465 (N_6465,N_6230,N_6390);
or U6466 (N_6466,N_6305,N_6254);
nor U6467 (N_6467,N_6351,N_6353);
nand U6468 (N_6468,N_6301,N_6220);
and U6469 (N_6469,N_6204,N_6356);
nand U6470 (N_6470,N_6286,N_6273);
nor U6471 (N_6471,N_6365,N_6294);
xnor U6472 (N_6472,N_6242,N_6284);
or U6473 (N_6473,N_6214,N_6227);
nor U6474 (N_6474,N_6354,N_6268);
xor U6475 (N_6475,N_6308,N_6203);
nand U6476 (N_6476,N_6226,N_6271);
nand U6477 (N_6477,N_6350,N_6282);
and U6478 (N_6478,N_6269,N_6215);
nand U6479 (N_6479,N_6359,N_6341);
or U6480 (N_6480,N_6283,N_6399);
xor U6481 (N_6481,N_6292,N_6261);
or U6482 (N_6482,N_6212,N_6329);
and U6483 (N_6483,N_6224,N_6381);
or U6484 (N_6484,N_6234,N_6231);
and U6485 (N_6485,N_6392,N_6348);
xor U6486 (N_6486,N_6318,N_6264);
nand U6487 (N_6487,N_6319,N_6244);
nand U6488 (N_6488,N_6236,N_6298);
and U6489 (N_6489,N_6287,N_6247);
and U6490 (N_6490,N_6290,N_6302);
and U6491 (N_6491,N_6314,N_6320);
and U6492 (N_6492,N_6370,N_6229);
nand U6493 (N_6493,N_6250,N_6288);
xnor U6494 (N_6494,N_6373,N_6343);
or U6495 (N_6495,N_6358,N_6285);
xnor U6496 (N_6496,N_6330,N_6303);
xnor U6497 (N_6497,N_6366,N_6272);
xor U6498 (N_6498,N_6221,N_6228);
xor U6499 (N_6499,N_6310,N_6331);
nor U6500 (N_6500,N_6276,N_6305);
or U6501 (N_6501,N_6370,N_6269);
nor U6502 (N_6502,N_6254,N_6375);
nand U6503 (N_6503,N_6360,N_6212);
xnor U6504 (N_6504,N_6251,N_6378);
nor U6505 (N_6505,N_6201,N_6271);
xor U6506 (N_6506,N_6321,N_6204);
xor U6507 (N_6507,N_6341,N_6241);
or U6508 (N_6508,N_6316,N_6320);
and U6509 (N_6509,N_6373,N_6387);
xor U6510 (N_6510,N_6217,N_6372);
nor U6511 (N_6511,N_6359,N_6249);
nor U6512 (N_6512,N_6325,N_6240);
xnor U6513 (N_6513,N_6287,N_6354);
and U6514 (N_6514,N_6248,N_6323);
nand U6515 (N_6515,N_6256,N_6276);
xor U6516 (N_6516,N_6248,N_6209);
and U6517 (N_6517,N_6385,N_6237);
or U6518 (N_6518,N_6310,N_6297);
or U6519 (N_6519,N_6217,N_6260);
nand U6520 (N_6520,N_6343,N_6395);
and U6521 (N_6521,N_6394,N_6239);
nand U6522 (N_6522,N_6355,N_6215);
xor U6523 (N_6523,N_6364,N_6200);
xor U6524 (N_6524,N_6328,N_6225);
nor U6525 (N_6525,N_6376,N_6235);
xnor U6526 (N_6526,N_6347,N_6282);
nor U6527 (N_6527,N_6347,N_6387);
and U6528 (N_6528,N_6329,N_6299);
and U6529 (N_6529,N_6305,N_6382);
or U6530 (N_6530,N_6300,N_6340);
nand U6531 (N_6531,N_6315,N_6240);
xnor U6532 (N_6532,N_6233,N_6311);
nand U6533 (N_6533,N_6256,N_6246);
or U6534 (N_6534,N_6322,N_6324);
or U6535 (N_6535,N_6265,N_6242);
or U6536 (N_6536,N_6326,N_6299);
xnor U6537 (N_6537,N_6205,N_6287);
nand U6538 (N_6538,N_6232,N_6303);
or U6539 (N_6539,N_6339,N_6220);
and U6540 (N_6540,N_6202,N_6246);
xnor U6541 (N_6541,N_6298,N_6332);
xor U6542 (N_6542,N_6313,N_6285);
nor U6543 (N_6543,N_6284,N_6302);
and U6544 (N_6544,N_6366,N_6248);
xor U6545 (N_6545,N_6254,N_6317);
nand U6546 (N_6546,N_6250,N_6222);
and U6547 (N_6547,N_6222,N_6291);
nor U6548 (N_6548,N_6301,N_6317);
nor U6549 (N_6549,N_6292,N_6371);
or U6550 (N_6550,N_6377,N_6386);
nand U6551 (N_6551,N_6393,N_6301);
nand U6552 (N_6552,N_6235,N_6273);
nand U6553 (N_6553,N_6217,N_6248);
nor U6554 (N_6554,N_6372,N_6384);
and U6555 (N_6555,N_6311,N_6378);
and U6556 (N_6556,N_6271,N_6356);
xor U6557 (N_6557,N_6295,N_6252);
nor U6558 (N_6558,N_6203,N_6291);
and U6559 (N_6559,N_6267,N_6276);
xor U6560 (N_6560,N_6395,N_6262);
nand U6561 (N_6561,N_6367,N_6200);
xor U6562 (N_6562,N_6313,N_6329);
nand U6563 (N_6563,N_6306,N_6316);
xor U6564 (N_6564,N_6235,N_6284);
nor U6565 (N_6565,N_6352,N_6343);
nor U6566 (N_6566,N_6351,N_6238);
nand U6567 (N_6567,N_6239,N_6391);
nor U6568 (N_6568,N_6304,N_6313);
or U6569 (N_6569,N_6243,N_6338);
nor U6570 (N_6570,N_6369,N_6363);
or U6571 (N_6571,N_6277,N_6259);
or U6572 (N_6572,N_6228,N_6301);
or U6573 (N_6573,N_6272,N_6363);
nor U6574 (N_6574,N_6391,N_6345);
nor U6575 (N_6575,N_6320,N_6273);
nand U6576 (N_6576,N_6286,N_6394);
nor U6577 (N_6577,N_6361,N_6308);
nor U6578 (N_6578,N_6314,N_6260);
nand U6579 (N_6579,N_6349,N_6217);
xor U6580 (N_6580,N_6390,N_6291);
and U6581 (N_6581,N_6259,N_6284);
nand U6582 (N_6582,N_6232,N_6245);
xor U6583 (N_6583,N_6283,N_6381);
and U6584 (N_6584,N_6244,N_6282);
and U6585 (N_6585,N_6232,N_6343);
or U6586 (N_6586,N_6386,N_6215);
nor U6587 (N_6587,N_6397,N_6217);
xnor U6588 (N_6588,N_6334,N_6395);
xnor U6589 (N_6589,N_6261,N_6341);
xor U6590 (N_6590,N_6366,N_6213);
nor U6591 (N_6591,N_6211,N_6357);
xnor U6592 (N_6592,N_6228,N_6248);
nor U6593 (N_6593,N_6298,N_6323);
or U6594 (N_6594,N_6273,N_6271);
or U6595 (N_6595,N_6294,N_6384);
or U6596 (N_6596,N_6367,N_6248);
xnor U6597 (N_6597,N_6254,N_6291);
and U6598 (N_6598,N_6297,N_6270);
or U6599 (N_6599,N_6336,N_6249);
xor U6600 (N_6600,N_6590,N_6459);
xor U6601 (N_6601,N_6588,N_6593);
or U6602 (N_6602,N_6527,N_6432);
nor U6603 (N_6603,N_6568,N_6472);
and U6604 (N_6604,N_6495,N_6484);
nor U6605 (N_6605,N_6445,N_6596);
xnor U6606 (N_6606,N_6507,N_6574);
or U6607 (N_6607,N_6439,N_6415);
xnor U6608 (N_6608,N_6514,N_6454);
nand U6609 (N_6609,N_6542,N_6558);
or U6610 (N_6610,N_6421,N_6429);
nand U6611 (N_6611,N_6523,N_6557);
or U6612 (N_6612,N_6570,N_6427);
xnor U6613 (N_6613,N_6576,N_6411);
xnor U6614 (N_6614,N_6425,N_6555);
xor U6615 (N_6615,N_6572,N_6410);
xor U6616 (N_6616,N_6506,N_6471);
and U6617 (N_6617,N_6450,N_6591);
or U6618 (N_6618,N_6573,N_6470);
or U6619 (N_6619,N_6420,N_6416);
or U6620 (N_6620,N_6577,N_6564);
nor U6621 (N_6621,N_6476,N_6456);
or U6622 (N_6622,N_6503,N_6419);
nand U6623 (N_6623,N_6464,N_6447);
nor U6624 (N_6624,N_6467,N_6404);
and U6625 (N_6625,N_6569,N_6547);
and U6626 (N_6626,N_6541,N_6442);
and U6627 (N_6627,N_6566,N_6468);
nand U6628 (N_6628,N_6430,N_6431);
nor U6629 (N_6629,N_6490,N_6553);
nand U6630 (N_6630,N_6441,N_6509);
xor U6631 (N_6631,N_6556,N_6453);
and U6632 (N_6632,N_6528,N_6538);
or U6633 (N_6633,N_6589,N_6455);
or U6634 (N_6634,N_6594,N_6409);
xnor U6635 (N_6635,N_6516,N_6436);
nor U6636 (N_6636,N_6504,N_6437);
nand U6637 (N_6637,N_6551,N_6497);
nor U6638 (N_6638,N_6510,N_6443);
xor U6639 (N_6639,N_6451,N_6537);
nor U6640 (N_6640,N_6480,N_6519);
nand U6641 (N_6641,N_6545,N_6444);
xor U6642 (N_6642,N_6406,N_6407);
and U6643 (N_6643,N_6483,N_6546);
xor U6644 (N_6644,N_6563,N_6525);
xnor U6645 (N_6645,N_6446,N_6440);
nor U6646 (N_6646,N_6486,N_6578);
nand U6647 (N_6647,N_6433,N_6599);
nand U6648 (N_6648,N_6526,N_6418);
nand U6649 (N_6649,N_6414,N_6493);
nand U6650 (N_6650,N_6482,N_6531);
or U6651 (N_6651,N_6561,N_6499);
or U6652 (N_6652,N_6417,N_6461);
nand U6653 (N_6653,N_6536,N_6428);
or U6654 (N_6654,N_6449,N_6540);
nand U6655 (N_6655,N_6422,N_6535);
xnor U6656 (N_6656,N_6582,N_6474);
xnor U6657 (N_6657,N_6462,N_6487);
xnor U6658 (N_6658,N_6579,N_6548);
and U6659 (N_6659,N_6508,N_6565);
xnor U6660 (N_6660,N_6585,N_6520);
and U6661 (N_6661,N_6452,N_6494);
or U6662 (N_6662,N_6597,N_6575);
or U6663 (N_6663,N_6400,N_6413);
or U6664 (N_6664,N_6550,N_6581);
xnor U6665 (N_6665,N_6544,N_6522);
and U6666 (N_6666,N_6457,N_6402);
xnor U6667 (N_6667,N_6435,N_6584);
xnor U6668 (N_6668,N_6466,N_6481);
nand U6669 (N_6669,N_6408,N_6517);
or U6670 (N_6670,N_6554,N_6571);
nand U6671 (N_6671,N_6539,N_6423);
nand U6672 (N_6672,N_6401,N_6448);
xor U6673 (N_6673,N_6534,N_6592);
nand U6674 (N_6674,N_6460,N_6586);
nor U6675 (N_6675,N_6598,N_6485);
nor U6676 (N_6676,N_6533,N_6515);
xnor U6677 (N_6677,N_6489,N_6412);
nand U6678 (N_6678,N_6583,N_6473);
and U6679 (N_6679,N_6426,N_6543);
xor U6680 (N_6680,N_6559,N_6463);
xnor U6681 (N_6681,N_6505,N_6502);
or U6682 (N_6682,N_6488,N_6511);
xnor U6683 (N_6683,N_6529,N_6475);
nand U6684 (N_6684,N_6501,N_6478);
nand U6685 (N_6685,N_6434,N_6562);
nor U6686 (N_6686,N_6469,N_6580);
and U6687 (N_6687,N_6518,N_6403);
nand U6688 (N_6688,N_6458,N_6552);
xnor U6689 (N_6689,N_6587,N_6424);
or U6690 (N_6690,N_6530,N_6491);
or U6691 (N_6691,N_6405,N_6479);
nand U6692 (N_6692,N_6549,N_6438);
or U6693 (N_6693,N_6498,N_6513);
xor U6694 (N_6694,N_6567,N_6532);
and U6695 (N_6695,N_6465,N_6595);
or U6696 (N_6696,N_6496,N_6512);
nand U6697 (N_6697,N_6560,N_6524);
nand U6698 (N_6698,N_6500,N_6477);
nand U6699 (N_6699,N_6492,N_6521);
or U6700 (N_6700,N_6594,N_6404);
nor U6701 (N_6701,N_6559,N_6478);
nor U6702 (N_6702,N_6575,N_6526);
or U6703 (N_6703,N_6524,N_6558);
nand U6704 (N_6704,N_6555,N_6504);
nor U6705 (N_6705,N_6507,N_6444);
nand U6706 (N_6706,N_6551,N_6426);
or U6707 (N_6707,N_6564,N_6519);
xnor U6708 (N_6708,N_6431,N_6450);
or U6709 (N_6709,N_6597,N_6413);
xor U6710 (N_6710,N_6480,N_6589);
nand U6711 (N_6711,N_6548,N_6450);
nand U6712 (N_6712,N_6525,N_6405);
nand U6713 (N_6713,N_6590,N_6538);
nand U6714 (N_6714,N_6426,N_6430);
nand U6715 (N_6715,N_6583,N_6513);
and U6716 (N_6716,N_6473,N_6403);
xor U6717 (N_6717,N_6557,N_6421);
nor U6718 (N_6718,N_6463,N_6584);
or U6719 (N_6719,N_6551,N_6594);
nor U6720 (N_6720,N_6579,N_6500);
nand U6721 (N_6721,N_6562,N_6549);
xor U6722 (N_6722,N_6471,N_6560);
xnor U6723 (N_6723,N_6546,N_6404);
nand U6724 (N_6724,N_6562,N_6529);
nand U6725 (N_6725,N_6556,N_6532);
nor U6726 (N_6726,N_6590,N_6579);
nand U6727 (N_6727,N_6587,N_6554);
xor U6728 (N_6728,N_6407,N_6539);
nand U6729 (N_6729,N_6457,N_6547);
nor U6730 (N_6730,N_6455,N_6537);
and U6731 (N_6731,N_6439,N_6529);
nor U6732 (N_6732,N_6420,N_6599);
or U6733 (N_6733,N_6417,N_6435);
xor U6734 (N_6734,N_6490,N_6449);
and U6735 (N_6735,N_6564,N_6517);
xnor U6736 (N_6736,N_6404,N_6522);
or U6737 (N_6737,N_6599,N_6401);
nor U6738 (N_6738,N_6526,N_6530);
nand U6739 (N_6739,N_6527,N_6510);
or U6740 (N_6740,N_6458,N_6434);
xor U6741 (N_6741,N_6430,N_6409);
xor U6742 (N_6742,N_6588,N_6564);
nand U6743 (N_6743,N_6470,N_6457);
or U6744 (N_6744,N_6538,N_6495);
nor U6745 (N_6745,N_6412,N_6446);
xnor U6746 (N_6746,N_6504,N_6406);
and U6747 (N_6747,N_6576,N_6588);
and U6748 (N_6748,N_6446,N_6448);
nor U6749 (N_6749,N_6485,N_6554);
nor U6750 (N_6750,N_6553,N_6508);
nor U6751 (N_6751,N_6438,N_6531);
and U6752 (N_6752,N_6519,N_6560);
nor U6753 (N_6753,N_6436,N_6478);
nor U6754 (N_6754,N_6589,N_6410);
and U6755 (N_6755,N_6565,N_6521);
and U6756 (N_6756,N_6466,N_6441);
nand U6757 (N_6757,N_6411,N_6409);
nand U6758 (N_6758,N_6571,N_6593);
or U6759 (N_6759,N_6456,N_6570);
nand U6760 (N_6760,N_6485,N_6522);
xor U6761 (N_6761,N_6524,N_6485);
xnor U6762 (N_6762,N_6436,N_6470);
or U6763 (N_6763,N_6503,N_6559);
xnor U6764 (N_6764,N_6424,N_6490);
xor U6765 (N_6765,N_6434,N_6406);
and U6766 (N_6766,N_6425,N_6532);
xor U6767 (N_6767,N_6476,N_6564);
xor U6768 (N_6768,N_6463,N_6555);
nor U6769 (N_6769,N_6423,N_6563);
or U6770 (N_6770,N_6521,N_6491);
nand U6771 (N_6771,N_6537,N_6445);
nand U6772 (N_6772,N_6536,N_6526);
xor U6773 (N_6773,N_6402,N_6432);
xor U6774 (N_6774,N_6503,N_6514);
nor U6775 (N_6775,N_6545,N_6573);
nor U6776 (N_6776,N_6480,N_6539);
and U6777 (N_6777,N_6419,N_6429);
and U6778 (N_6778,N_6443,N_6416);
xor U6779 (N_6779,N_6441,N_6568);
or U6780 (N_6780,N_6544,N_6483);
nor U6781 (N_6781,N_6423,N_6400);
and U6782 (N_6782,N_6536,N_6417);
and U6783 (N_6783,N_6473,N_6528);
nand U6784 (N_6784,N_6496,N_6440);
or U6785 (N_6785,N_6537,N_6526);
and U6786 (N_6786,N_6458,N_6592);
and U6787 (N_6787,N_6577,N_6487);
nor U6788 (N_6788,N_6590,N_6522);
nand U6789 (N_6789,N_6477,N_6549);
nor U6790 (N_6790,N_6461,N_6469);
xnor U6791 (N_6791,N_6404,N_6474);
or U6792 (N_6792,N_6480,N_6495);
or U6793 (N_6793,N_6446,N_6405);
nand U6794 (N_6794,N_6514,N_6444);
or U6795 (N_6795,N_6444,N_6404);
or U6796 (N_6796,N_6459,N_6429);
nor U6797 (N_6797,N_6541,N_6561);
or U6798 (N_6798,N_6447,N_6590);
xor U6799 (N_6799,N_6528,N_6492);
nor U6800 (N_6800,N_6641,N_6678);
or U6801 (N_6801,N_6790,N_6631);
or U6802 (N_6802,N_6771,N_6668);
nor U6803 (N_6803,N_6718,N_6603);
xnor U6804 (N_6804,N_6787,N_6647);
nand U6805 (N_6805,N_6646,N_6775);
nand U6806 (N_6806,N_6689,N_6770);
nor U6807 (N_6807,N_6757,N_6731);
or U6808 (N_6808,N_6773,N_6721);
and U6809 (N_6809,N_6791,N_6665);
and U6810 (N_6810,N_6758,N_6772);
xor U6811 (N_6811,N_6632,N_6685);
nor U6812 (N_6812,N_6763,N_6734);
nand U6813 (N_6813,N_6635,N_6760);
or U6814 (N_6814,N_6616,N_6602);
nor U6815 (N_6815,N_6753,N_6686);
xnor U6816 (N_6816,N_6601,N_6710);
nand U6817 (N_6817,N_6722,N_6769);
xor U6818 (N_6818,N_6680,N_6756);
and U6819 (N_6819,N_6645,N_6673);
xor U6820 (N_6820,N_6747,N_6626);
or U6821 (N_6821,N_6767,N_6614);
or U6822 (N_6822,N_6794,N_6785);
and U6823 (N_6823,N_6677,N_6611);
nor U6824 (N_6824,N_6792,N_6666);
nor U6825 (N_6825,N_6630,N_6779);
nor U6826 (N_6826,N_6783,N_6743);
or U6827 (N_6827,N_6663,N_6740);
nor U6828 (N_6828,N_6713,N_6788);
xnor U6829 (N_6829,N_6654,N_6674);
nand U6830 (N_6830,N_6617,N_6634);
nand U6831 (N_6831,N_6711,N_6717);
nor U6832 (N_6832,N_6762,N_6662);
and U6833 (N_6833,N_6620,N_6607);
nor U6834 (N_6834,N_6606,N_6608);
or U6835 (N_6835,N_6719,N_6732);
nor U6836 (N_6836,N_6676,N_6728);
and U6837 (N_6837,N_6696,N_6781);
nor U6838 (N_6838,N_6797,N_6730);
and U6839 (N_6839,N_6667,N_6741);
or U6840 (N_6840,N_6733,N_6774);
xnor U6841 (N_6841,N_6701,N_6746);
and U6842 (N_6842,N_6642,N_6752);
and U6843 (N_6843,N_6604,N_6690);
nor U6844 (N_6844,N_6729,N_6660);
and U6845 (N_6845,N_6652,N_6796);
and U6846 (N_6846,N_6671,N_6655);
nor U6847 (N_6847,N_6633,N_6782);
xnor U6848 (N_6848,N_6789,N_6727);
and U6849 (N_6849,N_6703,N_6681);
nor U6850 (N_6850,N_6610,N_6776);
nor U6851 (N_6851,N_6738,N_6709);
nand U6852 (N_6852,N_6750,N_6748);
and U6853 (N_6853,N_6765,N_6720);
or U6854 (N_6854,N_6777,N_6636);
xor U6855 (N_6855,N_6749,N_6697);
xnor U6856 (N_6856,N_6708,N_6623);
nor U6857 (N_6857,N_6609,N_6798);
nand U6858 (N_6858,N_6659,N_6694);
or U6859 (N_6859,N_6692,N_6651);
xnor U6860 (N_6860,N_6656,N_6695);
nor U6861 (N_6861,N_6706,N_6622);
xnor U6862 (N_6862,N_6736,N_6698);
or U6863 (N_6863,N_6629,N_6640);
xor U6864 (N_6864,N_6702,N_6688);
or U6865 (N_6865,N_6745,N_6742);
nor U6866 (N_6866,N_6764,N_6795);
and U6867 (N_6867,N_6657,N_6786);
nor U6868 (N_6868,N_6682,N_6618);
nor U6869 (N_6869,N_6724,N_6799);
or U6870 (N_6870,N_6683,N_6687);
nor U6871 (N_6871,N_6675,N_6723);
nand U6872 (N_6872,N_6761,N_6715);
xor U6873 (N_6873,N_6613,N_6600);
xor U6874 (N_6874,N_6725,N_6705);
and U6875 (N_6875,N_6670,N_6628);
xnor U6876 (N_6876,N_6637,N_6605);
and U6877 (N_6877,N_6664,N_6625);
xor U6878 (N_6878,N_6627,N_6707);
or U6879 (N_6879,N_6759,N_6704);
and U6880 (N_6880,N_6624,N_6739);
xor U6881 (N_6881,N_6653,N_6621);
xor U6882 (N_6882,N_6693,N_6737);
xor U6883 (N_6883,N_6712,N_6699);
nand U6884 (N_6884,N_6672,N_6755);
nand U6885 (N_6885,N_6639,N_6619);
or U6886 (N_6886,N_6643,N_6780);
nand U6887 (N_6887,N_6615,N_6751);
or U6888 (N_6888,N_6649,N_6754);
nor U6889 (N_6889,N_6644,N_6744);
or U6890 (N_6890,N_6716,N_6714);
nand U6891 (N_6891,N_6612,N_6778);
xor U6892 (N_6892,N_6768,N_6793);
nor U6893 (N_6893,N_6784,N_6661);
nand U6894 (N_6894,N_6658,N_6766);
nand U6895 (N_6895,N_6735,N_6726);
and U6896 (N_6896,N_6700,N_6669);
and U6897 (N_6897,N_6679,N_6691);
nor U6898 (N_6898,N_6650,N_6684);
xor U6899 (N_6899,N_6648,N_6638);
nor U6900 (N_6900,N_6623,N_6633);
nor U6901 (N_6901,N_6639,N_6791);
or U6902 (N_6902,N_6673,N_6608);
nand U6903 (N_6903,N_6696,N_6796);
or U6904 (N_6904,N_6775,N_6796);
or U6905 (N_6905,N_6755,N_6630);
xor U6906 (N_6906,N_6624,N_6617);
xor U6907 (N_6907,N_6605,N_6744);
nand U6908 (N_6908,N_6786,N_6669);
xnor U6909 (N_6909,N_6657,N_6677);
and U6910 (N_6910,N_6752,N_6726);
xor U6911 (N_6911,N_6779,N_6746);
or U6912 (N_6912,N_6610,N_6695);
nor U6913 (N_6913,N_6619,N_6628);
or U6914 (N_6914,N_6764,N_6601);
nor U6915 (N_6915,N_6776,N_6718);
or U6916 (N_6916,N_6673,N_6629);
and U6917 (N_6917,N_6640,N_6637);
and U6918 (N_6918,N_6732,N_6760);
nand U6919 (N_6919,N_6647,N_6712);
or U6920 (N_6920,N_6632,N_6628);
xnor U6921 (N_6921,N_6703,N_6612);
and U6922 (N_6922,N_6761,N_6766);
xor U6923 (N_6923,N_6639,N_6692);
and U6924 (N_6924,N_6775,N_6700);
and U6925 (N_6925,N_6669,N_6668);
nor U6926 (N_6926,N_6737,N_6642);
nand U6927 (N_6927,N_6793,N_6773);
nor U6928 (N_6928,N_6731,N_6760);
and U6929 (N_6929,N_6733,N_6692);
nor U6930 (N_6930,N_6760,N_6775);
and U6931 (N_6931,N_6768,N_6716);
or U6932 (N_6932,N_6763,N_6742);
or U6933 (N_6933,N_6637,N_6740);
nor U6934 (N_6934,N_6618,N_6683);
nand U6935 (N_6935,N_6726,N_6793);
nor U6936 (N_6936,N_6711,N_6668);
xnor U6937 (N_6937,N_6680,N_6709);
xnor U6938 (N_6938,N_6782,N_6777);
nand U6939 (N_6939,N_6746,N_6724);
nor U6940 (N_6940,N_6788,N_6708);
xnor U6941 (N_6941,N_6758,N_6751);
nor U6942 (N_6942,N_6610,N_6690);
nand U6943 (N_6943,N_6627,N_6769);
nor U6944 (N_6944,N_6668,N_6783);
nor U6945 (N_6945,N_6725,N_6793);
and U6946 (N_6946,N_6632,N_6773);
or U6947 (N_6947,N_6672,N_6699);
nor U6948 (N_6948,N_6731,N_6655);
and U6949 (N_6949,N_6659,N_6784);
nor U6950 (N_6950,N_6700,N_6752);
nand U6951 (N_6951,N_6666,N_6700);
nand U6952 (N_6952,N_6751,N_6711);
nor U6953 (N_6953,N_6748,N_6638);
and U6954 (N_6954,N_6719,N_6709);
and U6955 (N_6955,N_6781,N_6705);
nand U6956 (N_6956,N_6625,N_6672);
or U6957 (N_6957,N_6793,N_6743);
and U6958 (N_6958,N_6626,N_6659);
nand U6959 (N_6959,N_6712,N_6667);
nand U6960 (N_6960,N_6754,N_6632);
and U6961 (N_6961,N_6653,N_6776);
nand U6962 (N_6962,N_6674,N_6663);
or U6963 (N_6963,N_6619,N_6617);
nand U6964 (N_6964,N_6758,N_6632);
or U6965 (N_6965,N_6695,N_6672);
or U6966 (N_6966,N_6667,N_6652);
xor U6967 (N_6967,N_6699,N_6654);
nor U6968 (N_6968,N_6688,N_6693);
nand U6969 (N_6969,N_6765,N_6623);
nor U6970 (N_6970,N_6758,N_6642);
xnor U6971 (N_6971,N_6793,N_6739);
nand U6972 (N_6972,N_6788,N_6729);
and U6973 (N_6973,N_6679,N_6624);
xor U6974 (N_6974,N_6699,N_6767);
or U6975 (N_6975,N_6604,N_6730);
xor U6976 (N_6976,N_6763,N_6633);
or U6977 (N_6977,N_6792,N_6610);
and U6978 (N_6978,N_6615,N_6795);
and U6979 (N_6979,N_6782,N_6657);
nor U6980 (N_6980,N_6624,N_6707);
nand U6981 (N_6981,N_6728,N_6776);
nor U6982 (N_6982,N_6681,N_6654);
nand U6983 (N_6983,N_6642,N_6640);
nand U6984 (N_6984,N_6640,N_6776);
nand U6985 (N_6985,N_6792,N_6798);
xor U6986 (N_6986,N_6770,N_6646);
nand U6987 (N_6987,N_6735,N_6728);
xor U6988 (N_6988,N_6729,N_6780);
nor U6989 (N_6989,N_6784,N_6792);
and U6990 (N_6990,N_6662,N_6614);
nor U6991 (N_6991,N_6642,N_6750);
nand U6992 (N_6992,N_6780,N_6602);
nor U6993 (N_6993,N_6602,N_6771);
and U6994 (N_6994,N_6722,N_6736);
nor U6995 (N_6995,N_6745,N_6628);
nand U6996 (N_6996,N_6685,N_6679);
and U6997 (N_6997,N_6771,N_6738);
nand U6998 (N_6998,N_6629,N_6771);
or U6999 (N_6999,N_6754,N_6727);
or U7000 (N_7000,N_6911,N_6960);
or U7001 (N_7001,N_6848,N_6991);
nor U7002 (N_7002,N_6937,N_6861);
nor U7003 (N_7003,N_6899,N_6948);
or U7004 (N_7004,N_6831,N_6995);
and U7005 (N_7005,N_6976,N_6808);
nor U7006 (N_7006,N_6977,N_6913);
nand U7007 (N_7007,N_6971,N_6845);
nor U7008 (N_7008,N_6920,N_6890);
xor U7009 (N_7009,N_6879,N_6873);
or U7010 (N_7010,N_6804,N_6961);
nand U7011 (N_7011,N_6823,N_6963);
xnor U7012 (N_7012,N_6984,N_6935);
nor U7013 (N_7013,N_6933,N_6968);
nor U7014 (N_7014,N_6939,N_6998);
nor U7015 (N_7015,N_6851,N_6989);
and U7016 (N_7016,N_6875,N_6802);
or U7017 (N_7017,N_6815,N_6865);
nand U7018 (N_7018,N_6840,N_6950);
nand U7019 (N_7019,N_6938,N_6807);
nor U7020 (N_7020,N_6874,N_6943);
or U7021 (N_7021,N_6979,N_6908);
nor U7022 (N_7022,N_6967,N_6830);
nor U7023 (N_7023,N_6929,N_6853);
nand U7024 (N_7024,N_6826,N_6932);
nand U7025 (N_7025,N_6816,N_6922);
nand U7026 (N_7026,N_6819,N_6858);
nand U7027 (N_7027,N_6863,N_6942);
nor U7028 (N_7028,N_6949,N_6872);
nand U7029 (N_7029,N_6966,N_6842);
or U7030 (N_7030,N_6849,N_6891);
and U7031 (N_7031,N_6959,N_6994);
xor U7032 (N_7032,N_6981,N_6941);
xor U7033 (N_7033,N_6850,N_6987);
and U7034 (N_7034,N_6925,N_6944);
nor U7035 (N_7035,N_6878,N_6887);
xnor U7036 (N_7036,N_6917,N_6889);
and U7037 (N_7037,N_6880,N_6818);
and U7038 (N_7038,N_6962,N_6864);
nand U7039 (N_7039,N_6817,N_6806);
nand U7040 (N_7040,N_6870,N_6951);
or U7041 (N_7041,N_6834,N_6857);
nand U7042 (N_7042,N_6829,N_6919);
nor U7043 (N_7043,N_6956,N_6847);
nand U7044 (N_7044,N_6869,N_6876);
xor U7045 (N_7045,N_6901,N_6954);
and U7046 (N_7046,N_6905,N_6983);
xnor U7047 (N_7047,N_6997,N_6982);
xor U7048 (N_7048,N_6820,N_6985);
nor U7049 (N_7049,N_6953,N_6811);
nor U7050 (N_7050,N_6996,N_6838);
and U7051 (N_7051,N_6885,N_6900);
nand U7052 (N_7052,N_6812,N_6852);
and U7053 (N_7053,N_6800,N_6821);
nor U7054 (N_7054,N_6973,N_6881);
nor U7055 (N_7055,N_6914,N_6912);
xor U7056 (N_7056,N_6964,N_6980);
nor U7057 (N_7057,N_6888,N_6921);
nand U7058 (N_7058,N_6892,N_6813);
and U7059 (N_7059,N_6945,N_6803);
nor U7060 (N_7060,N_6839,N_6940);
and U7061 (N_7061,N_6836,N_6988);
nand U7062 (N_7062,N_6810,N_6930);
and U7063 (N_7063,N_6934,N_6822);
nor U7064 (N_7064,N_6931,N_6972);
or U7065 (N_7065,N_6978,N_6975);
or U7066 (N_7066,N_6928,N_6859);
nand U7067 (N_7067,N_6906,N_6896);
xnor U7068 (N_7068,N_6832,N_6915);
or U7069 (N_7069,N_6918,N_6936);
nor U7070 (N_7070,N_6801,N_6862);
or U7071 (N_7071,N_6833,N_6986);
nand U7072 (N_7072,N_6814,N_6877);
nand U7073 (N_7073,N_6886,N_6946);
nand U7074 (N_7074,N_6894,N_6805);
or U7075 (N_7075,N_6947,N_6825);
and U7076 (N_7076,N_6824,N_6927);
nor U7077 (N_7077,N_6999,N_6837);
nor U7078 (N_7078,N_6867,N_6882);
nor U7079 (N_7079,N_6957,N_6893);
and U7080 (N_7080,N_6952,N_6854);
or U7081 (N_7081,N_6841,N_6909);
nand U7082 (N_7082,N_6844,N_6898);
and U7083 (N_7083,N_6926,N_6827);
nor U7084 (N_7084,N_6866,N_6907);
or U7085 (N_7085,N_6855,N_6902);
nand U7086 (N_7086,N_6992,N_6843);
or U7087 (N_7087,N_6897,N_6895);
nand U7088 (N_7088,N_6846,N_6904);
nand U7089 (N_7089,N_6993,N_6828);
and U7090 (N_7090,N_6856,N_6809);
or U7091 (N_7091,N_6969,N_6883);
nor U7092 (N_7092,N_6884,N_6910);
or U7093 (N_7093,N_6970,N_6868);
nand U7094 (N_7094,N_6965,N_6974);
and U7095 (N_7095,N_6958,N_6916);
nand U7096 (N_7096,N_6924,N_6835);
nand U7097 (N_7097,N_6923,N_6903);
xor U7098 (N_7098,N_6860,N_6990);
or U7099 (N_7099,N_6955,N_6871);
or U7100 (N_7100,N_6848,N_6993);
nand U7101 (N_7101,N_6913,N_6877);
and U7102 (N_7102,N_6813,N_6931);
or U7103 (N_7103,N_6856,N_6945);
xnor U7104 (N_7104,N_6844,N_6912);
xnor U7105 (N_7105,N_6903,N_6803);
nand U7106 (N_7106,N_6889,N_6908);
nand U7107 (N_7107,N_6820,N_6821);
or U7108 (N_7108,N_6857,N_6931);
nand U7109 (N_7109,N_6968,N_6815);
xor U7110 (N_7110,N_6829,N_6983);
nand U7111 (N_7111,N_6874,N_6953);
xnor U7112 (N_7112,N_6920,N_6880);
and U7113 (N_7113,N_6899,N_6885);
nand U7114 (N_7114,N_6875,N_6828);
or U7115 (N_7115,N_6934,N_6975);
nand U7116 (N_7116,N_6950,N_6865);
or U7117 (N_7117,N_6974,N_6835);
and U7118 (N_7118,N_6892,N_6863);
xnor U7119 (N_7119,N_6959,N_6851);
or U7120 (N_7120,N_6995,N_6898);
nor U7121 (N_7121,N_6996,N_6963);
and U7122 (N_7122,N_6977,N_6921);
xor U7123 (N_7123,N_6974,N_6855);
or U7124 (N_7124,N_6866,N_6961);
nand U7125 (N_7125,N_6913,N_6864);
nand U7126 (N_7126,N_6936,N_6904);
xor U7127 (N_7127,N_6815,N_6989);
and U7128 (N_7128,N_6942,N_6974);
xor U7129 (N_7129,N_6907,N_6972);
or U7130 (N_7130,N_6983,N_6815);
xnor U7131 (N_7131,N_6961,N_6927);
and U7132 (N_7132,N_6984,N_6801);
nor U7133 (N_7133,N_6824,N_6810);
nand U7134 (N_7134,N_6832,N_6974);
nor U7135 (N_7135,N_6803,N_6860);
and U7136 (N_7136,N_6878,N_6949);
nor U7137 (N_7137,N_6822,N_6861);
and U7138 (N_7138,N_6885,N_6803);
nor U7139 (N_7139,N_6833,N_6980);
and U7140 (N_7140,N_6864,N_6984);
xor U7141 (N_7141,N_6906,N_6928);
and U7142 (N_7142,N_6882,N_6940);
and U7143 (N_7143,N_6870,N_6850);
nand U7144 (N_7144,N_6820,N_6871);
and U7145 (N_7145,N_6831,N_6926);
nand U7146 (N_7146,N_6877,N_6848);
nand U7147 (N_7147,N_6858,N_6903);
nand U7148 (N_7148,N_6818,N_6934);
nand U7149 (N_7149,N_6847,N_6981);
xnor U7150 (N_7150,N_6813,N_6822);
xor U7151 (N_7151,N_6877,N_6900);
nand U7152 (N_7152,N_6891,N_6960);
and U7153 (N_7153,N_6960,N_6983);
nor U7154 (N_7154,N_6831,N_6813);
xor U7155 (N_7155,N_6896,N_6868);
xnor U7156 (N_7156,N_6975,N_6838);
or U7157 (N_7157,N_6932,N_6981);
nand U7158 (N_7158,N_6950,N_6885);
nand U7159 (N_7159,N_6824,N_6827);
nand U7160 (N_7160,N_6865,N_6883);
nor U7161 (N_7161,N_6970,N_6932);
nor U7162 (N_7162,N_6961,N_6889);
nand U7163 (N_7163,N_6803,N_6872);
nand U7164 (N_7164,N_6909,N_6852);
nor U7165 (N_7165,N_6850,N_6993);
nor U7166 (N_7166,N_6901,N_6917);
nand U7167 (N_7167,N_6871,N_6984);
nor U7168 (N_7168,N_6942,N_6986);
nor U7169 (N_7169,N_6889,N_6969);
nand U7170 (N_7170,N_6844,N_6969);
or U7171 (N_7171,N_6844,N_6884);
xor U7172 (N_7172,N_6890,N_6932);
nand U7173 (N_7173,N_6816,N_6963);
nand U7174 (N_7174,N_6848,N_6936);
nand U7175 (N_7175,N_6990,N_6845);
nand U7176 (N_7176,N_6842,N_6901);
nor U7177 (N_7177,N_6855,N_6895);
or U7178 (N_7178,N_6888,N_6815);
nand U7179 (N_7179,N_6956,N_6995);
nand U7180 (N_7180,N_6988,N_6830);
and U7181 (N_7181,N_6995,N_6838);
nor U7182 (N_7182,N_6926,N_6970);
nand U7183 (N_7183,N_6945,N_6888);
nand U7184 (N_7184,N_6803,N_6929);
or U7185 (N_7185,N_6837,N_6930);
nand U7186 (N_7186,N_6899,N_6801);
or U7187 (N_7187,N_6904,N_6856);
and U7188 (N_7188,N_6869,N_6868);
nor U7189 (N_7189,N_6847,N_6869);
nand U7190 (N_7190,N_6884,N_6946);
nand U7191 (N_7191,N_6990,N_6868);
nand U7192 (N_7192,N_6971,N_6840);
and U7193 (N_7193,N_6906,N_6850);
nand U7194 (N_7194,N_6850,N_6823);
or U7195 (N_7195,N_6854,N_6997);
xnor U7196 (N_7196,N_6827,N_6935);
xnor U7197 (N_7197,N_6837,N_6992);
nor U7198 (N_7198,N_6876,N_6870);
and U7199 (N_7199,N_6892,N_6990);
nor U7200 (N_7200,N_7017,N_7130);
or U7201 (N_7201,N_7099,N_7118);
nor U7202 (N_7202,N_7088,N_7176);
nand U7203 (N_7203,N_7036,N_7152);
xnor U7204 (N_7204,N_7081,N_7103);
nand U7205 (N_7205,N_7133,N_7053);
xnor U7206 (N_7206,N_7199,N_7027);
and U7207 (N_7207,N_7054,N_7187);
nor U7208 (N_7208,N_7158,N_7097);
and U7209 (N_7209,N_7094,N_7167);
and U7210 (N_7210,N_7083,N_7125);
or U7211 (N_7211,N_7191,N_7020);
xor U7212 (N_7212,N_7196,N_7104);
nand U7213 (N_7213,N_7008,N_7038);
nor U7214 (N_7214,N_7040,N_7122);
or U7215 (N_7215,N_7032,N_7164);
nand U7216 (N_7216,N_7163,N_7136);
nor U7217 (N_7217,N_7064,N_7166);
xor U7218 (N_7218,N_7126,N_7043);
and U7219 (N_7219,N_7102,N_7135);
nand U7220 (N_7220,N_7010,N_7114);
and U7221 (N_7221,N_7192,N_7044);
nand U7222 (N_7222,N_7095,N_7145);
or U7223 (N_7223,N_7091,N_7073);
nand U7224 (N_7224,N_7194,N_7084);
nand U7225 (N_7225,N_7170,N_7089);
nand U7226 (N_7226,N_7157,N_7162);
and U7227 (N_7227,N_7108,N_7177);
xor U7228 (N_7228,N_7056,N_7023);
xor U7229 (N_7229,N_7079,N_7068);
or U7230 (N_7230,N_7193,N_7026);
xnor U7231 (N_7231,N_7065,N_7172);
and U7232 (N_7232,N_7110,N_7061);
and U7233 (N_7233,N_7171,N_7077);
nor U7234 (N_7234,N_7144,N_7123);
nand U7235 (N_7235,N_7074,N_7087);
or U7236 (N_7236,N_7060,N_7030);
nor U7237 (N_7237,N_7150,N_7139);
nor U7238 (N_7238,N_7055,N_7034);
nand U7239 (N_7239,N_7117,N_7012);
xnor U7240 (N_7240,N_7076,N_7131);
and U7241 (N_7241,N_7051,N_7180);
and U7242 (N_7242,N_7156,N_7189);
xnor U7243 (N_7243,N_7041,N_7190);
xnor U7244 (N_7244,N_7132,N_7016);
nand U7245 (N_7245,N_7165,N_7039);
nor U7246 (N_7246,N_7086,N_7022);
nor U7247 (N_7247,N_7174,N_7121);
and U7248 (N_7248,N_7119,N_7113);
and U7249 (N_7249,N_7195,N_7042);
nor U7250 (N_7250,N_7151,N_7109);
and U7251 (N_7251,N_7025,N_7072);
nand U7252 (N_7252,N_7120,N_7063);
or U7253 (N_7253,N_7147,N_7128);
or U7254 (N_7254,N_7045,N_7070);
nand U7255 (N_7255,N_7138,N_7050);
and U7256 (N_7256,N_7052,N_7037);
or U7257 (N_7257,N_7080,N_7127);
or U7258 (N_7258,N_7059,N_7067);
or U7259 (N_7259,N_7029,N_7005);
or U7260 (N_7260,N_7159,N_7015);
nor U7261 (N_7261,N_7071,N_7003);
and U7262 (N_7262,N_7024,N_7137);
nor U7263 (N_7263,N_7149,N_7141);
nor U7264 (N_7264,N_7018,N_7153);
or U7265 (N_7265,N_7142,N_7112);
or U7266 (N_7266,N_7046,N_7000);
or U7267 (N_7267,N_7078,N_7134);
xnor U7268 (N_7268,N_7090,N_7178);
nor U7269 (N_7269,N_7182,N_7093);
xor U7270 (N_7270,N_7154,N_7085);
and U7271 (N_7271,N_7013,N_7111);
nand U7272 (N_7272,N_7011,N_7019);
and U7273 (N_7273,N_7069,N_7098);
or U7274 (N_7274,N_7066,N_7175);
nand U7275 (N_7275,N_7129,N_7004);
and U7276 (N_7276,N_7002,N_7105);
or U7277 (N_7277,N_7007,N_7148);
xor U7278 (N_7278,N_7062,N_7198);
nor U7279 (N_7279,N_7009,N_7047);
xor U7280 (N_7280,N_7106,N_7082);
xor U7281 (N_7281,N_7115,N_7049);
xor U7282 (N_7282,N_7031,N_7186);
or U7283 (N_7283,N_7101,N_7075);
nand U7284 (N_7284,N_7161,N_7116);
nand U7285 (N_7285,N_7096,N_7124);
xor U7286 (N_7286,N_7160,N_7014);
nor U7287 (N_7287,N_7183,N_7057);
nand U7288 (N_7288,N_7155,N_7033);
and U7289 (N_7289,N_7140,N_7188);
and U7290 (N_7290,N_7021,N_7146);
and U7291 (N_7291,N_7028,N_7100);
nor U7292 (N_7292,N_7092,N_7181);
nor U7293 (N_7293,N_7168,N_7048);
or U7294 (N_7294,N_7169,N_7107);
nand U7295 (N_7295,N_7185,N_7184);
nor U7296 (N_7296,N_7173,N_7035);
or U7297 (N_7297,N_7006,N_7143);
nand U7298 (N_7298,N_7058,N_7001);
xnor U7299 (N_7299,N_7197,N_7179);
nand U7300 (N_7300,N_7043,N_7089);
and U7301 (N_7301,N_7047,N_7045);
or U7302 (N_7302,N_7175,N_7067);
nand U7303 (N_7303,N_7002,N_7063);
xnor U7304 (N_7304,N_7142,N_7064);
and U7305 (N_7305,N_7081,N_7140);
or U7306 (N_7306,N_7053,N_7142);
or U7307 (N_7307,N_7022,N_7010);
nand U7308 (N_7308,N_7042,N_7132);
xnor U7309 (N_7309,N_7179,N_7067);
and U7310 (N_7310,N_7103,N_7039);
or U7311 (N_7311,N_7185,N_7180);
nor U7312 (N_7312,N_7197,N_7164);
nand U7313 (N_7313,N_7150,N_7159);
xnor U7314 (N_7314,N_7014,N_7062);
nand U7315 (N_7315,N_7146,N_7095);
xnor U7316 (N_7316,N_7018,N_7066);
xor U7317 (N_7317,N_7070,N_7023);
xnor U7318 (N_7318,N_7045,N_7166);
nor U7319 (N_7319,N_7144,N_7000);
or U7320 (N_7320,N_7010,N_7046);
nand U7321 (N_7321,N_7191,N_7003);
xor U7322 (N_7322,N_7006,N_7144);
and U7323 (N_7323,N_7163,N_7185);
or U7324 (N_7324,N_7173,N_7051);
xnor U7325 (N_7325,N_7006,N_7001);
nor U7326 (N_7326,N_7193,N_7092);
and U7327 (N_7327,N_7146,N_7012);
xnor U7328 (N_7328,N_7181,N_7154);
nand U7329 (N_7329,N_7032,N_7102);
nor U7330 (N_7330,N_7131,N_7189);
nor U7331 (N_7331,N_7075,N_7116);
nand U7332 (N_7332,N_7032,N_7061);
xor U7333 (N_7333,N_7130,N_7026);
nand U7334 (N_7334,N_7111,N_7032);
nand U7335 (N_7335,N_7027,N_7091);
xnor U7336 (N_7336,N_7152,N_7151);
xor U7337 (N_7337,N_7195,N_7099);
xor U7338 (N_7338,N_7112,N_7069);
or U7339 (N_7339,N_7010,N_7067);
nand U7340 (N_7340,N_7135,N_7123);
xnor U7341 (N_7341,N_7168,N_7149);
and U7342 (N_7342,N_7121,N_7041);
nor U7343 (N_7343,N_7075,N_7011);
or U7344 (N_7344,N_7084,N_7078);
xor U7345 (N_7345,N_7139,N_7167);
xnor U7346 (N_7346,N_7005,N_7095);
and U7347 (N_7347,N_7153,N_7006);
and U7348 (N_7348,N_7107,N_7193);
and U7349 (N_7349,N_7094,N_7042);
nand U7350 (N_7350,N_7045,N_7170);
xor U7351 (N_7351,N_7153,N_7143);
nand U7352 (N_7352,N_7002,N_7153);
nand U7353 (N_7353,N_7179,N_7078);
nor U7354 (N_7354,N_7125,N_7163);
and U7355 (N_7355,N_7132,N_7175);
xor U7356 (N_7356,N_7087,N_7078);
or U7357 (N_7357,N_7055,N_7030);
nand U7358 (N_7358,N_7196,N_7010);
nor U7359 (N_7359,N_7180,N_7127);
or U7360 (N_7360,N_7006,N_7080);
or U7361 (N_7361,N_7149,N_7019);
or U7362 (N_7362,N_7044,N_7029);
or U7363 (N_7363,N_7015,N_7154);
or U7364 (N_7364,N_7149,N_7163);
xnor U7365 (N_7365,N_7059,N_7177);
and U7366 (N_7366,N_7191,N_7012);
nor U7367 (N_7367,N_7016,N_7171);
or U7368 (N_7368,N_7001,N_7054);
nor U7369 (N_7369,N_7019,N_7069);
or U7370 (N_7370,N_7024,N_7140);
nand U7371 (N_7371,N_7016,N_7003);
or U7372 (N_7372,N_7134,N_7109);
xor U7373 (N_7373,N_7097,N_7110);
xor U7374 (N_7374,N_7138,N_7145);
and U7375 (N_7375,N_7011,N_7137);
nor U7376 (N_7376,N_7191,N_7016);
xor U7377 (N_7377,N_7145,N_7003);
nor U7378 (N_7378,N_7154,N_7036);
xnor U7379 (N_7379,N_7008,N_7061);
or U7380 (N_7380,N_7146,N_7104);
nand U7381 (N_7381,N_7061,N_7097);
xor U7382 (N_7382,N_7047,N_7161);
and U7383 (N_7383,N_7098,N_7074);
nor U7384 (N_7384,N_7030,N_7058);
xor U7385 (N_7385,N_7058,N_7085);
xnor U7386 (N_7386,N_7181,N_7029);
nor U7387 (N_7387,N_7151,N_7057);
xnor U7388 (N_7388,N_7120,N_7072);
or U7389 (N_7389,N_7130,N_7180);
or U7390 (N_7390,N_7053,N_7192);
xor U7391 (N_7391,N_7118,N_7151);
and U7392 (N_7392,N_7019,N_7018);
and U7393 (N_7393,N_7017,N_7075);
and U7394 (N_7394,N_7021,N_7043);
and U7395 (N_7395,N_7190,N_7144);
nand U7396 (N_7396,N_7080,N_7183);
nor U7397 (N_7397,N_7152,N_7142);
nor U7398 (N_7398,N_7072,N_7196);
or U7399 (N_7399,N_7068,N_7186);
nand U7400 (N_7400,N_7333,N_7286);
nor U7401 (N_7401,N_7255,N_7299);
xor U7402 (N_7402,N_7360,N_7384);
or U7403 (N_7403,N_7395,N_7387);
xor U7404 (N_7404,N_7232,N_7262);
nand U7405 (N_7405,N_7369,N_7338);
xnor U7406 (N_7406,N_7371,N_7319);
nor U7407 (N_7407,N_7249,N_7204);
nand U7408 (N_7408,N_7259,N_7241);
and U7409 (N_7409,N_7270,N_7296);
and U7410 (N_7410,N_7326,N_7356);
nand U7411 (N_7411,N_7378,N_7322);
xnor U7412 (N_7412,N_7372,N_7252);
nand U7413 (N_7413,N_7389,N_7287);
and U7414 (N_7414,N_7201,N_7355);
nand U7415 (N_7415,N_7240,N_7317);
nor U7416 (N_7416,N_7272,N_7218);
and U7417 (N_7417,N_7373,N_7233);
nor U7418 (N_7418,N_7350,N_7311);
xnor U7419 (N_7419,N_7254,N_7244);
or U7420 (N_7420,N_7264,N_7330);
nor U7421 (N_7421,N_7275,N_7346);
nor U7422 (N_7422,N_7344,N_7279);
and U7423 (N_7423,N_7375,N_7250);
nand U7424 (N_7424,N_7261,N_7238);
nor U7425 (N_7425,N_7283,N_7305);
or U7426 (N_7426,N_7285,N_7392);
xor U7427 (N_7427,N_7353,N_7293);
or U7428 (N_7428,N_7328,N_7376);
nor U7429 (N_7429,N_7208,N_7382);
and U7430 (N_7430,N_7303,N_7300);
nand U7431 (N_7431,N_7205,N_7325);
or U7432 (N_7432,N_7341,N_7214);
xor U7433 (N_7433,N_7273,N_7234);
and U7434 (N_7434,N_7267,N_7298);
nor U7435 (N_7435,N_7245,N_7314);
nor U7436 (N_7436,N_7237,N_7291);
xnor U7437 (N_7437,N_7324,N_7334);
and U7438 (N_7438,N_7331,N_7381);
and U7439 (N_7439,N_7390,N_7246);
or U7440 (N_7440,N_7256,N_7310);
and U7441 (N_7441,N_7301,N_7271);
nand U7442 (N_7442,N_7370,N_7380);
and U7443 (N_7443,N_7327,N_7394);
nand U7444 (N_7444,N_7242,N_7351);
nor U7445 (N_7445,N_7231,N_7239);
and U7446 (N_7446,N_7203,N_7363);
xor U7447 (N_7447,N_7225,N_7397);
and U7448 (N_7448,N_7290,N_7251);
nor U7449 (N_7449,N_7348,N_7359);
and U7450 (N_7450,N_7318,N_7398);
nor U7451 (N_7451,N_7294,N_7307);
nand U7452 (N_7452,N_7302,N_7221);
xor U7453 (N_7453,N_7329,N_7399);
nand U7454 (N_7454,N_7364,N_7361);
or U7455 (N_7455,N_7282,N_7385);
nor U7456 (N_7456,N_7253,N_7345);
nor U7457 (N_7457,N_7257,N_7202);
xnor U7458 (N_7458,N_7349,N_7347);
nor U7459 (N_7459,N_7321,N_7343);
nand U7460 (N_7460,N_7222,N_7217);
and U7461 (N_7461,N_7263,N_7223);
and U7462 (N_7462,N_7247,N_7374);
nand U7463 (N_7463,N_7243,N_7352);
nor U7464 (N_7464,N_7269,N_7391);
xnor U7465 (N_7465,N_7268,N_7228);
nand U7466 (N_7466,N_7288,N_7226);
xor U7467 (N_7467,N_7277,N_7332);
nor U7468 (N_7468,N_7278,N_7216);
and U7469 (N_7469,N_7362,N_7377);
nand U7470 (N_7470,N_7368,N_7211);
nand U7471 (N_7471,N_7213,N_7393);
xor U7472 (N_7472,N_7207,N_7340);
xnor U7473 (N_7473,N_7236,N_7336);
nor U7474 (N_7474,N_7337,N_7366);
nor U7475 (N_7475,N_7312,N_7306);
nor U7476 (N_7476,N_7365,N_7280);
nand U7477 (N_7477,N_7274,N_7335);
nand U7478 (N_7478,N_7309,N_7212);
xor U7479 (N_7479,N_7396,N_7383);
nor U7480 (N_7480,N_7266,N_7292);
or U7481 (N_7481,N_7206,N_7295);
nor U7482 (N_7482,N_7227,N_7276);
xor U7483 (N_7483,N_7386,N_7358);
nand U7484 (N_7484,N_7320,N_7367);
nand U7485 (N_7485,N_7200,N_7219);
nand U7486 (N_7486,N_7258,N_7209);
nand U7487 (N_7487,N_7379,N_7281);
and U7488 (N_7488,N_7342,N_7308);
nor U7489 (N_7489,N_7339,N_7248);
and U7490 (N_7490,N_7315,N_7357);
and U7491 (N_7491,N_7220,N_7224);
and U7492 (N_7492,N_7316,N_7215);
nand U7493 (N_7493,N_7260,N_7235);
and U7494 (N_7494,N_7297,N_7304);
or U7495 (N_7495,N_7313,N_7323);
or U7496 (N_7496,N_7388,N_7289);
or U7497 (N_7497,N_7229,N_7265);
and U7498 (N_7498,N_7354,N_7230);
or U7499 (N_7499,N_7284,N_7210);
xor U7500 (N_7500,N_7237,N_7223);
nor U7501 (N_7501,N_7317,N_7348);
xor U7502 (N_7502,N_7209,N_7263);
xor U7503 (N_7503,N_7397,N_7211);
or U7504 (N_7504,N_7306,N_7309);
xnor U7505 (N_7505,N_7314,N_7205);
nor U7506 (N_7506,N_7216,N_7211);
and U7507 (N_7507,N_7378,N_7392);
and U7508 (N_7508,N_7267,N_7292);
nor U7509 (N_7509,N_7203,N_7249);
and U7510 (N_7510,N_7388,N_7224);
nor U7511 (N_7511,N_7397,N_7254);
nor U7512 (N_7512,N_7360,N_7261);
nor U7513 (N_7513,N_7322,N_7303);
and U7514 (N_7514,N_7349,N_7367);
xnor U7515 (N_7515,N_7315,N_7212);
xnor U7516 (N_7516,N_7209,N_7277);
nand U7517 (N_7517,N_7323,N_7345);
nand U7518 (N_7518,N_7226,N_7326);
or U7519 (N_7519,N_7327,N_7382);
nor U7520 (N_7520,N_7242,N_7311);
nand U7521 (N_7521,N_7343,N_7356);
xor U7522 (N_7522,N_7334,N_7336);
xor U7523 (N_7523,N_7219,N_7292);
nand U7524 (N_7524,N_7381,N_7279);
nor U7525 (N_7525,N_7237,N_7397);
nor U7526 (N_7526,N_7339,N_7358);
xnor U7527 (N_7527,N_7334,N_7220);
xnor U7528 (N_7528,N_7317,N_7232);
nor U7529 (N_7529,N_7258,N_7285);
nor U7530 (N_7530,N_7245,N_7278);
or U7531 (N_7531,N_7312,N_7395);
or U7532 (N_7532,N_7295,N_7287);
xor U7533 (N_7533,N_7221,N_7335);
xor U7534 (N_7534,N_7343,N_7274);
and U7535 (N_7535,N_7351,N_7283);
or U7536 (N_7536,N_7353,N_7301);
or U7537 (N_7537,N_7263,N_7321);
nand U7538 (N_7538,N_7244,N_7292);
nor U7539 (N_7539,N_7251,N_7259);
nor U7540 (N_7540,N_7271,N_7394);
or U7541 (N_7541,N_7205,N_7201);
and U7542 (N_7542,N_7365,N_7222);
xnor U7543 (N_7543,N_7222,N_7315);
nand U7544 (N_7544,N_7352,N_7237);
and U7545 (N_7545,N_7237,N_7346);
and U7546 (N_7546,N_7373,N_7240);
xnor U7547 (N_7547,N_7336,N_7374);
or U7548 (N_7548,N_7215,N_7204);
nand U7549 (N_7549,N_7280,N_7297);
and U7550 (N_7550,N_7237,N_7355);
or U7551 (N_7551,N_7369,N_7287);
nand U7552 (N_7552,N_7275,N_7316);
nor U7553 (N_7553,N_7398,N_7246);
nand U7554 (N_7554,N_7346,N_7314);
or U7555 (N_7555,N_7270,N_7242);
or U7556 (N_7556,N_7232,N_7340);
xor U7557 (N_7557,N_7230,N_7296);
nor U7558 (N_7558,N_7396,N_7282);
or U7559 (N_7559,N_7231,N_7214);
and U7560 (N_7560,N_7325,N_7228);
or U7561 (N_7561,N_7277,N_7261);
xor U7562 (N_7562,N_7241,N_7222);
or U7563 (N_7563,N_7285,N_7394);
nor U7564 (N_7564,N_7277,N_7288);
xnor U7565 (N_7565,N_7286,N_7353);
or U7566 (N_7566,N_7330,N_7338);
nand U7567 (N_7567,N_7324,N_7336);
nor U7568 (N_7568,N_7356,N_7215);
nand U7569 (N_7569,N_7389,N_7228);
nor U7570 (N_7570,N_7291,N_7306);
xor U7571 (N_7571,N_7255,N_7329);
xnor U7572 (N_7572,N_7339,N_7210);
nand U7573 (N_7573,N_7365,N_7392);
and U7574 (N_7574,N_7342,N_7228);
xnor U7575 (N_7575,N_7364,N_7237);
and U7576 (N_7576,N_7213,N_7292);
xnor U7577 (N_7577,N_7332,N_7340);
and U7578 (N_7578,N_7316,N_7337);
and U7579 (N_7579,N_7223,N_7240);
and U7580 (N_7580,N_7389,N_7248);
xnor U7581 (N_7581,N_7349,N_7319);
and U7582 (N_7582,N_7285,N_7341);
and U7583 (N_7583,N_7357,N_7380);
xor U7584 (N_7584,N_7362,N_7263);
xnor U7585 (N_7585,N_7250,N_7247);
xor U7586 (N_7586,N_7377,N_7241);
and U7587 (N_7587,N_7228,N_7398);
and U7588 (N_7588,N_7341,N_7305);
nor U7589 (N_7589,N_7356,N_7294);
xor U7590 (N_7590,N_7330,N_7392);
xnor U7591 (N_7591,N_7270,N_7233);
xnor U7592 (N_7592,N_7341,N_7209);
xnor U7593 (N_7593,N_7312,N_7368);
nor U7594 (N_7594,N_7395,N_7211);
and U7595 (N_7595,N_7246,N_7352);
nand U7596 (N_7596,N_7336,N_7323);
and U7597 (N_7597,N_7396,N_7350);
nand U7598 (N_7598,N_7247,N_7366);
or U7599 (N_7599,N_7308,N_7328);
nand U7600 (N_7600,N_7527,N_7541);
or U7601 (N_7601,N_7538,N_7518);
or U7602 (N_7602,N_7532,N_7597);
nand U7603 (N_7603,N_7529,N_7592);
or U7604 (N_7604,N_7520,N_7453);
and U7605 (N_7605,N_7584,N_7514);
and U7606 (N_7606,N_7556,N_7588);
nor U7607 (N_7607,N_7410,N_7501);
and U7608 (N_7608,N_7544,N_7446);
nand U7609 (N_7609,N_7579,N_7516);
xnor U7610 (N_7610,N_7562,N_7484);
nand U7611 (N_7611,N_7573,N_7472);
or U7612 (N_7612,N_7593,N_7507);
nor U7613 (N_7613,N_7533,N_7517);
and U7614 (N_7614,N_7425,N_7409);
xnor U7615 (N_7615,N_7582,N_7452);
nand U7616 (N_7616,N_7439,N_7570);
and U7617 (N_7617,N_7436,N_7508);
or U7618 (N_7618,N_7447,N_7531);
xor U7619 (N_7619,N_7408,N_7500);
nand U7620 (N_7620,N_7450,N_7553);
and U7621 (N_7621,N_7581,N_7441);
and U7622 (N_7622,N_7568,N_7539);
nand U7623 (N_7623,N_7525,N_7576);
or U7624 (N_7624,N_7481,N_7542);
nor U7625 (N_7625,N_7534,N_7572);
xor U7626 (N_7626,N_7402,N_7459);
xnor U7627 (N_7627,N_7565,N_7415);
or U7628 (N_7628,N_7435,N_7404);
or U7629 (N_7629,N_7543,N_7423);
nor U7630 (N_7630,N_7455,N_7463);
nand U7631 (N_7631,N_7526,N_7523);
and U7632 (N_7632,N_7401,N_7471);
and U7633 (N_7633,N_7434,N_7443);
or U7634 (N_7634,N_7462,N_7496);
nand U7635 (N_7635,N_7480,N_7515);
xnor U7636 (N_7636,N_7492,N_7440);
nand U7637 (N_7637,N_7557,N_7468);
xor U7638 (N_7638,N_7598,N_7499);
xor U7639 (N_7639,N_7438,N_7586);
xnor U7640 (N_7640,N_7420,N_7577);
and U7641 (N_7641,N_7444,N_7550);
nand U7642 (N_7642,N_7491,N_7546);
and U7643 (N_7643,N_7460,N_7449);
or U7644 (N_7644,N_7521,N_7405);
and U7645 (N_7645,N_7416,N_7485);
or U7646 (N_7646,N_7494,N_7596);
or U7647 (N_7647,N_7421,N_7403);
and U7648 (N_7648,N_7571,N_7495);
nand U7649 (N_7649,N_7473,N_7512);
or U7650 (N_7650,N_7498,N_7406);
and U7651 (N_7651,N_7490,N_7413);
xor U7652 (N_7652,N_7424,N_7591);
xnor U7653 (N_7653,N_7427,N_7476);
and U7654 (N_7654,N_7575,N_7564);
xor U7655 (N_7655,N_7547,N_7426);
or U7656 (N_7656,N_7551,N_7545);
nor U7657 (N_7657,N_7549,N_7554);
and U7658 (N_7658,N_7589,N_7563);
nand U7659 (N_7659,N_7535,N_7555);
nand U7660 (N_7660,N_7431,N_7411);
nor U7661 (N_7661,N_7478,N_7530);
xor U7662 (N_7662,N_7457,N_7552);
or U7663 (N_7663,N_7407,N_7493);
nand U7664 (N_7664,N_7497,N_7430);
or U7665 (N_7665,N_7437,N_7519);
nor U7666 (N_7666,N_7400,N_7456);
and U7667 (N_7667,N_7467,N_7432);
nand U7668 (N_7668,N_7505,N_7445);
nand U7669 (N_7669,N_7590,N_7558);
or U7670 (N_7670,N_7482,N_7509);
nor U7671 (N_7671,N_7566,N_7536);
and U7672 (N_7672,N_7418,N_7442);
nor U7673 (N_7673,N_7464,N_7537);
xnor U7674 (N_7674,N_7466,N_7475);
xor U7675 (N_7675,N_7412,N_7448);
and U7676 (N_7676,N_7433,N_7599);
nor U7677 (N_7677,N_7422,N_7574);
and U7678 (N_7678,N_7511,N_7585);
or U7679 (N_7679,N_7506,N_7474);
and U7680 (N_7680,N_7595,N_7528);
nand U7681 (N_7681,N_7548,N_7428);
and U7682 (N_7682,N_7569,N_7479);
xnor U7683 (N_7683,N_7540,N_7487);
xor U7684 (N_7684,N_7417,N_7503);
xor U7685 (N_7685,N_7594,N_7504);
or U7686 (N_7686,N_7522,N_7483);
xnor U7687 (N_7687,N_7580,N_7477);
nand U7688 (N_7688,N_7489,N_7510);
and U7689 (N_7689,N_7559,N_7470);
nor U7690 (N_7690,N_7561,N_7488);
or U7691 (N_7691,N_7451,N_7567);
nor U7692 (N_7692,N_7578,N_7560);
nand U7693 (N_7693,N_7513,N_7454);
or U7694 (N_7694,N_7469,N_7429);
nor U7695 (N_7695,N_7587,N_7465);
nor U7696 (N_7696,N_7524,N_7458);
nor U7697 (N_7697,N_7414,N_7461);
nand U7698 (N_7698,N_7419,N_7486);
nand U7699 (N_7699,N_7583,N_7502);
nand U7700 (N_7700,N_7449,N_7448);
or U7701 (N_7701,N_7402,N_7444);
nand U7702 (N_7702,N_7477,N_7439);
and U7703 (N_7703,N_7529,N_7493);
or U7704 (N_7704,N_7430,N_7453);
nand U7705 (N_7705,N_7419,N_7588);
nor U7706 (N_7706,N_7515,N_7446);
nand U7707 (N_7707,N_7580,N_7588);
or U7708 (N_7708,N_7593,N_7596);
xor U7709 (N_7709,N_7440,N_7429);
or U7710 (N_7710,N_7506,N_7512);
nor U7711 (N_7711,N_7571,N_7529);
and U7712 (N_7712,N_7522,N_7430);
nand U7713 (N_7713,N_7562,N_7591);
and U7714 (N_7714,N_7420,N_7409);
or U7715 (N_7715,N_7483,N_7468);
or U7716 (N_7716,N_7584,N_7412);
or U7717 (N_7717,N_7417,N_7576);
nand U7718 (N_7718,N_7439,N_7423);
nor U7719 (N_7719,N_7424,N_7434);
nor U7720 (N_7720,N_7459,N_7566);
nand U7721 (N_7721,N_7565,N_7419);
or U7722 (N_7722,N_7589,N_7593);
xnor U7723 (N_7723,N_7490,N_7468);
nand U7724 (N_7724,N_7406,N_7537);
or U7725 (N_7725,N_7458,N_7529);
or U7726 (N_7726,N_7572,N_7516);
or U7727 (N_7727,N_7400,N_7434);
nor U7728 (N_7728,N_7492,N_7418);
and U7729 (N_7729,N_7453,N_7441);
and U7730 (N_7730,N_7548,N_7519);
nor U7731 (N_7731,N_7470,N_7495);
and U7732 (N_7732,N_7581,N_7426);
and U7733 (N_7733,N_7440,N_7468);
or U7734 (N_7734,N_7504,N_7522);
xnor U7735 (N_7735,N_7487,N_7580);
or U7736 (N_7736,N_7507,N_7553);
nor U7737 (N_7737,N_7590,N_7568);
and U7738 (N_7738,N_7450,N_7599);
nor U7739 (N_7739,N_7478,N_7584);
xor U7740 (N_7740,N_7468,N_7504);
xor U7741 (N_7741,N_7516,N_7491);
xnor U7742 (N_7742,N_7537,N_7458);
and U7743 (N_7743,N_7564,N_7442);
xnor U7744 (N_7744,N_7467,N_7463);
or U7745 (N_7745,N_7495,N_7557);
nand U7746 (N_7746,N_7518,N_7437);
nand U7747 (N_7747,N_7494,N_7513);
or U7748 (N_7748,N_7495,N_7467);
nor U7749 (N_7749,N_7439,N_7550);
nor U7750 (N_7750,N_7451,N_7436);
nor U7751 (N_7751,N_7563,N_7491);
xnor U7752 (N_7752,N_7575,N_7423);
nand U7753 (N_7753,N_7444,N_7477);
xor U7754 (N_7754,N_7413,N_7494);
and U7755 (N_7755,N_7514,N_7454);
nor U7756 (N_7756,N_7489,N_7409);
nand U7757 (N_7757,N_7465,N_7437);
nor U7758 (N_7758,N_7463,N_7465);
or U7759 (N_7759,N_7441,N_7520);
nand U7760 (N_7760,N_7485,N_7509);
or U7761 (N_7761,N_7547,N_7584);
nand U7762 (N_7762,N_7462,N_7579);
xor U7763 (N_7763,N_7567,N_7575);
and U7764 (N_7764,N_7573,N_7580);
or U7765 (N_7765,N_7426,N_7432);
or U7766 (N_7766,N_7492,N_7414);
nor U7767 (N_7767,N_7557,N_7525);
nand U7768 (N_7768,N_7450,N_7507);
nor U7769 (N_7769,N_7568,N_7412);
or U7770 (N_7770,N_7462,N_7476);
or U7771 (N_7771,N_7505,N_7452);
or U7772 (N_7772,N_7493,N_7478);
and U7773 (N_7773,N_7511,N_7522);
or U7774 (N_7774,N_7512,N_7530);
and U7775 (N_7775,N_7571,N_7488);
nand U7776 (N_7776,N_7429,N_7516);
nor U7777 (N_7777,N_7404,N_7447);
and U7778 (N_7778,N_7499,N_7476);
nor U7779 (N_7779,N_7554,N_7525);
or U7780 (N_7780,N_7495,N_7435);
nor U7781 (N_7781,N_7427,N_7546);
nor U7782 (N_7782,N_7539,N_7449);
and U7783 (N_7783,N_7443,N_7558);
xnor U7784 (N_7784,N_7557,N_7506);
and U7785 (N_7785,N_7453,N_7535);
nand U7786 (N_7786,N_7410,N_7510);
or U7787 (N_7787,N_7552,N_7467);
xor U7788 (N_7788,N_7490,N_7409);
xor U7789 (N_7789,N_7554,N_7535);
or U7790 (N_7790,N_7409,N_7559);
xor U7791 (N_7791,N_7557,N_7412);
and U7792 (N_7792,N_7554,N_7495);
xor U7793 (N_7793,N_7412,N_7477);
and U7794 (N_7794,N_7558,N_7589);
nand U7795 (N_7795,N_7560,N_7445);
nor U7796 (N_7796,N_7528,N_7459);
nor U7797 (N_7797,N_7572,N_7533);
nor U7798 (N_7798,N_7443,N_7503);
and U7799 (N_7799,N_7481,N_7501);
nand U7800 (N_7800,N_7730,N_7698);
or U7801 (N_7801,N_7636,N_7654);
nor U7802 (N_7802,N_7761,N_7768);
and U7803 (N_7803,N_7621,N_7799);
or U7804 (N_7804,N_7655,N_7700);
nand U7805 (N_7805,N_7696,N_7784);
or U7806 (N_7806,N_7732,N_7684);
nor U7807 (N_7807,N_7720,N_7733);
nor U7808 (N_7808,N_7633,N_7686);
xor U7809 (N_7809,N_7744,N_7786);
xnor U7810 (N_7810,N_7779,N_7797);
and U7811 (N_7811,N_7674,N_7618);
nand U7812 (N_7812,N_7665,N_7702);
nor U7813 (N_7813,N_7602,N_7752);
or U7814 (N_7814,N_7650,N_7731);
nand U7815 (N_7815,N_7652,N_7782);
xor U7816 (N_7816,N_7662,N_7699);
or U7817 (N_7817,N_7787,N_7685);
or U7818 (N_7818,N_7758,N_7689);
nor U7819 (N_7819,N_7697,N_7634);
or U7820 (N_7820,N_7766,N_7717);
or U7821 (N_7821,N_7760,N_7794);
nand U7822 (N_7822,N_7785,N_7748);
nor U7823 (N_7823,N_7695,N_7675);
and U7824 (N_7824,N_7656,N_7663);
or U7825 (N_7825,N_7676,N_7778);
nor U7826 (N_7826,N_7745,N_7795);
nor U7827 (N_7827,N_7642,N_7707);
nor U7828 (N_7828,N_7788,N_7764);
xnor U7829 (N_7829,N_7737,N_7666);
nand U7830 (N_7830,N_7770,N_7694);
nor U7831 (N_7831,N_7793,N_7688);
nor U7832 (N_7832,N_7739,N_7701);
nor U7833 (N_7833,N_7651,N_7791);
nor U7834 (N_7834,N_7657,N_7624);
xor U7835 (N_7835,N_7661,N_7678);
nor U7836 (N_7836,N_7783,N_7660);
xnor U7837 (N_7837,N_7682,N_7756);
xnor U7838 (N_7838,N_7677,N_7780);
nor U7839 (N_7839,N_7713,N_7625);
nor U7840 (N_7840,N_7610,N_7798);
or U7841 (N_7841,N_7643,N_7711);
and U7842 (N_7842,N_7723,N_7776);
or U7843 (N_7843,N_7603,N_7635);
and U7844 (N_7844,N_7692,N_7648);
xor U7845 (N_7845,N_7734,N_7749);
xnor U7846 (N_7846,N_7613,N_7743);
nand U7847 (N_7847,N_7637,N_7658);
and U7848 (N_7848,N_7775,N_7649);
nand U7849 (N_7849,N_7726,N_7740);
and U7850 (N_7850,N_7703,N_7769);
nand U7851 (N_7851,N_7659,N_7710);
or U7852 (N_7852,N_7763,N_7622);
nand U7853 (N_7853,N_7600,N_7693);
xnor U7854 (N_7854,N_7691,N_7709);
nand U7855 (N_7855,N_7773,N_7722);
nor U7856 (N_7856,N_7708,N_7690);
xnor U7857 (N_7857,N_7683,N_7771);
nand U7858 (N_7858,N_7774,N_7646);
xor U7859 (N_7859,N_7705,N_7750);
nor U7860 (N_7860,N_7607,N_7746);
nor U7861 (N_7861,N_7647,N_7747);
or U7862 (N_7862,N_7712,N_7605);
xor U7863 (N_7863,N_7725,N_7772);
and U7864 (N_7864,N_7781,N_7606);
nand U7865 (N_7865,N_7653,N_7738);
or U7866 (N_7866,N_7608,N_7753);
or U7867 (N_7867,N_7704,N_7790);
nand U7868 (N_7868,N_7626,N_7792);
or U7869 (N_7869,N_7673,N_7617);
and U7870 (N_7870,N_7714,N_7741);
nand U7871 (N_7871,N_7640,N_7755);
nor U7872 (N_7872,N_7638,N_7757);
nor U7873 (N_7873,N_7718,N_7727);
xor U7874 (N_7874,N_7706,N_7628);
or U7875 (N_7875,N_7614,N_7632);
xor U7876 (N_7876,N_7616,N_7670);
and U7877 (N_7877,N_7631,N_7728);
nand U7878 (N_7878,N_7627,N_7645);
xnor U7879 (N_7879,N_7623,N_7668);
nand U7880 (N_7880,N_7751,N_7664);
nor U7881 (N_7881,N_7762,N_7630);
nor U7882 (N_7882,N_7620,N_7629);
or U7883 (N_7883,N_7767,N_7680);
and U7884 (N_7884,N_7777,N_7619);
and U7885 (N_7885,N_7789,N_7724);
nor U7886 (N_7886,N_7641,N_7601);
nor U7887 (N_7887,N_7609,N_7796);
or U7888 (N_7888,N_7729,N_7735);
nor U7889 (N_7889,N_7765,N_7639);
nor U7890 (N_7890,N_7669,N_7721);
or U7891 (N_7891,N_7719,N_7612);
nor U7892 (N_7892,N_7679,N_7687);
xnor U7893 (N_7893,N_7604,N_7759);
xor U7894 (N_7894,N_7615,N_7672);
and U7895 (N_7895,N_7671,N_7611);
and U7896 (N_7896,N_7754,N_7736);
nor U7897 (N_7897,N_7644,N_7681);
or U7898 (N_7898,N_7742,N_7715);
nor U7899 (N_7899,N_7716,N_7667);
nor U7900 (N_7900,N_7784,N_7798);
nor U7901 (N_7901,N_7676,N_7655);
nor U7902 (N_7902,N_7745,N_7793);
or U7903 (N_7903,N_7718,N_7760);
nand U7904 (N_7904,N_7774,N_7606);
or U7905 (N_7905,N_7642,N_7697);
xor U7906 (N_7906,N_7630,N_7734);
nand U7907 (N_7907,N_7720,N_7677);
and U7908 (N_7908,N_7650,N_7616);
and U7909 (N_7909,N_7659,N_7750);
xnor U7910 (N_7910,N_7757,N_7707);
or U7911 (N_7911,N_7729,N_7646);
nor U7912 (N_7912,N_7628,N_7686);
or U7913 (N_7913,N_7691,N_7771);
nand U7914 (N_7914,N_7751,N_7642);
xnor U7915 (N_7915,N_7779,N_7633);
nand U7916 (N_7916,N_7654,N_7600);
nor U7917 (N_7917,N_7649,N_7749);
nand U7918 (N_7918,N_7742,N_7611);
and U7919 (N_7919,N_7651,N_7782);
nand U7920 (N_7920,N_7618,N_7666);
nor U7921 (N_7921,N_7778,N_7707);
or U7922 (N_7922,N_7619,N_7690);
nor U7923 (N_7923,N_7653,N_7788);
or U7924 (N_7924,N_7673,N_7645);
xnor U7925 (N_7925,N_7714,N_7786);
nand U7926 (N_7926,N_7755,N_7643);
nor U7927 (N_7927,N_7631,N_7635);
nor U7928 (N_7928,N_7742,N_7691);
and U7929 (N_7929,N_7707,N_7709);
or U7930 (N_7930,N_7651,N_7683);
and U7931 (N_7931,N_7657,N_7601);
nand U7932 (N_7932,N_7690,N_7664);
nor U7933 (N_7933,N_7792,N_7613);
nand U7934 (N_7934,N_7701,N_7638);
and U7935 (N_7935,N_7609,N_7728);
and U7936 (N_7936,N_7632,N_7768);
nor U7937 (N_7937,N_7722,N_7775);
and U7938 (N_7938,N_7757,N_7769);
xnor U7939 (N_7939,N_7619,N_7663);
xor U7940 (N_7940,N_7721,N_7743);
nand U7941 (N_7941,N_7795,N_7723);
or U7942 (N_7942,N_7779,N_7664);
nor U7943 (N_7943,N_7695,N_7752);
nand U7944 (N_7944,N_7731,N_7740);
nor U7945 (N_7945,N_7653,N_7706);
xor U7946 (N_7946,N_7677,N_7765);
nor U7947 (N_7947,N_7632,N_7792);
nor U7948 (N_7948,N_7638,N_7641);
and U7949 (N_7949,N_7638,N_7784);
or U7950 (N_7950,N_7610,N_7650);
and U7951 (N_7951,N_7777,N_7785);
or U7952 (N_7952,N_7650,N_7774);
xnor U7953 (N_7953,N_7786,N_7664);
and U7954 (N_7954,N_7720,N_7640);
or U7955 (N_7955,N_7761,N_7754);
xnor U7956 (N_7956,N_7682,N_7642);
or U7957 (N_7957,N_7613,N_7782);
and U7958 (N_7958,N_7718,N_7796);
and U7959 (N_7959,N_7605,N_7754);
xnor U7960 (N_7960,N_7731,N_7687);
nor U7961 (N_7961,N_7770,N_7759);
nor U7962 (N_7962,N_7742,N_7653);
and U7963 (N_7963,N_7705,N_7742);
xnor U7964 (N_7964,N_7655,N_7735);
xnor U7965 (N_7965,N_7797,N_7764);
nor U7966 (N_7966,N_7781,N_7778);
and U7967 (N_7967,N_7611,N_7643);
xor U7968 (N_7968,N_7666,N_7683);
nand U7969 (N_7969,N_7789,N_7790);
nor U7970 (N_7970,N_7781,N_7752);
xnor U7971 (N_7971,N_7716,N_7731);
xnor U7972 (N_7972,N_7766,N_7626);
xor U7973 (N_7973,N_7713,N_7749);
nand U7974 (N_7974,N_7793,N_7729);
xnor U7975 (N_7975,N_7670,N_7792);
and U7976 (N_7976,N_7685,N_7639);
and U7977 (N_7977,N_7712,N_7600);
nor U7978 (N_7978,N_7681,N_7762);
nand U7979 (N_7979,N_7691,N_7662);
or U7980 (N_7980,N_7720,N_7681);
nand U7981 (N_7981,N_7676,N_7649);
nor U7982 (N_7982,N_7763,N_7600);
nand U7983 (N_7983,N_7759,N_7637);
nand U7984 (N_7984,N_7627,N_7757);
nor U7985 (N_7985,N_7666,N_7785);
xnor U7986 (N_7986,N_7659,N_7650);
xnor U7987 (N_7987,N_7691,N_7778);
and U7988 (N_7988,N_7626,N_7676);
nand U7989 (N_7989,N_7696,N_7707);
nor U7990 (N_7990,N_7755,N_7698);
and U7991 (N_7991,N_7644,N_7623);
nand U7992 (N_7992,N_7697,N_7782);
nor U7993 (N_7993,N_7660,N_7786);
and U7994 (N_7994,N_7707,N_7647);
or U7995 (N_7995,N_7637,N_7639);
nor U7996 (N_7996,N_7656,N_7734);
nor U7997 (N_7997,N_7714,N_7606);
nand U7998 (N_7998,N_7668,N_7706);
nand U7999 (N_7999,N_7775,N_7780);
and U8000 (N_8000,N_7866,N_7950);
or U8001 (N_8001,N_7869,N_7846);
or U8002 (N_8002,N_7999,N_7968);
and U8003 (N_8003,N_7962,N_7826);
xor U8004 (N_8004,N_7851,N_7803);
or U8005 (N_8005,N_7888,N_7900);
nand U8006 (N_8006,N_7832,N_7971);
nor U8007 (N_8007,N_7849,N_7923);
nand U8008 (N_8008,N_7981,N_7853);
or U8009 (N_8009,N_7895,N_7877);
nand U8010 (N_8010,N_7997,N_7912);
and U8011 (N_8011,N_7899,N_7914);
xor U8012 (N_8012,N_7865,N_7953);
nor U8013 (N_8013,N_7985,N_7967);
xnor U8014 (N_8014,N_7878,N_7938);
or U8015 (N_8015,N_7945,N_7990);
and U8016 (N_8016,N_7887,N_7951);
xnor U8017 (N_8017,N_7830,N_7860);
or U8018 (N_8018,N_7863,N_7802);
and U8019 (N_8019,N_7933,N_7913);
nand U8020 (N_8020,N_7905,N_7867);
nor U8021 (N_8021,N_7819,N_7848);
nand U8022 (N_8022,N_7957,N_7906);
nand U8023 (N_8023,N_7845,N_7904);
nand U8024 (N_8024,N_7955,N_7822);
xor U8025 (N_8025,N_7874,N_7934);
and U8026 (N_8026,N_7844,N_7927);
nor U8027 (N_8027,N_7935,N_7976);
xor U8028 (N_8028,N_7908,N_7987);
xnor U8029 (N_8029,N_7811,N_7944);
nand U8030 (N_8030,N_7894,N_7902);
nand U8031 (N_8031,N_7804,N_7931);
nand U8032 (N_8032,N_7966,N_7886);
nor U8033 (N_8033,N_7861,N_7806);
xnor U8034 (N_8034,N_7816,N_7831);
xnor U8035 (N_8035,N_7838,N_7864);
nand U8036 (N_8036,N_7977,N_7964);
nand U8037 (N_8037,N_7954,N_7871);
or U8038 (N_8038,N_7858,N_7898);
xnor U8039 (N_8039,N_7984,N_7883);
and U8040 (N_8040,N_7920,N_7921);
or U8041 (N_8041,N_7947,N_7928);
nor U8042 (N_8042,N_7841,N_7896);
nor U8043 (N_8043,N_7907,N_7943);
nor U8044 (N_8044,N_7855,N_7929);
nand U8045 (N_8045,N_7821,N_7918);
nor U8046 (N_8046,N_7872,N_7909);
nand U8047 (N_8047,N_7809,N_7989);
and U8048 (N_8048,N_7959,N_7975);
nor U8049 (N_8049,N_7965,N_7850);
or U8050 (N_8050,N_7972,N_7970);
or U8051 (N_8051,N_7993,N_7926);
nand U8052 (N_8052,N_7979,N_7847);
xnor U8053 (N_8053,N_7857,N_7817);
or U8054 (N_8054,N_7842,N_7910);
or U8055 (N_8055,N_7801,N_7818);
nand U8056 (N_8056,N_7889,N_7949);
or U8057 (N_8057,N_7884,N_7924);
nor U8058 (N_8058,N_7942,N_7958);
and U8059 (N_8059,N_7829,N_7862);
nand U8060 (N_8060,N_7892,N_7882);
xor U8061 (N_8061,N_7805,N_7901);
xnor U8062 (N_8062,N_7880,N_7939);
or U8063 (N_8063,N_7996,N_7808);
xnor U8064 (N_8064,N_7807,N_7988);
or U8065 (N_8065,N_7919,N_7952);
or U8066 (N_8066,N_7856,N_7982);
and U8067 (N_8067,N_7890,N_7941);
nand U8068 (N_8068,N_7814,N_7936);
xor U8069 (N_8069,N_7911,N_7881);
nand U8070 (N_8070,N_7917,N_7946);
or U8071 (N_8071,N_7813,N_7916);
nor U8072 (N_8072,N_7852,N_7932);
and U8073 (N_8073,N_7891,N_7825);
and U8074 (N_8074,N_7980,N_7870);
and U8075 (N_8075,N_7991,N_7983);
and U8076 (N_8076,N_7978,N_7834);
xnor U8077 (N_8077,N_7828,N_7915);
nand U8078 (N_8078,N_7956,N_7961);
xor U8079 (N_8079,N_7820,N_7812);
or U8080 (N_8080,N_7800,N_7995);
nand U8081 (N_8081,N_7837,N_7925);
or U8082 (N_8082,N_7835,N_7973);
or U8083 (N_8083,N_7986,N_7815);
or U8084 (N_8084,N_7974,N_7843);
or U8085 (N_8085,N_7998,N_7937);
and U8086 (N_8086,N_7827,N_7948);
nor U8087 (N_8087,N_7810,N_7836);
nand U8088 (N_8088,N_7893,N_7994);
and U8089 (N_8089,N_7873,N_7854);
nor U8090 (N_8090,N_7940,N_7875);
nor U8091 (N_8091,N_7859,N_7839);
xnor U8092 (N_8092,N_7897,N_7876);
xnor U8093 (N_8093,N_7930,N_7960);
nor U8094 (N_8094,N_7840,N_7969);
and U8095 (N_8095,N_7963,N_7903);
xnor U8096 (N_8096,N_7879,N_7823);
or U8097 (N_8097,N_7824,N_7868);
or U8098 (N_8098,N_7885,N_7992);
or U8099 (N_8099,N_7922,N_7833);
xor U8100 (N_8100,N_7943,N_7995);
nor U8101 (N_8101,N_7863,N_7895);
nand U8102 (N_8102,N_7870,N_7933);
nor U8103 (N_8103,N_7972,N_7881);
nand U8104 (N_8104,N_7906,N_7831);
or U8105 (N_8105,N_7998,N_7832);
or U8106 (N_8106,N_7946,N_7863);
nor U8107 (N_8107,N_7962,N_7815);
and U8108 (N_8108,N_7979,N_7861);
nand U8109 (N_8109,N_7821,N_7959);
xnor U8110 (N_8110,N_7900,N_7913);
and U8111 (N_8111,N_7811,N_7939);
nor U8112 (N_8112,N_7955,N_7818);
and U8113 (N_8113,N_7935,N_7893);
nor U8114 (N_8114,N_7810,N_7802);
and U8115 (N_8115,N_7855,N_7847);
nand U8116 (N_8116,N_7930,N_7915);
and U8117 (N_8117,N_7869,N_7831);
or U8118 (N_8118,N_7811,N_7963);
and U8119 (N_8119,N_7909,N_7929);
and U8120 (N_8120,N_7846,N_7991);
nor U8121 (N_8121,N_7999,N_7962);
xnor U8122 (N_8122,N_7918,N_7866);
and U8123 (N_8123,N_7947,N_7952);
and U8124 (N_8124,N_7979,N_7903);
nor U8125 (N_8125,N_7847,N_7987);
and U8126 (N_8126,N_7945,N_7976);
nand U8127 (N_8127,N_7994,N_7878);
xor U8128 (N_8128,N_7963,N_7979);
and U8129 (N_8129,N_7824,N_7937);
and U8130 (N_8130,N_7869,N_7844);
or U8131 (N_8131,N_7939,N_7995);
xor U8132 (N_8132,N_7992,N_7962);
nand U8133 (N_8133,N_7908,N_7929);
nor U8134 (N_8134,N_7806,N_7902);
or U8135 (N_8135,N_7870,N_7963);
xnor U8136 (N_8136,N_7839,N_7802);
xor U8137 (N_8137,N_7881,N_7900);
or U8138 (N_8138,N_7832,N_7979);
or U8139 (N_8139,N_7905,N_7864);
or U8140 (N_8140,N_7970,N_7958);
and U8141 (N_8141,N_7824,N_7896);
or U8142 (N_8142,N_7901,N_7852);
nand U8143 (N_8143,N_7814,N_7941);
nor U8144 (N_8144,N_7851,N_7801);
xor U8145 (N_8145,N_7960,N_7812);
or U8146 (N_8146,N_7842,N_7967);
and U8147 (N_8147,N_7915,N_7972);
xor U8148 (N_8148,N_7819,N_7820);
nor U8149 (N_8149,N_7943,N_7972);
and U8150 (N_8150,N_7803,N_7957);
nor U8151 (N_8151,N_7893,N_7907);
nand U8152 (N_8152,N_7830,N_7960);
nand U8153 (N_8153,N_7829,N_7850);
nand U8154 (N_8154,N_7913,N_7944);
nor U8155 (N_8155,N_7875,N_7933);
xor U8156 (N_8156,N_7850,N_7943);
nor U8157 (N_8157,N_7803,N_7863);
nand U8158 (N_8158,N_7917,N_7973);
nand U8159 (N_8159,N_7851,N_7905);
xnor U8160 (N_8160,N_7802,N_7871);
or U8161 (N_8161,N_7881,N_7891);
or U8162 (N_8162,N_7814,N_7905);
and U8163 (N_8163,N_7874,N_7999);
or U8164 (N_8164,N_7814,N_7929);
and U8165 (N_8165,N_7886,N_7894);
nor U8166 (N_8166,N_7813,N_7966);
nor U8167 (N_8167,N_7980,N_7932);
and U8168 (N_8168,N_7933,N_7834);
nand U8169 (N_8169,N_7972,N_7969);
nor U8170 (N_8170,N_7880,N_7920);
nand U8171 (N_8171,N_7904,N_7867);
or U8172 (N_8172,N_7809,N_7872);
or U8173 (N_8173,N_7912,N_7901);
or U8174 (N_8174,N_7839,N_7806);
nand U8175 (N_8175,N_7921,N_7959);
nand U8176 (N_8176,N_7922,N_7977);
xnor U8177 (N_8177,N_7852,N_7906);
and U8178 (N_8178,N_7977,N_7826);
nor U8179 (N_8179,N_7985,N_7868);
or U8180 (N_8180,N_7995,N_7814);
and U8181 (N_8181,N_7891,N_7984);
nand U8182 (N_8182,N_7944,N_7800);
nor U8183 (N_8183,N_7838,N_7980);
or U8184 (N_8184,N_7965,N_7996);
nor U8185 (N_8185,N_7850,N_7983);
xnor U8186 (N_8186,N_7874,N_7851);
xor U8187 (N_8187,N_7938,N_7932);
nand U8188 (N_8188,N_7996,N_7978);
nor U8189 (N_8189,N_7988,N_7960);
or U8190 (N_8190,N_7838,N_7863);
nand U8191 (N_8191,N_7864,N_7998);
and U8192 (N_8192,N_7870,N_7808);
nand U8193 (N_8193,N_7908,N_7824);
and U8194 (N_8194,N_7881,N_7838);
xnor U8195 (N_8195,N_7825,N_7988);
nor U8196 (N_8196,N_7857,N_7871);
or U8197 (N_8197,N_7852,N_7915);
nor U8198 (N_8198,N_7920,N_7837);
and U8199 (N_8199,N_7926,N_7998);
and U8200 (N_8200,N_8049,N_8039);
or U8201 (N_8201,N_8190,N_8088);
and U8202 (N_8202,N_8196,N_8022);
nand U8203 (N_8203,N_8185,N_8090);
xor U8204 (N_8204,N_8146,N_8063);
xnor U8205 (N_8205,N_8105,N_8015);
or U8206 (N_8206,N_8149,N_8156);
and U8207 (N_8207,N_8113,N_8059);
nor U8208 (N_8208,N_8037,N_8019);
xor U8209 (N_8209,N_8081,N_8013);
nand U8210 (N_8210,N_8048,N_8045);
and U8211 (N_8211,N_8099,N_8128);
or U8212 (N_8212,N_8000,N_8136);
nor U8213 (N_8213,N_8165,N_8121);
nand U8214 (N_8214,N_8100,N_8023);
nor U8215 (N_8215,N_8009,N_8135);
or U8216 (N_8216,N_8043,N_8192);
and U8217 (N_8217,N_8032,N_8166);
nor U8218 (N_8218,N_8142,N_8034);
or U8219 (N_8219,N_8064,N_8096);
nor U8220 (N_8220,N_8132,N_8016);
and U8221 (N_8221,N_8069,N_8175);
and U8222 (N_8222,N_8057,N_8127);
and U8223 (N_8223,N_8078,N_8199);
and U8224 (N_8224,N_8044,N_8188);
nand U8225 (N_8225,N_8062,N_8024);
xnor U8226 (N_8226,N_8020,N_8038);
nand U8227 (N_8227,N_8066,N_8179);
nor U8228 (N_8228,N_8089,N_8193);
xnor U8229 (N_8229,N_8046,N_8082);
nor U8230 (N_8230,N_8126,N_8195);
or U8231 (N_8231,N_8076,N_8180);
and U8232 (N_8232,N_8012,N_8025);
nor U8233 (N_8233,N_8083,N_8047);
or U8234 (N_8234,N_8040,N_8182);
nand U8235 (N_8235,N_8055,N_8177);
or U8236 (N_8236,N_8129,N_8116);
or U8237 (N_8237,N_8007,N_8031);
and U8238 (N_8238,N_8005,N_8109);
or U8239 (N_8239,N_8001,N_8077);
xor U8240 (N_8240,N_8178,N_8115);
xor U8241 (N_8241,N_8150,N_8094);
or U8242 (N_8242,N_8004,N_8067);
nand U8243 (N_8243,N_8120,N_8098);
nand U8244 (N_8244,N_8060,N_8189);
xnor U8245 (N_8245,N_8042,N_8041);
nor U8246 (N_8246,N_8006,N_8137);
and U8247 (N_8247,N_8071,N_8170);
or U8248 (N_8248,N_8052,N_8107);
nand U8249 (N_8249,N_8187,N_8171);
nor U8250 (N_8250,N_8065,N_8134);
nand U8251 (N_8251,N_8173,N_8075);
nor U8252 (N_8252,N_8161,N_8079);
nand U8253 (N_8253,N_8144,N_8035);
or U8254 (N_8254,N_8140,N_8074);
nor U8255 (N_8255,N_8036,N_8027);
nor U8256 (N_8256,N_8124,N_8097);
nand U8257 (N_8257,N_8111,N_8160);
or U8258 (N_8258,N_8017,N_8086);
nor U8259 (N_8259,N_8174,N_8104);
and U8260 (N_8260,N_8114,N_8197);
nor U8261 (N_8261,N_8151,N_8084);
nor U8262 (N_8262,N_8145,N_8085);
nand U8263 (N_8263,N_8147,N_8158);
or U8264 (N_8264,N_8125,N_8010);
or U8265 (N_8265,N_8021,N_8110);
nand U8266 (N_8266,N_8053,N_8153);
and U8267 (N_8267,N_8108,N_8058);
or U8268 (N_8268,N_8117,N_8148);
xnor U8269 (N_8269,N_8186,N_8139);
and U8270 (N_8270,N_8061,N_8183);
and U8271 (N_8271,N_8159,N_8131);
nor U8272 (N_8272,N_8051,N_8008);
xor U8273 (N_8273,N_8068,N_8154);
nand U8274 (N_8274,N_8181,N_8162);
nand U8275 (N_8275,N_8123,N_8091);
and U8276 (N_8276,N_8092,N_8080);
or U8277 (N_8277,N_8033,N_8164);
xnor U8278 (N_8278,N_8102,N_8169);
and U8279 (N_8279,N_8026,N_8141);
nor U8280 (N_8280,N_8029,N_8018);
nor U8281 (N_8281,N_8130,N_8198);
or U8282 (N_8282,N_8103,N_8003);
xor U8283 (N_8283,N_8176,N_8106);
nor U8284 (N_8284,N_8157,N_8070);
and U8285 (N_8285,N_8028,N_8112);
nor U8286 (N_8286,N_8030,N_8133);
or U8287 (N_8287,N_8118,N_8087);
and U8288 (N_8288,N_8073,N_8163);
nand U8289 (N_8289,N_8050,N_8093);
xor U8290 (N_8290,N_8072,N_8054);
nor U8291 (N_8291,N_8101,N_8191);
or U8292 (N_8292,N_8168,N_8138);
nor U8293 (N_8293,N_8143,N_8184);
or U8294 (N_8294,N_8119,N_8014);
nand U8295 (N_8295,N_8002,N_8011);
and U8296 (N_8296,N_8152,N_8056);
nor U8297 (N_8297,N_8167,N_8122);
nor U8298 (N_8298,N_8095,N_8155);
nand U8299 (N_8299,N_8194,N_8172);
and U8300 (N_8300,N_8172,N_8104);
xor U8301 (N_8301,N_8087,N_8036);
nor U8302 (N_8302,N_8178,N_8092);
nor U8303 (N_8303,N_8038,N_8024);
nand U8304 (N_8304,N_8184,N_8025);
nor U8305 (N_8305,N_8094,N_8041);
and U8306 (N_8306,N_8087,N_8102);
and U8307 (N_8307,N_8022,N_8119);
or U8308 (N_8308,N_8114,N_8018);
or U8309 (N_8309,N_8107,N_8190);
nor U8310 (N_8310,N_8183,N_8189);
and U8311 (N_8311,N_8116,N_8073);
xor U8312 (N_8312,N_8011,N_8149);
or U8313 (N_8313,N_8176,N_8033);
nor U8314 (N_8314,N_8194,N_8079);
nor U8315 (N_8315,N_8082,N_8173);
and U8316 (N_8316,N_8134,N_8064);
and U8317 (N_8317,N_8169,N_8183);
nand U8318 (N_8318,N_8011,N_8135);
and U8319 (N_8319,N_8045,N_8130);
or U8320 (N_8320,N_8145,N_8110);
nor U8321 (N_8321,N_8143,N_8055);
and U8322 (N_8322,N_8071,N_8133);
and U8323 (N_8323,N_8024,N_8183);
nor U8324 (N_8324,N_8118,N_8089);
nand U8325 (N_8325,N_8123,N_8011);
nor U8326 (N_8326,N_8141,N_8030);
or U8327 (N_8327,N_8140,N_8197);
nor U8328 (N_8328,N_8176,N_8066);
and U8329 (N_8329,N_8182,N_8090);
or U8330 (N_8330,N_8096,N_8029);
nand U8331 (N_8331,N_8015,N_8009);
xnor U8332 (N_8332,N_8153,N_8064);
xor U8333 (N_8333,N_8168,N_8053);
xnor U8334 (N_8334,N_8143,N_8002);
or U8335 (N_8335,N_8026,N_8066);
or U8336 (N_8336,N_8025,N_8084);
nor U8337 (N_8337,N_8157,N_8004);
xor U8338 (N_8338,N_8023,N_8064);
nand U8339 (N_8339,N_8172,N_8128);
and U8340 (N_8340,N_8080,N_8013);
nand U8341 (N_8341,N_8150,N_8108);
or U8342 (N_8342,N_8142,N_8108);
or U8343 (N_8343,N_8003,N_8109);
nand U8344 (N_8344,N_8015,N_8068);
xor U8345 (N_8345,N_8188,N_8136);
or U8346 (N_8346,N_8060,N_8156);
nor U8347 (N_8347,N_8084,N_8105);
xor U8348 (N_8348,N_8079,N_8100);
or U8349 (N_8349,N_8072,N_8025);
and U8350 (N_8350,N_8163,N_8043);
xnor U8351 (N_8351,N_8136,N_8079);
nor U8352 (N_8352,N_8146,N_8178);
nor U8353 (N_8353,N_8060,N_8103);
xnor U8354 (N_8354,N_8150,N_8071);
or U8355 (N_8355,N_8029,N_8147);
or U8356 (N_8356,N_8092,N_8180);
nand U8357 (N_8357,N_8081,N_8160);
nand U8358 (N_8358,N_8033,N_8145);
and U8359 (N_8359,N_8198,N_8053);
nand U8360 (N_8360,N_8158,N_8142);
or U8361 (N_8361,N_8148,N_8018);
nand U8362 (N_8362,N_8008,N_8157);
and U8363 (N_8363,N_8003,N_8029);
or U8364 (N_8364,N_8001,N_8010);
xor U8365 (N_8365,N_8117,N_8064);
nand U8366 (N_8366,N_8001,N_8189);
or U8367 (N_8367,N_8051,N_8093);
or U8368 (N_8368,N_8007,N_8111);
nand U8369 (N_8369,N_8120,N_8038);
xnor U8370 (N_8370,N_8094,N_8101);
xor U8371 (N_8371,N_8041,N_8083);
xor U8372 (N_8372,N_8121,N_8044);
xnor U8373 (N_8373,N_8062,N_8059);
or U8374 (N_8374,N_8166,N_8074);
xor U8375 (N_8375,N_8017,N_8158);
xor U8376 (N_8376,N_8078,N_8032);
nor U8377 (N_8377,N_8030,N_8054);
xor U8378 (N_8378,N_8173,N_8146);
nor U8379 (N_8379,N_8046,N_8149);
and U8380 (N_8380,N_8002,N_8052);
nand U8381 (N_8381,N_8160,N_8146);
nand U8382 (N_8382,N_8184,N_8167);
xor U8383 (N_8383,N_8149,N_8120);
and U8384 (N_8384,N_8130,N_8007);
or U8385 (N_8385,N_8056,N_8003);
nor U8386 (N_8386,N_8185,N_8153);
nand U8387 (N_8387,N_8154,N_8083);
or U8388 (N_8388,N_8148,N_8054);
or U8389 (N_8389,N_8118,N_8140);
or U8390 (N_8390,N_8126,N_8112);
nand U8391 (N_8391,N_8003,N_8131);
or U8392 (N_8392,N_8057,N_8054);
nand U8393 (N_8393,N_8169,N_8035);
xnor U8394 (N_8394,N_8159,N_8148);
nand U8395 (N_8395,N_8113,N_8002);
or U8396 (N_8396,N_8090,N_8027);
nand U8397 (N_8397,N_8083,N_8071);
or U8398 (N_8398,N_8098,N_8096);
and U8399 (N_8399,N_8000,N_8188);
nand U8400 (N_8400,N_8200,N_8338);
and U8401 (N_8401,N_8318,N_8366);
nor U8402 (N_8402,N_8252,N_8357);
nand U8403 (N_8403,N_8327,N_8394);
or U8404 (N_8404,N_8364,N_8291);
or U8405 (N_8405,N_8323,N_8233);
nor U8406 (N_8406,N_8339,N_8363);
nor U8407 (N_8407,N_8345,N_8232);
nand U8408 (N_8408,N_8230,N_8287);
nand U8409 (N_8409,N_8375,N_8313);
or U8410 (N_8410,N_8263,N_8242);
or U8411 (N_8411,N_8206,N_8373);
nor U8412 (N_8412,N_8332,N_8380);
or U8413 (N_8413,N_8308,N_8222);
nand U8414 (N_8414,N_8259,N_8255);
or U8415 (N_8415,N_8223,N_8274);
or U8416 (N_8416,N_8271,N_8336);
xor U8417 (N_8417,N_8299,N_8306);
xnor U8418 (N_8418,N_8254,N_8387);
xnor U8419 (N_8419,N_8326,N_8335);
nor U8420 (N_8420,N_8353,N_8283);
xnor U8421 (N_8421,N_8304,N_8293);
nor U8422 (N_8422,N_8292,N_8272);
nand U8423 (N_8423,N_8212,N_8214);
or U8424 (N_8424,N_8302,N_8238);
nand U8425 (N_8425,N_8205,N_8378);
nor U8426 (N_8426,N_8239,N_8278);
and U8427 (N_8427,N_8286,N_8359);
and U8428 (N_8428,N_8248,N_8325);
and U8429 (N_8429,N_8307,N_8265);
nor U8430 (N_8430,N_8352,N_8340);
nor U8431 (N_8431,N_8221,N_8280);
and U8432 (N_8432,N_8393,N_8386);
and U8433 (N_8433,N_8371,N_8321);
xnor U8434 (N_8434,N_8319,N_8273);
or U8435 (N_8435,N_8396,N_8243);
or U8436 (N_8436,N_8281,N_8389);
nand U8437 (N_8437,N_8354,N_8276);
or U8438 (N_8438,N_8294,N_8253);
or U8439 (N_8439,N_8365,N_8289);
nand U8440 (N_8440,N_8324,N_8368);
xnor U8441 (N_8441,N_8225,N_8210);
xnor U8442 (N_8442,N_8330,N_8303);
or U8443 (N_8443,N_8268,N_8329);
and U8444 (N_8444,N_8342,N_8370);
nand U8445 (N_8445,N_8297,N_8215);
nor U8446 (N_8446,N_8240,N_8337);
and U8447 (N_8447,N_8320,N_8282);
or U8448 (N_8448,N_8305,N_8213);
nor U8449 (N_8449,N_8229,N_8395);
and U8450 (N_8450,N_8256,N_8350);
xor U8451 (N_8451,N_8262,N_8250);
or U8452 (N_8452,N_8237,N_8360);
and U8453 (N_8453,N_8235,N_8257);
xnor U8454 (N_8454,N_8385,N_8367);
xor U8455 (N_8455,N_8301,N_8391);
xor U8456 (N_8456,N_8295,N_8203);
nor U8457 (N_8457,N_8201,N_8270);
or U8458 (N_8458,N_8290,N_8267);
or U8459 (N_8459,N_8346,N_8249);
or U8460 (N_8460,N_8236,N_8220);
or U8461 (N_8461,N_8241,N_8261);
nand U8462 (N_8462,N_8376,N_8316);
xnor U8463 (N_8463,N_8341,N_8382);
and U8464 (N_8464,N_8227,N_8343);
and U8465 (N_8465,N_8234,N_8349);
xnor U8466 (N_8466,N_8369,N_8298);
nand U8467 (N_8467,N_8275,N_8314);
or U8468 (N_8468,N_8355,N_8388);
nand U8469 (N_8469,N_8202,N_8269);
or U8470 (N_8470,N_8392,N_8296);
and U8471 (N_8471,N_8204,N_8361);
and U8472 (N_8472,N_8315,N_8399);
and U8473 (N_8473,N_8356,N_8217);
nand U8474 (N_8474,N_8383,N_8310);
nor U8475 (N_8475,N_8288,N_8266);
and U8476 (N_8476,N_8251,N_8208);
nor U8477 (N_8477,N_8300,N_8219);
nor U8478 (N_8478,N_8247,N_8351);
nand U8479 (N_8479,N_8284,N_8398);
nand U8480 (N_8480,N_8328,N_8231);
xor U8481 (N_8481,N_8379,N_8264);
or U8482 (N_8482,N_8216,N_8362);
nand U8483 (N_8483,N_8279,N_8344);
or U8484 (N_8484,N_8211,N_8333);
or U8485 (N_8485,N_8374,N_8244);
or U8486 (N_8486,N_8331,N_8384);
xnor U8487 (N_8487,N_8311,N_8218);
xor U8488 (N_8488,N_8277,N_8348);
nand U8489 (N_8489,N_8312,N_8358);
nor U8490 (N_8490,N_8245,N_8334);
nand U8491 (N_8491,N_8347,N_8309);
or U8492 (N_8492,N_8322,N_8390);
and U8493 (N_8493,N_8258,N_8285);
nor U8494 (N_8494,N_8397,N_8377);
and U8495 (N_8495,N_8372,N_8246);
xnor U8496 (N_8496,N_8207,N_8228);
or U8497 (N_8497,N_8381,N_8226);
xor U8498 (N_8498,N_8260,N_8224);
nand U8499 (N_8499,N_8317,N_8209);
or U8500 (N_8500,N_8267,N_8224);
nand U8501 (N_8501,N_8348,N_8300);
xnor U8502 (N_8502,N_8366,N_8271);
xnor U8503 (N_8503,N_8288,N_8273);
and U8504 (N_8504,N_8300,N_8390);
and U8505 (N_8505,N_8253,N_8380);
or U8506 (N_8506,N_8208,N_8332);
nor U8507 (N_8507,N_8297,N_8397);
nor U8508 (N_8508,N_8247,N_8226);
or U8509 (N_8509,N_8359,N_8308);
or U8510 (N_8510,N_8345,N_8348);
nand U8511 (N_8511,N_8217,N_8374);
nor U8512 (N_8512,N_8362,N_8337);
xnor U8513 (N_8513,N_8202,N_8320);
nand U8514 (N_8514,N_8266,N_8339);
or U8515 (N_8515,N_8351,N_8355);
nand U8516 (N_8516,N_8365,N_8320);
nor U8517 (N_8517,N_8281,N_8345);
or U8518 (N_8518,N_8313,N_8355);
or U8519 (N_8519,N_8389,N_8250);
nand U8520 (N_8520,N_8366,N_8254);
nor U8521 (N_8521,N_8389,N_8289);
xor U8522 (N_8522,N_8394,N_8320);
xor U8523 (N_8523,N_8295,N_8316);
and U8524 (N_8524,N_8249,N_8257);
nor U8525 (N_8525,N_8257,N_8361);
xor U8526 (N_8526,N_8371,N_8330);
xor U8527 (N_8527,N_8218,N_8344);
or U8528 (N_8528,N_8363,N_8221);
xnor U8529 (N_8529,N_8296,N_8328);
nor U8530 (N_8530,N_8396,N_8384);
nor U8531 (N_8531,N_8354,N_8280);
or U8532 (N_8532,N_8399,N_8262);
and U8533 (N_8533,N_8361,N_8381);
or U8534 (N_8534,N_8202,N_8261);
nand U8535 (N_8535,N_8340,N_8336);
and U8536 (N_8536,N_8380,N_8393);
nand U8537 (N_8537,N_8360,N_8349);
nand U8538 (N_8538,N_8249,N_8238);
nand U8539 (N_8539,N_8271,N_8209);
nor U8540 (N_8540,N_8269,N_8315);
nor U8541 (N_8541,N_8352,N_8365);
and U8542 (N_8542,N_8207,N_8200);
or U8543 (N_8543,N_8243,N_8264);
nand U8544 (N_8544,N_8330,N_8226);
nor U8545 (N_8545,N_8389,N_8265);
or U8546 (N_8546,N_8306,N_8241);
and U8547 (N_8547,N_8325,N_8245);
or U8548 (N_8548,N_8317,N_8285);
xor U8549 (N_8549,N_8258,N_8289);
xnor U8550 (N_8550,N_8374,N_8397);
nand U8551 (N_8551,N_8290,N_8368);
xnor U8552 (N_8552,N_8363,N_8373);
nand U8553 (N_8553,N_8371,N_8254);
and U8554 (N_8554,N_8251,N_8254);
or U8555 (N_8555,N_8370,N_8389);
nand U8556 (N_8556,N_8213,N_8231);
or U8557 (N_8557,N_8338,N_8354);
nand U8558 (N_8558,N_8203,N_8388);
and U8559 (N_8559,N_8250,N_8398);
or U8560 (N_8560,N_8300,N_8232);
nand U8561 (N_8561,N_8213,N_8208);
and U8562 (N_8562,N_8212,N_8216);
nor U8563 (N_8563,N_8381,N_8202);
nand U8564 (N_8564,N_8381,N_8287);
nor U8565 (N_8565,N_8336,N_8373);
nor U8566 (N_8566,N_8238,N_8307);
xor U8567 (N_8567,N_8217,N_8239);
nand U8568 (N_8568,N_8306,N_8319);
xnor U8569 (N_8569,N_8287,N_8356);
and U8570 (N_8570,N_8221,N_8342);
and U8571 (N_8571,N_8261,N_8327);
and U8572 (N_8572,N_8235,N_8269);
and U8573 (N_8573,N_8279,N_8274);
and U8574 (N_8574,N_8245,N_8252);
nor U8575 (N_8575,N_8213,N_8276);
nand U8576 (N_8576,N_8395,N_8398);
nand U8577 (N_8577,N_8298,N_8276);
nand U8578 (N_8578,N_8273,N_8337);
nor U8579 (N_8579,N_8352,N_8399);
and U8580 (N_8580,N_8220,N_8382);
xnor U8581 (N_8581,N_8390,N_8223);
nor U8582 (N_8582,N_8319,N_8240);
nand U8583 (N_8583,N_8295,N_8273);
xor U8584 (N_8584,N_8348,N_8389);
and U8585 (N_8585,N_8225,N_8354);
nor U8586 (N_8586,N_8392,N_8235);
xor U8587 (N_8587,N_8202,N_8286);
or U8588 (N_8588,N_8308,N_8337);
xor U8589 (N_8589,N_8245,N_8277);
or U8590 (N_8590,N_8259,N_8241);
xor U8591 (N_8591,N_8347,N_8317);
nor U8592 (N_8592,N_8321,N_8227);
and U8593 (N_8593,N_8261,N_8367);
nor U8594 (N_8594,N_8390,N_8316);
or U8595 (N_8595,N_8259,N_8337);
nand U8596 (N_8596,N_8308,N_8399);
or U8597 (N_8597,N_8303,N_8343);
xnor U8598 (N_8598,N_8290,N_8229);
nand U8599 (N_8599,N_8294,N_8243);
nor U8600 (N_8600,N_8439,N_8442);
or U8601 (N_8601,N_8473,N_8554);
and U8602 (N_8602,N_8425,N_8549);
and U8603 (N_8603,N_8577,N_8523);
nor U8604 (N_8604,N_8500,N_8487);
and U8605 (N_8605,N_8515,N_8597);
xnor U8606 (N_8606,N_8415,N_8548);
nand U8607 (N_8607,N_8513,N_8453);
xor U8608 (N_8608,N_8585,N_8519);
nor U8609 (N_8609,N_8593,N_8591);
nand U8610 (N_8610,N_8531,N_8480);
or U8611 (N_8611,N_8551,N_8509);
or U8612 (N_8612,N_8466,N_8405);
xnor U8613 (N_8613,N_8595,N_8403);
and U8614 (N_8614,N_8458,N_8502);
nand U8615 (N_8615,N_8534,N_8482);
or U8616 (N_8616,N_8481,N_8493);
or U8617 (N_8617,N_8556,N_8430);
and U8618 (N_8618,N_8573,N_8533);
and U8619 (N_8619,N_8579,N_8465);
xor U8620 (N_8620,N_8525,N_8555);
xor U8621 (N_8621,N_8567,N_8488);
nand U8622 (N_8622,N_8505,N_8566);
xor U8623 (N_8623,N_8431,N_8529);
and U8624 (N_8624,N_8535,N_8436);
or U8625 (N_8625,N_8448,N_8434);
and U8626 (N_8626,N_8572,N_8557);
nor U8627 (N_8627,N_8428,N_8569);
xnor U8628 (N_8628,N_8451,N_8552);
or U8629 (N_8629,N_8478,N_8537);
xor U8630 (N_8630,N_8543,N_8412);
nor U8631 (N_8631,N_8497,N_8524);
nor U8632 (N_8632,N_8401,N_8564);
and U8633 (N_8633,N_8475,N_8414);
xor U8634 (N_8634,N_8553,N_8514);
xnor U8635 (N_8635,N_8528,N_8459);
nand U8636 (N_8636,N_8558,N_8402);
nor U8637 (N_8637,N_8445,N_8446);
and U8638 (N_8638,N_8574,N_8449);
xor U8639 (N_8639,N_8588,N_8545);
and U8640 (N_8640,N_8450,N_8501);
nor U8641 (N_8641,N_8507,N_8526);
nor U8642 (N_8642,N_8464,N_8594);
xnor U8643 (N_8643,N_8454,N_8580);
nor U8644 (N_8644,N_8444,N_8433);
or U8645 (N_8645,N_8489,N_8527);
and U8646 (N_8646,N_8438,N_8485);
and U8647 (N_8647,N_8592,N_8578);
nor U8648 (N_8648,N_8440,N_8492);
xnor U8649 (N_8649,N_8581,N_8472);
nand U8650 (N_8650,N_8499,N_8599);
or U8651 (N_8651,N_8544,N_8496);
xnor U8652 (N_8652,N_8484,N_8441);
and U8653 (N_8653,N_8469,N_8471);
nor U8654 (N_8654,N_8586,N_8421);
and U8655 (N_8655,N_8538,N_8536);
xor U8656 (N_8656,N_8483,N_8559);
xnor U8657 (N_8657,N_8568,N_8443);
nor U8658 (N_8658,N_8565,N_8511);
nor U8659 (N_8659,N_8530,N_8419);
and U8660 (N_8660,N_8495,N_8447);
or U8661 (N_8661,N_8463,N_8455);
nand U8662 (N_8662,N_8437,N_8486);
xnor U8663 (N_8663,N_8432,N_8409);
and U8664 (N_8664,N_8503,N_8418);
or U8665 (N_8665,N_8521,N_8498);
nand U8666 (N_8666,N_8476,N_8490);
or U8667 (N_8667,N_8512,N_8504);
xnor U8668 (N_8668,N_8570,N_8456);
xnor U8669 (N_8669,N_8510,N_8470);
and U8670 (N_8670,N_8462,N_8474);
xor U8671 (N_8671,N_8479,N_8406);
nand U8672 (N_8672,N_8540,N_8452);
and U8673 (N_8673,N_8584,N_8461);
or U8674 (N_8674,N_8420,N_8571);
xor U8675 (N_8675,N_8541,N_8516);
xor U8676 (N_8676,N_8435,N_8561);
and U8677 (N_8677,N_8491,N_8598);
nor U8678 (N_8678,N_8583,N_8422);
and U8679 (N_8679,N_8427,N_8457);
nand U8680 (N_8680,N_8575,N_8589);
and U8681 (N_8681,N_8407,N_8404);
nand U8682 (N_8682,N_8517,N_8429);
nand U8683 (N_8683,N_8423,N_8546);
or U8684 (N_8684,N_8410,N_8596);
xnor U8685 (N_8685,N_8550,N_8468);
nor U8686 (N_8686,N_8408,N_8522);
xnor U8687 (N_8687,N_8411,N_8518);
xnor U8688 (N_8688,N_8426,N_8520);
or U8689 (N_8689,N_8590,N_8547);
xnor U8690 (N_8690,N_8560,N_8467);
or U8691 (N_8691,N_8587,N_8582);
xnor U8692 (N_8692,N_8539,N_8506);
or U8693 (N_8693,N_8494,N_8413);
nor U8694 (N_8694,N_8417,N_8416);
nor U8695 (N_8695,N_8542,N_8562);
or U8696 (N_8696,N_8460,N_8576);
nor U8697 (N_8697,N_8508,N_8563);
xor U8698 (N_8698,N_8477,N_8400);
nand U8699 (N_8699,N_8424,N_8532);
xnor U8700 (N_8700,N_8483,N_8475);
or U8701 (N_8701,N_8411,N_8558);
xor U8702 (N_8702,N_8435,N_8418);
or U8703 (N_8703,N_8433,N_8453);
xor U8704 (N_8704,N_8484,N_8581);
xor U8705 (N_8705,N_8442,N_8467);
or U8706 (N_8706,N_8414,N_8532);
xor U8707 (N_8707,N_8400,N_8430);
xor U8708 (N_8708,N_8467,N_8589);
or U8709 (N_8709,N_8598,N_8522);
and U8710 (N_8710,N_8562,N_8422);
nand U8711 (N_8711,N_8564,N_8435);
nor U8712 (N_8712,N_8439,N_8561);
or U8713 (N_8713,N_8465,N_8580);
xnor U8714 (N_8714,N_8501,N_8468);
nor U8715 (N_8715,N_8585,N_8446);
or U8716 (N_8716,N_8558,N_8442);
or U8717 (N_8717,N_8448,N_8483);
and U8718 (N_8718,N_8491,N_8411);
or U8719 (N_8719,N_8485,N_8459);
or U8720 (N_8720,N_8437,N_8588);
nand U8721 (N_8721,N_8524,N_8479);
xnor U8722 (N_8722,N_8485,N_8580);
nand U8723 (N_8723,N_8504,N_8534);
or U8724 (N_8724,N_8473,N_8442);
xor U8725 (N_8725,N_8413,N_8441);
xor U8726 (N_8726,N_8435,N_8424);
nor U8727 (N_8727,N_8425,N_8573);
nor U8728 (N_8728,N_8450,N_8511);
or U8729 (N_8729,N_8457,N_8454);
or U8730 (N_8730,N_8584,N_8455);
or U8731 (N_8731,N_8454,N_8434);
nor U8732 (N_8732,N_8580,N_8416);
xnor U8733 (N_8733,N_8467,N_8502);
nand U8734 (N_8734,N_8501,N_8414);
nor U8735 (N_8735,N_8550,N_8539);
nand U8736 (N_8736,N_8567,N_8400);
and U8737 (N_8737,N_8582,N_8506);
and U8738 (N_8738,N_8439,N_8412);
xnor U8739 (N_8739,N_8565,N_8536);
xnor U8740 (N_8740,N_8426,N_8553);
or U8741 (N_8741,N_8524,N_8409);
nor U8742 (N_8742,N_8440,N_8503);
xor U8743 (N_8743,N_8439,N_8512);
nand U8744 (N_8744,N_8488,N_8484);
xnor U8745 (N_8745,N_8400,N_8442);
and U8746 (N_8746,N_8457,N_8506);
or U8747 (N_8747,N_8561,N_8575);
and U8748 (N_8748,N_8536,N_8408);
nor U8749 (N_8749,N_8575,N_8551);
nor U8750 (N_8750,N_8525,N_8439);
xnor U8751 (N_8751,N_8422,N_8538);
or U8752 (N_8752,N_8475,N_8530);
nand U8753 (N_8753,N_8498,N_8524);
xor U8754 (N_8754,N_8567,N_8497);
or U8755 (N_8755,N_8420,N_8502);
and U8756 (N_8756,N_8503,N_8424);
nor U8757 (N_8757,N_8530,N_8527);
or U8758 (N_8758,N_8520,N_8566);
and U8759 (N_8759,N_8426,N_8579);
nand U8760 (N_8760,N_8474,N_8432);
and U8761 (N_8761,N_8596,N_8425);
nor U8762 (N_8762,N_8458,N_8549);
and U8763 (N_8763,N_8553,N_8503);
xor U8764 (N_8764,N_8592,N_8448);
nand U8765 (N_8765,N_8549,N_8597);
xnor U8766 (N_8766,N_8444,N_8515);
xnor U8767 (N_8767,N_8527,N_8410);
nand U8768 (N_8768,N_8429,N_8436);
or U8769 (N_8769,N_8436,N_8512);
xor U8770 (N_8770,N_8568,N_8419);
nor U8771 (N_8771,N_8409,N_8405);
nor U8772 (N_8772,N_8517,N_8457);
and U8773 (N_8773,N_8425,N_8597);
and U8774 (N_8774,N_8424,N_8582);
or U8775 (N_8775,N_8442,N_8409);
nor U8776 (N_8776,N_8577,N_8512);
and U8777 (N_8777,N_8503,N_8467);
xor U8778 (N_8778,N_8432,N_8500);
and U8779 (N_8779,N_8518,N_8584);
or U8780 (N_8780,N_8562,N_8593);
and U8781 (N_8781,N_8421,N_8536);
nand U8782 (N_8782,N_8509,N_8514);
xor U8783 (N_8783,N_8440,N_8589);
or U8784 (N_8784,N_8410,N_8413);
nand U8785 (N_8785,N_8445,N_8574);
xor U8786 (N_8786,N_8519,N_8425);
xnor U8787 (N_8787,N_8547,N_8548);
nor U8788 (N_8788,N_8489,N_8566);
and U8789 (N_8789,N_8498,N_8575);
or U8790 (N_8790,N_8450,N_8417);
and U8791 (N_8791,N_8432,N_8562);
nand U8792 (N_8792,N_8509,N_8538);
xnor U8793 (N_8793,N_8533,N_8461);
nor U8794 (N_8794,N_8526,N_8496);
nand U8795 (N_8795,N_8423,N_8441);
xor U8796 (N_8796,N_8487,N_8499);
nor U8797 (N_8797,N_8418,N_8431);
and U8798 (N_8798,N_8524,N_8552);
or U8799 (N_8799,N_8566,N_8567);
xor U8800 (N_8800,N_8626,N_8758);
nand U8801 (N_8801,N_8637,N_8622);
and U8802 (N_8802,N_8633,N_8649);
nor U8803 (N_8803,N_8636,N_8690);
nor U8804 (N_8804,N_8785,N_8739);
and U8805 (N_8805,N_8604,N_8650);
nor U8806 (N_8806,N_8621,N_8699);
nand U8807 (N_8807,N_8673,N_8760);
and U8808 (N_8808,N_8679,N_8705);
or U8809 (N_8809,N_8600,N_8668);
or U8810 (N_8810,N_8646,N_8745);
nor U8811 (N_8811,N_8607,N_8769);
nand U8812 (N_8812,N_8770,N_8789);
xnor U8813 (N_8813,N_8714,N_8670);
nand U8814 (N_8814,N_8677,N_8783);
xor U8815 (N_8815,N_8721,N_8779);
xnor U8816 (N_8816,N_8795,N_8708);
xnor U8817 (N_8817,N_8755,N_8618);
nand U8818 (N_8818,N_8645,N_8704);
and U8819 (N_8819,N_8691,N_8609);
and U8820 (N_8820,N_8759,N_8630);
and U8821 (N_8821,N_8615,N_8632);
nand U8822 (N_8822,N_8778,N_8667);
or U8823 (N_8823,N_8792,N_8753);
nor U8824 (N_8824,N_8798,N_8654);
nand U8825 (N_8825,N_8711,N_8735);
and U8826 (N_8826,N_8659,N_8794);
xor U8827 (N_8827,N_8611,N_8757);
nand U8828 (N_8828,N_8723,N_8742);
nor U8829 (N_8829,N_8702,N_8661);
or U8830 (N_8830,N_8799,N_8703);
or U8831 (N_8831,N_8692,N_8734);
and U8832 (N_8832,N_8719,N_8655);
and U8833 (N_8833,N_8675,N_8698);
or U8834 (N_8834,N_8652,N_8602);
xor U8835 (N_8835,N_8762,N_8674);
nand U8836 (N_8836,N_8763,N_8747);
and U8837 (N_8837,N_8623,N_8644);
or U8838 (N_8838,N_8712,N_8641);
and U8839 (N_8839,N_8638,N_8730);
or U8840 (N_8840,N_8606,N_8766);
xnor U8841 (N_8841,N_8726,N_8696);
nand U8842 (N_8842,N_8715,N_8648);
xor U8843 (N_8843,N_8631,N_8693);
nor U8844 (N_8844,N_8685,N_8660);
or U8845 (N_8845,N_8743,N_8634);
and U8846 (N_8846,N_8748,N_8643);
and U8847 (N_8847,N_8788,N_8780);
nor U8848 (N_8848,N_8772,N_8790);
nand U8849 (N_8849,N_8706,N_8603);
nand U8850 (N_8850,N_8737,N_8687);
and U8851 (N_8851,N_8786,N_8664);
nand U8852 (N_8852,N_8671,N_8700);
xnor U8853 (N_8853,N_8680,N_8776);
nand U8854 (N_8854,N_8695,N_8710);
nand U8855 (N_8855,N_8731,N_8740);
nand U8856 (N_8856,N_8665,N_8746);
nor U8857 (N_8857,N_8686,N_8732);
or U8858 (N_8858,N_8754,N_8777);
xnor U8859 (N_8859,N_8752,N_8716);
nor U8860 (N_8860,N_8647,N_8640);
nand U8861 (N_8861,N_8744,N_8749);
nand U8862 (N_8862,N_8628,N_8771);
xnor U8863 (N_8863,N_8656,N_8727);
nand U8864 (N_8864,N_8681,N_8773);
and U8865 (N_8865,N_8793,N_8614);
or U8866 (N_8866,N_8796,N_8733);
and U8867 (N_8867,N_8717,N_8782);
and U8868 (N_8868,N_8768,N_8718);
nor U8869 (N_8869,N_8639,N_8750);
or U8870 (N_8870,N_8775,N_8774);
xnor U8871 (N_8871,N_8713,N_8608);
nand U8872 (N_8872,N_8694,N_8765);
nand U8873 (N_8873,N_8738,N_8625);
nand U8874 (N_8874,N_8624,N_8651);
nor U8875 (N_8875,N_8657,N_8797);
or U8876 (N_8876,N_8627,N_8707);
or U8877 (N_8877,N_8761,N_8613);
nand U8878 (N_8878,N_8689,N_8764);
and U8879 (N_8879,N_8620,N_8605);
and U8880 (N_8880,N_8709,N_8781);
nor U8881 (N_8881,N_8672,N_8662);
and U8882 (N_8882,N_8683,N_8725);
or U8883 (N_8883,N_8617,N_8724);
and U8884 (N_8884,N_8658,N_8666);
xnor U8885 (N_8885,N_8756,N_8619);
xor U8886 (N_8886,N_8663,N_8601);
and U8887 (N_8887,N_8791,N_8767);
nor U8888 (N_8888,N_8697,N_8642);
nor U8889 (N_8889,N_8610,N_8682);
nand U8890 (N_8890,N_8635,N_8728);
nor U8891 (N_8891,N_8736,N_8676);
and U8892 (N_8892,N_8629,N_8701);
nand U8893 (N_8893,N_8741,N_8616);
xnor U8894 (N_8894,N_8612,N_8784);
nand U8895 (N_8895,N_8722,N_8729);
nor U8896 (N_8896,N_8678,N_8684);
or U8897 (N_8897,N_8653,N_8669);
or U8898 (N_8898,N_8720,N_8787);
xnor U8899 (N_8899,N_8751,N_8688);
and U8900 (N_8900,N_8653,N_8607);
nor U8901 (N_8901,N_8607,N_8721);
nor U8902 (N_8902,N_8644,N_8646);
nand U8903 (N_8903,N_8679,N_8608);
nor U8904 (N_8904,N_8670,N_8656);
nand U8905 (N_8905,N_8738,N_8706);
or U8906 (N_8906,N_8617,N_8685);
nor U8907 (N_8907,N_8733,N_8621);
nand U8908 (N_8908,N_8799,N_8680);
and U8909 (N_8909,N_8664,N_8600);
and U8910 (N_8910,N_8749,N_8605);
nand U8911 (N_8911,N_8756,N_8695);
nor U8912 (N_8912,N_8664,N_8794);
nand U8913 (N_8913,N_8613,N_8656);
nand U8914 (N_8914,N_8689,N_8791);
nor U8915 (N_8915,N_8641,N_8668);
xnor U8916 (N_8916,N_8648,N_8789);
nand U8917 (N_8917,N_8661,N_8740);
or U8918 (N_8918,N_8673,N_8717);
or U8919 (N_8919,N_8622,N_8785);
xnor U8920 (N_8920,N_8683,N_8733);
or U8921 (N_8921,N_8737,N_8717);
or U8922 (N_8922,N_8715,N_8719);
nor U8923 (N_8923,N_8770,N_8688);
or U8924 (N_8924,N_8648,N_8773);
or U8925 (N_8925,N_8721,N_8650);
nor U8926 (N_8926,N_8668,N_8626);
nand U8927 (N_8927,N_8702,N_8777);
xnor U8928 (N_8928,N_8712,N_8758);
nand U8929 (N_8929,N_8676,N_8767);
and U8930 (N_8930,N_8785,N_8790);
xnor U8931 (N_8931,N_8750,N_8771);
nand U8932 (N_8932,N_8616,N_8788);
xor U8933 (N_8933,N_8696,N_8690);
and U8934 (N_8934,N_8608,N_8781);
nand U8935 (N_8935,N_8603,N_8715);
nand U8936 (N_8936,N_8703,N_8787);
and U8937 (N_8937,N_8603,N_8726);
xnor U8938 (N_8938,N_8640,N_8791);
and U8939 (N_8939,N_8751,N_8735);
or U8940 (N_8940,N_8745,N_8628);
nand U8941 (N_8941,N_8751,N_8626);
or U8942 (N_8942,N_8648,N_8786);
nand U8943 (N_8943,N_8693,N_8682);
nand U8944 (N_8944,N_8673,N_8709);
or U8945 (N_8945,N_8688,N_8631);
and U8946 (N_8946,N_8667,N_8780);
and U8947 (N_8947,N_8675,N_8656);
and U8948 (N_8948,N_8728,N_8634);
nor U8949 (N_8949,N_8642,N_8726);
and U8950 (N_8950,N_8705,N_8681);
nor U8951 (N_8951,N_8632,N_8685);
or U8952 (N_8952,N_8713,N_8710);
nand U8953 (N_8953,N_8764,N_8725);
and U8954 (N_8954,N_8618,N_8715);
or U8955 (N_8955,N_8604,N_8671);
or U8956 (N_8956,N_8639,N_8679);
nand U8957 (N_8957,N_8799,N_8626);
nor U8958 (N_8958,N_8749,N_8654);
and U8959 (N_8959,N_8617,N_8757);
or U8960 (N_8960,N_8637,N_8692);
and U8961 (N_8961,N_8772,N_8722);
nor U8962 (N_8962,N_8788,N_8704);
or U8963 (N_8963,N_8630,N_8670);
and U8964 (N_8964,N_8620,N_8679);
nand U8965 (N_8965,N_8693,N_8730);
or U8966 (N_8966,N_8612,N_8788);
xor U8967 (N_8967,N_8641,N_8783);
and U8968 (N_8968,N_8761,N_8638);
and U8969 (N_8969,N_8799,N_8739);
and U8970 (N_8970,N_8758,N_8752);
and U8971 (N_8971,N_8677,N_8666);
nor U8972 (N_8972,N_8787,N_8789);
nor U8973 (N_8973,N_8785,N_8781);
or U8974 (N_8974,N_8642,N_8730);
and U8975 (N_8975,N_8645,N_8739);
nand U8976 (N_8976,N_8646,N_8713);
nor U8977 (N_8977,N_8616,N_8670);
and U8978 (N_8978,N_8644,N_8609);
or U8979 (N_8979,N_8616,N_8793);
or U8980 (N_8980,N_8773,N_8600);
nor U8981 (N_8981,N_8670,N_8742);
xor U8982 (N_8982,N_8624,N_8616);
nor U8983 (N_8983,N_8604,N_8796);
or U8984 (N_8984,N_8779,N_8638);
and U8985 (N_8985,N_8784,N_8742);
xor U8986 (N_8986,N_8607,N_8739);
or U8987 (N_8987,N_8660,N_8617);
nor U8988 (N_8988,N_8757,N_8770);
and U8989 (N_8989,N_8695,N_8602);
nor U8990 (N_8990,N_8688,N_8679);
nor U8991 (N_8991,N_8760,N_8719);
and U8992 (N_8992,N_8774,N_8618);
and U8993 (N_8993,N_8795,N_8601);
nand U8994 (N_8994,N_8796,N_8640);
or U8995 (N_8995,N_8772,N_8727);
or U8996 (N_8996,N_8640,N_8638);
nand U8997 (N_8997,N_8692,N_8600);
nand U8998 (N_8998,N_8622,N_8726);
xnor U8999 (N_8999,N_8761,N_8698);
xor U9000 (N_9000,N_8881,N_8975);
nand U9001 (N_9001,N_8913,N_8989);
nand U9002 (N_9002,N_8951,N_8803);
nor U9003 (N_9003,N_8812,N_8841);
xnor U9004 (N_9004,N_8979,N_8959);
or U9005 (N_9005,N_8946,N_8904);
and U9006 (N_9006,N_8875,N_8949);
or U9007 (N_9007,N_8825,N_8831);
nor U9008 (N_9008,N_8867,N_8856);
xnor U9009 (N_9009,N_8916,N_8935);
nand U9010 (N_9010,N_8871,N_8894);
or U9011 (N_9011,N_8837,N_8864);
xnor U9012 (N_9012,N_8983,N_8858);
and U9013 (N_9013,N_8836,N_8847);
nor U9014 (N_9014,N_8919,N_8879);
and U9015 (N_9015,N_8905,N_8948);
nand U9016 (N_9016,N_8990,N_8839);
and U9017 (N_9017,N_8971,N_8824);
and U9018 (N_9018,N_8911,N_8986);
nor U9019 (N_9019,N_8830,N_8827);
nor U9020 (N_9020,N_8941,N_8994);
xnor U9021 (N_9021,N_8802,N_8832);
nand U9022 (N_9022,N_8815,N_8886);
nand U9023 (N_9023,N_8902,N_8835);
nand U9024 (N_9024,N_8876,N_8929);
and U9025 (N_9025,N_8823,N_8923);
and U9026 (N_9026,N_8931,N_8819);
xnor U9027 (N_9027,N_8993,N_8906);
xor U9028 (N_9028,N_8992,N_8887);
or U9029 (N_9029,N_8954,N_8922);
or U9030 (N_9030,N_8897,N_8927);
and U9031 (N_9031,N_8901,N_8848);
nor U9032 (N_9032,N_8885,N_8842);
and U9033 (N_9033,N_8843,N_8991);
or U9034 (N_9034,N_8890,N_8960);
or U9035 (N_9035,N_8829,N_8899);
nand U9036 (N_9036,N_8855,N_8817);
or U9037 (N_9037,N_8809,N_8878);
and U9038 (N_9038,N_8840,N_8987);
nand U9039 (N_9039,N_8961,N_8888);
or U9040 (N_9040,N_8995,N_8883);
nor U9041 (N_9041,N_8988,N_8976);
nor U9042 (N_9042,N_8877,N_8972);
and U9043 (N_9043,N_8973,N_8985);
nand U9044 (N_9044,N_8943,N_8806);
nand U9045 (N_9045,N_8965,N_8914);
or U9046 (N_9046,N_8944,N_8999);
nor U9047 (N_9047,N_8964,N_8925);
xor U9048 (N_9048,N_8912,N_8918);
nand U9049 (N_9049,N_8953,N_8958);
nand U9050 (N_9050,N_8818,N_8863);
and U9051 (N_9051,N_8851,N_8850);
or U9052 (N_9052,N_8821,N_8966);
xor U9053 (N_9053,N_8908,N_8828);
nor U9054 (N_9054,N_8893,N_8945);
or U9055 (N_9055,N_8865,N_8822);
nand U9056 (N_9056,N_8816,N_8924);
or U9057 (N_9057,N_8873,N_8860);
xnor U9058 (N_9058,N_8869,N_8997);
or U9059 (N_9059,N_8955,N_8996);
nand U9060 (N_9060,N_8872,N_8981);
nor U9061 (N_9061,N_8920,N_8820);
xor U9062 (N_9062,N_8880,N_8882);
xnor U9063 (N_9063,N_8947,N_8942);
nand U9064 (N_9064,N_8852,N_8844);
or U9065 (N_9065,N_8956,N_8891);
nor U9066 (N_9066,N_8866,N_8853);
or U9067 (N_9067,N_8892,N_8967);
nor U9068 (N_9068,N_8940,N_8933);
xnor U9069 (N_9069,N_8810,N_8921);
or U9070 (N_9070,N_8910,N_8868);
nand U9071 (N_9071,N_8854,N_8898);
and U9072 (N_9072,N_8896,N_8811);
xnor U9073 (N_9073,N_8807,N_8861);
nand U9074 (N_9074,N_8982,N_8846);
nor U9075 (N_9075,N_8926,N_8978);
nor U9076 (N_9076,N_8909,N_8962);
nor U9077 (N_9077,N_8859,N_8814);
xnor U9078 (N_9078,N_8838,N_8862);
nor U9079 (N_9079,N_8968,N_8969);
nor U9080 (N_9080,N_8952,N_8800);
and U9081 (N_9081,N_8801,N_8804);
or U9082 (N_9082,N_8970,N_8833);
nor U9083 (N_9083,N_8903,N_8915);
nand U9084 (N_9084,N_8808,N_8984);
or U9085 (N_9085,N_8849,N_8937);
nor U9086 (N_9086,N_8977,N_8938);
xor U9087 (N_9087,N_8950,N_8805);
nor U9088 (N_9088,N_8998,N_8930);
xor U9089 (N_9089,N_8974,N_8963);
xor U9090 (N_9090,N_8857,N_8932);
and U9091 (N_9091,N_8845,N_8936);
nor U9092 (N_9092,N_8884,N_8870);
xnor U9093 (N_9093,N_8957,N_8826);
xnor U9094 (N_9094,N_8917,N_8928);
nor U9095 (N_9095,N_8889,N_8895);
or U9096 (N_9096,N_8900,N_8874);
and U9097 (N_9097,N_8907,N_8939);
or U9098 (N_9098,N_8834,N_8934);
xnor U9099 (N_9099,N_8980,N_8813);
xor U9100 (N_9100,N_8951,N_8990);
nor U9101 (N_9101,N_8823,N_8850);
xor U9102 (N_9102,N_8876,N_8884);
or U9103 (N_9103,N_8978,N_8843);
nor U9104 (N_9104,N_8948,N_8907);
nor U9105 (N_9105,N_8871,N_8872);
and U9106 (N_9106,N_8884,N_8893);
or U9107 (N_9107,N_8888,N_8956);
or U9108 (N_9108,N_8955,N_8849);
and U9109 (N_9109,N_8924,N_8981);
or U9110 (N_9110,N_8950,N_8825);
xor U9111 (N_9111,N_8892,N_8834);
or U9112 (N_9112,N_8939,N_8951);
nor U9113 (N_9113,N_8900,N_8944);
and U9114 (N_9114,N_8894,N_8956);
and U9115 (N_9115,N_8912,N_8853);
xor U9116 (N_9116,N_8852,N_8806);
nand U9117 (N_9117,N_8991,N_8942);
or U9118 (N_9118,N_8834,N_8911);
nor U9119 (N_9119,N_8949,N_8998);
and U9120 (N_9120,N_8852,N_8811);
and U9121 (N_9121,N_8802,N_8982);
nor U9122 (N_9122,N_8985,N_8882);
xnor U9123 (N_9123,N_8842,N_8972);
xnor U9124 (N_9124,N_8970,N_8939);
nor U9125 (N_9125,N_8881,N_8868);
nand U9126 (N_9126,N_8955,N_8991);
nor U9127 (N_9127,N_8992,N_8877);
nor U9128 (N_9128,N_8861,N_8958);
and U9129 (N_9129,N_8968,N_8813);
xnor U9130 (N_9130,N_8869,N_8881);
nand U9131 (N_9131,N_8986,N_8954);
and U9132 (N_9132,N_8908,N_8910);
nor U9133 (N_9133,N_8827,N_8987);
and U9134 (N_9134,N_8906,N_8811);
and U9135 (N_9135,N_8942,N_8822);
or U9136 (N_9136,N_8945,N_8927);
xnor U9137 (N_9137,N_8870,N_8880);
nor U9138 (N_9138,N_8917,N_8951);
xnor U9139 (N_9139,N_8903,N_8811);
or U9140 (N_9140,N_8918,N_8919);
nor U9141 (N_9141,N_8874,N_8924);
nor U9142 (N_9142,N_8818,N_8930);
nor U9143 (N_9143,N_8899,N_8916);
xnor U9144 (N_9144,N_8859,N_8874);
nor U9145 (N_9145,N_8859,N_8953);
and U9146 (N_9146,N_8950,N_8863);
xnor U9147 (N_9147,N_8865,N_8944);
nor U9148 (N_9148,N_8892,N_8846);
xnor U9149 (N_9149,N_8816,N_8851);
xor U9150 (N_9150,N_8954,N_8847);
or U9151 (N_9151,N_8947,N_8989);
nor U9152 (N_9152,N_8888,N_8804);
xnor U9153 (N_9153,N_8985,N_8896);
or U9154 (N_9154,N_8816,N_8870);
xor U9155 (N_9155,N_8899,N_8810);
xor U9156 (N_9156,N_8867,N_8855);
nor U9157 (N_9157,N_8856,N_8889);
nand U9158 (N_9158,N_8837,N_8829);
nor U9159 (N_9159,N_8947,N_8960);
xor U9160 (N_9160,N_8930,N_8936);
nor U9161 (N_9161,N_8993,N_8859);
nor U9162 (N_9162,N_8815,N_8889);
and U9163 (N_9163,N_8979,N_8892);
nor U9164 (N_9164,N_8818,N_8914);
xnor U9165 (N_9165,N_8816,N_8944);
or U9166 (N_9166,N_8991,N_8908);
nor U9167 (N_9167,N_8988,N_8982);
or U9168 (N_9168,N_8963,N_8873);
xor U9169 (N_9169,N_8846,N_8818);
nand U9170 (N_9170,N_8965,N_8812);
or U9171 (N_9171,N_8874,N_8864);
or U9172 (N_9172,N_8902,N_8939);
and U9173 (N_9173,N_8802,N_8968);
xor U9174 (N_9174,N_8949,N_8851);
nand U9175 (N_9175,N_8929,N_8954);
nor U9176 (N_9176,N_8825,N_8835);
nand U9177 (N_9177,N_8896,N_8812);
and U9178 (N_9178,N_8865,N_8975);
xnor U9179 (N_9179,N_8872,N_8939);
nor U9180 (N_9180,N_8904,N_8901);
nand U9181 (N_9181,N_8897,N_8969);
xnor U9182 (N_9182,N_8822,N_8925);
nand U9183 (N_9183,N_8988,N_8947);
xor U9184 (N_9184,N_8817,N_8813);
nor U9185 (N_9185,N_8801,N_8993);
xor U9186 (N_9186,N_8963,N_8938);
xnor U9187 (N_9187,N_8851,N_8866);
xnor U9188 (N_9188,N_8836,N_8917);
and U9189 (N_9189,N_8840,N_8966);
nor U9190 (N_9190,N_8868,N_8815);
xor U9191 (N_9191,N_8935,N_8979);
or U9192 (N_9192,N_8961,N_8831);
or U9193 (N_9193,N_8888,N_8865);
or U9194 (N_9194,N_8897,N_8965);
xor U9195 (N_9195,N_8856,N_8979);
or U9196 (N_9196,N_8886,N_8948);
nand U9197 (N_9197,N_8898,N_8892);
xnor U9198 (N_9198,N_8864,N_8883);
and U9199 (N_9199,N_8822,N_8819);
or U9200 (N_9200,N_9167,N_9025);
or U9201 (N_9201,N_9175,N_9002);
or U9202 (N_9202,N_9178,N_9046);
nand U9203 (N_9203,N_9019,N_9003);
xor U9204 (N_9204,N_9101,N_9068);
or U9205 (N_9205,N_9181,N_9058);
xor U9206 (N_9206,N_9157,N_9054);
nor U9207 (N_9207,N_9116,N_9090);
or U9208 (N_9208,N_9184,N_9111);
nand U9209 (N_9209,N_9089,N_9134);
nand U9210 (N_9210,N_9166,N_9071);
nand U9211 (N_9211,N_9142,N_9149);
nand U9212 (N_9212,N_9044,N_9008);
nor U9213 (N_9213,N_9107,N_9189);
and U9214 (N_9214,N_9183,N_9159);
and U9215 (N_9215,N_9162,N_9145);
or U9216 (N_9216,N_9047,N_9093);
or U9217 (N_9217,N_9153,N_9196);
nor U9218 (N_9218,N_9198,N_9027);
and U9219 (N_9219,N_9126,N_9190);
xor U9220 (N_9220,N_9079,N_9000);
xor U9221 (N_9221,N_9085,N_9033);
or U9222 (N_9222,N_9004,N_9014);
xnor U9223 (N_9223,N_9173,N_9154);
and U9224 (N_9224,N_9199,N_9006);
and U9225 (N_9225,N_9034,N_9036);
and U9226 (N_9226,N_9032,N_9061);
and U9227 (N_9227,N_9031,N_9059);
nor U9228 (N_9228,N_9050,N_9092);
nor U9229 (N_9229,N_9007,N_9103);
and U9230 (N_9230,N_9038,N_9155);
xnor U9231 (N_9231,N_9146,N_9094);
xor U9232 (N_9232,N_9096,N_9125);
nand U9233 (N_9233,N_9077,N_9188);
nand U9234 (N_9234,N_9057,N_9066);
or U9235 (N_9235,N_9122,N_9087);
or U9236 (N_9236,N_9164,N_9078);
and U9237 (N_9237,N_9072,N_9193);
or U9238 (N_9238,N_9192,N_9040);
nor U9239 (N_9239,N_9049,N_9098);
xnor U9240 (N_9240,N_9091,N_9097);
nand U9241 (N_9241,N_9165,N_9115);
and U9242 (N_9242,N_9023,N_9135);
nor U9243 (N_9243,N_9130,N_9106);
or U9244 (N_9244,N_9185,N_9124);
nor U9245 (N_9245,N_9132,N_9052);
xnor U9246 (N_9246,N_9172,N_9139);
xnor U9247 (N_9247,N_9011,N_9104);
and U9248 (N_9248,N_9114,N_9037);
nand U9249 (N_9249,N_9070,N_9067);
and U9250 (N_9250,N_9084,N_9076);
nor U9251 (N_9251,N_9156,N_9075);
nand U9252 (N_9252,N_9169,N_9062);
and U9253 (N_9253,N_9194,N_9133);
or U9254 (N_9254,N_9137,N_9105);
nand U9255 (N_9255,N_9051,N_9024);
nand U9256 (N_9256,N_9021,N_9191);
nand U9257 (N_9257,N_9095,N_9118);
and U9258 (N_9258,N_9144,N_9174);
xnor U9259 (N_9259,N_9069,N_9171);
nor U9260 (N_9260,N_9112,N_9120);
or U9261 (N_9261,N_9158,N_9029);
or U9262 (N_9262,N_9138,N_9168);
nand U9263 (N_9263,N_9005,N_9151);
xor U9264 (N_9264,N_9053,N_9017);
nor U9265 (N_9265,N_9110,N_9088);
xor U9266 (N_9266,N_9015,N_9018);
nor U9267 (N_9267,N_9176,N_9086);
nor U9268 (N_9268,N_9020,N_9186);
xnor U9269 (N_9269,N_9082,N_9197);
or U9270 (N_9270,N_9009,N_9143);
and U9271 (N_9271,N_9128,N_9163);
xnor U9272 (N_9272,N_9045,N_9182);
xor U9273 (N_9273,N_9141,N_9148);
xor U9274 (N_9274,N_9043,N_9041);
xor U9275 (N_9275,N_9195,N_9180);
or U9276 (N_9276,N_9160,N_9056);
nand U9277 (N_9277,N_9109,N_9039);
nor U9278 (N_9278,N_9147,N_9010);
nand U9279 (N_9279,N_9129,N_9055);
or U9280 (N_9280,N_9042,N_9127);
nor U9281 (N_9281,N_9035,N_9022);
or U9282 (N_9282,N_9119,N_9030);
nor U9283 (N_9283,N_9177,N_9100);
or U9284 (N_9284,N_9016,N_9108);
xor U9285 (N_9285,N_9048,N_9099);
and U9286 (N_9286,N_9187,N_9131);
nand U9287 (N_9287,N_9170,N_9063);
xor U9288 (N_9288,N_9073,N_9028);
and U9289 (N_9289,N_9179,N_9080);
nor U9290 (N_9290,N_9113,N_9001);
nand U9291 (N_9291,N_9081,N_9140);
and U9292 (N_9292,N_9060,N_9065);
nor U9293 (N_9293,N_9026,N_9136);
and U9294 (N_9294,N_9123,N_9117);
nor U9295 (N_9295,N_9161,N_9150);
or U9296 (N_9296,N_9012,N_9102);
xor U9297 (N_9297,N_9074,N_9083);
nand U9298 (N_9298,N_9152,N_9064);
or U9299 (N_9299,N_9013,N_9121);
and U9300 (N_9300,N_9067,N_9164);
xor U9301 (N_9301,N_9139,N_9177);
nand U9302 (N_9302,N_9116,N_9170);
nor U9303 (N_9303,N_9018,N_9043);
nand U9304 (N_9304,N_9023,N_9168);
and U9305 (N_9305,N_9079,N_9173);
nand U9306 (N_9306,N_9104,N_9134);
nand U9307 (N_9307,N_9195,N_9057);
or U9308 (N_9308,N_9079,N_9129);
or U9309 (N_9309,N_9056,N_9119);
and U9310 (N_9310,N_9104,N_9112);
nand U9311 (N_9311,N_9001,N_9132);
nor U9312 (N_9312,N_9038,N_9093);
nand U9313 (N_9313,N_9116,N_9110);
or U9314 (N_9314,N_9156,N_9132);
nor U9315 (N_9315,N_9114,N_9101);
nand U9316 (N_9316,N_9144,N_9083);
or U9317 (N_9317,N_9130,N_9101);
nor U9318 (N_9318,N_9031,N_9166);
xor U9319 (N_9319,N_9113,N_9025);
nand U9320 (N_9320,N_9082,N_9199);
or U9321 (N_9321,N_9017,N_9162);
and U9322 (N_9322,N_9100,N_9164);
xor U9323 (N_9323,N_9199,N_9018);
xnor U9324 (N_9324,N_9142,N_9184);
nand U9325 (N_9325,N_9190,N_9015);
nor U9326 (N_9326,N_9090,N_9162);
and U9327 (N_9327,N_9113,N_9156);
nand U9328 (N_9328,N_9131,N_9059);
nand U9329 (N_9329,N_9105,N_9168);
xor U9330 (N_9330,N_9051,N_9011);
and U9331 (N_9331,N_9184,N_9023);
or U9332 (N_9332,N_9106,N_9180);
nor U9333 (N_9333,N_9076,N_9188);
xor U9334 (N_9334,N_9107,N_9181);
nor U9335 (N_9335,N_9111,N_9158);
nand U9336 (N_9336,N_9135,N_9152);
and U9337 (N_9337,N_9079,N_9094);
nor U9338 (N_9338,N_9069,N_9087);
or U9339 (N_9339,N_9139,N_9127);
and U9340 (N_9340,N_9175,N_9179);
nand U9341 (N_9341,N_9041,N_9017);
xor U9342 (N_9342,N_9189,N_9039);
or U9343 (N_9343,N_9034,N_9171);
or U9344 (N_9344,N_9147,N_9121);
and U9345 (N_9345,N_9010,N_9105);
nor U9346 (N_9346,N_9192,N_9175);
and U9347 (N_9347,N_9158,N_9117);
or U9348 (N_9348,N_9072,N_9039);
nand U9349 (N_9349,N_9126,N_9162);
nand U9350 (N_9350,N_9006,N_9043);
and U9351 (N_9351,N_9165,N_9021);
nor U9352 (N_9352,N_9064,N_9188);
nor U9353 (N_9353,N_9072,N_9195);
or U9354 (N_9354,N_9006,N_9197);
nand U9355 (N_9355,N_9009,N_9010);
or U9356 (N_9356,N_9046,N_9119);
or U9357 (N_9357,N_9187,N_9135);
or U9358 (N_9358,N_9000,N_9177);
nand U9359 (N_9359,N_9108,N_9080);
and U9360 (N_9360,N_9156,N_9122);
and U9361 (N_9361,N_9028,N_9150);
nor U9362 (N_9362,N_9117,N_9196);
xor U9363 (N_9363,N_9123,N_9177);
and U9364 (N_9364,N_9043,N_9058);
nand U9365 (N_9365,N_9075,N_9121);
and U9366 (N_9366,N_9024,N_9136);
xor U9367 (N_9367,N_9055,N_9079);
nand U9368 (N_9368,N_9053,N_9099);
and U9369 (N_9369,N_9149,N_9170);
nand U9370 (N_9370,N_9090,N_9007);
xor U9371 (N_9371,N_9037,N_9025);
xnor U9372 (N_9372,N_9067,N_9182);
xor U9373 (N_9373,N_9090,N_9099);
and U9374 (N_9374,N_9174,N_9069);
xnor U9375 (N_9375,N_9104,N_9142);
xnor U9376 (N_9376,N_9003,N_9052);
nor U9377 (N_9377,N_9171,N_9043);
nand U9378 (N_9378,N_9150,N_9185);
xor U9379 (N_9379,N_9008,N_9031);
and U9380 (N_9380,N_9002,N_9141);
nor U9381 (N_9381,N_9007,N_9125);
xnor U9382 (N_9382,N_9082,N_9085);
xor U9383 (N_9383,N_9097,N_9059);
or U9384 (N_9384,N_9084,N_9060);
and U9385 (N_9385,N_9037,N_9078);
nand U9386 (N_9386,N_9150,N_9055);
nand U9387 (N_9387,N_9040,N_9139);
nand U9388 (N_9388,N_9065,N_9054);
and U9389 (N_9389,N_9024,N_9154);
nand U9390 (N_9390,N_9082,N_9136);
nor U9391 (N_9391,N_9054,N_9008);
and U9392 (N_9392,N_9134,N_9075);
or U9393 (N_9393,N_9166,N_9048);
and U9394 (N_9394,N_9197,N_9195);
or U9395 (N_9395,N_9112,N_9158);
and U9396 (N_9396,N_9098,N_9118);
or U9397 (N_9397,N_9171,N_9028);
xnor U9398 (N_9398,N_9000,N_9063);
nand U9399 (N_9399,N_9018,N_9116);
or U9400 (N_9400,N_9235,N_9275);
xnor U9401 (N_9401,N_9208,N_9319);
or U9402 (N_9402,N_9318,N_9306);
xnor U9403 (N_9403,N_9392,N_9343);
nand U9404 (N_9404,N_9227,N_9292);
nand U9405 (N_9405,N_9236,N_9379);
xor U9406 (N_9406,N_9320,N_9377);
or U9407 (N_9407,N_9255,N_9201);
xnor U9408 (N_9408,N_9209,N_9311);
xor U9409 (N_9409,N_9358,N_9220);
nand U9410 (N_9410,N_9229,N_9252);
xor U9411 (N_9411,N_9272,N_9370);
xnor U9412 (N_9412,N_9294,N_9291);
nand U9413 (N_9413,N_9317,N_9363);
nand U9414 (N_9414,N_9248,N_9212);
xnor U9415 (N_9415,N_9300,N_9387);
or U9416 (N_9416,N_9359,N_9205);
xnor U9417 (N_9417,N_9330,N_9265);
and U9418 (N_9418,N_9398,N_9224);
xnor U9419 (N_9419,N_9341,N_9380);
nand U9420 (N_9420,N_9213,N_9226);
nand U9421 (N_9421,N_9301,N_9378);
nor U9422 (N_9422,N_9242,N_9304);
nand U9423 (N_9423,N_9296,N_9207);
xor U9424 (N_9424,N_9303,N_9267);
nand U9425 (N_9425,N_9316,N_9218);
nand U9426 (N_9426,N_9222,N_9234);
and U9427 (N_9427,N_9225,N_9285);
nand U9428 (N_9428,N_9355,N_9271);
xnor U9429 (N_9429,N_9273,N_9257);
nor U9430 (N_9430,N_9269,N_9231);
or U9431 (N_9431,N_9356,N_9314);
nand U9432 (N_9432,N_9245,N_9324);
xnor U9433 (N_9433,N_9354,N_9390);
xor U9434 (N_9434,N_9366,N_9323);
nor U9435 (N_9435,N_9381,N_9263);
or U9436 (N_9436,N_9253,N_9282);
nand U9437 (N_9437,N_9289,N_9246);
nor U9438 (N_9438,N_9375,N_9206);
nand U9439 (N_9439,N_9388,N_9249);
nor U9440 (N_9440,N_9276,N_9260);
and U9441 (N_9441,N_9337,N_9277);
nand U9442 (N_9442,N_9335,N_9345);
xor U9443 (N_9443,N_9293,N_9254);
or U9444 (N_9444,N_9389,N_9279);
xnor U9445 (N_9445,N_9256,N_9351);
nor U9446 (N_9446,N_9262,N_9283);
or U9447 (N_9447,N_9384,N_9307);
nand U9448 (N_9448,N_9251,N_9210);
xor U9449 (N_9449,N_9346,N_9281);
xnor U9450 (N_9450,N_9393,N_9399);
xnor U9451 (N_9451,N_9340,N_9211);
nor U9452 (N_9452,N_9313,N_9237);
nor U9453 (N_9453,N_9362,N_9250);
and U9454 (N_9454,N_9348,N_9395);
xor U9455 (N_9455,N_9298,N_9396);
and U9456 (N_9456,N_9312,N_9299);
xor U9457 (N_9457,N_9374,N_9357);
and U9458 (N_9458,N_9350,N_9240);
and U9459 (N_9459,N_9243,N_9287);
or U9460 (N_9460,N_9328,N_9244);
nand U9461 (N_9461,N_9230,N_9365);
or U9462 (N_9462,N_9264,N_9325);
nor U9463 (N_9463,N_9247,N_9385);
and U9464 (N_9464,N_9332,N_9238);
and U9465 (N_9465,N_9368,N_9344);
nor U9466 (N_9466,N_9361,N_9373);
nand U9467 (N_9467,N_9367,N_9241);
xor U9468 (N_9468,N_9372,N_9309);
and U9469 (N_9469,N_9347,N_9394);
and U9470 (N_9470,N_9228,N_9302);
or U9471 (N_9471,N_9391,N_9329);
nand U9472 (N_9472,N_9203,N_9270);
or U9473 (N_9473,N_9214,N_9326);
or U9474 (N_9474,N_9295,N_9360);
nand U9475 (N_9475,N_9336,N_9315);
and U9476 (N_9476,N_9339,N_9278);
nand U9477 (N_9477,N_9288,N_9334);
xnor U9478 (N_9478,N_9280,N_9268);
nand U9479 (N_9479,N_9327,N_9386);
or U9480 (N_9480,N_9376,N_9219);
nor U9481 (N_9481,N_9371,N_9290);
xnor U9482 (N_9482,N_9383,N_9308);
nand U9483 (N_9483,N_9297,N_9305);
and U9484 (N_9484,N_9310,N_9233);
xor U9485 (N_9485,N_9331,N_9202);
and U9486 (N_9486,N_9239,N_9200);
nor U9487 (N_9487,N_9274,N_9322);
xnor U9488 (N_9488,N_9221,N_9333);
nand U9489 (N_9489,N_9352,N_9259);
or U9490 (N_9490,N_9382,N_9397);
nand U9491 (N_9491,N_9369,N_9266);
or U9492 (N_9492,N_9342,N_9353);
and U9493 (N_9493,N_9349,N_9258);
nor U9494 (N_9494,N_9232,N_9364);
or U9495 (N_9495,N_9284,N_9215);
xor U9496 (N_9496,N_9321,N_9286);
xnor U9497 (N_9497,N_9204,N_9338);
nor U9498 (N_9498,N_9261,N_9217);
and U9499 (N_9499,N_9223,N_9216);
nor U9500 (N_9500,N_9335,N_9339);
or U9501 (N_9501,N_9389,N_9222);
xor U9502 (N_9502,N_9351,N_9320);
xor U9503 (N_9503,N_9292,N_9279);
and U9504 (N_9504,N_9283,N_9264);
xor U9505 (N_9505,N_9301,N_9342);
xor U9506 (N_9506,N_9396,N_9370);
or U9507 (N_9507,N_9264,N_9287);
xnor U9508 (N_9508,N_9301,N_9260);
nand U9509 (N_9509,N_9353,N_9220);
nand U9510 (N_9510,N_9223,N_9342);
and U9511 (N_9511,N_9377,N_9244);
and U9512 (N_9512,N_9378,N_9209);
xor U9513 (N_9513,N_9366,N_9227);
and U9514 (N_9514,N_9278,N_9342);
and U9515 (N_9515,N_9315,N_9372);
nand U9516 (N_9516,N_9311,N_9347);
nand U9517 (N_9517,N_9212,N_9243);
and U9518 (N_9518,N_9231,N_9241);
and U9519 (N_9519,N_9214,N_9268);
or U9520 (N_9520,N_9230,N_9377);
or U9521 (N_9521,N_9301,N_9317);
nor U9522 (N_9522,N_9210,N_9341);
xor U9523 (N_9523,N_9300,N_9349);
xor U9524 (N_9524,N_9367,N_9377);
nand U9525 (N_9525,N_9334,N_9220);
nand U9526 (N_9526,N_9216,N_9340);
nand U9527 (N_9527,N_9296,N_9224);
nor U9528 (N_9528,N_9299,N_9218);
xor U9529 (N_9529,N_9255,N_9285);
and U9530 (N_9530,N_9377,N_9325);
nor U9531 (N_9531,N_9368,N_9287);
or U9532 (N_9532,N_9368,N_9340);
and U9533 (N_9533,N_9384,N_9204);
nor U9534 (N_9534,N_9336,N_9249);
and U9535 (N_9535,N_9324,N_9373);
nand U9536 (N_9536,N_9378,N_9210);
nand U9537 (N_9537,N_9285,N_9287);
xor U9538 (N_9538,N_9315,N_9222);
and U9539 (N_9539,N_9276,N_9333);
xnor U9540 (N_9540,N_9390,N_9208);
nor U9541 (N_9541,N_9385,N_9266);
xnor U9542 (N_9542,N_9397,N_9272);
nand U9543 (N_9543,N_9397,N_9238);
or U9544 (N_9544,N_9269,N_9307);
nor U9545 (N_9545,N_9274,N_9311);
xor U9546 (N_9546,N_9316,N_9269);
and U9547 (N_9547,N_9224,N_9370);
or U9548 (N_9548,N_9242,N_9302);
or U9549 (N_9549,N_9254,N_9328);
nor U9550 (N_9550,N_9285,N_9282);
or U9551 (N_9551,N_9357,N_9333);
nor U9552 (N_9552,N_9286,N_9221);
or U9553 (N_9553,N_9289,N_9335);
xor U9554 (N_9554,N_9352,N_9313);
xnor U9555 (N_9555,N_9276,N_9360);
xnor U9556 (N_9556,N_9370,N_9201);
or U9557 (N_9557,N_9304,N_9232);
xor U9558 (N_9558,N_9213,N_9354);
nor U9559 (N_9559,N_9232,N_9264);
or U9560 (N_9560,N_9375,N_9372);
or U9561 (N_9561,N_9271,N_9253);
nor U9562 (N_9562,N_9231,N_9395);
nand U9563 (N_9563,N_9331,N_9393);
nor U9564 (N_9564,N_9217,N_9225);
and U9565 (N_9565,N_9318,N_9275);
or U9566 (N_9566,N_9208,N_9265);
nor U9567 (N_9567,N_9220,N_9201);
nor U9568 (N_9568,N_9243,N_9373);
nor U9569 (N_9569,N_9366,N_9325);
xor U9570 (N_9570,N_9349,N_9257);
xor U9571 (N_9571,N_9331,N_9274);
and U9572 (N_9572,N_9271,N_9218);
or U9573 (N_9573,N_9242,N_9375);
nand U9574 (N_9574,N_9368,N_9362);
and U9575 (N_9575,N_9250,N_9285);
nand U9576 (N_9576,N_9261,N_9367);
nor U9577 (N_9577,N_9397,N_9333);
nor U9578 (N_9578,N_9273,N_9321);
and U9579 (N_9579,N_9246,N_9392);
nor U9580 (N_9580,N_9275,N_9315);
and U9581 (N_9581,N_9327,N_9262);
xor U9582 (N_9582,N_9227,N_9207);
nor U9583 (N_9583,N_9302,N_9314);
and U9584 (N_9584,N_9370,N_9390);
and U9585 (N_9585,N_9317,N_9234);
xnor U9586 (N_9586,N_9233,N_9395);
nand U9587 (N_9587,N_9223,N_9380);
nor U9588 (N_9588,N_9333,N_9384);
or U9589 (N_9589,N_9388,N_9317);
xnor U9590 (N_9590,N_9325,N_9293);
nor U9591 (N_9591,N_9303,N_9248);
nor U9592 (N_9592,N_9269,N_9223);
nand U9593 (N_9593,N_9307,N_9267);
nand U9594 (N_9594,N_9227,N_9328);
nand U9595 (N_9595,N_9218,N_9395);
nand U9596 (N_9596,N_9270,N_9272);
or U9597 (N_9597,N_9253,N_9241);
or U9598 (N_9598,N_9284,N_9372);
nand U9599 (N_9599,N_9337,N_9265);
and U9600 (N_9600,N_9528,N_9586);
or U9601 (N_9601,N_9588,N_9599);
nor U9602 (N_9602,N_9418,N_9442);
nor U9603 (N_9603,N_9511,N_9436);
xnor U9604 (N_9604,N_9474,N_9456);
nor U9605 (N_9605,N_9517,N_9550);
and U9606 (N_9606,N_9504,N_9541);
and U9607 (N_9607,N_9408,N_9489);
and U9608 (N_9608,N_9476,N_9443);
nand U9609 (N_9609,N_9593,N_9400);
or U9610 (N_9610,N_9404,N_9457);
or U9611 (N_9611,N_9486,N_9546);
and U9612 (N_9612,N_9585,N_9577);
and U9613 (N_9613,N_9407,N_9596);
nand U9614 (N_9614,N_9507,N_9576);
nand U9615 (N_9615,N_9477,N_9464);
xor U9616 (N_9616,N_9402,N_9462);
and U9617 (N_9617,N_9472,N_9427);
and U9618 (N_9618,N_9512,N_9547);
or U9619 (N_9619,N_9426,N_9557);
nand U9620 (N_9620,N_9467,N_9409);
xnor U9621 (N_9621,N_9564,N_9582);
and U9622 (N_9622,N_9548,N_9565);
and U9623 (N_9623,N_9411,N_9510);
xor U9624 (N_9624,N_9452,N_9578);
nand U9625 (N_9625,N_9433,N_9539);
or U9626 (N_9626,N_9424,N_9495);
and U9627 (N_9627,N_9532,N_9447);
or U9628 (N_9628,N_9590,N_9497);
nor U9629 (N_9629,N_9479,N_9566);
xor U9630 (N_9630,N_9439,N_9549);
nand U9631 (N_9631,N_9429,N_9534);
nor U9632 (N_9632,N_9563,N_9525);
nand U9633 (N_9633,N_9570,N_9449);
nand U9634 (N_9634,N_9491,N_9494);
or U9635 (N_9635,N_9551,N_9513);
and U9636 (N_9636,N_9468,N_9567);
and U9637 (N_9637,N_9560,N_9401);
nor U9638 (N_9638,N_9591,N_9453);
nor U9639 (N_9639,N_9448,N_9482);
xor U9640 (N_9640,N_9434,N_9473);
and U9641 (N_9641,N_9417,N_9422);
nor U9642 (N_9642,N_9581,N_9415);
and U9643 (N_9643,N_9441,N_9580);
nand U9644 (N_9644,N_9544,N_9420);
xnor U9645 (N_9645,N_9553,N_9431);
nor U9646 (N_9646,N_9554,N_9543);
nor U9647 (N_9647,N_9587,N_9555);
nor U9648 (N_9648,N_9579,N_9592);
nor U9649 (N_9649,N_9446,N_9505);
nor U9650 (N_9650,N_9561,N_9536);
or U9651 (N_9651,N_9527,N_9460);
nor U9652 (N_9652,N_9583,N_9562);
nor U9653 (N_9653,N_9481,N_9416);
or U9654 (N_9654,N_9465,N_9405);
xnor U9655 (N_9655,N_9530,N_9597);
and U9656 (N_9656,N_9503,N_9595);
and U9657 (N_9657,N_9538,N_9425);
xor U9658 (N_9658,N_9529,N_9435);
xor U9659 (N_9659,N_9501,N_9455);
nor U9660 (N_9660,N_9521,N_9545);
or U9661 (N_9661,N_9438,N_9499);
xor U9662 (N_9662,N_9522,N_9461);
or U9663 (N_9663,N_9569,N_9428);
nand U9664 (N_9664,N_9444,N_9535);
or U9665 (N_9665,N_9573,N_9502);
nand U9666 (N_9666,N_9594,N_9437);
nand U9667 (N_9667,N_9423,N_9493);
xor U9668 (N_9668,N_9552,N_9484);
nand U9669 (N_9669,N_9450,N_9478);
xor U9670 (N_9670,N_9440,N_9531);
or U9671 (N_9671,N_9537,N_9403);
xor U9672 (N_9672,N_9412,N_9589);
xor U9673 (N_9673,N_9483,N_9575);
nor U9674 (N_9674,N_9598,N_9518);
nor U9675 (N_9675,N_9413,N_9523);
or U9676 (N_9676,N_9533,N_9542);
nand U9677 (N_9677,N_9540,N_9524);
or U9678 (N_9678,N_9500,N_9520);
xnor U9679 (N_9679,N_9556,N_9506);
or U9680 (N_9680,N_9572,N_9519);
and U9681 (N_9681,N_9414,N_9559);
nand U9682 (N_9682,N_9516,N_9432);
nand U9683 (N_9683,N_9475,N_9454);
nor U9684 (N_9684,N_9471,N_9470);
and U9685 (N_9685,N_9469,N_9421);
xnor U9686 (N_9686,N_9466,N_9526);
and U9687 (N_9687,N_9458,N_9558);
or U9688 (N_9688,N_9514,N_9584);
and U9689 (N_9689,N_9509,N_9498);
and U9690 (N_9690,N_9410,N_9490);
nor U9691 (N_9691,N_9496,N_9568);
nand U9692 (N_9692,N_9485,N_9430);
nand U9693 (N_9693,N_9445,N_9487);
or U9694 (N_9694,N_9574,N_9406);
or U9695 (N_9695,N_9459,N_9451);
nor U9696 (N_9696,N_9571,N_9492);
and U9697 (N_9697,N_9480,N_9488);
and U9698 (N_9698,N_9419,N_9463);
nand U9699 (N_9699,N_9515,N_9508);
xor U9700 (N_9700,N_9561,N_9509);
and U9701 (N_9701,N_9516,N_9491);
and U9702 (N_9702,N_9485,N_9579);
and U9703 (N_9703,N_9452,N_9443);
nor U9704 (N_9704,N_9598,N_9523);
and U9705 (N_9705,N_9521,N_9520);
nor U9706 (N_9706,N_9443,N_9505);
or U9707 (N_9707,N_9544,N_9553);
xor U9708 (N_9708,N_9507,N_9492);
nand U9709 (N_9709,N_9463,N_9529);
xnor U9710 (N_9710,N_9408,N_9538);
xnor U9711 (N_9711,N_9489,N_9439);
or U9712 (N_9712,N_9505,N_9426);
or U9713 (N_9713,N_9463,N_9433);
nand U9714 (N_9714,N_9592,N_9479);
nand U9715 (N_9715,N_9567,N_9411);
xnor U9716 (N_9716,N_9592,N_9577);
nor U9717 (N_9717,N_9573,N_9505);
xor U9718 (N_9718,N_9555,N_9406);
nor U9719 (N_9719,N_9524,N_9484);
nor U9720 (N_9720,N_9561,N_9431);
nand U9721 (N_9721,N_9535,N_9495);
or U9722 (N_9722,N_9555,N_9530);
nor U9723 (N_9723,N_9536,N_9456);
and U9724 (N_9724,N_9546,N_9506);
or U9725 (N_9725,N_9581,N_9505);
and U9726 (N_9726,N_9597,N_9522);
and U9727 (N_9727,N_9492,N_9426);
and U9728 (N_9728,N_9425,N_9583);
nor U9729 (N_9729,N_9479,N_9422);
nor U9730 (N_9730,N_9567,N_9550);
or U9731 (N_9731,N_9457,N_9576);
and U9732 (N_9732,N_9443,N_9402);
or U9733 (N_9733,N_9520,N_9444);
or U9734 (N_9734,N_9559,N_9437);
or U9735 (N_9735,N_9545,N_9459);
or U9736 (N_9736,N_9535,N_9577);
nand U9737 (N_9737,N_9552,N_9492);
and U9738 (N_9738,N_9416,N_9419);
nand U9739 (N_9739,N_9453,N_9486);
nor U9740 (N_9740,N_9560,N_9476);
nor U9741 (N_9741,N_9516,N_9430);
xnor U9742 (N_9742,N_9512,N_9418);
and U9743 (N_9743,N_9414,N_9498);
xnor U9744 (N_9744,N_9530,N_9553);
and U9745 (N_9745,N_9516,N_9504);
xnor U9746 (N_9746,N_9408,N_9459);
and U9747 (N_9747,N_9459,N_9434);
and U9748 (N_9748,N_9501,N_9460);
and U9749 (N_9749,N_9428,N_9442);
and U9750 (N_9750,N_9493,N_9407);
nand U9751 (N_9751,N_9480,N_9523);
and U9752 (N_9752,N_9405,N_9482);
or U9753 (N_9753,N_9549,N_9479);
nor U9754 (N_9754,N_9511,N_9503);
or U9755 (N_9755,N_9500,N_9488);
or U9756 (N_9756,N_9471,N_9527);
nor U9757 (N_9757,N_9539,N_9595);
or U9758 (N_9758,N_9577,N_9579);
nor U9759 (N_9759,N_9562,N_9573);
or U9760 (N_9760,N_9482,N_9478);
xor U9761 (N_9761,N_9441,N_9475);
xnor U9762 (N_9762,N_9509,N_9517);
nor U9763 (N_9763,N_9444,N_9476);
xor U9764 (N_9764,N_9463,N_9570);
nor U9765 (N_9765,N_9520,N_9508);
nor U9766 (N_9766,N_9514,N_9458);
nor U9767 (N_9767,N_9558,N_9596);
or U9768 (N_9768,N_9475,N_9572);
nor U9769 (N_9769,N_9429,N_9427);
and U9770 (N_9770,N_9514,N_9575);
xor U9771 (N_9771,N_9541,N_9486);
nand U9772 (N_9772,N_9587,N_9575);
and U9773 (N_9773,N_9592,N_9480);
xor U9774 (N_9774,N_9471,N_9511);
xnor U9775 (N_9775,N_9545,N_9525);
or U9776 (N_9776,N_9405,N_9568);
nor U9777 (N_9777,N_9419,N_9464);
or U9778 (N_9778,N_9538,N_9523);
xor U9779 (N_9779,N_9551,N_9477);
nor U9780 (N_9780,N_9448,N_9449);
xnor U9781 (N_9781,N_9508,N_9533);
xnor U9782 (N_9782,N_9565,N_9516);
or U9783 (N_9783,N_9434,N_9527);
or U9784 (N_9784,N_9443,N_9574);
xor U9785 (N_9785,N_9535,N_9501);
nand U9786 (N_9786,N_9582,N_9562);
and U9787 (N_9787,N_9464,N_9550);
and U9788 (N_9788,N_9444,N_9403);
nor U9789 (N_9789,N_9460,N_9538);
xnor U9790 (N_9790,N_9532,N_9511);
xnor U9791 (N_9791,N_9591,N_9501);
nor U9792 (N_9792,N_9577,N_9536);
and U9793 (N_9793,N_9504,N_9540);
nor U9794 (N_9794,N_9529,N_9599);
nand U9795 (N_9795,N_9459,N_9449);
nand U9796 (N_9796,N_9459,N_9490);
nor U9797 (N_9797,N_9570,N_9514);
or U9798 (N_9798,N_9423,N_9596);
and U9799 (N_9799,N_9542,N_9505);
and U9800 (N_9800,N_9625,N_9622);
xnor U9801 (N_9801,N_9673,N_9715);
xnor U9802 (N_9802,N_9763,N_9638);
xor U9803 (N_9803,N_9693,N_9672);
nand U9804 (N_9804,N_9692,N_9703);
nand U9805 (N_9805,N_9781,N_9761);
or U9806 (N_9806,N_9769,N_9795);
nand U9807 (N_9807,N_9608,N_9647);
xnor U9808 (N_9808,N_9753,N_9752);
and U9809 (N_9809,N_9780,N_9728);
and U9810 (N_9810,N_9727,N_9605);
or U9811 (N_9811,N_9745,N_9774);
nor U9812 (N_9812,N_9686,N_9737);
nand U9813 (N_9813,N_9704,N_9792);
and U9814 (N_9814,N_9600,N_9661);
and U9815 (N_9815,N_9614,N_9716);
nor U9816 (N_9816,N_9665,N_9734);
or U9817 (N_9817,N_9666,N_9682);
and U9818 (N_9818,N_9687,N_9617);
and U9819 (N_9819,N_9644,N_9615);
and U9820 (N_9820,N_9705,N_9604);
nand U9821 (N_9821,N_9607,N_9711);
nand U9822 (N_9822,N_9697,N_9675);
and U9823 (N_9823,N_9739,N_9751);
or U9824 (N_9824,N_9606,N_9710);
xor U9825 (N_9825,N_9725,N_9790);
nand U9826 (N_9826,N_9629,N_9655);
and U9827 (N_9827,N_9740,N_9779);
xnor U9828 (N_9828,N_9624,N_9755);
nor U9829 (N_9829,N_9764,N_9729);
nand U9830 (N_9830,N_9713,N_9791);
or U9831 (N_9831,N_9632,N_9640);
nor U9832 (N_9832,N_9771,N_9766);
or U9833 (N_9833,N_9707,N_9639);
xor U9834 (N_9834,N_9700,N_9690);
or U9835 (N_9835,N_9793,N_9656);
or U9836 (N_9836,N_9699,N_9775);
xnor U9837 (N_9837,N_9748,N_9799);
or U9838 (N_9838,N_9654,N_9749);
and U9839 (N_9839,N_9694,N_9797);
or U9840 (N_9840,N_9721,N_9626);
nand U9841 (N_9841,N_9601,N_9696);
nor U9842 (N_9842,N_9668,N_9735);
or U9843 (N_9843,N_9663,N_9657);
xnor U9844 (N_9844,N_9714,N_9630);
and U9845 (N_9845,N_9648,N_9635);
xor U9846 (N_9846,N_9743,N_9603);
nor U9847 (N_9847,N_9720,N_9768);
or U9848 (N_9848,N_9623,N_9789);
nand U9849 (N_9849,N_9760,N_9733);
nand U9850 (N_9850,N_9645,N_9689);
nor U9851 (N_9851,N_9679,N_9784);
xnor U9852 (N_9852,N_9754,N_9650);
xor U9853 (N_9853,N_9620,N_9765);
nor U9854 (N_9854,N_9747,N_9712);
nor U9855 (N_9855,N_9643,N_9702);
and U9856 (N_9856,N_9723,N_9613);
or U9857 (N_9857,N_9724,N_9683);
and U9858 (N_9858,N_9610,N_9612);
nor U9859 (N_9859,N_9742,N_9641);
nand U9860 (N_9860,N_9738,N_9688);
or U9861 (N_9861,N_9762,N_9651);
or U9862 (N_9862,N_9787,N_9636);
and U9863 (N_9863,N_9649,N_9756);
nor U9864 (N_9864,N_9627,N_9678);
xnor U9865 (N_9865,N_9684,N_9767);
xnor U9866 (N_9866,N_9619,N_9646);
nand U9867 (N_9867,N_9770,N_9776);
xor U9868 (N_9868,N_9691,N_9709);
nand U9869 (N_9869,N_9746,N_9653);
nand U9870 (N_9870,N_9732,N_9621);
or U9871 (N_9871,N_9731,N_9680);
nand U9872 (N_9872,N_9685,N_9759);
or U9873 (N_9873,N_9677,N_9676);
or U9874 (N_9874,N_9772,N_9744);
and U9875 (N_9875,N_9718,N_9695);
xnor U9876 (N_9876,N_9777,N_9796);
nand U9877 (N_9877,N_9664,N_9782);
xor U9878 (N_9878,N_9637,N_9750);
nand U9879 (N_9879,N_9788,N_9634);
nand U9880 (N_9880,N_9662,N_9659);
xor U9881 (N_9881,N_9741,N_9794);
nor U9882 (N_9882,N_9786,N_9757);
and U9883 (N_9883,N_9631,N_9652);
nand U9884 (N_9884,N_9660,N_9628);
nor U9885 (N_9885,N_9609,N_9726);
and U9886 (N_9886,N_9706,N_9669);
or U9887 (N_9887,N_9708,N_9717);
nand U9888 (N_9888,N_9719,N_9658);
xor U9889 (N_9889,N_9698,N_9611);
or U9890 (N_9890,N_9633,N_9778);
or U9891 (N_9891,N_9773,N_9758);
nor U9892 (N_9892,N_9785,N_9642);
and U9893 (N_9893,N_9736,N_9670);
nor U9894 (N_9894,N_9602,N_9798);
and U9895 (N_9895,N_9671,N_9722);
or U9896 (N_9896,N_9616,N_9667);
nand U9897 (N_9897,N_9783,N_9681);
and U9898 (N_9898,N_9730,N_9701);
nor U9899 (N_9899,N_9618,N_9674);
nor U9900 (N_9900,N_9754,N_9679);
or U9901 (N_9901,N_9627,N_9695);
nand U9902 (N_9902,N_9767,N_9753);
and U9903 (N_9903,N_9695,N_9614);
and U9904 (N_9904,N_9639,N_9629);
nand U9905 (N_9905,N_9795,N_9786);
and U9906 (N_9906,N_9613,N_9673);
xor U9907 (N_9907,N_9696,N_9651);
xnor U9908 (N_9908,N_9722,N_9677);
and U9909 (N_9909,N_9684,N_9621);
and U9910 (N_9910,N_9637,N_9630);
or U9911 (N_9911,N_9743,N_9704);
xor U9912 (N_9912,N_9658,N_9768);
nor U9913 (N_9913,N_9600,N_9786);
nand U9914 (N_9914,N_9786,N_9652);
xnor U9915 (N_9915,N_9745,N_9770);
nand U9916 (N_9916,N_9713,N_9775);
and U9917 (N_9917,N_9700,N_9640);
nor U9918 (N_9918,N_9738,N_9746);
nand U9919 (N_9919,N_9657,N_9629);
or U9920 (N_9920,N_9649,N_9670);
nor U9921 (N_9921,N_9750,N_9790);
or U9922 (N_9922,N_9644,N_9708);
and U9923 (N_9923,N_9692,N_9701);
nand U9924 (N_9924,N_9674,N_9778);
or U9925 (N_9925,N_9790,N_9683);
and U9926 (N_9926,N_9737,N_9666);
xnor U9927 (N_9927,N_9677,N_9674);
and U9928 (N_9928,N_9637,N_9615);
nand U9929 (N_9929,N_9690,N_9600);
nor U9930 (N_9930,N_9746,N_9727);
nor U9931 (N_9931,N_9634,N_9731);
nand U9932 (N_9932,N_9607,N_9731);
nor U9933 (N_9933,N_9789,N_9645);
nand U9934 (N_9934,N_9785,N_9685);
or U9935 (N_9935,N_9639,N_9664);
and U9936 (N_9936,N_9705,N_9672);
or U9937 (N_9937,N_9716,N_9695);
nand U9938 (N_9938,N_9620,N_9708);
and U9939 (N_9939,N_9644,N_9772);
and U9940 (N_9940,N_9707,N_9778);
and U9941 (N_9941,N_9643,N_9637);
or U9942 (N_9942,N_9695,N_9740);
or U9943 (N_9943,N_9796,N_9651);
or U9944 (N_9944,N_9675,N_9717);
nand U9945 (N_9945,N_9723,N_9758);
and U9946 (N_9946,N_9784,N_9745);
and U9947 (N_9947,N_9796,N_9639);
xnor U9948 (N_9948,N_9617,N_9644);
nor U9949 (N_9949,N_9764,N_9672);
xnor U9950 (N_9950,N_9740,N_9792);
xnor U9951 (N_9951,N_9741,N_9624);
nand U9952 (N_9952,N_9634,N_9717);
and U9953 (N_9953,N_9680,N_9766);
xor U9954 (N_9954,N_9602,N_9741);
nand U9955 (N_9955,N_9727,N_9711);
nand U9956 (N_9956,N_9789,N_9671);
or U9957 (N_9957,N_9776,N_9655);
xor U9958 (N_9958,N_9737,N_9753);
and U9959 (N_9959,N_9602,N_9770);
xor U9960 (N_9960,N_9733,N_9687);
or U9961 (N_9961,N_9623,N_9643);
and U9962 (N_9962,N_9603,N_9762);
nor U9963 (N_9963,N_9647,N_9752);
nor U9964 (N_9964,N_9762,N_9700);
xnor U9965 (N_9965,N_9711,N_9715);
and U9966 (N_9966,N_9664,N_9612);
nand U9967 (N_9967,N_9679,N_9615);
or U9968 (N_9968,N_9757,N_9641);
xor U9969 (N_9969,N_9662,N_9703);
nand U9970 (N_9970,N_9759,N_9614);
or U9971 (N_9971,N_9766,N_9716);
nor U9972 (N_9972,N_9664,N_9700);
or U9973 (N_9973,N_9630,N_9651);
nand U9974 (N_9974,N_9778,N_9695);
nor U9975 (N_9975,N_9642,N_9641);
xnor U9976 (N_9976,N_9723,N_9614);
and U9977 (N_9977,N_9775,N_9694);
nand U9978 (N_9978,N_9680,N_9743);
nor U9979 (N_9979,N_9745,N_9692);
xnor U9980 (N_9980,N_9619,N_9726);
nor U9981 (N_9981,N_9744,N_9606);
and U9982 (N_9982,N_9755,N_9767);
nand U9983 (N_9983,N_9700,N_9604);
and U9984 (N_9984,N_9657,N_9683);
or U9985 (N_9985,N_9721,N_9729);
nand U9986 (N_9986,N_9786,N_9758);
nor U9987 (N_9987,N_9649,N_9615);
nor U9988 (N_9988,N_9752,N_9784);
xor U9989 (N_9989,N_9610,N_9767);
xor U9990 (N_9990,N_9729,N_9771);
nand U9991 (N_9991,N_9646,N_9624);
nand U9992 (N_9992,N_9722,N_9695);
and U9993 (N_9993,N_9794,N_9610);
nand U9994 (N_9994,N_9709,N_9701);
nor U9995 (N_9995,N_9724,N_9619);
nand U9996 (N_9996,N_9789,N_9767);
nor U9997 (N_9997,N_9761,N_9759);
or U9998 (N_9998,N_9618,N_9694);
or U9999 (N_9999,N_9793,N_9664);
xnor U10000 (N_10000,N_9990,N_9994);
or U10001 (N_10001,N_9867,N_9888);
nor U10002 (N_10002,N_9881,N_9808);
xnor U10003 (N_10003,N_9998,N_9807);
and U10004 (N_10004,N_9918,N_9912);
or U10005 (N_10005,N_9909,N_9925);
nand U10006 (N_10006,N_9898,N_9855);
nand U10007 (N_10007,N_9906,N_9955);
and U10008 (N_10008,N_9956,N_9938);
nor U10009 (N_10009,N_9966,N_9852);
xnor U10010 (N_10010,N_9907,N_9826);
nor U10011 (N_10011,N_9838,N_9854);
xnor U10012 (N_10012,N_9819,N_9839);
or U10013 (N_10013,N_9823,N_9857);
and U10014 (N_10014,N_9983,N_9922);
xor U10015 (N_10015,N_9978,N_9962);
nand U10016 (N_10016,N_9836,N_9833);
nand U10017 (N_10017,N_9902,N_9970);
nor U10018 (N_10018,N_9940,N_9976);
xor U10019 (N_10019,N_9841,N_9917);
nand U10020 (N_10020,N_9911,N_9923);
xnor U10021 (N_10021,N_9893,N_9952);
nor U10022 (N_10022,N_9934,N_9860);
xor U10023 (N_10023,N_9827,N_9942);
nor U10024 (N_10024,N_9984,N_9948);
and U10025 (N_10025,N_9943,N_9930);
nor U10026 (N_10026,N_9992,N_9968);
or U10027 (N_10027,N_9979,N_9862);
nand U10028 (N_10028,N_9928,N_9964);
or U10029 (N_10029,N_9802,N_9886);
or U10030 (N_10030,N_9818,N_9878);
nor U10031 (N_10031,N_9961,N_9870);
nand U10032 (N_10032,N_9832,N_9879);
and U10033 (N_10033,N_9863,N_9971);
and U10034 (N_10034,N_9959,N_9829);
xnor U10035 (N_10035,N_9908,N_9900);
nor U10036 (N_10036,N_9828,N_9884);
nor U10037 (N_10037,N_9965,N_9865);
nor U10038 (N_10038,N_9859,N_9946);
or U10039 (N_10039,N_9873,N_9901);
and U10040 (N_10040,N_9931,N_9840);
nor U10041 (N_10041,N_9920,N_9847);
and U10042 (N_10042,N_9866,N_9844);
or U10043 (N_10043,N_9945,N_9896);
or U10044 (N_10044,N_9825,N_9805);
nor U10045 (N_10045,N_9846,N_9835);
and U10046 (N_10046,N_9939,N_9915);
nor U10047 (N_10047,N_9861,N_9989);
xor U10048 (N_10048,N_9877,N_9820);
and U10049 (N_10049,N_9985,N_9975);
or U10050 (N_10050,N_9895,N_9916);
nor U10051 (N_10051,N_9951,N_9837);
xnor U10052 (N_10052,N_9967,N_9804);
and U10053 (N_10053,N_9980,N_9949);
nand U10054 (N_10054,N_9894,N_9813);
nand U10055 (N_10055,N_9914,N_9972);
xor U10056 (N_10056,N_9904,N_9811);
or U10057 (N_10057,N_9995,N_9815);
nor U10058 (N_10058,N_9817,N_9876);
nand U10059 (N_10059,N_9927,N_9868);
nand U10060 (N_10060,N_9869,N_9999);
xnor U10061 (N_10061,N_9803,N_9889);
or U10062 (N_10062,N_9988,N_9801);
or U10063 (N_10063,N_9899,N_9848);
and U10064 (N_10064,N_9882,N_9973);
nand U10065 (N_10065,N_9822,N_9937);
and U10066 (N_10066,N_9842,N_9806);
or U10067 (N_10067,N_9903,N_9834);
or U10068 (N_10068,N_9821,N_9814);
nand U10069 (N_10069,N_9850,N_9987);
or U10070 (N_10070,N_9875,N_9885);
and U10071 (N_10071,N_9947,N_9977);
and U10072 (N_10072,N_9810,N_9974);
and U10073 (N_10073,N_9933,N_9864);
xnor U10074 (N_10074,N_9872,N_9996);
nand U10075 (N_10075,N_9953,N_9809);
xnor U10076 (N_10076,N_9892,N_9874);
nor U10077 (N_10077,N_9880,N_9891);
nand U10078 (N_10078,N_9849,N_9929);
and U10079 (N_10079,N_9831,N_9845);
nor U10080 (N_10080,N_9944,N_9887);
xnor U10081 (N_10081,N_9986,N_9991);
nor U10082 (N_10082,N_9812,N_9883);
or U10083 (N_10083,N_9816,N_9910);
nand U10084 (N_10084,N_9969,N_9800);
nand U10085 (N_10085,N_9957,N_9851);
or U10086 (N_10086,N_9993,N_9932);
nor U10087 (N_10087,N_9871,N_9924);
or U10088 (N_10088,N_9926,N_9935);
and U10089 (N_10089,N_9950,N_9897);
nand U10090 (N_10090,N_9824,N_9905);
and U10091 (N_10091,N_9919,N_9997);
xnor U10092 (N_10092,N_9960,N_9936);
nor U10093 (N_10093,N_9856,N_9941);
nor U10094 (N_10094,N_9981,N_9858);
nor U10095 (N_10095,N_9963,N_9843);
and U10096 (N_10096,N_9958,N_9913);
nor U10097 (N_10097,N_9954,N_9982);
nor U10098 (N_10098,N_9853,N_9921);
and U10099 (N_10099,N_9890,N_9830);
nand U10100 (N_10100,N_9966,N_9894);
xor U10101 (N_10101,N_9910,N_9883);
nor U10102 (N_10102,N_9994,N_9827);
xnor U10103 (N_10103,N_9828,N_9982);
xnor U10104 (N_10104,N_9936,N_9860);
nand U10105 (N_10105,N_9946,N_9987);
nor U10106 (N_10106,N_9913,N_9814);
xnor U10107 (N_10107,N_9823,N_9902);
or U10108 (N_10108,N_9920,N_9953);
nor U10109 (N_10109,N_9853,N_9951);
xor U10110 (N_10110,N_9865,N_9800);
xor U10111 (N_10111,N_9998,N_9970);
and U10112 (N_10112,N_9830,N_9914);
or U10113 (N_10113,N_9998,N_9826);
and U10114 (N_10114,N_9801,N_9891);
or U10115 (N_10115,N_9894,N_9957);
and U10116 (N_10116,N_9979,N_9945);
or U10117 (N_10117,N_9880,N_9930);
xor U10118 (N_10118,N_9951,N_9901);
and U10119 (N_10119,N_9859,N_9936);
or U10120 (N_10120,N_9979,N_9853);
nand U10121 (N_10121,N_9931,N_9902);
xnor U10122 (N_10122,N_9956,N_9957);
or U10123 (N_10123,N_9930,N_9800);
or U10124 (N_10124,N_9885,N_9838);
or U10125 (N_10125,N_9920,N_9841);
nand U10126 (N_10126,N_9835,N_9824);
or U10127 (N_10127,N_9861,N_9937);
xor U10128 (N_10128,N_9803,N_9905);
nor U10129 (N_10129,N_9812,N_9857);
or U10130 (N_10130,N_9841,N_9829);
and U10131 (N_10131,N_9807,N_9852);
nor U10132 (N_10132,N_9840,N_9979);
nand U10133 (N_10133,N_9916,N_9913);
nand U10134 (N_10134,N_9829,N_9878);
xnor U10135 (N_10135,N_9952,N_9874);
xnor U10136 (N_10136,N_9966,N_9953);
nand U10137 (N_10137,N_9931,N_9824);
or U10138 (N_10138,N_9952,N_9929);
and U10139 (N_10139,N_9881,N_9927);
nand U10140 (N_10140,N_9950,N_9884);
xnor U10141 (N_10141,N_9932,N_9814);
xor U10142 (N_10142,N_9948,N_9893);
nand U10143 (N_10143,N_9913,N_9829);
and U10144 (N_10144,N_9948,N_9867);
nand U10145 (N_10145,N_9905,N_9935);
xor U10146 (N_10146,N_9917,N_9973);
and U10147 (N_10147,N_9994,N_9876);
nor U10148 (N_10148,N_9803,N_9834);
and U10149 (N_10149,N_9901,N_9933);
and U10150 (N_10150,N_9879,N_9944);
or U10151 (N_10151,N_9946,N_9842);
nand U10152 (N_10152,N_9942,N_9998);
nand U10153 (N_10153,N_9988,N_9897);
or U10154 (N_10154,N_9853,N_9843);
nand U10155 (N_10155,N_9800,N_9923);
xnor U10156 (N_10156,N_9831,N_9827);
xnor U10157 (N_10157,N_9844,N_9939);
nor U10158 (N_10158,N_9882,N_9917);
xor U10159 (N_10159,N_9844,N_9986);
or U10160 (N_10160,N_9953,N_9839);
and U10161 (N_10161,N_9886,N_9953);
xor U10162 (N_10162,N_9916,N_9872);
xor U10163 (N_10163,N_9904,N_9800);
xnor U10164 (N_10164,N_9993,N_9826);
nor U10165 (N_10165,N_9990,N_9872);
nand U10166 (N_10166,N_9950,N_9832);
or U10167 (N_10167,N_9949,N_9806);
and U10168 (N_10168,N_9830,N_9846);
nor U10169 (N_10169,N_9917,N_9946);
nand U10170 (N_10170,N_9971,N_9968);
nand U10171 (N_10171,N_9968,N_9833);
nand U10172 (N_10172,N_9810,N_9891);
nand U10173 (N_10173,N_9894,N_9819);
nor U10174 (N_10174,N_9968,N_9919);
and U10175 (N_10175,N_9884,N_9859);
nor U10176 (N_10176,N_9919,N_9825);
nand U10177 (N_10177,N_9856,N_9936);
and U10178 (N_10178,N_9841,N_9986);
nor U10179 (N_10179,N_9854,N_9911);
and U10180 (N_10180,N_9959,N_9897);
or U10181 (N_10181,N_9984,N_9817);
and U10182 (N_10182,N_9813,N_9918);
nand U10183 (N_10183,N_9916,N_9848);
nand U10184 (N_10184,N_9958,N_9849);
xor U10185 (N_10185,N_9829,N_9988);
nand U10186 (N_10186,N_9836,N_9802);
nor U10187 (N_10187,N_9830,N_9868);
and U10188 (N_10188,N_9890,N_9853);
and U10189 (N_10189,N_9943,N_9848);
and U10190 (N_10190,N_9895,N_9950);
and U10191 (N_10191,N_9860,N_9951);
nand U10192 (N_10192,N_9809,N_9948);
nand U10193 (N_10193,N_9802,N_9923);
xor U10194 (N_10194,N_9917,N_9979);
and U10195 (N_10195,N_9837,N_9947);
or U10196 (N_10196,N_9993,N_9938);
and U10197 (N_10197,N_9808,N_9980);
xor U10198 (N_10198,N_9805,N_9814);
nand U10199 (N_10199,N_9949,N_9925);
nor U10200 (N_10200,N_10131,N_10021);
nand U10201 (N_10201,N_10026,N_10061);
xnor U10202 (N_10202,N_10135,N_10060);
and U10203 (N_10203,N_10162,N_10035);
and U10204 (N_10204,N_10157,N_10041);
or U10205 (N_10205,N_10175,N_10125);
xnor U10206 (N_10206,N_10111,N_10073);
nor U10207 (N_10207,N_10070,N_10112);
or U10208 (N_10208,N_10142,N_10078);
nor U10209 (N_10209,N_10055,N_10039);
xnor U10210 (N_10210,N_10056,N_10120);
or U10211 (N_10211,N_10161,N_10119);
nand U10212 (N_10212,N_10168,N_10109);
nand U10213 (N_10213,N_10054,N_10134);
or U10214 (N_10214,N_10029,N_10046);
xor U10215 (N_10215,N_10100,N_10025);
nor U10216 (N_10216,N_10133,N_10190);
xor U10217 (N_10217,N_10185,N_10079);
nor U10218 (N_10218,N_10163,N_10166);
and U10219 (N_10219,N_10178,N_10167);
xnor U10220 (N_10220,N_10186,N_10188);
or U10221 (N_10221,N_10030,N_10053);
nor U10222 (N_10222,N_10118,N_10152);
nor U10223 (N_10223,N_10144,N_10095);
and U10224 (N_10224,N_10007,N_10031);
or U10225 (N_10225,N_10011,N_10067);
nor U10226 (N_10226,N_10148,N_10003);
or U10227 (N_10227,N_10088,N_10004);
and U10228 (N_10228,N_10065,N_10108);
nand U10229 (N_10229,N_10027,N_10128);
and U10230 (N_10230,N_10172,N_10158);
or U10231 (N_10231,N_10138,N_10034);
nor U10232 (N_10232,N_10075,N_10000);
nand U10233 (N_10233,N_10062,N_10001);
nor U10234 (N_10234,N_10040,N_10082);
or U10235 (N_10235,N_10077,N_10022);
xor U10236 (N_10236,N_10193,N_10028);
or U10237 (N_10237,N_10182,N_10098);
and U10238 (N_10238,N_10023,N_10057);
xnor U10239 (N_10239,N_10006,N_10038);
nor U10240 (N_10240,N_10071,N_10103);
xor U10241 (N_10241,N_10149,N_10124);
nand U10242 (N_10242,N_10094,N_10192);
and U10243 (N_10243,N_10130,N_10066);
nor U10244 (N_10244,N_10009,N_10008);
nor U10245 (N_10245,N_10197,N_10147);
and U10246 (N_10246,N_10123,N_10129);
and U10247 (N_10247,N_10116,N_10164);
xnor U10248 (N_10248,N_10020,N_10086);
nor U10249 (N_10249,N_10052,N_10084);
nand U10250 (N_10250,N_10195,N_10102);
and U10251 (N_10251,N_10110,N_10083);
xnor U10252 (N_10252,N_10187,N_10101);
xor U10253 (N_10253,N_10154,N_10136);
xnor U10254 (N_10254,N_10173,N_10177);
and U10255 (N_10255,N_10032,N_10151);
nand U10256 (N_10256,N_10005,N_10159);
or U10257 (N_10257,N_10170,N_10146);
nor U10258 (N_10258,N_10018,N_10132);
xor U10259 (N_10259,N_10122,N_10097);
nand U10260 (N_10260,N_10194,N_10051);
nand U10261 (N_10261,N_10155,N_10012);
or U10262 (N_10262,N_10064,N_10181);
and U10263 (N_10263,N_10196,N_10019);
nand U10264 (N_10264,N_10050,N_10127);
or U10265 (N_10265,N_10092,N_10099);
xnor U10266 (N_10266,N_10198,N_10069);
nor U10267 (N_10267,N_10015,N_10013);
xor U10268 (N_10268,N_10081,N_10121);
nand U10269 (N_10269,N_10063,N_10058);
and U10270 (N_10270,N_10180,N_10091);
nor U10271 (N_10271,N_10150,N_10089);
nand U10272 (N_10272,N_10080,N_10036);
or U10273 (N_10273,N_10010,N_10113);
xor U10274 (N_10274,N_10165,N_10105);
nor U10275 (N_10275,N_10059,N_10114);
or U10276 (N_10276,N_10044,N_10183);
or U10277 (N_10277,N_10139,N_10047);
nor U10278 (N_10278,N_10087,N_10153);
nor U10279 (N_10279,N_10107,N_10143);
nor U10280 (N_10280,N_10085,N_10106);
and U10281 (N_10281,N_10072,N_10191);
xnor U10282 (N_10282,N_10045,N_10117);
nand U10283 (N_10283,N_10189,N_10016);
xor U10284 (N_10284,N_10068,N_10043);
nand U10285 (N_10285,N_10093,N_10174);
nand U10286 (N_10286,N_10141,N_10137);
nor U10287 (N_10287,N_10199,N_10037);
xor U10288 (N_10288,N_10048,N_10156);
nor U10289 (N_10289,N_10033,N_10104);
xnor U10290 (N_10290,N_10014,N_10145);
nor U10291 (N_10291,N_10074,N_10042);
nor U10292 (N_10292,N_10140,N_10076);
and U10293 (N_10293,N_10017,N_10184);
xnor U10294 (N_10294,N_10179,N_10160);
nor U10295 (N_10295,N_10171,N_10176);
or U10296 (N_10296,N_10049,N_10024);
or U10297 (N_10297,N_10126,N_10115);
nor U10298 (N_10298,N_10169,N_10002);
and U10299 (N_10299,N_10090,N_10096);
xor U10300 (N_10300,N_10009,N_10180);
or U10301 (N_10301,N_10091,N_10041);
and U10302 (N_10302,N_10112,N_10017);
and U10303 (N_10303,N_10047,N_10065);
nor U10304 (N_10304,N_10089,N_10166);
xor U10305 (N_10305,N_10111,N_10114);
and U10306 (N_10306,N_10016,N_10004);
or U10307 (N_10307,N_10052,N_10066);
nor U10308 (N_10308,N_10172,N_10031);
nor U10309 (N_10309,N_10005,N_10050);
nand U10310 (N_10310,N_10037,N_10171);
nor U10311 (N_10311,N_10194,N_10184);
xnor U10312 (N_10312,N_10154,N_10113);
nor U10313 (N_10313,N_10045,N_10074);
nor U10314 (N_10314,N_10084,N_10174);
and U10315 (N_10315,N_10167,N_10019);
nand U10316 (N_10316,N_10180,N_10001);
or U10317 (N_10317,N_10114,N_10096);
or U10318 (N_10318,N_10017,N_10105);
nand U10319 (N_10319,N_10165,N_10194);
nor U10320 (N_10320,N_10076,N_10123);
nor U10321 (N_10321,N_10147,N_10115);
xnor U10322 (N_10322,N_10135,N_10116);
nor U10323 (N_10323,N_10014,N_10026);
xnor U10324 (N_10324,N_10191,N_10024);
nand U10325 (N_10325,N_10174,N_10117);
nand U10326 (N_10326,N_10175,N_10157);
xor U10327 (N_10327,N_10146,N_10143);
nor U10328 (N_10328,N_10074,N_10116);
nor U10329 (N_10329,N_10182,N_10185);
nor U10330 (N_10330,N_10101,N_10094);
nor U10331 (N_10331,N_10059,N_10168);
and U10332 (N_10332,N_10190,N_10019);
nor U10333 (N_10333,N_10177,N_10011);
nor U10334 (N_10334,N_10094,N_10070);
xnor U10335 (N_10335,N_10116,N_10015);
nand U10336 (N_10336,N_10029,N_10170);
nor U10337 (N_10337,N_10125,N_10168);
nor U10338 (N_10338,N_10125,N_10035);
or U10339 (N_10339,N_10136,N_10158);
and U10340 (N_10340,N_10158,N_10046);
and U10341 (N_10341,N_10156,N_10027);
xnor U10342 (N_10342,N_10005,N_10026);
nor U10343 (N_10343,N_10095,N_10078);
nand U10344 (N_10344,N_10196,N_10108);
or U10345 (N_10345,N_10072,N_10178);
xor U10346 (N_10346,N_10130,N_10188);
or U10347 (N_10347,N_10090,N_10137);
or U10348 (N_10348,N_10096,N_10109);
xnor U10349 (N_10349,N_10014,N_10083);
nand U10350 (N_10350,N_10065,N_10146);
and U10351 (N_10351,N_10126,N_10049);
xnor U10352 (N_10352,N_10140,N_10024);
or U10353 (N_10353,N_10060,N_10187);
nand U10354 (N_10354,N_10194,N_10010);
nand U10355 (N_10355,N_10198,N_10121);
or U10356 (N_10356,N_10059,N_10039);
xnor U10357 (N_10357,N_10046,N_10045);
or U10358 (N_10358,N_10005,N_10013);
xor U10359 (N_10359,N_10053,N_10023);
xor U10360 (N_10360,N_10039,N_10057);
nand U10361 (N_10361,N_10070,N_10106);
and U10362 (N_10362,N_10064,N_10156);
or U10363 (N_10363,N_10038,N_10133);
or U10364 (N_10364,N_10014,N_10065);
nor U10365 (N_10365,N_10056,N_10114);
and U10366 (N_10366,N_10197,N_10090);
nand U10367 (N_10367,N_10159,N_10070);
nand U10368 (N_10368,N_10114,N_10192);
xnor U10369 (N_10369,N_10105,N_10168);
nor U10370 (N_10370,N_10182,N_10179);
nand U10371 (N_10371,N_10004,N_10062);
and U10372 (N_10372,N_10177,N_10167);
nand U10373 (N_10373,N_10156,N_10147);
and U10374 (N_10374,N_10040,N_10119);
xnor U10375 (N_10375,N_10124,N_10198);
nor U10376 (N_10376,N_10120,N_10023);
or U10377 (N_10377,N_10174,N_10006);
xor U10378 (N_10378,N_10038,N_10114);
nor U10379 (N_10379,N_10044,N_10037);
nor U10380 (N_10380,N_10196,N_10185);
xnor U10381 (N_10381,N_10069,N_10046);
and U10382 (N_10382,N_10077,N_10199);
nor U10383 (N_10383,N_10135,N_10113);
or U10384 (N_10384,N_10050,N_10008);
nand U10385 (N_10385,N_10160,N_10116);
nand U10386 (N_10386,N_10104,N_10187);
nand U10387 (N_10387,N_10150,N_10168);
nor U10388 (N_10388,N_10093,N_10151);
nand U10389 (N_10389,N_10007,N_10078);
nor U10390 (N_10390,N_10047,N_10110);
nand U10391 (N_10391,N_10119,N_10096);
or U10392 (N_10392,N_10038,N_10040);
xor U10393 (N_10393,N_10185,N_10103);
or U10394 (N_10394,N_10129,N_10101);
nand U10395 (N_10395,N_10099,N_10163);
nand U10396 (N_10396,N_10184,N_10118);
and U10397 (N_10397,N_10130,N_10024);
and U10398 (N_10398,N_10098,N_10089);
nand U10399 (N_10399,N_10112,N_10065);
nand U10400 (N_10400,N_10239,N_10385);
nand U10401 (N_10401,N_10247,N_10215);
and U10402 (N_10402,N_10356,N_10233);
xnor U10403 (N_10403,N_10321,N_10200);
nand U10404 (N_10404,N_10294,N_10302);
or U10405 (N_10405,N_10228,N_10201);
xnor U10406 (N_10406,N_10389,N_10382);
nor U10407 (N_10407,N_10358,N_10284);
and U10408 (N_10408,N_10292,N_10384);
and U10409 (N_10409,N_10353,N_10315);
xor U10410 (N_10410,N_10261,N_10216);
xnor U10411 (N_10411,N_10330,N_10311);
xnor U10412 (N_10412,N_10269,N_10245);
nor U10413 (N_10413,N_10285,N_10367);
nor U10414 (N_10414,N_10300,N_10303);
nand U10415 (N_10415,N_10364,N_10256);
xnor U10416 (N_10416,N_10307,N_10267);
or U10417 (N_10417,N_10249,N_10281);
and U10418 (N_10418,N_10386,N_10318);
xnor U10419 (N_10419,N_10243,N_10263);
and U10420 (N_10420,N_10211,N_10387);
nand U10421 (N_10421,N_10255,N_10209);
xnor U10422 (N_10422,N_10277,N_10316);
or U10423 (N_10423,N_10238,N_10324);
xnor U10424 (N_10424,N_10378,N_10348);
nand U10425 (N_10425,N_10399,N_10379);
nor U10426 (N_10426,N_10349,N_10250);
xnor U10427 (N_10427,N_10363,N_10271);
nor U10428 (N_10428,N_10212,N_10265);
or U10429 (N_10429,N_10217,N_10373);
and U10430 (N_10430,N_10388,N_10397);
nand U10431 (N_10431,N_10394,N_10288);
xor U10432 (N_10432,N_10213,N_10275);
nor U10433 (N_10433,N_10381,N_10383);
nor U10434 (N_10434,N_10246,N_10357);
or U10435 (N_10435,N_10334,N_10237);
and U10436 (N_10436,N_10227,N_10225);
or U10437 (N_10437,N_10396,N_10337);
or U10438 (N_10438,N_10231,N_10323);
and U10439 (N_10439,N_10343,N_10322);
nand U10440 (N_10440,N_10219,N_10359);
or U10441 (N_10441,N_10205,N_10398);
or U10442 (N_10442,N_10308,N_10347);
or U10443 (N_10443,N_10258,N_10214);
nand U10444 (N_10444,N_10224,N_10362);
xnor U10445 (N_10445,N_10289,N_10360);
and U10446 (N_10446,N_10262,N_10346);
or U10447 (N_10447,N_10276,N_10336);
xnor U10448 (N_10448,N_10366,N_10248);
xnor U10449 (N_10449,N_10369,N_10242);
xnor U10450 (N_10450,N_10203,N_10293);
nor U10451 (N_10451,N_10327,N_10236);
or U10452 (N_10452,N_10344,N_10391);
and U10453 (N_10453,N_10232,N_10376);
xnor U10454 (N_10454,N_10314,N_10319);
nand U10455 (N_10455,N_10352,N_10226);
or U10456 (N_10456,N_10222,N_10368);
and U10457 (N_10457,N_10331,N_10280);
xor U10458 (N_10458,N_10260,N_10342);
or U10459 (N_10459,N_10374,N_10234);
nand U10460 (N_10460,N_10204,N_10371);
xor U10461 (N_10461,N_10370,N_10392);
or U10462 (N_10462,N_10361,N_10230);
or U10463 (N_10463,N_10305,N_10220);
or U10464 (N_10464,N_10268,N_10393);
nand U10465 (N_10465,N_10241,N_10320);
and U10466 (N_10466,N_10341,N_10372);
nor U10467 (N_10467,N_10264,N_10339);
or U10468 (N_10468,N_10351,N_10287);
nor U10469 (N_10469,N_10253,N_10340);
and U10470 (N_10470,N_10229,N_10333);
or U10471 (N_10471,N_10345,N_10286);
xor U10472 (N_10472,N_10251,N_10283);
nand U10473 (N_10473,N_10208,N_10335);
nor U10474 (N_10474,N_10240,N_10291);
nor U10475 (N_10475,N_10355,N_10202);
nor U10476 (N_10476,N_10252,N_10221);
or U10477 (N_10477,N_10325,N_10254);
or U10478 (N_10478,N_10328,N_10354);
and U10479 (N_10479,N_10298,N_10282);
and U10480 (N_10480,N_10375,N_10279);
nor U10481 (N_10481,N_10312,N_10304);
xor U10482 (N_10482,N_10235,N_10272);
nor U10483 (N_10483,N_10206,N_10297);
xor U10484 (N_10484,N_10329,N_10338);
or U10485 (N_10485,N_10207,N_10309);
and U10486 (N_10486,N_10218,N_10301);
nand U10487 (N_10487,N_10274,N_10259);
or U10488 (N_10488,N_10295,N_10257);
or U10489 (N_10489,N_10326,N_10395);
xor U10490 (N_10490,N_10306,N_10380);
nor U10491 (N_10491,N_10210,N_10310);
or U10492 (N_10492,N_10270,N_10390);
nor U10493 (N_10493,N_10313,N_10317);
xnor U10494 (N_10494,N_10332,N_10290);
nand U10495 (N_10495,N_10244,N_10273);
or U10496 (N_10496,N_10278,N_10365);
nand U10497 (N_10497,N_10377,N_10350);
and U10498 (N_10498,N_10223,N_10266);
nand U10499 (N_10499,N_10296,N_10299);
nand U10500 (N_10500,N_10214,N_10350);
xor U10501 (N_10501,N_10380,N_10242);
nand U10502 (N_10502,N_10340,N_10252);
nand U10503 (N_10503,N_10320,N_10324);
xnor U10504 (N_10504,N_10254,N_10282);
or U10505 (N_10505,N_10224,N_10265);
xnor U10506 (N_10506,N_10200,N_10319);
xnor U10507 (N_10507,N_10247,N_10341);
or U10508 (N_10508,N_10339,N_10356);
nor U10509 (N_10509,N_10211,N_10259);
xnor U10510 (N_10510,N_10225,N_10236);
and U10511 (N_10511,N_10358,N_10340);
nor U10512 (N_10512,N_10284,N_10281);
nor U10513 (N_10513,N_10251,N_10356);
nand U10514 (N_10514,N_10245,N_10398);
xnor U10515 (N_10515,N_10252,N_10251);
nand U10516 (N_10516,N_10326,N_10288);
and U10517 (N_10517,N_10224,N_10268);
xor U10518 (N_10518,N_10223,N_10284);
nand U10519 (N_10519,N_10314,N_10257);
or U10520 (N_10520,N_10253,N_10202);
nand U10521 (N_10521,N_10290,N_10393);
and U10522 (N_10522,N_10394,N_10210);
nand U10523 (N_10523,N_10336,N_10216);
and U10524 (N_10524,N_10296,N_10270);
and U10525 (N_10525,N_10219,N_10226);
nand U10526 (N_10526,N_10314,N_10393);
nand U10527 (N_10527,N_10295,N_10281);
nand U10528 (N_10528,N_10242,N_10253);
nor U10529 (N_10529,N_10244,N_10220);
xor U10530 (N_10530,N_10242,N_10316);
nor U10531 (N_10531,N_10386,N_10282);
xnor U10532 (N_10532,N_10294,N_10393);
or U10533 (N_10533,N_10203,N_10216);
and U10534 (N_10534,N_10207,N_10399);
nor U10535 (N_10535,N_10219,N_10205);
nand U10536 (N_10536,N_10230,N_10227);
or U10537 (N_10537,N_10237,N_10372);
or U10538 (N_10538,N_10253,N_10284);
and U10539 (N_10539,N_10397,N_10307);
xor U10540 (N_10540,N_10362,N_10210);
and U10541 (N_10541,N_10238,N_10327);
or U10542 (N_10542,N_10211,N_10399);
nor U10543 (N_10543,N_10253,N_10322);
nand U10544 (N_10544,N_10346,N_10320);
xnor U10545 (N_10545,N_10287,N_10254);
xor U10546 (N_10546,N_10348,N_10299);
xnor U10547 (N_10547,N_10286,N_10328);
and U10548 (N_10548,N_10278,N_10336);
nand U10549 (N_10549,N_10306,N_10270);
or U10550 (N_10550,N_10201,N_10262);
nor U10551 (N_10551,N_10254,N_10338);
nand U10552 (N_10552,N_10300,N_10374);
nor U10553 (N_10553,N_10340,N_10307);
or U10554 (N_10554,N_10296,N_10211);
and U10555 (N_10555,N_10396,N_10276);
nor U10556 (N_10556,N_10212,N_10320);
nor U10557 (N_10557,N_10300,N_10366);
xor U10558 (N_10558,N_10370,N_10395);
nand U10559 (N_10559,N_10352,N_10278);
or U10560 (N_10560,N_10349,N_10347);
xor U10561 (N_10561,N_10392,N_10368);
or U10562 (N_10562,N_10282,N_10339);
and U10563 (N_10563,N_10227,N_10286);
nor U10564 (N_10564,N_10389,N_10293);
and U10565 (N_10565,N_10256,N_10390);
xnor U10566 (N_10566,N_10376,N_10336);
and U10567 (N_10567,N_10232,N_10380);
nand U10568 (N_10568,N_10397,N_10267);
and U10569 (N_10569,N_10225,N_10310);
xnor U10570 (N_10570,N_10395,N_10364);
or U10571 (N_10571,N_10271,N_10300);
or U10572 (N_10572,N_10329,N_10267);
xnor U10573 (N_10573,N_10253,N_10392);
or U10574 (N_10574,N_10329,N_10377);
xnor U10575 (N_10575,N_10366,N_10265);
and U10576 (N_10576,N_10319,N_10371);
and U10577 (N_10577,N_10270,N_10264);
and U10578 (N_10578,N_10359,N_10337);
nor U10579 (N_10579,N_10356,N_10357);
and U10580 (N_10580,N_10384,N_10222);
nand U10581 (N_10581,N_10236,N_10234);
and U10582 (N_10582,N_10324,N_10298);
xnor U10583 (N_10583,N_10380,N_10296);
xnor U10584 (N_10584,N_10326,N_10273);
and U10585 (N_10585,N_10236,N_10224);
or U10586 (N_10586,N_10254,N_10208);
nor U10587 (N_10587,N_10312,N_10248);
nor U10588 (N_10588,N_10344,N_10334);
or U10589 (N_10589,N_10342,N_10350);
and U10590 (N_10590,N_10203,N_10279);
or U10591 (N_10591,N_10215,N_10311);
or U10592 (N_10592,N_10307,N_10371);
nand U10593 (N_10593,N_10208,N_10274);
nand U10594 (N_10594,N_10255,N_10249);
nor U10595 (N_10595,N_10303,N_10386);
and U10596 (N_10596,N_10331,N_10210);
xor U10597 (N_10597,N_10276,N_10242);
nand U10598 (N_10598,N_10228,N_10211);
nand U10599 (N_10599,N_10363,N_10257);
nand U10600 (N_10600,N_10495,N_10435);
xor U10601 (N_10601,N_10523,N_10477);
and U10602 (N_10602,N_10588,N_10479);
or U10603 (N_10603,N_10563,N_10455);
or U10604 (N_10604,N_10529,N_10522);
or U10605 (N_10605,N_10545,N_10508);
xnor U10606 (N_10606,N_10587,N_10473);
nor U10607 (N_10607,N_10555,N_10505);
xor U10608 (N_10608,N_10461,N_10576);
or U10609 (N_10609,N_10440,N_10472);
xnor U10610 (N_10610,N_10598,N_10497);
nand U10611 (N_10611,N_10415,N_10401);
or U10612 (N_10612,N_10542,N_10402);
xnor U10613 (N_10613,N_10426,N_10492);
xnor U10614 (N_10614,N_10457,N_10501);
xor U10615 (N_10615,N_10458,N_10411);
xor U10616 (N_10616,N_10570,N_10488);
xnor U10617 (N_10617,N_10417,N_10575);
xnor U10618 (N_10618,N_10527,N_10447);
nor U10619 (N_10619,N_10443,N_10595);
nand U10620 (N_10620,N_10537,N_10424);
nand U10621 (N_10621,N_10483,N_10528);
xnor U10622 (N_10622,N_10553,N_10539);
xor U10623 (N_10623,N_10552,N_10400);
nor U10624 (N_10624,N_10409,N_10407);
nand U10625 (N_10625,N_10408,N_10504);
nand U10626 (N_10626,N_10583,N_10487);
nand U10627 (N_10627,N_10469,N_10464);
and U10628 (N_10628,N_10590,N_10456);
xnor U10629 (N_10629,N_10574,N_10466);
or U10630 (N_10630,N_10470,N_10453);
nor U10631 (N_10631,N_10586,N_10511);
nand U10632 (N_10632,N_10538,N_10556);
nor U10633 (N_10633,N_10571,N_10494);
and U10634 (N_10634,N_10418,N_10599);
and U10635 (N_10635,N_10549,N_10567);
nor U10636 (N_10636,N_10413,N_10503);
and U10637 (N_10637,N_10580,N_10450);
xor U10638 (N_10638,N_10547,N_10510);
and U10639 (N_10639,N_10517,N_10565);
nor U10640 (N_10640,N_10568,N_10428);
nor U10641 (N_10641,N_10582,N_10591);
or U10642 (N_10642,N_10405,N_10442);
nand U10643 (N_10643,N_10560,N_10467);
and U10644 (N_10644,N_10445,N_10562);
and U10645 (N_10645,N_10515,N_10481);
xnor U10646 (N_10646,N_10584,N_10451);
nand U10647 (N_10647,N_10500,N_10594);
and U10648 (N_10648,N_10530,N_10578);
nor U10649 (N_10649,N_10577,N_10536);
xor U10650 (N_10650,N_10403,N_10437);
or U10651 (N_10651,N_10518,N_10564);
xnor U10652 (N_10652,N_10410,N_10533);
nand U10653 (N_10653,N_10558,N_10439);
nand U10654 (N_10654,N_10434,N_10561);
or U10655 (N_10655,N_10532,N_10507);
and U10656 (N_10656,N_10460,N_10416);
or U10657 (N_10657,N_10482,N_10448);
and U10658 (N_10658,N_10454,N_10490);
nor U10659 (N_10659,N_10573,N_10569);
or U10660 (N_10660,N_10420,N_10431);
and U10661 (N_10661,N_10513,N_10412);
or U10662 (N_10662,N_10491,N_10476);
nor U10663 (N_10663,N_10519,N_10592);
xnor U10664 (N_10664,N_10444,N_10496);
nor U10665 (N_10665,N_10534,N_10452);
nor U10666 (N_10666,N_10463,N_10572);
xor U10667 (N_10667,N_10535,N_10581);
nand U10668 (N_10668,N_10579,N_10484);
nand U10669 (N_10669,N_10478,N_10512);
nand U10670 (N_10670,N_10526,N_10427);
xor U10671 (N_10671,N_10414,N_10548);
nand U10672 (N_10672,N_10421,N_10429);
and U10673 (N_10673,N_10589,N_10433);
and U10674 (N_10674,N_10502,N_10509);
and U10675 (N_10675,N_10459,N_10471);
or U10676 (N_10676,N_10506,N_10546);
nand U10677 (N_10677,N_10423,N_10551);
or U10678 (N_10678,N_10499,N_10449);
and U10679 (N_10679,N_10468,N_10486);
nand U10680 (N_10680,N_10430,N_10525);
xor U10681 (N_10681,N_10489,N_10566);
xor U10682 (N_10682,N_10465,N_10485);
nor U10683 (N_10683,N_10446,N_10480);
and U10684 (N_10684,N_10540,N_10543);
nand U10685 (N_10685,N_10531,N_10554);
or U10686 (N_10686,N_10593,N_10550);
nand U10687 (N_10687,N_10425,N_10514);
and U10688 (N_10688,N_10521,N_10475);
nor U10689 (N_10689,N_10438,N_10432);
and U10690 (N_10690,N_10544,N_10419);
xor U10691 (N_10691,N_10436,N_10498);
xnor U10692 (N_10692,N_10524,N_10493);
xnor U10693 (N_10693,N_10516,N_10404);
nand U10694 (N_10694,N_10462,N_10422);
nand U10695 (N_10695,N_10585,N_10520);
nand U10696 (N_10696,N_10559,N_10597);
nand U10697 (N_10697,N_10441,N_10596);
nor U10698 (N_10698,N_10474,N_10557);
and U10699 (N_10699,N_10406,N_10541);
or U10700 (N_10700,N_10443,N_10579);
nand U10701 (N_10701,N_10422,N_10565);
or U10702 (N_10702,N_10460,N_10540);
or U10703 (N_10703,N_10503,N_10599);
and U10704 (N_10704,N_10510,N_10447);
and U10705 (N_10705,N_10564,N_10541);
nand U10706 (N_10706,N_10425,N_10436);
nand U10707 (N_10707,N_10498,N_10400);
nand U10708 (N_10708,N_10575,N_10452);
and U10709 (N_10709,N_10474,N_10465);
nor U10710 (N_10710,N_10422,N_10513);
xor U10711 (N_10711,N_10568,N_10569);
and U10712 (N_10712,N_10571,N_10486);
and U10713 (N_10713,N_10449,N_10514);
or U10714 (N_10714,N_10493,N_10446);
nor U10715 (N_10715,N_10486,N_10563);
xor U10716 (N_10716,N_10496,N_10508);
nor U10717 (N_10717,N_10535,N_10465);
nor U10718 (N_10718,N_10507,N_10588);
and U10719 (N_10719,N_10536,N_10497);
nand U10720 (N_10720,N_10426,N_10448);
nand U10721 (N_10721,N_10432,N_10568);
nand U10722 (N_10722,N_10451,N_10596);
xor U10723 (N_10723,N_10458,N_10457);
or U10724 (N_10724,N_10476,N_10474);
nand U10725 (N_10725,N_10558,N_10404);
xor U10726 (N_10726,N_10438,N_10447);
xor U10727 (N_10727,N_10570,N_10551);
and U10728 (N_10728,N_10503,N_10554);
nor U10729 (N_10729,N_10491,N_10445);
and U10730 (N_10730,N_10408,N_10498);
xor U10731 (N_10731,N_10424,N_10430);
or U10732 (N_10732,N_10404,N_10461);
and U10733 (N_10733,N_10579,N_10536);
nand U10734 (N_10734,N_10405,N_10489);
or U10735 (N_10735,N_10449,N_10573);
nand U10736 (N_10736,N_10599,N_10583);
and U10737 (N_10737,N_10437,N_10460);
nand U10738 (N_10738,N_10480,N_10562);
nand U10739 (N_10739,N_10593,N_10592);
xor U10740 (N_10740,N_10507,N_10448);
nor U10741 (N_10741,N_10430,N_10562);
and U10742 (N_10742,N_10472,N_10414);
and U10743 (N_10743,N_10499,N_10402);
xnor U10744 (N_10744,N_10491,N_10453);
nor U10745 (N_10745,N_10464,N_10567);
xor U10746 (N_10746,N_10544,N_10467);
or U10747 (N_10747,N_10447,N_10405);
and U10748 (N_10748,N_10480,N_10452);
nor U10749 (N_10749,N_10568,N_10514);
nand U10750 (N_10750,N_10585,N_10535);
nor U10751 (N_10751,N_10466,N_10544);
and U10752 (N_10752,N_10412,N_10564);
or U10753 (N_10753,N_10451,N_10416);
xnor U10754 (N_10754,N_10570,N_10546);
and U10755 (N_10755,N_10516,N_10466);
or U10756 (N_10756,N_10412,N_10515);
and U10757 (N_10757,N_10577,N_10461);
nand U10758 (N_10758,N_10547,N_10577);
nor U10759 (N_10759,N_10466,N_10533);
and U10760 (N_10760,N_10596,N_10564);
nor U10761 (N_10761,N_10535,N_10491);
xnor U10762 (N_10762,N_10464,N_10570);
xnor U10763 (N_10763,N_10466,N_10416);
xnor U10764 (N_10764,N_10417,N_10469);
xor U10765 (N_10765,N_10494,N_10550);
xnor U10766 (N_10766,N_10428,N_10517);
nand U10767 (N_10767,N_10506,N_10545);
nand U10768 (N_10768,N_10560,N_10565);
xor U10769 (N_10769,N_10559,N_10507);
and U10770 (N_10770,N_10581,N_10437);
nor U10771 (N_10771,N_10589,N_10463);
nand U10772 (N_10772,N_10464,N_10414);
nor U10773 (N_10773,N_10416,N_10518);
and U10774 (N_10774,N_10527,N_10569);
nor U10775 (N_10775,N_10449,N_10595);
nand U10776 (N_10776,N_10444,N_10423);
xor U10777 (N_10777,N_10479,N_10524);
and U10778 (N_10778,N_10518,N_10500);
and U10779 (N_10779,N_10589,N_10554);
nor U10780 (N_10780,N_10491,N_10401);
nand U10781 (N_10781,N_10582,N_10586);
or U10782 (N_10782,N_10423,N_10493);
nand U10783 (N_10783,N_10455,N_10501);
or U10784 (N_10784,N_10474,N_10592);
or U10785 (N_10785,N_10479,N_10473);
or U10786 (N_10786,N_10429,N_10550);
nor U10787 (N_10787,N_10401,N_10468);
xor U10788 (N_10788,N_10484,N_10458);
nand U10789 (N_10789,N_10502,N_10430);
nor U10790 (N_10790,N_10458,N_10468);
nor U10791 (N_10791,N_10483,N_10557);
xnor U10792 (N_10792,N_10525,N_10556);
nand U10793 (N_10793,N_10474,N_10532);
and U10794 (N_10794,N_10531,N_10595);
nand U10795 (N_10795,N_10447,N_10422);
nor U10796 (N_10796,N_10492,N_10475);
nor U10797 (N_10797,N_10544,N_10532);
nand U10798 (N_10798,N_10532,N_10522);
xnor U10799 (N_10799,N_10433,N_10460);
and U10800 (N_10800,N_10723,N_10625);
and U10801 (N_10801,N_10765,N_10712);
or U10802 (N_10802,N_10793,N_10711);
nand U10803 (N_10803,N_10717,N_10745);
nor U10804 (N_10804,N_10726,N_10718);
nand U10805 (N_10805,N_10725,N_10759);
xnor U10806 (N_10806,N_10611,N_10747);
or U10807 (N_10807,N_10630,N_10710);
xor U10808 (N_10808,N_10665,N_10795);
xnor U10809 (N_10809,N_10781,N_10637);
nand U10810 (N_10810,N_10790,N_10771);
xor U10811 (N_10811,N_10691,N_10604);
nor U10812 (N_10812,N_10758,N_10743);
or U10813 (N_10813,N_10640,N_10739);
and U10814 (N_10814,N_10660,N_10748);
and U10815 (N_10815,N_10667,N_10621);
nor U10816 (N_10816,N_10693,N_10638);
or U10817 (N_10817,N_10688,N_10609);
nor U10818 (N_10818,N_10624,N_10680);
xor U10819 (N_10819,N_10631,N_10618);
nand U10820 (N_10820,N_10794,N_10755);
or U10821 (N_10821,N_10720,N_10656);
xor U10822 (N_10822,N_10735,N_10601);
xor U10823 (N_10823,N_10605,N_10746);
or U10824 (N_10824,N_10686,N_10700);
or U10825 (N_10825,N_10616,N_10778);
nand U10826 (N_10826,N_10791,N_10713);
nand U10827 (N_10827,N_10756,N_10652);
or U10828 (N_10828,N_10776,N_10669);
xor U10829 (N_10829,N_10732,N_10648);
and U10830 (N_10830,N_10753,N_10751);
xor U10831 (N_10831,N_10600,N_10785);
or U10832 (N_10832,N_10639,N_10658);
and U10833 (N_10833,N_10727,N_10644);
nor U10834 (N_10834,N_10788,N_10699);
or U10835 (N_10835,N_10768,N_10733);
nand U10836 (N_10836,N_10608,N_10653);
or U10837 (N_10837,N_10615,N_10642);
or U10838 (N_10838,N_10687,N_10650);
xnor U10839 (N_10839,N_10606,N_10602);
nand U10840 (N_10840,N_10620,N_10729);
xor U10841 (N_10841,N_10782,N_10709);
nand U10842 (N_10842,N_10666,N_10623);
nand U10843 (N_10843,N_10626,N_10744);
or U10844 (N_10844,N_10677,N_10654);
and U10845 (N_10845,N_10651,N_10668);
xnor U10846 (N_10846,N_10766,N_10634);
nand U10847 (N_10847,N_10610,N_10683);
nand U10848 (N_10848,N_10672,N_10730);
xnor U10849 (N_10849,N_10645,N_10731);
nor U10850 (N_10850,N_10749,N_10622);
nand U10851 (N_10851,N_10689,N_10763);
nand U10852 (N_10852,N_10724,N_10646);
nor U10853 (N_10853,N_10603,N_10696);
xor U10854 (N_10854,N_10772,N_10673);
xnor U10855 (N_10855,N_10767,N_10780);
or U10856 (N_10856,N_10679,N_10722);
or U10857 (N_10857,N_10671,N_10742);
xor U10858 (N_10858,N_10779,N_10761);
xor U10859 (N_10859,N_10705,N_10787);
and U10860 (N_10860,N_10789,N_10632);
and U10861 (N_10861,N_10777,N_10760);
and U10862 (N_10862,N_10773,N_10738);
nand U10863 (N_10863,N_10786,N_10661);
or U10864 (N_10864,N_10647,N_10714);
nand U10865 (N_10865,N_10670,N_10678);
xnor U10866 (N_10866,N_10681,N_10614);
or U10867 (N_10867,N_10757,N_10784);
xor U10868 (N_10868,N_10641,N_10740);
xnor U10869 (N_10869,N_10764,N_10702);
nor U10870 (N_10870,N_10697,N_10690);
nand U10871 (N_10871,N_10792,N_10701);
xor U10872 (N_10872,N_10741,N_10695);
or U10873 (N_10873,N_10685,N_10635);
nand U10874 (N_10874,N_10612,N_10694);
nand U10875 (N_10875,N_10775,N_10704);
or U10876 (N_10876,N_10716,N_10662);
or U10877 (N_10877,N_10675,N_10737);
and U10878 (N_10878,N_10736,N_10728);
and U10879 (N_10879,N_10796,N_10770);
xor U10880 (N_10880,N_10798,N_10762);
xor U10881 (N_10881,N_10684,N_10707);
xnor U10882 (N_10882,N_10643,N_10636);
xnor U10883 (N_10883,N_10628,N_10619);
or U10884 (N_10884,N_10674,N_10692);
nor U10885 (N_10885,N_10719,N_10715);
nor U10886 (N_10886,N_10657,N_10783);
or U10887 (N_10887,N_10613,N_10698);
or U10888 (N_10888,N_10734,N_10708);
or U10889 (N_10889,N_10633,N_10655);
nand U10890 (N_10890,N_10752,N_10721);
or U10891 (N_10891,N_10797,N_10703);
and U10892 (N_10892,N_10676,N_10617);
or U10893 (N_10893,N_10769,N_10664);
nor U10894 (N_10894,N_10750,N_10774);
nor U10895 (N_10895,N_10706,N_10627);
or U10896 (N_10896,N_10607,N_10663);
nor U10897 (N_10897,N_10659,N_10754);
xor U10898 (N_10898,N_10682,N_10629);
nand U10899 (N_10899,N_10799,N_10649);
and U10900 (N_10900,N_10762,N_10677);
nor U10901 (N_10901,N_10647,N_10614);
and U10902 (N_10902,N_10785,N_10797);
nor U10903 (N_10903,N_10729,N_10647);
xnor U10904 (N_10904,N_10777,N_10695);
xnor U10905 (N_10905,N_10681,N_10698);
nand U10906 (N_10906,N_10745,N_10708);
and U10907 (N_10907,N_10718,N_10732);
and U10908 (N_10908,N_10766,N_10781);
xnor U10909 (N_10909,N_10600,N_10730);
xnor U10910 (N_10910,N_10653,N_10615);
xor U10911 (N_10911,N_10767,N_10732);
xnor U10912 (N_10912,N_10682,N_10723);
xor U10913 (N_10913,N_10790,N_10688);
nor U10914 (N_10914,N_10721,N_10676);
nand U10915 (N_10915,N_10704,N_10780);
nor U10916 (N_10916,N_10661,N_10714);
xor U10917 (N_10917,N_10616,N_10766);
or U10918 (N_10918,N_10774,N_10730);
nand U10919 (N_10919,N_10615,N_10744);
nand U10920 (N_10920,N_10767,N_10638);
nor U10921 (N_10921,N_10686,N_10757);
nand U10922 (N_10922,N_10758,N_10733);
or U10923 (N_10923,N_10714,N_10611);
xnor U10924 (N_10924,N_10678,N_10640);
xnor U10925 (N_10925,N_10761,N_10728);
nand U10926 (N_10926,N_10786,N_10688);
and U10927 (N_10927,N_10705,N_10759);
and U10928 (N_10928,N_10759,N_10651);
and U10929 (N_10929,N_10669,N_10795);
or U10930 (N_10930,N_10704,N_10680);
xor U10931 (N_10931,N_10792,N_10697);
or U10932 (N_10932,N_10680,N_10636);
and U10933 (N_10933,N_10715,N_10700);
nand U10934 (N_10934,N_10769,N_10771);
nand U10935 (N_10935,N_10670,N_10611);
and U10936 (N_10936,N_10742,N_10789);
nand U10937 (N_10937,N_10642,N_10681);
nand U10938 (N_10938,N_10784,N_10680);
or U10939 (N_10939,N_10759,N_10672);
xnor U10940 (N_10940,N_10643,N_10764);
or U10941 (N_10941,N_10704,N_10762);
nor U10942 (N_10942,N_10687,N_10751);
and U10943 (N_10943,N_10663,N_10711);
or U10944 (N_10944,N_10650,N_10717);
or U10945 (N_10945,N_10728,N_10629);
nor U10946 (N_10946,N_10794,N_10685);
nor U10947 (N_10947,N_10762,N_10676);
and U10948 (N_10948,N_10671,N_10633);
or U10949 (N_10949,N_10761,N_10644);
nand U10950 (N_10950,N_10646,N_10601);
xnor U10951 (N_10951,N_10786,N_10680);
and U10952 (N_10952,N_10662,N_10617);
nand U10953 (N_10953,N_10606,N_10695);
nor U10954 (N_10954,N_10792,N_10612);
xnor U10955 (N_10955,N_10626,N_10714);
nand U10956 (N_10956,N_10659,N_10643);
xnor U10957 (N_10957,N_10617,N_10780);
or U10958 (N_10958,N_10685,N_10713);
nand U10959 (N_10959,N_10719,N_10780);
nand U10960 (N_10960,N_10745,N_10615);
xnor U10961 (N_10961,N_10796,N_10716);
xnor U10962 (N_10962,N_10633,N_10791);
nand U10963 (N_10963,N_10697,N_10740);
nand U10964 (N_10964,N_10719,N_10659);
xor U10965 (N_10965,N_10686,N_10620);
nand U10966 (N_10966,N_10604,N_10666);
and U10967 (N_10967,N_10734,N_10658);
xnor U10968 (N_10968,N_10704,N_10690);
xnor U10969 (N_10969,N_10733,N_10629);
or U10970 (N_10970,N_10790,N_10613);
nor U10971 (N_10971,N_10739,N_10787);
xnor U10972 (N_10972,N_10786,N_10757);
or U10973 (N_10973,N_10624,N_10658);
nand U10974 (N_10974,N_10735,N_10747);
nor U10975 (N_10975,N_10792,N_10750);
nor U10976 (N_10976,N_10606,N_10680);
and U10977 (N_10977,N_10612,N_10624);
or U10978 (N_10978,N_10681,N_10765);
and U10979 (N_10979,N_10645,N_10688);
nor U10980 (N_10980,N_10613,N_10634);
xnor U10981 (N_10981,N_10630,N_10768);
or U10982 (N_10982,N_10791,N_10653);
xnor U10983 (N_10983,N_10605,N_10781);
nor U10984 (N_10984,N_10760,N_10694);
or U10985 (N_10985,N_10673,N_10659);
or U10986 (N_10986,N_10744,N_10777);
xnor U10987 (N_10987,N_10798,N_10745);
xnor U10988 (N_10988,N_10759,N_10631);
nor U10989 (N_10989,N_10777,N_10609);
nand U10990 (N_10990,N_10759,N_10778);
xnor U10991 (N_10991,N_10703,N_10627);
and U10992 (N_10992,N_10643,N_10674);
nor U10993 (N_10993,N_10664,N_10658);
nor U10994 (N_10994,N_10733,N_10690);
xnor U10995 (N_10995,N_10757,N_10795);
nand U10996 (N_10996,N_10615,N_10711);
and U10997 (N_10997,N_10654,N_10777);
or U10998 (N_10998,N_10755,N_10696);
nor U10999 (N_10999,N_10787,N_10729);
or U11000 (N_11000,N_10877,N_10830);
xor U11001 (N_11001,N_10868,N_10976);
nor U11002 (N_11002,N_10948,N_10867);
and U11003 (N_11003,N_10930,N_10824);
or U11004 (N_11004,N_10869,N_10981);
and U11005 (N_11005,N_10967,N_10907);
or U11006 (N_11006,N_10841,N_10968);
and U11007 (N_11007,N_10989,N_10982);
nor U11008 (N_11008,N_10875,N_10939);
and U11009 (N_11009,N_10924,N_10984);
and U11010 (N_11010,N_10823,N_10935);
xor U11011 (N_11011,N_10918,N_10892);
nand U11012 (N_11012,N_10912,N_10945);
nor U11013 (N_11013,N_10958,N_10896);
nor U11014 (N_11014,N_10931,N_10809);
and U11015 (N_11015,N_10842,N_10920);
xnor U11016 (N_11016,N_10906,N_10897);
nor U11017 (N_11017,N_10942,N_10934);
nor U11018 (N_11018,N_10946,N_10847);
and U11019 (N_11019,N_10802,N_10940);
and U11020 (N_11020,N_10889,N_10966);
nand U11021 (N_11021,N_10998,N_10825);
nand U11022 (N_11022,N_10890,N_10969);
nand U11023 (N_11023,N_10900,N_10804);
or U11024 (N_11024,N_10808,N_10941);
nor U11025 (N_11025,N_10950,N_10929);
and U11026 (N_11026,N_10973,N_10836);
xor U11027 (N_11027,N_10947,N_10944);
and U11028 (N_11028,N_10811,N_10894);
or U11029 (N_11029,N_10840,N_10974);
nor U11030 (N_11030,N_10845,N_10937);
nor U11031 (N_11031,N_10972,N_10881);
and U11032 (N_11032,N_10904,N_10844);
and U11033 (N_11033,N_10949,N_10861);
and U11034 (N_11034,N_10835,N_10990);
and U11035 (N_11035,N_10873,N_10913);
and U11036 (N_11036,N_10880,N_10905);
nor U11037 (N_11037,N_10848,N_10955);
nor U11038 (N_11038,N_10843,N_10957);
nand U11039 (N_11039,N_10870,N_10928);
or U11040 (N_11040,N_10985,N_10916);
and U11041 (N_11041,N_10908,N_10979);
xnor U11042 (N_11042,N_10999,N_10882);
xnor U11043 (N_11043,N_10962,N_10895);
xnor U11044 (N_11044,N_10864,N_10862);
or U11045 (N_11045,N_10991,N_10986);
or U11046 (N_11046,N_10883,N_10810);
and U11047 (N_11047,N_10860,N_10901);
xor U11048 (N_11048,N_10997,N_10954);
nand U11049 (N_11049,N_10878,N_10884);
xor U11050 (N_11050,N_10831,N_10938);
and U11051 (N_11051,N_10888,N_10933);
xnor U11052 (N_11052,N_10874,N_10837);
nand U11053 (N_11053,N_10826,N_10818);
nor U11054 (N_11054,N_10953,N_10995);
or U11055 (N_11055,N_10801,N_10885);
or U11056 (N_11056,N_10866,N_10872);
nor U11057 (N_11057,N_10812,N_10978);
nor U11058 (N_11058,N_10876,N_10919);
nor U11059 (N_11059,N_10932,N_10921);
and U11060 (N_11060,N_10980,N_10850);
and U11061 (N_11061,N_10902,N_10983);
and U11062 (N_11062,N_10816,N_10909);
nand U11063 (N_11063,N_10833,N_10800);
nor U11064 (N_11064,N_10926,N_10923);
or U11065 (N_11065,N_10858,N_10822);
xor U11066 (N_11066,N_10834,N_10846);
and U11067 (N_11067,N_10956,N_10879);
and U11068 (N_11068,N_10917,N_10815);
or U11069 (N_11069,N_10855,N_10849);
and U11070 (N_11070,N_10922,N_10857);
xor U11071 (N_11071,N_10887,N_10854);
xor U11072 (N_11072,N_10893,N_10963);
and U11073 (N_11073,N_10865,N_10817);
nor U11074 (N_11074,N_10915,N_10829);
nor U11075 (N_11075,N_10975,N_10851);
or U11076 (N_11076,N_10853,N_10961);
or U11077 (N_11077,N_10891,N_10943);
nand U11078 (N_11078,N_10988,N_10952);
nor U11079 (N_11079,N_10993,N_10838);
nor U11080 (N_11080,N_10960,N_10959);
nand U11081 (N_11081,N_10820,N_10827);
xnor U11082 (N_11082,N_10936,N_10898);
nor U11083 (N_11083,N_10852,N_10821);
or U11084 (N_11084,N_10911,N_10806);
or U11085 (N_11085,N_10992,N_10927);
xnor U11086 (N_11086,N_10925,N_10828);
xor U11087 (N_11087,N_10977,N_10805);
nor U11088 (N_11088,N_10871,N_10832);
nand U11089 (N_11089,N_10863,N_10859);
nor U11090 (N_11090,N_10951,N_10856);
and U11091 (N_11091,N_10839,N_10814);
nor U11092 (N_11092,N_10914,N_10886);
or U11093 (N_11093,N_10994,N_10971);
xnor U11094 (N_11094,N_10813,N_10819);
xnor U11095 (N_11095,N_10964,N_10965);
and U11096 (N_11096,N_10899,N_10903);
and U11097 (N_11097,N_10996,N_10987);
or U11098 (N_11098,N_10910,N_10970);
and U11099 (N_11099,N_10803,N_10807);
nor U11100 (N_11100,N_10884,N_10951);
xor U11101 (N_11101,N_10892,N_10945);
or U11102 (N_11102,N_10808,N_10880);
and U11103 (N_11103,N_10865,N_10926);
and U11104 (N_11104,N_10979,N_10954);
or U11105 (N_11105,N_10890,N_10868);
and U11106 (N_11106,N_10910,N_10964);
xnor U11107 (N_11107,N_10944,N_10885);
nor U11108 (N_11108,N_10817,N_10910);
xor U11109 (N_11109,N_10940,N_10925);
nand U11110 (N_11110,N_10965,N_10827);
and U11111 (N_11111,N_10848,N_10947);
nand U11112 (N_11112,N_10849,N_10966);
and U11113 (N_11113,N_10914,N_10860);
and U11114 (N_11114,N_10886,N_10912);
nor U11115 (N_11115,N_10837,N_10890);
and U11116 (N_11116,N_10912,N_10889);
and U11117 (N_11117,N_10962,N_10804);
nand U11118 (N_11118,N_10924,N_10881);
nor U11119 (N_11119,N_10835,N_10974);
nor U11120 (N_11120,N_10860,N_10975);
nand U11121 (N_11121,N_10812,N_10899);
or U11122 (N_11122,N_10830,N_10867);
and U11123 (N_11123,N_10878,N_10838);
nand U11124 (N_11124,N_10857,N_10865);
or U11125 (N_11125,N_10921,N_10928);
nand U11126 (N_11126,N_10968,N_10862);
nand U11127 (N_11127,N_10893,N_10928);
xor U11128 (N_11128,N_10891,N_10918);
nand U11129 (N_11129,N_10879,N_10848);
nor U11130 (N_11130,N_10881,N_10839);
or U11131 (N_11131,N_10936,N_10960);
xor U11132 (N_11132,N_10883,N_10862);
nor U11133 (N_11133,N_10866,N_10865);
and U11134 (N_11134,N_10993,N_10980);
nand U11135 (N_11135,N_10839,N_10810);
or U11136 (N_11136,N_10937,N_10855);
nor U11137 (N_11137,N_10827,N_10991);
and U11138 (N_11138,N_10946,N_10871);
nand U11139 (N_11139,N_10936,N_10849);
or U11140 (N_11140,N_10844,N_10936);
nand U11141 (N_11141,N_10857,N_10877);
nand U11142 (N_11142,N_10951,N_10875);
xnor U11143 (N_11143,N_10927,N_10856);
nand U11144 (N_11144,N_10994,N_10906);
nand U11145 (N_11145,N_10932,N_10901);
nand U11146 (N_11146,N_10958,N_10801);
and U11147 (N_11147,N_10895,N_10873);
nor U11148 (N_11148,N_10816,N_10994);
and U11149 (N_11149,N_10973,N_10810);
xor U11150 (N_11150,N_10825,N_10833);
or U11151 (N_11151,N_10807,N_10907);
and U11152 (N_11152,N_10932,N_10969);
nor U11153 (N_11153,N_10857,N_10946);
nor U11154 (N_11154,N_10945,N_10981);
and U11155 (N_11155,N_10817,N_10978);
and U11156 (N_11156,N_10979,N_10815);
or U11157 (N_11157,N_10920,N_10959);
nor U11158 (N_11158,N_10874,N_10984);
nand U11159 (N_11159,N_10998,N_10888);
and U11160 (N_11160,N_10949,N_10924);
or U11161 (N_11161,N_10964,N_10841);
xor U11162 (N_11162,N_10930,N_10915);
or U11163 (N_11163,N_10937,N_10948);
or U11164 (N_11164,N_10975,N_10973);
xnor U11165 (N_11165,N_10807,N_10877);
and U11166 (N_11166,N_10904,N_10952);
xnor U11167 (N_11167,N_10956,N_10915);
and U11168 (N_11168,N_10860,N_10909);
nand U11169 (N_11169,N_10942,N_10958);
xnor U11170 (N_11170,N_10938,N_10986);
or U11171 (N_11171,N_10984,N_10858);
or U11172 (N_11172,N_10976,N_10826);
or U11173 (N_11173,N_10859,N_10815);
nand U11174 (N_11174,N_10989,N_10818);
and U11175 (N_11175,N_10995,N_10810);
or U11176 (N_11176,N_10921,N_10948);
nand U11177 (N_11177,N_10898,N_10820);
nand U11178 (N_11178,N_10996,N_10971);
or U11179 (N_11179,N_10907,N_10864);
or U11180 (N_11180,N_10831,N_10983);
nand U11181 (N_11181,N_10842,N_10915);
xor U11182 (N_11182,N_10886,N_10844);
nor U11183 (N_11183,N_10967,N_10906);
nor U11184 (N_11184,N_10954,N_10910);
and U11185 (N_11185,N_10937,N_10930);
and U11186 (N_11186,N_10975,N_10903);
nor U11187 (N_11187,N_10921,N_10855);
or U11188 (N_11188,N_10883,N_10828);
and U11189 (N_11189,N_10962,N_10844);
nor U11190 (N_11190,N_10954,N_10820);
or U11191 (N_11191,N_10974,N_10843);
xnor U11192 (N_11192,N_10848,N_10840);
nor U11193 (N_11193,N_10813,N_10995);
nand U11194 (N_11194,N_10880,N_10833);
nor U11195 (N_11195,N_10806,N_10803);
xor U11196 (N_11196,N_10806,N_10809);
or U11197 (N_11197,N_10908,N_10832);
and U11198 (N_11198,N_10857,N_10916);
xnor U11199 (N_11199,N_10865,N_10955);
and U11200 (N_11200,N_11000,N_11051);
xor U11201 (N_11201,N_11168,N_11067);
nor U11202 (N_11202,N_11006,N_11043);
nand U11203 (N_11203,N_11106,N_11027);
nor U11204 (N_11204,N_11145,N_11012);
xnor U11205 (N_11205,N_11198,N_11116);
or U11206 (N_11206,N_11005,N_11050);
xnor U11207 (N_11207,N_11034,N_11042);
and U11208 (N_11208,N_11079,N_11010);
or U11209 (N_11209,N_11008,N_11038);
or U11210 (N_11210,N_11192,N_11171);
or U11211 (N_11211,N_11052,N_11100);
nor U11212 (N_11212,N_11046,N_11133);
or U11213 (N_11213,N_11189,N_11071);
or U11214 (N_11214,N_11144,N_11172);
nor U11215 (N_11215,N_11176,N_11056);
and U11216 (N_11216,N_11011,N_11124);
nor U11217 (N_11217,N_11064,N_11066);
nor U11218 (N_11218,N_11199,N_11140);
nand U11219 (N_11219,N_11060,N_11151);
nand U11220 (N_11220,N_11030,N_11069);
xnor U11221 (N_11221,N_11161,N_11036);
nor U11222 (N_11222,N_11091,N_11016);
nand U11223 (N_11223,N_11033,N_11087);
nand U11224 (N_11224,N_11125,N_11021);
nand U11225 (N_11225,N_11175,N_11196);
nor U11226 (N_11226,N_11102,N_11024);
or U11227 (N_11227,N_11132,N_11174);
and U11228 (N_11228,N_11009,N_11096);
or U11229 (N_11229,N_11049,N_11197);
nand U11230 (N_11230,N_11081,N_11154);
or U11231 (N_11231,N_11156,N_11029);
nand U11232 (N_11232,N_11022,N_11111);
xnor U11233 (N_11233,N_11083,N_11099);
nand U11234 (N_11234,N_11195,N_11084);
or U11235 (N_11235,N_11184,N_11004);
nand U11236 (N_11236,N_11044,N_11028);
or U11237 (N_11237,N_11191,N_11164);
xor U11238 (N_11238,N_11138,N_11158);
nor U11239 (N_11239,N_11101,N_11163);
xor U11240 (N_11240,N_11026,N_11153);
or U11241 (N_11241,N_11186,N_11014);
or U11242 (N_11242,N_11058,N_11020);
nor U11243 (N_11243,N_11182,N_11121);
and U11244 (N_11244,N_11115,N_11035);
nor U11245 (N_11245,N_11090,N_11107);
nand U11246 (N_11246,N_11147,N_11047);
or U11247 (N_11247,N_11041,N_11149);
or U11248 (N_11248,N_11135,N_11080);
xnor U11249 (N_11249,N_11003,N_11025);
nor U11250 (N_11250,N_11007,N_11037);
nand U11251 (N_11251,N_11122,N_11159);
or U11252 (N_11252,N_11190,N_11136);
xor U11253 (N_11253,N_11039,N_11059);
nor U11254 (N_11254,N_11155,N_11150);
nand U11255 (N_11255,N_11188,N_11181);
and U11256 (N_11256,N_11131,N_11143);
nor U11257 (N_11257,N_11119,N_11180);
nor U11258 (N_11258,N_11166,N_11097);
nor U11259 (N_11259,N_11194,N_11086);
nand U11260 (N_11260,N_11117,N_11193);
and U11261 (N_11261,N_11109,N_11078);
xor U11262 (N_11262,N_11183,N_11152);
and U11263 (N_11263,N_11141,N_11054);
or U11264 (N_11264,N_11173,N_11123);
xor U11265 (N_11265,N_11085,N_11075);
xor U11266 (N_11266,N_11105,N_11061);
and U11267 (N_11267,N_11178,N_11165);
or U11268 (N_11268,N_11095,N_11092);
and U11269 (N_11269,N_11048,N_11118);
xnor U11270 (N_11270,N_11162,N_11094);
or U11271 (N_11271,N_11113,N_11142);
xnor U11272 (N_11272,N_11139,N_11169);
and U11273 (N_11273,N_11134,N_11074);
nor U11274 (N_11274,N_11018,N_11177);
nor U11275 (N_11275,N_11077,N_11104);
nor U11276 (N_11276,N_11112,N_11103);
nor U11277 (N_11277,N_11031,N_11110);
xor U11278 (N_11278,N_11070,N_11137);
xor U11279 (N_11279,N_11126,N_11160);
or U11280 (N_11280,N_11023,N_11072);
nor U11281 (N_11281,N_11032,N_11098);
nor U11282 (N_11282,N_11179,N_11082);
and U11283 (N_11283,N_11019,N_11057);
or U11284 (N_11284,N_11062,N_11170);
and U11285 (N_11285,N_11017,N_11053);
and U11286 (N_11286,N_11063,N_11120);
xnor U11287 (N_11287,N_11076,N_11128);
xor U11288 (N_11288,N_11001,N_11129);
nand U11289 (N_11289,N_11127,N_11093);
and U11290 (N_11290,N_11013,N_11130);
or U11291 (N_11291,N_11185,N_11065);
nand U11292 (N_11292,N_11167,N_11002);
xor U11293 (N_11293,N_11148,N_11073);
xor U11294 (N_11294,N_11157,N_11068);
and U11295 (N_11295,N_11187,N_11146);
or U11296 (N_11296,N_11088,N_11108);
xor U11297 (N_11297,N_11015,N_11055);
nand U11298 (N_11298,N_11045,N_11114);
nor U11299 (N_11299,N_11089,N_11040);
xnor U11300 (N_11300,N_11102,N_11013);
xnor U11301 (N_11301,N_11130,N_11011);
nor U11302 (N_11302,N_11199,N_11188);
and U11303 (N_11303,N_11053,N_11087);
and U11304 (N_11304,N_11155,N_11034);
and U11305 (N_11305,N_11043,N_11161);
or U11306 (N_11306,N_11083,N_11047);
nor U11307 (N_11307,N_11097,N_11046);
nor U11308 (N_11308,N_11174,N_11001);
nand U11309 (N_11309,N_11102,N_11195);
xor U11310 (N_11310,N_11119,N_11134);
or U11311 (N_11311,N_11079,N_11126);
and U11312 (N_11312,N_11138,N_11031);
or U11313 (N_11313,N_11194,N_11170);
and U11314 (N_11314,N_11059,N_11151);
nor U11315 (N_11315,N_11129,N_11060);
nor U11316 (N_11316,N_11035,N_11106);
nor U11317 (N_11317,N_11048,N_11000);
or U11318 (N_11318,N_11015,N_11162);
xor U11319 (N_11319,N_11009,N_11140);
nor U11320 (N_11320,N_11011,N_11118);
xnor U11321 (N_11321,N_11061,N_11025);
and U11322 (N_11322,N_11163,N_11021);
xnor U11323 (N_11323,N_11066,N_11021);
or U11324 (N_11324,N_11051,N_11031);
or U11325 (N_11325,N_11122,N_11079);
nor U11326 (N_11326,N_11122,N_11194);
xnor U11327 (N_11327,N_11164,N_11135);
or U11328 (N_11328,N_11059,N_11043);
or U11329 (N_11329,N_11147,N_11053);
nand U11330 (N_11330,N_11081,N_11043);
nand U11331 (N_11331,N_11152,N_11061);
nand U11332 (N_11332,N_11112,N_11116);
nor U11333 (N_11333,N_11055,N_11000);
nor U11334 (N_11334,N_11178,N_11181);
xor U11335 (N_11335,N_11029,N_11141);
nor U11336 (N_11336,N_11187,N_11138);
nor U11337 (N_11337,N_11021,N_11078);
or U11338 (N_11338,N_11041,N_11021);
nor U11339 (N_11339,N_11080,N_11018);
nand U11340 (N_11340,N_11037,N_11102);
and U11341 (N_11341,N_11078,N_11107);
or U11342 (N_11342,N_11141,N_11099);
or U11343 (N_11343,N_11068,N_11189);
nor U11344 (N_11344,N_11029,N_11113);
nor U11345 (N_11345,N_11057,N_11100);
nor U11346 (N_11346,N_11034,N_11192);
and U11347 (N_11347,N_11059,N_11082);
and U11348 (N_11348,N_11166,N_11085);
xnor U11349 (N_11349,N_11088,N_11105);
xnor U11350 (N_11350,N_11120,N_11045);
nand U11351 (N_11351,N_11109,N_11123);
or U11352 (N_11352,N_11065,N_11123);
xor U11353 (N_11353,N_11124,N_11067);
xor U11354 (N_11354,N_11088,N_11073);
nand U11355 (N_11355,N_11152,N_11133);
and U11356 (N_11356,N_11171,N_11108);
and U11357 (N_11357,N_11122,N_11042);
nor U11358 (N_11358,N_11185,N_11151);
nand U11359 (N_11359,N_11168,N_11009);
and U11360 (N_11360,N_11147,N_11185);
nand U11361 (N_11361,N_11185,N_11141);
nand U11362 (N_11362,N_11015,N_11052);
xnor U11363 (N_11363,N_11030,N_11080);
nor U11364 (N_11364,N_11173,N_11020);
nor U11365 (N_11365,N_11075,N_11072);
and U11366 (N_11366,N_11003,N_11004);
nand U11367 (N_11367,N_11143,N_11088);
and U11368 (N_11368,N_11118,N_11181);
or U11369 (N_11369,N_11038,N_11020);
nor U11370 (N_11370,N_11085,N_11195);
nor U11371 (N_11371,N_11190,N_11063);
or U11372 (N_11372,N_11039,N_11038);
and U11373 (N_11373,N_11034,N_11158);
xor U11374 (N_11374,N_11035,N_11181);
nor U11375 (N_11375,N_11049,N_11185);
xor U11376 (N_11376,N_11066,N_11194);
xnor U11377 (N_11377,N_11198,N_11016);
or U11378 (N_11378,N_11168,N_11043);
and U11379 (N_11379,N_11066,N_11086);
nor U11380 (N_11380,N_11017,N_11040);
nand U11381 (N_11381,N_11073,N_11124);
and U11382 (N_11382,N_11165,N_11086);
xnor U11383 (N_11383,N_11081,N_11134);
and U11384 (N_11384,N_11065,N_11134);
nand U11385 (N_11385,N_11126,N_11102);
xnor U11386 (N_11386,N_11079,N_11067);
xor U11387 (N_11387,N_11136,N_11099);
or U11388 (N_11388,N_11157,N_11037);
nor U11389 (N_11389,N_11090,N_11102);
nor U11390 (N_11390,N_11081,N_11002);
xor U11391 (N_11391,N_11092,N_11034);
xor U11392 (N_11392,N_11014,N_11156);
xor U11393 (N_11393,N_11176,N_11037);
or U11394 (N_11394,N_11026,N_11061);
and U11395 (N_11395,N_11072,N_11046);
xnor U11396 (N_11396,N_11044,N_11070);
nand U11397 (N_11397,N_11179,N_11188);
and U11398 (N_11398,N_11094,N_11157);
nor U11399 (N_11399,N_11024,N_11198);
or U11400 (N_11400,N_11302,N_11290);
or U11401 (N_11401,N_11255,N_11241);
nand U11402 (N_11402,N_11279,N_11217);
nor U11403 (N_11403,N_11354,N_11372);
and U11404 (N_11404,N_11394,N_11208);
xor U11405 (N_11405,N_11390,N_11306);
nor U11406 (N_11406,N_11223,N_11203);
and U11407 (N_11407,N_11305,N_11285);
xor U11408 (N_11408,N_11325,N_11288);
nand U11409 (N_11409,N_11393,N_11281);
and U11410 (N_11410,N_11384,N_11259);
nand U11411 (N_11411,N_11368,N_11339);
xnor U11412 (N_11412,N_11278,N_11249);
nand U11413 (N_11413,N_11301,N_11369);
or U11414 (N_11414,N_11320,N_11231);
nand U11415 (N_11415,N_11352,N_11373);
nand U11416 (N_11416,N_11219,N_11221);
or U11417 (N_11417,N_11271,N_11361);
nor U11418 (N_11418,N_11389,N_11298);
nor U11419 (N_11419,N_11370,N_11353);
nor U11420 (N_11420,N_11265,N_11381);
and U11421 (N_11421,N_11233,N_11287);
nand U11422 (N_11422,N_11210,N_11299);
and U11423 (N_11423,N_11258,N_11309);
or U11424 (N_11424,N_11211,N_11310);
and U11425 (N_11425,N_11216,N_11378);
or U11426 (N_11426,N_11234,N_11206);
and U11427 (N_11427,N_11350,N_11292);
nand U11428 (N_11428,N_11311,N_11282);
and U11429 (N_11429,N_11204,N_11209);
and U11430 (N_11430,N_11360,N_11345);
and U11431 (N_11431,N_11340,N_11229);
or U11432 (N_11432,N_11395,N_11242);
nor U11433 (N_11433,N_11263,N_11230);
nand U11434 (N_11434,N_11245,N_11387);
nand U11435 (N_11435,N_11379,N_11296);
nand U11436 (N_11436,N_11335,N_11371);
nand U11437 (N_11437,N_11222,N_11256);
or U11438 (N_11438,N_11382,N_11396);
nand U11439 (N_11439,N_11253,N_11254);
nor U11440 (N_11440,N_11348,N_11383);
or U11441 (N_11441,N_11270,N_11272);
and U11442 (N_11442,N_11261,N_11375);
nor U11443 (N_11443,N_11347,N_11262);
nor U11444 (N_11444,N_11313,N_11248);
xnor U11445 (N_11445,N_11334,N_11266);
and U11446 (N_11446,N_11228,N_11257);
or U11447 (N_11447,N_11332,N_11338);
xor U11448 (N_11448,N_11386,N_11236);
nor U11449 (N_11449,N_11226,N_11201);
or U11450 (N_11450,N_11391,N_11247);
nor U11451 (N_11451,N_11363,N_11326);
nor U11452 (N_11452,N_11377,N_11239);
and U11453 (N_11453,N_11362,N_11304);
nand U11454 (N_11454,N_11235,N_11202);
and U11455 (N_11455,N_11398,N_11349);
nor U11456 (N_11456,N_11355,N_11225);
nand U11457 (N_11457,N_11359,N_11397);
xor U11458 (N_11458,N_11273,N_11275);
xor U11459 (N_11459,N_11341,N_11358);
nor U11460 (N_11460,N_11246,N_11321);
nor U11461 (N_11461,N_11342,N_11289);
nand U11462 (N_11462,N_11252,N_11330);
nor U11463 (N_11463,N_11323,N_11251);
and U11464 (N_11464,N_11200,N_11220);
xnor U11465 (N_11465,N_11205,N_11250);
nand U11466 (N_11466,N_11260,N_11264);
xor U11467 (N_11467,N_11344,N_11357);
and U11468 (N_11468,N_11244,N_11367);
nor U11469 (N_11469,N_11308,N_11276);
and U11470 (N_11470,N_11237,N_11294);
xor U11471 (N_11471,N_11295,N_11215);
nor U11472 (N_11472,N_11322,N_11224);
nor U11473 (N_11473,N_11392,N_11327);
nor U11474 (N_11474,N_11399,N_11286);
nor U11475 (N_11475,N_11374,N_11337);
and U11476 (N_11476,N_11351,N_11284);
xor U11477 (N_11477,N_11293,N_11212);
nor U11478 (N_11478,N_11274,N_11328);
and U11479 (N_11479,N_11319,N_11227);
nand U11480 (N_11480,N_11297,N_11218);
or U11481 (N_11481,N_11207,N_11376);
nor U11482 (N_11482,N_11214,N_11346);
and U11483 (N_11483,N_11317,N_11315);
nor U11484 (N_11484,N_11336,N_11312);
nand U11485 (N_11485,N_11316,N_11329);
nor U11486 (N_11486,N_11243,N_11356);
and U11487 (N_11487,N_11307,N_11303);
or U11488 (N_11488,N_11267,N_11213);
nand U11489 (N_11489,N_11331,N_11232);
or U11490 (N_11490,N_11343,N_11333);
and U11491 (N_11491,N_11324,N_11300);
nand U11492 (N_11492,N_11291,N_11364);
xor U11493 (N_11493,N_11380,N_11318);
nand U11494 (N_11494,N_11238,N_11240);
and U11495 (N_11495,N_11277,N_11283);
xnor U11496 (N_11496,N_11268,N_11280);
nand U11497 (N_11497,N_11314,N_11269);
or U11498 (N_11498,N_11388,N_11385);
and U11499 (N_11499,N_11366,N_11365);
and U11500 (N_11500,N_11332,N_11363);
nand U11501 (N_11501,N_11342,N_11232);
nor U11502 (N_11502,N_11290,N_11331);
or U11503 (N_11503,N_11279,N_11364);
and U11504 (N_11504,N_11208,N_11337);
nand U11505 (N_11505,N_11280,N_11388);
or U11506 (N_11506,N_11394,N_11279);
nor U11507 (N_11507,N_11391,N_11220);
nor U11508 (N_11508,N_11353,N_11244);
xnor U11509 (N_11509,N_11248,N_11286);
nor U11510 (N_11510,N_11380,N_11274);
or U11511 (N_11511,N_11264,N_11214);
nand U11512 (N_11512,N_11215,N_11263);
and U11513 (N_11513,N_11274,N_11325);
and U11514 (N_11514,N_11378,N_11211);
nand U11515 (N_11515,N_11224,N_11335);
and U11516 (N_11516,N_11275,N_11292);
xnor U11517 (N_11517,N_11334,N_11240);
xnor U11518 (N_11518,N_11356,N_11383);
or U11519 (N_11519,N_11232,N_11353);
xor U11520 (N_11520,N_11271,N_11227);
and U11521 (N_11521,N_11328,N_11309);
and U11522 (N_11522,N_11225,N_11214);
xnor U11523 (N_11523,N_11255,N_11231);
nor U11524 (N_11524,N_11381,N_11310);
and U11525 (N_11525,N_11290,N_11208);
and U11526 (N_11526,N_11392,N_11330);
and U11527 (N_11527,N_11387,N_11203);
nor U11528 (N_11528,N_11219,N_11291);
and U11529 (N_11529,N_11311,N_11241);
and U11530 (N_11530,N_11276,N_11299);
nor U11531 (N_11531,N_11368,N_11382);
nor U11532 (N_11532,N_11281,N_11267);
xnor U11533 (N_11533,N_11275,N_11379);
xnor U11534 (N_11534,N_11331,N_11378);
xnor U11535 (N_11535,N_11344,N_11215);
and U11536 (N_11536,N_11281,N_11248);
and U11537 (N_11537,N_11267,N_11233);
nand U11538 (N_11538,N_11291,N_11259);
xnor U11539 (N_11539,N_11276,N_11342);
nand U11540 (N_11540,N_11249,N_11308);
nand U11541 (N_11541,N_11262,N_11281);
nand U11542 (N_11542,N_11251,N_11270);
or U11543 (N_11543,N_11229,N_11222);
or U11544 (N_11544,N_11397,N_11288);
nor U11545 (N_11545,N_11224,N_11353);
or U11546 (N_11546,N_11365,N_11208);
and U11547 (N_11547,N_11213,N_11288);
and U11548 (N_11548,N_11291,N_11388);
or U11549 (N_11549,N_11379,N_11249);
nor U11550 (N_11550,N_11284,N_11340);
or U11551 (N_11551,N_11312,N_11276);
nand U11552 (N_11552,N_11234,N_11366);
xnor U11553 (N_11553,N_11287,N_11235);
or U11554 (N_11554,N_11294,N_11396);
xnor U11555 (N_11555,N_11383,N_11254);
nor U11556 (N_11556,N_11302,N_11371);
or U11557 (N_11557,N_11255,N_11324);
nand U11558 (N_11558,N_11341,N_11394);
nor U11559 (N_11559,N_11254,N_11362);
nand U11560 (N_11560,N_11327,N_11366);
nand U11561 (N_11561,N_11224,N_11217);
nand U11562 (N_11562,N_11388,N_11203);
xnor U11563 (N_11563,N_11384,N_11249);
and U11564 (N_11564,N_11360,N_11273);
nand U11565 (N_11565,N_11305,N_11395);
nand U11566 (N_11566,N_11302,N_11244);
xor U11567 (N_11567,N_11253,N_11264);
or U11568 (N_11568,N_11316,N_11232);
nand U11569 (N_11569,N_11231,N_11343);
or U11570 (N_11570,N_11284,N_11342);
and U11571 (N_11571,N_11234,N_11322);
nor U11572 (N_11572,N_11259,N_11316);
xnor U11573 (N_11573,N_11229,N_11371);
xor U11574 (N_11574,N_11399,N_11264);
or U11575 (N_11575,N_11209,N_11315);
and U11576 (N_11576,N_11207,N_11277);
nor U11577 (N_11577,N_11246,N_11302);
or U11578 (N_11578,N_11363,N_11287);
or U11579 (N_11579,N_11372,N_11222);
xor U11580 (N_11580,N_11223,N_11378);
nor U11581 (N_11581,N_11263,N_11245);
or U11582 (N_11582,N_11281,N_11332);
nor U11583 (N_11583,N_11340,N_11302);
xnor U11584 (N_11584,N_11345,N_11317);
and U11585 (N_11585,N_11260,N_11365);
nand U11586 (N_11586,N_11279,N_11322);
or U11587 (N_11587,N_11334,N_11282);
or U11588 (N_11588,N_11262,N_11399);
nor U11589 (N_11589,N_11342,N_11328);
nand U11590 (N_11590,N_11216,N_11386);
nor U11591 (N_11591,N_11362,N_11205);
xor U11592 (N_11592,N_11274,N_11364);
xnor U11593 (N_11593,N_11276,N_11302);
and U11594 (N_11594,N_11207,N_11249);
or U11595 (N_11595,N_11297,N_11315);
or U11596 (N_11596,N_11245,N_11312);
and U11597 (N_11597,N_11222,N_11254);
and U11598 (N_11598,N_11219,N_11320);
nor U11599 (N_11599,N_11351,N_11207);
nand U11600 (N_11600,N_11585,N_11512);
nand U11601 (N_11601,N_11471,N_11488);
nor U11602 (N_11602,N_11451,N_11558);
and U11603 (N_11603,N_11570,N_11591);
nor U11604 (N_11604,N_11485,N_11427);
and U11605 (N_11605,N_11475,N_11448);
or U11606 (N_11606,N_11514,N_11523);
and U11607 (N_11607,N_11455,N_11513);
nor U11608 (N_11608,N_11564,N_11435);
and U11609 (N_11609,N_11550,N_11571);
or U11610 (N_11610,N_11548,N_11426);
xnor U11611 (N_11611,N_11461,N_11587);
nand U11612 (N_11612,N_11495,N_11486);
xnor U11613 (N_11613,N_11439,N_11510);
and U11614 (N_11614,N_11480,N_11506);
or U11615 (N_11615,N_11560,N_11420);
and U11616 (N_11616,N_11563,N_11578);
and U11617 (N_11617,N_11476,N_11458);
nand U11618 (N_11618,N_11419,N_11519);
nand U11619 (N_11619,N_11532,N_11579);
and U11620 (N_11620,N_11528,N_11531);
and U11621 (N_11621,N_11406,N_11567);
nor U11622 (N_11622,N_11540,N_11421);
nand U11623 (N_11623,N_11598,N_11539);
nand U11624 (N_11624,N_11457,N_11559);
and U11625 (N_11625,N_11518,N_11580);
and U11626 (N_11626,N_11590,N_11584);
nand U11627 (N_11627,N_11418,N_11544);
or U11628 (N_11628,N_11487,N_11556);
nor U11629 (N_11629,N_11589,N_11465);
or U11630 (N_11630,N_11401,N_11469);
nand U11631 (N_11631,N_11482,N_11542);
nor U11632 (N_11632,N_11562,N_11416);
nand U11633 (N_11633,N_11569,N_11505);
xnor U11634 (N_11634,N_11561,N_11454);
or U11635 (N_11635,N_11545,N_11450);
and U11636 (N_11636,N_11509,N_11430);
or U11637 (N_11637,N_11400,N_11446);
nor U11638 (N_11638,N_11463,N_11489);
nand U11639 (N_11639,N_11565,N_11557);
or U11640 (N_11640,N_11520,N_11552);
or U11641 (N_11641,N_11515,N_11445);
or U11642 (N_11642,N_11497,N_11459);
xnor U11643 (N_11643,N_11516,N_11404);
nor U11644 (N_11644,N_11588,N_11534);
xnor U11645 (N_11645,N_11527,N_11555);
nor U11646 (N_11646,N_11408,N_11483);
and U11647 (N_11647,N_11462,N_11425);
or U11648 (N_11648,N_11592,N_11575);
nor U11649 (N_11649,N_11581,N_11549);
xor U11650 (N_11650,N_11440,N_11524);
or U11651 (N_11651,N_11507,N_11444);
nand U11652 (N_11652,N_11496,N_11547);
nor U11653 (N_11653,N_11503,N_11521);
xnor U11654 (N_11654,N_11599,N_11583);
nand U11655 (N_11655,N_11594,N_11405);
xnor U11656 (N_11656,N_11452,N_11597);
nand U11657 (N_11657,N_11478,N_11402);
nor U11658 (N_11658,N_11538,N_11508);
and U11659 (N_11659,N_11428,N_11566);
nand U11660 (N_11660,N_11413,N_11494);
nor U11661 (N_11661,N_11525,N_11554);
nand U11662 (N_11662,N_11474,N_11442);
nor U11663 (N_11663,N_11412,N_11436);
xor U11664 (N_11664,N_11410,N_11537);
nand U11665 (N_11665,N_11526,N_11573);
and U11666 (N_11666,N_11491,N_11511);
nand U11667 (N_11667,N_11504,N_11414);
or U11668 (N_11668,N_11437,N_11477);
nand U11669 (N_11669,N_11453,N_11484);
nand U11670 (N_11670,N_11568,N_11467);
and U11671 (N_11671,N_11431,N_11535);
nand U11672 (N_11672,N_11464,N_11481);
nor U11673 (N_11673,N_11551,N_11577);
and U11674 (N_11674,N_11502,N_11470);
xnor U11675 (N_11675,N_11596,N_11574);
or U11676 (N_11676,N_11582,N_11411);
and U11677 (N_11677,N_11553,N_11403);
nand U11678 (N_11678,N_11586,N_11546);
nor U11679 (N_11679,N_11499,N_11407);
nand U11680 (N_11680,N_11543,N_11493);
and U11681 (N_11681,N_11536,N_11498);
and U11682 (N_11682,N_11429,N_11529);
xor U11683 (N_11683,N_11595,N_11533);
nand U11684 (N_11684,N_11422,N_11441);
xor U11685 (N_11685,N_11572,N_11517);
nor U11686 (N_11686,N_11472,N_11443);
nor U11687 (N_11687,N_11432,N_11423);
and U11688 (N_11688,N_11490,N_11449);
and U11689 (N_11689,N_11473,N_11424);
nor U11690 (N_11690,N_11434,N_11433);
nand U11691 (N_11691,N_11492,N_11417);
and U11692 (N_11692,N_11530,N_11541);
nand U11693 (N_11693,N_11576,N_11593);
nand U11694 (N_11694,N_11466,N_11460);
xor U11695 (N_11695,N_11501,N_11409);
or U11696 (N_11696,N_11415,N_11456);
xnor U11697 (N_11697,N_11438,N_11522);
or U11698 (N_11698,N_11447,N_11500);
or U11699 (N_11699,N_11468,N_11479);
and U11700 (N_11700,N_11543,N_11506);
xor U11701 (N_11701,N_11496,N_11499);
nand U11702 (N_11702,N_11446,N_11521);
nand U11703 (N_11703,N_11444,N_11453);
or U11704 (N_11704,N_11441,N_11503);
nor U11705 (N_11705,N_11525,N_11514);
and U11706 (N_11706,N_11442,N_11405);
nand U11707 (N_11707,N_11493,N_11488);
xor U11708 (N_11708,N_11478,N_11432);
and U11709 (N_11709,N_11494,N_11597);
xor U11710 (N_11710,N_11498,N_11594);
or U11711 (N_11711,N_11533,N_11519);
nand U11712 (N_11712,N_11432,N_11422);
xnor U11713 (N_11713,N_11518,N_11486);
nand U11714 (N_11714,N_11456,N_11424);
nand U11715 (N_11715,N_11453,N_11531);
nor U11716 (N_11716,N_11568,N_11482);
nor U11717 (N_11717,N_11556,N_11532);
or U11718 (N_11718,N_11580,N_11541);
xor U11719 (N_11719,N_11414,N_11493);
nand U11720 (N_11720,N_11582,N_11506);
xnor U11721 (N_11721,N_11530,N_11485);
nor U11722 (N_11722,N_11410,N_11422);
nor U11723 (N_11723,N_11562,N_11498);
nor U11724 (N_11724,N_11485,N_11578);
nor U11725 (N_11725,N_11412,N_11588);
xnor U11726 (N_11726,N_11546,N_11596);
or U11727 (N_11727,N_11542,N_11423);
and U11728 (N_11728,N_11408,N_11400);
and U11729 (N_11729,N_11571,N_11468);
xnor U11730 (N_11730,N_11572,N_11533);
nand U11731 (N_11731,N_11559,N_11460);
or U11732 (N_11732,N_11451,N_11513);
or U11733 (N_11733,N_11491,N_11474);
nor U11734 (N_11734,N_11582,N_11416);
nor U11735 (N_11735,N_11548,N_11409);
xor U11736 (N_11736,N_11550,N_11543);
xnor U11737 (N_11737,N_11561,N_11532);
and U11738 (N_11738,N_11599,N_11562);
nor U11739 (N_11739,N_11527,N_11467);
xor U11740 (N_11740,N_11412,N_11509);
xor U11741 (N_11741,N_11504,N_11512);
or U11742 (N_11742,N_11574,N_11489);
or U11743 (N_11743,N_11428,N_11420);
nand U11744 (N_11744,N_11515,N_11543);
nor U11745 (N_11745,N_11512,N_11568);
xnor U11746 (N_11746,N_11410,N_11419);
nor U11747 (N_11747,N_11404,N_11549);
or U11748 (N_11748,N_11592,N_11507);
nand U11749 (N_11749,N_11596,N_11532);
xor U11750 (N_11750,N_11520,N_11531);
or U11751 (N_11751,N_11472,N_11457);
and U11752 (N_11752,N_11403,N_11523);
or U11753 (N_11753,N_11532,N_11480);
or U11754 (N_11754,N_11433,N_11524);
nand U11755 (N_11755,N_11497,N_11477);
or U11756 (N_11756,N_11484,N_11415);
or U11757 (N_11757,N_11456,N_11560);
or U11758 (N_11758,N_11504,N_11425);
nand U11759 (N_11759,N_11443,N_11517);
xor U11760 (N_11760,N_11425,N_11432);
nand U11761 (N_11761,N_11505,N_11472);
or U11762 (N_11762,N_11404,N_11470);
nand U11763 (N_11763,N_11432,N_11547);
or U11764 (N_11764,N_11412,N_11464);
nor U11765 (N_11765,N_11412,N_11489);
nand U11766 (N_11766,N_11485,N_11458);
nor U11767 (N_11767,N_11506,N_11496);
and U11768 (N_11768,N_11538,N_11575);
xor U11769 (N_11769,N_11524,N_11436);
and U11770 (N_11770,N_11467,N_11515);
and U11771 (N_11771,N_11537,N_11563);
xnor U11772 (N_11772,N_11414,N_11531);
and U11773 (N_11773,N_11432,N_11418);
xnor U11774 (N_11774,N_11511,N_11452);
and U11775 (N_11775,N_11413,N_11561);
or U11776 (N_11776,N_11463,N_11520);
or U11777 (N_11777,N_11413,N_11426);
nor U11778 (N_11778,N_11596,N_11431);
xor U11779 (N_11779,N_11564,N_11524);
nand U11780 (N_11780,N_11510,N_11448);
xor U11781 (N_11781,N_11459,N_11584);
nor U11782 (N_11782,N_11512,N_11518);
xor U11783 (N_11783,N_11564,N_11508);
nand U11784 (N_11784,N_11509,N_11433);
nand U11785 (N_11785,N_11592,N_11504);
or U11786 (N_11786,N_11418,N_11586);
or U11787 (N_11787,N_11451,N_11539);
nand U11788 (N_11788,N_11585,N_11547);
nand U11789 (N_11789,N_11501,N_11496);
xnor U11790 (N_11790,N_11598,N_11504);
and U11791 (N_11791,N_11519,N_11445);
or U11792 (N_11792,N_11592,N_11440);
nand U11793 (N_11793,N_11530,N_11595);
or U11794 (N_11794,N_11465,N_11422);
and U11795 (N_11795,N_11529,N_11414);
nor U11796 (N_11796,N_11493,N_11495);
or U11797 (N_11797,N_11479,N_11524);
nor U11798 (N_11798,N_11539,N_11521);
xor U11799 (N_11799,N_11511,N_11563);
nand U11800 (N_11800,N_11637,N_11735);
xnor U11801 (N_11801,N_11636,N_11686);
or U11802 (N_11802,N_11659,N_11749);
nand U11803 (N_11803,N_11691,N_11611);
nor U11804 (N_11804,N_11662,N_11603);
or U11805 (N_11805,N_11709,N_11633);
or U11806 (N_11806,N_11678,N_11625);
xor U11807 (N_11807,N_11688,N_11604);
xnor U11808 (N_11808,N_11738,N_11660);
or U11809 (N_11809,N_11729,N_11793);
nor U11810 (N_11810,N_11671,N_11797);
nor U11811 (N_11811,N_11742,N_11654);
nor U11812 (N_11812,N_11646,N_11799);
xnor U11813 (N_11813,N_11672,N_11619);
and U11814 (N_11814,N_11798,N_11669);
nor U11815 (N_11815,N_11668,N_11683);
or U11816 (N_11816,N_11763,N_11605);
nor U11817 (N_11817,N_11717,N_11730);
and U11818 (N_11818,N_11631,N_11700);
nand U11819 (N_11819,N_11701,N_11716);
or U11820 (N_11820,N_11706,N_11705);
nand U11821 (N_11821,N_11682,N_11724);
nand U11822 (N_11822,N_11677,N_11769);
nor U11823 (N_11823,N_11609,N_11777);
or U11824 (N_11824,N_11721,N_11634);
xor U11825 (N_11825,N_11759,N_11737);
nand U11826 (N_11826,N_11630,N_11788);
and U11827 (N_11827,N_11756,N_11783);
xor U11828 (N_11828,N_11658,N_11685);
nand U11829 (N_11829,N_11789,N_11612);
or U11830 (N_11830,N_11695,N_11621);
or U11831 (N_11831,N_11618,N_11667);
xnor U11832 (N_11832,N_11649,N_11762);
and U11833 (N_11833,N_11698,N_11702);
nor U11834 (N_11834,N_11725,N_11727);
or U11835 (N_11835,N_11676,N_11656);
nand U11836 (N_11836,N_11773,N_11720);
or U11837 (N_11837,N_11616,N_11746);
and U11838 (N_11838,N_11774,N_11650);
nor U11839 (N_11839,N_11684,N_11606);
nor U11840 (N_11840,N_11750,N_11786);
and U11841 (N_11841,N_11670,N_11647);
and U11842 (N_11842,N_11692,N_11714);
xnor U11843 (N_11843,N_11745,N_11610);
nor U11844 (N_11844,N_11718,N_11719);
and U11845 (N_11845,N_11644,N_11743);
nor U11846 (N_11846,N_11780,N_11600);
or U11847 (N_11847,N_11771,N_11794);
xor U11848 (N_11848,N_11694,N_11744);
xor U11849 (N_11849,N_11664,N_11766);
nor U11850 (N_11850,N_11657,N_11753);
nor U11851 (N_11851,N_11734,N_11768);
and U11852 (N_11852,N_11687,N_11728);
nor U11853 (N_11853,N_11617,N_11639);
or U11854 (N_11854,N_11641,N_11772);
xor U11855 (N_11855,N_11602,N_11758);
or U11856 (N_11856,N_11632,N_11748);
nand U11857 (N_11857,N_11733,N_11697);
or U11858 (N_11858,N_11615,N_11628);
xor U11859 (N_11859,N_11674,N_11689);
nor U11860 (N_11860,N_11693,N_11652);
or U11861 (N_11861,N_11732,N_11601);
xor U11862 (N_11862,N_11764,N_11747);
and U11863 (N_11863,N_11627,N_11715);
xor U11864 (N_11864,N_11623,N_11741);
xnor U11865 (N_11865,N_11648,N_11779);
nand U11866 (N_11866,N_11736,N_11711);
nor U11867 (N_11867,N_11760,N_11626);
or U11868 (N_11868,N_11761,N_11699);
nand U11869 (N_11869,N_11731,N_11638);
nand U11870 (N_11870,N_11651,N_11781);
nand U11871 (N_11871,N_11673,N_11643);
xnor U11872 (N_11872,N_11782,N_11613);
and U11873 (N_11873,N_11755,N_11787);
xor U11874 (N_11874,N_11792,N_11754);
or U11875 (N_11875,N_11795,N_11752);
and U11876 (N_11876,N_11740,N_11723);
nand U11877 (N_11877,N_11712,N_11640);
and U11878 (N_11878,N_11726,N_11655);
nand U11879 (N_11879,N_11713,N_11665);
xnor U11880 (N_11880,N_11790,N_11653);
or U11881 (N_11881,N_11703,N_11681);
nor U11882 (N_11882,N_11607,N_11767);
and U11883 (N_11883,N_11622,N_11791);
or U11884 (N_11884,N_11679,N_11775);
nor U11885 (N_11885,N_11629,N_11635);
nor U11886 (N_11886,N_11680,N_11784);
xnor U11887 (N_11887,N_11710,N_11757);
xnor U11888 (N_11888,N_11624,N_11675);
xor U11889 (N_11889,N_11696,N_11770);
nor U11890 (N_11890,N_11608,N_11707);
nand U11891 (N_11891,N_11722,N_11796);
nor U11892 (N_11892,N_11661,N_11776);
nand U11893 (N_11893,N_11614,N_11765);
xor U11894 (N_11894,N_11620,N_11663);
nor U11895 (N_11895,N_11645,N_11690);
or U11896 (N_11896,N_11708,N_11642);
nor U11897 (N_11897,N_11751,N_11666);
or U11898 (N_11898,N_11778,N_11704);
or U11899 (N_11899,N_11739,N_11785);
xnor U11900 (N_11900,N_11632,N_11653);
xnor U11901 (N_11901,N_11650,N_11613);
and U11902 (N_11902,N_11612,N_11615);
nand U11903 (N_11903,N_11781,N_11732);
nor U11904 (N_11904,N_11743,N_11782);
nor U11905 (N_11905,N_11691,N_11724);
xor U11906 (N_11906,N_11670,N_11677);
nor U11907 (N_11907,N_11762,N_11606);
and U11908 (N_11908,N_11686,N_11726);
xor U11909 (N_11909,N_11607,N_11666);
nor U11910 (N_11910,N_11674,N_11623);
nor U11911 (N_11911,N_11762,N_11641);
xnor U11912 (N_11912,N_11776,N_11665);
xnor U11913 (N_11913,N_11607,N_11749);
or U11914 (N_11914,N_11624,N_11740);
and U11915 (N_11915,N_11765,N_11684);
nor U11916 (N_11916,N_11797,N_11751);
nor U11917 (N_11917,N_11651,N_11718);
and U11918 (N_11918,N_11675,N_11756);
nand U11919 (N_11919,N_11728,N_11766);
and U11920 (N_11920,N_11765,N_11772);
and U11921 (N_11921,N_11738,N_11761);
nand U11922 (N_11922,N_11669,N_11794);
nand U11923 (N_11923,N_11761,N_11726);
or U11924 (N_11924,N_11667,N_11784);
xnor U11925 (N_11925,N_11617,N_11603);
or U11926 (N_11926,N_11621,N_11741);
or U11927 (N_11927,N_11704,N_11787);
nand U11928 (N_11928,N_11656,N_11609);
or U11929 (N_11929,N_11746,N_11605);
xor U11930 (N_11930,N_11737,N_11651);
nand U11931 (N_11931,N_11628,N_11790);
and U11932 (N_11932,N_11605,N_11601);
xnor U11933 (N_11933,N_11780,N_11756);
or U11934 (N_11934,N_11700,N_11741);
xor U11935 (N_11935,N_11685,N_11728);
nand U11936 (N_11936,N_11713,N_11670);
nand U11937 (N_11937,N_11758,N_11637);
nand U11938 (N_11938,N_11790,N_11662);
nand U11939 (N_11939,N_11651,N_11771);
and U11940 (N_11940,N_11784,N_11692);
nor U11941 (N_11941,N_11786,N_11698);
and U11942 (N_11942,N_11616,N_11614);
and U11943 (N_11943,N_11784,N_11709);
nor U11944 (N_11944,N_11642,N_11696);
nand U11945 (N_11945,N_11701,N_11621);
and U11946 (N_11946,N_11634,N_11779);
or U11947 (N_11947,N_11680,N_11756);
nand U11948 (N_11948,N_11753,N_11690);
xor U11949 (N_11949,N_11796,N_11766);
nand U11950 (N_11950,N_11613,N_11616);
nand U11951 (N_11951,N_11669,N_11628);
nor U11952 (N_11952,N_11602,N_11626);
or U11953 (N_11953,N_11737,N_11639);
nand U11954 (N_11954,N_11762,N_11605);
xnor U11955 (N_11955,N_11744,N_11633);
nor U11956 (N_11956,N_11679,N_11690);
or U11957 (N_11957,N_11707,N_11763);
or U11958 (N_11958,N_11607,N_11678);
nor U11959 (N_11959,N_11608,N_11777);
nand U11960 (N_11960,N_11766,N_11732);
and U11961 (N_11961,N_11646,N_11755);
nand U11962 (N_11962,N_11747,N_11787);
or U11963 (N_11963,N_11768,N_11733);
nor U11964 (N_11964,N_11700,N_11616);
nand U11965 (N_11965,N_11611,N_11757);
and U11966 (N_11966,N_11670,N_11706);
xor U11967 (N_11967,N_11632,N_11750);
or U11968 (N_11968,N_11736,N_11783);
xor U11969 (N_11969,N_11792,N_11727);
xnor U11970 (N_11970,N_11767,N_11636);
nand U11971 (N_11971,N_11632,N_11723);
nor U11972 (N_11972,N_11735,N_11606);
nor U11973 (N_11973,N_11629,N_11698);
or U11974 (N_11974,N_11691,N_11688);
nand U11975 (N_11975,N_11660,N_11680);
xnor U11976 (N_11976,N_11666,N_11645);
xor U11977 (N_11977,N_11606,N_11748);
or U11978 (N_11978,N_11687,N_11718);
nor U11979 (N_11979,N_11655,N_11648);
xor U11980 (N_11980,N_11759,N_11632);
nor U11981 (N_11981,N_11655,N_11795);
xnor U11982 (N_11982,N_11767,N_11786);
or U11983 (N_11983,N_11675,N_11631);
nand U11984 (N_11984,N_11761,N_11713);
nand U11985 (N_11985,N_11606,N_11694);
xor U11986 (N_11986,N_11603,N_11654);
nor U11987 (N_11987,N_11747,N_11794);
xor U11988 (N_11988,N_11698,N_11647);
nor U11989 (N_11989,N_11694,N_11723);
nor U11990 (N_11990,N_11791,N_11682);
nor U11991 (N_11991,N_11745,N_11706);
or U11992 (N_11992,N_11794,N_11654);
nand U11993 (N_11993,N_11630,N_11610);
nor U11994 (N_11994,N_11712,N_11611);
or U11995 (N_11995,N_11774,N_11655);
xor U11996 (N_11996,N_11638,N_11755);
nor U11997 (N_11997,N_11639,N_11768);
and U11998 (N_11998,N_11691,N_11782);
or U11999 (N_11999,N_11644,N_11754);
nand U12000 (N_12000,N_11912,N_11815);
nor U12001 (N_12001,N_11972,N_11897);
nor U12002 (N_12002,N_11914,N_11866);
xor U12003 (N_12003,N_11863,N_11818);
nand U12004 (N_12004,N_11885,N_11852);
nand U12005 (N_12005,N_11814,N_11958);
nor U12006 (N_12006,N_11881,N_11903);
nand U12007 (N_12007,N_11981,N_11869);
and U12008 (N_12008,N_11947,N_11865);
and U12009 (N_12009,N_11828,N_11944);
nor U12010 (N_12010,N_11998,N_11884);
nor U12011 (N_12011,N_11970,N_11997);
nor U12012 (N_12012,N_11831,N_11960);
nand U12013 (N_12013,N_11816,N_11977);
nor U12014 (N_12014,N_11837,N_11900);
nand U12015 (N_12015,N_11849,N_11949);
xor U12016 (N_12016,N_11982,N_11834);
nor U12017 (N_12017,N_11820,N_11800);
xnor U12018 (N_12018,N_11833,N_11938);
nor U12019 (N_12019,N_11882,N_11811);
nor U12020 (N_12020,N_11813,N_11995);
nor U12021 (N_12021,N_11999,N_11971);
nand U12022 (N_12022,N_11943,N_11907);
nor U12023 (N_12023,N_11855,N_11948);
and U12024 (N_12024,N_11939,N_11892);
nor U12025 (N_12025,N_11827,N_11821);
and U12026 (N_12026,N_11965,N_11803);
and U12027 (N_12027,N_11874,N_11929);
nor U12028 (N_12028,N_11942,N_11986);
or U12029 (N_12029,N_11919,N_11893);
nand U12030 (N_12030,N_11807,N_11975);
nor U12031 (N_12031,N_11952,N_11926);
xnor U12032 (N_12032,N_11812,N_11924);
or U12033 (N_12033,N_11851,N_11842);
nand U12034 (N_12034,N_11940,N_11941);
nand U12035 (N_12035,N_11802,N_11930);
nand U12036 (N_12036,N_11902,N_11911);
xnor U12037 (N_12037,N_11898,N_11936);
xor U12038 (N_12038,N_11966,N_11878);
xnor U12039 (N_12039,N_11886,N_11961);
or U12040 (N_12040,N_11857,N_11826);
and U12041 (N_12041,N_11973,N_11910);
or U12042 (N_12042,N_11809,N_11860);
nand U12043 (N_12043,N_11850,N_11959);
nor U12044 (N_12044,N_11808,N_11937);
and U12045 (N_12045,N_11935,N_11921);
and U12046 (N_12046,N_11984,N_11861);
and U12047 (N_12047,N_11953,N_11905);
nand U12048 (N_12048,N_11950,N_11899);
xnor U12049 (N_12049,N_11810,N_11932);
nand U12050 (N_12050,N_11859,N_11916);
or U12051 (N_12051,N_11870,N_11896);
nand U12052 (N_12052,N_11945,N_11844);
or U12053 (N_12053,N_11979,N_11962);
xor U12054 (N_12054,N_11846,N_11832);
nand U12055 (N_12055,N_11987,N_11909);
or U12056 (N_12056,N_11817,N_11906);
and U12057 (N_12057,N_11880,N_11858);
xnor U12058 (N_12058,N_11963,N_11923);
and U12059 (N_12059,N_11891,N_11951);
nor U12060 (N_12060,N_11967,N_11883);
and U12061 (N_12061,N_11908,N_11848);
or U12062 (N_12062,N_11877,N_11913);
and U12063 (N_12063,N_11875,N_11829);
nand U12064 (N_12064,N_11835,N_11801);
and U12065 (N_12065,N_11990,N_11978);
nand U12066 (N_12066,N_11934,N_11838);
xor U12067 (N_12067,N_11954,N_11804);
nor U12068 (N_12068,N_11927,N_11819);
and U12069 (N_12069,N_11805,N_11806);
and U12070 (N_12070,N_11876,N_11969);
xnor U12071 (N_12071,N_11964,N_11991);
or U12072 (N_12072,N_11904,N_11894);
nor U12073 (N_12073,N_11974,N_11901);
nand U12074 (N_12074,N_11889,N_11841);
or U12075 (N_12075,N_11996,N_11955);
xnor U12076 (N_12076,N_11993,N_11956);
nor U12077 (N_12077,N_11957,N_11946);
or U12078 (N_12078,N_11853,N_11895);
and U12079 (N_12079,N_11825,N_11856);
and U12080 (N_12080,N_11976,N_11928);
nor U12081 (N_12081,N_11918,N_11871);
nor U12082 (N_12082,N_11879,N_11985);
and U12083 (N_12083,N_11988,N_11920);
or U12084 (N_12084,N_11847,N_11862);
nand U12085 (N_12085,N_11824,N_11839);
xor U12086 (N_12086,N_11868,N_11922);
xnor U12087 (N_12087,N_11836,N_11933);
nand U12088 (N_12088,N_11887,N_11925);
nor U12089 (N_12089,N_11822,N_11917);
or U12090 (N_12090,N_11864,N_11890);
and U12091 (N_12091,N_11830,N_11968);
xor U12092 (N_12092,N_11980,N_11989);
or U12093 (N_12093,N_11854,N_11915);
or U12094 (N_12094,N_11931,N_11888);
nand U12095 (N_12095,N_11994,N_11843);
nand U12096 (N_12096,N_11992,N_11845);
or U12097 (N_12097,N_11983,N_11873);
or U12098 (N_12098,N_11867,N_11872);
nand U12099 (N_12099,N_11840,N_11823);
and U12100 (N_12100,N_11953,N_11893);
and U12101 (N_12101,N_11913,N_11942);
and U12102 (N_12102,N_11877,N_11970);
nor U12103 (N_12103,N_11911,N_11943);
nand U12104 (N_12104,N_11814,N_11959);
or U12105 (N_12105,N_11872,N_11986);
and U12106 (N_12106,N_11921,N_11993);
xnor U12107 (N_12107,N_11859,N_11971);
nand U12108 (N_12108,N_11947,N_11965);
nand U12109 (N_12109,N_11813,N_11984);
and U12110 (N_12110,N_11892,N_11913);
or U12111 (N_12111,N_11820,N_11912);
xnor U12112 (N_12112,N_11998,N_11873);
nor U12113 (N_12113,N_11954,N_11999);
nor U12114 (N_12114,N_11968,N_11853);
and U12115 (N_12115,N_11987,N_11966);
xnor U12116 (N_12116,N_11865,N_11827);
and U12117 (N_12117,N_11952,N_11826);
and U12118 (N_12118,N_11983,N_11948);
xnor U12119 (N_12119,N_11801,N_11920);
nand U12120 (N_12120,N_11849,N_11825);
and U12121 (N_12121,N_11923,N_11984);
or U12122 (N_12122,N_11813,N_11824);
and U12123 (N_12123,N_11851,N_11839);
xor U12124 (N_12124,N_11877,N_11952);
xnor U12125 (N_12125,N_11914,N_11810);
xor U12126 (N_12126,N_11820,N_11846);
nand U12127 (N_12127,N_11901,N_11813);
and U12128 (N_12128,N_11864,N_11980);
nor U12129 (N_12129,N_11921,N_11896);
nand U12130 (N_12130,N_11930,N_11967);
xnor U12131 (N_12131,N_11880,N_11938);
nand U12132 (N_12132,N_11982,N_11806);
and U12133 (N_12133,N_11823,N_11907);
nand U12134 (N_12134,N_11831,N_11968);
xnor U12135 (N_12135,N_11859,N_11909);
or U12136 (N_12136,N_11981,N_11838);
nand U12137 (N_12137,N_11945,N_11982);
and U12138 (N_12138,N_11979,N_11978);
nor U12139 (N_12139,N_11899,N_11928);
or U12140 (N_12140,N_11825,N_11852);
or U12141 (N_12141,N_11884,N_11815);
or U12142 (N_12142,N_11891,N_11976);
nor U12143 (N_12143,N_11868,N_11992);
nand U12144 (N_12144,N_11886,N_11945);
nor U12145 (N_12145,N_11842,N_11979);
nor U12146 (N_12146,N_11910,N_11895);
nor U12147 (N_12147,N_11875,N_11844);
xnor U12148 (N_12148,N_11929,N_11919);
or U12149 (N_12149,N_11845,N_11857);
nor U12150 (N_12150,N_11991,N_11901);
and U12151 (N_12151,N_11873,N_11974);
nand U12152 (N_12152,N_11992,N_11805);
xnor U12153 (N_12153,N_11856,N_11839);
or U12154 (N_12154,N_11858,N_11825);
nor U12155 (N_12155,N_11994,N_11882);
nor U12156 (N_12156,N_11874,N_11853);
nor U12157 (N_12157,N_11876,N_11973);
nor U12158 (N_12158,N_11876,N_11964);
or U12159 (N_12159,N_11998,N_11951);
and U12160 (N_12160,N_11876,N_11932);
nor U12161 (N_12161,N_11921,N_11832);
and U12162 (N_12162,N_11839,N_11869);
nand U12163 (N_12163,N_11852,N_11890);
nor U12164 (N_12164,N_11923,N_11970);
nand U12165 (N_12165,N_11847,N_11914);
or U12166 (N_12166,N_11969,N_11978);
and U12167 (N_12167,N_11932,N_11849);
xor U12168 (N_12168,N_11923,N_11830);
xor U12169 (N_12169,N_11944,N_11820);
nand U12170 (N_12170,N_11803,N_11863);
and U12171 (N_12171,N_11877,N_11896);
nand U12172 (N_12172,N_11862,N_11951);
xnor U12173 (N_12173,N_11932,N_11905);
nor U12174 (N_12174,N_11869,N_11966);
and U12175 (N_12175,N_11987,N_11846);
xor U12176 (N_12176,N_11831,N_11867);
nand U12177 (N_12177,N_11948,N_11854);
nor U12178 (N_12178,N_11802,N_11977);
or U12179 (N_12179,N_11939,N_11968);
nor U12180 (N_12180,N_11934,N_11835);
xor U12181 (N_12181,N_11842,N_11806);
xnor U12182 (N_12182,N_11925,N_11920);
or U12183 (N_12183,N_11843,N_11875);
nor U12184 (N_12184,N_11851,N_11865);
and U12185 (N_12185,N_11915,N_11814);
xor U12186 (N_12186,N_11848,N_11922);
or U12187 (N_12187,N_11987,N_11852);
or U12188 (N_12188,N_11998,N_11960);
nand U12189 (N_12189,N_11995,N_11900);
nand U12190 (N_12190,N_11954,N_11988);
nor U12191 (N_12191,N_11961,N_11914);
xnor U12192 (N_12192,N_11966,N_11863);
and U12193 (N_12193,N_11923,N_11870);
nand U12194 (N_12194,N_11952,N_11949);
xor U12195 (N_12195,N_11913,N_11944);
or U12196 (N_12196,N_11900,N_11846);
nand U12197 (N_12197,N_11805,N_11855);
or U12198 (N_12198,N_11834,N_11950);
nand U12199 (N_12199,N_11947,N_11820);
xnor U12200 (N_12200,N_12193,N_12086);
or U12201 (N_12201,N_12014,N_12174);
nand U12202 (N_12202,N_12082,N_12033);
and U12203 (N_12203,N_12142,N_12066);
or U12204 (N_12204,N_12047,N_12010);
xnor U12205 (N_12205,N_12091,N_12121);
and U12206 (N_12206,N_12016,N_12058);
nor U12207 (N_12207,N_12188,N_12129);
xor U12208 (N_12208,N_12131,N_12099);
and U12209 (N_12209,N_12022,N_12029);
and U12210 (N_12210,N_12006,N_12171);
nor U12211 (N_12211,N_12081,N_12197);
or U12212 (N_12212,N_12049,N_12113);
and U12213 (N_12213,N_12028,N_12153);
xor U12214 (N_12214,N_12177,N_12013);
and U12215 (N_12215,N_12190,N_12187);
and U12216 (N_12216,N_12196,N_12125);
or U12217 (N_12217,N_12094,N_12052);
nand U12218 (N_12218,N_12191,N_12128);
and U12219 (N_12219,N_12007,N_12057);
nand U12220 (N_12220,N_12186,N_12036);
and U12221 (N_12221,N_12070,N_12048);
nor U12222 (N_12222,N_12141,N_12062);
and U12223 (N_12223,N_12011,N_12067);
or U12224 (N_12224,N_12021,N_12064);
xor U12225 (N_12225,N_12164,N_12076);
or U12226 (N_12226,N_12023,N_12110);
xnor U12227 (N_12227,N_12127,N_12103);
xor U12228 (N_12228,N_12000,N_12092);
nor U12229 (N_12229,N_12138,N_12192);
or U12230 (N_12230,N_12182,N_12104);
xnor U12231 (N_12231,N_12194,N_12156);
and U12232 (N_12232,N_12140,N_12150);
nand U12233 (N_12233,N_12001,N_12050);
xor U12234 (N_12234,N_12089,N_12105);
xnor U12235 (N_12235,N_12137,N_12163);
xor U12236 (N_12236,N_12080,N_12046);
and U12237 (N_12237,N_12043,N_12002);
nand U12238 (N_12238,N_12026,N_12195);
and U12239 (N_12239,N_12093,N_12040);
xnor U12240 (N_12240,N_12199,N_12118);
xor U12241 (N_12241,N_12189,N_12119);
xnor U12242 (N_12242,N_12005,N_12148);
xnor U12243 (N_12243,N_12060,N_12176);
nor U12244 (N_12244,N_12123,N_12095);
or U12245 (N_12245,N_12151,N_12157);
and U12246 (N_12246,N_12160,N_12063);
nor U12247 (N_12247,N_12100,N_12087);
nor U12248 (N_12248,N_12146,N_12068);
or U12249 (N_12249,N_12096,N_12117);
and U12250 (N_12250,N_12008,N_12154);
xor U12251 (N_12251,N_12126,N_12136);
nor U12252 (N_12252,N_12009,N_12030);
nor U12253 (N_12253,N_12085,N_12079);
and U12254 (N_12254,N_12003,N_12069);
and U12255 (N_12255,N_12071,N_12054);
or U12256 (N_12256,N_12149,N_12143);
or U12257 (N_12257,N_12175,N_12165);
and U12258 (N_12258,N_12032,N_12020);
and U12259 (N_12259,N_12098,N_12116);
or U12260 (N_12260,N_12044,N_12097);
nor U12261 (N_12261,N_12162,N_12161);
and U12262 (N_12262,N_12155,N_12139);
nand U12263 (N_12263,N_12132,N_12145);
and U12264 (N_12264,N_12055,N_12042);
or U12265 (N_12265,N_12041,N_12078);
nor U12266 (N_12266,N_12147,N_12166);
and U12267 (N_12267,N_12111,N_12122);
xor U12268 (N_12268,N_12039,N_12077);
nor U12269 (N_12269,N_12124,N_12038);
xnor U12270 (N_12270,N_12073,N_12159);
xor U12271 (N_12271,N_12181,N_12167);
xor U12272 (N_12272,N_12065,N_12061);
nand U12273 (N_12273,N_12072,N_12185);
xnor U12274 (N_12274,N_12180,N_12112);
xor U12275 (N_12275,N_12133,N_12004);
xor U12276 (N_12276,N_12059,N_12088);
xnor U12277 (N_12277,N_12019,N_12018);
nor U12278 (N_12278,N_12090,N_12179);
or U12279 (N_12279,N_12172,N_12115);
nand U12280 (N_12280,N_12144,N_12027);
nor U12281 (N_12281,N_12075,N_12056);
nand U12282 (N_12282,N_12135,N_12102);
nand U12283 (N_12283,N_12045,N_12170);
xor U12284 (N_12284,N_12024,N_12035);
nand U12285 (N_12285,N_12109,N_12130);
nor U12286 (N_12286,N_12169,N_12084);
nor U12287 (N_12287,N_12025,N_12152);
xor U12288 (N_12288,N_12012,N_12178);
nand U12289 (N_12289,N_12114,N_12015);
nand U12290 (N_12290,N_12107,N_12158);
and U12291 (N_12291,N_12101,N_12051);
and U12292 (N_12292,N_12083,N_12053);
and U12293 (N_12293,N_12168,N_12198);
nor U12294 (N_12294,N_12017,N_12183);
xor U12295 (N_12295,N_12120,N_12031);
nand U12296 (N_12296,N_12134,N_12108);
nand U12297 (N_12297,N_12106,N_12037);
xor U12298 (N_12298,N_12034,N_12184);
and U12299 (N_12299,N_12074,N_12173);
xnor U12300 (N_12300,N_12197,N_12173);
xor U12301 (N_12301,N_12024,N_12171);
and U12302 (N_12302,N_12162,N_12053);
and U12303 (N_12303,N_12070,N_12166);
and U12304 (N_12304,N_12123,N_12164);
nor U12305 (N_12305,N_12159,N_12082);
nand U12306 (N_12306,N_12145,N_12129);
and U12307 (N_12307,N_12017,N_12087);
or U12308 (N_12308,N_12199,N_12021);
xor U12309 (N_12309,N_12123,N_12113);
xor U12310 (N_12310,N_12162,N_12029);
xor U12311 (N_12311,N_12190,N_12167);
nand U12312 (N_12312,N_12096,N_12170);
nand U12313 (N_12313,N_12099,N_12148);
or U12314 (N_12314,N_12029,N_12140);
nand U12315 (N_12315,N_12159,N_12122);
and U12316 (N_12316,N_12101,N_12057);
or U12317 (N_12317,N_12083,N_12164);
nor U12318 (N_12318,N_12149,N_12139);
and U12319 (N_12319,N_12164,N_12079);
and U12320 (N_12320,N_12165,N_12092);
nor U12321 (N_12321,N_12144,N_12062);
nand U12322 (N_12322,N_12178,N_12136);
nand U12323 (N_12323,N_12150,N_12044);
nor U12324 (N_12324,N_12089,N_12013);
xor U12325 (N_12325,N_12070,N_12159);
xnor U12326 (N_12326,N_12105,N_12015);
or U12327 (N_12327,N_12069,N_12071);
xor U12328 (N_12328,N_12028,N_12007);
or U12329 (N_12329,N_12009,N_12052);
nand U12330 (N_12330,N_12069,N_12124);
nor U12331 (N_12331,N_12169,N_12132);
or U12332 (N_12332,N_12102,N_12091);
or U12333 (N_12333,N_12102,N_12126);
and U12334 (N_12334,N_12163,N_12050);
or U12335 (N_12335,N_12139,N_12100);
and U12336 (N_12336,N_12149,N_12087);
nor U12337 (N_12337,N_12161,N_12141);
and U12338 (N_12338,N_12188,N_12173);
nand U12339 (N_12339,N_12117,N_12087);
or U12340 (N_12340,N_12104,N_12039);
nor U12341 (N_12341,N_12020,N_12014);
xor U12342 (N_12342,N_12182,N_12134);
nor U12343 (N_12343,N_12147,N_12163);
and U12344 (N_12344,N_12165,N_12007);
nor U12345 (N_12345,N_12096,N_12162);
nand U12346 (N_12346,N_12014,N_12117);
or U12347 (N_12347,N_12069,N_12117);
and U12348 (N_12348,N_12060,N_12102);
nand U12349 (N_12349,N_12116,N_12070);
nor U12350 (N_12350,N_12123,N_12177);
and U12351 (N_12351,N_12102,N_12000);
or U12352 (N_12352,N_12194,N_12144);
or U12353 (N_12353,N_12030,N_12142);
xnor U12354 (N_12354,N_12153,N_12174);
nor U12355 (N_12355,N_12164,N_12105);
and U12356 (N_12356,N_12139,N_12153);
nand U12357 (N_12357,N_12166,N_12163);
nor U12358 (N_12358,N_12058,N_12101);
or U12359 (N_12359,N_12194,N_12029);
and U12360 (N_12360,N_12126,N_12162);
nor U12361 (N_12361,N_12003,N_12027);
or U12362 (N_12362,N_12060,N_12024);
nor U12363 (N_12363,N_12032,N_12027);
or U12364 (N_12364,N_12119,N_12144);
nor U12365 (N_12365,N_12095,N_12183);
and U12366 (N_12366,N_12031,N_12131);
or U12367 (N_12367,N_12059,N_12039);
nand U12368 (N_12368,N_12140,N_12043);
or U12369 (N_12369,N_12120,N_12074);
and U12370 (N_12370,N_12146,N_12011);
nand U12371 (N_12371,N_12116,N_12199);
or U12372 (N_12372,N_12091,N_12150);
nand U12373 (N_12373,N_12101,N_12083);
nand U12374 (N_12374,N_12172,N_12150);
or U12375 (N_12375,N_12023,N_12089);
nor U12376 (N_12376,N_12109,N_12177);
nor U12377 (N_12377,N_12125,N_12175);
nand U12378 (N_12378,N_12192,N_12042);
nand U12379 (N_12379,N_12079,N_12076);
xnor U12380 (N_12380,N_12052,N_12115);
xor U12381 (N_12381,N_12045,N_12111);
or U12382 (N_12382,N_12091,N_12131);
nor U12383 (N_12383,N_12063,N_12042);
nor U12384 (N_12384,N_12094,N_12170);
nand U12385 (N_12385,N_12015,N_12135);
and U12386 (N_12386,N_12163,N_12072);
and U12387 (N_12387,N_12058,N_12060);
or U12388 (N_12388,N_12021,N_12118);
and U12389 (N_12389,N_12048,N_12194);
nor U12390 (N_12390,N_12007,N_12133);
xnor U12391 (N_12391,N_12043,N_12095);
nor U12392 (N_12392,N_12038,N_12025);
nor U12393 (N_12393,N_12009,N_12093);
nand U12394 (N_12394,N_12033,N_12019);
nor U12395 (N_12395,N_12140,N_12157);
or U12396 (N_12396,N_12146,N_12085);
nand U12397 (N_12397,N_12142,N_12181);
or U12398 (N_12398,N_12031,N_12045);
nand U12399 (N_12399,N_12145,N_12191);
nand U12400 (N_12400,N_12393,N_12223);
and U12401 (N_12401,N_12205,N_12243);
nand U12402 (N_12402,N_12224,N_12231);
xnor U12403 (N_12403,N_12322,N_12278);
nor U12404 (N_12404,N_12359,N_12274);
or U12405 (N_12405,N_12375,N_12284);
nand U12406 (N_12406,N_12289,N_12303);
nor U12407 (N_12407,N_12396,N_12313);
or U12408 (N_12408,N_12387,N_12291);
nor U12409 (N_12409,N_12225,N_12228);
or U12410 (N_12410,N_12360,N_12294);
nor U12411 (N_12411,N_12269,N_12301);
and U12412 (N_12412,N_12255,N_12370);
nor U12413 (N_12413,N_12250,N_12397);
nand U12414 (N_12414,N_12212,N_12352);
or U12415 (N_12415,N_12342,N_12209);
xor U12416 (N_12416,N_12325,N_12238);
nand U12417 (N_12417,N_12221,N_12249);
and U12418 (N_12418,N_12245,N_12367);
or U12419 (N_12419,N_12229,N_12399);
nand U12420 (N_12420,N_12283,N_12297);
xor U12421 (N_12421,N_12389,N_12200);
xnor U12422 (N_12422,N_12395,N_12383);
nor U12423 (N_12423,N_12390,N_12234);
nand U12424 (N_12424,N_12203,N_12295);
xnor U12425 (N_12425,N_12305,N_12353);
and U12426 (N_12426,N_12333,N_12369);
and U12427 (N_12427,N_12252,N_12279);
xnor U12428 (N_12428,N_12201,N_12320);
and U12429 (N_12429,N_12288,N_12363);
nor U12430 (N_12430,N_12332,N_12233);
nor U12431 (N_12431,N_12371,N_12351);
nand U12432 (N_12432,N_12366,N_12327);
nor U12433 (N_12433,N_12323,N_12207);
or U12434 (N_12434,N_12385,N_12246);
or U12435 (N_12435,N_12334,N_12382);
nor U12436 (N_12436,N_12347,N_12237);
and U12437 (N_12437,N_12258,N_12319);
nor U12438 (N_12438,N_12378,N_12208);
or U12439 (N_12439,N_12275,N_12310);
nor U12440 (N_12440,N_12321,N_12253);
or U12441 (N_12441,N_12242,N_12247);
xnor U12442 (N_12442,N_12287,N_12339);
nor U12443 (N_12443,N_12219,N_12316);
nor U12444 (N_12444,N_12248,N_12299);
or U12445 (N_12445,N_12239,N_12230);
and U12446 (N_12446,N_12391,N_12376);
and U12447 (N_12447,N_12309,N_12286);
and U12448 (N_12448,N_12361,N_12394);
nand U12449 (N_12449,N_12356,N_12314);
nor U12450 (N_12450,N_12236,N_12348);
nand U12451 (N_12451,N_12218,N_12335);
xnor U12452 (N_12452,N_12285,N_12256);
xnor U12453 (N_12453,N_12254,N_12271);
or U12454 (N_12454,N_12273,N_12340);
xnor U12455 (N_12455,N_12210,N_12355);
or U12456 (N_12456,N_12392,N_12226);
and U12457 (N_12457,N_12280,N_12276);
xor U12458 (N_12458,N_12270,N_12317);
nor U12459 (N_12459,N_12324,N_12337);
nand U12460 (N_12460,N_12222,N_12338);
xnor U12461 (N_12461,N_12341,N_12268);
or U12462 (N_12462,N_12377,N_12331);
and U12463 (N_12463,N_12272,N_12262);
or U12464 (N_12464,N_12257,N_12315);
nor U12465 (N_12465,N_12267,N_12344);
nor U12466 (N_12466,N_12251,N_12362);
nand U12467 (N_12467,N_12346,N_12306);
xor U12468 (N_12468,N_12282,N_12307);
nor U12469 (N_12469,N_12241,N_12296);
or U12470 (N_12470,N_12281,N_12227);
and U12471 (N_12471,N_12350,N_12368);
and U12472 (N_12472,N_12326,N_12345);
and U12473 (N_12473,N_12318,N_12330);
or U12474 (N_12474,N_12343,N_12204);
and U12475 (N_12475,N_12336,N_12213);
or U12476 (N_12476,N_12311,N_12384);
and U12477 (N_12477,N_12398,N_12259);
or U12478 (N_12478,N_12215,N_12232);
and U12479 (N_12479,N_12261,N_12365);
nand U12480 (N_12480,N_12372,N_12386);
or U12481 (N_12481,N_12380,N_12349);
or U12482 (N_12482,N_12308,N_12214);
nor U12483 (N_12483,N_12302,N_12293);
nand U12484 (N_12484,N_12217,N_12374);
xnor U12485 (N_12485,N_12300,N_12373);
nor U12486 (N_12486,N_12292,N_12329);
or U12487 (N_12487,N_12364,N_12235);
or U12488 (N_12488,N_12304,N_12328);
nand U12489 (N_12489,N_12354,N_12381);
nand U12490 (N_12490,N_12211,N_12216);
nor U12491 (N_12491,N_12277,N_12379);
and U12492 (N_12492,N_12220,N_12312);
nor U12493 (N_12493,N_12202,N_12264);
or U12494 (N_12494,N_12358,N_12298);
nor U12495 (N_12495,N_12206,N_12290);
and U12496 (N_12496,N_12263,N_12266);
or U12497 (N_12497,N_12265,N_12260);
nand U12498 (N_12498,N_12244,N_12357);
xnor U12499 (N_12499,N_12240,N_12388);
and U12500 (N_12500,N_12299,N_12315);
nor U12501 (N_12501,N_12200,N_12342);
nand U12502 (N_12502,N_12314,N_12323);
nand U12503 (N_12503,N_12264,N_12358);
and U12504 (N_12504,N_12263,N_12338);
and U12505 (N_12505,N_12249,N_12384);
nor U12506 (N_12506,N_12353,N_12377);
nor U12507 (N_12507,N_12249,N_12211);
xor U12508 (N_12508,N_12358,N_12375);
or U12509 (N_12509,N_12316,N_12325);
nor U12510 (N_12510,N_12397,N_12389);
and U12511 (N_12511,N_12375,N_12252);
nor U12512 (N_12512,N_12388,N_12309);
nand U12513 (N_12513,N_12218,N_12376);
and U12514 (N_12514,N_12327,N_12218);
xor U12515 (N_12515,N_12223,N_12335);
nor U12516 (N_12516,N_12246,N_12202);
and U12517 (N_12517,N_12362,N_12267);
or U12518 (N_12518,N_12217,N_12213);
xor U12519 (N_12519,N_12340,N_12281);
xor U12520 (N_12520,N_12234,N_12223);
and U12521 (N_12521,N_12335,N_12259);
xor U12522 (N_12522,N_12321,N_12322);
or U12523 (N_12523,N_12399,N_12303);
nor U12524 (N_12524,N_12370,N_12394);
or U12525 (N_12525,N_12220,N_12322);
and U12526 (N_12526,N_12302,N_12353);
or U12527 (N_12527,N_12322,N_12237);
nand U12528 (N_12528,N_12276,N_12331);
or U12529 (N_12529,N_12300,N_12286);
nor U12530 (N_12530,N_12217,N_12360);
or U12531 (N_12531,N_12279,N_12327);
xnor U12532 (N_12532,N_12383,N_12241);
nand U12533 (N_12533,N_12261,N_12315);
nand U12534 (N_12534,N_12319,N_12253);
nor U12535 (N_12535,N_12225,N_12363);
and U12536 (N_12536,N_12388,N_12372);
and U12537 (N_12537,N_12312,N_12320);
nand U12538 (N_12538,N_12272,N_12200);
and U12539 (N_12539,N_12307,N_12274);
xor U12540 (N_12540,N_12390,N_12393);
or U12541 (N_12541,N_12343,N_12323);
nor U12542 (N_12542,N_12217,N_12263);
xor U12543 (N_12543,N_12260,N_12378);
nor U12544 (N_12544,N_12393,N_12250);
xnor U12545 (N_12545,N_12343,N_12287);
nor U12546 (N_12546,N_12304,N_12371);
nand U12547 (N_12547,N_12234,N_12258);
xor U12548 (N_12548,N_12367,N_12276);
nor U12549 (N_12549,N_12297,N_12372);
and U12550 (N_12550,N_12352,N_12371);
and U12551 (N_12551,N_12326,N_12238);
xor U12552 (N_12552,N_12248,N_12353);
nor U12553 (N_12553,N_12247,N_12330);
nand U12554 (N_12554,N_12247,N_12296);
or U12555 (N_12555,N_12275,N_12387);
or U12556 (N_12556,N_12315,N_12241);
nor U12557 (N_12557,N_12247,N_12273);
and U12558 (N_12558,N_12318,N_12349);
xor U12559 (N_12559,N_12292,N_12221);
nor U12560 (N_12560,N_12287,N_12384);
nor U12561 (N_12561,N_12242,N_12263);
and U12562 (N_12562,N_12332,N_12365);
xnor U12563 (N_12563,N_12206,N_12237);
and U12564 (N_12564,N_12212,N_12332);
nor U12565 (N_12565,N_12319,N_12385);
or U12566 (N_12566,N_12291,N_12272);
xor U12567 (N_12567,N_12325,N_12221);
xnor U12568 (N_12568,N_12335,N_12263);
and U12569 (N_12569,N_12345,N_12275);
and U12570 (N_12570,N_12205,N_12347);
or U12571 (N_12571,N_12370,N_12240);
nand U12572 (N_12572,N_12242,N_12346);
nand U12573 (N_12573,N_12384,N_12327);
nand U12574 (N_12574,N_12368,N_12265);
and U12575 (N_12575,N_12216,N_12299);
nor U12576 (N_12576,N_12206,N_12250);
nand U12577 (N_12577,N_12380,N_12216);
nand U12578 (N_12578,N_12256,N_12346);
xnor U12579 (N_12579,N_12326,N_12272);
or U12580 (N_12580,N_12232,N_12386);
or U12581 (N_12581,N_12367,N_12359);
and U12582 (N_12582,N_12317,N_12256);
and U12583 (N_12583,N_12217,N_12204);
and U12584 (N_12584,N_12223,N_12327);
nor U12585 (N_12585,N_12296,N_12214);
xnor U12586 (N_12586,N_12243,N_12204);
nand U12587 (N_12587,N_12329,N_12361);
nand U12588 (N_12588,N_12373,N_12367);
nor U12589 (N_12589,N_12281,N_12210);
and U12590 (N_12590,N_12334,N_12365);
nor U12591 (N_12591,N_12328,N_12330);
or U12592 (N_12592,N_12389,N_12333);
nand U12593 (N_12593,N_12338,N_12299);
nor U12594 (N_12594,N_12358,N_12397);
nand U12595 (N_12595,N_12246,N_12342);
xnor U12596 (N_12596,N_12343,N_12309);
nor U12597 (N_12597,N_12350,N_12286);
and U12598 (N_12598,N_12395,N_12203);
or U12599 (N_12599,N_12262,N_12250);
xor U12600 (N_12600,N_12549,N_12584);
nor U12601 (N_12601,N_12466,N_12494);
or U12602 (N_12602,N_12412,N_12437);
xor U12603 (N_12603,N_12527,N_12583);
nand U12604 (N_12604,N_12535,N_12409);
and U12605 (N_12605,N_12483,N_12586);
nand U12606 (N_12606,N_12468,N_12480);
nor U12607 (N_12607,N_12434,N_12533);
nor U12608 (N_12608,N_12499,N_12554);
xor U12609 (N_12609,N_12457,N_12514);
or U12610 (N_12610,N_12492,N_12574);
xor U12611 (N_12611,N_12576,N_12534);
xor U12612 (N_12612,N_12579,N_12495);
or U12613 (N_12613,N_12500,N_12442);
nor U12614 (N_12614,N_12532,N_12454);
xor U12615 (N_12615,N_12530,N_12581);
nor U12616 (N_12616,N_12551,N_12544);
or U12617 (N_12617,N_12450,N_12570);
xor U12618 (N_12618,N_12585,N_12526);
nor U12619 (N_12619,N_12587,N_12496);
and U12620 (N_12620,N_12593,N_12519);
nand U12621 (N_12621,N_12546,N_12426);
and U12622 (N_12622,N_12595,N_12591);
or U12623 (N_12623,N_12474,N_12473);
xnor U12624 (N_12624,N_12522,N_12565);
or U12625 (N_12625,N_12511,N_12460);
nor U12626 (N_12626,N_12540,N_12517);
or U12627 (N_12627,N_12420,N_12542);
nor U12628 (N_12628,N_12582,N_12571);
xor U12629 (N_12629,N_12577,N_12408);
nor U12630 (N_12630,N_12589,N_12558);
xor U12631 (N_12631,N_12413,N_12529);
nor U12632 (N_12632,N_12539,N_12553);
and U12633 (N_12633,N_12507,N_12493);
and U12634 (N_12634,N_12520,N_12428);
or U12635 (N_12635,N_12518,N_12489);
nand U12636 (N_12636,N_12566,N_12599);
nand U12637 (N_12637,N_12485,N_12464);
xnor U12638 (N_12638,N_12543,N_12438);
xnor U12639 (N_12639,N_12567,N_12479);
nor U12640 (N_12640,N_12557,N_12417);
nor U12641 (N_12641,N_12404,N_12429);
and U12642 (N_12642,N_12537,N_12422);
xor U12643 (N_12643,N_12451,N_12509);
and U12644 (N_12644,N_12431,N_12414);
nor U12645 (N_12645,N_12564,N_12555);
xor U12646 (N_12646,N_12508,N_12447);
nand U12647 (N_12647,N_12559,N_12596);
or U12648 (N_12648,N_12419,N_12456);
nand U12649 (N_12649,N_12590,N_12427);
nor U12650 (N_12650,N_12523,N_12401);
or U12651 (N_12651,N_12580,N_12594);
nand U12652 (N_12652,N_12488,N_12424);
or U12653 (N_12653,N_12563,N_12423);
and U12654 (N_12654,N_12503,N_12512);
xnor U12655 (N_12655,N_12405,N_12575);
or U12656 (N_12656,N_12536,N_12418);
nor U12657 (N_12657,N_12463,N_12562);
nand U12658 (N_12658,N_12446,N_12421);
and U12659 (N_12659,N_12545,N_12505);
nor U12660 (N_12660,N_12462,N_12498);
or U12661 (N_12661,N_12455,N_12504);
nand U12662 (N_12662,N_12547,N_12502);
nand U12663 (N_12663,N_12470,N_12541);
xnor U12664 (N_12664,N_12550,N_12400);
xor U12665 (N_12665,N_12482,N_12432);
and U12666 (N_12666,N_12449,N_12531);
xor U12667 (N_12667,N_12411,N_12588);
and U12668 (N_12668,N_12556,N_12516);
nand U12669 (N_12669,N_12416,N_12469);
and U12670 (N_12670,N_12406,N_12441);
nand U12671 (N_12671,N_12436,N_12524);
and U12672 (N_12672,N_12458,N_12445);
nor U12673 (N_12673,N_12528,N_12501);
nor U12674 (N_12674,N_12568,N_12578);
nand U12675 (N_12675,N_12439,N_12475);
or U12676 (N_12676,N_12476,N_12515);
or U12677 (N_12677,N_12561,N_12425);
xnor U12678 (N_12678,N_12560,N_12403);
and U12679 (N_12679,N_12448,N_12435);
and U12680 (N_12680,N_12513,N_12478);
nor U12681 (N_12681,N_12452,N_12459);
xor U12682 (N_12682,N_12402,N_12490);
nor U12683 (N_12683,N_12597,N_12444);
nand U12684 (N_12684,N_12486,N_12491);
nand U12685 (N_12685,N_12465,N_12471);
nand U12686 (N_12686,N_12453,N_12472);
nand U12687 (N_12687,N_12484,N_12481);
xor U12688 (N_12688,N_12497,N_12430);
nand U12689 (N_12689,N_12552,N_12407);
nand U12690 (N_12690,N_12506,N_12433);
nand U12691 (N_12691,N_12598,N_12410);
xor U12692 (N_12692,N_12487,N_12510);
or U12693 (N_12693,N_12467,N_12440);
nand U12694 (N_12694,N_12572,N_12525);
xor U12695 (N_12695,N_12521,N_12443);
nor U12696 (N_12696,N_12461,N_12592);
xnor U12697 (N_12697,N_12548,N_12573);
and U12698 (N_12698,N_12538,N_12415);
or U12699 (N_12699,N_12569,N_12477);
xnor U12700 (N_12700,N_12545,N_12574);
and U12701 (N_12701,N_12540,N_12590);
xnor U12702 (N_12702,N_12509,N_12581);
nand U12703 (N_12703,N_12562,N_12523);
or U12704 (N_12704,N_12536,N_12508);
xnor U12705 (N_12705,N_12483,N_12402);
nor U12706 (N_12706,N_12450,N_12597);
nand U12707 (N_12707,N_12481,N_12434);
and U12708 (N_12708,N_12557,N_12574);
or U12709 (N_12709,N_12484,N_12477);
or U12710 (N_12710,N_12512,N_12524);
xnor U12711 (N_12711,N_12418,N_12406);
xor U12712 (N_12712,N_12500,N_12531);
nor U12713 (N_12713,N_12515,N_12570);
or U12714 (N_12714,N_12472,N_12564);
nor U12715 (N_12715,N_12506,N_12508);
and U12716 (N_12716,N_12560,N_12587);
or U12717 (N_12717,N_12544,N_12407);
or U12718 (N_12718,N_12439,N_12534);
and U12719 (N_12719,N_12587,N_12479);
nand U12720 (N_12720,N_12533,N_12466);
nor U12721 (N_12721,N_12599,N_12460);
or U12722 (N_12722,N_12433,N_12403);
xnor U12723 (N_12723,N_12505,N_12407);
nor U12724 (N_12724,N_12595,N_12474);
nor U12725 (N_12725,N_12449,N_12483);
or U12726 (N_12726,N_12446,N_12567);
or U12727 (N_12727,N_12515,N_12528);
xnor U12728 (N_12728,N_12546,N_12473);
or U12729 (N_12729,N_12519,N_12465);
and U12730 (N_12730,N_12553,N_12484);
nand U12731 (N_12731,N_12586,N_12562);
nand U12732 (N_12732,N_12533,N_12547);
xnor U12733 (N_12733,N_12554,N_12473);
and U12734 (N_12734,N_12547,N_12468);
nand U12735 (N_12735,N_12531,N_12465);
xor U12736 (N_12736,N_12470,N_12562);
nand U12737 (N_12737,N_12407,N_12468);
nor U12738 (N_12738,N_12539,N_12521);
xnor U12739 (N_12739,N_12446,N_12451);
nand U12740 (N_12740,N_12506,N_12570);
xor U12741 (N_12741,N_12513,N_12402);
xnor U12742 (N_12742,N_12574,N_12444);
xor U12743 (N_12743,N_12449,N_12511);
nand U12744 (N_12744,N_12558,N_12576);
and U12745 (N_12745,N_12450,N_12560);
and U12746 (N_12746,N_12596,N_12598);
nand U12747 (N_12747,N_12475,N_12570);
or U12748 (N_12748,N_12499,N_12566);
and U12749 (N_12749,N_12520,N_12542);
or U12750 (N_12750,N_12514,N_12594);
or U12751 (N_12751,N_12486,N_12412);
and U12752 (N_12752,N_12440,N_12404);
nor U12753 (N_12753,N_12458,N_12523);
or U12754 (N_12754,N_12570,N_12562);
nor U12755 (N_12755,N_12576,N_12578);
and U12756 (N_12756,N_12424,N_12401);
or U12757 (N_12757,N_12427,N_12484);
xor U12758 (N_12758,N_12585,N_12494);
and U12759 (N_12759,N_12479,N_12530);
nor U12760 (N_12760,N_12488,N_12498);
or U12761 (N_12761,N_12481,N_12407);
nand U12762 (N_12762,N_12478,N_12471);
or U12763 (N_12763,N_12534,N_12429);
and U12764 (N_12764,N_12481,N_12457);
and U12765 (N_12765,N_12511,N_12480);
xor U12766 (N_12766,N_12531,N_12479);
nand U12767 (N_12767,N_12512,N_12499);
and U12768 (N_12768,N_12418,N_12496);
or U12769 (N_12769,N_12462,N_12548);
nor U12770 (N_12770,N_12561,N_12436);
xnor U12771 (N_12771,N_12545,N_12530);
nor U12772 (N_12772,N_12426,N_12441);
xnor U12773 (N_12773,N_12593,N_12549);
and U12774 (N_12774,N_12468,N_12552);
nor U12775 (N_12775,N_12499,N_12401);
or U12776 (N_12776,N_12426,N_12525);
nand U12777 (N_12777,N_12546,N_12488);
and U12778 (N_12778,N_12404,N_12412);
or U12779 (N_12779,N_12529,N_12418);
nand U12780 (N_12780,N_12548,N_12523);
nand U12781 (N_12781,N_12432,N_12461);
xor U12782 (N_12782,N_12409,N_12425);
xor U12783 (N_12783,N_12461,N_12539);
or U12784 (N_12784,N_12500,N_12598);
nand U12785 (N_12785,N_12570,N_12595);
xor U12786 (N_12786,N_12413,N_12573);
or U12787 (N_12787,N_12584,N_12466);
and U12788 (N_12788,N_12496,N_12561);
nand U12789 (N_12789,N_12532,N_12512);
or U12790 (N_12790,N_12513,N_12539);
and U12791 (N_12791,N_12515,N_12411);
and U12792 (N_12792,N_12568,N_12431);
and U12793 (N_12793,N_12467,N_12486);
and U12794 (N_12794,N_12556,N_12507);
xnor U12795 (N_12795,N_12455,N_12568);
and U12796 (N_12796,N_12516,N_12572);
xor U12797 (N_12797,N_12498,N_12448);
or U12798 (N_12798,N_12448,N_12593);
xor U12799 (N_12799,N_12446,N_12493);
nor U12800 (N_12800,N_12620,N_12661);
and U12801 (N_12801,N_12700,N_12645);
and U12802 (N_12802,N_12657,N_12693);
xor U12803 (N_12803,N_12626,N_12696);
xnor U12804 (N_12804,N_12612,N_12779);
or U12805 (N_12805,N_12793,N_12778);
xnor U12806 (N_12806,N_12752,N_12791);
xnor U12807 (N_12807,N_12738,N_12601);
nand U12808 (N_12808,N_12756,N_12740);
or U12809 (N_12809,N_12745,N_12730);
or U12810 (N_12810,N_12610,N_12634);
or U12811 (N_12811,N_12753,N_12721);
or U12812 (N_12812,N_12616,N_12695);
xnor U12813 (N_12813,N_12764,N_12703);
nand U12814 (N_12814,N_12788,N_12751);
xnor U12815 (N_12815,N_12602,N_12706);
or U12816 (N_12816,N_12773,N_12650);
and U12817 (N_12817,N_12737,N_12698);
xnor U12818 (N_12818,N_12609,N_12614);
and U12819 (N_12819,N_12799,N_12600);
nand U12820 (N_12820,N_12789,N_12760);
xnor U12821 (N_12821,N_12627,N_12763);
or U12822 (N_12822,N_12683,N_12794);
nor U12823 (N_12823,N_12603,N_12750);
nand U12824 (N_12824,N_12735,N_12783);
xnor U12825 (N_12825,N_12605,N_12649);
xnor U12826 (N_12826,N_12767,N_12618);
or U12827 (N_12827,N_12734,N_12708);
and U12828 (N_12828,N_12632,N_12728);
or U12829 (N_12829,N_12727,N_12768);
xor U12830 (N_12830,N_12607,N_12687);
nand U12831 (N_12831,N_12672,N_12654);
nand U12832 (N_12832,N_12670,N_12772);
or U12833 (N_12833,N_12784,N_12686);
xnor U12834 (N_12834,N_12780,N_12655);
xor U12835 (N_12835,N_12606,N_12682);
and U12836 (N_12836,N_12613,N_12786);
nand U12837 (N_12837,N_12717,N_12676);
xor U12838 (N_12838,N_12771,N_12795);
or U12839 (N_12839,N_12642,N_12707);
xnor U12840 (N_12840,N_12675,N_12688);
or U12841 (N_12841,N_12636,N_12774);
nand U12842 (N_12842,N_12665,N_12662);
and U12843 (N_12843,N_12684,N_12619);
or U12844 (N_12844,N_12705,N_12736);
and U12845 (N_12845,N_12625,N_12630);
nor U12846 (N_12846,N_12716,N_12726);
xnor U12847 (N_12847,N_12741,N_12617);
or U12848 (N_12848,N_12658,N_12622);
or U12849 (N_12849,N_12667,N_12638);
nor U12850 (N_12850,N_12790,N_12798);
xor U12851 (N_12851,N_12785,N_12694);
and U12852 (N_12852,N_12690,N_12781);
nor U12853 (N_12853,N_12673,N_12663);
nor U12854 (N_12854,N_12646,N_12651);
or U12855 (N_12855,N_12758,N_12677);
or U12856 (N_12856,N_12724,N_12787);
or U12857 (N_12857,N_12608,N_12628);
and U12858 (N_12858,N_12635,N_12719);
xor U12859 (N_12859,N_12762,N_12692);
xnor U12860 (N_12860,N_12659,N_12652);
xnor U12861 (N_12861,N_12797,N_12742);
and U12862 (N_12862,N_12680,N_12660);
nand U12863 (N_12863,N_12713,N_12715);
nor U12864 (N_12864,N_12776,N_12624);
or U12865 (N_12865,N_12639,N_12647);
or U12866 (N_12866,N_12664,N_12669);
nor U12867 (N_12867,N_12744,N_12621);
and U12868 (N_12868,N_12691,N_12748);
or U12869 (N_12869,N_12743,N_12729);
or U12870 (N_12870,N_12754,N_12711);
xnor U12871 (N_12871,N_12689,N_12701);
nand U12872 (N_12872,N_12604,N_12653);
nor U12873 (N_12873,N_12755,N_12770);
nor U12874 (N_12874,N_12666,N_12709);
or U12875 (N_12875,N_12641,N_12629);
and U12876 (N_12876,N_12796,N_12759);
nor U12877 (N_12877,N_12697,N_12777);
nand U12878 (N_12878,N_12674,N_12656);
xnor U12879 (N_12879,N_12668,N_12643);
or U12880 (N_12880,N_12723,N_12681);
or U12881 (N_12881,N_12765,N_12733);
or U12882 (N_12882,N_12704,N_12633);
and U12883 (N_12883,N_12637,N_12611);
nand U12884 (N_12884,N_12761,N_12766);
nand U12885 (N_12885,N_12747,N_12648);
and U12886 (N_12886,N_12644,N_12749);
or U12887 (N_12887,N_12722,N_12720);
and U12888 (N_12888,N_12710,N_12782);
nand U12889 (N_12889,N_12640,N_12731);
xnor U12890 (N_12890,N_12769,N_12623);
nor U12891 (N_12891,N_12746,N_12725);
xor U12892 (N_12892,N_12699,N_12792);
nand U12893 (N_12893,N_12775,N_12615);
or U12894 (N_12894,N_12702,N_12714);
or U12895 (N_12895,N_12718,N_12712);
nor U12896 (N_12896,N_12739,N_12732);
xnor U12897 (N_12897,N_12631,N_12757);
and U12898 (N_12898,N_12679,N_12678);
nor U12899 (N_12899,N_12685,N_12671);
xnor U12900 (N_12900,N_12745,N_12744);
nand U12901 (N_12901,N_12755,N_12749);
and U12902 (N_12902,N_12792,N_12668);
nor U12903 (N_12903,N_12709,N_12692);
or U12904 (N_12904,N_12727,N_12741);
xnor U12905 (N_12905,N_12637,N_12778);
nand U12906 (N_12906,N_12748,N_12695);
and U12907 (N_12907,N_12621,N_12728);
nor U12908 (N_12908,N_12619,N_12663);
xnor U12909 (N_12909,N_12708,N_12658);
or U12910 (N_12910,N_12679,N_12697);
or U12911 (N_12911,N_12789,N_12672);
nor U12912 (N_12912,N_12658,N_12628);
nor U12913 (N_12913,N_12752,N_12693);
nand U12914 (N_12914,N_12692,N_12719);
and U12915 (N_12915,N_12661,N_12724);
or U12916 (N_12916,N_12725,N_12763);
nand U12917 (N_12917,N_12638,N_12697);
nand U12918 (N_12918,N_12754,N_12660);
or U12919 (N_12919,N_12726,N_12678);
or U12920 (N_12920,N_12750,N_12726);
or U12921 (N_12921,N_12653,N_12674);
or U12922 (N_12922,N_12603,N_12712);
nor U12923 (N_12923,N_12606,N_12612);
nor U12924 (N_12924,N_12626,N_12768);
nor U12925 (N_12925,N_12761,N_12750);
or U12926 (N_12926,N_12697,N_12609);
nand U12927 (N_12927,N_12684,N_12780);
xnor U12928 (N_12928,N_12676,N_12602);
nand U12929 (N_12929,N_12755,N_12759);
or U12930 (N_12930,N_12690,N_12609);
nand U12931 (N_12931,N_12685,N_12665);
nand U12932 (N_12932,N_12616,N_12772);
and U12933 (N_12933,N_12634,N_12741);
nor U12934 (N_12934,N_12671,N_12620);
or U12935 (N_12935,N_12601,N_12749);
nor U12936 (N_12936,N_12670,N_12612);
nor U12937 (N_12937,N_12623,N_12784);
xor U12938 (N_12938,N_12786,N_12601);
and U12939 (N_12939,N_12771,N_12754);
xor U12940 (N_12940,N_12765,N_12773);
xnor U12941 (N_12941,N_12665,N_12687);
nor U12942 (N_12942,N_12702,N_12740);
xor U12943 (N_12943,N_12700,N_12761);
xnor U12944 (N_12944,N_12612,N_12691);
and U12945 (N_12945,N_12738,N_12757);
nand U12946 (N_12946,N_12651,N_12683);
nor U12947 (N_12947,N_12677,N_12691);
and U12948 (N_12948,N_12732,N_12677);
xor U12949 (N_12949,N_12622,N_12695);
or U12950 (N_12950,N_12655,N_12789);
and U12951 (N_12951,N_12796,N_12676);
nand U12952 (N_12952,N_12605,N_12722);
nor U12953 (N_12953,N_12706,N_12744);
or U12954 (N_12954,N_12696,N_12708);
nand U12955 (N_12955,N_12724,N_12652);
xnor U12956 (N_12956,N_12784,N_12709);
and U12957 (N_12957,N_12632,N_12704);
nor U12958 (N_12958,N_12752,N_12783);
and U12959 (N_12959,N_12603,N_12687);
and U12960 (N_12960,N_12741,N_12733);
xnor U12961 (N_12961,N_12675,N_12620);
and U12962 (N_12962,N_12715,N_12708);
nand U12963 (N_12963,N_12795,N_12627);
xnor U12964 (N_12964,N_12606,N_12635);
nor U12965 (N_12965,N_12730,N_12633);
or U12966 (N_12966,N_12618,N_12736);
xor U12967 (N_12967,N_12620,N_12799);
and U12968 (N_12968,N_12763,N_12672);
nor U12969 (N_12969,N_12763,N_12607);
nand U12970 (N_12970,N_12796,N_12664);
nor U12971 (N_12971,N_12686,N_12675);
nand U12972 (N_12972,N_12778,N_12617);
and U12973 (N_12973,N_12659,N_12715);
nand U12974 (N_12974,N_12728,N_12654);
nand U12975 (N_12975,N_12705,N_12617);
and U12976 (N_12976,N_12748,N_12620);
nor U12977 (N_12977,N_12660,N_12635);
nor U12978 (N_12978,N_12674,N_12632);
and U12979 (N_12979,N_12663,N_12660);
and U12980 (N_12980,N_12768,N_12760);
and U12981 (N_12981,N_12728,N_12740);
xnor U12982 (N_12982,N_12622,N_12778);
nand U12983 (N_12983,N_12649,N_12643);
nand U12984 (N_12984,N_12622,N_12790);
and U12985 (N_12985,N_12748,N_12736);
or U12986 (N_12986,N_12695,N_12646);
nor U12987 (N_12987,N_12625,N_12783);
nor U12988 (N_12988,N_12789,N_12633);
nor U12989 (N_12989,N_12799,N_12739);
nor U12990 (N_12990,N_12677,N_12602);
nor U12991 (N_12991,N_12759,N_12688);
or U12992 (N_12992,N_12677,N_12641);
or U12993 (N_12993,N_12791,N_12636);
xor U12994 (N_12994,N_12661,N_12672);
or U12995 (N_12995,N_12645,N_12682);
and U12996 (N_12996,N_12633,N_12715);
or U12997 (N_12997,N_12614,N_12773);
or U12998 (N_12998,N_12747,N_12687);
xor U12999 (N_12999,N_12624,N_12638);
nand U13000 (N_13000,N_12956,N_12808);
nor U13001 (N_13001,N_12957,N_12961);
or U13002 (N_13002,N_12828,N_12915);
nand U13003 (N_13003,N_12998,N_12891);
nand U13004 (N_13004,N_12838,N_12805);
or U13005 (N_13005,N_12860,N_12960);
and U13006 (N_13006,N_12879,N_12898);
and U13007 (N_13007,N_12839,N_12804);
xor U13008 (N_13008,N_12917,N_12883);
or U13009 (N_13009,N_12858,N_12822);
nand U13010 (N_13010,N_12945,N_12938);
and U13011 (N_13011,N_12921,N_12829);
xnor U13012 (N_13012,N_12847,N_12834);
xnor U13013 (N_13013,N_12918,N_12954);
xor U13014 (N_13014,N_12888,N_12959);
nand U13015 (N_13015,N_12920,N_12801);
or U13016 (N_13016,N_12992,N_12859);
xor U13017 (N_13017,N_12955,N_12984);
xnor U13018 (N_13018,N_12977,N_12873);
and U13019 (N_13019,N_12816,N_12867);
xor U13020 (N_13020,N_12999,N_12944);
nor U13021 (N_13021,N_12884,N_12963);
and U13022 (N_13022,N_12830,N_12856);
and U13023 (N_13023,N_12831,N_12893);
xnor U13024 (N_13024,N_12866,N_12901);
and U13025 (N_13025,N_12947,N_12911);
or U13026 (N_13026,N_12827,N_12853);
nor U13027 (N_13027,N_12833,N_12979);
nand U13028 (N_13028,N_12933,N_12800);
nand U13029 (N_13029,N_12820,N_12973);
nand U13030 (N_13030,N_12880,N_12906);
nand U13031 (N_13031,N_12872,N_12824);
or U13032 (N_13032,N_12912,N_12886);
xnor U13033 (N_13033,N_12821,N_12807);
and U13034 (N_13034,N_12812,N_12953);
nand U13035 (N_13035,N_12882,N_12836);
or U13036 (N_13036,N_12842,N_12975);
or U13037 (N_13037,N_12892,N_12943);
or U13038 (N_13038,N_12934,N_12914);
xnor U13039 (N_13039,N_12994,N_12976);
nand U13040 (N_13040,N_12810,N_12923);
nor U13041 (N_13041,N_12855,N_12935);
or U13042 (N_13042,N_12857,N_12925);
or U13043 (N_13043,N_12968,N_12826);
or U13044 (N_13044,N_12815,N_12969);
nand U13045 (N_13045,N_12970,N_12889);
xor U13046 (N_13046,N_12835,N_12930);
nor U13047 (N_13047,N_12868,N_12951);
or U13048 (N_13048,N_12817,N_12991);
or U13049 (N_13049,N_12851,N_12907);
or U13050 (N_13050,N_12978,N_12997);
xnor U13051 (N_13051,N_12983,N_12927);
and U13052 (N_13052,N_12931,N_12908);
or U13053 (N_13053,N_12965,N_12878);
and U13054 (N_13054,N_12809,N_12823);
nand U13055 (N_13055,N_12940,N_12926);
nor U13056 (N_13056,N_12967,N_12982);
nand U13057 (N_13057,N_12950,N_12952);
xor U13058 (N_13058,N_12871,N_12900);
or U13059 (N_13059,N_12837,N_12806);
nand U13060 (N_13060,N_12895,N_12985);
nand U13061 (N_13061,N_12802,N_12845);
xor U13062 (N_13062,N_12894,N_12850);
nor U13063 (N_13063,N_12986,N_12971);
xor U13064 (N_13064,N_12864,N_12885);
nor U13065 (N_13065,N_12819,N_12863);
xnor U13066 (N_13066,N_12928,N_12877);
and U13067 (N_13067,N_12909,N_12936);
or U13068 (N_13068,N_12876,N_12814);
and U13069 (N_13069,N_12966,N_12870);
or U13070 (N_13070,N_12903,N_12843);
xnor U13071 (N_13071,N_12958,N_12840);
nand U13072 (N_13072,N_12993,N_12916);
or U13073 (N_13073,N_12846,N_12939);
and U13074 (N_13074,N_12854,N_12989);
and U13075 (N_13075,N_12913,N_12905);
nor U13076 (N_13076,N_12813,N_12881);
xnor U13077 (N_13077,N_12988,N_12841);
nor U13078 (N_13078,N_12972,N_12910);
and U13079 (N_13079,N_12981,N_12896);
xor U13080 (N_13080,N_12849,N_12904);
or U13081 (N_13081,N_12941,N_12890);
and U13082 (N_13082,N_12832,N_12937);
nand U13083 (N_13083,N_12932,N_12990);
nand U13084 (N_13084,N_12811,N_12869);
xor U13085 (N_13085,N_12803,N_12922);
xnor U13086 (N_13086,N_12980,N_12862);
nand U13087 (N_13087,N_12962,N_12848);
nor U13088 (N_13088,N_12865,N_12818);
and U13089 (N_13089,N_12996,N_12924);
nand U13090 (N_13090,N_12987,N_12995);
or U13091 (N_13091,N_12887,N_12861);
nand U13092 (N_13092,N_12948,N_12946);
xnor U13093 (N_13093,N_12875,N_12899);
and U13094 (N_13094,N_12919,N_12942);
and U13095 (N_13095,N_12825,N_12844);
or U13096 (N_13096,N_12897,N_12974);
xor U13097 (N_13097,N_12949,N_12964);
xnor U13098 (N_13098,N_12929,N_12852);
nand U13099 (N_13099,N_12874,N_12902);
or U13100 (N_13100,N_12943,N_12905);
and U13101 (N_13101,N_12989,N_12901);
nor U13102 (N_13102,N_12907,N_12933);
and U13103 (N_13103,N_12880,N_12986);
nand U13104 (N_13104,N_12904,N_12887);
xor U13105 (N_13105,N_12970,N_12821);
nor U13106 (N_13106,N_12836,N_12852);
or U13107 (N_13107,N_12949,N_12914);
and U13108 (N_13108,N_12883,N_12946);
or U13109 (N_13109,N_12978,N_12957);
xor U13110 (N_13110,N_12819,N_12890);
nor U13111 (N_13111,N_12824,N_12802);
nand U13112 (N_13112,N_12873,N_12842);
xor U13113 (N_13113,N_12862,N_12998);
nor U13114 (N_13114,N_12903,N_12985);
and U13115 (N_13115,N_12889,N_12829);
nand U13116 (N_13116,N_12985,N_12846);
and U13117 (N_13117,N_12941,N_12979);
nor U13118 (N_13118,N_12886,N_12868);
or U13119 (N_13119,N_12896,N_12876);
xnor U13120 (N_13120,N_12875,N_12825);
and U13121 (N_13121,N_12826,N_12827);
xor U13122 (N_13122,N_12907,N_12892);
nand U13123 (N_13123,N_12919,N_12983);
nor U13124 (N_13124,N_12985,N_12935);
nor U13125 (N_13125,N_12932,N_12839);
nor U13126 (N_13126,N_12975,N_12937);
or U13127 (N_13127,N_12994,N_12986);
nand U13128 (N_13128,N_12826,N_12993);
nand U13129 (N_13129,N_12851,N_12929);
xnor U13130 (N_13130,N_12922,N_12970);
or U13131 (N_13131,N_12942,N_12924);
or U13132 (N_13132,N_12862,N_12918);
and U13133 (N_13133,N_12886,N_12988);
or U13134 (N_13134,N_12932,N_12957);
or U13135 (N_13135,N_12997,N_12839);
nor U13136 (N_13136,N_12816,N_12817);
nand U13137 (N_13137,N_12906,N_12912);
xor U13138 (N_13138,N_12997,N_12836);
nand U13139 (N_13139,N_12905,N_12895);
or U13140 (N_13140,N_12801,N_12845);
nor U13141 (N_13141,N_12915,N_12819);
nand U13142 (N_13142,N_12842,N_12800);
nand U13143 (N_13143,N_12992,N_12882);
xor U13144 (N_13144,N_12891,N_12871);
nor U13145 (N_13145,N_12862,N_12817);
nor U13146 (N_13146,N_12868,N_12998);
nor U13147 (N_13147,N_12955,N_12959);
nor U13148 (N_13148,N_12848,N_12941);
nand U13149 (N_13149,N_12848,N_12895);
or U13150 (N_13150,N_12999,N_12927);
or U13151 (N_13151,N_12828,N_12886);
nand U13152 (N_13152,N_12982,N_12800);
and U13153 (N_13153,N_12818,N_12888);
or U13154 (N_13154,N_12905,N_12936);
xnor U13155 (N_13155,N_12955,N_12975);
and U13156 (N_13156,N_12848,N_12832);
nand U13157 (N_13157,N_12853,N_12804);
and U13158 (N_13158,N_12988,N_12805);
xnor U13159 (N_13159,N_12953,N_12929);
nor U13160 (N_13160,N_12867,N_12989);
or U13161 (N_13161,N_12864,N_12919);
xor U13162 (N_13162,N_12945,N_12970);
nand U13163 (N_13163,N_12978,N_12804);
xnor U13164 (N_13164,N_12945,N_12914);
nand U13165 (N_13165,N_12830,N_12902);
and U13166 (N_13166,N_12848,N_12936);
nand U13167 (N_13167,N_12849,N_12958);
and U13168 (N_13168,N_12919,N_12896);
nand U13169 (N_13169,N_12928,N_12836);
nor U13170 (N_13170,N_12805,N_12992);
xor U13171 (N_13171,N_12993,N_12978);
or U13172 (N_13172,N_12964,N_12895);
xnor U13173 (N_13173,N_12891,N_12814);
or U13174 (N_13174,N_12926,N_12952);
nor U13175 (N_13175,N_12845,N_12966);
nor U13176 (N_13176,N_12867,N_12980);
nand U13177 (N_13177,N_12947,N_12878);
or U13178 (N_13178,N_12930,N_12877);
and U13179 (N_13179,N_12830,N_12883);
or U13180 (N_13180,N_12999,N_12930);
xnor U13181 (N_13181,N_12821,N_12941);
nor U13182 (N_13182,N_12999,N_12863);
xnor U13183 (N_13183,N_12864,N_12972);
and U13184 (N_13184,N_12994,N_12907);
nand U13185 (N_13185,N_12957,N_12835);
nand U13186 (N_13186,N_12954,N_12949);
or U13187 (N_13187,N_12856,N_12963);
or U13188 (N_13188,N_12875,N_12969);
xnor U13189 (N_13189,N_12994,N_12873);
nand U13190 (N_13190,N_12956,N_12914);
or U13191 (N_13191,N_12814,N_12829);
xor U13192 (N_13192,N_12891,N_12863);
xnor U13193 (N_13193,N_12845,N_12895);
or U13194 (N_13194,N_12957,N_12997);
or U13195 (N_13195,N_12853,N_12919);
or U13196 (N_13196,N_12990,N_12826);
nand U13197 (N_13197,N_12883,N_12928);
xor U13198 (N_13198,N_12810,N_12981);
nor U13199 (N_13199,N_12834,N_12848);
xnor U13200 (N_13200,N_13136,N_13043);
or U13201 (N_13201,N_13147,N_13013);
and U13202 (N_13202,N_13022,N_13027);
and U13203 (N_13203,N_13011,N_13128);
nor U13204 (N_13204,N_13140,N_13187);
and U13205 (N_13205,N_13077,N_13132);
nor U13206 (N_13206,N_13113,N_13193);
nand U13207 (N_13207,N_13095,N_13196);
or U13208 (N_13208,N_13165,N_13081);
nor U13209 (N_13209,N_13171,N_13084);
or U13210 (N_13210,N_13024,N_13007);
nand U13211 (N_13211,N_13110,N_13180);
nand U13212 (N_13212,N_13177,N_13099);
nor U13213 (N_13213,N_13109,N_13048);
xor U13214 (N_13214,N_13032,N_13191);
and U13215 (N_13215,N_13160,N_13061);
or U13216 (N_13216,N_13037,N_13148);
nand U13217 (N_13217,N_13133,N_13166);
nor U13218 (N_13218,N_13112,N_13069);
nor U13219 (N_13219,N_13195,N_13044);
or U13220 (N_13220,N_13145,N_13130);
and U13221 (N_13221,N_13121,N_13129);
or U13222 (N_13222,N_13036,N_13010);
xnor U13223 (N_13223,N_13019,N_13008);
or U13224 (N_13224,N_13197,N_13068);
nor U13225 (N_13225,N_13033,N_13015);
and U13226 (N_13226,N_13003,N_13001);
nand U13227 (N_13227,N_13038,N_13065);
xnor U13228 (N_13228,N_13163,N_13098);
nand U13229 (N_13229,N_13073,N_13169);
xor U13230 (N_13230,N_13137,N_13090);
nor U13231 (N_13231,N_13017,N_13067);
xnor U13232 (N_13232,N_13083,N_13192);
nor U13233 (N_13233,N_13086,N_13035);
or U13234 (N_13234,N_13088,N_13093);
or U13235 (N_13235,N_13190,N_13047);
and U13236 (N_13236,N_13114,N_13164);
and U13237 (N_13237,N_13054,N_13102);
nor U13238 (N_13238,N_13025,N_13118);
and U13239 (N_13239,N_13080,N_13091);
or U13240 (N_13240,N_13076,N_13006);
nand U13241 (N_13241,N_13143,N_13116);
and U13242 (N_13242,N_13170,N_13012);
xor U13243 (N_13243,N_13018,N_13058);
nand U13244 (N_13244,N_13146,N_13066);
xor U13245 (N_13245,N_13049,N_13153);
or U13246 (N_13246,N_13052,N_13167);
or U13247 (N_13247,N_13004,N_13138);
xor U13248 (N_13248,N_13123,N_13060);
xnor U13249 (N_13249,N_13087,N_13016);
nand U13250 (N_13250,N_13055,N_13040);
and U13251 (N_13251,N_13174,N_13021);
or U13252 (N_13252,N_13152,N_13030);
or U13253 (N_13253,N_13062,N_13135);
nand U13254 (N_13254,N_13131,N_13141);
or U13255 (N_13255,N_13119,N_13186);
nor U13256 (N_13256,N_13057,N_13176);
xor U13257 (N_13257,N_13199,N_13059);
nor U13258 (N_13258,N_13162,N_13009);
and U13259 (N_13259,N_13144,N_13026);
nand U13260 (N_13260,N_13126,N_13155);
nor U13261 (N_13261,N_13074,N_13103);
and U13262 (N_13262,N_13122,N_13082);
and U13263 (N_13263,N_13000,N_13188);
xnor U13264 (N_13264,N_13161,N_13168);
xor U13265 (N_13265,N_13184,N_13002);
xor U13266 (N_13266,N_13064,N_13101);
xor U13267 (N_13267,N_13127,N_13031);
and U13268 (N_13268,N_13142,N_13106);
nand U13269 (N_13269,N_13178,N_13120);
or U13270 (N_13270,N_13124,N_13045);
and U13271 (N_13271,N_13089,N_13046);
nand U13272 (N_13272,N_13117,N_13014);
nor U13273 (N_13273,N_13149,N_13151);
nand U13274 (N_13274,N_13198,N_13154);
xnor U13275 (N_13275,N_13042,N_13039);
nand U13276 (N_13276,N_13096,N_13071);
xnor U13277 (N_13277,N_13105,N_13183);
and U13278 (N_13278,N_13097,N_13150);
nor U13279 (N_13279,N_13023,N_13051);
and U13280 (N_13280,N_13053,N_13005);
nor U13281 (N_13281,N_13063,N_13029);
nand U13282 (N_13282,N_13108,N_13107);
xnor U13283 (N_13283,N_13079,N_13050);
nand U13284 (N_13284,N_13182,N_13085);
and U13285 (N_13285,N_13034,N_13104);
and U13286 (N_13286,N_13075,N_13041);
xnor U13287 (N_13287,N_13158,N_13092);
nand U13288 (N_13288,N_13156,N_13072);
nand U13289 (N_13289,N_13157,N_13179);
or U13290 (N_13290,N_13078,N_13185);
or U13291 (N_13291,N_13175,N_13056);
nor U13292 (N_13292,N_13139,N_13111);
nor U13293 (N_13293,N_13194,N_13189);
nor U13294 (N_13294,N_13125,N_13173);
nor U13295 (N_13295,N_13181,N_13100);
and U13296 (N_13296,N_13115,N_13028);
nor U13297 (N_13297,N_13134,N_13159);
nor U13298 (N_13298,N_13094,N_13172);
or U13299 (N_13299,N_13070,N_13020);
nand U13300 (N_13300,N_13136,N_13195);
nor U13301 (N_13301,N_13039,N_13197);
nor U13302 (N_13302,N_13086,N_13045);
xnor U13303 (N_13303,N_13061,N_13050);
nor U13304 (N_13304,N_13139,N_13196);
nand U13305 (N_13305,N_13093,N_13084);
nor U13306 (N_13306,N_13199,N_13040);
nor U13307 (N_13307,N_13047,N_13172);
nand U13308 (N_13308,N_13024,N_13188);
xor U13309 (N_13309,N_13043,N_13169);
nand U13310 (N_13310,N_13171,N_13110);
nor U13311 (N_13311,N_13134,N_13161);
xnor U13312 (N_13312,N_13119,N_13100);
and U13313 (N_13313,N_13046,N_13085);
nand U13314 (N_13314,N_13071,N_13130);
or U13315 (N_13315,N_13063,N_13124);
or U13316 (N_13316,N_13113,N_13114);
nor U13317 (N_13317,N_13028,N_13017);
nor U13318 (N_13318,N_13141,N_13151);
nor U13319 (N_13319,N_13105,N_13050);
nand U13320 (N_13320,N_13051,N_13041);
and U13321 (N_13321,N_13186,N_13120);
nor U13322 (N_13322,N_13016,N_13081);
or U13323 (N_13323,N_13109,N_13007);
xnor U13324 (N_13324,N_13114,N_13146);
nand U13325 (N_13325,N_13105,N_13113);
and U13326 (N_13326,N_13001,N_13158);
nand U13327 (N_13327,N_13161,N_13074);
xnor U13328 (N_13328,N_13034,N_13128);
nand U13329 (N_13329,N_13129,N_13028);
and U13330 (N_13330,N_13141,N_13025);
or U13331 (N_13331,N_13137,N_13121);
nor U13332 (N_13332,N_13116,N_13135);
or U13333 (N_13333,N_13035,N_13133);
nor U13334 (N_13334,N_13180,N_13149);
xor U13335 (N_13335,N_13004,N_13198);
and U13336 (N_13336,N_13118,N_13112);
nor U13337 (N_13337,N_13138,N_13103);
nor U13338 (N_13338,N_13029,N_13037);
or U13339 (N_13339,N_13060,N_13181);
xnor U13340 (N_13340,N_13026,N_13046);
nor U13341 (N_13341,N_13137,N_13136);
nand U13342 (N_13342,N_13189,N_13164);
nor U13343 (N_13343,N_13004,N_13062);
nand U13344 (N_13344,N_13100,N_13178);
nor U13345 (N_13345,N_13170,N_13177);
nor U13346 (N_13346,N_13069,N_13061);
xor U13347 (N_13347,N_13130,N_13147);
and U13348 (N_13348,N_13004,N_13039);
and U13349 (N_13349,N_13057,N_13075);
xor U13350 (N_13350,N_13003,N_13077);
and U13351 (N_13351,N_13071,N_13036);
xnor U13352 (N_13352,N_13017,N_13000);
nand U13353 (N_13353,N_13016,N_13002);
xor U13354 (N_13354,N_13135,N_13111);
and U13355 (N_13355,N_13159,N_13024);
or U13356 (N_13356,N_13185,N_13164);
nand U13357 (N_13357,N_13078,N_13137);
nand U13358 (N_13358,N_13096,N_13141);
xor U13359 (N_13359,N_13178,N_13038);
nand U13360 (N_13360,N_13010,N_13100);
and U13361 (N_13361,N_13194,N_13072);
nor U13362 (N_13362,N_13110,N_13041);
nor U13363 (N_13363,N_13033,N_13075);
and U13364 (N_13364,N_13165,N_13189);
and U13365 (N_13365,N_13077,N_13086);
and U13366 (N_13366,N_13094,N_13013);
xor U13367 (N_13367,N_13166,N_13021);
or U13368 (N_13368,N_13144,N_13027);
or U13369 (N_13369,N_13140,N_13173);
xor U13370 (N_13370,N_13080,N_13172);
and U13371 (N_13371,N_13026,N_13124);
or U13372 (N_13372,N_13169,N_13118);
nor U13373 (N_13373,N_13182,N_13031);
nor U13374 (N_13374,N_13040,N_13025);
and U13375 (N_13375,N_13181,N_13179);
xor U13376 (N_13376,N_13007,N_13176);
or U13377 (N_13377,N_13044,N_13094);
nand U13378 (N_13378,N_13159,N_13140);
nor U13379 (N_13379,N_13178,N_13196);
nor U13380 (N_13380,N_13022,N_13047);
nor U13381 (N_13381,N_13133,N_13026);
xor U13382 (N_13382,N_13169,N_13156);
nand U13383 (N_13383,N_13098,N_13106);
nor U13384 (N_13384,N_13148,N_13020);
xor U13385 (N_13385,N_13009,N_13063);
or U13386 (N_13386,N_13089,N_13177);
nand U13387 (N_13387,N_13197,N_13055);
nor U13388 (N_13388,N_13198,N_13005);
or U13389 (N_13389,N_13008,N_13160);
xor U13390 (N_13390,N_13104,N_13132);
nand U13391 (N_13391,N_13029,N_13114);
nor U13392 (N_13392,N_13190,N_13100);
xnor U13393 (N_13393,N_13111,N_13150);
nand U13394 (N_13394,N_13097,N_13144);
nand U13395 (N_13395,N_13112,N_13081);
xor U13396 (N_13396,N_13056,N_13006);
or U13397 (N_13397,N_13100,N_13136);
xor U13398 (N_13398,N_13039,N_13062);
nand U13399 (N_13399,N_13184,N_13166);
and U13400 (N_13400,N_13364,N_13282);
xor U13401 (N_13401,N_13226,N_13341);
and U13402 (N_13402,N_13200,N_13324);
nand U13403 (N_13403,N_13399,N_13307);
nor U13404 (N_13404,N_13333,N_13369);
xor U13405 (N_13405,N_13367,N_13280);
nor U13406 (N_13406,N_13394,N_13286);
xor U13407 (N_13407,N_13207,N_13291);
xor U13408 (N_13408,N_13326,N_13386);
nand U13409 (N_13409,N_13295,N_13330);
nor U13410 (N_13410,N_13398,N_13372);
or U13411 (N_13411,N_13297,N_13213);
nand U13412 (N_13412,N_13331,N_13285);
and U13413 (N_13413,N_13222,N_13340);
nor U13414 (N_13414,N_13262,N_13270);
or U13415 (N_13415,N_13377,N_13316);
or U13416 (N_13416,N_13206,N_13254);
and U13417 (N_13417,N_13352,N_13240);
and U13418 (N_13418,N_13313,N_13283);
or U13419 (N_13419,N_13247,N_13299);
nor U13420 (N_13420,N_13237,N_13265);
and U13421 (N_13421,N_13378,N_13217);
xor U13422 (N_13422,N_13231,N_13290);
or U13423 (N_13423,N_13312,N_13379);
xor U13424 (N_13424,N_13343,N_13298);
xor U13425 (N_13425,N_13355,N_13287);
xnor U13426 (N_13426,N_13245,N_13309);
nor U13427 (N_13427,N_13366,N_13246);
nor U13428 (N_13428,N_13278,N_13243);
nand U13429 (N_13429,N_13232,N_13274);
or U13430 (N_13430,N_13224,N_13203);
nor U13431 (N_13431,N_13396,N_13211);
xor U13432 (N_13432,N_13271,N_13362);
nand U13433 (N_13433,N_13381,N_13261);
or U13434 (N_13434,N_13393,N_13281);
nor U13435 (N_13435,N_13248,N_13300);
xnor U13436 (N_13436,N_13373,N_13337);
or U13437 (N_13437,N_13370,N_13269);
or U13438 (N_13438,N_13252,N_13277);
nand U13439 (N_13439,N_13392,N_13215);
and U13440 (N_13440,N_13253,N_13228);
xor U13441 (N_13441,N_13223,N_13360);
or U13442 (N_13442,N_13348,N_13250);
xor U13443 (N_13443,N_13389,N_13235);
and U13444 (N_13444,N_13391,N_13344);
or U13445 (N_13445,N_13242,N_13227);
and U13446 (N_13446,N_13305,N_13284);
or U13447 (N_13447,N_13259,N_13339);
or U13448 (N_13448,N_13332,N_13395);
xnor U13449 (N_13449,N_13202,N_13383);
and U13450 (N_13450,N_13201,N_13338);
nor U13451 (N_13451,N_13314,N_13325);
and U13452 (N_13452,N_13236,N_13329);
xnor U13453 (N_13453,N_13216,N_13288);
and U13454 (N_13454,N_13279,N_13327);
or U13455 (N_13455,N_13257,N_13251);
or U13456 (N_13456,N_13249,N_13268);
or U13457 (N_13457,N_13380,N_13342);
xnor U13458 (N_13458,N_13204,N_13276);
xor U13459 (N_13459,N_13365,N_13239);
and U13460 (N_13460,N_13371,N_13357);
or U13461 (N_13461,N_13230,N_13387);
and U13462 (N_13462,N_13345,N_13294);
and U13463 (N_13463,N_13384,N_13234);
or U13464 (N_13464,N_13349,N_13323);
xnor U13465 (N_13465,N_13205,N_13315);
or U13466 (N_13466,N_13221,N_13255);
nand U13467 (N_13467,N_13328,N_13210);
nand U13468 (N_13468,N_13318,N_13376);
nor U13469 (N_13469,N_13359,N_13354);
xnor U13470 (N_13470,N_13267,N_13351);
nand U13471 (N_13471,N_13302,N_13275);
and U13472 (N_13472,N_13320,N_13303);
xnor U13473 (N_13473,N_13310,N_13272);
xnor U13474 (N_13474,N_13289,N_13266);
or U13475 (N_13475,N_13397,N_13292);
or U13476 (N_13476,N_13220,N_13346);
xor U13477 (N_13477,N_13208,N_13212);
and U13478 (N_13478,N_13256,N_13263);
and U13479 (N_13479,N_13350,N_13321);
nand U13480 (N_13480,N_13363,N_13214);
and U13481 (N_13481,N_13336,N_13358);
nor U13482 (N_13482,N_13308,N_13317);
or U13483 (N_13483,N_13375,N_13382);
nand U13484 (N_13484,N_13306,N_13388);
or U13485 (N_13485,N_13385,N_13264);
nor U13486 (N_13486,N_13374,N_13335);
xor U13487 (N_13487,N_13296,N_13334);
or U13488 (N_13488,N_13260,N_13244);
or U13489 (N_13489,N_13311,N_13304);
nand U13490 (N_13490,N_13347,N_13238);
or U13491 (N_13491,N_13361,N_13368);
xor U13492 (N_13492,N_13233,N_13322);
or U13493 (N_13493,N_13229,N_13356);
or U13494 (N_13494,N_13218,N_13353);
nor U13495 (N_13495,N_13301,N_13273);
xnor U13496 (N_13496,N_13258,N_13209);
nand U13497 (N_13497,N_13241,N_13219);
nor U13498 (N_13498,N_13319,N_13293);
or U13499 (N_13499,N_13390,N_13225);
nor U13500 (N_13500,N_13304,N_13333);
nor U13501 (N_13501,N_13310,N_13301);
and U13502 (N_13502,N_13234,N_13351);
and U13503 (N_13503,N_13323,N_13249);
and U13504 (N_13504,N_13208,N_13331);
xnor U13505 (N_13505,N_13221,N_13262);
and U13506 (N_13506,N_13289,N_13393);
and U13507 (N_13507,N_13328,N_13277);
nand U13508 (N_13508,N_13232,N_13304);
nor U13509 (N_13509,N_13205,N_13313);
nor U13510 (N_13510,N_13308,N_13228);
xnor U13511 (N_13511,N_13204,N_13258);
or U13512 (N_13512,N_13377,N_13331);
nand U13513 (N_13513,N_13287,N_13341);
nand U13514 (N_13514,N_13208,N_13216);
xnor U13515 (N_13515,N_13392,N_13394);
xor U13516 (N_13516,N_13309,N_13275);
and U13517 (N_13517,N_13382,N_13371);
or U13518 (N_13518,N_13398,N_13350);
xnor U13519 (N_13519,N_13258,N_13329);
and U13520 (N_13520,N_13375,N_13370);
nor U13521 (N_13521,N_13366,N_13315);
xnor U13522 (N_13522,N_13248,N_13383);
or U13523 (N_13523,N_13384,N_13279);
or U13524 (N_13524,N_13306,N_13271);
and U13525 (N_13525,N_13201,N_13279);
and U13526 (N_13526,N_13327,N_13282);
and U13527 (N_13527,N_13232,N_13201);
nand U13528 (N_13528,N_13320,N_13226);
and U13529 (N_13529,N_13318,N_13389);
and U13530 (N_13530,N_13250,N_13253);
and U13531 (N_13531,N_13231,N_13274);
xnor U13532 (N_13532,N_13245,N_13344);
and U13533 (N_13533,N_13210,N_13221);
and U13534 (N_13534,N_13353,N_13268);
nand U13535 (N_13535,N_13281,N_13384);
nor U13536 (N_13536,N_13244,N_13347);
nor U13537 (N_13537,N_13278,N_13334);
nor U13538 (N_13538,N_13347,N_13202);
or U13539 (N_13539,N_13267,N_13314);
or U13540 (N_13540,N_13337,N_13202);
nand U13541 (N_13541,N_13376,N_13313);
xnor U13542 (N_13542,N_13266,N_13329);
nor U13543 (N_13543,N_13223,N_13365);
or U13544 (N_13544,N_13349,N_13240);
xnor U13545 (N_13545,N_13321,N_13233);
or U13546 (N_13546,N_13266,N_13263);
nand U13547 (N_13547,N_13261,N_13244);
nor U13548 (N_13548,N_13374,N_13212);
xor U13549 (N_13549,N_13344,N_13214);
nor U13550 (N_13550,N_13373,N_13360);
xnor U13551 (N_13551,N_13292,N_13374);
or U13552 (N_13552,N_13216,N_13287);
nor U13553 (N_13553,N_13204,N_13326);
nand U13554 (N_13554,N_13306,N_13314);
xnor U13555 (N_13555,N_13365,N_13337);
xor U13556 (N_13556,N_13301,N_13338);
and U13557 (N_13557,N_13388,N_13265);
and U13558 (N_13558,N_13280,N_13336);
and U13559 (N_13559,N_13336,N_13201);
nor U13560 (N_13560,N_13245,N_13392);
nand U13561 (N_13561,N_13367,N_13246);
or U13562 (N_13562,N_13361,N_13393);
nand U13563 (N_13563,N_13379,N_13200);
nor U13564 (N_13564,N_13343,N_13275);
or U13565 (N_13565,N_13290,N_13265);
nor U13566 (N_13566,N_13307,N_13330);
or U13567 (N_13567,N_13269,N_13355);
xor U13568 (N_13568,N_13220,N_13237);
xnor U13569 (N_13569,N_13234,N_13240);
nand U13570 (N_13570,N_13378,N_13313);
nand U13571 (N_13571,N_13291,N_13287);
nor U13572 (N_13572,N_13204,N_13228);
xor U13573 (N_13573,N_13272,N_13385);
nor U13574 (N_13574,N_13320,N_13213);
or U13575 (N_13575,N_13253,N_13230);
nand U13576 (N_13576,N_13388,N_13300);
and U13577 (N_13577,N_13227,N_13371);
or U13578 (N_13578,N_13213,N_13227);
nand U13579 (N_13579,N_13327,N_13261);
and U13580 (N_13580,N_13363,N_13381);
or U13581 (N_13581,N_13318,N_13370);
nand U13582 (N_13582,N_13389,N_13347);
or U13583 (N_13583,N_13363,N_13290);
and U13584 (N_13584,N_13263,N_13335);
and U13585 (N_13585,N_13240,N_13340);
and U13586 (N_13586,N_13357,N_13353);
nor U13587 (N_13587,N_13217,N_13342);
and U13588 (N_13588,N_13387,N_13288);
or U13589 (N_13589,N_13385,N_13360);
nand U13590 (N_13590,N_13349,N_13231);
or U13591 (N_13591,N_13340,N_13300);
or U13592 (N_13592,N_13310,N_13222);
or U13593 (N_13593,N_13384,N_13383);
and U13594 (N_13594,N_13209,N_13390);
nor U13595 (N_13595,N_13264,N_13215);
nor U13596 (N_13596,N_13274,N_13209);
nand U13597 (N_13597,N_13359,N_13207);
and U13598 (N_13598,N_13244,N_13323);
and U13599 (N_13599,N_13216,N_13266);
nand U13600 (N_13600,N_13555,N_13407);
nor U13601 (N_13601,N_13495,N_13422);
nor U13602 (N_13602,N_13503,N_13545);
xor U13603 (N_13603,N_13451,N_13448);
nor U13604 (N_13604,N_13530,N_13590);
nor U13605 (N_13605,N_13491,N_13426);
nor U13606 (N_13606,N_13476,N_13415);
xnor U13607 (N_13607,N_13431,N_13484);
or U13608 (N_13608,N_13570,N_13517);
nor U13609 (N_13609,N_13411,N_13583);
or U13610 (N_13610,N_13447,N_13443);
nor U13611 (N_13611,N_13487,N_13507);
or U13612 (N_13612,N_13474,N_13512);
xor U13613 (N_13613,N_13571,N_13598);
nand U13614 (N_13614,N_13592,N_13478);
nand U13615 (N_13615,N_13556,N_13542);
and U13616 (N_13616,N_13565,N_13466);
nand U13617 (N_13617,N_13524,N_13456);
or U13618 (N_13618,N_13505,N_13498);
xor U13619 (N_13619,N_13421,N_13471);
nor U13620 (N_13620,N_13497,N_13551);
nor U13621 (N_13621,N_13461,N_13467);
xor U13622 (N_13622,N_13549,N_13402);
nor U13623 (N_13623,N_13423,N_13409);
xor U13624 (N_13624,N_13435,N_13534);
or U13625 (N_13625,N_13532,N_13473);
nand U13626 (N_13626,N_13433,N_13404);
xor U13627 (N_13627,N_13541,N_13424);
and U13628 (N_13628,N_13574,N_13539);
xor U13629 (N_13629,N_13492,N_13531);
nor U13630 (N_13630,N_13501,N_13518);
nor U13631 (N_13631,N_13483,N_13405);
nor U13632 (N_13632,N_13526,N_13490);
and U13633 (N_13633,N_13416,N_13525);
xor U13634 (N_13634,N_13544,N_13579);
nor U13635 (N_13635,N_13504,N_13566);
xnor U13636 (N_13636,N_13464,N_13557);
nor U13637 (N_13637,N_13403,N_13414);
or U13638 (N_13638,N_13514,N_13516);
and U13639 (N_13639,N_13513,N_13442);
nor U13640 (N_13640,N_13477,N_13500);
nand U13641 (N_13641,N_13455,N_13536);
or U13642 (N_13642,N_13578,N_13577);
and U13643 (N_13643,N_13439,N_13520);
xnor U13644 (N_13644,N_13440,N_13538);
or U13645 (N_13645,N_13463,N_13521);
xor U13646 (N_13646,N_13420,N_13569);
and U13647 (N_13647,N_13596,N_13438);
nand U13648 (N_13648,N_13499,N_13564);
nor U13649 (N_13649,N_13417,N_13581);
and U13650 (N_13650,N_13535,N_13418);
and U13651 (N_13651,N_13591,N_13552);
nor U13652 (N_13652,N_13588,N_13462);
nand U13653 (N_13653,N_13595,N_13546);
and U13654 (N_13654,N_13468,N_13406);
and U13655 (N_13655,N_13509,N_13527);
xor U13656 (N_13656,N_13529,N_13446);
and U13657 (N_13657,N_13410,N_13472);
or U13658 (N_13658,N_13519,N_13401);
xnor U13659 (N_13659,N_13425,N_13568);
or U13660 (N_13660,N_13452,N_13515);
or U13661 (N_13661,N_13444,N_13599);
and U13662 (N_13662,N_13434,N_13413);
nor U13663 (N_13663,N_13528,N_13450);
nor U13664 (N_13664,N_13586,N_13482);
nand U13665 (N_13665,N_13475,N_13584);
xor U13666 (N_13666,N_13575,N_13589);
nand U13667 (N_13667,N_13585,N_13436);
xor U13668 (N_13668,N_13412,N_13465);
xor U13669 (N_13669,N_13453,N_13480);
and U13670 (N_13670,N_13562,N_13441);
or U13671 (N_13671,N_13428,N_13489);
nor U13672 (N_13672,N_13479,N_13563);
or U13673 (N_13673,N_13548,N_13594);
nor U13674 (N_13674,N_13537,N_13567);
xnor U13675 (N_13675,N_13430,N_13408);
and U13676 (N_13676,N_13488,N_13494);
nor U13677 (N_13677,N_13580,N_13511);
or U13678 (N_13678,N_13522,N_13496);
and U13679 (N_13679,N_13506,N_13470);
nand U13680 (N_13680,N_13427,N_13587);
or U13681 (N_13681,N_13540,N_13510);
nor U13682 (N_13682,N_13533,N_13432);
xnor U13683 (N_13683,N_13486,N_13508);
or U13684 (N_13684,N_13593,N_13553);
nand U13685 (N_13685,N_13576,N_13547);
and U13686 (N_13686,N_13429,N_13457);
xor U13687 (N_13687,N_13573,N_13419);
nor U13688 (N_13688,N_13481,N_13558);
xor U13689 (N_13689,N_13502,N_13459);
and U13690 (N_13690,N_13458,N_13572);
xnor U13691 (N_13691,N_13597,N_13460);
xor U13692 (N_13692,N_13469,N_13493);
or U13693 (N_13693,N_13559,N_13449);
or U13694 (N_13694,N_13554,N_13523);
and U13695 (N_13695,N_13437,N_13445);
xnor U13696 (N_13696,N_13550,N_13400);
nand U13697 (N_13697,N_13543,N_13582);
nand U13698 (N_13698,N_13561,N_13485);
nor U13699 (N_13699,N_13454,N_13560);
nor U13700 (N_13700,N_13468,N_13571);
or U13701 (N_13701,N_13416,N_13468);
nand U13702 (N_13702,N_13405,N_13436);
xnor U13703 (N_13703,N_13444,N_13431);
and U13704 (N_13704,N_13481,N_13408);
xor U13705 (N_13705,N_13529,N_13410);
or U13706 (N_13706,N_13597,N_13442);
xnor U13707 (N_13707,N_13491,N_13431);
nand U13708 (N_13708,N_13519,N_13548);
xor U13709 (N_13709,N_13589,N_13543);
and U13710 (N_13710,N_13446,N_13480);
and U13711 (N_13711,N_13430,N_13535);
nor U13712 (N_13712,N_13458,N_13477);
or U13713 (N_13713,N_13444,N_13557);
and U13714 (N_13714,N_13554,N_13518);
or U13715 (N_13715,N_13487,N_13445);
nand U13716 (N_13716,N_13592,N_13523);
nand U13717 (N_13717,N_13587,N_13542);
nor U13718 (N_13718,N_13496,N_13511);
nor U13719 (N_13719,N_13536,N_13460);
and U13720 (N_13720,N_13408,N_13571);
or U13721 (N_13721,N_13400,N_13593);
xor U13722 (N_13722,N_13470,N_13402);
xnor U13723 (N_13723,N_13437,N_13436);
or U13724 (N_13724,N_13563,N_13496);
xor U13725 (N_13725,N_13444,N_13570);
nor U13726 (N_13726,N_13522,N_13551);
nand U13727 (N_13727,N_13416,N_13404);
or U13728 (N_13728,N_13445,N_13457);
and U13729 (N_13729,N_13560,N_13475);
nand U13730 (N_13730,N_13586,N_13510);
nor U13731 (N_13731,N_13584,N_13482);
or U13732 (N_13732,N_13537,N_13500);
and U13733 (N_13733,N_13527,N_13463);
nand U13734 (N_13734,N_13463,N_13596);
nand U13735 (N_13735,N_13582,N_13448);
and U13736 (N_13736,N_13407,N_13533);
xnor U13737 (N_13737,N_13488,N_13570);
or U13738 (N_13738,N_13417,N_13598);
nand U13739 (N_13739,N_13483,N_13422);
nand U13740 (N_13740,N_13430,N_13559);
xor U13741 (N_13741,N_13469,N_13454);
xnor U13742 (N_13742,N_13549,N_13582);
xnor U13743 (N_13743,N_13513,N_13493);
nand U13744 (N_13744,N_13548,N_13552);
xor U13745 (N_13745,N_13503,N_13563);
or U13746 (N_13746,N_13513,N_13481);
and U13747 (N_13747,N_13462,N_13549);
nor U13748 (N_13748,N_13566,N_13429);
or U13749 (N_13749,N_13402,N_13557);
or U13750 (N_13750,N_13496,N_13452);
and U13751 (N_13751,N_13447,N_13502);
and U13752 (N_13752,N_13418,N_13452);
and U13753 (N_13753,N_13456,N_13483);
nand U13754 (N_13754,N_13498,N_13465);
xnor U13755 (N_13755,N_13436,N_13414);
and U13756 (N_13756,N_13508,N_13598);
nor U13757 (N_13757,N_13435,N_13403);
and U13758 (N_13758,N_13421,N_13417);
nor U13759 (N_13759,N_13548,N_13589);
nand U13760 (N_13760,N_13513,N_13408);
and U13761 (N_13761,N_13404,N_13420);
nor U13762 (N_13762,N_13578,N_13404);
nand U13763 (N_13763,N_13429,N_13517);
nor U13764 (N_13764,N_13516,N_13544);
xnor U13765 (N_13765,N_13415,N_13450);
nand U13766 (N_13766,N_13502,N_13501);
xor U13767 (N_13767,N_13401,N_13475);
or U13768 (N_13768,N_13511,N_13553);
nand U13769 (N_13769,N_13554,N_13504);
xnor U13770 (N_13770,N_13516,N_13546);
and U13771 (N_13771,N_13532,N_13537);
nor U13772 (N_13772,N_13510,N_13518);
or U13773 (N_13773,N_13427,N_13405);
xor U13774 (N_13774,N_13539,N_13497);
nand U13775 (N_13775,N_13417,N_13509);
xnor U13776 (N_13776,N_13595,N_13458);
nand U13777 (N_13777,N_13568,N_13520);
nor U13778 (N_13778,N_13481,N_13487);
or U13779 (N_13779,N_13546,N_13418);
nor U13780 (N_13780,N_13585,N_13402);
nand U13781 (N_13781,N_13518,N_13524);
or U13782 (N_13782,N_13530,N_13598);
or U13783 (N_13783,N_13488,N_13417);
and U13784 (N_13784,N_13476,N_13559);
nor U13785 (N_13785,N_13550,N_13575);
and U13786 (N_13786,N_13586,N_13556);
nor U13787 (N_13787,N_13557,N_13501);
xor U13788 (N_13788,N_13401,N_13585);
and U13789 (N_13789,N_13545,N_13460);
xor U13790 (N_13790,N_13420,N_13595);
nor U13791 (N_13791,N_13582,N_13596);
or U13792 (N_13792,N_13563,N_13560);
nand U13793 (N_13793,N_13465,N_13517);
or U13794 (N_13794,N_13462,N_13567);
or U13795 (N_13795,N_13551,N_13404);
xor U13796 (N_13796,N_13477,N_13542);
nor U13797 (N_13797,N_13555,N_13467);
nand U13798 (N_13798,N_13594,N_13523);
nor U13799 (N_13799,N_13555,N_13564);
xor U13800 (N_13800,N_13794,N_13692);
nand U13801 (N_13801,N_13660,N_13756);
nand U13802 (N_13802,N_13765,N_13787);
xor U13803 (N_13803,N_13704,N_13786);
nand U13804 (N_13804,N_13659,N_13623);
or U13805 (N_13805,N_13687,N_13754);
nand U13806 (N_13806,N_13686,N_13769);
xor U13807 (N_13807,N_13766,N_13797);
nand U13808 (N_13808,N_13682,N_13655);
or U13809 (N_13809,N_13725,N_13670);
nand U13810 (N_13810,N_13683,N_13711);
nand U13811 (N_13811,N_13770,N_13742);
nand U13812 (N_13812,N_13762,N_13796);
or U13813 (N_13813,N_13728,N_13701);
or U13814 (N_13814,N_13789,N_13689);
nand U13815 (N_13815,N_13740,N_13668);
xnor U13816 (N_13816,N_13696,N_13675);
nand U13817 (N_13817,N_13707,N_13680);
nor U13818 (N_13818,N_13662,N_13615);
nor U13819 (N_13819,N_13671,N_13705);
xor U13820 (N_13820,N_13674,N_13730);
nor U13821 (N_13821,N_13720,N_13753);
or U13822 (N_13822,N_13639,N_13643);
and U13823 (N_13823,N_13719,N_13798);
nand U13824 (N_13824,N_13637,N_13748);
nor U13825 (N_13825,N_13613,N_13635);
or U13826 (N_13826,N_13724,N_13758);
nand U13827 (N_13827,N_13644,N_13627);
nand U13828 (N_13828,N_13733,N_13774);
or U13829 (N_13829,N_13647,N_13710);
nor U13830 (N_13830,N_13784,N_13633);
and U13831 (N_13831,N_13661,N_13642);
and U13832 (N_13832,N_13792,N_13717);
nand U13833 (N_13833,N_13620,N_13630);
or U13834 (N_13834,N_13666,N_13695);
nand U13835 (N_13835,N_13614,N_13777);
and U13836 (N_13836,N_13743,N_13712);
nor U13837 (N_13837,N_13658,N_13793);
and U13838 (N_13838,N_13601,N_13732);
nor U13839 (N_13839,N_13773,N_13771);
nor U13840 (N_13840,N_13657,N_13638);
and U13841 (N_13841,N_13760,N_13678);
xor U13842 (N_13842,N_13763,N_13738);
or U13843 (N_13843,N_13757,N_13799);
nand U13844 (N_13844,N_13729,N_13772);
or U13845 (N_13845,N_13721,N_13636);
nand U13846 (N_13846,N_13782,N_13795);
and U13847 (N_13847,N_13788,N_13616);
or U13848 (N_13848,N_13746,N_13741);
xnor U13849 (N_13849,N_13649,N_13669);
nand U13850 (N_13850,N_13652,N_13656);
xnor U13851 (N_13851,N_13654,N_13681);
or U13852 (N_13852,N_13667,N_13673);
nand U13853 (N_13853,N_13735,N_13603);
nand U13854 (N_13854,N_13611,N_13672);
or U13855 (N_13855,N_13734,N_13684);
or U13856 (N_13856,N_13708,N_13628);
xor U13857 (N_13857,N_13602,N_13648);
nand U13858 (N_13858,N_13767,N_13755);
nand U13859 (N_13859,N_13731,N_13619);
nand U13860 (N_13860,N_13785,N_13706);
and U13861 (N_13861,N_13610,N_13700);
and U13862 (N_13862,N_13702,N_13718);
nand U13863 (N_13863,N_13749,N_13791);
nor U13864 (N_13864,N_13618,N_13607);
or U13865 (N_13865,N_13703,N_13750);
nor U13866 (N_13866,N_13641,N_13690);
xnor U13867 (N_13867,N_13715,N_13646);
xnor U13868 (N_13868,N_13693,N_13699);
or U13869 (N_13869,N_13676,N_13650);
nor U13870 (N_13870,N_13722,N_13775);
or U13871 (N_13871,N_13737,N_13698);
xnor U13872 (N_13872,N_13779,N_13752);
xor U13873 (N_13873,N_13697,N_13609);
or U13874 (N_13874,N_13679,N_13739);
xor U13875 (N_13875,N_13790,N_13745);
xor U13876 (N_13876,N_13626,N_13606);
nor U13877 (N_13877,N_13622,N_13694);
nand U13878 (N_13878,N_13600,N_13685);
and U13879 (N_13879,N_13640,N_13688);
nand U13880 (N_13880,N_13624,N_13629);
nor U13881 (N_13881,N_13713,N_13634);
nor U13882 (N_13882,N_13709,N_13612);
nor U13883 (N_13883,N_13723,N_13776);
nand U13884 (N_13884,N_13744,N_13605);
or U13885 (N_13885,N_13768,N_13691);
xnor U13886 (N_13886,N_13677,N_13663);
xnor U13887 (N_13887,N_13651,N_13604);
or U13888 (N_13888,N_13726,N_13747);
or U13889 (N_13889,N_13653,N_13714);
nor U13890 (N_13890,N_13664,N_13761);
nand U13891 (N_13891,N_13759,N_13665);
and U13892 (N_13892,N_13631,N_13645);
nand U13893 (N_13893,N_13625,N_13621);
xnor U13894 (N_13894,N_13608,N_13716);
or U13895 (N_13895,N_13736,N_13617);
nor U13896 (N_13896,N_13778,N_13764);
and U13897 (N_13897,N_13780,N_13632);
nand U13898 (N_13898,N_13751,N_13727);
nand U13899 (N_13899,N_13781,N_13783);
or U13900 (N_13900,N_13700,N_13678);
or U13901 (N_13901,N_13751,N_13654);
nor U13902 (N_13902,N_13756,N_13722);
xnor U13903 (N_13903,N_13684,N_13703);
xor U13904 (N_13904,N_13681,N_13712);
nor U13905 (N_13905,N_13703,N_13700);
xor U13906 (N_13906,N_13681,N_13732);
nand U13907 (N_13907,N_13639,N_13631);
nor U13908 (N_13908,N_13605,N_13644);
nand U13909 (N_13909,N_13772,N_13641);
nand U13910 (N_13910,N_13776,N_13771);
or U13911 (N_13911,N_13754,N_13792);
xor U13912 (N_13912,N_13737,N_13669);
or U13913 (N_13913,N_13757,N_13678);
nand U13914 (N_13914,N_13652,N_13701);
nand U13915 (N_13915,N_13611,N_13647);
or U13916 (N_13916,N_13704,N_13631);
xor U13917 (N_13917,N_13683,N_13742);
nor U13918 (N_13918,N_13747,N_13663);
or U13919 (N_13919,N_13679,N_13651);
xnor U13920 (N_13920,N_13609,N_13789);
nor U13921 (N_13921,N_13744,N_13713);
and U13922 (N_13922,N_13774,N_13779);
nand U13923 (N_13923,N_13795,N_13765);
and U13924 (N_13924,N_13753,N_13708);
nor U13925 (N_13925,N_13758,N_13717);
xor U13926 (N_13926,N_13675,N_13755);
nand U13927 (N_13927,N_13684,N_13683);
or U13928 (N_13928,N_13782,N_13648);
nand U13929 (N_13929,N_13740,N_13616);
nand U13930 (N_13930,N_13633,N_13641);
and U13931 (N_13931,N_13767,N_13731);
xor U13932 (N_13932,N_13700,N_13798);
nor U13933 (N_13933,N_13645,N_13754);
xnor U13934 (N_13934,N_13701,N_13761);
xor U13935 (N_13935,N_13619,N_13798);
xor U13936 (N_13936,N_13618,N_13600);
xor U13937 (N_13937,N_13724,N_13657);
or U13938 (N_13938,N_13711,N_13626);
nand U13939 (N_13939,N_13671,N_13716);
xor U13940 (N_13940,N_13719,N_13682);
and U13941 (N_13941,N_13694,N_13698);
nand U13942 (N_13942,N_13796,N_13709);
xnor U13943 (N_13943,N_13700,N_13708);
nor U13944 (N_13944,N_13755,N_13753);
or U13945 (N_13945,N_13779,N_13623);
nand U13946 (N_13946,N_13706,N_13759);
and U13947 (N_13947,N_13642,N_13732);
nor U13948 (N_13948,N_13702,N_13796);
and U13949 (N_13949,N_13654,N_13790);
xnor U13950 (N_13950,N_13792,N_13686);
and U13951 (N_13951,N_13644,N_13729);
and U13952 (N_13952,N_13738,N_13733);
nand U13953 (N_13953,N_13789,N_13625);
nand U13954 (N_13954,N_13685,N_13689);
or U13955 (N_13955,N_13723,N_13714);
or U13956 (N_13956,N_13618,N_13625);
nor U13957 (N_13957,N_13609,N_13665);
xor U13958 (N_13958,N_13740,N_13653);
nand U13959 (N_13959,N_13606,N_13781);
or U13960 (N_13960,N_13796,N_13729);
nor U13961 (N_13961,N_13608,N_13742);
nand U13962 (N_13962,N_13726,N_13745);
nand U13963 (N_13963,N_13675,N_13684);
xor U13964 (N_13964,N_13626,N_13740);
or U13965 (N_13965,N_13658,N_13683);
or U13966 (N_13966,N_13775,N_13693);
and U13967 (N_13967,N_13621,N_13755);
xor U13968 (N_13968,N_13635,N_13602);
and U13969 (N_13969,N_13602,N_13787);
nor U13970 (N_13970,N_13785,N_13724);
and U13971 (N_13971,N_13656,N_13627);
and U13972 (N_13972,N_13603,N_13639);
or U13973 (N_13973,N_13776,N_13778);
and U13974 (N_13974,N_13777,N_13604);
xnor U13975 (N_13975,N_13711,N_13677);
or U13976 (N_13976,N_13776,N_13775);
xnor U13977 (N_13977,N_13642,N_13641);
xor U13978 (N_13978,N_13784,N_13700);
or U13979 (N_13979,N_13624,N_13665);
and U13980 (N_13980,N_13689,N_13767);
nor U13981 (N_13981,N_13634,N_13798);
nor U13982 (N_13982,N_13712,N_13601);
and U13983 (N_13983,N_13641,N_13756);
nand U13984 (N_13984,N_13770,N_13666);
or U13985 (N_13985,N_13711,N_13740);
nor U13986 (N_13986,N_13700,N_13642);
and U13987 (N_13987,N_13730,N_13731);
and U13988 (N_13988,N_13671,N_13695);
nand U13989 (N_13989,N_13638,N_13755);
nor U13990 (N_13990,N_13626,N_13612);
nand U13991 (N_13991,N_13706,N_13750);
nand U13992 (N_13992,N_13617,N_13677);
or U13993 (N_13993,N_13707,N_13746);
nand U13994 (N_13994,N_13644,N_13664);
nand U13995 (N_13995,N_13739,N_13644);
or U13996 (N_13996,N_13653,N_13760);
xnor U13997 (N_13997,N_13771,N_13665);
nand U13998 (N_13998,N_13620,N_13711);
or U13999 (N_13999,N_13755,N_13610);
xnor U14000 (N_14000,N_13925,N_13881);
nor U14001 (N_14001,N_13937,N_13868);
nor U14002 (N_14002,N_13973,N_13869);
or U14003 (N_14003,N_13862,N_13900);
nand U14004 (N_14004,N_13980,N_13842);
nand U14005 (N_14005,N_13971,N_13995);
nor U14006 (N_14006,N_13871,N_13952);
and U14007 (N_14007,N_13891,N_13954);
and U14008 (N_14008,N_13944,N_13874);
xor U14009 (N_14009,N_13808,N_13837);
xnor U14010 (N_14010,N_13844,N_13846);
and U14011 (N_14011,N_13916,N_13850);
or U14012 (N_14012,N_13910,N_13929);
nor U14013 (N_14013,N_13974,N_13939);
xnor U14014 (N_14014,N_13807,N_13964);
xor U14015 (N_14015,N_13985,N_13813);
xnor U14016 (N_14016,N_13998,N_13911);
xnor U14017 (N_14017,N_13931,N_13854);
or U14018 (N_14018,N_13930,N_13986);
nand U14019 (N_14019,N_13924,N_13904);
nor U14020 (N_14020,N_13926,N_13969);
and U14021 (N_14021,N_13899,N_13901);
or U14022 (N_14022,N_13962,N_13981);
and U14023 (N_14023,N_13909,N_13913);
nand U14024 (N_14024,N_13912,N_13861);
xnor U14025 (N_14025,N_13923,N_13878);
or U14026 (N_14026,N_13920,N_13825);
and U14027 (N_14027,N_13997,N_13864);
nor U14028 (N_14028,N_13857,N_13801);
nor U14029 (N_14029,N_13953,N_13961);
and U14030 (N_14030,N_13814,N_13988);
nand U14031 (N_14031,N_13940,N_13826);
and U14032 (N_14032,N_13815,N_13840);
nor U14033 (N_14033,N_13992,N_13804);
nor U14034 (N_14034,N_13820,N_13938);
or U14035 (N_14035,N_13816,N_13963);
or U14036 (N_14036,N_13890,N_13976);
xnor U14037 (N_14037,N_13896,N_13841);
and U14038 (N_14038,N_13987,N_13927);
nor U14039 (N_14039,N_13918,N_13852);
xor U14040 (N_14040,N_13991,N_13893);
or U14041 (N_14041,N_13809,N_13829);
or U14042 (N_14042,N_13830,N_13897);
xor U14043 (N_14043,N_13977,N_13824);
nand U14044 (N_14044,N_13892,N_13875);
xnor U14045 (N_14045,N_13818,N_13999);
nand U14046 (N_14046,N_13903,N_13989);
nand U14047 (N_14047,N_13905,N_13888);
xor U14048 (N_14048,N_13873,N_13885);
nand U14049 (N_14049,N_13984,N_13955);
or U14050 (N_14050,N_13957,N_13908);
nand U14051 (N_14051,N_13928,N_13994);
nand U14052 (N_14052,N_13949,N_13956);
nand U14053 (N_14053,N_13835,N_13932);
or U14054 (N_14054,N_13884,N_13802);
nor U14055 (N_14055,N_13847,N_13979);
nand U14056 (N_14056,N_13823,N_13810);
nand U14057 (N_14057,N_13921,N_13860);
xor U14058 (N_14058,N_13948,N_13836);
nor U14059 (N_14059,N_13941,N_13880);
xor U14060 (N_14060,N_13831,N_13805);
nand U14061 (N_14061,N_13917,N_13883);
nand U14062 (N_14062,N_13855,N_13895);
xnor U14063 (N_14063,N_13817,N_13843);
nor U14064 (N_14064,N_13978,N_13922);
and U14065 (N_14065,N_13915,N_13993);
and U14066 (N_14066,N_13856,N_13959);
xnor U14067 (N_14067,N_13972,N_13828);
nand U14068 (N_14068,N_13967,N_13821);
xnor U14069 (N_14069,N_13966,N_13945);
xor U14070 (N_14070,N_13851,N_13943);
nand U14071 (N_14071,N_13919,N_13907);
xor U14072 (N_14072,N_13811,N_13866);
nor U14073 (N_14073,N_13849,N_13858);
or U14074 (N_14074,N_13902,N_13975);
nand U14075 (N_14075,N_13935,N_13845);
nor U14076 (N_14076,N_13872,N_13832);
xor U14077 (N_14077,N_13947,N_13936);
nand U14078 (N_14078,N_13886,N_13965);
nand U14079 (N_14079,N_13946,N_13838);
nor U14080 (N_14080,N_13803,N_13876);
xor U14081 (N_14081,N_13889,N_13834);
and U14082 (N_14082,N_13894,N_13882);
or U14083 (N_14083,N_13914,N_13827);
xnor U14084 (N_14084,N_13990,N_13839);
or U14085 (N_14085,N_13819,N_13867);
or U14086 (N_14086,N_13859,N_13870);
nand U14087 (N_14087,N_13887,N_13983);
nand U14088 (N_14088,N_13950,N_13933);
nor U14089 (N_14089,N_13934,N_13898);
and U14090 (N_14090,N_13958,N_13942);
nand U14091 (N_14091,N_13812,N_13970);
and U14092 (N_14092,N_13877,N_13960);
and U14093 (N_14093,N_13806,N_13982);
and U14094 (N_14094,N_13853,N_13879);
and U14095 (N_14095,N_13996,N_13863);
and U14096 (N_14096,N_13800,N_13906);
xnor U14097 (N_14097,N_13848,N_13968);
and U14098 (N_14098,N_13865,N_13833);
xnor U14099 (N_14099,N_13822,N_13951);
xor U14100 (N_14100,N_13869,N_13845);
or U14101 (N_14101,N_13940,N_13844);
and U14102 (N_14102,N_13814,N_13964);
xnor U14103 (N_14103,N_13852,N_13928);
xor U14104 (N_14104,N_13837,N_13941);
nor U14105 (N_14105,N_13953,N_13915);
nor U14106 (N_14106,N_13843,N_13942);
nand U14107 (N_14107,N_13899,N_13823);
xor U14108 (N_14108,N_13832,N_13984);
nand U14109 (N_14109,N_13978,N_13880);
nor U14110 (N_14110,N_13937,N_13957);
nand U14111 (N_14111,N_13893,N_13964);
or U14112 (N_14112,N_13902,N_13946);
nand U14113 (N_14113,N_13828,N_13832);
nor U14114 (N_14114,N_13839,N_13898);
xor U14115 (N_14115,N_13972,N_13804);
or U14116 (N_14116,N_13919,N_13868);
or U14117 (N_14117,N_13838,N_13913);
and U14118 (N_14118,N_13876,N_13952);
nand U14119 (N_14119,N_13826,N_13927);
or U14120 (N_14120,N_13957,N_13960);
nor U14121 (N_14121,N_13951,N_13825);
or U14122 (N_14122,N_13873,N_13961);
xnor U14123 (N_14123,N_13913,N_13991);
nor U14124 (N_14124,N_13853,N_13964);
nand U14125 (N_14125,N_13833,N_13915);
xor U14126 (N_14126,N_13998,N_13990);
nand U14127 (N_14127,N_13839,N_13979);
or U14128 (N_14128,N_13930,N_13914);
nor U14129 (N_14129,N_13878,N_13949);
or U14130 (N_14130,N_13830,N_13839);
nor U14131 (N_14131,N_13806,N_13897);
xor U14132 (N_14132,N_13934,N_13963);
and U14133 (N_14133,N_13954,N_13830);
nand U14134 (N_14134,N_13903,N_13889);
xnor U14135 (N_14135,N_13873,N_13990);
nor U14136 (N_14136,N_13982,N_13932);
nor U14137 (N_14137,N_13993,N_13828);
xnor U14138 (N_14138,N_13812,N_13848);
nor U14139 (N_14139,N_13809,N_13934);
nor U14140 (N_14140,N_13930,N_13849);
nand U14141 (N_14141,N_13843,N_13990);
xor U14142 (N_14142,N_13815,N_13913);
nor U14143 (N_14143,N_13874,N_13838);
nand U14144 (N_14144,N_13964,N_13833);
nor U14145 (N_14145,N_13804,N_13823);
nand U14146 (N_14146,N_13806,N_13816);
nor U14147 (N_14147,N_13928,N_13956);
or U14148 (N_14148,N_13877,N_13979);
xnor U14149 (N_14149,N_13933,N_13850);
xor U14150 (N_14150,N_13919,N_13897);
and U14151 (N_14151,N_13904,N_13898);
nor U14152 (N_14152,N_13961,N_13946);
nand U14153 (N_14153,N_13922,N_13857);
and U14154 (N_14154,N_13960,N_13870);
nor U14155 (N_14155,N_13854,N_13932);
xor U14156 (N_14156,N_13994,N_13946);
or U14157 (N_14157,N_13928,N_13995);
or U14158 (N_14158,N_13891,N_13907);
nor U14159 (N_14159,N_13843,N_13888);
nand U14160 (N_14160,N_13878,N_13912);
and U14161 (N_14161,N_13827,N_13904);
nand U14162 (N_14162,N_13801,N_13892);
and U14163 (N_14163,N_13810,N_13848);
xor U14164 (N_14164,N_13882,N_13968);
xnor U14165 (N_14165,N_13804,N_13908);
nor U14166 (N_14166,N_13849,N_13998);
nand U14167 (N_14167,N_13838,N_13903);
or U14168 (N_14168,N_13869,N_13834);
nor U14169 (N_14169,N_13977,N_13841);
nand U14170 (N_14170,N_13887,N_13938);
and U14171 (N_14171,N_13980,N_13949);
nor U14172 (N_14172,N_13808,N_13915);
or U14173 (N_14173,N_13861,N_13994);
xnor U14174 (N_14174,N_13852,N_13807);
xnor U14175 (N_14175,N_13819,N_13945);
nand U14176 (N_14176,N_13832,N_13926);
nor U14177 (N_14177,N_13826,N_13875);
nand U14178 (N_14178,N_13806,N_13878);
or U14179 (N_14179,N_13928,N_13889);
xnor U14180 (N_14180,N_13803,N_13859);
or U14181 (N_14181,N_13940,N_13935);
nand U14182 (N_14182,N_13808,N_13996);
nand U14183 (N_14183,N_13872,N_13845);
nand U14184 (N_14184,N_13839,N_13989);
or U14185 (N_14185,N_13804,N_13828);
nand U14186 (N_14186,N_13816,N_13958);
nor U14187 (N_14187,N_13995,N_13859);
nand U14188 (N_14188,N_13967,N_13896);
xnor U14189 (N_14189,N_13953,N_13918);
xor U14190 (N_14190,N_13819,N_13878);
nor U14191 (N_14191,N_13922,N_13822);
nand U14192 (N_14192,N_13975,N_13814);
xor U14193 (N_14193,N_13941,N_13963);
xnor U14194 (N_14194,N_13974,N_13994);
nor U14195 (N_14195,N_13856,N_13909);
nor U14196 (N_14196,N_13970,N_13800);
nor U14197 (N_14197,N_13879,N_13893);
xor U14198 (N_14198,N_13952,N_13986);
or U14199 (N_14199,N_13822,N_13886);
nand U14200 (N_14200,N_14125,N_14171);
xor U14201 (N_14201,N_14064,N_14118);
nor U14202 (N_14202,N_14043,N_14065);
xor U14203 (N_14203,N_14031,N_14109);
nor U14204 (N_14204,N_14158,N_14060);
nand U14205 (N_14205,N_14154,N_14101);
nor U14206 (N_14206,N_14067,N_14013);
and U14207 (N_14207,N_14046,N_14077);
and U14208 (N_14208,N_14147,N_14083);
nand U14209 (N_14209,N_14194,N_14198);
nor U14210 (N_14210,N_14135,N_14119);
and U14211 (N_14211,N_14032,N_14052);
xnor U14212 (N_14212,N_14112,N_14131);
nor U14213 (N_14213,N_14104,N_14170);
xnor U14214 (N_14214,N_14041,N_14011);
and U14215 (N_14215,N_14184,N_14076);
or U14216 (N_14216,N_14029,N_14102);
xor U14217 (N_14217,N_14062,N_14003);
nand U14218 (N_14218,N_14089,N_14163);
and U14219 (N_14219,N_14017,N_14074);
xnor U14220 (N_14220,N_14020,N_14082);
nand U14221 (N_14221,N_14040,N_14183);
nor U14222 (N_14222,N_14026,N_14001);
or U14223 (N_14223,N_14140,N_14116);
nor U14224 (N_14224,N_14162,N_14161);
nor U14225 (N_14225,N_14004,N_14189);
nor U14226 (N_14226,N_14037,N_14096);
nor U14227 (N_14227,N_14137,N_14010);
and U14228 (N_14228,N_14055,N_14128);
or U14229 (N_14229,N_14008,N_14036);
xor U14230 (N_14230,N_14053,N_14068);
xnor U14231 (N_14231,N_14092,N_14034);
xnor U14232 (N_14232,N_14193,N_14059);
xnor U14233 (N_14233,N_14000,N_14025);
nor U14234 (N_14234,N_14054,N_14009);
or U14235 (N_14235,N_14091,N_14002);
nand U14236 (N_14236,N_14038,N_14063);
or U14237 (N_14237,N_14132,N_14190);
or U14238 (N_14238,N_14093,N_14086);
or U14239 (N_14239,N_14196,N_14103);
or U14240 (N_14240,N_14151,N_14022);
nor U14241 (N_14241,N_14095,N_14061);
nor U14242 (N_14242,N_14129,N_14106);
or U14243 (N_14243,N_14182,N_14006);
nand U14244 (N_14244,N_14090,N_14085);
or U14245 (N_14245,N_14072,N_14197);
nor U14246 (N_14246,N_14152,N_14175);
and U14247 (N_14247,N_14172,N_14153);
nor U14248 (N_14248,N_14111,N_14127);
and U14249 (N_14249,N_14039,N_14117);
and U14250 (N_14250,N_14097,N_14018);
xnor U14251 (N_14251,N_14051,N_14113);
xnor U14252 (N_14252,N_14044,N_14126);
nor U14253 (N_14253,N_14148,N_14110);
nor U14254 (N_14254,N_14150,N_14179);
nor U14255 (N_14255,N_14075,N_14165);
or U14256 (N_14256,N_14045,N_14167);
nor U14257 (N_14257,N_14164,N_14049);
or U14258 (N_14258,N_14199,N_14159);
xor U14259 (N_14259,N_14176,N_14073);
and U14260 (N_14260,N_14007,N_14107);
nand U14261 (N_14261,N_14160,N_14035);
and U14262 (N_14262,N_14155,N_14069);
nor U14263 (N_14263,N_14138,N_14005);
nor U14264 (N_14264,N_14122,N_14174);
and U14265 (N_14265,N_14188,N_14178);
xor U14266 (N_14266,N_14195,N_14185);
xnor U14267 (N_14267,N_14180,N_14187);
and U14268 (N_14268,N_14169,N_14120);
nor U14269 (N_14269,N_14057,N_14166);
nand U14270 (N_14270,N_14136,N_14094);
nor U14271 (N_14271,N_14100,N_14149);
xor U14272 (N_14272,N_14115,N_14181);
nor U14273 (N_14273,N_14177,N_14014);
nand U14274 (N_14274,N_14134,N_14133);
xnor U14275 (N_14275,N_14144,N_14078);
nor U14276 (N_14276,N_14123,N_14081);
xnor U14277 (N_14277,N_14056,N_14050);
nor U14278 (N_14278,N_14087,N_14030);
nor U14279 (N_14279,N_14124,N_14156);
nand U14280 (N_14280,N_14173,N_14191);
xnor U14281 (N_14281,N_14157,N_14024);
nand U14282 (N_14282,N_14021,N_14027);
nand U14283 (N_14283,N_14042,N_14088);
nand U14284 (N_14284,N_14105,N_14058);
xor U14285 (N_14285,N_14066,N_14186);
xnor U14286 (N_14286,N_14070,N_14012);
xor U14287 (N_14287,N_14192,N_14080);
nor U14288 (N_14288,N_14084,N_14028);
nand U14289 (N_14289,N_14019,N_14130);
and U14290 (N_14290,N_14047,N_14071);
and U14291 (N_14291,N_14048,N_14098);
or U14292 (N_14292,N_14015,N_14139);
nand U14293 (N_14293,N_14121,N_14079);
xnor U14294 (N_14294,N_14146,N_14141);
and U14295 (N_14295,N_14114,N_14145);
and U14296 (N_14296,N_14143,N_14033);
and U14297 (N_14297,N_14099,N_14168);
and U14298 (N_14298,N_14016,N_14108);
nand U14299 (N_14299,N_14023,N_14142);
and U14300 (N_14300,N_14049,N_14078);
nor U14301 (N_14301,N_14138,N_14148);
nand U14302 (N_14302,N_14071,N_14033);
xor U14303 (N_14303,N_14086,N_14036);
or U14304 (N_14304,N_14133,N_14131);
and U14305 (N_14305,N_14100,N_14154);
nor U14306 (N_14306,N_14151,N_14190);
or U14307 (N_14307,N_14108,N_14167);
and U14308 (N_14308,N_14082,N_14083);
nand U14309 (N_14309,N_14179,N_14076);
and U14310 (N_14310,N_14081,N_14016);
nand U14311 (N_14311,N_14042,N_14174);
nor U14312 (N_14312,N_14156,N_14192);
nand U14313 (N_14313,N_14006,N_14102);
xor U14314 (N_14314,N_14143,N_14010);
nor U14315 (N_14315,N_14180,N_14163);
nor U14316 (N_14316,N_14037,N_14084);
nand U14317 (N_14317,N_14180,N_14067);
and U14318 (N_14318,N_14157,N_14096);
and U14319 (N_14319,N_14029,N_14168);
xnor U14320 (N_14320,N_14055,N_14092);
or U14321 (N_14321,N_14059,N_14105);
and U14322 (N_14322,N_14161,N_14154);
nand U14323 (N_14323,N_14068,N_14137);
xor U14324 (N_14324,N_14063,N_14181);
xor U14325 (N_14325,N_14160,N_14188);
nor U14326 (N_14326,N_14029,N_14101);
nand U14327 (N_14327,N_14064,N_14173);
and U14328 (N_14328,N_14161,N_14160);
and U14329 (N_14329,N_14027,N_14064);
or U14330 (N_14330,N_14137,N_14065);
or U14331 (N_14331,N_14016,N_14122);
and U14332 (N_14332,N_14046,N_14089);
xnor U14333 (N_14333,N_14077,N_14168);
and U14334 (N_14334,N_14038,N_14097);
nor U14335 (N_14335,N_14111,N_14021);
xnor U14336 (N_14336,N_14070,N_14175);
and U14337 (N_14337,N_14007,N_14172);
nand U14338 (N_14338,N_14010,N_14083);
nor U14339 (N_14339,N_14145,N_14102);
nand U14340 (N_14340,N_14065,N_14179);
nand U14341 (N_14341,N_14185,N_14104);
nor U14342 (N_14342,N_14095,N_14069);
or U14343 (N_14343,N_14159,N_14106);
xor U14344 (N_14344,N_14199,N_14007);
or U14345 (N_14345,N_14190,N_14178);
or U14346 (N_14346,N_14190,N_14140);
or U14347 (N_14347,N_14025,N_14053);
nand U14348 (N_14348,N_14058,N_14167);
and U14349 (N_14349,N_14144,N_14121);
or U14350 (N_14350,N_14072,N_14005);
nor U14351 (N_14351,N_14038,N_14159);
nor U14352 (N_14352,N_14134,N_14126);
nor U14353 (N_14353,N_14043,N_14150);
nor U14354 (N_14354,N_14144,N_14183);
nand U14355 (N_14355,N_14069,N_14068);
xnor U14356 (N_14356,N_14082,N_14157);
or U14357 (N_14357,N_14149,N_14198);
or U14358 (N_14358,N_14071,N_14127);
and U14359 (N_14359,N_14096,N_14182);
xnor U14360 (N_14360,N_14008,N_14045);
or U14361 (N_14361,N_14104,N_14065);
nand U14362 (N_14362,N_14119,N_14004);
xnor U14363 (N_14363,N_14037,N_14017);
and U14364 (N_14364,N_14026,N_14040);
nor U14365 (N_14365,N_14088,N_14107);
or U14366 (N_14366,N_14128,N_14111);
nor U14367 (N_14367,N_14038,N_14020);
or U14368 (N_14368,N_14136,N_14134);
nor U14369 (N_14369,N_14142,N_14053);
or U14370 (N_14370,N_14093,N_14049);
xor U14371 (N_14371,N_14169,N_14187);
or U14372 (N_14372,N_14003,N_14011);
and U14373 (N_14373,N_14168,N_14011);
nand U14374 (N_14374,N_14045,N_14102);
or U14375 (N_14375,N_14045,N_14186);
xor U14376 (N_14376,N_14133,N_14142);
nand U14377 (N_14377,N_14058,N_14022);
xor U14378 (N_14378,N_14175,N_14083);
or U14379 (N_14379,N_14186,N_14077);
xnor U14380 (N_14380,N_14096,N_14171);
or U14381 (N_14381,N_14146,N_14178);
nor U14382 (N_14382,N_14180,N_14125);
xor U14383 (N_14383,N_14195,N_14125);
nor U14384 (N_14384,N_14090,N_14180);
nor U14385 (N_14385,N_14125,N_14122);
xor U14386 (N_14386,N_14143,N_14030);
xor U14387 (N_14387,N_14002,N_14101);
or U14388 (N_14388,N_14199,N_14171);
and U14389 (N_14389,N_14149,N_14114);
and U14390 (N_14390,N_14022,N_14008);
nand U14391 (N_14391,N_14057,N_14168);
nor U14392 (N_14392,N_14191,N_14076);
xnor U14393 (N_14393,N_14179,N_14121);
or U14394 (N_14394,N_14168,N_14178);
or U14395 (N_14395,N_14150,N_14101);
xnor U14396 (N_14396,N_14103,N_14101);
nor U14397 (N_14397,N_14030,N_14129);
nor U14398 (N_14398,N_14019,N_14165);
nand U14399 (N_14399,N_14086,N_14101);
and U14400 (N_14400,N_14296,N_14212);
or U14401 (N_14401,N_14289,N_14259);
xor U14402 (N_14402,N_14325,N_14365);
and U14403 (N_14403,N_14266,N_14388);
nand U14404 (N_14404,N_14341,N_14260);
or U14405 (N_14405,N_14337,N_14340);
nand U14406 (N_14406,N_14338,N_14243);
and U14407 (N_14407,N_14369,N_14330);
or U14408 (N_14408,N_14229,N_14327);
xnor U14409 (N_14409,N_14252,N_14247);
xnor U14410 (N_14410,N_14233,N_14262);
and U14411 (N_14411,N_14227,N_14223);
and U14412 (N_14412,N_14258,N_14257);
or U14413 (N_14413,N_14274,N_14367);
nor U14414 (N_14414,N_14228,N_14348);
nor U14415 (N_14415,N_14333,N_14209);
or U14416 (N_14416,N_14372,N_14214);
nand U14417 (N_14417,N_14270,N_14271);
or U14418 (N_14418,N_14359,N_14235);
nand U14419 (N_14419,N_14349,N_14332);
and U14420 (N_14420,N_14217,N_14383);
nor U14421 (N_14421,N_14384,N_14371);
xor U14422 (N_14422,N_14215,N_14208);
nor U14423 (N_14423,N_14292,N_14336);
and U14424 (N_14424,N_14361,N_14297);
nand U14425 (N_14425,N_14353,N_14393);
nand U14426 (N_14426,N_14366,N_14385);
nand U14427 (N_14427,N_14310,N_14394);
and U14428 (N_14428,N_14277,N_14392);
nor U14429 (N_14429,N_14350,N_14263);
xnor U14430 (N_14430,N_14304,N_14397);
nand U14431 (N_14431,N_14313,N_14302);
and U14432 (N_14432,N_14276,N_14249);
nand U14433 (N_14433,N_14379,N_14205);
and U14434 (N_14434,N_14275,N_14246);
nor U14435 (N_14435,N_14354,N_14206);
xor U14436 (N_14436,N_14295,N_14202);
nand U14437 (N_14437,N_14281,N_14334);
xnor U14438 (N_14438,N_14375,N_14381);
xor U14439 (N_14439,N_14207,N_14343);
or U14440 (N_14440,N_14329,N_14219);
or U14441 (N_14441,N_14244,N_14387);
nor U14442 (N_14442,N_14299,N_14237);
nand U14443 (N_14443,N_14267,N_14238);
and U14444 (N_14444,N_14374,N_14324);
or U14445 (N_14445,N_14222,N_14314);
xnor U14446 (N_14446,N_14345,N_14294);
nand U14447 (N_14447,N_14323,N_14358);
or U14448 (N_14448,N_14328,N_14288);
nand U14449 (N_14449,N_14278,N_14390);
or U14450 (N_14450,N_14220,N_14221);
nor U14451 (N_14451,N_14355,N_14253);
xnor U14452 (N_14452,N_14380,N_14261);
and U14453 (N_14453,N_14396,N_14320);
or U14454 (N_14454,N_14346,N_14268);
xor U14455 (N_14455,N_14342,N_14357);
or U14456 (N_14456,N_14315,N_14290);
and U14457 (N_14457,N_14286,N_14213);
xnor U14458 (N_14458,N_14264,N_14285);
and U14459 (N_14459,N_14232,N_14225);
and U14460 (N_14460,N_14256,N_14200);
nand U14461 (N_14461,N_14210,N_14382);
nor U14462 (N_14462,N_14203,N_14368);
xnor U14463 (N_14463,N_14298,N_14318);
nor U14464 (N_14464,N_14224,N_14201);
xor U14465 (N_14465,N_14360,N_14326);
and U14466 (N_14466,N_14245,N_14284);
nand U14467 (N_14467,N_14236,N_14347);
xor U14468 (N_14468,N_14306,N_14226);
nor U14469 (N_14469,N_14352,N_14216);
nand U14470 (N_14470,N_14335,N_14398);
nor U14471 (N_14471,N_14287,N_14218);
xnor U14472 (N_14472,N_14364,N_14311);
nor U14473 (N_14473,N_14362,N_14282);
and U14474 (N_14474,N_14242,N_14377);
nand U14475 (N_14475,N_14240,N_14250);
or U14476 (N_14476,N_14331,N_14269);
nor U14477 (N_14477,N_14312,N_14351);
xnor U14478 (N_14478,N_14303,N_14376);
nor U14479 (N_14479,N_14251,N_14378);
nand U14480 (N_14480,N_14309,N_14265);
and U14481 (N_14481,N_14280,N_14273);
or U14482 (N_14482,N_14399,N_14321);
and U14483 (N_14483,N_14344,N_14241);
and U14484 (N_14484,N_14254,N_14317);
nor U14485 (N_14485,N_14395,N_14293);
nand U14486 (N_14486,N_14356,N_14231);
nor U14487 (N_14487,N_14230,N_14291);
nand U14488 (N_14488,N_14248,N_14389);
nand U14489 (N_14489,N_14322,N_14204);
nand U14490 (N_14490,N_14373,N_14279);
nand U14491 (N_14491,N_14255,N_14386);
nor U14492 (N_14492,N_14391,N_14319);
and U14493 (N_14493,N_14339,N_14316);
nand U14494 (N_14494,N_14283,N_14305);
xor U14495 (N_14495,N_14307,N_14300);
or U14496 (N_14496,N_14301,N_14272);
nor U14497 (N_14497,N_14239,N_14363);
nor U14498 (N_14498,N_14308,N_14234);
nand U14499 (N_14499,N_14370,N_14211);
xnor U14500 (N_14500,N_14370,N_14272);
and U14501 (N_14501,N_14352,N_14277);
nand U14502 (N_14502,N_14329,N_14328);
xor U14503 (N_14503,N_14205,N_14305);
nor U14504 (N_14504,N_14223,N_14234);
nor U14505 (N_14505,N_14333,N_14256);
nand U14506 (N_14506,N_14252,N_14212);
xnor U14507 (N_14507,N_14293,N_14375);
xnor U14508 (N_14508,N_14298,N_14225);
nor U14509 (N_14509,N_14260,N_14287);
and U14510 (N_14510,N_14204,N_14216);
nor U14511 (N_14511,N_14202,N_14215);
or U14512 (N_14512,N_14267,N_14317);
nor U14513 (N_14513,N_14216,N_14208);
xnor U14514 (N_14514,N_14278,N_14389);
and U14515 (N_14515,N_14358,N_14278);
nor U14516 (N_14516,N_14206,N_14213);
and U14517 (N_14517,N_14375,N_14291);
or U14518 (N_14518,N_14362,N_14260);
nand U14519 (N_14519,N_14284,N_14273);
and U14520 (N_14520,N_14212,N_14214);
nor U14521 (N_14521,N_14222,N_14383);
and U14522 (N_14522,N_14376,N_14338);
nor U14523 (N_14523,N_14233,N_14283);
or U14524 (N_14524,N_14346,N_14340);
xor U14525 (N_14525,N_14344,N_14310);
or U14526 (N_14526,N_14295,N_14318);
xnor U14527 (N_14527,N_14396,N_14241);
nor U14528 (N_14528,N_14308,N_14259);
nor U14529 (N_14529,N_14294,N_14339);
nand U14530 (N_14530,N_14301,N_14375);
nand U14531 (N_14531,N_14237,N_14371);
or U14532 (N_14532,N_14360,N_14316);
nor U14533 (N_14533,N_14356,N_14340);
nand U14534 (N_14534,N_14300,N_14312);
or U14535 (N_14535,N_14330,N_14255);
and U14536 (N_14536,N_14374,N_14271);
nand U14537 (N_14537,N_14221,N_14261);
nand U14538 (N_14538,N_14356,N_14234);
nor U14539 (N_14539,N_14295,N_14375);
nand U14540 (N_14540,N_14282,N_14252);
nand U14541 (N_14541,N_14283,N_14280);
nor U14542 (N_14542,N_14250,N_14201);
nor U14543 (N_14543,N_14350,N_14277);
or U14544 (N_14544,N_14283,N_14321);
xnor U14545 (N_14545,N_14253,N_14394);
xnor U14546 (N_14546,N_14359,N_14361);
or U14547 (N_14547,N_14205,N_14299);
xnor U14548 (N_14548,N_14213,N_14244);
nand U14549 (N_14549,N_14266,N_14354);
and U14550 (N_14550,N_14387,N_14261);
xnor U14551 (N_14551,N_14271,N_14301);
xor U14552 (N_14552,N_14239,N_14355);
nand U14553 (N_14553,N_14295,N_14377);
nand U14554 (N_14554,N_14263,N_14204);
nor U14555 (N_14555,N_14329,N_14341);
and U14556 (N_14556,N_14206,N_14357);
or U14557 (N_14557,N_14251,N_14345);
xor U14558 (N_14558,N_14248,N_14352);
nand U14559 (N_14559,N_14244,N_14272);
or U14560 (N_14560,N_14329,N_14267);
nor U14561 (N_14561,N_14399,N_14328);
xor U14562 (N_14562,N_14320,N_14347);
nor U14563 (N_14563,N_14352,N_14398);
or U14564 (N_14564,N_14365,N_14310);
and U14565 (N_14565,N_14385,N_14331);
nor U14566 (N_14566,N_14388,N_14379);
or U14567 (N_14567,N_14308,N_14232);
and U14568 (N_14568,N_14247,N_14298);
nor U14569 (N_14569,N_14373,N_14290);
or U14570 (N_14570,N_14262,N_14368);
and U14571 (N_14571,N_14210,N_14290);
xnor U14572 (N_14572,N_14214,N_14306);
nand U14573 (N_14573,N_14290,N_14240);
nor U14574 (N_14574,N_14260,N_14241);
xor U14575 (N_14575,N_14277,N_14289);
nand U14576 (N_14576,N_14306,N_14321);
nor U14577 (N_14577,N_14380,N_14329);
xor U14578 (N_14578,N_14399,N_14357);
or U14579 (N_14579,N_14226,N_14341);
or U14580 (N_14580,N_14215,N_14276);
and U14581 (N_14581,N_14275,N_14257);
xnor U14582 (N_14582,N_14284,N_14399);
nand U14583 (N_14583,N_14370,N_14395);
xnor U14584 (N_14584,N_14254,N_14276);
nor U14585 (N_14585,N_14285,N_14376);
nand U14586 (N_14586,N_14276,N_14333);
or U14587 (N_14587,N_14249,N_14365);
and U14588 (N_14588,N_14226,N_14272);
nor U14589 (N_14589,N_14294,N_14379);
or U14590 (N_14590,N_14331,N_14250);
and U14591 (N_14591,N_14203,N_14249);
xnor U14592 (N_14592,N_14229,N_14233);
nand U14593 (N_14593,N_14358,N_14271);
and U14594 (N_14594,N_14351,N_14241);
or U14595 (N_14595,N_14383,N_14211);
and U14596 (N_14596,N_14373,N_14357);
nand U14597 (N_14597,N_14232,N_14222);
and U14598 (N_14598,N_14259,N_14316);
xor U14599 (N_14599,N_14364,N_14234);
nor U14600 (N_14600,N_14537,N_14539);
and U14601 (N_14601,N_14513,N_14594);
or U14602 (N_14602,N_14545,N_14592);
and U14603 (N_14603,N_14487,N_14588);
nor U14604 (N_14604,N_14485,N_14428);
xnor U14605 (N_14605,N_14526,N_14480);
or U14606 (N_14606,N_14585,N_14484);
or U14607 (N_14607,N_14430,N_14549);
and U14608 (N_14608,N_14451,N_14449);
and U14609 (N_14609,N_14412,N_14503);
nor U14610 (N_14610,N_14577,N_14536);
xor U14611 (N_14611,N_14534,N_14597);
xor U14612 (N_14612,N_14595,N_14570);
xnor U14613 (N_14613,N_14574,N_14510);
or U14614 (N_14614,N_14550,N_14483);
xnor U14615 (N_14615,N_14524,N_14468);
xor U14616 (N_14616,N_14509,N_14414);
or U14617 (N_14617,N_14421,N_14425);
or U14618 (N_14618,N_14482,N_14472);
nor U14619 (N_14619,N_14532,N_14481);
xnor U14620 (N_14620,N_14411,N_14465);
nand U14621 (N_14621,N_14567,N_14471);
xor U14622 (N_14622,N_14438,N_14402);
and U14623 (N_14623,N_14488,N_14562);
and U14624 (N_14624,N_14456,N_14401);
xnor U14625 (N_14625,N_14533,N_14467);
nor U14626 (N_14626,N_14400,N_14464);
nand U14627 (N_14627,N_14437,N_14598);
nor U14628 (N_14628,N_14500,N_14419);
or U14629 (N_14629,N_14426,N_14543);
xor U14630 (N_14630,N_14552,N_14590);
or U14631 (N_14631,N_14554,N_14440);
nor U14632 (N_14632,N_14519,N_14409);
or U14633 (N_14633,N_14501,N_14442);
nand U14634 (N_14634,N_14593,N_14494);
and U14635 (N_14635,N_14457,N_14497);
nand U14636 (N_14636,N_14455,N_14436);
nor U14637 (N_14637,N_14478,N_14517);
or U14638 (N_14638,N_14568,N_14529);
xnor U14639 (N_14639,N_14518,N_14540);
and U14640 (N_14640,N_14558,N_14572);
nor U14641 (N_14641,N_14427,N_14406);
xnor U14642 (N_14642,N_14542,N_14466);
nand U14643 (N_14643,N_14523,N_14458);
xnor U14644 (N_14644,N_14499,N_14505);
and U14645 (N_14645,N_14564,N_14506);
and U14646 (N_14646,N_14424,N_14553);
nand U14647 (N_14647,N_14420,N_14565);
xor U14648 (N_14648,N_14535,N_14515);
or U14649 (N_14649,N_14528,N_14446);
xor U14650 (N_14650,N_14569,N_14418);
or U14651 (N_14651,N_14511,N_14447);
or U14652 (N_14652,N_14559,N_14434);
nor U14653 (N_14653,N_14495,N_14583);
nor U14654 (N_14654,N_14450,N_14561);
xor U14655 (N_14655,N_14514,N_14453);
and U14656 (N_14656,N_14445,N_14433);
or U14657 (N_14657,N_14498,N_14454);
or U14658 (N_14658,N_14448,N_14582);
and U14659 (N_14659,N_14435,N_14573);
xor U14660 (N_14660,N_14462,N_14596);
xnor U14661 (N_14661,N_14416,N_14516);
nand U14662 (N_14662,N_14473,N_14551);
and U14663 (N_14663,N_14492,N_14439);
nand U14664 (N_14664,N_14520,N_14555);
nand U14665 (N_14665,N_14566,N_14407);
xnor U14666 (N_14666,N_14415,N_14504);
nor U14667 (N_14667,N_14479,N_14544);
or U14668 (N_14668,N_14474,N_14486);
or U14669 (N_14669,N_14563,N_14452);
and U14670 (N_14670,N_14477,N_14441);
xor U14671 (N_14671,N_14429,N_14548);
and U14672 (N_14672,N_14591,N_14489);
nand U14673 (N_14673,N_14413,N_14493);
xnor U14674 (N_14674,N_14538,N_14576);
nor U14675 (N_14675,N_14580,N_14512);
and U14676 (N_14676,N_14417,N_14490);
and U14677 (N_14677,N_14475,N_14422);
or U14678 (N_14678,N_14546,N_14470);
nor U14679 (N_14679,N_14507,N_14404);
and U14680 (N_14680,N_14599,N_14541);
nand U14681 (N_14681,N_14530,N_14423);
nand U14682 (N_14682,N_14431,N_14589);
and U14683 (N_14683,N_14579,N_14586);
nor U14684 (N_14684,N_14432,N_14531);
nand U14685 (N_14685,N_14496,N_14557);
nand U14686 (N_14686,N_14581,N_14578);
nor U14687 (N_14687,N_14461,N_14410);
xor U14688 (N_14688,N_14491,N_14476);
and U14689 (N_14689,N_14460,N_14527);
xnor U14690 (N_14690,N_14408,N_14459);
xor U14691 (N_14691,N_14571,N_14522);
nand U14692 (N_14692,N_14525,N_14443);
nand U14693 (N_14693,N_14584,N_14403);
nor U14694 (N_14694,N_14521,N_14444);
and U14695 (N_14695,N_14508,N_14469);
nand U14696 (N_14696,N_14587,N_14556);
xor U14697 (N_14697,N_14502,N_14560);
xor U14698 (N_14698,N_14575,N_14547);
nand U14699 (N_14699,N_14463,N_14405);
xnor U14700 (N_14700,N_14599,N_14516);
xnor U14701 (N_14701,N_14409,N_14423);
or U14702 (N_14702,N_14541,N_14565);
nand U14703 (N_14703,N_14541,N_14455);
nand U14704 (N_14704,N_14483,N_14447);
or U14705 (N_14705,N_14595,N_14505);
nor U14706 (N_14706,N_14546,N_14441);
nor U14707 (N_14707,N_14512,N_14414);
or U14708 (N_14708,N_14511,N_14524);
or U14709 (N_14709,N_14581,N_14413);
nand U14710 (N_14710,N_14496,N_14469);
nand U14711 (N_14711,N_14583,N_14599);
xor U14712 (N_14712,N_14529,N_14587);
and U14713 (N_14713,N_14561,N_14573);
nor U14714 (N_14714,N_14473,N_14444);
nor U14715 (N_14715,N_14453,N_14473);
xor U14716 (N_14716,N_14433,N_14470);
xnor U14717 (N_14717,N_14499,N_14498);
or U14718 (N_14718,N_14593,N_14530);
nor U14719 (N_14719,N_14430,N_14517);
nand U14720 (N_14720,N_14590,N_14480);
xnor U14721 (N_14721,N_14568,N_14565);
and U14722 (N_14722,N_14514,N_14589);
and U14723 (N_14723,N_14502,N_14511);
xnor U14724 (N_14724,N_14439,N_14535);
and U14725 (N_14725,N_14420,N_14414);
nand U14726 (N_14726,N_14562,N_14531);
xnor U14727 (N_14727,N_14403,N_14441);
and U14728 (N_14728,N_14423,N_14495);
nor U14729 (N_14729,N_14431,N_14459);
xnor U14730 (N_14730,N_14480,N_14409);
and U14731 (N_14731,N_14483,N_14548);
nand U14732 (N_14732,N_14593,N_14527);
nand U14733 (N_14733,N_14572,N_14578);
nand U14734 (N_14734,N_14546,N_14568);
nand U14735 (N_14735,N_14528,N_14433);
xor U14736 (N_14736,N_14584,N_14457);
or U14737 (N_14737,N_14421,N_14533);
nand U14738 (N_14738,N_14471,N_14441);
nand U14739 (N_14739,N_14451,N_14445);
nor U14740 (N_14740,N_14518,N_14536);
nand U14741 (N_14741,N_14454,N_14466);
or U14742 (N_14742,N_14564,N_14597);
or U14743 (N_14743,N_14403,N_14573);
nor U14744 (N_14744,N_14530,N_14426);
and U14745 (N_14745,N_14555,N_14540);
nand U14746 (N_14746,N_14538,N_14569);
nor U14747 (N_14747,N_14566,N_14435);
nor U14748 (N_14748,N_14491,N_14497);
nor U14749 (N_14749,N_14574,N_14563);
xor U14750 (N_14750,N_14468,N_14409);
nand U14751 (N_14751,N_14523,N_14435);
nor U14752 (N_14752,N_14430,N_14458);
or U14753 (N_14753,N_14526,N_14556);
xnor U14754 (N_14754,N_14598,N_14538);
nand U14755 (N_14755,N_14551,N_14493);
xor U14756 (N_14756,N_14536,N_14467);
and U14757 (N_14757,N_14512,N_14511);
or U14758 (N_14758,N_14557,N_14480);
nand U14759 (N_14759,N_14534,N_14516);
and U14760 (N_14760,N_14523,N_14547);
or U14761 (N_14761,N_14545,N_14564);
or U14762 (N_14762,N_14547,N_14486);
or U14763 (N_14763,N_14425,N_14474);
xor U14764 (N_14764,N_14408,N_14412);
or U14765 (N_14765,N_14437,N_14432);
or U14766 (N_14766,N_14440,N_14488);
or U14767 (N_14767,N_14595,N_14512);
nand U14768 (N_14768,N_14481,N_14476);
nor U14769 (N_14769,N_14442,N_14439);
nor U14770 (N_14770,N_14401,N_14427);
nor U14771 (N_14771,N_14556,N_14487);
xnor U14772 (N_14772,N_14505,N_14407);
nand U14773 (N_14773,N_14406,N_14555);
nor U14774 (N_14774,N_14477,N_14560);
nor U14775 (N_14775,N_14560,N_14444);
and U14776 (N_14776,N_14484,N_14430);
and U14777 (N_14777,N_14457,N_14411);
nor U14778 (N_14778,N_14523,N_14432);
xnor U14779 (N_14779,N_14583,N_14432);
nand U14780 (N_14780,N_14486,N_14408);
nor U14781 (N_14781,N_14565,N_14489);
nor U14782 (N_14782,N_14499,N_14506);
and U14783 (N_14783,N_14514,N_14596);
xor U14784 (N_14784,N_14473,N_14575);
xnor U14785 (N_14785,N_14489,N_14441);
nand U14786 (N_14786,N_14482,N_14477);
nand U14787 (N_14787,N_14478,N_14541);
or U14788 (N_14788,N_14526,N_14456);
nor U14789 (N_14789,N_14415,N_14593);
xnor U14790 (N_14790,N_14416,N_14461);
or U14791 (N_14791,N_14552,N_14454);
nand U14792 (N_14792,N_14402,N_14465);
and U14793 (N_14793,N_14401,N_14490);
nor U14794 (N_14794,N_14466,N_14538);
xor U14795 (N_14795,N_14482,N_14479);
or U14796 (N_14796,N_14552,N_14586);
and U14797 (N_14797,N_14401,N_14498);
or U14798 (N_14798,N_14476,N_14482);
nand U14799 (N_14799,N_14548,N_14475);
nor U14800 (N_14800,N_14628,N_14780);
nand U14801 (N_14801,N_14751,N_14776);
xor U14802 (N_14802,N_14755,N_14789);
and U14803 (N_14803,N_14699,N_14785);
and U14804 (N_14804,N_14795,N_14786);
nor U14805 (N_14805,N_14706,N_14792);
and U14806 (N_14806,N_14668,N_14689);
or U14807 (N_14807,N_14770,N_14667);
nand U14808 (N_14808,N_14700,N_14688);
xor U14809 (N_14809,N_14680,N_14767);
xor U14810 (N_14810,N_14763,N_14744);
and U14811 (N_14811,N_14707,N_14708);
or U14812 (N_14812,N_14606,N_14656);
and U14813 (N_14813,N_14794,N_14641);
nor U14814 (N_14814,N_14650,N_14748);
and U14815 (N_14815,N_14727,N_14649);
or U14816 (N_14816,N_14670,N_14690);
nand U14817 (N_14817,N_14623,N_14711);
and U14818 (N_14818,N_14791,N_14798);
and U14819 (N_14819,N_14716,N_14626);
or U14820 (N_14820,N_14646,N_14730);
or U14821 (N_14821,N_14639,N_14788);
nor U14822 (N_14822,N_14677,N_14603);
or U14823 (N_14823,N_14745,N_14790);
or U14824 (N_14824,N_14671,N_14661);
nand U14825 (N_14825,N_14771,N_14600);
nand U14826 (N_14826,N_14756,N_14613);
or U14827 (N_14827,N_14753,N_14681);
nor U14828 (N_14828,N_14718,N_14799);
and U14829 (N_14829,N_14651,N_14724);
xor U14830 (N_14830,N_14666,N_14608);
and U14831 (N_14831,N_14679,N_14741);
or U14832 (N_14832,N_14652,N_14687);
nand U14833 (N_14833,N_14634,N_14750);
xor U14834 (N_14834,N_14728,N_14775);
nand U14835 (N_14835,N_14635,N_14622);
nand U14836 (N_14836,N_14644,N_14604);
or U14837 (N_14837,N_14605,N_14709);
nand U14838 (N_14838,N_14740,N_14697);
nor U14839 (N_14839,N_14781,N_14654);
xor U14840 (N_14840,N_14673,N_14778);
and U14841 (N_14841,N_14637,N_14682);
nor U14842 (N_14842,N_14742,N_14645);
xor U14843 (N_14843,N_14643,N_14664);
xor U14844 (N_14844,N_14692,N_14705);
xor U14845 (N_14845,N_14787,N_14624);
or U14846 (N_14846,N_14746,N_14659);
and U14847 (N_14847,N_14757,N_14675);
nor U14848 (N_14848,N_14616,N_14638);
xnor U14849 (N_14849,N_14734,N_14725);
and U14850 (N_14850,N_14717,N_14760);
nand U14851 (N_14851,N_14738,N_14607);
nand U14852 (N_14852,N_14683,N_14722);
or U14853 (N_14853,N_14739,N_14618);
and U14854 (N_14854,N_14769,N_14774);
nand U14855 (N_14855,N_14632,N_14721);
nor U14856 (N_14856,N_14797,N_14733);
nor U14857 (N_14857,N_14630,N_14715);
or U14858 (N_14858,N_14619,N_14658);
xnor U14859 (N_14859,N_14768,N_14636);
or U14860 (N_14860,N_14676,N_14601);
nor U14861 (N_14861,N_14633,N_14698);
nand U14862 (N_14862,N_14719,N_14762);
or U14863 (N_14863,N_14761,N_14653);
or U14864 (N_14864,N_14640,N_14696);
xor U14865 (N_14865,N_14686,N_14726);
nand U14866 (N_14866,N_14758,N_14735);
xnor U14867 (N_14867,N_14627,N_14710);
or U14868 (N_14868,N_14737,N_14684);
nor U14869 (N_14869,N_14796,N_14663);
nand U14870 (N_14870,N_14783,N_14609);
xnor U14871 (N_14871,N_14747,N_14703);
and U14872 (N_14872,N_14779,N_14772);
xnor U14873 (N_14873,N_14773,N_14648);
or U14874 (N_14874,N_14702,N_14691);
xor U14875 (N_14875,N_14615,N_14665);
or U14876 (N_14876,N_14713,N_14701);
nor U14877 (N_14877,N_14610,N_14612);
nand U14878 (N_14878,N_14731,N_14662);
or U14879 (N_14879,N_14712,N_14629);
or U14880 (N_14880,N_14620,N_14749);
and U14881 (N_14881,N_14611,N_14660);
and U14882 (N_14882,N_14631,N_14759);
nor U14883 (N_14883,N_14655,N_14723);
nor U14884 (N_14884,N_14694,N_14782);
nand U14885 (N_14885,N_14704,N_14765);
nor U14886 (N_14886,N_14678,N_14642);
or U14887 (N_14887,N_14647,N_14766);
nand U14888 (N_14888,N_14685,N_14714);
nand U14889 (N_14889,N_14674,N_14784);
and U14890 (N_14890,N_14617,N_14754);
nor U14891 (N_14891,N_14720,N_14793);
nand U14892 (N_14892,N_14621,N_14752);
or U14893 (N_14893,N_14625,N_14669);
nor U14894 (N_14894,N_14602,N_14732);
and U14895 (N_14895,N_14614,N_14693);
nand U14896 (N_14896,N_14764,N_14777);
or U14897 (N_14897,N_14672,N_14657);
nor U14898 (N_14898,N_14695,N_14729);
or U14899 (N_14899,N_14736,N_14743);
nor U14900 (N_14900,N_14664,N_14701);
or U14901 (N_14901,N_14683,N_14785);
nor U14902 (N_14902,N_14608,N_14636);
and U14903 (N_14903,N_14661,N_14636);
xnor U14904 (N_14904,N_14651,N_14730);
or U14905 (N_14905,N_14692,N_14677);
or U14906 (N_14906,N_14635,N_14697);
nand U14907 (N_14907,N_14714,N_14655);
xor U14908 (N_14908,N_14754,N_14784);
nor U14909 (N_14909,N_14672,N_14601);
nand U14910 (N_14910,N_14731,N_14712);
and U14911 (N_14911,N_14760,N_14783);
nor U14912 (N_14912,N_14764,N_14603);
nand U14913 (N_14913,N_14685,N_14679);
nor U14914 (N_14914,N_14631,N_14660);
nor U14915 (N_14915,N_14776,N_14672);
nand U14916 (N_14916,N_14713,N_14602);
or U14917 (N_14917,N_14671,N_14795);
xor U14918 (N_14918,N_14691,N_14779);
or U14919 (N_14919,N_14696,N_14651);
nor U14920 (N_14920,N_14666,N_14618);
xor U14921 (N_14921,N_14712,N_14795);
or U14922 (N_14922,N_14642,N_14621);
xor U14923 (N_14923,N_14717,N_14767);
or U14924 (N_14924,N_14678,N_14704);
or U14925 (N_14925,N_14725,N_14629);
and U14926 (N_14926,N_14686,N_14608);
or U14927 (N_14927,N_14654,N_14766);
nand U14928 (N_14928,N_14709,N_14630);
xnor U14929 (N_14929,N_14798,N_14726);
nand U14930 (N_14930,N_14616,N_14678);
and U14931 (N_14931,N_14624,N_14670);
xnor U14932 (N_14932,N_14724,N_14716);
nor U14933 (N_14933,N_14775,N_14798);
or U14934 (N_14934,N_14662,N_14795);
xnor U14935 (N_14935,N_14751,N_14724);
nor U14936 (N_14936,N_14640,N_14791);
xor U14937 (N_14937,N_14737,N_14600);
and U14938 (N_14938,N_14660,N_14690);
nor U14939 (N_14939,N_14691,N_14670);
nor U14940 (N_14940,N_14794,N_14741);
xnor U14941 (N_14941,N_14736,N_14735);
nor U14942 (N_14942,N_14770,N_14630);
xor U14943 (N_14943,N_14654,N_14772);
and U14944 (N_14944,N_14755,N_14796);
and U14945 (N_14945,N_14688,N_14656);
nand U14946 (N_14946,N_14771,N_14701);
and U14947 (N_14947,N_14796,N_14730);
xnor U14948 (N_14948,N_14630,N_14690);
and U14949 (N_14949,N_14612,N_14720);
xor U14950 (N_14950,N_14760,N_14766);
and U14951 (N_14951,N_14610,N_14726);
or U14952 (N_14952,N_14625,N_14681);
nand U14953 (N_14953,N_14735,N_14616);
nand U14954 (N_14954,N_14682,N_14772);
nor U14955 (N_14955,N_14660,N_14722);
xor U14956 (N_14956,N_14633,N_14687);
nor U14957 (N_14957,N_14610,N_14664);
or U14958 (N_14958,N_14739,N_14690);
nor U14959 (N_14959,N_14767,N_14705);
xor U14960 (N_14960,N_14607,N_14797);
and U14961 (N_14961,N_14644,N_14600);
or U14962 (N_14962,N_14759,N_14640);
and U14963 (N_14963,N_14755,N_14729);
or U14964 (N_14964,N_14701,N_14748);
and U14965 (N_14965,N_14643,N_14749);
xor U14966 (N_14966,N_14698,N_14724);
nor U14967 (N_14967,N_14726,N_14790);
nand U14968 (N_14968,N_14779,N_14654);
nand U14969 (N_14969,N_14675,N_14782);
or U14970 (N_14970,N_14754,N_14757);
xor U14971 (N_14971,N_14786,N_14725);
nand U14972 (N_14972,N_14799,N_14659);
or U14973 (N_14973,N_14617,N_14616);
nor U14974 (N_14974,N_14708,N_14649);
xor U14975 (N_14975,N_14658,N_14787);
nor U14976 (N_14976,N_14605,N_14660);
xor U14977 (N_14977,N_14627,N_14703);
and U14978 (N_14978,N_14789,N_14612);
nor U14979 (N_14979,N_14734,N_14730);
nand U14980 (N_14980,N_14718,N_14749);
xnor U14981 (N_14981,N_14769,N_14659);
nor U14982 (N_14982,N_14706,N_14610);
nor U14983 (N_14983,N_14774,N_14704);
or U14984 (N_14984,N_14741,N_14650);
xnor U14985 (N_14985,N_14775,N_14781);
nand U14986 (N_14986,N_14651,N_14741);
and U14987 (N_14987,N_14610,N_14701);
or U14988 (N_14988,N_14704,N_14659);
xnor U14989 (N_14989,N_14778,N_14622);
nand U14990 (N_14990,N_14661,N_14699);
nand U14991 (N_14991,N_14795,N_14797);
or U14992 (N_14992,N_14755,N_14684);
xor U14993 (N_14993,N_14762,N_14760);
nand U14994 (N_14994,N_14718,N_14737);
nor U14995 (N_14995,N_14745,N_14644);
or U14996 (N_14996,N_14732,N_14692);
nor U14997 (N_14997,N_14742,N_14612);
xor U14998 (N_14998,N_14717,N_14644);
nor U14999 (N_14999,N_14758,N_14668);
and U15000 (N_15000,N_14858,N_14964);
xnor U15001 (N_15001,N_14843,N_14856);
and U15002 (N_15002,N_14851,N_14966);
xnor U15003 (N_15003,N_14854,N_14979);
xor U15004 (N_15004,N_14880,N_14951);
nor U15005 (N_15005,N_14827,N_14803);
and U15006 (N_15006,N_14848,N_14958);
xor U15007 (N_15007,N_14907,N_14932);
or U15008 (N_15008,N_14996,N_14938);
nor U15009 (N_15009,N_14894,N_14929);
nand U15010 (N_15010,N_14835,N_14896);
and U15011 (N_15011,N_14837,N_14826);
nand U15012 (N_15012,N_14988,N_14899);
or U15013 (N_15013,N_14949,N_14847);
nand U15014 (N_15014,N_14945,N_14865);
nand U15015 (N_15015,N_14961,N_14992);
and U15016 (N_15016,N_14860,N_14890);
and U15017 (N_15017,N_14902,N_14963);
or U15018 (N_15018,N_14942,N_14967);
xnor U15019 (N_15019,N_14886,N_14972);
nand U15020 (N_15020,N_14874,N_14838);
or U15021 (N_15021,N_14940,N_14878);
or U15022 (N_15022,N_14864,N_14937);
nor U15023 (N_15023,N_14823,N_14813);
nand U15024 (N_15024,N_14871,N_14916);
xor U15025 (N_15025,N_14849,N_14872);
and U15026 (N_15026,N_14859,N_14946);
xor U15027 (N_15027,N_14959,N_14834);
nand U15028 (N_15028,N_14952,N_14881);
or U15029 (N_15029,N_14810,N_14926);
nor U15030 (N_15030,N_14917,N_14969);
xor U15031 (N_15031,N_14876,N_14804);
nand U15032 (N_15032,N_14825,N_14944);
xor U15033 (N_15033,N_14831,N_14844);
xor U15034 (N_15034,N_14913,N_14976);
and U15035 (N_15035,N_14805,N_14820);
nand U15036 (N_15036,N_14889,N_14869);
and U15037 (N_15037,N_14991,N_14978);
or U15038 (N_15038,N_14891,N_14863);
xnor U15039 (N_15039,N_14850,N_14960);
nor U15040 (N_15040,N_14806,N_14822);
nand U15041 (N_15041,N_14846,N_14955);
nor U15042 (N_15042,N_14885,N_14883);
nand U15043 (N_15043,N_14971,N_14970);
nand U15044 (N_15044,N_14909,N_14857);
or U15045 (N_15045,N_14931,N_14974);
xnor U15046 (N_15046,N_14832,N_14948);
nand U15047 (N_15047,N_14947,N_14898);
nand U15048 (N_15048,N_14817,N_14953);
or U15049 (N_15049,N_14918,N_14998);
or U15050 (N_15050,N_14980,N_14830);
and U15051 (N_15051,N_14892,N_14845);
nand U15052 (N_15052,N_14868,N_14995);
xnor U15053 (N_15053,N_14914,N_14954);
and U15054 (N_15054,N_14939,N_14919);
and U15055 (N_15055,N_14920,N_14922);
nor U15056 (N_15056,N_14809,N_14821);
or U15057 (N_15057,N_14866,N_14815);
xnor U15058 (N_15058,N_14893,N_14906);
nor U15059 (N_15059,N_14936,N_14841);
nor U15060 (N_15060,N_14957,N_14997);
xor U15061 (N_15061,N_14875,N_14927);
or U15062 (N_15062,N_14994,N_14956);
and U15063 (N_15063,N_14903,N_14839);
and U15064 (N_15064,N_14819,N_14867);
nand U15065 (N_15065,N_14877,N_14836);
nor U15066 (N_15066,N_14814,N_14811);
or U15067 (N_15067,N_14925,N_14816);
and U15068 (N_15068,N_14853,N_14862);
nor U15069 (N_15069,N_14879,N_14924);
nor U15070 (N_15070,N_14829,N_14905);
nand U15071 (N_15071,N_14983,N_14928);
or U15072 (N_15072,N_14812,N_14808);
and U15073 (N_15073,N_14873,N_14887);
xor U15074 (N_15074,N_14912,N_14934);
xor U15075 (N_15075,N_14982,N_14977);
and U15076 (N_15076,N_14973,N_14842);
xnor U15077 (N_15077,N_14968,N_14824);
or U15078 (N_15078,N_14900,N_14802);
nand U15079 (N_15079,N_14915,N_14870);
xor U15080 (N_15080,N_14807,N_14990);
nor U15081 (N_15081,N_14950,N_14941);
xnor U15082 (N_15082,N_14975,N_14933);
nor U15083 (N_15083,N_14828,N_14908);
or U15084 (N_15084,N_14855,N_14861);
nand U15085 (N_15085,N_14910,N_14943);
xnor U15086 (N_15086,N_14901,N_14989);
nor U15087 (N_15087,N_14962,N_14930);
xor U15088 (N_15088,N_14852,N_14904);
nand U15089 (N_15089,N_14999,N_14888);
and U15090 (N_15090,N_14935,N_14801);
or U15091 (N_15091,N_14921,N_14993);
xnor U15092 (N_15092,N_14987,N_14965);
or U15093 (N_15093,N_14911,N_14800);
or U15094 (N_15094,N_14984,N_14895);
or U15095 (N_15095,N_14884,N_14833);
nand U15096 (N_15096,N_14923,N_14986);
xnor U15097 (N_15097,N_14818,N_14840);
and U15098 (N_15098,N_14882,N_14897);
xor U15099 (N_15099,N_14985,N_14981);
nor U15100 (N_15100,N_14965,N_14904);
nand U15101 (N_15101,N_14989,N_14920);
and U15102 (N_15102,N_14846,N_14872);
nand U15103 (N_15103,N_14876,N_14943);
nor U15104 (N_15104,N_14818,N_14940);
or U15105 (N_15105,N_14992,N_14965);
and U15106 (N_15106,N_14995,N_14916);
nor U15107 (N_15107,N_14864,N_14905);
xor U15108 (N_15108,N_14947,N_14820);
xnor U15109 (N_15109,N_14837,N_14817);
xor U15110 (N_15110,N_14809,N_14971);
nand U15111 (N_15111,N_14897,N_14831);
xor U15112 (N_15112,N_14846,N_14849);
and U15113 (N_15113,N_14810,N_14820);
nor U15114 (N_15114,N_14969,N_14939);
or U15115 (N_15115,N_14951,N_14836);
xnor U15116 (N_15116,N_14918,N_14867);
nand U15117 (N_15117,N_14889,N_14986);
or U15118 (N_15118,N_14941,N_14860);
nand U15119 (N_15119,N_14844,N_14812);
xnor U15120 (N_15120,N_14831,N_14944);
nor U15121 (N_15121,N_14852,N_14895);
or U15122 (N_15122,N_14807,N_14890);
and U15123 (N_15123,N_14947,N_14915);
nand U15124 (N_15124,N_14943,N_14988);
nor U15125 (N_15125,N_14989,N_14948);
nor U15126 (N_15126,N_14948,N_14888);
nor U15127 (N_15127,N_14840,N_14849);
nor U15128 (N_15128,N_14972,N_14949);
xnor U15129 (N_15129,N_14999,N_14855);
xor U15130 (N_15130,N_14942,N_14922);
nand U15131 (N_15131,N_14878,N_14900);
nand U15132 (N_15132,N_14825,N_14818);
or U15133 (N_15133,N_14843,N_14948);
nand U15134 (N_15134,N_14885,N_14935);
xnor U15135 (N_15135,N_14894,N_14910);
nor U15136 (N_15136,N_14974,N_14830);
nand U15137 (N_15137,N_14877,N_14961);
nand U15138 (N_15138,N_14927,N_14830);
or U15139 (N_15139,N_14956,N_14816);
nor U15140 (N_15140,N_14861,N_14894);
nand U15141 (N_15141,N_14913,N_14848);
or U15142 (N_15142,N_14935,N_14891);
and U15143 (N_15143,N_14802,N_14951);
xnor U15144 (N_15144,N_14820,N_14890);
or U15145 (N_15145,N_14885,N_14856);
nand U15146 (N_15146,N_14895,N_14893);
nor U15147 (N_15147,N_14932,N_14988);
nor U15148 (N_15148,N_14890,N_14937);
and U15149 (N_15149,N_14935,N_14948);
or U15150 (N_15150,N_14830,N_14990);
or U15151 (N_15151,N_14835,N_14879);
xnor U15152 (N_15152,N_14824,N_14802);
and U15153 (N_15153,N_14994,N_14841);
and U15154 (N_15154,N_14879,N_14923);
nand U15155 (N_15155,N_14982,N_14851);
xor U15156 (N_15156,N_14917,N_14999);
nand U15157 (N_15157,N_14908,N_14904);
nor U15158 (N_15158,N_14991,N_14950);
nor U15159 (N_15159,N_14881,N_14826);
or U15160 (N_15160,N_14810,N_14861);
and U15161 (N_15161,N_14863,N_14819);
xnor U15162 (N_15162,N_14930,N_14990);
or U15163 (N_15163,N_14867,N_14853);
nand U15164 (N_15164,N_14953,N_14841);
xor U15165 (N_15165,N_14997,N_14996);
xor U15166 (N_15166,N_14963,N_14908);
nand U15167 (N_15167,N_14982,N_14847);
nand U15168 (N_15168,N_14980,N_14958);
nor U15169 (N_15169,N_14931,N_14855);
nor U15170 (N_15170,N_14849,N_14805);
nor U15171 (N_15171,N_14925,N_14911);
nand U15172 (N_15172,N_14872,N_14988);
or U15173 (N_15173,N_14874,N_14904);
or U15174 (N_15174,N_14951,N_14949);
nand U15175 (N_15175,N_14829,N_14953);
and U15176 (N_15176,N_14869,N_14900);
nand U15177 (N_15177,N_14844,N_14852);
nand U15178 (N_15178,N_14905,N_14995);
nand U15179 (N_15179,N_14992,N_14810);
nand U15180 (N_15180,N_14972,N_14806);
nor U15181 (N_15181,N_14819,N_14978);
xnor U15182 (N_15182,N_14922,N_14833);
nand U15183 (N_15183,N_14933,N_14853);
or U15184 (N_15184,N_14989,N_14955);
nand U15185 (N_15185,N_14911,N_14973);
nand U15186 (N_15186,N_14958,N_14921);
and U15187 (N_15187,N_14970,N_14892);
nand U15188 (N_15188,N_14818,N_14838);
nor U15189 (N_15189,N_14801,N_14959);
or U15190 (N_15190,N_14883,N_14915);
nand U15191 (N_15191,N_14900,N_14810);
or U15192 (N_15192,N_14959,N_14933);
nor U15193 (N_15193,N_14957,N_14872);
or U15194 (N_15194,N_14960,N_14961);
or U15195 (N_15195,N_14816,N_14946);
xor U15196 (N_15196,N_14837,N_14866);
and U15197 (N_15197,N_14861,N_14836);
or U15198 (N_15198,N_14998,N_14882);
and U15199 (N_15199,N_14820,N_14930);
and U15200 (N_15200,N_15086,N_15123);
nor U15201 (N_15201,N_15143,N_15000);
and U15202 (N_15202,N_15008,N_15190);
and U15203 (N_15203,N_15195,N_15130);
or U15204 (N_15204,N_15129,N_15041);
and U15205 (N_15205,N_15074,N_15018);
nand U15206 (N_15206,N_15128,N_15030);
nor U15207 (N_15207,N_15025,N_15164);
or U15208 (N_15208,N_15159,N_15026);
xor U15209 (N_15209,N_15015,N_15133);
nor U15210 (N_15210,N_15078,N_15155);
and U15211 (N_15211,N_15055,N_15170);
or U15212 (N_15212,N_15101,N_15099);
xor U15213 (N_15213,N_15047,N_15140);
xnor U15214 (N_15214,N_15134,N_15196);
nand U15215 (N_15215,N_15161,N_15027);
and U15216 (N_15216,N_15031,N_15070);
or U15217 (N_15217,N_15131,N_15054);
or U15218 (N_15218,N_15023,N_15189);
nand U15219 (N_15219,N_15034,N_15036);
xnor U15220 (N_15220,N_15142,N_15186);
nand U15221 (N_15221,N_15158,N_15040);
xor U15222 (N_15222,N_15132,N_15057);
nand U15223 (N_15223,N_15029,N_15028);
and U15224 (N_15224,N_15065,N_15084);
nand U15225 (N_15225,N_15184,N_15137);
and U15226 (N_15226,N_15092,N_15192);
and U15227 (N_15227,N_15116,N_15096);
nand U15228 (N_15228,N_15004,N_15177);
and U15229 (N_15229,N_15061,N_15102);
xor U15230 (N_15230,N_15194,N_15156);
nand U15231 (N_15231,N_15067,N_15037);
nor U15232 (N_15232,N_15012,N_15060);
and U15233 (N_15233,N_15112,N_15151);
and U15234 (N_15234,N_15089,N_15022);
xnor U15235 (N_15235,N_15197,N_15064);
or U15236 (N_15236,N_15149,N_15066);
or U15237 (N_15237,N_15139,N_15111);
or U15238 (N_15238,N_15152,N_15162);
xnor U15239 (N_15239,N_15125,N_15021);
nor U15240 (N_15240,N_15010,N_15183);
or U15241 (N_15241,N_15188,N_15006);
nand U15242 (N_15242,N_15119,N_15051);
xnor U15243 (N_15243,N_15135,N_15053);
and U15244 (N_15244,N_15115,N_15114);
nor U15245 (N_15245,N_15118,N_15091);
xor U15246 (N_15246,N_15165,N_15087);
nor U15247 (N_15247,N_15168,N_15174);
xor U15248 (N_15248,N_15069,N_15154);
xnor U15249 (N_15249,N_15124,N_15150);
or U15250 (N_15250,N_15083,N_15059);
nand U15251 (N_15251,N_15014,N_15146);
nand U15252 (N_15252,N_15182,N_15173);
xor U15253 (N_15253,N_15180,N_15056);
and U15254 (N_15254,N_15121,N_15003);
and U15255 (N_15255,N_15082,N_15122);
nor U15256 (N_15256,N_15153,N_15043);
nor U15257 (N_15257,N_15163,N_15048);
or U15258 (N_15258,N_15079,N_15073);
nor U15259 (N_15259,N_15167,N_15058);
nor U15260 (N_15260,N_15032,N_15001);
nand U15261 (N_15261,N_15024,N_15016);
nand U15262 (N_15262,N_15094,N_15002);
nor U15263 (N_15263,N_15103,N_15166);
xor U15264 (N_15264,N_15187,N_15080);
nand U15265 (N_15265,N_15068,N_15093);
nor U15266 (N_15266,N_15105,N_15100);
nor U15267 (N_15267,N_15108,N_15145);
nor U15268 (N_15268,N_15088,N_15045);
nand U15269 (N_15269,N_15160,N_15020);
nand U15270 (N_15270,N_15178,N_15141);
and U15271 (N_15271,N_15193,N_15097);
and U15272 (N_15272,N_15052,N_15181);
nand U15273 (N_15273,N_15148,N_15157);
xor U15274 (N_15274,N_15042,N_15090);
or U15275 (N_15275,N_15138,N_15147);
nor U15276 (N_15276,N_15107,N_15172);
nand U15277 (N_15277,N_15179,N_15198);
nor U15278 (N_15278,N_15169,N_15106);
or U15279 (N_15279,N_15110,N_15171);
and U15280 (N_15280,N_15019,N_15009);
xor U15281 (N_15281,N_15185,N_15176);
or U15282 (N_15282,N_15113,N_15136);
nand U15283 (N_15283,N_15039,N_15062);
and U15284 (N_15284,N_15117,N_15081);
and U15285 (N_15285,N_15085,N_15199);
nor U15286 (N_15286,N_15175,N_15127);
nand U15287 (N_15287,N_15076,N_15098);
or U15288 (N_15288,N_15007,N_15038);
or U15289 (N_15289,N_15126,N_15044);
nor U15290 (N_15290,N_15005,N_15013);
and U15291 (N_15291,N_15144,N_15049);
or U15292 (N_15292,N_15095,N_15077);
nand U15293 (N_15293,N_15063,N_15046);
nand U15294 (N_15294,N_15011,N_15109);
xor U15295 (N_15295,N_15035,N_15075);
nor U15296 (N_15296,N_15072,N_15120);
nor U15297 (N_15297,N_15017,N_15071);
nor U15298 (N_15298,N_15104,N_15191);
nand U15299 (N_15299,N_15050,N_15033);
or U15300 (N_15300,N_15035,N_15148);
nor U15301 (N_15301,N_15080,N_15136);
or U15302 (N_15302,N_15168,N_15082);
and U15303 (N_15303,N_15101,N_15156);
nor U15304 (N_15304,N_15038,N_15130);
xnor U15305 (N_15305,N_15189,N_15016);
and U15306 (N_15306,N_15033,N_15076);
xor U15307 (N_15307,N_15115,N_15194);
or U15308 (N_15308,N_15182,N_15172);
and U15309 (N_15309,N_15185,N_15000);
or U15310 (N_15310,N_15094,N_15073);
nor U15311 (N_15311,N_15125,N_15158);
nor U15312 (N_15312,N_15006,N_15068);
nand U15313 (N_15313,N_15085,N_15013);
or U15314 (N_15314,N_15066,N_15115);
nor U15315 (N_15315,N_15074,N_15177);
and U15316 (N_15316,N_15013,N_15140);
and U15317 (N_15317,N_15132,N_15116);
xnor U15318 (N_15318,N_15126,N_15195);
nor U15319 (N_15319,N_15039,N_15032);
nand U15320 (N_15320,N_15014,N_15133);
and U15321 (N_15321,N_15147,N_15113);
and U15322 (N_15322,N_15173,N_15039);
nand U15323 (N_15323,N_15109,N_15026);
nor U15324 (N_15324,N_15058,N_15076);
xnor U15325 (N_15325,N_15062,N_15187);
and U15326 (N_15326,N_15125,N_15193);
or U15327 (N_15327,N_15189,N_15168);
xor U15328 (N_15328,N_15046,N_15007);
nand U15329 (N_15329,N_15129,N_15006);
xor U15330 (N_15330,N_15040,N_15146);
xnor U15331 (N_15331,N_15117,N_15190);
and U15332 (N_15332,N_15071,N_15131);
and U15333 (N_15333,N_15114,N_15033);
or U15334 (N_15334,N_15145,N_15162);
nand U15335 (N_15335,N_15100,N_15111);
nand U15336 (N_15336,N_15148,N_15120);
nor U15337 (N_15337,N_15169,N_15152);
and U15338 (N_15338,N_15108,N_15074);
and U15339 (N_15339,N_15162,N_15081);
and U15340 (N_15340,N_15086,N_15060);
xor U15341 (N_15341,N_15111,N_15052);
or U15342 (N_15342,N_15008,N_15084);
and U15343 (N_15343,N_15174,N_15106);
or U15344 (N_15344,N_15110,N_15157);
and U15345 (N_15345,N_15100,N_15149);
nor U15346 (N_15346,N_15103,N_15198);
and U15347 (N_15347,N_15132,N_15166);
nor U15348 (N_15348,N_15035,N_15109);
and U15349 (N_15349,N_15009,N_15049);
and U15350 (N_15350,N_15129,N_15034);
or U15351 (N_15351,N_15011,N_15037);
nand U15352 (N_15352,N_15090,N_15115);
nor U15353 (N_15353,N_15113,N_15089);
and U15354 (N_15354,N_15146,N_15170);
nand U15355 (N_15355,N_15157,N_15109);
and U15356 (N_15356,N_15004,N_15126);
and U15357 (N_15357,N_15172,N_15001);
nor U15358 (N_15358,N_15150,N_15074);
nor U15359 (N_15359,N_15116,N_15046);
nor U15360 (N_15360,N_15147,N_15176);
nor U15361 (N_15361,N_15091,N_15187);
nor U15362 (N_15362,N_15023,N_15113);
or U15363 (N_15363,N_15189,N_15156);
xnor U15364 (N_15364,N_15124,N_15007);
and U15365 (N_15365,N_15022,N_15093);
and U15366 (N_15366,N_15105,N_15074);
nand U15367 (N_15367,N_15071,N_15021);
and U15368 (N_15368,N_15132,N_15015);
xor U15369 (N_15369,N_15109,N_15002);
or U15370 (N_15370,N_15005,N_15148);
nand U15371 (N_15371,N_15032,N_15150);
nor U15372 (N_15372,N_15082,N_15145);
nand U15373 (N_15373,N_15121,N_15188);
and U15374 (N_15374,N_15065,N_15131);
nor U15375 (N_15375,N_15035,N_15122);
nor U15376 (N_15376,N_15076,N_15183);
nand U15377 (N_15377,N_15094,N_15035);
nand U15378 (N_15378,N_15046,N_15170);
nor U15379 (N_15379,N_15003,N_15168);
xnor U15380 (N_15380,N_15084,N_15195);
xnor U15381 (N_15381,N_15164,N_15041);
xnor U15382 (N_15382,N_15198,N_15180);
or U15383 (N_15383,N_15016,N_15192);
nand U15384 (N_15384,N_15085,N_15176);
and U15385 (N_15385,N_15034,N_15006);
or U15386 (N_15386,N_15140,N_15180);
xor U15387 (N_15387,N_15075,N_15077);
or U15388 (N_15388,N_15063,N_15058);
nor U15389 (N_15389,N_15156,N_15132);
nand U15390 (N_15390,N_15134,N_15159);
xor U15391 (N_15391,N_15108,N_15034);
or U15392 (N_15392,N_15033,N_15027);
xnor U15393 (N_15393,N_15074,N_15163);
nand U15394 (N_15394,N_15094,N_15104);
or U15395 (N_15395,N_15127,N_15014);
nor U15396 (N_15396,N_15107,N_15018);
nand U15397 (N_15397,N_15026,N_15066);
or U15398 (N_15398,N_15082,N_15129);
nor U15399 (N_15399,N_15098,N_15025);
nand U15400 (N_15400,N_15243,N_15372);
nor U15401 (N_15401,N_15292,N_15227);
nand U15402 (N_15402,N_15310,N_15321);
or U15403 (N_15403,N_15380,N_15350);
nor U15404 (N_15404,N_15211,N_15327);
or U15405 (N_15405,N_15214,N_15363);
nor U15406 (N_15406,N_15242,N_15283);
xor U15407 (N_15407,N_15273,N_15257);
xor U15408 (N_15408,N_15232,N_15376);
nor U15409 (N_15409,N_15276,N_15396);
or U15410 (N_15410,N_15342,N_15397);
xnor U15411 (N_15411,N_15209,N_15244);
nor U15412 (N_15412,N_15255,N_15216);
or U15413 (N_15413,N_15375,N_15371);
nor U15414 (N_15414,N_15382,N_15364);
nand U15415 (N_15415,N_15277,N_15206);
and U15416 (N_15416,N_15296,N_15381);
nand U15417 (N_15417,N_15286,N_15252);
nand U15418 (N_15418,N_15210,N_15305);
nor U15419 (N_15419,N_15339,N_15355);
nor U15420 (N_15420,N_15302,N_15308);
nor U15421 (N_15421,N_15386,N_15217);
and U15422 (N_15422,N_15278,N_15203);
or U15423 (N_15423,N_15299,N_15240);
nand U15424 (N_15424,N_15306,N_15247);
xnor U15425 (N_15425,N_15239,N_15220);
xnor U15426 (N_15426,N_15347,N_15314);
and U15427 (N_15427,N_15218,N_15204);
nor U15428 (N_15428,N_15213,N_15205);
nor U15429 (N_15429,N_15212,N_15280);
nor U15430 (N_15430,N_15236,N_15219);
and U15431 (N_15431,N_15285,N_15331);
or U15432 (N_15432,N_15329,N_15366);
xnor U15433 (N_15433,N_15361,N_15295);
xnor U15434 (N_15434,N_15266,N_15333);
nand U15435 (N_15435,N_15328,N_15385);
xnor U15436 (N_15436,N_15341,N_15313);
xnor U15437 (N_15437,N_15265,N_15332);
and U15438 (N_15438,N_15200,N_15297);
or U15439 (N_15439,N_15362,N_15369);
and U15440 (N_15440,N_15250,N_15245);
nand U15441 (N_15441,N_15272,N_15288);
nand U15442 (N_15442,N_15340,N_15323);
xor U15443 (N_15443,N_15222,N_15393);
and U15444 (N_15444,N_15330,N_15387);
xnor U15445 (N_15445,N_15258,N_15264);
nor U15446 (N_15446,N_15359,N_15253);
xnor U15447 (N_15447,N_15383,N_15298);
and U15448 (N_15448,N_15357,N_15399);
and U15449 (N_15449,N_15343,N_15263);
nand U15450 (N_15450,N_15349,N_15259);
xnor U15451 (N_15451,N_15237,N_15289);
and U15452 (N_15452,N_15368,N_15261);
or U15453 (N_15453,N_15307,N_15279);
or U15454 (N_15454,N_15300,N_15241);
or U15455 (N_15455,N_15284,N_15208);
nor U15456 (N_15456,N_15230,N_15224);
and U15457 (N_15457,N_15215,N_15294);
xor U15458 (N_15458,N_15271,N_15291);
and U15459 (N_15459,N_15377,N_15354);
nand U15460 (N_15460,N_15238,N_15389);
and U15461 (N_15461,N_15324,N_15390);
nor U15462 (N_15462,N_15348,N_15318);
nand U15463 (N_15463,N_15358,N_15351);
xnor U15464 (N_15464,N_15248,N_15246);
xnor U15465 (N_15465,N_15309,N_15353);
nor U15466 (N_15466,N_15326,N_15334);
and U15467 (N_15467,N_15370,N_15344);
nor U15468 (N_15468,N_15262,N_15225);
nor U15469 (N_15469,N_15395,N_15260);
or U15470 (N_15470,N_15202,N_15233);
nand U15471 (N_15471,N_15367,N_15269);
or U15472 (N_15472,N_15392,N_15378);
xnor U15473 (N_15473,N_15356,N_15394);
nor U15474 (N_15474,N_15228,N_15360);
nand U15475 (N_15475,N_15388,N_15384);
and U15476 (N_15476,N_15249,N_15274);
nor U15477 (N_15477,N_15398,N_15374);
nor U15478 (N_15478,N_15315,N_15293);
xnor U15479 (N_15479,N_15231,N_15322);
xnor U15480 (N_15480,N_15290,N_15270);
or U15481 (N_15481,N_15325,N_15320);
nand U15482 (N_15482,N_15336,N_15365);
xnor U15483 (N_15483,N_15235,N_15201);
and U15484 (N_15484,N_15223,N_15352);
nand U15485 (N_15485,N_15281,N_15345);
nor U15486 (N_15486,N_15256,N_15254);
nand U15487 (N_15487,N_15304,N_15373);
nand U15488 (N_15488,N_15303,N_15312);
or U15489 (N_15489,N_15335,N_15267);
nor U15490 (N_15490,N_15207,N_15268);
or U15491 (N_15491,N_15316,N_15226);
nor U15492 (N_15492,N_15229,N_15337);
xor U15493 (N_15493,N_15319,N_15251);
xnor U15494 (N_15494,N_15338,N_15391);
or U15495 (N_15495,N_15282,N_15287);
xnor U15496 (N_15496,N_15317,N_15301);
and U15497 (N_15497,N_15379,N_15346);
nor U15498 (N_15498,N_15311,N_15234);
nand U15499 (N_15499,N_15221,N_15275);
xnor U15500 (N_15500,N_15301,N_15322);
nor U15501 (N_15501,N_15352,N_15301);
or U15502 (N_15502,N_15324,N_15203);
and U15503 (N_15503,N_15306,N_15337);
nor U15504 (N_15504,N_15379,N_15307);
and U15505 (N_15505,N_15239,N_15397);
nor U15506 (N_15506,N_15394,N_15257);
or U15507 (N_15507,N_15370,N_15311);
xor U15508 (N_15508,N_15226,N_15285);
nand U15509 (N_15509,N_15331,N_15237);
and U15510 (N_15510,N_15345,N_15319);
xnor U15511 (N_15511,N_15399,N_15395);
nor U15512 (N_15512,N_15381,N_15352);
nor U15513 (N_15513,N_15347,N_15258);
or U15514 (N_15514,N_15371,N_15219);
nand U15515 (N_15515,N_15289,N_15234);
nand U15516 (N_15516,N_15217,N_15219);
nor U15517 (N_15517,N_15339,N_15279);
xnor U15518 (N_15518,N_15339,N_15310);
xor U15519 (N_15519,N_15392,N_15245);
xor U15520 (N_15520,N_15248,N_15282);
nor U15521 (N_15521,N_15287,N_15236);
and U15522 (N_15522,N_15248,N_15399);
and U15523 (N_15523,N_15247,N_15217);
or U15524 (N_15524,N_15294,N_15230);
xor U15525 (N_15525,N_15258,N_15232);
nor U15526 (N_15526,N_15278,N_15250);
and U15527 (N_15527,N_15307,N_15295);
nand U15528 (N_15528,N_15267,N_15323);
or U15529 (N_15529,N_15203,N_15316);
nand U15530 (N_15530,N_15284,N_15325);
nand U15531 (N_15531,N_15327,N_15305);
nor U15532 (N_15532,N_15312,N_15321);
nor U15533 (N_15533,N_15209,N_15395);
nor U15534 (N_15534,N_15220,N_15208);
xor U15535 (N_15535,N_15209,N_15333);
xnor U15536 (N_15536,N_15343,N_15271);
nand U15537 (N_15537,N_15216,N_15288);
nand U15538 (N_15538,N_15234,N_15384);
nand U15539 (N_15539,N_15376,N_15216);
or U15540 (N_15540,N_15241,N_15337);
and U15541 (N_15541,N_15364,N_15275);
nor U15542 (N_15542,N_15324,N_15386);
or U15543 (N_15543,N_15361,N_15364);
and U15544 (N_15544,N_15242,N_15378);
nand U15545 (N_15545,N_15324,N_15353);
and U15546 (N_15546,N_15210,N_15201);
xnor U15547 (N_15547,N_15247,N_15346);
xnor U15548 (N_15548,N_15276,N_15259);
and U15549 (N_15549,N_15254,N_15306);
or U15550 (N_15550,N_15260,N_15339);
nor U15551 (N_15551,N_15230,N_15395);
xor U15552 (N_15552,N_15251,N_15230);
nand U15553 (N_15553,N_15247,N_15261);
xnor U15554 (N_15554,N_15285,N_15262);
xnor U15555 (N_15555,N_15234,N_15387);
or U15556 (N_15556,N_15390,N_15341);
nand U15557 (N_15557,N_15340,N_15305);
and U15558 (N_15558,N_15370,N_15225);
xnor U15559 (N_15559,N_15311,N_15385);
and U15560 (N_15560,N_15399,N_15359);
xnor U15561 (N_15561,N_15378,N_15377);
or U15562 (N_15562,N_15382,N_15208);
or U15563 (N_15563,N_15344,N_15345);
and U15564 (N_15564,N_15200,N_15228);
or U15565 (N_15565,N_15345,N_15375);
xor U15566 (N_15566,N_15314,N_15286);
nor U15567 (N_15567,N_15325,N_15259);
or U15568 (N_15568,N_15385,N_15227);
nor U15569 (N_15569,N_15343,N_15319);
or U15570 (N_15570,N_15377,N_15267);
and U15571 (N_15571,N_15210,N_15311);
nand U15572 (N_15572,N_15338,N_15351);
and U15573 (N_15573,N_15284,N_15215);
nand U15574 (N_15574,N_15342,N_15328);
or U15575 (N_15575,N_15349,N_15325);
nand U15576 (N_15576,N_15360,N_15313);
and U15577 (N_15577,N_15397,N_15352);
or U15578 (N_15578,N_15308,N_15240);
and U15579 (N_15579,N_15382,N_15265);
nand U15580 (N_15580,N_15252,N_15265);
nor U15581 (N_15581,N_15354,N_15226);
or U15582 (N_15582,N_15238,N_15394);
nand U15583 (N_15583,N_15200,N_15204);
nand U15584 (N_15584,N_15299,N_15290);
xnor U15585 (N_15585,N_15247,N_15289);
nand U15586 (N_15586,N_15311,N_15294);
nor U15587 (N_15587,N_15318,N_15261);
nand U15588 (N_15588,N_15277,N_15337);
nand U15589 (N_15589,N_15379,N_15287);
xor U15590 (N_15590,N_15307,N_15255);
nor U15591 (N_15591,N_15337,N_15296);
or U15592 (N_15592,N_15201,N_15270);
nand U15593 (N_15593,N_15388,N_15253);
nor U15594 (N_15594,N_15314,N_15254);
or U15595 (N_15595,N_15263,N_15297);
or U15596 (N_15596,N_15241,N_15236);
and U15597 (N_15597,N_15232,N_15392);
xnor U15598 (N_15598,N_15256,N_15311);
nor U15599 (N_15599,N_15231,N_15281);
nand U15600 (N_15600,N_15432,N_15409);
xnor U15601 (N_15601,N_15537,N_15469);
nand U15602 (N_15602,N_15584,N_15587);
and U15603 (N_15603,N_15456,N_15549);
xnor U15604 (N_15604,N_15582,N_15402);
nor U15605 (N_15605,N_15408,N_15412);
nand U15606 (N_15606,N_15514,N_15555);
nand U15607 (N_15607,N_15489,N_15573);
and U15608 (N_15608,N_15506,N_15591);
and U15609 (N_15609,N_15400,N_15499);
and U15610 (N_15610,N_15422,N_15428);
xnor U15611 (N_15611,N_15517,N_15507);
and U15612 (N_15612,N_15566,N_15540);
or U15613 (N_15613,N_15501,N_15518);
nand U15614 (N_15614,N_15553,N_15521);
or U15615 (N_15615,N_15420,N_15453);
nor U15616 (N_15616,N_15597,N_15559);
xor U15617 (N_15617,N_15538,N_15568);
nand U15618 (N_15618,N_15472,N_15439);
and U15619 (N_15619,N_15438,N_15450);
or U15620 (N_15620,N_15416,N_15404);
nor U15621 (N_15621,N_15545,N_15570);
nor U15622 (N_15622,N_15505,N_15580);
nor U15623 (N_15623,N_15476,N_15547);
and U15624 (N_15624,N_15561,N_15473);
or U15625 (N_15625,N_15542,N_15579);
nor U15626 (N_15626,N_15467,N_15485);
nand U15627 (N_15627,N_15554,N_15403);
or U15628 (N_15628,N_15434,N_15433);
nand U15629 (N_15629,N_15425,N_15449);
nand U15630 (N_15630,N_15464,N_15520);
nand U15631 (N_15631,N_15497,N_15511);
or U15632 (N_15632,N_15446,N_15572);
nand U15633 (N_15633,N_15415,N_15430);
nand U15634 (N_15634,N_15503,N_15574);
or U15635 (N_15635,N_15552,N_15541);
or U15636 (N_15636,N_15411,N_15492);
and U15637 (N_15637,N_15526,N_15534);
xor U15638 (N_15638,N_15576,N_15525);
and U15639 (N_15639,N_15471,N_15444);
nand U15640 (N_15640,N_15481,N_15460);
or U15641 (N_15641,N_15483,N_15480);
and U15642 (N_15642,N_15457,N_15458);
or U15643 (N_15643,N_15583,N_15596);
nand U15644 (N_15644,N_15586,N_15590);
or U15645 (N_15645,N_15585,N_15441);
xor U15646 (N_15646,N_15593,N_15468);
and U15647 (N_15647,N_15494,N_15567);
xnor U15648 (N_15648,N_15474,N_15565);
nor U15649 (N_15649,N_15482,N_15592);
or U15650 (N_15650,N_15510,N_15571);
or U15651 (N_15651,N_15478,N_15528);
and U15652 (N_15652,N_15595,N_15410);
or U15653 (N_15653,N_15564,N_15429);
nand U15654 (N_15654,N_15533,N_15419);
and U15655 (N_15655,N_15594,N_15519);
and U15656 (N_15656,N_15431,N_15448);
nor U15657 (N_15657,N_15445,N_15466);
nor U15658 (N_15658,N_15470,N_15447);
nor U15659 (N_15659,N_15413,N_15423);
and U15660 (N_15660,N_15569,N_15527);
nor U15661 (N_15661,N_15440,N_15508);
and U15662 (N_15662,N_15509,N_15484);
and U15663 (N_15663,N_15421,N_15454);
xnor U15664 (N_15664,N_15486,N_15546);
nand U15665 (N_15665,N_15407,N_15459);
or U15666 (N_15666,N_15550,N_15502);
nand U15667 (N_15667,N_15556,N_15577);
and U15668 (N_15668,N_15475,N_15455);
or U15669 (N_15669,N_15512,N_15529);
and U15670 (N_15670,N_15451,N_15491);
and U15671 (N_15671,N_15578,N_15493);
or U15672 (N_15672,N_15436,N_15513);
xor U15673 (N_15673,N_15543,N_15548);
and U15674 (N_15674,N_15498,N_15598);
or U15675 (N_15675,N_15414,N_15599);
and U15676 (N_15676,N_15424,N_15487);
xor U15677 (N_15677,N_15524,N_15522);
nor U15678 (N_15678,N_15530,N_15465);
nand U15679 (N_15679,N_15516,N_15532);
and U15680 (N_15680,N_15452,N_15418);
nor U15681 (N_15681,N_15461,N_15462);
xnor U15682 (N_15682,N_15490,N_15535);
or U15683 (N_15683,N_15560,N_15588);
xor U15684 (N_15684,N_15463,N_15536);
nand U15685 (N_15685,N_15442,N_15479);
or U15686 (N_15686,N_15427,N_15562);
nor U15687 (N_15687,N_15435,N_15495);
nor U15688 (N_15688,N_15477,N_15496);
xnor U15689 (N_15689,N_15515,N_15544);
and U15690 (N_15690,N_15563,N_15551);
xor U15691 (N_15691,N_15443,N_15531);
nand U15692 (N_15692,N_15589,N_15539);
nand U15693 (N_15693,N_15575,N_15405);
xor U15694 (N_15694,N_15523,N_15504);
nor U15695 (N_15695,N_15581,N_15437);
nor U15696 (N_15696,N_15426,N_15557);
or U15697 (N_15697,N_15401,N_15500);
and U15698 (N_15698,N_15406,N_15558);
nand U15699 (N_15699,N_15417,N_15488);
xor U15700 (N_15700,N_15477,N_15572);
or U15701 (N_15701,N_15464,N_15541);
nor U15702 (N_15702,N_15588,N_15487);
and U15703 (N_15703,N_15564,N_15515);
nand U15704 (N_15704,N_15454,N_15522);
nand U15705 (N_15705,N_15587,N_15534);
nor U15706 (N_15706,N_15419,N_15580);
or U15707 (N_15707,N_15470,N_15588);
or U15708 (N_15708,N_15576,N_15592);
and U15709 (N_15709,N_15410,N_15590);
xnor U15710 (N_15710,N_15572,N_15448);
or U15711 (N_15711,N_15421,N_15456);
or U15712 (N_15712,N_15508,N_15480);
nor U15713 (N_15713,N_15543,N_15411);
xor U15714 (N_15714,N_15482,N_15518);
xor U15715 (N_15715,N_15563,N_15432);
or U15716 (N_15716,N_15500,N_15470);
nor U15717 (N_15717,N_15492,N_15427);
nand U15718 (N_15718,N_15586,N_15411);
and U15719 (N_15719,N_15582,N_15429);
or U15720 (N_15720,N_15488,N_15553);
and U15721 (N_15721,N_15437,N_15422);
nand U15722 (N_15722,N_15450,N_15518);
and U15723 (N_15723,N_15469,N_15499);
nand U15724 (N_15724,N_15456,N_15401);
nand U15725 (N_15725,N_15446,N_15561);
or U15726 (N_15726,N_15506,N_15412);
and U15727 (N_15727,N_15518,N_15480);
or U15728 (N_15728,N_15433,N_15518);
and U15729 (N_15729,N_15545,N_15583);
or U15730 (N_15730,N_15483,N_15428);
and U15731 (N_15731,N_15527,N_15577);
nor U15732 (N_15732,N_15589,N_15495);
and U15733 (N_15733,N_15461,N_15559);
nand U15734 (N_15734,N_15583,N_15421);
or U15735 (N_15735,N_15472,N_15573);
and U15736 (N_15736,N_15483,N_15560);
nand U15737 (N_15737,N_15422,N_15501);
and U15738 (N_15738,N_15512,N_15507);
xor U15739 (N_15739,N_15418,N_15595);
nor U15740 (N_15740,N_15552,N_15514);
or U15741 (N_15741,N_15585,N_15506);
xor U15742 (N_15742,N_15502,N_15552);
xor U15743 (N_15743,N_15402,N_15583);
or U15744 (N_15744,N_15445,N_15469);
or U15745 (N_15745,N_15570,N_15511);
or U15746 (N_15746,N_15434,N_15522);
nor U15747 (N_15747,N_15477,N_15400);
nand U15748 (N_15748,N_15445,N_15531);
nor U15749 (N_15749,N_15467,N_15407);
and U15750 (N_15750,N_15402,N_15437);
and U15751 (N_15751,N_15420,N_15469);
nor U15752 (N_15752,N_15463,N_15422);
nand U15753 (N_15753,N_15495,N_15425);
and U15754 (N_15754,N_15492,N_15410);
nand U15755 (N_15755,N_15562,N_15488);
xnor U15756 (N_15756,N_15444,N_15439);
and U15757 (N_15757,N_15506,N_15570);
and U15758 (N_15758,N_15583,N_15488);
nand U15759 (N_15759,N_15483,N_15565);
xor U15760 (N_15760,N_15476,N_15486);
xnor U15761 (N_15761,N_15598,N_15461);
nor U15762 (N_15762,N_15468,N_15515);
nor U15763 (N_15763,N_15543,N_15404);
xnor U15764 (N_15764,N_15585,N_15429);
xor U15765 (N_15765,N_15431,N_15595);
or U15766 (N_15766,N_15400,N_15510);
xnor U15767 (N_15767,N_15571,N_15538);
nand U15768 (N_15768,N_15469,N_15507);
nor U15769 (N_15769,N_15413,N_15508);
nand U15770 (N_15770,N_15588,N_15460);
xnor U15771 (N_15771,N_15582,N_15520);
or U15772 (N_15772,N_15590,N_15544);
and U15773 (N_15773,N_15526,N_15548);
and U15774 (N_15774,N_15416,N_15566);
nor U15775 (N_15775,N_15463,N_15515);
and U15776 (N_15776,N_15473,N_15599);
and U15777 (N_15777,N_15543,N_15560);
or U15778 (N_15778,N_15560,N_15531);
nor U15779 (N_15779,N_15448,N_15513);
nand U15780 (N_15780,N_15413,N_15595);
or U15781 (N_15781,N_15457,N_15545);
xnor U15782 (N_15782,N_15588,N_15500);
nor U15783 (N_15783,N_15550,N_15441);
nand U15784 (N_15784,N_15485,N_15589);
nor U15785 (N_15785,N_15479,N_15417);
and U15786 (N_15786,N_15584,N_15596);
and U15787 (N_15787,N_15460,N_15512);
and U15788 (N_15788,N_15521,N_15544);
nand U15789 (N_15789,N_15504,N_15550);
or U15790 (N_15790,N_15435,N_15445);
nand U15791 (N_15791,N_15416,N_15493);
and U15792 (N_15792,N_15525,N_15505);
xnor U15793 (N_15793,N_15437,N_15572);
nand U15794 (N_15794,N_15579,N_15543);
or U15795 (N_15795,N_15489,N_15429);
or U15796 (N_15796,N_15549,N_15502);
or U15797 (N_15797,N_15549,N_15448);
xnor U15798 (N_15798,N_15425,N_15434);
and U15799 (N_15799,N_15497,N_15553);
xnor U15800 (N_15800,N_15639,N_15683);
nand U15801 (N_15801,N_15748,N_15652);
xnor U15802 (N_15802,N_15749,N_15774);
or U15803 (N_15803,N_15750,N_15737);
nor U15804 (N_15804,N_15787,N_15667);
nor U15805 (N_15805,N_15718,N_15719);
nor U15806 (N_15806,N_15689,N_15744);
or U15807 (N_15807,N_15640,N_15691);
or U15808 (N_15808,N_15673,N_15605);
xor U15809 (N_15809,N_15740,N_15675);
and U15810 (N_15810,N_15708,N_15717);
and U15811 (N_15811,N_15734,N_15789);
or U15812 (N_15812,N_15730,N_15658);
nand U15813 (N_15813,N_15797,N_15726);
nor U15814 (N_15814,N_15761,N_15759);
and U15815 (N_15815,N_15742,N_15615);
and U15816 (N_15816,N_15745,N_15733);
nand U15817 (N_15817,N_15782,N_15692);
xnor U15818 (N_15818,N_15693,N_15649);
nand U15819 (N_15819,N_15709,N_15739);
and U15820 (N_15820,N_15765,N_15790);
nand U15821 (N_15821,N_15612,N_15636);
and U15822 (N_15822,N_15610,N_15729);
or U15823 (N_15823,N_15614,N_15713);
nor U15824 (N_15824,N_15619,N_15657);
or U15825 (N_15825,N_15766,N_15668);
or U15826 (N_15826,N_15724,N_15715);
and U15827 (N_15827,N_15677,N_15736);
and U15828 (N_15828,N_15798,N_15743);
or U15829 (N_15829,N_15635,N_15676);
and U15830 (N_15830,N_15779,N_15747);
or U15831 (N_15831,N_15776,N_15603);
nor U15832 (N_15832,N_15627,N_15613);
or U15833 (N_15833,N_15767,N_15799);
nor U15834 (N_15834,N_15775,N_15783);
or U15835 (N_15835,N_15786,N_15707);
and U15836 (N_15836,N_15638,N_15617);
or U15837 (N_15837,N_15651,N_15633);
and U15838 (N_15838,N_15792,N_15778);
nor U15839 (N_15839,N_15671,N_15780);
and U15840 (N_15840,N_15630,N_15696);
or U15841 (N_15841,N_15752,N_15662);
nand U15842 (N_15842,N_15629,N_15731);
xor U15843 (N_15843,N_15769,N_15637);
nor U15844 (N_15844,N_15757,N_15661);
or U15845 (N_15845,N_15654,N_15660);
and U15846 (N_15846,N_15681,N_15656);
nand U15847 (N_15847,N_15704,N_15723);
xor U15848 (N_15848,N_15687,N_15622);
nor U15849 (N_15849,N_15702,N_15710);
or U15850 (N_15850,N_15753,N_15760);
nand U15851 (N_15851,N_15678,N_15621);
nor U15852 (N_15852,N_15793,N_15795);
nand U15853 (N_15853,N_15646,N_15669);
xor U15854 (N_15854,N_15728,N_15722);
nand U15855 (N_15855,N_15791,N_15644);
or U15856 (N_15856,N_15694,N_15698);
and U15857 (N_15857,N_15674,N_15645);
and U15858 (N_15858,N_15631,N_15642);
nand U15859 (N_15859,N_15794,N_15624);
and U15860 (N_15860,N_15618,N_15773);
or U15861 (N_15861,N_15751,N_15714);
nor U15862 (N_15862,N_15699,N_15628);
or U15863 (N_15863,N_15626,N_15700);
and U15864 (N_15864,N_15684,N_15690);
nor U15865 (N_15865,N_15720,N_15620);
xnor U15866 (N_15866,N_15682,N_15721);
nand U15867 (N_15867,N_15788,N_15607);
or U15868 (N_15868,N_15706,N_15768);
xnor U15869 (N_15869,N_15711,N_15712);
xnor U15870 (N_15870,N_15685,N_15725);
nor U15871 (N_15871,N_15616,N_15643);
xnor U15872 (N_15872,N_15716,N_15602);
or U15873 (N_15873,N_15679,N_15705);
or U15874 (N_15874,N_15735,N_15672);
nand U15875 (N_15875,N_15701,N_15732);
nand U15876 (N_15876,N_15663,N_15697);
xor U15877 (N_15877,N_15611,N_15606);
xor U15878 (N_15878,N_15755,N_15727);
and U15879 (N_15879,N_15796,N_15688);
nand U15880 (N_15880,N_15648,N_15680);
xnor U15881 (N_15881,N_15746,N_15625);
xnor U15882 (N_15882,N_15600,N_15609);
nand U15883 (N_15883,N_15763,N_15634);
and U15884 (N_15884,N_15741,N_15653);
xnor U15885 (N_15885,N_15772,N_15686);
or U15886 (N_15886,N_15641,N_15664);
or U15887 (N_15887,N_15655,N_15785);
nand U15888 (N_15888,N_15754,N_15647);
xor U15889 (N_15889,N_15756,N_15784);
nor U15890 (N_15890,N_15777,N_15695);
or U15891 (N_15891,N_15632,N_15762);
or U15892 (N_15892,N_15738,N_15659);
and U15893 (N_15893,N_15758,N_15770);
or U15894 (N_15894,N_15703,N_15764);
or U15895 (N_15895,N_15666,N_15670);
nand U15896 (N_15896,N_15781,N_15608);
and U15897 (N_15897,N_15604,N_15771);
or U15898 (N_15898,N_15665,N_15601);
xnor U15899 (N_15899,N_15650,N_15623);
and U15900 (N_15900,N_15771,N_15701);
nor U15901 (N_15901,N_15744,N_15795);
nand U15902 (N_15902,N_15624,N_15631);
nand U15903 (N_15903,N_15673,N_15705);
nor U15904 (N_15904,N_15778,N_15714);
nor U15905 (N_15905,N_15652,N_15751);
or U15906 (N_15906,N_15609,N_15746);
nor U15907 (N_15907,N_15768,N_15691);
xnor U15908 (N_15908,N_15641,N_15786);
or U15909 (N_15909,N_15638,N_15770);
or U15910 (N_15910,N_15752,N_15727);
or U15911 (N_15911,N_15687,N_15713);
and U15912 (N_15912,N_15625,N_15638);
nor U15913 (N_15913,N_15622,N_15717);
and U15914 (N_15914,N_15720,N_15773);
nor U15915 (N_15915,N_15755,N_15669);
nor U15916 (N_15916,N_15660,N_15752);
nand U15917 (N_15917,N_15778,N_15706);
and U15918 (N_15918,N_15644,N_15643);
nor U15919 (N_15919,N_15764,N_15629);
or U15920 (N_15920,N_15643,N_15737);
nand U15921 (N_15921,N_15606,N_15717);
xnor U15922 (N_15922,N_15787,N_15719);
or U15923 (N_15923,N_15682,N_15743);
xnor U15924 (N_15924,N_15625,N_15601);
xor U15925 (N_15925,N_15765,N_15613);
and U15926 (N_15926,N_15732,N_15662);
and U15927 (N_15927,N_15706,N_15607);
and U15928 (N_15928,N_15748,N_15613);
nor U15929 (N_15929,N_15710,N_15662);
or U15930 (N_15930,N_15656,N_15673);
xnor U15931 (N_15931,N_15675,N_15622);
nand U15932 (N_15932,N_15633,N_15731);
xnor U15933 (N_15933,N_15620,N_15689);
nor U15934 (N_15934,N_15773,N_15608);
or U15935 (N_15935,N_15680,N_15772);
xnor U15936 (N_15936,N_15766,N_15777);
xor U15937 (N_15937,N_15654,N_15692);
nand U15938 (N_15938,N_15681,N_15745);
nor U15939 (N_15939,N_15663,N_15758);
nand U15940 (N_15940,N_15657,N_15666);
nor U15941 (N_15941,N_15635,N_15745);
nand U15942 (N_15942,N_15730,N_15607);
or U15943 (N_15943,N_15739,N_15699);
nand U15944 (N_15944,N_15719,N_15612);
or U15945 (N_15945,N_15630,N_15624);
and U15946 (N_15946,N_15793,N_15749);
xnor U15947 (N_15947,N_15749,N_15637);
xnor U15948 (N_15948,N_15724,N_15649);
and U15949 (N_15949,N_15640,N_15704);
xnor U15950 (N_15950,N_15703,N_15640);
nand U15951 (N_15951,N_15723,N_15667);
xnor U15952 (N_15952,N_15666,N_15620);
xnor U15953 (N_15953,N_15741,N_15703);
nor U15954 (N_15954,N_15758,N_15658);
xor U15955 (N_15955,N_15792,N_15798);
or U15956 (N_15956,N_15755,N_15766);
or U15957 (N_15957,N_15775,N_15749);
xor U15958 (N_15958,N_15609,N_15625);
xnor U15959 (N_15959,N_15600,N_15752);
or U15960 (N_15960,N_15685,N_15717);
xor U15961 (N_15961,N_15627,N_15674);
or U15962 (N_15962,N_15759,N_15750);
xor U15963 (N_15963,N_15641,N_15769);
nand U15964 (N_15964,N_15643,N_15673);
and U15965 (N_15965,N_15717,N_15744);
nor U15966 (N_15966,N_15653,N_15650);
xnor U15967 (N_15967,N_15769,N_15702);
xor U15968 (N_15968,N_15742,N_15632);
nor U15969 (N_15969,N_15724,N_15609);
xor U15970 (N_15970,N_15707,N_15698);
nor U15971 (N_15971,N_15745,N_15688);
or U15972 (N_15972,N_15659,N_15720);
nor U15973 (N_15973,N_15718,N_15713);
nand U15974 (N_15974,N_15792,N_15724);
and U15975 (N_15975,N_15765,N_15650);
and U15976 (N_15976,N_15701,N_15747);
or U15977 (N_15977,N_15708,N_15770);
or U15978 (N_15978,N_15647,N_15697);
or U15979 (N_15979,N_15632,N_15702);
and U15980 (N_15980,N_15602,N_15752);
nand U15981 (N_15981,N_15678,N_15713);
xnor U15982 (N_15982,N_15720,N_15641);
and U15983 (N_15983,N_15641,N_15768);
xor U15984 (N_15984,N_15638,N_15604);
xnor U15985 (N_15985,N_15655,N_15611);
nand U15986 (N_15986,N_15698,N_15668);
and U15987 (N_15987,N_15698,N_15704);
nand U15988 (N_15988,N_15725,N_15615);
nor U15989 (N_15989,N_15649,N_15752);
nand U15990 (N_15990,N_15708,N_15628);
or U15991 (N_15991,N_15647,N_15698);
and U15992 (N_15992,N_15674,N_15776);
or U15993 (N_15993,N_15613,N_15779);
nand U15994 (N_15994,N_15669,N_15649);
and U15995 (N_15995,N_15722,N_15783);
and U15996 (N_15996,N_15730,N_15619);
nand U15997 (N_15997,N_15604,N_15731);
or U15998 (N_15998,N_15719,N_15621);
nor U15999 (N_15999,N_15762,N_15706);
xor U16000 (N_16000,N_15915,N_15828);
nand U16001 (N_16001,N_15999,N_15889);
nand U16002 (N_16002,N_15904,N_15948);
or U16003 (N_16003,N_15928,N_15805);
nor U16004 (N_16004,N_15975,N_15842);
nand U16005 (N_16005,N_15987,N_15818);
or U16006 (N_16006,N_15868,N_15974);
and U16007 (N_16007,N_15838,N_15959);
nor U16008 (N_16008,N_15991,N_15916);
xnor U16009 (N_16009,N_15854,N_15874);
and U16010 (N_16010,N_15850,N_15815);
or U16011 (N_16011,N_15851,N_15953);
nand U16012 (N_16012,N_15812,N_15907);
xor U16013 (N_16013,N_15962,N_15871);
xnor U16014 (N_16014,N_15971,N_15813);
or U16015 (N_16015,N_15817,N_15966);
nand U16016 (N_16016,N_15964,N_15914);
and U16017 (N_16017,N_15943,N_15827);
nor U16018 (N_16018,N_15908,N_15918);
nor U16019 (N_16019,N_15855,N_15940);
xor U16020 (N_16020,N_15963,N_15806);
xor U16021 (N_16021,N_15829,N_15988);
xnor U16022 (N_16022,N_15899,N_15937);
nor U16023 (N_16023,N_15882,N_15996);
nand U16024 (N_16024,N_15826,N_15912);
nor U16025 (N_16025,N_15867,N_15824);
xor U16026 (N_16026,N_15832,N_15910);
nand U16027 (N_16027,N_15917,N_15836);
or U16028 (N_16028,N_15969,N_15950);
nand U16029 (N_16029,N_15891,N_15835);
or U16030 (N_16030,N_15994,N_15906);
xor U16031 (N_16031,N_15861,N_15927);
and U16032 (N_16032,N_15951,N_15905);
and U16033 (N_16033,N_15923,N_15968);
nor U16034 (N_16034,N_15848,N_15841);
xor U16035 (N_16035,N_15958,N_15839);
and U16036 (N_16036,N_15955,N_15823);
nor U16037 (N_16037,N_15981,N_15877);
or U16038 (N_16038,N_15886,N_15941);
and U16039 (N_16039,N_15863,N_15894);
and U16040 (N_16040,N_15849,N_15972);
nand U16041 (N_16041,N_15961,N_15831);
xnor U16042 (N_16042,N_15881,N_15834);
xor U16043 (N_16043,N_15847,N_15960);
and U16044 (N_16044,N_15909,N_15935);
nor U16045 (N_16045,N_15872,N_15875);
and U16046 (N_16046,N_15985,N_15986);
or U16047 (N_16047,N_15807,N_15819);
or U16048 (N_16048,N_15913,N_15803);
nand U16049 (N_16049,N_15862,N_15938);
or U16050 (N_16050,N_15885,N_15924);
xor U16051 (N_16051,N_15995,N_15825);
xor U16052 (N_16052,N_15814,N_15840);
nand U16053 (N_16053,N_15957,N_15998);
or U16054 (N_16054,N_15952,N_15865);
xor U16055 (N_16055,N_15859,N_15900);
or U16056 (N_16056,N_15926,N_15852);
xor U16057 (N_16057,N_15833,N_15801);
or U16058 (N_16058,N_15808,N_15934);
or U16059 (N_16059,N_15897,N_15880);
nor U16060 (N_16060,N_15816,N_15920);
or U16061 (N_16061,N_15980,N_15903);
xnor U16062 (N_16062,N_15933,N_15878);
xnor U16063 (N_16063,N_15876,N_15919);
and U16064 (N_16064,N_15967,N_15896);
xor U16065 (N_16065,N_15947,N_15984);
nand U16066 (N_16066,N_15921,N_15979);
or U16067 (N_16067,N_15883,N_15932);
nor U16068 (N_16068,N_15802,N_15978);
or U16069 (N_16069,N_15911,N_15990);
nand U16070 (N_16070,N_15997,N_15965);
and U16071 (N_16071,N_15857,N_15949);
and U16072 (N_16072,N_15892,N_15869);
nand U16073 (N_16073,N_15946,N_15929);
nor U16074 (N_16074,N_15989,N_15890);
and U16075 (N_16075,N_15800,N_15804);
xnor U16076 (N_16076,N_15809,N_15837);
and U16077 (N_16077,N_15895,N_15843);
nand U16078 (N_16078,N_15866,N_15884);
nor U16079 (N_16079,N_15922,N_15956);
or U16080 (N_16080,N_15939,N_15870);
xor U16081 (N_16081,N_15973,N_15853);
xor U16082 (N_16082,N_15888,N_15970);
nor U16083 (N_16083,N_15864,N_15820);
nand U16084 (N_16084,N_15931,N_15976);
or U16085 (N_16085,N_15898,N_15811);
nor U16086 (N_16086,N_15810,N_15992);
nor U16087 (N_16087,N_15936,N_15942);
and U16088 (N_16088,N_15983,N_15944);
or U16089 (N_16089,N_15930,N_15860);
nor U16090 (N_16090,N_15993,N_15977);
xnor U16091 (N_16091,N_15982,N_15858);
nor U16092 (N_16092,N_15954,N_15902);
nand U16093 (N_16093,N_15879,N_15844);
nor U16094 (N_16094,N_15845,N_15822);
nand U16095 (N_16095,N_15846,N_15901);
or U16096 (N_16096,N_15925,N_15830);
and U16097 (N_16097,N_15873,N_15887);
and U16098 (N_16098,N_15821,N_15856);
nand U16099 (N_16099,N_15893,N_15945);
or U16100 (N_16100,N_15990,N_15925);
nor U16101 (N_16101,N_15962,N_15979);
or U16102 (N_16102,N_15980,N_15871);
xnor U16103 (N_16103,N_15803,N_15957);
xor U16104 (N_16104,N_15970,N_15831);
and U16105 (N_16105,N_15908,N_15898);
nor U16106 (N_16106,N_15911,N_15909);
and U16107 (N_16107,N_15856,N_15823);
or U16108 (N_16108,N_15890,N_15874);
nor U16109 (N_16109,N_15995,N_15984);
xnor U16110 (N_16110,N_15846,N_15917);
and U16111 (N_16111,N_15841,N_15924);
xor U16112 (N_16112,N_15831,N_15909);
and U16113 (N_16113,N_15865,N_15870);
nor U16114 (N_16114,N_15972,N_15845);
xor U16115 (N_16115,N_15969,N_15835);
and U16116 (N_16116,N_15980,N_15861);
and U16117 (N_16117,N_15877,N_15988);
nand U16118 (N_16118,N_15863,N_15855);
xor U16119 (N_16119,N_15971,N_15943);
nor U16120 (N_16120,N_15901,N_15939);
and U16121 (N_16121,N_15893,N_15921);
nand U16122 (N_16122,N_15880,N_15965);
and U16123 (N_16123,N_15934,N_15863);
xor U16124 (N_16124,N_15917,N_15963);
xor U16125 (N_16125,N_15904,N_15811);
xor U16126 (N_16126,N_15870,N_15867);
and U16127 (N_16127,N_15895,N_15868);
nand U16128 (N_16128,N_15812,N_15904);
nand U16129 (N_16129,N_15923,N_15972);
nand U16130 (N_16130,N_15870,N_15918);
nor U16131 (N_16131,N_15845,N_15958);
xnor U16132 (N_16132,N_15923,N_15858);
nand U16133 (N_16133,N_15995,N_15981);
nand U16134 (N_16134,N_15836,N_15973);
xor U16135 (N_16135,N_15948,N_15816);
nor U16136 (N_16136,N_15823,N_15865);
nand U16137 (N_16137,N_15896,N_15828);
nand U16138 (N_16138,N_15883,N_15823);
nand U16139 (N_16139,N_15928,N_15942);
and U16140 (N_16140,N_15859,N_15883);
xor U16141 (N_16141,N_15942,N_15864);
or U16142 (N_16142,N_15810,N_15964);
and U16143 (N_16143,N_15811,N_15934);
or U16144 (N_16144,N_15831,N_15967);
nand U16145 (N_16145,N_15829,N_15892);
xnor U16146 (N_16146,N_15970,N_15899);
xnor U16147 (N_16147,N_15847,N_15808);
nor U16148 (N_16148,N_15940,N_15877);
nand U16149 (N_16149,N_15813,N_15808);
or U16150 (N_16150,N_15879,N_15815);
nand U16151 (N_16151,N_15945,N_15818);
nor U16152 (N_16152,N_15888,N_15948);
and U16153 (N_16153,N_15885,N_15806);
and U16154 (N_16154,N_15801,N_15960);
and U16155 (N_16155,N_15847,N_15871);
nor U16156 (N_16156,N_15829,N_15970);
and U16157 (N_16157,N_15835,N_15876);
and U16158 (N_16158,N_15837,N_15925);
nor U16159 (N_16159,N_15879,N_15857);
and U16160 (N_16160,N_15931,N_15816);
and U16161 (N_16161,N_15992,N_15888);
nor U16162 (N_16162,N_15827,N_15821);
and U16163 (N_16163,N_15812,N_15921);
nor U16164 (N_16164,N_15989,N_15955);
or U16165 (N_16165,N_15997,N_15956);
nand U16166 (N_16166,N_15979,N_15978);
and U16167 (N_16167,N_15932,N_15907);
nand U16168 (N_16168,N_15835,N_15821);
or U16169 (N_16169,N_15968,N_15832);
xnor U16170 (N_16170,N_15811,N_15855);
and U16171 (N_16171,N_15833,N_15880);
and U16172 (N_16172,N_15871,N_15872);
xor U16173 (N_16173,N_15977,N_15999);
and U16174 (N_16174,N_15843,N_15804);
xor U16175 (N_16175,N_15894,N_15837);
nor U16176 (N_16176,N_15984,N_15838);
nand U16177 (N_16177,N_15937,N_15968);
nor U16178 (N_16178,N_15930,N_15973);
nor U16179 (N_16179,N_15909,N_15993);
or U16180 (N_16180,N_15930,N_15994);
or U16181 (N_16181,N_15916,N_15951);
xnor U16182 (N_16182,N_15993,N_15989);
nor U16183 (N_16183,N_15965,N_15892);
and U16184 (N_16184,N_15928,N_15967);
nor U16185 (N_16185,N_15993,N_15830);
nor U16186 (N_16186,N_15905,N_15803);
or U16187 (N_16187,N_15846,N_15958);
or U16188 (N_16188,N_15868,N_15987);
nor U16189 (N_16189,N_15842,N_15929);
nor U16190 (N_16190,N_15915,N_15893);
xnor U16191 (N_16191,N_15927,N_15993);
xnor U16192 (N_16192,N_15846,N_15926);
and U16193 (N_16193,N_15825,N_15914);
or U16194 (N_16194,N_15819,N_15919);
xor U16195 (N_16195,N_15804,N_15828);
nand U16196 (N_16196,N_15939,N_15932);
nor U16197 (N_16197,N_15965,N_15979);
and U16198 (N_16198,N_15985,N_15815);
or U16199 (N_16199,N_15807,N_15865);
or U16200 (N_16200,N_16143,N_16138);
nand U16201 (N_16201,N_16198,N_16156);
or U16202 (N_16202,N_16136,N_16082);
nand U16203 (N_16203,N_16161,N_16030);
nor U16204 (N_16204,N_16053,N_16023);
xnor U16205 (N_16205,N_16058,N_16095);
or U16206 (N_16206,N_16061,N_16105);
nand U16207 (N_16207,N_16078,N_16113);
xor U16208 (N_16208,N_16024,N_16182);
nand U16209 (N_16209,N_16016,N_16097);
nand U16210 (N_16210,N_16141,N_16004);
xnor U16211 (N_16211,N_16149,N_16032);
and U16212 (N_16212,N_16154,N_16017);
or U16213 (N_16213,N_16140,N_16075);
or U16214 (N_16214,N_16002,N_16015);
nor U16215 (N_16215,N_16196,N_16035);
nand U16216 (N_16216,N_16081,N_16114);
nand U16217 (N_16217,N_16162,N_16009);
nor U16218 (N_16218,N_16008,N_16070);
or U16219 (N_16219,N_16067,N_16028);
or U16220 (N_16220,N_16007,N_16103);
nor U16221 (N_16221,N_16124,N_16107);
and U16222 (N_16222,N_16066,N_16025);
xor U16223 (N_16223,N_16014,N_16049);
nor U16224 (N_16224,N_16121,N_16189);
nor U16225 (N_16225,N_16045,N_16171);
and U16226 (N_16226,N_16133,N_16115);
nor U16227 (N_16227,N_16047,N_16064);
xor U16228 (N_16228,N_16089,N_16038);
and U16229 (N_16229,N_16037,N_16046);
nor U16230 (N_16230,N_16057,N_16164);
or U16231 (N_16231,N_16163,N_16068);
xnor U16232 (N_16232,N_16001,N_16056);
or U16233 (N_16233,N_16010,N_16074);
and U16234 (N_16234,N_16191,N_16181);
nor U16235 (N_16235,N_16020,N_16022);
nand U16236 (N_16236,N_16117,N_16073);
nand U16237 (N_16237,N_16027,N_16160);
nand U16238 (N_16238,N_16013,N_16118);
nor U16239 (N_16239,N_16085,N_16019);
or U16240 (N_16240,N_16129,N_16029);
nand U16241 (N_16241,N_16060,N_16135);
and U16242 (N_16242,N_16090,N_16127);
and U16243 (N_16243,N_16031,N_16192);
nor U16244 (N_16244,N_16128,N_16176);
nor U16245 (N_16245,N_16100,N_16165);
or U16246 (N_16246,N_16072,N_16190);
and U16247 (N_16247,N_16083,N_16033);
and U16248 (N_16248,N_16173,N_16126);
and U16249 (N_16249,N_16087,N_16144);
and U16250 (N_16250,N_16018,N_16119);
or U16251 (N_16251,N_16186,N_16112);
or U16252 (N_16252,N_16051,N_16077);
and U16253 (N_16253,N_16000,N_16054);
nor U16254 (N_16254,N_16110,N_16188);
xor U16255 (N_16255,N_16088,N_16079);
nand U16256 (N_16256,N_16134,N_16101);
and U16257 (N_16257,N_16034,N_16178);
nand U16258 (N_16258,N_16197,N_16116);
nand U16259 (N_16259,N_16169,N_16183);
or U16260 (N_16260,N_16142,N_16042);
nand U16261 (N_16261,N_16125,N_16076);
xnor U16262 (N_16262,N_16145,N_16153);
and U16263 (N_16263,N_16052,N_16059);
xnor U16264 (N_16264,N_16040,N_16044);
nor U16265 (N_16265,N_16177,N_16166);
or U16266 (N_16266,N_16055,N_16096);
or U16267 (N_16267,N_16012,N_16131);
nand U16268 (N_16268,N_16065,N_16102);
nor U16269 (N_16269,N_16109,N_16194);
nor U16270 (N_16270,N_16043,N_16167);
xnor U16271 (N_16271,N_16174,N_16108);
and U16272 (N_16272,N_16104,N_16021);
nor U16273 (N_16273,N_16111,N_16069);
and U16274 (N_16274,N_16179,N_16006);
or U16275 (N_16275,N_16184,N_16193);
xnor U16276 (N_16276,N_16084,N_16147);
or U16277 (N_16277,N_16130,N_16152);
and U16278 (N_16278,N_16172,N_16011);
xnor U16279 (N_16279,N_16063,N_16048);
nand U16280 (N_16280,N_16139,N_16170);
nor U16281 (N_16281,N_16195,N_16180);
xnor U16282 (N_16282,N_16041,N_16148);
nor U16283 (N_16283,N_16093,N_16062);
xor U16284 (N_16284,N_16098,N_16091);
nand U16285 (N_16285,N_16150,N_16099);
xnor U16286 (N_16286,N_16080,N_16175);
and U16287 (N_16287,N_16159,N_16151);
nand U16288 (N_16288,N_16132,N_16094);
and U16289 (N_16289,N_16036,N_16026);
and U16290 (N_16290,N_16137,N_16106);
nor U16291 (N_16291,N_16155,N_16185);
nor U16292 (N_16292,N_16123,N_16157);
and U16293 (N_16293,N_16187,N_16071);
or U16294 (N_16294,N_16199,N_16158);
or U16295 (N_16295,N_16039,N_16005);
nand U16296 (N_16296,N_16086,N_16122);
nor U16297 (N_16297,N_16120,N_16050);
or U16298 (N_16298,N_16146,N_16168);
and U16299 (N_16299,N_16003,N_16092);
nor U16300 (N_16300,N_16125,N_16041);
or U16301 (N_16301,N_16071,N_16046);
and U16302 (N_16302,N_16194,N_16117);
xor U16303 (N_16303,N_16153,N_16163);
xnor U16304 (N_16304,N_16038,N_16058);
or U16305 (N_16305,N_16098,N_16093);
and U16306 (N_16306,N_16074,N_16075);
and U16307 (N_16307,N_16018,N_16189);
xor U16308 (N_16308,N_16134,N_16023);
or U16309 (N_16309,N_16116,N_16091);
nor U16310 (N_16310,N_16120,N_16063);
xnor U16311 (N_16311,N_16065,N_16183);
or U16312 (N_16312,N_16143,N_16126);
nor U16313 (N_16313,N_16043,N_16084);
or U16314 (N_16314,N_16069,N_16053);
nor U16315 (N_16315,N_16008,N_16129);
and U16316 (N_16316,N_16130,N_16087);
nor U16317 (N_16317,N_16078,N_16059);
nor U16318 (N_16318,N_16152,N_16019);
and U16319 (N_16319,N_16181,N_16135);
nor U16320 (N_16320,N_16021,N_16177);
nand U16321 (N_16321,N_16100,N_16174);
and U16322 (N_16322,N_16151,N_16090);
or U16323 (N_16323,N_16005,N_16169);
and U16324 (N_16324,N_16183,N_16164);
nand U16325 (N_16325,N_16111,N_16015);
nor U16326 (N_16326,N_16099,N_16097);
nand U16327 (N_16327,N_16034,N_16035);
and U16328 (N_16328,N_16127,N_16151);
and U16329 (N_16329,N_16055,N_16103);
nand U16330 (N_16330,N_16087,N_16024);
or U16331 (N_16331,N_16134,N_16126);
nand U16332 (N_16332,N_16062,N_16018);
xor U16333 (N_16333,N_16034,N_16183);
nor U16334 (N_16334,N_16035,N_16091);
or U16335 (N_16335,N_16198,N_16054);
xor U16336 (N_16336,N_16194,N_16001);
nand U16337 (N_16337,N_16046,N_16135);
and U16338 (N_16338,N_16145,N_16047);
nor U16339 (N_16339,N_16133,N_16156);
nand U16340 (N_16340,N_16146,N_16123);
nor U16341 (N_16341,N_16159,N_16145);
or U16342 (N_16342,N_16056,N_16086);
nor U16343 (N_16343,N_16011,N_16028);
and U16344 (N_16344,N_16074,N_16040);
or U16345 (N_16345,N_16132,N_16007);
or U16346 (N_16346,N_16097,N_16157);
nor U16347 (N_16347,N_16121,N_16168);
nor U16348 (N_16348,N_16169,N_16184);
nand U16349 (N_16349,N_16116,N_16016);
xnor U16350 (N_16350,N_16081,N_16157);
nand U16351 (N_16351,N_16080,N_16038);
or U16352 (N_16352,N_16064,N_16160);
or U16353 (N_16353,N_16101,N_16063);
or U16354 (N_16354,N_16006,N_16132);
or U16355 (N_16355,N_16044,N_16120);
nand U16356 (N_16356,N_16168,N_16039);
xor U16357 (N_16357,N_16187,N_16061);
or U16358 (N_16358,N_16141,N_16150);
nand U16359 (N_16359,N_16118,N_16167);
or U16360 (N_16360,N_16014,N_16168);
xor U16361 (N_16361,N_16049,N_16035);
and U16362 (N_16362,N_16198,N_16152);
and U16363 (N_16363,N_16064,N_16103);
xnor U16364 (N_16364,N_16106,N_16131);
xnor U16365 (N_16365,N_16193,N_16131);
and U16366 (N_16366,N_16173,N_16097);
nor U16367 (N_16367,N_16029,N_16119);
and U16368 (N_16368,N_16028,N_16033);
nand U16369 (N_16369,N_16160,N_16187);
xnor U16370 (N_16370,N_16149,N_16043);
or U16371 (N_16371,N_16027,N_16199);
xnor U16372 (N_16372,N_16008,N_16144);
xnor U16373 (N_16373,N_16021,N_16091);
and U16374 (N_16374,N_16045,N_16040);
nor U16375 (N_16375,N_16192,N_16140);
and U16376 (N_16376,N_16014,N_16108);
nand U16377 (N_16377,N_16052,N_16184);
nand U16378 (N_16378,N_16036,N_16060);
or U16379 (N_16379,N_16050,N_16017);
nor U16380 (N_16380,N_16141,N_16166);
and U16381 (N_16381,N_16135,N_16147);
nor U16382 (N_16382,N_16059,N_16123);
nand U16383 (N_16383,N_16085,N_16043);
or U16384 (N_16384,N_16161,N_16136);
nand U16385 (N_16385,N_16179,N_16170);
and U16386 (N_16386,N_16090,N_16100);
or U16387 (N_16387,N_16147,N_16040);
nand U16388 (N_16388,N_16186,N_16103);
xor U16389 (N_16389,N_16016,N_16192);
and U16390 (N_16390,N_16156,N_16041);
or U16391 (N_16391,N_16160,N_16195);
nor U16392 (N_16392,N_16191,N_16028);
nor U16393 (N_16393,N_16180,N_16081);
xor U16394 (N_16394,N_16042,N_16195);
and U16395 (N_16395,N_16101,N_16190);
nor U16396 (N_16396,N_16065,N_16115);
xnor U16397 (N_16397,N_16176,N_16143);
and U16398 (N_16398,N_16022,N_16188);
nor U16399 (N_16399,N_16031,N_16145);
nand U16400 (N_16400,N_16273,N_16396);
and U16401 (N_16401,N_16327,N_16237);
or U16402 (N_16402,N_16302,N_16323);
or U16403 (N_16403,N_16317,N_16384);
xor U16404 (N_16404,N_16374,N_16314);
or U16405 (N_16405,N_16257,N_16263);
or U16406 (N_16406,N_16255,N_16256);
xnor U16407 (N_16407,N_16217,N_16218);
nand U16408 (N_16408,N_16297,N_16215);
xor U16409 (N_16409,N_16346,N_16310);
xnor U16410 (N_16410,N_16348,N_16210);
nor U16411 (N_16411,N_16363,N_16253);
or U16412 (N_16412,N_16324,N_16308);
xnor U16413 (N_16413,N_16204,N_16219);
or U16414 (N_16414,N_16393,N_16392);
nand U16415 (N_16415,N_16272,N_16258);
nor U16416 (N_16416,N_16207,N_16252);
xor U16417 (N_16417,N_16389,N_16285);
or U16418 (N_16418,N_16360,N_16288);
or U16419 (N_16419,N_16300,N_16343);
and U16420 (N_16420,N_16330,N_16299);
xor U16421 (N_16421,N_16292,N_16245);
or U16422 (N_16422,N_16301,N_16345);
xor U16423 (N_16423,N_16304,N_16238);
or U16424 (N_16424,N_16376,N_16329);
nor U16425 (N_16425,N_16201,N_16313);
and U16426 (N_16426,N_16349,N_16391);
nor U16427 (N_16427,N_16373,N_16259);
nor U16428 (N_16428,N_16286,N_16298);
nand U16429 (N_16429,N_16395,N_16332);
nand U16430 (N_16430,N_16249,N_16228);
nand U16431 (N_16431,N_16351,N_16379);
or U16432 (N_16432,N_16388,N_16338);
xnor U16433 (N_16433,N_16326,N_16251);
xnor U16434 (N_16434,N_16377,N_16381);
nand U16435 (N_16435,N_16365,N_16387);
or U16436 (N_16436,N_16340,N_16293);
nor U16437 (N_16437,N_16331,N_16295);
or U16438 (N_16438,N_16378,N_16276);
xor U16439 (N_16439,N_16235,N_16320);
nand U16440 (N_16440,N_16341,N_16278);
and U16441 (N_16441,N_16335,N_16397);
nor U16442 (N_16442,N_16352,N_16386);
or U16443 (N_16443,N_16268,N_16284);
nor U16444 (N_16444,N_16282,N_16208);
nor U16445 (N_16445,N_16220,N_16281);
nor U16446 (N_16446,N_16354,N_16312);
xnor U16447 (N_16447,N_16342,N_16212);
nand U16448 (N_16448,N_16309,N_16280);
nor U16449 (N_16449,N_16380,N_16367);
nand U16450 (N_16450,N_16226,N_16221);
xnor U16451 (N_16451,N_16321,N_16216);
xor U16452 (N_16452,N_16232,N_16394);
xnor U16453 (N_16453,N_16356,N_16369);
nand U16454 (N_16454,N_16211,N_16372);
nand U16455 (N_16455,N_16224,N_16230);
xnor U16456 (N_16456,N_16291,N_16289);
xor U16457 (N_16457,N_16279,N_16205);
nor U16458 (N_16458,N_16315,N_16385);
nand U16459 (N_16459,N_16262,N_16311);
or U16460 (N_16460,N_16347,N_16260);
or U16461 (N_16461,N_16333,N_16294);
xnor U16462 (N_16462,N_16261,N_16274);
nor U16463 (N_16463,N_16240,N_16206);
xor U16464 (N_16464,N_16334,N_16366);
xor U16465 (N_16465,N_16318,N_16227);
and U16466 (N_16466,N_16209,N_16271);
or U16467 (N_16467,N_16339,N_16350);
nor U16468 (N_16468,N_16390,N_16359);
xor U16469 (N_16469,N_16364,N_16242);
nor U16470 (N_16470,N_16306,N_16244);
xnor U16471 (N_16471,N_16353,N_16275);
or U16472 (N_16472,N_16277,N_16248);
nand U16473 (N_16473,N_16358,N_16241);
nor U16474 (N_16474,N_16213,N_16305);
and U16475 (N_16475,N_16371,N_16319);
or U16476 (N_16476,N_16246,N_16265);
nor U16477 (N_16477,N_16283,N_16325);
and U16478 (N_16478,N_16266,N_16344);
or U16479 (N_16479,N_16382,N_16370);
xnor U16480 (N_16480,N_16355,N_16336);
xnor U16481 (N_16481,N_16264,N_16269);
nand U16482 (N_16482,N_16214,N_16222);
and U16483 (N_16483,N_16236,N_16399);
and U16484 (N_16484,N_16239,N_16322);
nor U16485 (N_16485,N_16375,N_16398);
xor U16486 (N_16486,N_16231,N_16233);
nor U16487 (N_16487,N_16247,N_16296);
nor U16488 (N_16488,N_16234,N_16229);
or U16489 (N_16489,N_16243,N_16361);
or U16490 (N_16490,N_16287,N_16307);
xnor U16491 (N_16491,N_16290,N_16383);
nor U16492 (N_16492,N_16337,N_16202);
and U16493 (N_16493,N_16303,N_16267);
xnor U16494 (N_16494,N_16357,N_16368);
nand U16495 (N_16495,N_16225,N_16250);
nand U16496 (N_16496,N_16203,N_16316);
and U16497 (N_16497,N_16328,N_16223);
nand U16498 (N_16498,N_16254,N_16270);
nand U16499 (N_16499,N_16200,N_16362);
or U16500 (N_16500,N_16314,N_16368);
and U16501 (N_16501,N_16304,N_16393);
or U16502 (N_16502,N_16335,N_16247);
nor U16503 (N_16503,N_16212,N_16206);
nor U16504 (N_16504,N_16215,N_16239);
or U16505 (N_16505,N_16367,N_16291);
nor U16506 (N_16506,N_16222,N_16302);
and U16507 (N_16507,N_16356,N_16319);
xnor U16508 (N_16508,N_16252,N_16238);
or U16509 (N_16509,N_16321,N_16381);
or U16510 (N_16510,N_16389,N_16275);
xnor U16511 (N_16511,N_16387,N_16330);
and U16512 (N_16512,N_16380,N_16253);
and U16513 (N_16513,N_16301,N_16237);
and U16514 (N_16514,N_16209,N_16391);
and U16515 (N_16515,N_16225,N_16207);
and U16516 (N_16516,N_16208,N_16259);
and U16517 (N_16517,N_16399,N_16361);
and U16518 (N_16518,N_16211,N_16309);
xnor U16519 (N_16519,N_16346,N_16364);
xor U16520 (N_16520,N_16248,N_16361);
and U16521 (N_16521,N_16334,N_16374);
nand U16522 (N_16522,N_16207,N_16258);
or U16523 (N_16523,N_16238,N_16203);
nand U16524 (N_16524,N_16270,N_16375);
xnor U16525 (N_16525,N_16382,N_16394);
nand U16526 (N_16526,N_16262,N_16309);
nor U16527 (N_16527,N_16269,N_16330);
and U16528 (N_16528,N_16284,N_16277);
nand U16529 (N_16529,N_16394,N_16351);
nand U16530 (N_16530,N_16365,N_16235);
or U16531 (N_16531,N_16287,N_16313);
nor U16532 (N_16532,N_16377,N_16334);
xnor U16533 (N_16533,N_16378,N_16240);
nand U16534 (N_16534,N_16393,N_16206);
xor U16535 (N_16535,N_16252,N_16255);
nor U16536 (N_16536,N_16202,N_16274);
and U16537 (N_16537,N_16305,N_16227);
xnor U16538 (N_16538,N_16378,N_16271);
and U16539 (N_16539,N_16345,N_16203);
nand U16540 (N_16540,N_16282,N_16292);
nor U16541 (N_16541,N_16345,N_16242);
and U16542 (N_16542,N_16216,N_16325);
or U16543 (N_16543,N_16261,N_16245);
nor U16544 (N_16544,N_16368,N_16287);
nand U16545 (N_16545,N_16399,N_16226);
or U16546 (N_16546,N_16335,N_16317);
nand U16547 (N_16547,N_16300,N_16273);
and U16548 (N_16548,N_16351,N_16330);
nor U16549 (N_16549,N_16298,N_16294);
nand U16550 (N_16550,N_16265,N_16278);
nand U16551 (N_16551,N_16260,N_16277);
nor U16552 (N_16552,N_16240,N_16387);
and U16553 (N_16553,N_16200,N_16386);
nor U16554 (N_16554,N_16311,N_16279);
and U16555 (N_16555,N_16397,N_16388);
xor U16556 (N_16556,N_16282,N_16231);
xnor U16557 (N_16557,N_16271,N_16277);
xor U16558 (N_16558,N_16382,N_16397);
and U16559 (N_16559,N_16358,N_16345);
or U16560 (N_16560,N_16239,N_16296);
nand U16561 (N_16561,N_16230,N_16384);
nor U16562 (N_16562,N_16270,N_16261);
nand U16563 (N_16563,N_16287,N_16365);
nand U16564 (N_16564,N_16263,N_16234);
xnor U16565 (N_16565,N_16256,N_16287);
nand U16566 (N_16566,N_16241,N_16383);
or U16567 (N_16567,N_16317,N_16208);
or U16568 (N_16568,N_16398,N_16355);
xor U16569 (N_16569,N_16246,N_16357);
nand U16570 (N_16570,N_16284,N_16382);
nor U16571 (N_16571,N_16349,N_16326);
or U16572 (N_16572,N_16347,N_16319);
nor U16573 (N_16573,N_16227,N_16368);
xor U16574 (N_16574,N_16224,N_16239);
or U16575 (N_16575,N_16236,N_16290);
xnor U16576 (N_16576,N_16354,N_16223);
or U16577 (N_16577,N_16307,N_16248);
or U16578 (N_16578,N_16250,N_16208);
or U16579 (N_16579,N_16339,N_16290);
and U16580 (N_16580,N_16283,N_16284);
nor U16581 (N_16581,N_16314,N_16321);
nor U16582 (N_16582,N_16328,N_16353);
and U16583 (N_16583,N_16320,N_16303);
xnor U16584 (N_16584,N_16308,N_16353);
and U16585 (N_16585,N_16375,N_16305);
xnor U16586 (N_16586,N_16229,N_16373);
and U16587 (N_16587,N_16383,N_16267);
and U16588 (N_16588,N_16330,N_16304);
nand U16589 (N_16589,N_16347,N_16269);
and U16590 (N_16590,N_16395,N_16272);
and U16591 (N_16591,N_16346,N_16259);
nor U16592 (N_16592,N_16254,N_16338);
nand U16593 (N_16593,N_16297,N_16206);
nand U16594 (N_16594,N_16369,N_16225);
or U16595 (N_16595,N_16358,N_16330);
or U16596 (N_16596,N_16399,N_16258);
or U16597 (N_16597,N_16219,N_16353);
nor U16598 (N_16598,N_16393,N_16370);
or U16599 (N_16599,N_16239,N_16207);
nand U16600 (N_16600,N_16425,N_16413);
and U16601 (N_16601,N_16529,N_16436);
and U16602 (N_16602,N_16426,N_16499);
nand U16603 (N_16603,N_16581,N_16420);
or U16604 (N_16604,N_16447,N_16592);
and U16605 (N_16605,N_16500,N_16411);
or U16606 (N_16606,N_16463,N_16518);
or U16607 (N_16607,N_16474,N_16594);
nand U16608 (N_16608,N_16487,N_16446);
nand U16609 (N_16609,N_16403,N_16492);
and U16610 (N_16610,N_16458,N_16490);
or U16611 (N_16611,N_16464,N_16541);
or U16612 (N_16612,N_16596,N_16408);
xor U16613 (N_16613,N_16489,N_16442);
nor U16614 (N_16614,N_16506,N_16514);
xnor U16615 (N_16615,N_16418,N_16577);
and U16616 (N_16616,N_16488,N_16575);
nand U16617 (N_16617,N_16445,N_16502);
or U16618 (N_16618,N_16407,N_16462);
xnor U16619 (N_16619,N_16466,N_16497);
xor U16620 (N_16620,N_16475,N_16574);
xor U16621 (N_16621,N_16531,N_16556);
or U16622 (N_16622,N_16562,N_16591);
xor U16623 (N_16623,N_16435,N_16473);
and U16624 (N_16624,N_16522,N_16482);
xor U16625 (N_16625,N_16516,N_16595);
nor U16626 (N_16626,N_16479,N_16599);
and U16627 (N_16627,N_16528,N_16544);
and U16628 (N_16628,N_16477,N_16587);
xnor U16629 (N_16629,N_16467,N_16437);
nand U16630 (N_16630,N_16461,N_16583);
xor U16631 (N_16631,N_16557,N_16576);
xor U16632 (N_16632,N_16553,N_16443);
xor U16633 (N_16633,N_16555,N_16417);
nor U16634 (N_16634,N_16448,N_16476);
xor U16635 (N_16635,N_16554,N_16414);
nand U16636 (N_16636,N_16505,N_16427);
nand U16637 (N_16637,N_16540,N_16512);
nor U16638 (N_16638,N_16547,N_16504);
xnor U16639 (N_16639,N_16455,N_16585);
or U16640 (N_16640,N_16432,N_16478);
nor U16641 (N_16641,N_16412,N_16523);
and U16642 (N_16642,N_16586,N_16539);
xor U16643 (N_16643,N_16496,N_16580);
or U16644 (N_16644,N_16501,N_16422);
or U16645 (N_16645,N_16508,N_16548);
nand U16646 (N_16646,N_16451,N_16551);
and U16647 (N_16647,N_16483,N_16563);
nand U16648 (N_16648,N_16573,N_16578);
nor U16649 (N_16649,N_16517,N_16532);
xor U16650 (N_16650,N_16525,N_16400);
and U16651 (N_16651,N_16570,N_16493);
nand U16652 (N_16652,N_16579,N_16530);
or U16653 (N_16653,N_16569,N_16515);
or U16654 (N_16654,N_16566,N_16441);
and U16655 (N_16655,N_16421,N_16460);
and U16656 (N_16656,N_16589,N_16444);
nor U16657 (N_16657,N_16485,N_16453);
nand U16658 (N_16658,N_16439,N_16537);
nor U16659 (N_16659,N_16538,N_16495);
xor U16660 (N_16660,N_16519,N_16564);
nand U16661 (N_16661,N_16484,N_16560);
and U16662 (N_16662,N_16456,N_16567);
nor U16663 (N_16663,N_16428,N_16565);
or U16664 (N_16664,N_16481,N_16542);
xor U16665 (N_16665,N_16597,N_16533);
xor U16666 (N_16666,N_16521,N_16429);
xor U16667 (N_16667,N_16568,N_16526);
and U16668 (N_16668,N_16438,N_16434);
nand U16669 (N_16669,N_16423,N_16598);
or U16670 (N_16670,N_16494,N_16543);
nand U16671 (N_16671,N_16449,N_16405);
or U16672 (N_16672,N_16559,N_16450);
and U16673 (N_16673,N_16430,N_16498);
or U16674 (N_16674,N_16454,N_16433);
or U16675 (N_16675,N_16416,N_16470);
nor U16676 (N_16676,N_16410,N_16536);
or U16677 (N_16677,N_16457,N_16584);
nor U16678 (N_16678,N_16409,N_16561);
and U16679 (N_16679,N_16507,N_16491);
and U16680 (N_16680,N_16588,N_16503);
nand U16681 (N_16681,N_16510,N_16558);
xnor U16682 (N_16682,N_16486,N_16459);
or U16683 (N_16683,N_16590,N_16571);
and U16684 (N_16684,N_16545,N_16549);
xnor U16685 (N_16685,N_16469,N_16468);
nand U16686 (N_16686,N_16572,N_16513);
xor U16687 (N_16687,N_16552,N_16440);
nand U16688 (N_16688,N_16465,N_16471);
xor U16689 (N_16689,N_16535,N_16480);
or U16690 (N_16690,N_16404,N_16431);
xor U16691 (N_16691,N_16406,N_16527);
and U16692 (N_16692,N_16472,N_16524);
xnor U16693 (N_16693,N_16402,N_16401);
and U16694 (N_16694,N_16415,N_16546);
or U16695 (N_16695,N_16582,N_16520);
or U16696 (N_16696,N_16511,N_16534);
xnor U16697 (N_16697,N_16452,N_16419);
or U16698 (N_16698,N_16424,N_16550);
or U16699 (N_16699,N_16593,N_16509);
or U16700 (N_16700,N_16486,N_16549);
and U16701 (N_16701,N_16520,N_16483);
nand U16702 (N_16702,N_16594,N_16580);
and U16703 (N_16703,N_16522,N_16404);
and U16704 (N_16704,N_16578,N_16465);
nor U16705 (N_16705,N_16510,N_16407);
nor U16706 (N_16706,N_16408,N_16477);
xnor U16707 (N_16707,N_16511,N_16566);
xor U16708 (N_16708,N_16509,N_16582);
nand U16709 (N_16709,N_16491,N_16480);
nor U16710 (N_16710,N_16452,N_16488);
nand U16711 (N_16711,N_16571,N_16422);
nor U16712 (N_16712,N_16559,N_16582);
xnor U16713 (N_16713,N_16457,N_16425);
and U16714 (N_16714,N_16560,N_16594);
nand U16715 (N_16715,N_16456,N_16594);
or U16716 (N_16716,N_16537,N_16409);
and U16717 (N_16717,N_16503,N_16461);
or U16718 (N_16718,N_16589,N_16548);
nor U16719 (N_16719,N_16409,N_16496);
or U16720 (N_16720,N_16476,N_16564);
or U16721 (N_16721,N_16520,N_16541);
or U16722 (N_16722,N_16509,N_16404);
xnor U16723 (N_16723,N_16514,N_16562);
xor U16724 (N_16724,N_16595,N_16464);
xor U16725 (N_16725,N_16412,N_16463);
and U16726 (N_16726,N_16546,N_16559);
xnor U16727 (N_16727,N_16425,N_16572);
xor U16728 (N_16728,N_16498,N_16411);
nand U16729 (N_16729,N_16535,N_16532);
and U16730 (N_16730,N_16445,N_16574);
or U16731 (N_16731,N_16489,N_16453);
nand U16732 (N_16732,N_16446,N_16596);
and U16733 (N_16733,N_16456,N_16595);
and U16734 (N_16734,N_16554,N_16476);
or U16735 (N_16735,N_16534,N_16559);
nand U16736 (N_16736,N_16590,N_16445);
and U16737 (N_16737,N_16595,N_16544);
nor U16738 (N_16738,N_16574,N_16532);
and U16739 (N_16739,N_16555,N_16502);
nor U16740 (N_16740,N_16580,N_16519);
nor U16741 (N_16741,N_16515,N_16594);
and U16742 (N_16742,N_16564,N_16491);
nor U16743 (N_16743,N_16568,N_16443);
nand U16744 (N_16744,N_16525,N_16511);
or U16745 (N_16745,N_16507,N_16594);
nor U16746 (N_16746,N_16570,N_16497);
or U16747 (N_16747,N_16453,N_16428);
nor U16748 (N_16748,N_16491,N_16439);
nand U16749 (N_16749,N_16400,N_16512);
and U16750 (N_16750,N_16552,N_16554);
or U16751 (N_16751,N_16546,N_16467);
and U16752 (N_16752,N_16537,N_16598);
nor U16753 (N_16753,N_16563,N_16556);
or U16754 (N_16754,N_16590,N_16470);
nand U16755 (N_16755,N_16491,N_16483);
xor U16756 (N_16756,N_16493,N_16461);
or U16757 (N_16757,N_16477,N_16492);
xor U16758 (N_16758,N_16426,N_16403);
nand U16759 (N_16759,N_16522,N_16515);
and U16760 (N_16760,N_16436,N_16508);
nor U16761 (N_16761,N_16481,N_16577);
nand U16762 (N_16762,N_16566,N_16543);
nor U16763 (N_16763,N_16492,N_16592);
and U16764 (N_16764,N_16497,N_16437);
xnor U16765 (N_16765,N_16599,N_16496);
nor U16766 (N_16766,N_16400,N_16446);
nand U16767 (N_16767,N_16475,N_16496);
and U16768 (N_16768,N_16447,N_16475);
nand U16769 (N_16769,N_16462,N_16402);
or U16770 (N_16770,N_16514,N_16572);
or U16771 (N_16771,N_16525,N_16439);
or U16772 (N_16772,N_16526,N_16577);
and U16773 (N_16773,N_16428,N_16458);
and U16774 (N_16774,N_16557,N_16410);
nand U16775 (N_16775,N_16417,N_16443);
xor U16776 (N_16776,N_16427,N_16422);
xor U16777 (N_16777,N_16489,N_16519);
or U16778 (N_16778,N_16514,N_16453);
nor U16779 (N_16779,N_16576,N_16505);
xor U16780 (N_16780,N_16599,N_16537);
nand U16781 (N_16781,N_16457,N_16504);
nand U16782 (N_16782,N_16439,N_16428);
nor U16783 (N_16783,N_16497,N_16599);
nor U16784 (N_16784,N_16553,N_16497);
nand U16785 (N_16785,N_16505,N_16543);
or U16786 (N_16786,N_16441,N_16531);
xnor U16787 (N_16787,N_16415,N_16423);
and U16788 (N_16788,N_16450,N_16539);
nor U16789 (N_16789,N_16523,N_16559);
nand U16790 (N_16790,N_16452,N_16537);
nor U16791 (N_16791,N_16478,N_16551);
or U16792 (N_16792,N_16543,N_16410);
xor U16793 (N_16793,N_16537,N_16549);
nor U16794 (N_16794,N_16539,N_16428);
nand U16795 (N_16795,N_16497,N_16577);
xnor U16796 (N_16796,N_16482,N_16497);
xor U16797 (N_16797,N_16577,N_16423);
nand U16798 (N_16798,N_16500,N_16586);
or U16799 (N_16799,N_16456,N_16506);
and U16800 (N_16800,N_16761,N_16720);
and U16801 (N_16801,N_16658,N_16775);
xor U16802 (N_16802,N_16625,N_16749);
and U16803 (N_16803,N_16696,N_16771);
and U16804 (N_16804,N_16676,N_16624);
nand U16805 (N_16805,N_16763,N_16770);
or U16806 (N_16806,N_16693,N_16772);
xnor U16807 (N_16807,N_16641,N_16683);
nor U16808 (N_16808,N_16726,N_16681);
and U16809 (N_16809,N_16774,N_16785);
xor U16810 (N_16810,N_16606,N_16661);
xor U16811 (N_16811,N_16751,N_16666);
and U16812 (N_16812,N_16668,N_16782);
xor U16813 (N_16813,N_16732,N_16787);
nand U16814 (N_16814,N_16753,N_16791);
xor U16815 (N_16815,N_16619,N_16691);
and U16816 (N_16816,N_16750,N_16703);
xor U16817 (N_16817,N_16780,N_16685);
xnor U16818 (N_16818,N_16605,N_16620);
or U16819 (N_16819,N_16739,N_16737);
and U16820 (N_16820,N_16645,N_16764);
xor U16821 (N_16821,N_16776,N_16613);
and U16822 (N_16822,N_16628,N_16712);
nor U16823 (N_16823,N_16632,N_16610);
and U16824 (N_16824,N_16724,N_16657);
and U16825 (N_16825,N_16649,N_16690);
or U16826 (N_16826,N_16654,N_16626);
nand U16827 (N_16827,N_16783,N_16653);
nand U16828 (N_16828,N_16634,N_16752);
nand U16829 (N_16829,N_16600,N_16794);
xor U16830 (N_16830,N_16709,N_16798);
or U16831 (N_16831,N_16621,N_16665);
or U16832 (N_16832,N_16730,N_16615);
nor U16833 (N_16833,N_16638,N_16677);
and U16834 (N_16834,N_16741,N_16722);
and U16835 (N_16835,N_16707,N_16652);
xor U16836 (N_16836,N_16686,N_16740);
and U16837 (N_16837,N_16612,N_16779);
or U16838 (N_16838,N_16608,N_16748);
nor U16839 (N_16839,N_16742,N_16604);
nor U16840 (N_16840,N_16717,N_16663);
nor U16841 (N_16841,N_16797,N_16680);
nand U16842 (N_16842,N_16647,N_16727);
nand U16843 (N_16843,N_16799,N_16725);
nor U16844 (N_16844,N_16640,N_16644);
nand U16845 (N_16845,N_16679,N_16745);
and U16846 (N_16846,N_16614,N_16602);
or U16847 (N_16847,N_16788,N_16646);
nand U16848 (N_16848,N_16762,N_16689);
nor U16849 (N_16849,N_16639,N_16656);
xnor U16850 (N_16850,N_16682,N_16684);
and U16851 (N_16851,N_16719,N_16757);
nor U16852 (N_16852,N_16714,N_16786);
nand U16853 (N_16853,N_16767,N_16735);
and U16854 (N_16854,N_16678,N_16754);
nand U16855 (N_16855,N_16773,N_16659);
xnor U16856 (N_16856,N_16708,N_16630);
xnor U16857 (N_16857,N_16700,N_16711);
nand U16858 (N_16858,N_16781,N_16702);
nand U16859 (N_16859,N_16631,N_16738);
and U16860 (N_16860,N_16705,N_16784);
nand U16861 (N_16861,N_16746,N_16721);
nor U16862 (N_16862,N_16716,N_16674);
and U16863 (N_16863,N_16651,N_16642);
and U16864 (N_16864,N_16672,N_16664);
nand U16865 (N_16865,N_16733,N_16671);
and U16866 (N_16866,N_16728,N_16694);
or U16867 (N_16867,N_16795,N_16636);
nor U16868 (N_16868,N_16760,N_16743);
or U16869 (N_16869,N_16777,N_16611);
xor U16870 (N_16870,N_16758,N_16796);
or U16871 (N_16871,N_16736,N_16697);
and U16872 (N_16872,N_16669,N_16650);
xnor U16873 (N_16873,N_16723,N_16789);
and U16874 (N_16874,N_16609,N_16765);
or U16875 (N_16875,N_16715,N_16759);
and U16876 (N_16876,N_16633,N_16643);
xor U16877 (N_16877,N_16718,N_16731);
nor U16878 (N_16878,N_16603,N_16687);
nor U16879 (N_16879,N_16637,N_16747);
or U16880 (N_16880,N_16635,N_16706);
and U16881 (N_16881,N_16692,N_16792);
and U16882 (N_16882,N_16618,N_16793);
and U16883 (N_16883,N_16698,N_16627);
xnor U16884 (N_16884,N_16673,N_16667);
or U16885 (N_16885,N_16701,N_16660);
or U16886 (N_16886,N_16734,N_16769);
and U16887 (N_16887,N_16713,N_16790);
xnor U16888 (N_16888,N_16675,N_16710);
and U16889 (N_16889,N_16622,N_16778);
or U16890 (N_16890,N_16756,N_16607);
and U16891 (N_16891,N_16768,N_16704);
and U16892 (N_16892,N_16616,N_16623);
and U16893 (N_16893,N_16670,N_16655);
or U16894 (N_16894,N_16688,N_16766);
nand U16895 (N_16895,N_16601,N_16755);
xnor U16896 (N_16896,N_16629,N_16617);
xor U16897 (N_16897,N_16662,N_16695);
nand U16898 (N_16898,N_16729,N_16648);
xnor U16899 (N_16899,N_16744,N_16699);
xor U16900 (N_16900,N_16659,N_16690);
or U16901 (N_16901,N_16749,N_16742);
nor U16902 (N_16902,N_16776,N_16681);
nor U16903 (N_16903,N_16620,N_16715);
and U16904 (N_16904,N_16704,N_16702);
and U16905 (N_16905,N_16641,N_16605);
and U16906 (N_16906,N_16787,N_16657);
xor U16907 (N_16907,N_16758,N_16707);
xor U16908 (N_16908,N_16691,N_16627);
or U16909 (N_16909,N_16610,N_16662);
and U16910 (N_16910,N_16750,N_16616);
nor U16911 (N_16911,N_16649,N_16603);
or U16912 (N_16912,N_16610,N_16646);
nand U16913 (N_16913,N_16689,N_16629);
xor U16914 (N_16914,N_16723,N_16745);
nor U16915 (N_16915,N_16700,N_16713);
nor U16916 (N_16916,N_16689,N_16769);
xnor U16917 (N_16917,N_16693,N_16630);
and U16918 (N_16918,N_16647,N_16620);
xnor U16919 (N_16919,N_16604,N_16667);
xnor U16920 (N_16920,N_16729,N_16774);
nor U16921 (N_16921,N_16786,N_16779);
nor U16922 (N_16922,N_16653,N_16775);
or U16923 (N_16923,N_16625,N_16775);
or U16924 (N_16924,N_16715,N_16682);
or U16925 (N_16925,N_16627,N_16768);
xor U16926 (N_16926,N_16679,N_16619);
or U16927 (N_16927,N_16643,N_16662);
or U16928 (N_16928,N_16759,N_16797);
nand U16929 (N_16929,N_16624,N_16694);
xor U16930 (N_16930,N_16702,N_16663);
xnor U16931 (N_16931,N_16682,N_16766);
or U16932 (N_16932,N_16754,N_16701);
nand U16933 (N_16933,N_16685,N_16784);
or U16934 (N_16934,N_16775,N_16713);
or U16935 (N_16935,N_16675,N_16619);
and U16936 (N_16936,N_16719,N_16773);
nor U16937 (N_16937,N_16764,N_16753);
nand U16938 (N_16938,N_16739,N_16701);
and U16939 (N_16939,N_16655,N_16607);
and U16940 (N_16940,N_16791,N_16797);
nor U16941 (N_16941,N_16782,N_16647);
or U16942 (N_16942,N_16602,N_16715);
or U16943 (N_16943,N_16725,N_16680);
nor U16944 (N_16944,N_16727,N_16620);
nand U16945 (N_16945,N_16771,N_16615);
xor U16946 (N_16946,N_16754,N_16698);
nor U16947 (N_16947,N_16607,N_16636);
and U16948 (N_16948,N_16698,N_16795);
and U16949 (N_16949,N_16777,N_16694);
xor U16950 (N_16950,N_16679,N_16617);
xor U16951 (N_16951,N_16650,N_16755);
or U16952 (N_16952,N_16620,N_16775);
nor U16953 (N_16953,N_16747,N_16726);
xnor U16954 (N_16954,N_16783,N_16719);
and U16955 (N_16955,N_16696,N_16772);
and U16956 (N_16956,N_16794,N_16714);
or U16957 (N_16957,N_16763,N_16640);
nor U16958 (N_16958,N_16752,N_16754);
nor U16959 (N_16959,N_16662,N_16730);
xnor U16960 (N_16960,N_16620,N_16709);
nand U16961 (N_16961,N_16778,N_16767);
xor U16962 (N_16962,N_16757,N_16722);
or U16963 (N_16963,N_16683,N_16787);
nand U16964 (N_16964,N_16715,N_16686);
or U16965 (N_16965,N_16677,N_16774);
nand U16966 (N_16966,N_16776,N_16616);
or U16967 (N_16967,N_16799,N_16603);
or U16968 (N_16968,N_16685,N_16766);
nor U16969 (N_16969,N_16609,N_16770);
or U16970 (N_16970,N_16602,N_16637);
or U16971 (N_16971,N_16632,N_16791);
nand U16972 (N_16972,N_16634,N_16662);
nand U16973 (N_16973,N_16657,N_16736);
xor U16974 (N_16974,N_16795,N_16664);
xor U16975 (N_16975,N_16786,N_16693);
or U16976 (N_16976,N_16625,N_16783);
nand U16977 (N_16977,N_16711,N_16684);
and U16978 (N_16978,N_16698,N_16606);
nand U16979 (N_16979,N_16705,N_16715);
xnor U16980 (N_16980,N_16689,N_16644);
or U16981 (N_16981,N_16732,N_16761);
or U16982 (N_16982,N_16715,N_16755);
nor U16983 (N_16983,N_16669,N_16796);
and U16984 (N_16984,N_16746,N_16700);
and U16985 (N_16985,N_16753,N_16719);
xor U16986 (N_16986,N_16660,N_16723);
nor U16987 (N_16987,N_16648,N_16761);
and U16988 (N_16988,N_16727,N_16668);
xor U16989 (N_16989,N_16647,N_16751);
nand U16990 (N_16990,N_16699,N_16647);
or U16991 (N_16991,N_16628,N_16608);
nand U16992 (N_16992,N_16716,N_16696);
xnor U16993 (N_16993,N_16666,N_16704);
nand U16994 (N_16994,N_16618,N_16792);
xnor U16995 (N_16995,N_16763,N_16721);
and U16996 (N_16996,N_16663,N_16634);
nand U16997 (N_16997,N_16688,N_16715);
nor U16998 (N_16998,N_16647,N_16638);
xnor U16999 (N_16999,N_16723,N_16684);
or U17000 (N_17000,N_16829,N_16935);
nor U17001 (N_17001,N_16959,N_16843);
nand U17002 (N_17002,N_16905,N_16813);
nor U17003 (N_17003,N_16926,N_16877);
or U17004 (N_17004,N_16956,N_16974);
xnor U17005 (N_17005,N_16976,N_16846);
xnor U17006 (N_17006,N_16801,N_16975);
and U17007 (N_17007,N_16887,N_16897);
and U17008 (N_17008,N_16849,N_16853);
nand U17009 (N_17009,N_16873,N_16891);
nand U17010 (N_17010,N_16800,N_16864);
and U17011 (N_17011,N_16820,N_16874);
nor U17012 (N_17012,N_16941,N_16899);
nand U17013 (N_17013,N_16821,N_16988);
xor U17014 (N_17014,N_16922,N_16992);
or U17015 (N_17015,N_16819,N_16951);
and U17016 (N_17016,N_16945,N_16978);
xnor U17017 (N_17017,N_16869,N_16982);
and U17018 (N_17018,N_16972,N_16940);
nor U17019 (N_17019,N_16844,N_16930);
nand U17020 (N_17020,N_16909,N_16936);
and U17021 (N_17021,N_16997,N_16817);
nor U17022 (N_17022,N_16833,N_16840);
or U17023 (N_17023,N_16987,N_16831);
or U17024 (N_17024,N_16994,N_16923);
xor U17025 (N_17025,N_16943,N_16867);
or U17026 (N_17026,N_16968,N_16848);
or U17027 (N_17027,N_16952,N_16900);
or U17028 (N_17028,N_16863,N_16962);
and U17029 (N_17029,N_16805,N_16880);
nand U17030 (N_17030,N_16857,N_16870);
and U17031 (N_17031,N_16850,N_16865);
and U17032 (N_17032,N_16989,N_16802);
nand U17033 (N_17033,N_16889,N_16804);
nand U17034 (N_17034,N_16983,N_16845);
nand U17035 (N_17035,N_16810,N_16855);
xor U17036 (N_17036,N_16854,N_16823);
xor U17037 (N_17037,N_16852,N_16862);
or U17038 (N_17038,N_16929,N_16914);
xnor U17039 (N_17039,N_16841,N_16816);
nor U17040 (N_17040,N_16828,N_16910);
xnor U17041 (N_17041,N_16830,N_16898);
nand U17042 (N_17042,N_16868,N_16904);
and U17043 (N_17043,N_16902,N_16949);
xnor U17044 (N_17044,N_16859,N_16928);
or U17045 (N_17045,N_16826,N_16906);
nand U17046 (N_17046,N_16903,N_16937);
xnor U17047 (N_17047,N_16835,N_16993);
xnor U17048 (N_17048,N_16818,N_16856);
or U17049 (N_17049,N_16806,N_16851);
xor U17050 (N_17050,N_16916,N_16955);
and U17051 (N_17051,N_16832,N_16809);
and U17052 (N_17052,N_16999,N_16967);
nor U17053 (N_17053,N_16847,N_16969);
or U17054 (N_17054,N_16939,N_16883);
nor U17055 (N_17055,N_16932,N_16827);
xnor U17056 (N_17056,N_16811,N_16964);
nand U17057 (N_17057,N_16950,N_16915);
nor U17058 (N_17058,N_16957,N_16980);
nor U17059 (N_17059,N_16970,N_16825);
and U17060 (N_17060,N_16858,N_16958);
and U17061 (N_17061,N_16838,N_16907);
nand U17062 (N_17062,N_16996,N_16812);
and U17063 (N_17063,N_16885,N_16878);
nor U17064 (N_17064,N_16881,N_16913);
nor U17065 (N_17065,N_16979,N_16875);
and U17066 (N_17066,N_16925,N_16938);
xnor U17067 (N_17067,N_16918,N_16837);
nor U17068 (N_17068,N_16893,N_16971);
xor U17069 (N_17069,N_16924,N_16942);
xor U17070 (N_17070,N_16872,N_16966);
xnor U17071 (N_17071,N_16961,N_16998);
nor U17072 (N_17072,N_16836,N_16927);
nor U17073 (N_17073,N_16944,N_16803);
nand U17074 (N_17074,N_16963,N_16912);
or U17075 (N_17075,N_16888,N_16931);
and U17076 (N_17076,N_16953,N_16990);
nand U17077 (N_17077,N_16895,N_16985);
xor U17078 (N_17078,N_16921,N_16896);
xor U17079 (N_17079,N_16884,N_16842);
nand U17080 (N_17080,N_16876,N_16808);
xor U17081 (N_17081,N_16919,N_16894);
xor U17082 (N_17082,N_16947,N_16984);
or U17083 (N_17083,N_16965,N_16908);
nand U17084 (N_17084,N_16807,N_16901);
or U17085 (N_17085,N_16892,N_16861);
or U17086 (N_17086,N_16886,N_16890);
xnor U17087 (N_17087,N_16954,N_16920);
xnor U17088 (N_17088,N_16814,N_16860);
and U17089 (N_17089,N_16995,N_16948);
nor U17090 (N_17090,N_16834,N_16934);
or U17091 (N_17091,N_16986,N_16977);
nand U17092 (N_17092,N_16882,N_16933);
and U17093 (N_17093,N_16981,N_16973);
nor U17094 (N_17094,N_16879,N_16946);
and U17095 (N_17095,N_16824,N_16871);
nand U17096 (N_17096,N_16866,N_16839);
and U17097 (N_17097,N_16991,N_16917);
nand U17098 (N_17098,N_16815,N_16822);
and U17099 (N_17099,N_16960,N_16911);
xnor U17100 (N_17100,N_16800,N_16977);
or U17101 (N_17101,N_16909,N_16833);
xor U17102 (N_17102,N_16910,N_16836);
and U17103 (N_17103,N_16896,N_16955);
and U17104 (N_17104,N_16914,N_16811);
or U17105 (N_17105,N_16886,N_16972);
xnor U17106 (N_17106,N_16877,N_16840);
nor U17107 (N_17107,N_16825,N_16811);
xnor U17108 (N_17108,N_16999,N_16809);
or U17109 (N_17109,N_16942,N_16895);
or U17110 (N_17110,N_16981,N_16857);
or U17111 (N_17111,N_16910,N_16889);
xor U17112 (N_17112,N_16843,N_16947);
xnor U17113 (N_17113,N_16870,N_16899);
or U17114 (N_17114,N_16876,N_16922);
nand U17115 (N_17115,N_16812,N_16972);
nand U17116 (N_17116,N_16859,N_16940);
or U17117 (N_17117,N_16907,N_16928);
xnor U17118 (N_17118,N_16991,N_16876);
nor U17119 (N_17119,N_16907,N_16861);
and U17120 (N_17120,N_16958,N_16974);
xor U17121 (N_17121,N_16833,N_16891);
or U17122 (N_17122,N_16948,N_16992);
and U17123 (N_17123,N_16939,N_16871);
nor U17124 (N_17124,N_16928,N_16917);
nand U17125 (N_17125,N_16901,N_16847);
or U17126 (N_17126,N_16911,N_16820);
nor U17127 (N_17127,N_16915,N_16940);
and U17128 (N_17128,N_16883,N_16943);
nand U17129 (N_17129,N_16977,N_16998);
and U17130 (N_17130,N_16843,N_16904);
or U17131 (N_17131,N_16904,N_16962);
and U17132 (N_17132,N_16816,N_16975);
nand U17133 (N_17133,N_16866,N_16958);
and U17134 (N_17134,N_16915,N_16800);
nor U17135 (N_17135,N_16813,N_16857);
or U17136 (N_17136,N_16960,N_16916);
and U17137 (N_17137,N_16837,N_16835);
xnor U17138 (N_17138,N_16998,N_16814);
and U17139 (N_17139,N_16865,N_16887);
xor U17140 (N_17140,N_16874,N_16829);
and U17141 (N_17141,N_16977,N_16855);
nand U17142 (N_17142,N_16940,N_16890);
xor U17143 (N_17143,N_16917,N_16801);
nor U17144 (N_17144,N_16906,N_16843);
nand U17145 (N_17145,N_16884,N_16883);
or U17146 (N_17146,N_16831,N_16940);
xnor U17147 (N_17147,N_16981,N_16804);
and U17148 (N_17148,N_16977,N_16927);
xor U17149 (N_17149,N_16826,N_16806);
and U17150 (N_17150,N_16873,N_16934);
xnor U17151 (N_17151,N_16836,N_16885);
nor U17152 (N_17152,N_16960,N_16861);
or U17153 (N_17153,N_16883,N_16811);
and U17154 (N_17154,N_16887,N_16804);
nor U17155 (N_17155,N_16931,N_16980);
xnor U17156 (N_17156,N_16833,N_16879);
or U17157 (N_17157,N_16965,N_16866);
xor U17158 (N_17158,N_16927,N_16979);
xnor U17159 (N_17159,N_16912,N_16863);
or U17160 (N_17160,N_16855,N_16996);
or U17161 (N_17161,N_16852,N_16966);
and U17162 (N_17162,N_16999,N_16987);
and U17163 (N_17163,N_16932,N_16918);
or U17164 (N_17164,N_16880,N_16977);
nor U17165 (N_17165,N_16922,N_16963);
nand U17166 (N_17166,N_16859,N_16853);
or U17167 (N_17167,N_16951,N_16942);
nand U17168 (N_17168,N_16833,N_16827);
nor U17169 (N_17169,N_16900,N_16977);
nand U17170 (N_17170,N_16840,N_16898);
or U17171 (N_17171,N_16844,N_16965);
nor U17172 (N_17172,N_16809,N_16967);
xnor U17173 (N_17173,N_16982,N_16906);
and U17174 (N_17174,N_16963,N_16972);
or U17175 (N_17175,N_16980,N_16821);
or U17176 (N_17176,N_16816,N_16874);
nor U17177 (N_17177,N_16801,N_16886);
nand U17178 (N_17178,N_16945,N_16845);
and U17179 (N_17179,N_16981,N_16955);
nor U17180 (N_17180,N_16948,N_16944);
nor U17181 (N_17181,N_16969,N_16988);
and U17182 (N_17182,N_16932,N_16997);
nand U17183 (N_17183,N_16929,N_16846);
nor U17184 (N_17184,N_16800,N_16905);
xnor U17185 (N_17185,N_16819,N_16948);
nand U17186 (N_17186,N_16810,N_16962);
and U17187 (N_17187,N_16939,N_16999);
nor U17188 (N_17188,N_16977,N_16848);
or U17189 (N_17189,N_16890,N_16860);
nand U17190 (N_17190,N_16960,N_16915);
nand U17191 (N_17191,N_16932,N_16802);
and U17192 (N_17192,N_16820,N_16997);
nor U17193 (N_17193,N_16816,N_16954);
xor U17194 (N_17194,N_16852,N_16819);
xnor U17195 (N_17195,N_16825,N_16959);
or U17196 (N_17196,N_16835,N_16900);
nand U17197 (N_17197,N_16809,N_16990);
nor U17198 (N_17198,N_16894,N_16966);
and U17199 (N_17199,N_16939,N_16840);
and U17200 (N_17200,N_17180,N_17183);
or U17201 (N_17201,N_17007,N_17132);
and U17202 (N_17202,N_17095,N_17071);
or U17203 (N_17203,N_17032,N_17008);
nand U17204 (N_17204,N_17164,N_17063);
nand U17205 (N_17205,N_17060,N_17006);
and U17206 (N_17206,N_17177,N_17146);
xor U17207 (N_17207,N_17159,N_17004);
nor U17208 (N_17208,N_17139,N_17131);
nor U17209 (N_17209,N_17038,N_17124);
nand U17210 (N_17210,N_17072,N_17054);
and U17211 (N_17211,N_17112,N_17126);
nand U17212 (N_17212,N_17020,N_17107);
and U17213 (N_17213,N_17036,N_17024);
nor U17214 (N_17214,N_17044,N_17156);
xor U17215 (N_17215,N_17172,N_17040);
xnor U17216 (N_17216,N_17068,N_17161);
nor U17217 (N_17217,N_17053,N_17197);
xor U17218 (N_17218,N_17014,N_17144);
xnor U17219 (N_17219,N_17153,N_17078);
nand U17220 (N_17220,N_17151,N_17075);
nand U17221 (N_17221,N_17138,N_17002);
and U17222 (N_17222,N_17011,N_17001);
xnor U17223 (N_17223,N_17101,N_17152);
or U17224 (N_17224,N_17021,N_17149);
or U17225 (N_17225,N_17106,N_17099);
xor U17226 (N_17226,N_17086,N_17052);
and U17227 (N_17227,N_17034,N_17087);
and U17228 (N_17228,N_17176,N_17108);
or U17229 (N_17229,N_17080,N_17104);
or U17230 (N_17230,N_17188,N_17182);
nand U17231 (N_17231,N_17169,N_17154);
xnor U17232 (N_17232,N_17173,N_17179);
nand U17233 (N_17233,N_17118,N_17127);
and U17234 (N_17234,N_17171,N_17163);
nor U17235 (N_17235,N_17140,N_17082);
nand U17236 (N_17236,N_17074,N_17039);
xnor U17237 (N_17237,N_17057,N_17048);
and U17238 (N_17238,N_17025,N_17056);
or U17239 (N_17239,N_17062,N_17174);
xnor U17240 (N_17240,N_17026,N_17136);
xor U17241 (N_17241,N_17045,N_17166);
nand U17242 (N_17242,N_17186,N_17097);
or U17243 (N_17243,N_17184,N_17162);
and U17244 (N_17244,N_17134,N_17130);
nor U17245 (N_17245,N_17129,N_17155);
nor U17246 (N_17246,N_17102,N_17160);
nand U17247 (N_17247,N_17100,N_17192);
nor U17248 (N_17248,N_17181,N_17051);
nand U17249 (N_17249,N_17079,N_17195);
nor U17250 (N_17250,N_17046,N_17147);
or U17251 (N_17251,N_17058,N_17033);
or U17252 (N_17252,N_17199,N_17041);
or U17253 (N_17253,N_17114,N_17190);
nor U17254 (N_17254,N_17096,N_17084);
nand U17255 (N_17255,N_17150,N_17091);
or U17256 (N_17256,N_17141,N_17116);
xnor U17257 (N_17257,N_17073,N_17123);
nand U17258 (N_17258,N_17185,N_17010);
nor U17259 (N_17259,N_17030,N_17117);
nand U17260 (N_17260,N_17092,N_17022);
and U17261 (N_17261,N_17088,N_17083);
and U17262 (N_17262,N_17000,N_17037);
xor U17263 (N_17263,N_17081,N_17187);
or U17264 (N_17264,N_17050,N_17055);
or U17265 (N_17265,N_17145,N_17076);
and U17266 (N_17266,N_17023,N_17120);
and U17267 (N_17267,N_17135,N_17125);
or U17268 (N_17268,N_17194,N_17017);
and U17269 (N_17269,N_17047,N_17193);
nand U17270 (N_17270,N_17009,N_17028);
nor U17271 (N_17271,N_17067,N_17110);
nand U17272 (N_17272,N_17111,N_17069);
xor U17273 (N_17273,N_17165,N_17113);
nand U17274 (N_17274,N_17158,N_17064);
xor U17275 (N_17275,N_17128,N_17198);
nor U17276 (N_17276,N_17065,N_17031);
xor U17277 (N_17277,N_17003,N_17119);
nor U17278 (N_17278,N_17018,N_17089);
or U17279 (N_17279,N_17178,N_17143);
or U17280 (N_17280,N_17066,N_17167);
nor U17281 (N_17281,N_17157,N_17191);
xnor U17282 (N_17282,N_17090,N_17061);
nor U17283 (N_17283,N_17059,N_17094);
nor U17284 (N_17284,N_17105,N_17133);
xor U17285 (N_17285,N_17168,N_17093);
nor U17286 (N_17286,N_17013,N_17085);
nand U17287 (N_17287,N_17098,N_17148);
nand U17288 (N_17288,N_17049,N_17035);
nand U17289 (N_17289,N_17122,N_17043);
xnor U17290 (N_17290,N_17109,N_17170);
and U17291 (N_17291,N_17016,N_17019);
xor U17292 (N_17292,N_17077,N_17137);
or U17293 (N_17293,N_17121,N_17029);
nand U17294 (N_17294,N_17189,N_17115);
xnor U17295 (N_17295,N_17175,N_17027);
nor U17296 (N_17296,N_17070,N_17196);
and U17297 (N_17297,N_17005,N_17042);
and U17298 (N_17298,N_17015,N_17142);
nand U17299 (N_17299,N_17103,N_17012);
or U17300 (N_17300,N_17000,N_17089);
nor U17301 (N_17301,N_17058,N_17095);
or U17302 (N_17302,N_17159,N_17077);
and U17303 (N_17303,N_17169,N_17003);
nor U17304 (N_17304,N_17056,N_17058);
nor U17305 (N_17305,N_17181,N_17088);
or U17306 (N_17306,N_17159,N_17089);
and U17307 (N_17307,N_17052,N_17002);
and U17308 (N_17308,N_17029,N_17073);
and U17309 (N_17309,N_17015,N_17039);
xor U17310 (N_17310,N_17182,N_17070);
nor U17311 (N_17311,N_17120,N_17067);
and U17312 (N_17312,N_17022,N_17091);
nor U17313 (N_17313,N_17148,N_17182);
or U17314 (N_17314,N_17081,N_17031);
xor U17315 (N_17315,N_17013,N_17040);
xnor U17316 (N_17316,N_17107,N_17036);
nor U17317 (N_17317,N_17130,N_17182);
nor U17318 (N_17318,N_17001,N_17144);
nor U17319 (N_17319,N_17162,N_17039);
xnor U17320 (N_17320,N_17053,N_17101);
xor U17321 (N_17321,N_17138,N_17160);
or U17322 (N_17322,N_17144,N_17127);
xnor U17323 (N_17323,N_17016,N_17022);
nor U17324 (N_17324,N_17145,N_17135);
and U17325 (N_17325,N_17140,N_17028);
nand U17326 (N_17326,N_17152,N_17140);
xnor U17327 (N_17327,N_17128,N_17035);
xnor U17328 (N_17328,N_17133,N_17004);
or U17329 (N_17329,N_17172,N_17024);
nand U17330 (N_17330,N_17060,N_17172);
or U17331 (N_17331,N_17159,N_17085);
nor U17332 (N_17332,N_17037,N_17175);
nand U17333 (N_17333,N_17022,N_17128);
xnor U17334 (N_17334,N_17132,N_17045);
nand U17335 (N_17335,N_17053,N_17177);
nor U17336 (N_17336,N_17068,N_17109);
and U17337 (N_17337,N_17033,N_17013);
nand U17338 (N_17338,N_17102,N_17023);
nand U17339 (N_17339,N_17194,N_17197);
nand U17340 (N_17340,N_17181,N_17055);
nor U17341 (N_17341,N_17107,N_17049);
xor U17342 (N_17342,N_17186,N_17083);
xor U17343 (N_17343,N_17115,N_17105);
and U17344 (N_17344,N_17131,N_17025);
xnor U17345 (N_17345,N_17192,N_17157);
xnor U17346 (N_17346,N_17133,N_17056);
or U17347 (N_17347,N_17032,N_17075);
nand U17348 (N_17348,N_17154,N_17115);
nand U17349 (N_17349,N_17037,N_17144);
xnor U17350 (N_17350,N_17182,N_17022);
and U17351 (N_17351,N_17091,N_17054);
nand U17352 (N_17352,N_17116,N_17081);
xor U17353 (N_17353,N_17132,N_17117);
nand U17354 (N_17354,N_17093,N_17159);
or U17355 (N_17355,N_17100,N_17175);
nor U17356 (N_17356,N_17037,N_17176);
and U17357 (N_17357,N_17021,N_17098);
nand U17358 (N_17358,N_17011,N_17103);
nand U17359 (N_17359,N_17078,N_17191);
nor U17360 (N_17360,N_17022,N_17082);
xor U17361 (N_17361,N_17039,N_17070);
or U17362 (N_17362,N_17082,N_17135);
xor U17363 (N_17363,N_17029,N_17005);
nand U17364 (N_17364,N_17199,N_17029);
nand U17365 (N_17365,N_17184,N_17136);
nand U17366 (N_17366,N_17083,N_17199);
and U17367 (N_17367,N_17177,N_17119);
xnor U17368 (N_17368,N_17151,N_17034);
nand U17369 (N_17369,N_17103,N_17132);
xnor U17370 (N_17370,N_17145,N_17189);
nand U17371 (N_17371,N_17100,N_17084);
xor U17372 (N_17372,N_17051,N_17038);
or U17373 (N_17373,N_17071,N_17006);
nor U17374 (N_17374,N_17127,N_17095);
nor U17375 (N_17375,N_17133,N_17029);
or U17376 (N_17376,N_17001,N_17052);
or U17377 (N_17377,N_17083,N_17171);
xor U17378 (N_17378,N_17074,N_17124);
or U17379 (N_17379,N_17194,N_17109);
nor U17380 (N_17380,N_17089,N_17166);
nor U17381 (N_17381,N_17180,N_17148);
or U17382 (N_17382,N_17197,N_17011);
nor U17383 (N_17383,N_17108,N_17146);
nand U17384 (N_17384,N_17067,N_17044);
or U17385 (N_17385,N_17135,N_17131);
nand U17386 (N_17386,N_17027,N_17160);
nor U17387 (N_17387,N_17121,N_17169);
and U17388 (N_17388,N_17137,N_17050);
xor U17389 (N_17389,N_17150,N_17089);
and U17390 (N_17390,N_17076,N_17049);
xnor U17391 (N_17391,N_17122,N_17066);
nand U17392 (N_17392,N_17177,N_17079);
nor U17393 (N_17393,N_17107,N_17158);
nand U17394 (N_17394,N_17015,N_17104);
xor U17395 (N_17395,N_17055,N_17138);
nand U17396 (N_17396,N_17003,N_17066);
or U17397 (N_17397,N_17090,N_17152);
nor U17398 (N_17398,N_17081,N_17120);
and U17399 (N_17399,N_17079,N_17186);
nor U17400 (N_17400,N_17278,N_17384);
nor U17401 (N_17401,N_17363,N_17242);
nand U17402 (N_17402,N_17220,N_17292);
nor U17403 (N_17403,N_17263,N_17324);
and U17404 (N_17404,N_17217,N_17393);
or U17405 (N_17405,N_17276,N_17306);
nor U17406 (N_17406,N_17274,N_17244);
and U17407 (N_17407,N_17265,N_17219);
nand U17408 (N_17408,N_17389,N_17345);
and U17409 (N_17409,N_17218,N_17241);
nor U17410 (N_17410,N_17396,N_17320);
and U17411 (N_17411,N_17310,N_17299);
or U17412 (N_17412,N_17348,N_17300);
or U17413 (N_17413,N_17236,N_17235);
or U17414 (N_17414,N_17256,N_17346);
or U17415 (N_17415,N_17397,N_17333);
and U17416 (N_17416,N_17215,N_17286);
or U17417 (N_17417,N_17337,N_17291);
nand U17418 (N_17418,N_17270,N_17223);
nand U17419 (N_17419,N_17246,N_17309);
or U17420 (N_17420,N_17232,N_17332);
xnor U17421 (N_17421,N_17289,N_17204);
nor U17422 (N_17422,N_17296,N_17216);
nand U17423 (N_17423,N_17343,N_17255);
xnor U17424 (N_17424,N_17351,N_17248);
and U17425 (N_17425,N_17392,N_17264);
or U17426 (N_17426,N_17288,N_17212);
xor U17427 (N_17427,N_17383,N_17322);
or U17428 (N_17428,N_17326,N_17331);
nand U17429 (N_17429,N_17319,N_17386);
xnor U17430 (N_17430,N_17398,N_17349);
nor U17431 (N_17431,N_17374,N_17370);
or U17432 (N_17432,N_17275,N_17339);
nand U17433 (N_17433,N_17239,N_17234);
or U17434 (N_17434,N_17379,N_17302);
or U17435 (N_17435,N_17366,N_17279);
xor U17436 (N_17436,N_17237,N_17316);
or U17437 (N_17437,N_17243,N_17259);
and U17438 (N_17438,N_17224,N_17329);
and U17439 (N_17439,N_17352,N_17254);
nand U17440 (N_17440,N_17390,N_17338);
and U17441 (N_17441,N_17202,N_17284);
nand U17442 (N_17442,N_17210,N_17294);
and U17443 (N_17443,N_17283,N_17353);
nand U17444 (N_17444,N_17388,N_17376);
nor U17445 (N_17445,N_17305,N_17277);
xnor U17446 (N_17446,N_17377,N_17262);
and U17447 (N_17447,N_17260,N_17361);
and U17448 (N_17448,N_17231,N_17214);
nand U17449 (N_17449,N_17267,N_17372);
nor U17450 (N_17450,N_17325,N_17280);
nand U17451 (N_17451,N_17367,N_17301);
nand U17452 (N_17452,N_17240,N_17252);
xor U17453 (N_17453,N_17378,N_17371);
or U17454 (N_17454,N_17211,N_17272);
nor U17455 (N_17455,N_17250,N_17330);
nand U17456 (N_17456,N_17365,N_17381);
or U17457 (N_17457,N_17382,N_17362);
xnor U17458 (N_17458,N_17399,N_17249);
nand U17459 (N_17459,N_17209,N_17247);
nand U17460 (N_17460,N_17253,N_17341);
or U17461 (N_17461,N_17328,N_17287);
and U17462 (N_17462,N_17315,N_17281);
xnor U17463 (N_17463,N_17313,N_17230);
nor U17464 (N_17464,N_17227,N_17293);
and U17465 (N_17465,N_17228,N_17380);
xnor U17466 (N_17466,N_17303,N_17285);
nor U17467 (N_17467,N_17312,N_17307);
nor U17468 (N_17468,N_17257,N_17373);
or U17469 (N_17469,N_17323,N_17206);
or U17470 (N_17470,N_17354,N_17203);
nor U17471 (N_17471,N_17314,N_17200);
xor U17472 (N_17472,N_17271,N_17269);
nor U17473 (N_17473,N_17391,N_17201);
and U17474 (N_17474,N_17311,N_17334);
and U17475 (N_17475,N_17213,N_17266);
or U17476 (N_17476,N_17394,N_17360);
or U17477 (N_17477,N_17359,N_17295);
nor U17478 (N_17478,N_17273,N_17385);
and U17479 (N_17479,N_17225,N_17335);
nor U17480 (N_17480,N_17375,N_17229);
or U17481 (N_17481,N_17395,N_17207);
nand U17482 (N_17482,N_17290,N_17233);
or U17483 (N_17483,N_17387,N_17327);
and U17484 (N_17484,N_17356,N_17342);
nor U17485 (N_17485,N_17304,N_17317);
nor U17486 (N_17486,N_17347,N_17282);
or U17487 (N_17487,N_17355,N_17245);
xnor U17488 (N_17488,N_17222,N_17358);
nor U17489 (N_17489,N_17308,N_17340);
xor U17490 (N_17490,N_17226,N_17364);
nor U17491 (N_17491,N_17238,N_17221);
and U17492 (N_17492,N_17350,N_17368);
nor U17493 (N_17493,N_17298,N_17251);
nand U17494 (N_17494,N_17208,N_17258);
nor U17495 (N_17495,N_17369,N_17336);
nor U17496 (N_17496,N_17357,N_17318);
and U17497 (N_17497,N_17321,N_17297);
nor U17498 (N_17498,N_17268,N_17205);
nor U17499 (N_17499,N_17261,N_17344);
and U17500 (N_17500,N_17384,N_17268);
or U17501 (N_17501,N_17325,N_17382);
nor U17502 (N_17502,N_17280,N_17321);
and U17503 (N_17503,N_17259,N_17296);
nand U17504 (N_17504,N_17293,N_17254);
nor U17505 (N_17505,N_17257,N_17321);
or U17506 (N_17506,N_17243,N_17256);
xor U17507 (N_17507,N_17324,N_17339);
or U17508 (N_17508,N_17328,N_17301);
or U17509 (N_17509,N_17205,N_17237);
and U17510 (N_17510,N_17340,N_17334);
or U17511 (N_17511,N_17360,N_17293);
and U17512 (N_17512,N_17391,N_17346);
nor U17513 (N_17513,N_17222,N_17300);
nand U17514 (N_17514,N_17318,N_17367);
xor U17515 (N_17515,N_17295,N_17393);
nand U17516 (N_17516,N_17268,N_17288);
or U17517 (N_17517,N_17291,N_17259);
xor U17518 (N_17518,N_17326,N_17213);
nand U17519 (N_17519,N_17301,N_17339);
and U17520 (N_17520,N_17333,N_17318);
xnor U17521 (N_17521,N_17250,N_17353);
nand U17522 (N_17522,N_17242,N_17201);
xor U17523 (N_17523,N_17302,N_17338);
xnor U17524 (N_17524,N_17378,N_17395);
or U17525 (N_17525,N_17361,N_17353);
or U17526 (N_17526,N_17217,N_17208);
nand U17527 (N_17527,N_17271,N_17388);
nand U17528 (N_17528,N_17371,N_17392);
xor U17529 (N_17529,N_17366,N_17295);
xor U17530 (N_17530,N_17239,N_17387);
nor U17531 (N_17531,N_17318,N_17337);
xor U17532 (N_17532,N_17249,N_17377);
nand U17533 (N_17533,N_17346,N_17315);
or U17534 (N_17534,N_17299,N_17306);
nand U17535 (N_17535,N_17261,N_17272);
and U17536 (N_17536,N_17325,N_17387);
xnor U17537 (N_17537,N_17259,N_17363);
and U17538 (N_17538,N_17294,N_17337);
nor U17539 (N_17539,N_17328,N_17396);
nand U17540 (N_17540,N_17305,N_17238);
nand U17541 (N_17541,N_17311,N_17351);
nand U17542 (N_17542,N_17235,N_17251);
or U17543 (N_17543,N_17327,N_17277);
nand U17544 (N_17544,N_17364,N_17215);
and U17545 (N_17545,N_17373,N_17200);
and U17546 (N_17546,N_17236,N_17265);
nor U17547 (N_17547,N_17309,N_17230);
nand U17548 (N_17548,N_17382,N_17230);
and U17549 (N_17549,N_17295,N_17379);
nor U17550 (N_17550,N_17370,N_17321);
xor U17551 (N_17551,N_17243,N_17369);
nand U17552 (N_17552,N_17357,N_17370);
nor U17553 (N_17553,N_17218,N_17286);
nand U17554 (N_17554,N_17295,N_17330);
nor U17555 (N_17555,N_17235,N_17333);
nor U17556 (N_17556,N_17287,N_17311);
nand U17557 (N_17557,N_17344,N_17228);
and U17558 (N_17558,N_17281,N_17222);
and U17559 (N_17559,N_17257,N_17212);
xnor U17560 (N_17560,N_17308,N_17208);
or U17561 (N_17561,N_17206,N_17326);
or U17562 (N_17562,N_17261,N_17303);
nor U17563 (N_17563,N_17356,N_17351);
or U17564 (N_17564,N_17334,N_17394);
xnor U17565 (N_17565,N_17243,N_17332);
or U17566 (N_17566,N_17284,N_17269);
and U17567 (N_17567,N_17324,N_17397);
or U17568 (N_17568,N_17304,N_17231);
and U17569 (N_17569,N_17326,N_17215);
and U17570 (N_17570,N_17207,N_17362);
or U17571 (N_17571,N_17258,N_17334);
nand U17572 (N_17572,N_17208,N_17300);
nor U17573 (N_17573,N_17216,N_17379);
xnor U17574 (N_17574,N_17256,N_17324);
and U17575 (N_17575,N_17258,N_17354);
nand U17576 (N_17576,N_17330,N_17322);
nand U17577 (N_17577,N_17246,N_17265);
nor U17578 (N_17578,N_17287,N_17300);
nor U17579 (N_17579,N_17338,N_17216);
nand U17580 (N_17580,N_17284,N_17369);
and U17581 (N_17581,N_17341,N_17209);
nor U17582 (N_17582,N_17244,N_17306);
xor U17583 (N_17583,N_17399,N_17292);
nor U17584 (N_17584,N_17337,N_17286);
nand U17585 (N_17585,N_17315,N_17218);
xor U17586 (N_17586,N_17296,N_17239);
and U17587 (N_17587,N_17371,N_17266);
nor U17588 (N_17588,N_17348,N_17340);
and U17589 (N_17589,N_17299,N_17289);
nand U17590 (N_17590,N_17337,N_17242);
nor U17591 (N_17591,N_17342,N_17205);
xnor U17592 (N_17592,N_17319,N_17266);
and U17593 (N_17593,N_17313,N_17287);
xor U17594 (N_17594,N_17215,N_17335);
nor U17595 (N_17595,N_17262,N_17204);
nor U17596 (N_17596,N_17318,N_17308);
nor U17597 (N_17597,N_17336,N_17340);
xnor U17598 (N_17598,N_17201,N_17377);
nor U17599 (N_17599,N_17366,N_17284);
nor U17600 (N_17600,N_17439,N_17592);
or U17601 (N_17601,N_17447,N_17403);
and U17602 (N_17602,N_17417,N_17567);
and U17603 (N_17603,N_17553,N_17500);
or U17604 (N_17604,N_17452,N_17412);
or U17605 (N_17605,N_17560,N_17472);
and U17606 (N_17606,N_17585,N_17531);
nand U17607 (N_17607,N_17438,N_17404);
and U17608 (N_17608,N_17426,N_17428);
or U17609 (N_17609,N_17579,N_17483);
nand U17610 (N_17610,N_17487,N_17590);
xnor U17611 (N_17611,N_17532,N_17528);
and U17612 (N_17612,N_17406,N_17411);
nor U17613 (N_17613,N_17571,N_17449);
nand U17614 (N_17614,N_17557,N_17416);
or U17615 (N_17615,N_17517,N_17423);
xnor U17616 (N_17616,N_17454,N_17538);
or U17617 (N_17617,N_17505,N_17573);
xor U17618 (N_17618,N_17476,N_17494);
nor U17619 (N_17619,N_17424,N_17451);
nor U17620 (N_17620,N_17565,N_17501);
and U17621 (N_17621,N_17499,N_17556);
or U17622 (N_17622,N_17530,N_17470);
nor U17623 (N_17623,N_17486,N_17473);
or U17624 (N_17624,N_17455,N_17540);
nor U17625 (N_17625,N_17575,N_17461);
nand U17626 (N_17626,N_17562,N_17492);
nand U17627 (N_17627,N_17525,N_17506);
and U17628 (N_17628,N_17593,N_17588);
and U17629 (N_17629,N_17463,N_17552);
xor U17630 (N_17630,N_17547,N_17489);
or U17631 (N_17631,N_17468,N_17535);
and U17632 (N_17632,N_17570,N_17563);
and U17633 (N_17633,N_17495,N_17533);
and U17634 (N_17634,N_17453,N_17576);
xnor U17635 (N_17635,N_17441,N_17566);
and U17636 (N_17636,N_17539,N_17515);
nor U17637 (N_17637,N_17536,N_17543);
xnor U17638 (N_17638,N_17549,N_17509);
nand U17639 (N_17639,N_17521,N_17418);
nor U17640 (N_17640,N_17457,N_17497);
nand U17641 (N_17641,N_17523,N_17529);
and U17642 (N_17642,N_17581,N_17580);
xnor U17643 (N_17643,N_17559,N_17482);
xnor U17644 (N_17644,N_17450,N_17534);
and U17645 (N_17645,N_17503,N_17513);
or U17646 (N_17646,N_17443,N_17548);
or U17647 (N_17647,N_17440,N_17436);
nor U17648 (N_17648,N_17421,N_17555);
xor U17649 (N_17649,N_17572,N_17496);
nand U17650 (N_17650,N_17493,N_17401);
or U17651 (N_17651,N_17419,N_17577);
nor U17652 (N_17652,N_17545,N_17480);
and U17653 (N_17653,N_17542,N_17471);
and U17654 (N_17654,N_17448,N_17591);
xor U17655 (N_17655,N_17481,N_17522);
nor U17656 (N_17656,N_17554,N_17456);
nand U17657 (N_17657,N_17596,N_17582);
nand U17658 (N_17658,N_17475,N_17507);
and U17659 (N_17659,N_17598,N_17442);
and U17660 (N_17660,N_17408,N_17595);
nor U17661 (N_17661,N_17409,N_17498);
and U17662 (N_17662,N_17519,N_17478);
and U17663 (N_17663,N_17437,N_17479);
or U17664 (N_17664,N_17516,N_17512);
and U17665 (N_17665,N_17541,N_17527);
xor U17666 (N_17666,N_17510,N_17474);
nor U17667 (N_17667,N_17465,N_17508);
and U17668 (N_17668,N_17429,N_17558);
xnor U17669 (N_17669,N_17462,N_17413);
and U17670 (N_17670,N_17407,N_17414);
or U17671 (N_17671,N_17584,N_17551);
nand U17672 (N_17672,N_17432,N_17459);
or U17673 (N_17673,N_17415,N_17402);
and U17674 (N_17674,N_17410,N_17488);
nand U17675 (N_17675,N_17544,N_17561);
nor U17676 (N_17676,N_17550,N_17433);
nand U17677 (N_17677,N_17422,N_17520);
or U17678 (N_17678,N_17524,N_17594);
nand U17679 (N_17679,N_17469,N_17460);
nand U17680 (N_17680,N_17537,N_17587);
nand U17681 (N_17681,N_17502,N_17484);
or U17682 (N_17682,N_17434,N_17504);
and U17683 (N_17683,N_17583,N_17564);
nand U17684 (N_17684,N_17477,N_17569);
nor U17685 (N_17685,N_17400,N_17597);
nand U17686 (N_17686,N_17430,N_17446);
and U17687 (N_17687,N_17485,N_17467);
or U17688 (N_17688,N_17405,N_17589);
and U17689 (N_17689,N_17464,N_17574);
nand U17690 (N_17690,N_17578,N_17546);
nand U17691 (N_17691,N_17511,N_17514);
and U17692 (N_17692,N_17420,N_17490);
and U17693 (N_17693,N_17599,N_17435);
nand U17694 (N_17694,N_17431,N_17445);
xnor U17695 (N_17695,N_17466,N_17458);
and U17696 (N_17696,N_17518,N_17568);
or U17697 (N_17697,N_17491,N_17586);
nor U17698 (N_17698,N_17444,N_17427);
or U17699 (N_17699,N_17526,N_17425);
xnor U17700 (N_17700,N_17467,N_17581);
nor U17701 (N_17701,N_17574,N_17448);
nor U17702 (N_17702,N_17414,N_17493);
nand U17703 (N_17703,N_17481,N_17504);
xor U17704 (N_17704,N_17546,N_17504);
and U17705 (N_17705,N_17423,N_17443);
or U17706 (N_17706,N_17571,N_17458);
nand U17707 (N_17707,N_17463,N_17422);
xnor U17708 (N_17708,N_17432,N_17485);
nor U17709 (N_17709,N_17468,N_17505);
xor U17710 (N_17710,N_17402,N_17428);
xor U17711 (N_17711,N_17414,N_17579);
nor U17712 (N_17712,N_17512,N_17479);
nor U17713 (N_17713,N_17455,N_17517);
or U17714 (N_17714,N_17495,N_17569);
nand U17715 (N_17715,N_17446,N_17541);
or U17716 (N_17716,N_17409,N_17524);
and U17717 (N_17717,N_17533,N_17456);
nand U17718 (N_17718,N_17453,N_17401);
or U17719 (N_17719,N_17483,N_17547);
or U17720 (N_17720,N_17409,N_17597);
or U17721 (N_17721,N_17483,N_17469);
or U17722 (N_17722,N_17448,N_17528);
or U17723 (N_17723,N_17525,N_17439);
nor U17724 (N_17724,N_17593,N_17404);
xnor U17725 (N_17725,N_17403,N_17413);
nor U17726 (N_17726,N_17415,N_17480);
xnor U17727 (N_17727,N_17589,N_17421);
nor U17728 (N_17728,N_17432,N_17564);
nand U17729 (N_17729,N_17576,N_17464);
xor U17730 (N_17730,N_17421,N_17467);
nor U17731 (N_17731,N_17468,N_17551);
and U17732 (N_17732,N_17570,N_17423);
nand U17733 (N_17733,N_17558,N_17479);
xnor U17734 (N_17734,N_17484,N_17538);
and U17735 (N_17735,N_17540,N_17469);
nand U17736 (N_17736,N_17553,N_17559);
xor U17737 (N_17737,N_17510,N_17534);
and U17738 (N_17738,N_17416,N_17560);
xnor U17739 (N_17739,N_17577,N_17482);
nor U17740 (N_17740,N_17484,N_17403);
xnor U17741 (N_17741,N_17475,N_17569);
and U17742 (N_17742,N_17414,N_17560);
nand U17743 (N_17743,N_17585,N_17569);
and U17744 (N_17744,N_17455,N_17491);
xor U17745 (N_17745,N_17526,N_17418);
or U17746 (N_17746,N_17535,N_17477);
or U17747 (N_17747,N_17525,N_17566);
and U17748 (N_17748,N_17553,N_17591);
xor U17749 (N_17749,N_17575,N_17563);
and U17750 (N_17750,N_17538,N_17520);
nor U17751 (N_17751,N_17553,N_17577);
or U17752 (N_17752,N_17582,N_17444);
or U17753 (N_17753,N_17444,N_17537);
xnor U17754 (N_17754,N_17507,N_17575);
and U17755 (N_17755,N_17491,N_17469);
or U17756 (N_17756,N_17543,N_17510);
nand U17757 (N_17757,N_17481,N_17425);
nor U17758 (N_17758,N_17438,N_17472);
xnor U17759 (N_17759,N_17474,N_17537);
nand U17760 (N_17760,N_17568,N_17537);
nor U17761 (N_17761,N_17417,N_17484);
and U17762 (N_17762,N_17457,N_17416);
and U17763 (N_17763,N_17587,N_17593);
or U17764 (N_17764,N_17579,N_17496);
nand U17765 (N_17765,N_17552,N_17528);
xnor U17766 (N_17766,N_17492,N_17461);
nand U17767 (N_17767,N_17436,N_17497);
nand U17768 (N_17768,N_17481,N_17440);
or U17769 (N_17769,N_17480,N_17506);
nor U17770 (N_17770,N_17437,N_17554);
xor U17771 (N_17771,N_17576,N_17403);
nor U17772 (N_17772,N_17455,N_17501);
or U17773 (N_17773,N_17478,N_17539);
nand U17774 (N_17774,N_17591,N_17477);
xor U17775 (N_17775,N_17578,N_17550);
nor U17776 (N_17776,N_17494,N_17560);
nor U17777 (N_17777,N_17470,N_17460);
and U17778 (N_17778,N_17472,N_17539);
nor U17779 (N_17779,N_17519,N_17568);
nor U17780 (N_17780,N_17506,N_17472);
xor U17781 (N_17781,N_17425,N_17444);
or U17782 (N_17782,N_17591,N_17409);
nand U17783 (N_17783,N_17599,N_17459);
nand U17784 (N_17784,N_17495,N_17458);
nand U17785 (N_17785,N_17582,N_17413);
or U17786 (N_17786,N_17488,N_17588);
xor U17787 (N_17787,N_17576,N_17429);
or U17788 (N_17788,N_17599,N_17439);
xor U17789 (N_17789,N_17564,N_17503);
nand U17790 (N_17790,N_17418,N_17499);
and U17791 (N_17791,N_17560,N_17421);
nand U17792 (N_17792,N_17534,N_17424);
xor U17793 (N_17793,N_17409,N_17462);
nand U17794 (N_17794,N_17419,N_17516);
nor U17795 (N_17795,N_17464,N_17561);
or U17796 (N_17796,N_17485,N_17422);
nand U17797 (N_17797,N_17522,N_17498);
nor U17798 (N_17798,N_17559,N_17577);
or U17799 (N_17799,N_17529,N_17558);
and U17800 (N_17800,N_17754,N_17648);
and U17801 (N_17801,N_17660,N_17688);
nand U17802 (N_17802,N_17691,N_17743);
nor U17803 (N_17803,N_17636,N_17772);
xor U17804 (N_17804,N_17661,N_17645);
xor U17805 (N_17805,N_17638,N_17750);
and U17806 (N_17806,N_17668,N_17655);
xor U17807 (N_17807,N_17604,N_17781);
and U17808 (N_17808,N_17644,N_17608);
nand U17809 (N_17809,N_17744,N_17747);
nand U17810 (N_17810,N_17762,N_17721);
and U17811 (N_17811,N_17756,N_17605);
or U17812 (N_17812,N_17687,N_17639);
xor U17813 (N_17813,N_17615,N_17631);
nand U17814 (N_17814,N_17777,N_17713);
nand U17815 (N_17815,N_17704,N_17731);
xnor U17816 (N_17816,N_17725,N_17717);
and U17817 (N_17817,N_17726,N_17702);
xnor U17818 (N_17818,N_17658,N_17663);
nor U17819 (N_17819,N_17724,N_17764);
or U17820 (N_17820,N_17718,N_17775);
or U17821 (N_17821,N_17755,N_17742);
nor U17822 (N_17822,N_17703,N_17679);
nand U17823 (N_17823,N_17716,N_17649);
or U17824 (N_17824,N_17746,N_17791);
nor U17825 (N_17825,N_17758,N_17728);
nand U17826 (N_17826,N_17727,N_17795);
xor U17827 (N_17827,N_17619,N_17776);
xnor U17828 (N_17828,N_17642,N_17705);
nor U17829 (N_17829,N_17602,N_17771);
and U17830 (N_17830,N_17618,N_17629);
or U17831 (N_17831,N_17712,N_17774);
and U17832 (N_17832,N_17799,N_17613);
and U17833 (N_17833,N_17637,N_17601);
or U17834 (N_17834,N_17616,N_17690);
nor U17835 (N_17835,N_17697,N_17693);
nor U17836 (N_17836,N_17650,N_17790);
nor U17837 (N_17837,N_17741,N_17740);
nor U17838 (N_17838,N_17798,N_17662);
or U17839 (N_17839,N_17677,N_17665);
or U17840 (N_17840,N_17696,N_17792);
nor U17841 (N_17841,N_17752,N_17607);
and U17842 (N_17842,N_17617,N_17794);
nand U17843 (N_17843,N_17733,N_17643);
or U17844 (N_17844,N_17735,N_17610);
xnor U17845 (N_17845,N_17773,N_17673);
nor U17846 (N_17846,N_17694,N_17614);
nand U17847 (N_17847,N_17698,N_17768);
nor U17848 (N_17848,N_17783,N_17670);
nand U17849 (N_17849,N_17748,N_17757);
nand U17850 (N_17850,N_17715,N_17761);
nor U17851 (N_17851,N_17708,N_17782);
nor U17852 (N_17852,N_17736,N_17763);
nand U17853 (N_17853,N_17779,N_17681);
nand U17854 (N_17854,N_17667,N_17714);
or U17855 (N_17855,N_17706,N_17634);
and U17856 (N_17856,N_17709,N_17793);
and U17857 (N_17857,N_17719,N_17766);
xnor U17858 (N_17858,N_17641,N_17720);
nor U17859 (N_17859,N_17753,N_17699);
nor U17860 (N_17860,N_17695,N_17711);
and U17861 (N_17861,N_17684,N_17729);
nor U17862 (N_17862,N_17620,N_17797);
and U17863 (N_17863,N_17669,N_17787);
nor U17864 (N_17864,N_17785,N_17786);
or U17865 (N_17865,N_17751,N_17737);
nand U17866 (N_17866,N_17640,N_17760);
and U17867 (N_17867,N_17635,N_17653);
nor U17868 (N_17868,N_17674,N_17680);
and U17869 (N_17869,N_17678,N_17624);
nand U17870 (N_17870,N_17646,N_17672);
or U17871 (N_17871,N_17651,N_17611);
nor U17872 (N_17872,N_17780,N_17657);
or U17873 (N_17873,N_17652,N_17630);
and U17874 (N_17874,N_17778,N_17749);
nand U17875 (N_17875,N_17659,N_17700);
nor U17876 (N_17876,N_17784,N_17633);
nand U17877 (N_17877,N_17730,N_17623);
nand U17878 (N_17878,N_17770,N_17622);
and U17879 (N_17879,N_17745,N_17671);
and U17880 (N_17880,N_17621,N_17732);
xnor U17881 (N_17881,N_17710,N_17769);
nor U17882 (N_17882,N_17682,N_17689);
and U17883 (N_17883,N_17796,N_17656);
xnor U17884 (N_17884,N_17767,N_17738);
and U17885 (N_17885,N_17612,N_17686);
nand U17886 (N_17886,N_17685,N_17632);
nor U17887 (N_17887,N_17600,N_17666);
or U17888 (N_17888,N_17739,N_17603);
xor U17889 (N_17889,N_17647,N_17606);
nor U17890 (N_17890,N_17626,N_17788);
and U17891 (N_17891,N_17627,N_17701);
nor U17892 (N_17892,N_17759,N_17654);
nand U17893 (N_17893,N_17683,N_17675);
or U17894 (N_17894,N_17734,N_17722);
nor U17895 (N_17895,N_17676,N_17609);
and U17896 (N_17896,N_17789,N_17664);
or U17897 (N_17897,N_17628,N_17723);
nand U17898 (N_17898,N_17625,N_17692);
xnor U17899 (N_17899,N_17765,N_17707);
nand U17900 (N_17900,N_17669,N_17700);
or U17901 (N_17901,N_17666,N_17684);
nor U17902 (N_17902,N_17744,N_17720);
xor U17903 (N_17903,N_17664,N_17699);
xnor U17904 (N_17904,N_17789,N_17767);
or U17905 (N_17905,N_17773,N_17614);
and U17906 (N_17906,N_17651,N_17764);
and U17907 (N_17907,N_17643,N_17674);
xor U17908 (N_17908,N_17642,N_17637);
or U17909 (N_17909,N_17671,N_17623);
and U17910 (N_17910,N_17605,N_17768);
nor U17911 (N_17911,N_17610,N_17696);
xnor U17912 (N_17912,N_17757,N_17769);
and U17913 (N_17913,N_17757,N_17655);
nand U17914 (N_17914,N_17634,N_17605);
nand U17915 (N_17915,N_17724,N_17775);
or U17916 (N_17916,N_17706,N_17713);
nor U17917 (N_17917,N_17740,N_17776);
xor U17918 (N_17918,N_17685,N_17690);
nor U17919 (N_17919,N_17642,N_17607);
xnor U17920 (N_17920,N_17796,N_17629);
nor U17921 (N_17921,N_17683,N_17654);
nand U17922 (N_17922,N_17769,N_17703);
or U17923 (N_17923,N_17722,N_17631);
nand U17924 (N_17924,N_17635,N_17651);
and U17925 (N_17925,N_17741,N_17780);
or U17926 (N_17926,N_17702,N_17660);
and U17927 (N_17927,N_17691,N_17629);
and U17928 (N_17928,N_17787,N_17619);
and U17929 (N_17929,N_17733,N_17619);
nand U17930 (N_17930,N_17600,N_17750);
nand U17931 (N_17931,N_17768,N_17712);
and U17932 (N_17932,N_17625,N_17731);
nor U17933 (N_17933,N_17785,N_17704);
and U17934 (N_17934,N_17642,N_17760);
nor U17935 (N_17935,N_17609,N_17638);
or U17936 (N_17936,N_17740,N_17646);
and U17937 (N_17937,N_17770,N_17625);
nor U17938 (N_17938,N_17639,N_17668);
or U17939 (N_17939,N_17624,N_17635);
xnor U17940 (N_17940,N_17616,N_17720);
nand U17941 (N_17941,N_17738,N_17723);
and U17942 (N_17942,N_17729,N_17644);
xnor U17943 (N_17943,N_17716,N_17609);
and U17944 (N_17944,N_17622,N_17793);
xor U17945 (N_17945,N_17615,N_17757);
xnor U17946 (N_17946,N_17618,N_17686);
or U17947 (N_17947,N_17758,N_17703);
nor U17948 (N_17948,N_17750,N_17776);
and U17949 (N_17949,N_17676,N_17667);
xnor U17950 (N_17950,N_17744,N_17798);
and U17951 (N_17951,N_17661,N_17721);
and U17952 (N_17952,N_17689,N_17782);
xnor U17953 (N_17953,N_17658,N_17694);
nand U17954 (N_17954,N_17607,N_17627);
xnor U17955 (N_17955,N_17673,N_17762);
nand U17956 (N_17956,N_17617,N_17629);
and U17957 (N_17957,N_17631,N_17666);
nor U17958 (N_17958,N_17799,N_17711);
nor U17959 (N_17959,N_17639,N_17788);
nand U17960 (N_17960,N_17641,N_17640);
nor U17961 (N_17961,N_17717,N_17713);
nand U17962 (N_17962,N_17618,N_17789);
nor U17963 (N_17963,N_17761,N_17646);
or U17964 (N_17964,N_17706,N_17755);
nor U17965 (N_17965,N_17635,N_17662);
nor U17966 (N_17966,N_17790,N_17642);
nand U17967 (N_17967,N_17768,N_17754);
nor U17968 (N_17968,N_17713,N_17676);
or U17969 (N_17969,N_17629,N_17763);
nor U17970 (N_17970,N_17676,N_17780);
nor U17971 (N_17971,N_17631,N_17743);
nor U17972 (N_17972,N_17643,N_17646);
and U17973 (N_17973,N_17609,N_17780);
or U17974 (N_17974,N_17791,N_17646);
or U17975 (N_17975,N_17741,N_17676);
or U17976 (N_17976,N_17640,N_17619);
nor U17977 (N_17977,N_17627,N_17615);
and U17978 (N_17978,N_17603,N_17769);
nor U17979 (N_17979,N_17777,N_17687);
and U17980 (N_17980,N_17644,N_17667);
nand U17981 (N_17981,N_17759,N_17762);
nand U17982 (N_17982,N_17645,N_17646);
nor U17983 (N_17983,N_17628,N_17633);
or U17984 (N_17984,N_17629,N_17786);
nor U17985 (N_17985,N_17712,N_17658);
xnor U17986 (N_17986,N_17744,N_17752);
xnor U17987 (N_17987,N_17681,N_17776);
nor U17988 (N_17988,N_17669,N_17751);
and U17989 (N_17989,N_17672,N_17649);
nand U17990 (N_17990,N_17759,N_17627);
nor U17991 (N_17991,N_17658,N_17665);
nand U17992 (N_17992,N_17721,N_17726);
nor U17993 (N_17993,N_17629,N_17762);
nand U17994 (N_17994,N_17753,N_17726);
or U17995 (N_17995,N_17740,N_17616);
xor U17996 (N_17996,N_17692,N_17682);
or U17997 (N_17997,N_17712,N_17626);
nand U17998 (N_17998,N_17679,N_17752);
or U17999 (N_17999,N_17716,N_17641);
nor U18000 (N_18000,N_17994,N_17806);
nand U18001 (N_18001,N_17982,N_17971);
and U18002 (N_18002,N_17943,N_17898);
or U18003 (N_18003,N_17878,N_17966);
nor U18004 (N_18004,N_17895,N_17809);
xor U18005 (N_18005,N_17944,N_17822);
or U18006 (N_18006,N_17891,N_17808);
and U18007 (N_18007,N_17914,N_17950);
and U18008 (N_18008,N_17913,N_17807);
nand U18009 (N_18009,N_17932,N_17974);
nand U18010 (N_18010,N_17849,N_17868);
nor U18011 (N_18011,N_17866,N_17845);
xnor U18012 (N_18012,N_17864,N_17985);
and U18013 (N_18013,N_17955,N_17946);
nor U18014 (N_18014,N_17826,N_17968);
nor U18015 (N_18015,N_17896,N_17999);
and U18016 (N_18016,N_17803,N_17885);
nand U18017 (N_18017,N_17902,N_17859);
nor U18018 (N_18018,N_17897,N_17860);
and U18019 (N_18019,N_17963,N_17996);
and U18020 (N_18020,N_17837,N_17906);
or U18021 (N_18021,N_17981,N_17827);
xnor U18022 (N_18022,N_17912,N_17976);
and U18023 (N_18023,N_17997,N_17931);
or U18024 (N_18024,N_17867,N_17852);
nor U18025 (N_18025,N_17909,N_17858);
nand U18026 (N_18026,N_17984,N_17908);
nand U18027 (N_18027,N_17915,N_17830);
or U18028 (N_18028,N_17821,N_17964);
nor U18029 (N_18029,N_17887,N_17818);
nor U18030 (N_18030,N_17930,N_17831);
or U18031 (N_18031,N_17870,N_17857);
or U18032 (N_18032,N_17947,N_17936);
or U18033 (N_18033,N_17881,N_17977);
xor U18034 (N_18034,N_17841,N_17889);
and U18035 (N_18035,N_17907,N_17899);
nor U18036 (N_18036,N_17834,N_17817);
and U18037 (N_18037,N_17998,N_17823);
nand U18038 (N_18038,N_17957,N_17846);
nor U18039 (N_18039,N_17884,N_17813);
nor U18040 (N_18040,N_17855,N_17901);
nor U18041 (N_18041,N_17992,N_17939);
xor U18042 (N_18042,N_17980,N_17938);
and U18043 (N_18043,N_17816,N_17917);
xor U18044 (N_18044,N_17862,N_17967);
nor U18045 (N_18045,N_17865,N_17850);
or U18046 (N_18046,N_17802,N_17820);
nor U18047 (N_18047,N_17851,N_17833);
xor U18048 (N_18048,N_17972,N_17805);
nor U18049 (N_18049,N_17928,N_17843);
xor U18050 (N_18050,N_17880,N_17923);
or U18051 (N_18051,N_17904,N_17874);
nor U18052 (N_18052,N_17910,N_17920);
or U18053 (N_18053,N_17995,N_17934);
or U18054 (N_18054,N_17954,N_17991);
nor U18055 (N_18055,N_17988,N_17801);
nor U18056 (N_18056,N_17819,N_17979);
xor U18057 (N_18057,N_17848,N_17970);
nor U18058 (N_18058,N_17960,N_17911);
and U18059 (N_18059,N_17804,N_17829);
xnor U18060 (N_18060,N_17814,N_17892);
nor U18061 (N_18061,N_17986,N_17875);
or U18062 (N_18062,N_17836,N_17956);
or U18063 (N_18063,N_17842,N_17888);
and U18064 (N_18064,N_17879,N_17925);
nor U18065 (N_18065,N_17937,N_17800);
or U18066 (N_18066,N_17962,N_17840);
nor U18067 (N_18067,N_17924,N_17872);
or U18068 (N_18068,N_17853,N_17941);
nand U18069 (N_18069,N_17838,N_17978);
xnor U18070 (N_18070,N_17900,N_17945);
or U18071 (N_18071,N_17824,N_17927);
or U18072 (N_18072,N_17973,N_17975);
xor U18073 (N_18073,N_17883,N_17863);
nor U18074 (N_18074,N_17969,N_17916);
and U18075 (N_18075,N_17832,N_17993);
or U18076 (N_18076,N_17933,N_17894);
nor U18077 (N_18077,N_17869,N_17953);
nand U18078 (N_18078,N_17812,N_17926);
xnor U18079 (N_18079,N_17958,N_17989);
xnor U18080 (N_18080,N_17810,N_17921);
and U18081 (N_18081,N_17922,N_17940);
and U18082 (N_18082,N_17987,N_17825);
or U18083 (N_18083,N_17949,N_17815);
and U18084 (N_18084,N_17811,N_17918);
or U18085 (N_18085,N_17847,N_17903);
and U18086 (N_18086,N_17871,N_17990);
nand U18087 (N_18087,N_17929,N_17873);
nand U18088 (N_18088,N_17952,N_17856);
xnor U18089 (N_18089,N_17844,N_17905);
and U18090 (N_18090,N_17886,N_17948);
and U18091 (N_18091,N_17959,N_17961);
xnor U18092 (N_18092,N_17890,N_17835);
nand U18093 (N_18093,N_17876,N_17877);
nand U18094 (N_18094,N_17965,N_17882);
xor U18095 (N_18095,N_17839,N_17854);
xnor U18096 (N_18096,N_17935,N_17942);
or U18097 (N_18097,N_17893,N_17861);
nor U18098 (N_18098,N_17951,N_17919);
xor U18099 (N_18099,N_17983,N_17828);
nor U18100 (N_18100,N_17922,N_17936);
and U18101 (N_18101,N_17883,N_17830);
nor U18102 (N_18102,N_17873,N_17822);
nand U18103 (N_18103,N_17816,N_17963);
and U18104 (N_18104,N_17897,N_17859);
xor U18105 (N_18105,N_17957,N_17833);
or U18106 (N_18106,N_17983,N_17870);
nand U18107 (N_18107,N_17974,N_17927);
or U18108 (N_18108,N_17905,N_17836);
xor U18109 (N_18109,N_17943,N_17949);
and U18110 (N_18110,N_17868,N_17949);
and U18111 (N_18111,N_17800,N_17960);
or U18112 (N_18112,N_17992,N_17852);
and U18113 (N_18113,N_17874,N_17823);
xor U18114 (N_18114,N_17803,N_17934);
or U18115 (N_18115,N_17930,N_17955);
nor U18116 (N_18116,N_17848,N_17852);
nand U18117 (N_18117,N_17973,N_17838);
or U18118 (N_18118,N_17894,N_17839);
or U18119 (N_18119,N_17836,N_17848);
xor U18120 (N_18120,N_17874,N_17973);
xnor U18121 (N_18121,N_17910,N_17880);
and U18122 (N_18122,N_17857,N_17835);
and U18123 (N_18123,N_17984,N_17870);
and U18124 (N_18124,N_17860,N_17804);
xnor U18125 (N_18125,N_17865,N_17843);
or U18126 (N_18126,N_17842,N_17966);
nand U18127 (N_18127,N_17994,N_17902);
or U18128 (N_18128,N_17867,N_17918);
xnor U18129 (N_18129,N_17870,N_17966);
and U18130 (N_18130,N_17937,N_17806);
or U18131 (N_18131,N_17907,N_17815);
nor U18132 (N_18132,N_17845,N_17962);
or U18133 (N_18133,N_17849,N_17991);
nand U18134 (N_18134,N_17971,N_17802);
xnor U18135 (N_18135,N_17835,N_17855);
and U18136 (N_18136,N_17858,N_17888);
or U18137 (N_18137,N_17923,N_17862);
or U18138 (N_18138,N_17935,N_17870);
nand U18139 (N_18139,N_17869,N_17977);
and U18140 (N_18140,N_17961,N_17821);
and U18141 (N_18141,N_17996,N_17926);
and U18142 (N_18142,N_17859,N_17943);
and U18143 (N_18143,N_17824,N_17905);
xor U18144 (N_18144,N_17915,N_17850);
or U18145 (N_18145,N_17885,N_17976);
or U18146 (N_18146,N_17868,N_17984);
or U18147 (N_18147,N_17990,N_17940);
nand U18148 (N_18148,N_17804,N_17800);
xnor U18149 (N_18149,N_17832,N_17912);
and U18150 (N_18150,N_17877,N_17855);
nand U18151 (N_18151,N_17809,N_17982);
or U18152 (N_18152,N_17953,N_17923);
and U18153 (N_18153,N_17895,N_17862);
nor U18154 (N_18154,N_17884,N_17933);
nand U18155 (N_18155,N_17846,N_17986);
or U18156 (N_18156,N_17964,N_17948);
nand U18157 (N_18157,N_17868,N_17960);
nor U18158 (N_18158,N_17835,N_17911);
or U18159 (N_18159,N_17811,N_17951);
and U18160 (N_18160,N_17806,N_17831);
and U18161 (N_18161,N_17926,N_17995);
and U18162 (N_18162,N_17991,N_17924);
nor U18163 (N_18163,N_17928,N_17894);
and U18164 (N_18164,N_17841,N_17931);
and U18165 (N_18165,N_17802,N_17891);
xor U18166 (N_18166,N_17889,N_17957);
or U18167 (N_18167,N_17941,N_17982);
nor U18168 (N_18168,N_17921,N_17900);
nor U18169 (N_18169,N_17860,N_17824);
nand U18170 (N_18170,N_17913,N_17884);
nand U18171 (N_18171,N_17938,N_17979);
xnor U18172 (N_18172,N_17879,N_17800);
and U18173 (N_18173,N_17832,N_17810);
or U18174 (N_18174,N_17950,N_17912);
nor U18175 (N_18175,N_17827,N_17930);
xor U18176 (N_18176,N_17931,N_17936);
or U18177 (N_18177,N_17832,N_17970);
xor U18178 (N_18178,N_17993,N_17979);
or U18179 (N_18179,N_17948,N_17884);
and U18180 (N_18180,N_17899,N_17840);
xnor U18181 (N_18181,N_17916,N_17885);
nand U18182 (N_18182,N_17960,N_17870);
and U18183 (N_18183,N_17880,N_17986);
xnor U18184 (N_18184,N_17992,N_17847);
nor U18185 (N_18185,N_17821,N_17861);
nor U18186 (N_18186,N_17912,N_17834);
nor U18187 (N_18187,N_17927,N_17960);
nor U18188 (N_18188,N_17863,N_17946);
xor U18189 (N_18189,N_17842,N_17911);
nor U18190 (N_18190,N_17843,N_17822);
and U18191 (N_18191,N_17801,N_17833);
or U18192 (N_18192,N_17854,N_17820);
and U18193 (N_18193,N_17970,N_17961);
or U18194 (N_18194,N_17884,N_17967);
or U18195 (N_18195,N_17985,N_17912);
or U18196 (N_18196,N_17807,N_17958);
or U18197 (N_18197,N_17981,N_17894);
nor U18198 (N_18198,N_17856,N_17893);
xor U18199 (N_18199,N_17885,N_17849);
or U18200 (N_18200,N_18062,N_18071);
or U18201 (N_18201,N_18065,N_18067);
or U18202 (N_18202,N_18184,N_18151);
nand U18203 (N_18203,N_18015,N_18188);
and U18204 (N_18204,N_18050,N_18162);
and U18205 (N_18205,N_18131,N_18135);
nor U18206 (N_18206,N_18112,N_18099);
xnor U18207 (N_18207,N_18199,N_18011);
nand U18208 (N_18208,N_18069,N_18105);
and U18209 (N_18209,N_18157,N_18150);
xor U18210 (N_18210,N_18006,N_18111);
and U18211 (N_18211,N_18023,N_18160);
xor U18212 (N_18212,N_18073,N_18085);
nor U18213 (N_18213,N_18002,N_18174);
xor U18214 (N_18214,N_18140,N_18136);
nand U18215 (N_18215,N_18117,N_18074);
and U18216 (N_18216,N_18154,N_18142);
nor U18217 (N_18217,N_18144,N_18179);
or U18218 (N_18218,N_18124,N_18147);
or U18219 (N_18219,N_18031,N_18021);
xnor U18220 (N_18220,N_18094,N_18058);
xor U18221 (N_18221,N_18103,N_18026);
nor U18222 (N_18222,N_18053,N_18101);
or U18223 (N_18223,N_18166,N_18076);
and U18224 (N_18224,N_18185,N_18004);
nor U18225 (N_18225,N_18192,N_18091);
or U18226 (N_18226,N_18196,N_18138);
and U18227 (N_18227,N_18033,N_18178);
or U18228 (N_18228,N_18007,N_18032);
xor U18229 (N_18229,N_18128,N_18010);
and U18230 (N_18230,N_18182,N_18037);
or U18231 (N_18231,N_18109,N_18152);
or U18232 (N_18232,N_18098,N_18102);
or U18233 (N_18233,N_18119,N_18156);
xor U18234 (N_18234,N_18164,N_18046);
nand U18235 (N_18235,N_18039,N_18122);
nand U18236 (N_18236,N_18044,N_18027);
nor U18237 (N_18237,N_18000,N_18030);
and U18238 (N_18238,N_18163,N_18080);
nor U18239 (N_18239,N_18127,N_18063);
xor U18240 (N_18240,N_18107,N_18090);
or U18241 (N_18241,N_18025,N_18155);
and U18242 (N_18242,N_18095,N_18014);
nor U18243 (N_18243,N_18040,N_18034);
and U18244 (N_18244,N_18132,N_18186);
and U18245 (N_18245,N_18001,N_18024);
xnor U18246 (N_18246,N_18134,N_18077);
and U18247 (N_18247,N_18173,N_18104);
or U18248 (N_18248,N_18054,N_18035);
nor U18249 (N_18249,N_18191,N_18116);
nor U18250 (N_18250,N_18167,N_18038);
xnor U18251 (N_18251,N_18159,N_18060);
nor U18252 (N_18252,N_18115,N_18056);
or U18253 (N_18253,N_18059,N_18018);
or U18254 (N_18254,N_18008,N_18092);
or U18255 (N_18255,N_18070,N_18113);
or U18256 (N_18256,N_18120,N_18052);
xnor U18257 (N_18257,N_18153,N_18019);
or U18258 (N_18258,N_18180,N_18049);
nand U18259 (N_18259,N_18064,N_18137);
xnor U18260 (N_18260,N_18183,N_18100);
nand U18261 (N_18261,N_18083,N_18013);
or U18262 (N_18262,N_18012,N_18082);
nand U18263 (N_18263,N_18187,N_18110);
nor U18264 (N_18264,N_18168,N_18133);
nand U18265 (N_18265,N_18081,N_18078);
or U18266 (N_18266,N_18123,N_18042);
nand U18267 (N_18267,N_18016,N_18176);
and U18268 (N_18268,N_18029,N_18005);
xnor U18269 (N_18269,N_18009,N_18197);
nand U18270 (N_18270,N_18125,N_18108);
or U18271 (N_18271,N_18055,N_18088);
nor U18272 (N_18272,N_18177,N_18047);
or U18273 (N_18273,N_18193,N_18017);
xnor U18274 (N_18274,N_18189,N_18145);
xor U18275 (N_18275,N_18048,N_18087);
nand U18276 (N_18276,N_18161,N_18003);
or U18277 (N_18277,N_18169,N_18118);
or U18278 (N_18278,N_18148,N_18096);
nand U18279 (N_18279,N_18171,N_18181);
nor U18280 (N_18280,N_18121,N_18190);
xnor U18281 (N_18281,N_18061,N_18089);
nor U18282 (N_18282,N_18129,N_18097);
and U18283 (N_18283,N_18172,N_18139);
and U18284 (N_18284,N_18075,N_18175);
xor U18285 (N_18285,N_18146,N_18149);
nand U18286 (N_18286,N_18114,N_18022);
or U18287 (N_18287,N_18195,N_18051);
nor U18288 (N_18288,N_18036,N_18041);
or U18289 (N_18289,N_18143,N_18086);
nor U18290 (N_18290,N_18028,N_18158);
nand U18291 (N_18291,N_18170,N_18045);
xor U18292 (N_18292,N_18066,N_18198);
or U18293 (N_18293,N_18057,N_18141);
nor U18294 (N_18294,N_18126,N_18130);
xor U18295 (N_18295,N_18165,N_18043);
or U18296 (N_18296,N_18072,N_18106);
xor U18297 (N_18297,N_18068,N_18084);
nand U18298 (N_18298,N_18093,N_18020);
nor U18299 (N_18299,N_18079,N_18194);
nor U18300 (N_18300,N_18193,N_18145);
xor U18301 (N_18301,N_18167,N_18156);
nor U18302 (N_18302,N_18129,N_18021);
and U18303 (N_18303,N_18095,N_18005);
nand U18304 (N_18304,N_18054,N_18130);
nand U18305 (N_18305,N_18183,N_18002);
and U18306 (N_18306,N_18098,N_18117);
xnor U18307 (N_18307,N_18052,N_18009);
nor U18308 (N_18308,N_18039,N_18022);
nand U18309 (N_18309,N_18165,N_18050);
nor U18310 (N_18310,N_18111,N_18182);
xor U18311 (N_18311,N_18092,N_18056);
nor U18312 (N_18312,N_18084,N_18122);
and U18313 (N_18313,N_18043,N_18126);
xnor U18314 (N_18314,N_18042,N_18131);
nand U18315 (N_18315,N_18175,N_18048);
nor U18316 (N_18316,N_18017,N_18181);
nand U18317 (N_18317,N_18021,N_18184);
nor U18318 (N_18318,N_18125,N_18135);
xor U18319 (N_18319,N_18014,N_18196);
and U18320 (N_18320,N_18056,N_18123);
xor U18321 (N_18321,N_18081,N_18040);
or U18322 (N_18322,N_18153,N_18109);
nand U18323 (N_18323,N_18078,N_18000);
or U18324 (N_18324,N_18150,N_18164);
and U18325 (N_18325,N_18102,N_18163);
and U18326 (N_18326,N_18074,N_18130);
nand U18327 (N_18327,N_18011,N_18156);
nand U18328 (N_18328,N_18074,N_18030);
nor U18329 (N_18329,N_18147,N_18039);
or U18330 (N_18330,N_18178,N_18058);
or U18331 (N_18331,N_18129,N_18001);
nand U18332 (N_18332,N_18101,N_18067);
xor U18333 (N_18333,N_18158,N_18027);
xor U18334 (N_18334,N_18152,N_18075);
nand U18335 (N_18335,N_18157,N_18002);
nor U18336 (N_18336,N_18094,N_18039);
nand U18337 (N_18337,N_18123,N_18126);
nor U18338 (N_18338,N_18019,N_18196);
xnor U18339 (N_18339,N_18130,N_18103);
and U18340 (N_18340,N_18180,N_18046);
nand U18341 (N_18341,N_18194,N_18091);
nand U18342 (N_18342,N_18003,N_18164);
and U18343 (N_18343,N_18084,N_18056);
nand U18344 (N_18344,N_18068,N_18117);
and U18345 (N_18345,N_18008,N_18065);
nor U18346 (N_18346,N_18176,N_18087);
nand U18347 (N_18347,N_18144,N_18096);
or U18348 (N_18348,N_18192,N_18180);
or U18349 (N_18349,N_18031,N_18177);
nand U18350 (N_18350,N_18158,N_18121);
xor U18351 (N_18351,N_18032,N_18117);
nor U18352 (N_18352,N_18059,N_18191);
nor U18353 (N_18353,N_18002,N_18069);
nand U18354 (N_18354,N_18180,N_18033);
nor U18355 (N_18355,N_18139,N_18132);
nand U18356 (N_18356,N_18000,N_18149);
or U18357 (N_18357,N_18133,N_18057);
xnor U18358 (N_18358,N_18118,N_18160);
or U18359 (N_18359,N_18182,N_18160);
nor U18360 (N_18360,N_18111,N_18132);
or U18361 (N_18361,N_18161,N_18091);
xnor U18362 (N_18362,N_18114,N_18077);
xnor U18363 (N_18363,N_18193,N_18065);
and U18364 (N_18364,N_18065,N_18121);
xnor U18365 (N_18365,N_18131,N_18181);
nor U18366 (N_18366,N_18114,N_18153);
or U18367 (N_18367,N_18081,N_18155);
or U18368 (N_18368,N_18112,N_18034);
and U18369 (N_18369,N_18171,N_18031);
and U18370 (N_18370,N_18145,N_18183);
xnor U18371 (N_18371,N_18124,N_18009);
and U18372 (N_18372,N_18151,N_18061);
nor U18373 (N_18373,N_18016,N_18154);
nor U18374 (N_18374,N_18008,N_18078);
and U18375 (N_18375,N_18103,N_18149);
xnor U18376 (N_18376,N_18152,N_18021);
xor U18377 (N_18377,N_18032,N_18043);
nand U18378 (N_18378,N_18024,N_18036);
xor U18379 (N_18379,N_18150,N_18116);
xor U18380 (N_18380,N_18091,N_18113);
nor U18381 (N_18381,N_18119,N_18151);
or U18382 (N_18382,N_18065,N_18096);
and U18383 (N_18383,N_18069,N_18055);
xor U18384 (N_18384,N_18162,N_18192);
nor U18385 (N_18385,N_18185,N_18046);
nand U18386 (N_18386,N_18181,N_18169);
and U18387 (N_18387,N_18013,N_18075);
and U18388 (N_18388,N_18033,N_18030);
xnor U18389 (N_18389,N_18175,N_18031);
nand U18390 (N_18390,N_18034,N_18121);
and U18391 (N_18391,N_18104,N_18105);
nor U18392 (N_18392,N_18107,N_18196);
xnor U18393 (N_18393,N_18071,N_18106);
nor U18394 (N_18394,N_18158,N_18172);
and U18395 (N_18395,N_18008,N_18032);
or U18396 (N_18396,N_18191,N_18192);
xor U18397 (N_18397,N_18058,N_18007);
nand U18398 (N_18398,N_18162,N_18079);
nor U18399 (N_18399,N_18167,N_18153);
and U18400 (N_18400,N_18209,N_18372);
xnor U18401 (N_18401,N_18306,N_18271);
xor U18402 (N_18402,N_18395,N_18244);
nand U18403 (N_18403,N_18374,N_18207);
or U18404 (N_18404,N_18295,N_18370);
nand U18405 (N_18405,N_18344,N_18227);
nand U18406 (N_18406,N_18336,N_18368);
nand U18407 (N_18407,N_18280,N_18330);
xnor U18408 (N_18408,N_18215,N_18226);
nand U18409 (N_18409,N_18219,N_18254);
xor U18410 (N_18410,N_18356,N_18290);
nor U18411 (N_18411,N_18279,N_18283);
and U18412 (N_18412,N_18246,N_18314);
nand U18413 (N_18413,N_18338,N_18259);
nor U18414 (N_18414,N_18318,N_18339);
nand U18415 (N_18415,N_18363,N_18304);
nor U18416 (N_18416,N_18264,N_18276);
xnor U18417 (N_18417,N_18360,N_18203);
nor U18418 (N_18418,N_18221,N_18245);
xnor U18419 (N_18419,N_18265,N_18296);
or U18420 (N_18420,N_18206,N_18371);
nand U18421 (N_18421,N_18294,N_18373);
nand U18422 (N_18422,N_18255,N_18321);
nor U18423 (N_18423,N_18311,N_18323);
nor U18424 (N_18424,N_18386,N_18319);
or U18425 (N_18425,N_18358,N_18303);
or U18426 (N_18426,N_18224,N_18268);
nand U18427 (N_18427,N_18378,N_18345);
nor U18428 (N_18428,N_18377,N_18313);
and U18429 (N_18429,N_18217,N_18269);
or U18430 (N_18430,N_18223,N_18347);
nor U18431 (N_18431,N_18293,N_18352);
and U18432 (N_18432,N_18383,N_18392);
nor U18433 (N_18433,N_18301,N_18208);
or U18434 (N_18434,N_18212,N_18234);
nand U18435 (N_18435,N_18394,N_18309);
and U18436 (N_18436,N_18284,N_18243);
nor U18437 (N_18437,N_18385,N_18367);
or U18438 (N_18438,N_18278,N_18326);
or U18439 (N_18439,N_18220,N_18287);
nand U18440 (N_18440,N_18289,N_18351);
and U18441 (N_18441,N_18256,N_18300);
or U18442 (N_18442,N_18298,N_18364);
xnor U18443 (N_18443,N_18241,N_18362);
xnor U18444 (N_18444,N_18308,N_18361);
or U18445 (N_18445,N_18285,N_18382);
xor U18446 (N_18446,N_18355,N_18248);
nor U18447 (N_18447,N_18222,N_18216);
or U18448 (N_18448,N_18291,N_18365);
nor U18449 (N_18449,N_18266,N_18320);
or U18450 (N_18450,N_18307,N_18399);
nand U18451 (N_18451,N_18312,N_18349);
nor U18452 (N_18452,N_18263,N_18315);
or U18453 (N_18453,N_18282,N_18341);
nor U18454 (N_18454,N_18353,N_18390);
or U18455 (N_18455,N_18233,N_18334);
xnor U18456 (N_18456,N_18381,N_18327);
nor U18457 (N_18457,N_18350,N_18379);
xor U18458 (N_18458,N_18340,N_18229);
or U18459 (N_18459,N_18387,N_18249);
or U18460 (N_18460,N_18218,N_18204);
or U18461 (N_18461,N_18333,N_18302);
or U18462 (N_18462,N_18237,N_18346);
nor U18463 (N_18463,N_18260,N_18275);
xnor U18464 (N_18464,N_18316,N_18236);
xor U18465 (N_18465,N_18230,N_18232);
nor U18466 (N_18466,N_18239,N_18348);
nor U18467 (N_18467,N_18359,N_18317);
and U18468 (N_18468,N_18329,N_18288);
nor U18469 (N_18469,N_18342,N_18228);
nand U18470 (N_18470,N_18238,N_18354);
or U18471 (N_18471,N_18398,N_18240);
or U18472 (N_18472,N_18213,N_18366);
and U18473 (N_18473,N_18397,N_18286);
nand U18474 (N_18474,N_18270,N_18299);
nand U18475 (N_18475,N_18262,N_18389);
and U18476 (N_18476,N_18273,N_18375);
nor U18477 (N_18477,N_18332,N_18200);
xor U18478 (N_18478,N_18235,N_18337);
or U18479 (N_18479,N_18214,N_18274);
or U18480 (N_18480,N_18211,N_18201);
and U18481 (N_18481,N_18225,N_18252);
nand U18482 (N_18482,N_18310,N_18210);
xnor U18483 (N_18483,N_18277,N_18396);
xor U18484 (N_18484,N_18376,N_18325);
xnor U18485 (N_18485,N_18202,N_18328);
and U18486 (N_18486,N_18205,N_18305);
xnor U18487 (N_18487,N_18242,N_18384);
and U18488 (N_18488,N_18391,N_18247);
and U18489 (N_18489,N_18331,N_18324);
and U18490 (N_18490,N_18281,N_18380);
nand U18491 (N_18491,N_18250,N_18335);
nor U18492 (N_18492,N_18251,N_18343);
nand U18493 (N_18493,N_18261,N_18297);
and U18494 (N_18494,N_18257,N_18267);
or U18495 (N_18495,N_18272,N_18231);
xor U18496 (N_18496,N_18292,N_18369);
nand U18497 (N_18497,N_18322,N_18357);
xor U18498 (N_18498,N_18393,N_18253);
or U18499 (N_18499,N_18388,N_18258);
nand U18500 (N_18500,N_18219,N_18386);
nor U18501 (N_18501,N_18267,N_18327);
and U18502 (N_18502,N_18390,N_18232);
xor U18503 (N_18503,N_18339,N_18210);
nand U18504 (N_18504,N_18342,N_18284);
xnor U18505 (N_18505,N_18212,N_18330);
nand U18506 (N_18506,N_18229,N_18236);
xor U18507 (N_18507,N_18256,N_18377);
nor U18508 (N_18508,N_18217,N_18254);
or U18509 (N_18509,N_18288,N_18317);
nor U18510 (N_18510,N_18365,N_18379);
xnor U18511 (N_18511,N_18271,N_18217);
xor U18512 (N_18512,N_18288,N_18369);
nand U18513 (N_18513,N_18327,N_18235);
or U18514 (N_18514,N_18280,N_18218);
nand U18515 (N_18515,N_18254,N_18323);
xnor U18516 (N_18516,N_18313,N_18349);
nor U18517 (N_18517,N_18300,N_18292);
or U18518 (N_18518,N_18399,N_18359);
xor U18519 (N_18519,N_18231,N_18383);
nor U18520 (N_18520,N_18219,N_18343);
or U18521 (N_18521,N_18384,N_18276);
or U18522 (N_18522,N_18342,N_18275);
nor U18523 (N_18523,N_18231,N_18336);
and U18524 (N_18524,N_18309,N_18303);
nand U18525 (N_18525,N_18336,N_18345);
xnor U18526 (N_18526,N_18288,N_18348);
xor U18527 (N_18527,N_18282,N_18360);
nor U18528 (N_18528,N_18292,N_18396);
and U18529 (N_18529,N_18319,N_18381);
or U18530 (N_18530,N_18234,N_18207);
or U18531 (N_18531,N_18366,N_18292);
nand U18532 (N_18532,N_18377,N_18383);
xor U18533 (N_18533,N_18301,N_18270);
and U18534 (N_18534,N_18238,N_18268);
or U18535 (N_18535,N_18253,N_18380);
nand U18536 (N_18536,N_18331,N_18274);
nor U18537 (N_18537,N_18368,N_18200);
xor U18538 (N_18538,N_18299,N_18311);
and U18539 (N_18539,N_18337,N_18269);
nor U18540 (N_18540,N_18216,N_18304);
nand U18541 (N_18541,N_18246,N_18278);
nor U18542 (N_18542,N_18285,N_18232);
nand U18543 (N_18543,N_18229,N_18212);
nand U18544 (N_18544,N_18371,N_18309);
xnor U18545 (N_18545,N_18210,N_18276);
and U18546 (N_18546,N_18362,N_18238);
or U18547 (N_18547,N_18365,N_18329);
or U18548 (N_18548,N_18295,N_18395);
nand U18549 (N_18549,N_18207,N_18224);
or U18550 (N_18550,N_18358,N_18274);
xor U18551 (N_18551,N_18318,N_18231);
xnor U18552 (N_18552,N_18254,N_18236);
nand U18553 (N_18553,N_18244,N_18317);
or U18554 (N_18554,N_18215,N_18256);
nor U18555 (N_18555,N_18329,N_18366);
nand U18556 (N_18556,N_18238,N_18343);
or U18557 (N_18557,N_18319,N_18257);
and U18558 (N_18558,N_18214,N_18202);
xor U18559 (N_18559,N_18245,N_18363);
nand U18560 (N_18560,N_18339,N_18377);
nor U18561 (N_18561,N_18364,N_18312);
and U18562 (N_18562,N_18248,N_18349);
nor U18563 (N_18563,N_18233,N_18270);
nand U18564 (N_18564,N_18344,N_18316);
or U18565 (N_18565,N_18243,N_18329);
and U18566 (N_18566,N_18215,N_18277);
nor U18567 (N_18567,N_18374,N_18211);
and U18568 (N_18568,N_18288,N_18229);
xor U18569 (N_18569,N_18386,N_18293);
nand U18570 (N_18570,N_18276,N_18220);
nand U18571 (N_18571,N_18298,N_18211);
and U18572 (N_18572,N_18259,N_18363);
nor U18573 (N_18573,N_18323,N_18349);
xor U18574 (N_18574,N_18379,N_18354);
xnor U18575 (N_18575,N_18371,N_18324);
nor U18576 (N_18576,N_18354,N_18340);
xor U18577 (N_18577,N_18207,N_18275);
xnor U18578 (N_18578,N_18279,N_18238);
nand U18579 (N_18579,N_18262,N_18359);
or U18580 (N_18580,N_18211,N_18398);
or U18581 (N_18581,N_18311,N_18398);
nand U18582 (N_18582,N_18336,N_18383);
nand U18583 (N_18583,N_18224,N_18338);
and U18584 (N_18584,N_18297,N_18314);
nand U18585 (N_18585,N_18272,N_18253);
nand U18586 (N_18586,N_18266,N_18292);
or U18587 (N_18587,N_18242,N_18393);
nor U18588 (N_18588,N_18229,N_18315);
and U18589 (N_18589,N_18353,N_18269);
nand U18590 (N_18590,N_18259,N_18356);
nand U18591 (N_18591,N_18211,N_18301);
or U18592 (N_18592,N_18305,N_18308);
nor U18593 (N_18593,N_18310,N_18390);
nor U18594 (N_18594,N_18276,N_18296);
xnor U18595 (N_18595,N_18397,N_18288);
or U18596 (N_18596,N_18231,N_18345);
nor U18597 (N_18597,N_18387,N_18261);
nand U18598 (N_18598,N_18372,N_18266);
or U18599 (N_18599,N_18328,N_18201);
xor U18600 (N_18600,N_18509,N_18589);
xnor U18601 (N_18601,N_18555,N_18505);
nand U18602 (N_18602,N_18540,N_18450);
xor U18603 (N_18603,N_18438,N_18514);
and U18604 (N_18604,N_18506,N_18489);
and U18605 (N_18605,N_18585,N_18541);
and U18606 (N_18606,N_18404,N_18479);
and U18607 (N_18607,N_18430,N_18442);
and U18608 (N_18608,N_18467,N_18542);
xor U18609 (N_18609,N_18434,N_18448);
nand U18610 (N_18610,N_18465,N_18451);
nor U18611 (N_18611,N_18432,N_18452);
and U18612 (N_18612,N_18461,N_18576);
or U18613 (N_18613,N_18449,N_18419);
xnor U18614 (N_18614,N_18410,N_18460);
and U18615 (N_18615,N_18496,N_18469);
nand U18616 (N_18616,N_18497,N_18420);
and U18617 (N_18617,N_18582,N_18474);
nor U18618 (N_18618,N_18554,N_18443);
xnor U18619 (N_18619,N_18488,N_18539);
xnor U18620 (N_18620,N_18584,N_18548);
or U18621 (N_18621,N_18466,N_18447);
nor U18622 (N_18622,N_18490,N_18411);
nor U18623 (N_18623,N_18527,N_18519);
and U18624 (N_18624,N_18416,N_18441);
or U18625 (N_18625,N_18413,N_18545);
or U18626 (N_18626,N_18536,N_18493);
xnor U18627 (N_18627,N_18522,N_18501);
xor U18628 (N_18628,N_18526,N_18583);
nand U18629 (N_18629,N_18546,N_18512);
nor U18630 (N_18630,N_18486,N_18464);
xor U18631 (N_18631,N_18424,N_18552);
nor U18632 (N_18632,N_18445,N_18440);
or U18633 (N_18633,N_18455,N_18510);
nor U18634 (N_18634,N_18433,N_18568);
xnor U18635 (N_18635,N_18518,N_18556);
nand U18636 (N_18636,N_18503,N_18476);
or U18637 (N_18637,N_18567,N_18577);
xor U18638 (N_18638,N_18558,N_18483);
xor U18639 (N_18639,N_18453,N_18504);
or U18640 (N_18640,N_18477,N_18561);
or U18641 (N_18641,N_18588,N_18400);
nor U18642 (N_18642,N_18468,N_18470);
or U18643 (N_18643,N_18457,N_18431);
or U18644 (N_18644,N_18418,N_18507);
or U18645 (N_18645,N_18562,N_18482);
nand U18646 (N_18646,N_18528,N_18500);
nor U18647 (N_18647,N_18480,N_18459);
or U18648 (N_18648,N_18596,N_18487);
nor U18649 (N_18649,N_18529,N_18569);
xnor U18650 (N_18650,N_18566,N_18523);
xor U18651 (N_18651,N_18516,N_18439);
nor U18652 (N_18652,N_18508,N_18579);
and U18653 (N_18653,N_18428,N_18560);
xnor U18654 (N_18654,N_18520,N_18590);
or U18655 (N_18655,N_18533,N_18429);
nor U18656 (N_18656,N_18551,N_18543);
and U18657 (N_18657,N_18498,N_18573);
nand U18658 (N_18658,N_18415,N_18598);
nand U18659 (N_18659,N_18553,N_18499);
or U18660 (N_18660,N_18532,N_18580);
nand U18661 (N_18661,N_18407,N_18481);
nand U18662 (N_18662,N_18425,N_18594);
nand U18663 (N_18663,N_18494,N_18402);
or U18664 (N_18664,N_18409,N_18591);
xor U18665 (N_18665,N_18456,N_18571);
and U18666 (N_18666,N_18538,N_18570);
xor U18667 (N_18667,N_18587,N_18524);
nand U18668 (N_18668,N_18586,N_18534);
nand U18669 (N_18669,N_18427,N_18471);
xnor U18670 (N_18670,N_18511,N_18436);
xnor U18671 (N_18671,N_18537,N_18559);
and U18672 (N_18672,N_18525,N_18421);
and U18673 (N_18673,N_18595,N_18574);
xor U18674 (N_18674,N_18547,N_18401);
nor U18675 (N_18675,N_18414,N_18597);
or U18676 (N_18676,N_18423,N_18550);
and U18677 (N_18677,N_18412,N_18593);
and U18678 (N_18678,N_18564,N_18515);
xor U18679 (N_18679,N_18405,N_18426);
nor U18680 (N_18680,N_18484,N_18473);
or U18681 (N_18681,N_18485,N_18435);
or U18682 (N_18682,N_18463,N_18535);
or U18683 (N_18683,N_18565,N_18417);
xor U18684 (N_18684,N_18563,N_18408);
nand U18685 (N_18685,N_18572,N_18444);
nor U18686 (N_18686,N_18422,N_18592);
xor U18687 (N_18687,N_18454,N_18521);
or U18688 (N_18688,N_18472,N_18544);
and U18689 (N_18689,N_18495,N_18530);
nor U18690 (N_18690,N_18531,N_18403);
nor U18691 (N_18691,N_18513,N_18549);
nor U18692 (N_18692,N_18437,N_18557);
nor U18693 (N_18693,N_18406,N_18475);
xor U18694 (N_18694,N_18462,N_18492);
nand U18695 (N_18695,N_18578,N_18517);
and U18696 (N_18696,N_18581,N_18458);
xnor U18697 (N_18697,N_18575,N_18599);
and U18698 (N_18698,N_18491,N_18502);
nand U18699 (N_18699,N_18478,N_18446);
nor U18700 (N_18700,N_18416,N_18482);
nor U18701 (N_18701,N_18421,N_18505);
nand U18702 (N_18702,N_18427,N_18495);
or U18703 (N_18703,N_18554,N_18453);
xor U18704 (N_18704,N_18563,N_18410);
and U18705 (N_18705,N_18414,N_18590);
and U18706 (N_18706,N_18542,N_18591);
nor U18707 (N_18707,N_18596,N_18543);
xor U18708 (N_18708,N_18431,N_18506);
and U18709 (N_18709,N_18597,N_18418);
or U18710 (N_18710,N_18590,N_18403);
nor U18711 (N_18711,N_18553,N_18580);
and U18712 (N_18712,N_18503,N_18485);
or U18713 (N_18713,N_18500,N_18552);
and U18714 (N_18714,N_18535,N_18523);
or U18715 (N_18715,N_18480,N_18467);
and U18716 (N_18716,N_18450,N_18433);
nand U18717 (N_18717,N_18535,N_18441);
and U18718 (N_18718,N_18482,N_18510);
xnor U18719 (N_18719,N_18518,N_18484);
xor U18720 (N_18720,N_18451,N_18428);
nand U18721 (N_18721,N_18556,N_18432);
or U18722 (N_18722,N_18484,N_18459);
nand U18723 (N_18723,N_18534,N_18448);
xnor U18724 (N_18724,N_18417,N_18533);
nor U18725 (N_18725,N_18485,N_18557);
xor U18726 (N_18726,N_18407,N_18455);
nand U18727 (N_18727,N_18476,N_18471);
or U18728 (N_18728,N_18536,N_18585);
and U18729 (N_18729,N_18493,N_18586);
xor U18730 (N_18730,N_18584,N_18406);
or U18731 (N_18731,N_18562,N_18539);
nor U18732 (N_18732,N_18456,N_18412);
or U18733 (N_18733,N_18513,N_18536);
nor U18734 (N_18734,N_18476,N_18417);
xor U18735 (N_18735,N_18498,N_18520);
nor U18736 (N_18736,N_18484,N_18426);
or U18737 (N_18737,N_18554,N_18414);
and U18738 (N_18738,N_18529,N_18594);
nand U18739 (N_18739,N_18524,N_18522);
or U18740 (N_18740,N_18518,N_18470);
and U18741 (N_18741,N_18523,N_18414);
nor U18742 (N_18742,N_18553,N_18471);
and U18743 (N_18743,N_18430,N_18494);
or U18744 (N_18744,N_18560,N_18597);
nand U18745 (N_18745,N_18570,N_18430);
nor U18746 (N_18746,N_18478,N_18518);
and U18747 (N_18747,N_18425,N_18556);
xnor U18748 (N_18748,N_18588,N_18405);
and U18749 (N_18749,N_18540,N_18410);
nand U18750 (N_18750,N_18511,N_18541);
nor U18751 (N_18751,N_18489,N_18420);
or U18752 (N_18752,N_18479,N_18564);
and U18753 (N_18753,N_18580,N_18547);
or U18754 (N_18754,N_18448,N_18592);
and U18755 (N_18755,N_18553,N_18548);
and U18756 (N_18756,N_18548,N_18592);
or U18757 (N_18757,N_18401,N_18415);
or U18758 (N_18758,N_18438,N_18401);
nor U18759 (N_18759,N_18522,N_18508);
nor U18760 (N_18760,N_18565,N_18508);
xnor U18761 (N_18761,N_18571,N_18522);
or U18762 (N_18762,N_18419,N_18578);
xnor U18763 (N_18763,N_18569,N_18468);
nor U18764 (N_18764,N_18488,N_18516);
xor U18765 (N_18765,N_18455,N_18569);
nor U18766 (N_18766,N_18485,N_18481);
nor U18767 (N_18767,N_18566,N_18494);
xor U18768 (N_18768,N_18579,N_18471);
nor U18769 (N_18769,N_18575,N_18452);
nor U18770 (N_18770,N_18593,N_18482);
nand U18771 (N_18771,N_18466,N_18423);
nand U18772 (N_18772,N_18488,N_18444);
xnor U18773 (N_18773,N_18583,N_18420);
or U18774 (N_18774,N_18558,N_18486);
or U18775 (N_18775,N_18575,N_18596);
nand U18776 (N_18776,N_18466,N_18565);
xor U18777 (N_18777,N_18403,N_18477);
and U18778 (N_18778,N_18409,N_18554);
nor U18779 (N_18779,N_18403,N_18573);
nor U18780 (N_18780,N_18454,N_18492);
or U18781 (N_18781,N_18478,N_18448);
xor U18782 (N_18782,N_18417,N_18410);
nor U18783 (N_18783,N_18457,N_18421);
nand U18784 (N_18784,N_18500,N_18481);
and U18785 (N_18785,N_18417,N_18517);
nor U18786 (N_18786,N_18583,N_18548);
nand U18787 (N_18787,N_18543,N_18589);
nor U18788 (N_18788,N_18510,N_18556);
nor U18789 (N_18789,N_18455,N_18467);
nand U18790 (N_18790,N_18418,N_18465);
and U18791 (N_18791,N_18424,N_18455);
nor U18792 (N_18792,N_18498,N_18471);
nor U18793 (N_18793,N_18450,N_18466);
and U18794 (N_18794,N_18565,N_18493);
xor U18795 (N_18795,N_18546,N_18578);
or U18796 (N_18796,N_18448,N_18485);
nor U18797 (N_18797,N_18419,N_18482);
and U18798 (N_18798,N_18436,N_18420);
nand U18799 (N_18799,N_18517,N_18525);
and U18800 (N_18800,N_18732,N_18666);
nor U18801 (N_18801,N_18664,N_18641);
nor U18802 (N_18802,N_18736,N_18765);
nand U18803 (N_18803,N_18779,N_18730);
or U18804 (N_18804,N_18615,N_18760);
and U18805 (N_18805,N_18603,N_18771);
and U18806 (N_18806,N_18650,N_18616);
and U18807 (N_18807,N_18738,N_18624);
or U18808 (N_18808,N_18633,N_18661);
xor U18809 (N_18809,N_18635,N_18672);
xnor U18810 (N_18810,N_18627,N_18705);
or U18811 (N_18811,N_18734,N_18658);
or U18812 (N_18812,N_18646,N_18639);
and U18813 (N_18813,N_18785,N_18747);
or U18814 (N_18814,N_18695,N_18679);
xnor U18815 (N_18815,N_18723,N_18655);
and U18816 (N_18816,N_18698,N_18746);
and U18817 (N_18817,N_18786,N_18636);
xnor U18818 (N_18818,N_18689,N_18733);
nor U18819 (N_18819,N_18690,N_18634);
or U18820 (N_18820,N_18601,N_18715);
nand U18821 (N_18821,N_18716,N_18762);
and U18822 (N_18822,N_18799,N_18703);
nand U18823 (N_18823,N_18725,N_18788);
or U18824 (N_18824,N_18757,N_18741);
nand U18825 (N_18825,N_18739,N_18653);
xor U18826 (N_18826,N_18776,N_18791);
nor U18827 (N_18827,N_18640,N_18677);
and U18828 (N_18828,N_18637,N_18623);
and U18829 (N_18829,N_18629,N_18630);
and U18830 (N_18830,N_18613,N_18610);
and U18831 (N_18831,N_18673,N_18674);
nor U18832 (N_18832,N_18711,N_18729);
nor U18833 (N_18833,N_18767,N_18774);
and U18834 (N_18834,N_18777,N_18797);
or U18835 (N_18835,N_18647,N_18675);
nor U18836 (N_18836,N_18709,N_18770);
nand U18837 (N_18837,N_18671,N_18707);
nand U18838 (N_18838,N_18609,N_18753);
xor U18839 (N_18839,N_18780,N_18687);
nand U18840 (N_18840,N_18652,N_18778);
nand U18841 (N_18841,N_18745,N_18743);
and U18842 (N_18842,N_18704,N_18602);
nor U18843 (N_18843,N_18787,N_18728);
and U18844 (N_18844,N_18682,N_18714);
and U18845 (N_18845,N_18758,N_18626);
or U18846 (N_18846,N_18644,N_18683);
or U18847 (N_18847,N_18618,N_18724);
xnor U18848 (N_18848,N_18648,N_18717);
and U18849 (N_18849,N_18660,N_18676);
nand U18850 (N_18850,N_18727,N_18670);
nor U18851 (N_18851,N_18726,N_18798);
nor U18852 (N_18852,N_18604,N_18693);
nand U18853 (N_18853,N_18751,N_18608);
nor U18854 (N_18854,N_18792,N_18692);
and U18855 (N_18855,N_18606,N_18617);
nand U18856 (N_18856,N_18600,N_18669);
or U18857 (N_18857,N_18775,N_18710);
xor U18858 (N_18858,N_18701,N_18699);
nand U18859 (N_18859,N_18796,N_18789);
or U18860 (N_18860,N_18622,N_18620);
nor U18861 (N_18861,N_18749,N_18750);
xor U18862 (N_18862,N_18756,N_18688);
xnor U18863 (N_18863,N_18663,N_18612);
or U18864 (N_18864,N_18643,N_18656);
xnor U18865 (N_18865,N_18783,N_18735);
xnor U18866 (N_18866,N_18681,N_18654);
and U18867 (N_18867,N_18713,N_18694);
and U18868 (N_18868,N_18773,N_18719);
xor U18869 (N_18869,N_18625,N_18607);
and U18870 (N_18870,N_18769,N_18632);
and U18871 (N_18871,N_18697,N_18642);
and U18872 (N_18872,N_18754,N_18761);
xor U18873 (N_18873,N_18645,N_18702);
nand U18874 (N_18874,N_18721,N_18794);
nor U18875 (N_18875,N_18621,N_18718);
or U18876 (N_18876,N_18722,N_18657);
nor U18877 (N_18877,N_18619,N_18781);
nand U18878 (N_18878,N_18611,N_18708);
or U18879 (N_18879,N_18691,N_18667);
nand U18880 (N_18880,N_18784,N_18744);
nor U18881 (N_18881,N_18720,N_18790);
nor U18882 (N_18882,N_18649,N_18678);
nand U18883 (N_18883,N_18684,N_18668);
nand U18884 (N_18884,N_18659,N_18759);
nand U18885 (N_18885,N_18696,N_18748);
and U18886 (N_18886,N_18638,N_18766);
and U18887 (N_18887,N_18742,N_18651);
and U18888 (N_18888,N_18755,N_18628);
xnor U18889 (N_18889,N_18614,N_18782);
or U18890 (N_18890,N_18752,N_18665);
nor U18891 (N_18891,N_18795,N_18700);
and U18892 (N_18892,N_18772,N_18605);
xor U18893 (N_18893,N_18737,N_18662);
xnor U18894 (N_18894,N_18706,N_18631);
xnor U18895 (N_18895,N_18685,N_18763);
or U18896 (N_18896,N_18793,N_18768);
nor U18897 (N_18897,N_18740,N_18764);
and U18898 (N_18898,N_18680,N_18686);
or U18899 (N_18899,N_18731,N_18712);
xor U18900 (N_18900,N_18732,N_18625);
and U18901 (N_18901,N_18741,N_18748);
and U18902 (N_18902,N_18718,N_18669);
nand U18903 (N_18903,N_18613,N_18617);
xnor U18904 (N_18904,N_18774,N_18608);
xnor U18905 (N_18905,N_18673,N_18633);
nand U18906 (N_18906,N_18787,N_18615);
nand U18907 (N_18907,N_18680,N_18702);
nor U18908 (N_18908,N_18613,N_18600);
nor U18909 (N_18909,N_18638,N_18771);
xnor U18910 (N_18910,N_18689,N_18692);
or U18911 (N_18911,N_18606,N_18667);
nor U18912 (N_18912,N_18796,N_18777);
or U18913 (N_18913,N_18756,N_18733);
nand U18914 (N_18914,N_18701,N_18709);
and U18915 (N_18915,N_18624,N_18633);
or U18916 (N_18916,N_18615,N_18703);
or U18917 (N_18917,N_18715,N_18629);
and U18918 (N_18918,N_18643,N_18685);
or U18919 (N_18919,N_18767,N_18761);
and U18920 (N_18920,N_18726,N_18614);
and U18921 (N_18921,N_18752,N_18631);
and U18922 (N_18922,N_18797,N_18720);
nor U18923 (N_18923,N_18743,N_18718);
nor U18924 (N_18924,N_18654,N_18735);
and U18925 (N_18925,N_18745,N_18789);
xor U18926 (N_18926,N_18678,N_18768);
xor U18927 (N_18927,N_18678,N_18763);
xor U18928 (N_18928,N_18782,N_18753);
and U18929 (N_18929,N_18629,N_18753);
and U18930 (N_18930,N_18794,N_18731);
nand U18931 (N_18931,N_18689,N_18735);
nor U18932 (N_18932,N_18694,N_18673);
and U18933 (N_18933,N_18679,N_18757);
and U18934 (N_18934,N_18734,N_18692);
or U18935 (N_18935,N_18698,N_18761);
nor U18936 (N_18936,N_18728,N_18722);
or U18937 (N_18937,N_18657,N_18743);
nor U18938 (N_18938,N_18601,N_18600);
or U18939 (N_18939,N_18790,N_18706);
xnor U18940 (N_18940,N_18748,N_18631);
or U18941 (N_18941,N_18750,N_18728);
nor U18942 (N_18942,N_18609,N_18754);
nor U18943 (N_18943,N_18703,N_18602);
nor U18944 (N_18944,N_18677,N_18759);
or U18945 (N_18945,N_18766,N_18704);
and U18946 (N_18946,N_18774,N_18710);
and U18947 (N_18947,N_18607,N_18740);
xor U18948 (N_18948,N_18703,N_18772);
nor U18949 (N_18949,N_18748,N_18726);
or U18950 (N_18950,N_18746,N_18755);
nand U18951 (N_18951,N_18728,N_18701);
nor U18952 (N_18952,N_18601,N_18621);
and U18953 (N_18953,N_18732,N_18655);
nor U18954 (N_18954,N_18646,N_18680);
nor U18955 (N_18955,N_18761,N_18612);
xnor U18956 (N_18956,N_18700,N_18735);
nor U18957 (N_18957,N_18793,N_18752);
xor U18958 (N_18958,N_18755,N_18687);
nor U18959 (N_18959,N_18661,N_18673);
and U18960 (N_18960,N_18721,N_18753);
and U18961 (N_18961,N_18747,N_18608);
nand U18962 (N_18962,N_18769,N_18662);
or U18963 (N_18963,N_18730,N_18737);
nand U18964 (N_18964,N_18673,N_18663);
nor U18965 (N_18965,N_18630,N_18645);
nor U18966 (N_18966,N_18790,N_18781);
or U18967 (N_18967,N_18705,N_18755);
and U18968 (N_18968,N_18627,N_18739);
xor U18969 (N_18969,N_18759,N_18668);
nand U18970 (N_18970,N_18691,N_18751);
nand U18971 (N_18971,N_18753,N_18794);
and U18972 (N_18972,N_18724,N_18670);
nor U18973 (N_18973,N_18747,N_18602);
nor U18974 (N_18974,N_18751,N_18727);
and U18975 (N_18975,N_18753,N_18732);
and U18976 (N_18976,N_18684,N_18766);
xor U18977 (N_18977,N_18678,N_18652);
and U18978 (N_18978,N_18755,N_18678);
and U18979 (N_18979,N_18726,N_18743);
nor U18980 (N_18980,N_18610,N_18661);
nor U18981 (N_18981,N_18707,N_18647);
or U18982 (N_18982,N_18648,N_18668);
xor U18983 (N_18983,N_18719,N_18756);
nor U18984 (N_18984,N_18743,N_18600);
nor U18985 (N_18985,N_18640,N_18617);
nor U18986 (N_18986,N_18680,N_18651);
and U18987 (N_18987,N_18624,N_18695);
nand U18988 (N_18988,N_18619,N_18735);
and U18989 (N_18989,N_18732,N_18742);
and U18990 (N_18990,N_18791,N_18782);
nand U18991 (N_18991,N_18656,N_18707);
or U18992 (N_18992,N_18675,N_18722);
nor U18993 (N_18993,N_18791,N_18729);
nand U18994 (N_18994,N_18714,N_18626);
xnor U18995 (N_18995,N_18796,N_18644);
or U18996 (N_18996,N_18739,N_18668);
and U18997 (N_18997,N_18636,N_18731);
xnor U18998 (N_18998,N_18735,N_18696);
and U18999 (N_18999,N_18668,N_18691);
and U19000 (N_19000,N_18893,N_18934);
xor U19001 (N_19001,N_18879,N_18800);
and U19002 (N_19002,N_18949,N_18845);
nand U19003 (N_19003,N_18810,N_18908);
or U19004 (N_19004,N_18927,N_18942);
or U19005 (N_19005,N_18946,N_18903);
nand U19006 (N_19006,N_18914,N_18923);
nor U19007 (N_19007,N_18981,N_18905);
or U19008 (N_19008,N_18843,N_18972);
and U19009 (N_19009,N_18881,N_18888);
xnor U19010 (N_19010,N_18804,N_18867);
or U19011 (N_19011,N_18830,N_18988);
nor U19012 (N_19012,N_18877,N_18863);
nor U19013 (N_19013,N_18841,N_18994);
nand U19014 (N_19014,N_18890,N_18937);
nand U19015 (N_19015,N_18938,N_18955);
and U19016 (N_19016,N_18947,N_18873);
xor U19017 (N_19017,N_18939,N_18971);
nor U19018 (N_19018,N_18999,N_18885);
and U19019 (N_19019,N_18948,N_18980);
or U19020 (N_19020,N_18808,N_18814);
xor U19021 (N_19021,N_18857,N_18901);
nand U19022 (N_19022,N_18909,N_18957);
xnor U19023 (N_19023,N_18855,N_18926);
xnor U19024 (N_19024,N_18907,N_18811);
or U19025 (N_19025,N_18839,N_18828);
xor U19026 (N_19026,N_18862,N_18819);
xnor U19027 (N_19027,N_18996,N_18992);
and U19028 (N_19028,N_18967,N_18887);
nand U19029 (N_19029,N_18978,N_18991);
xnor U19030 (N_19030,N_18861,N_18858);
nor U19031 (N_19031,N_18812,N_18977);
nand U19032 (N_19032,N_18979,N_18920);
and U19033 (N_19033,N_18974,N_18835);
nor U19034 (N_19034,N_18961,N_18860);
xnor U19035 (N_19035,N_18899,N_18874);
nand U19036 (N_19036,N_18973,N_18989);
or U19037 (N_19037,N_18976,N_18878);
or U19038 (N_19038,N_18809,N_18986);
nor U19039 (N_19039,N_18823,N_18849);
and U19040 (N_19040,N_18990,N_18884);
nand U19041 (N_19041,N_18966,N_18825);
nor U19042 (N_19042,N_18856,N_18802);
nor U19043 (N_19043,N_18951,N_18834);
nand U19044 (N_19044,N_18913,N_18997);
xnor U19045 (N_19045,N_18806,N_18910);
nor U19046 (N_19046,N_18963,N_18985);
or U19047 (N_19047,N_18940,N_18842);
nand U19048 (N_19048,N_18965,N_18818);
nand U19049 (N_19049,N_18850,N_18936);
nand U19050 (N_19050,N_18822,N_18803);
xnor U19051 (N_19051,N_18801,N_18870);
or U19052 (N_19052,N_18959,N_18925);
xnor U19053 (N_19053,N_18928,N_18917);
nand U19054 (N_19054,N_18962,N_18827);
and U19055 (N_19055,N_18950,N_18866);
xnor U19056 (N_19056,N_18851,N_18898);
or U19057 (N_19057,N_18871,N_18848);
nor U19058 (N_19058,N_18895,N_18875);
and U19059 (N_19059,N_18886,N_18852);
or U19060 (N_19060,N_18838,N_18969);
nor U19061 (N_19061,N_18805,N_18826);
or U19062 (N_19062,N_18869,N_18970);
xor U19063 (N_19063,N_18817,N_18956);
and U19064 (N_19064,N_18984,N_18902);
nand U19065 (N_19065,N_18935,N_18915);
nand U19066 (N_19066,N_18987,N_18889);
and U19067 (N_19067,N_18912,N_18924);
nand U19068 (N_19068,N_18931,N_18837);
xnor U19069 (N_19069,N_18900,N_18918);
or U19070 (N_19070,N_18883,N_18820);
or U19071 (N_19071,N_18832,N_18998);
xor U19072 (N_19072,N_18847,N_18836);
nor U19073 (N_19073,N_18916,N_18880);
or U19074 (N_19074,N_18824,N_18864);
xor U19075 (N_19075,N_18896,N_18941);
nand U19076 (N_19076,N_18943,N_18868);
nor U19077 (N_19077,N_18807,N_18945);
or U19078 (N_19078,N_18944,N_18829);
xor U19079 (N_19079,N_18954,N_18854);
xor U19080 (N_19080,N_18975,N_18831);
and U19081 (N_19081,N_18853,N_18897);
xnor U19082 (N_19082,N_18892,N_18815);
xnor U19083 (N_19083,N_18929,N_18993);
or U19084 (N_19084,N_18911,N_18816);
nor U19085 (N_19085,N_18932,N_18846);
and U19086 (N_19086,N_18952,N_18876);
nand U19087 (N_19087,N_18960,N_18840);
and U19088 (N_19088,N_18872,N_18882);
xor U19089 (N_19089,N_18906,N_18964);
nor U19090 (N_19090,N_18859,N_18922);
nor U19091 (N_19091,N_18968,N_18958);
or U19092 (N_19092,N_18813,N_18894);
xnor U19093 (N_19093,N_18953,N_18982);
nand U19094 (N_19094,N_18904,N_18995);
or U19095 (N_19095,N_18933,N_18891);
nand U19096 (N_19096,N_18919,N_18983);
and U19097 (N_19097,N_18930,N_18844);
and U19098 (N_19098,N_18865,N_18833);
or U19099 (N_19099,N_18821,N_18921);
and U19100 (N_19100,N_18989,N_18815);
or U19101 (N_19101,N_18994,N_18862);
or U19102 (N_19102,N_18980,N_18998);
nor U19103 (N_19103,N_18874,N_18814);
and U19104 (N_19104,N_18809,N_18834);
or U19105 (N_19105,N_18943,N_18927);
nor U19106 (N_19106,N_18869,N_18966);
nand U19107 (N_19107,N_18898,N_18929);
or U19108 (N_19108,N_18808,N_18810);
or U19109 (N_19109,N_18854,N_18919);
xor U19110 (N_19110,N_18808,N_18804);
nand U19111 (N_19111,N_18849,N_18879);
or U19112 (N_19112,N_18918,N_18932);
nand U19113 (N_19113,N_18820,N_18902);
xor U19114 (N_19114,N_18889,N_18984);
xor U19115 (N_19115,N_18847,N_18899);
nand U19116 (N_19116,N_18963,N_18979);
or U19117 (N_19117,N_18852,N_18936);
and U19118 (N_19118,N_18904,N_18953);
nand U19119 (N_19119,N_18910,N_18831);
nand U19120 (N_19120,N_18986,N_18869);
and U19121 (N_19121,N_18900,N_18892);
nand U19122 (N_19122,N_18834,N_18993);
nand U19123 (N_19123,N_18906,N_18822);
nand U19124 (N_19124,N_18971,N_18960);
and U19125 (N_19125,N_18992,N_18822);
xnor U19126 (N_19126,N_18815,N_18858);
or U19127 (N_19127,N_18832,N_18957);
and U19128 (N_19128,N_18815,N_18895);
or U19129 (N_19129,N_18800,N_18894);
nand U19130 (N_19130,N_18973,N_18879);
nor U19131 (N_19131,N_18829,N_18900);
nand U19132 (N_19132,N_18828,N_18822);
nand U19133 (N_19133,N_18821,N_18801);
and U19134 (N_19134,N_18905,N_18862);
and U19135 (N_19135,N_18852,N_18904);
nand U19136 (N_19136,N_18834,N_18805);
nor U19137 (N_19137,N_18999,N_18841);
or U19138 (N_19138,N_18918,N_18850);
nand U19139 (N_19139,N_18806,N_18954);
xor U19140 (N_19140,N_18967,N_18998);
nor U19141 (N_19141,N_18830,N_18828);
xnor U19142 (N_19142,N_18803,N_18827);
xor U19143 (N_19143,N_18952,N_18992);
nor U19144 (N_19144,N_18864,N_18877);
xnor U19145 (N_19145,N_18832,N_18879);
nor U19146 (N_19146,N_18826,N_18885);
and U19147 (N_19147,N_18923,N_18959);
and U19148 (N_19148,N_18803,N_18956);
nor U19149 (N_19149,N_18925,N_18969);
nand U19150 (N_19150,N_18973,N_18958);
or U19151 (N_19151,N_18938,N_18806);
or U19152 (N_19152,N_18967,N_18870);
or U19153 (N_19153,N_18839,N_18884);
xor U19154 (N_19154,N_18816,N_18967);
or U19155 (N_19155,N_18848,N_18820);
xnor U19156 (N_19156,N_18939,N_18829);
nand U19157 (N_19157,N_18801,N_18993);
or U19158 (N_19158,N_18868,N_18979);
nor U19159 (N_19159,N_18981,N_18878);
nand U19160 (N_19160,N_18917,N_18886);
xnor U19161 (N_19161,N_18812,N_18885);
or U19162 (N_19162,N_18954,N_18995);
xnor U19163 (N_19163,N_18905,N_18809);
xnor U19164 (N_19164,N_18949,N_18837);
nand U19165 (N_19165,N_18923,N_18946);
xor U19166 (N_19166,N_18913,N_18822);
nor U19167 (N_19167,N_18885,N_18853);
xnor U19168 (N_19168,N_18820,N_18874);
nand U19169 (N_19169,N_18809,N_18825);
nand U19170 (N_19170,N_18962,N_18808);
or U19171 (N_19171,N_18957,N_18894);
and U19172 (N_19172,N_18989,N_18951);
nor U19173 (N_19173,N_18938,N_18964);
nor U19174 (N_19174,N_18811,N_18942);
nand U19175 (N_19175,N_18967,N_18968);
nand U19176 (N_19176,N_18808,N_18811);
and U19177 (N_19177,N_18918,N_18853);
and U19178 (N_19178,N_18982,N_18977);
and U19179 (N_19179,N_18830,N_18935);
xnor U19180 (N_19180,N_18990,N_18891);
or U19181 (N_19181,N_18937,N_18978);
and U19182 (N_19182,N_18936,N_18809);
xnor U19183 (N_19183,N_18840,N_18920);
or U19184 (N_19184,N_18911,N_18910);
and U19185 (N_19185,N_18825,N_18907);
nor U19186 (N_19186,N_18888,N_18846);
or U19187 (N_19187,N_18836,N_18810);
nor U19188 (N_19188,N_18896,N_18916);
nand U19189 (N_19189,N_18871,N_18888);
and U19190 (N_19190,N_18833,N_18909);
or U19191 (N_19191,N_18898,N_18976);
or U19192 (N_19192,N_18970,N_18944);
nand U19193 (N_19193,N_18999,N_18828);
and U19194 (N_19194,N_18875,N_18874);
nand U19195 (N_19195,N_18838,N_18992);
xor U19196 (N_19196,N_18819,N_18821);
nor U19197 (N_19197,N_18974,N_18990);
or U19198 (N_19198,N_18812,N_18896);
and U19199 (N_19199,N_18947,N_18986);
nor U19200 (N_19200,N_19058,N_19122);
xor U19201 (N_19201,N_19120,N_19097);
nand U19202 (N_19202,N_19003,N_19115);
nor U19203 (N_19203,N_19061,N_19106);
or U19204 (N_19204,N_19002,N_19132);
nor U19205 (N_19205,N_19063,N_19175);
nor U19206 (N_19206,N_19173,N_19111);
or U19207 (N_19207,N_19001,N_19186);
nand U19208 (N_19208,N_19188,N_19109);
or U19209 (N_19209,N_19059,N_19052);
nor U19210 (N_19210,N_19022,N_19043);
and U19211 (N_19211,N_19136,N_19070);
xor U19212 (N_19212,N_19050,N_19131);
nor U19213 (N_19213,N_19068,N_19133);
nand U19214 (N_19214,N_19194,N_19086);
xnor U19215 (N_19215,N_19191,N_19161);
and U19216 (N_19216,N_19174,N_19121);
xnor U19217 (N_19217,N_19148,N_19139);
or U19218 (N_19218,N_19184,N_19105);
nand U19219 (N_19219,N_19123,N_19033);
xnor U19220 (N_19220,N_19113,N_19099);
xnor U19221 (N_19221,N_19066,N_19041);
nand U19222 (N_19222,N_19124,N_19076);
nand U19223 (N_19223,N_19015,N_19075);
and U19224 (N_19224,N_19026,N_19170);
xnor U19225 (N_19225,N_19071,N_19053);
nand U19226 (N_19226,N_19198,N_19134);
and U19227 (N_19227,N_19110,N_19129);
or U19228 (N_19228,N_19038,N_19012);
nand U19229 (N_19229,N_19119,N_19056);
nand U19230 (N_19230,N_19144,N_19095);
xor U19231 (N_19231,N_19032,N_19128);
and U19232 (N_19232,N_19190,N_19158);
and U19233 (N_19233,N_19079,N_19080);
nor U19234 (N_19234,N_19000,N_19102);
xor U19235 (N_19235,N_19196,N_19009);
nand U19236 (N_19236,N_19163,N_19195);
and U19237 (N_19237,N_19065,N_19023);
nor U19238 (N_19238,N_19157,N_19085);
xor U19239 (N_19239,N_19137,N_19168);
nand U19240 (N_19240,N_19048,N_19118);
nor U19241 (N_19241,N_19062,N_19096);
nor U19242 (N_19242,N_19146,N_19060);
and U19243 (N_19243,N_19069,N_19073);
nor U19244 (N_19244,N_19077,N_19153);
and U19245 (N_19245,N_19074,N_19107);
nand U19246 (N_19246,N_19125,N_19145);
nor U19247 (N_19247,N_19135,N_19092);
nand U19248 (N_19248,N_19116,N_19176);
nor U19249 (N_19249,N_19027,N_19094);
nand U19250 (N_19250,N_19151,N_19087);
and U19251 (N_19251,N_19159,N_19082);
xnor U19252 (N_19252,N_19057,N_19181);
nand U19253 (N_19253,N_19182,N_19114);
or U19254 (N_19254,N_19141,N_19169);
nand U19255 (N_19255,N_19108,N_19013);
nor U19256 (N_19256,N_19127,N_19126);
and U19257 (N_19257,N_19185,N_19081);
nor U19258 (N_19258,N_19164,N_19171);
or U19259 (N_19259,N_19093,N_19177);
nand U19260 (N_19260,N_19101,N_19083);
nand U19261 (N_19261,N_19089,N_19192);
nor U19262 (N_19262,N_19078,N_19047);
nand U19263 (N_19263,N_19034,N_19091);
xor U19264 (N_19264,N_19055,N_19160);
nand U19265 (N_19265,N_19004,N_19143);
nand U19266 (N_19266,N_19042,N_19183);
nand U19267 (N_19267,N_19199,N_19103);
and U19268 (N_19268,N_19098,N_19044);
or U19269 (N_19269,N_19014,N_19037);
nand U19270 (N_19270,N_19028,N_19049);
or U19271 (N_19271,N_19035,N_19142);
and U19272 (N_19272,N_19166,N_19152);
and U19273 (N_19273,N_19030,N_19007);
xnor U19274 (N_19274,N_19112,N_19138);
and U19275 (N_19275,N_19088,N_19172);
nand U19276 (N_19276,N_19008,N_19193);
nand U19277 (N_19277,N_19011,N_19067);
nor U19278 (N_19278,N_19039,N_19046);
or U19279 (N_19279,N_19064,N_19147);
xnor U19280 (N_19280,N_19025,N_19189);
nand U19281 (N_19281,N_19016,N_19024);
and U19282 (N_19282,N_19187,N_19051);
nor U19283 (N_19283,N_19162,N_19021);
xor U19284 (N_19284,N_19149,N_19020);
nand U19285 (N_19285,N_19005,N_19040);
xnor U19286 (N_19286,N_19018,N_19130);
or U19287 (N_19287,N_19090,N_19084);
and U19288 (N_19288,N_19117,N_19029);
nor U19289 (N_19289,N_19140,N_19165);
nand U19290 (N_19290,N_19036,N_19156);
or U19291 (N_19291,N_19045,N_19100);
xor U19292 (N_19292,N_19031,N_19019);
nor U19293 (N_19293,N_19017,N_19155);
or U19294 (N_19294,N_19179,N_19154);
xor U19295 (N_19295,N_19104,N_19072);
and U19296 (N_19296,N_19006,N_19054);
and U19297 (N_19297,N_19197,N_19010);
or U19298 (N_19298,N_19167,N_19180);
nand U19299 (N_19299,N_19150,N_19178);
xor U19300 (N_19300,N_19001,N_19044);
nand U19301 (N_19301,N_19039,N_19079);
and U19302 (N_19302,N_19092,N_19175);
nor U19303 (N_19303,N_19182,N_19014);
and U19304 (N_19304,N_19160,N_19006);
xnor U19305 (N_19305,N_19065,N_19110);
and U19306 (N_19306,N_19069,N_19148);
and U19307 (N_19307,N_19165,N_19023);
or U19308 (N_19308,N_19188,N_19106);
nor U19309 (N_19309,N_19066,N_19101);
xor U19310 (N_19310,N_19156,N_19014);
and U19311 (N_19311,N_19075,N_19056);
and U19312 (N_19312,N_19119,N_19179);
nor U19313 (N_19313,N_19135,N_19118);
xor U19314 (N_19314,N_19184,N_19144);
or U19315 (N_19315,N_19077,N_19156);
xnor U19316 (N_19316,N_19159,N_19144);
xor U19317 (N_19317,N_19007,N_19143);
or U19318 (N_19318,N_19120,N_19082);
xnor U19319 (N_19319,N_19050,N_19176);
or U19320 (N_19320,N_19036,N_19192);
xor U19321 (N_19321,N_19069,N_19165);
xnor U19322 (N_19322,N_19141,N_19108);
and U19323 (N_19323,N_19052,N_19035);
or U19324 (N_19324,N_19135,N_19071);
xnor U19325 (N_19325,N_19103,N_19116);
or U19326 (N_19326,N_19146,N_19008);
xor U19327 (N_19327,N_19177,N_19045);
and U19328 (N_19328,N_19066,N_19005);
and U19329 (N_19329,N_19060,N_19085);
nor U19330 (N_19330,N_19178,N_19032);
nor U19331 (N_19331,N_19149,N_19117);
nor U19332 (N_19332,N_19039,N_19092);
nor U19333 (N_19333,N_19079,N_19178);
nand U19334 (N_19334,N_19104,N_19051);
nor U19335 (N_19335,N_19077,N_19131);
nand U19336 (N_19336,N_19032,N_19124);
nand U19337 (N_19337,N_19168,N_19022);
xor U19338 (N_19338,N_19088,N_19071);
and U19339 (N_19339,N_19055,N_19179);
xnor U19340 (N_19340,N_19067,N_19109);
xor U19341 (N_19341,N_19070,N_19118);
and U19342 (N_19342,N_19141,N_19061);
and U19343 (N_19343,N_19018,N_19051);
or U19344 (N_19344,N_19092,N_19120);
nand U19345 (N_19345,N_19136,N_19177);
nand U19346 (N_19346,N_19045,N_19157);
and U19347 (N_19347,N_19115,N_19159);
or U19348 (N_19348,N_19073,N_19142);
nand U19349 (N_19349,N_19021,N_19135);
nand U19350 (N_19350,N_19157,N_19028);
nand U19351 (N_19351,N_19177,N_19151);
nand U19352 (N_19352,N_19044,N_19069);
nand U19353 (N_19353,N_19065,N_19133);
or U19354 (N_19354,N_19020,N_19159);
xnor U19355 (N_19355,N_19196,N_19044);
or U19356 (N_19356,N_19101,N_19142);
xor U19357 (N_19357,N_19008,N_19051);
and U19358 (N_19358,N_19169,N_19049);
and U19359 (N_19359,N_19134,N_19006);
and U19360 (N_19360,N_19163,N_19014);
xor U19361 (N_19361,N_19018,N_19152);
nand U19362 (N_19362,N_19081,N_19099);
nor U19363 (N_19363,N_19019,N_19074);
xor U19364 (N_19364,N_19171,N_19142);
and U19365 (N_19365,N_19053,N_19189);
or U19366 (N_19366,N_19070,N_19082);
and U19367 (N_19367,N_19085,N_19130);
nor U19368 (N_19368,N_19115,N_19027);
xnor U19369 (N_19369,N_19090,N_19076);
nor U19370 (N_19370,N_19170,N_19025);
or U19371 (N_19371,N_19173,N_19142);
and U19372 (N_19372,N_19083,N_19014);
nor U19373 (N_19373,N_19097,N_19178);
nor U19374 (N_19374,N_19116,N_19079);
xnor U19375 (N_19375,N_19167,N_19064);
nand U19376 (N_19376,N_19195,N_19102);
xor U19377 (N_19377,N_19118,N_19103);
nand U19378 (N_19378,N_19058,N_19011);
xor U19379 (N_19379,N_19043,N_19139);
xnor U19380 (N_19380,N_19065,N_19010);
and U19381 (N_19381,N_19014,N_19099);
nor U19382 (N_19382,N_19040,N_19017);
xnor U19383 (N_19383,N_19100,N_19115);
nor U19384 (N_19384,N_19089,N_19088);
nand U19385 (N_19385,N_19149,N_19034);
and U19386 (N_19386,N_19186,N_19061);
and U19387 (N_19387,N_19194,N_19118);
and U19388 (N_19388,N_19133,N_19110);
or U19389 (N_19389,N_19058,N_19038);
xnor U19390 (N_19390,N_19065,N_19052);
nand U19391 (N_19391,N_19177,N_19139);
and U19392 (N_19392,N_19000,N_19061);
or U19393 (N_19393,N_19134,N_19028);
or U19394 (N_19394,N_19169,N_19021);
or U19395 (N_19395,N_19072,N_19010);
xor U19396 (N_19396,N_19193,N_19122);
nor U19397 (N_19397,N_19039,N_19007);
xor U19398 (N_19398,N_19052,N_19088);
nand U19399 (N_19399,N_19020,N_19099);
or U19400 (N_19400,N_19364,N_19323);
nor U19401 (N_19401,N_19206,N_19201);
xor U19402 (N_19402,N_19244,N_19236);
and U19403 (N_19403,N_19370,N_19222);
nor U19404 (N_19404,N_19286,N_19371);
nor U19405 (N_19405,N_19301,N_19391);
and U19406 (N_19406,N_19397,N_19294);
nand U19407 (N_19407,N_19232,N_19270);
xor U19408 (N_19408,N_19247,N_19309);
xor U19409 (N_19409,N_19275,N_19289);
nand U19410 (N_19410,N_19252,N_19385);
and U19411 (N_19411,N_19314,N_19225);
nand U19412 (N_19412,N_19234,N_19271);
xnor U19413 (N_19413,N_19280,N_19228);
nor U19414 (N_19414,N_19342,N_19398);
nor U19415 (N_19415,N_19369,N_19384);
xnor U19416 (N_19416,N_19372,N_19213);
xnor U19417 (N_19417,N_19359,N_19214);
nor U19418 (N_19418,N_19219,N_19302);
and U19419 (N_19419,N_19267,N_19217);
xor U19420 (N_19420,N_19368,N_19324);
or U19421 (N_19421,N_19262,N_19346);
nor U19422 (N_19422,N_19373,N_19258);
or U19423 (N_19423,N_19380,N_19282);
nor U19424 (N_19424,N_19290,N_19387);
nand U19425 (N_19425,N_19283,N_19345);
and U19426 (N_19426,N_19202,N_19325);
and U19427 (N_19427,N_19330,N_19204);
and U19428 (N_19428,N_19281,N_19308);
or U19429 (N_19429,N_19362,N_19320);
nand U19430 (N_19430,N_19200,N_19240);
xor U19431 (N_19431,N_19340,N_19210);
nand U19432 (N_19432,N_19221,N_19353);
nand U19433 (N_19433,N_19277,N_19241);
nand U19434 (N_19434,N_19375,N_19295);
nand U19435 (N_19435,N_19343,N_19207);
and U19436 (N_19436,N_19312,N_19205);
or U19437 (N_19437,N_19296,N_19284);
and U19438 (N_19438,N_19350,N_19399);
or U19439 (N_19439,N_19378,N_19336);
xor U19440 (N_19440,N_19263,N_19249);
xor U19441 (N_19441,N_19274,N_19321);
xor U19442 (N_19442,N_19276,N_19233);
and U19443 (N_19443,N_19208,N_19382);
or U19444 (N_19444,N_19355,N_19331);
and U19445 (N_19445,N_19297,N_19245);
and U19446 (N_19446,N_19278,N_19348);
and U19447 (N_19447,N_19253,N_19315);
nand U19448 (N_19448,N_19361,N_19363);
nor U19449 (N_19449,N_19332,N_19344);
and U19450 (N_19450,N_19335,N_19386);
or U19451 (N_19451,N_19215,N_19334);
nor U19452 (N_19452,N_19352,N_19231);
nor U19453 (N_19453,N_19269,N_19360);
and U19454 (N_19454,N_19227,N_19341);
nand U19455 (N_19455,N_19251,N_19326);
nor U19456 (N_19456,N_19310,N_19381);
or U19457 (N_19457,N_19260,N_19266);
or U19458 (N_19458,N_19379,N_19242);
and U19459 (N_19459,N_19351,N_19256);
xnor U19460 (N_19460,N_19216,N_19328);
nor U19461 (N_19461,N_19235,N_19261);
xor U19462 (N_19462,N_19272,N_19291);
or U19463 (N_19463,N_19238,N_19354);
and U19464 (N_19464,N_19376,N_19383);
nand U19465 (N_19465,N_19358,N_19300);
or U19466 (N_19466,N_19307,N_19224);
or U19467 (N_19467,N_19313,N_19306);
nor U19468 (N_19468,N_19367,N_19349);
or U19469 (N_19469,N_19357,N_19327);
or U19470 (N_19470,N_19264,N_19229);
and U19471 (N_19471,N_19318,N_19255);
or U19472 (N_19472,N_19239,N_19298);
xor U19473 (N_19473,N_19243,N_19259);
nor U19474 (N_19474,N_19246,N_19212);
and U19475 (N_19475,N_19377,N_19211);
nand U19476 (N_19476,N_19394,N_19288);
nor U19477 (N_19477,N_19396,N_19388);
nor U19478 (N_19478,N_19374,N_19365);
or U19479 (N_19479,N_19347,N_19395);
nand U19480 (N_19480,N_19322,N_19389);
nor U19481 (N_19481,N_19223,N_19305);
and U19482 (N_19482,N_19299,N_19254);
or U19483 (N_19483,N_19356,N_19311);
xnor U19484 (N_19484,N_19265,N_19304);
and U19485 (N_19485,N_19392,N_19303);
and U19486 (N_19486,N_19339,N_19390);
xor U19487 (N_19487,N_19237,N_19218);
or U19488 (N_19488,N_19203,N_19257);
nand U19489 (N_19489,N_19329,N_19273);
nor U19490 (N_19490,N_19366,N_19393);
nand U19491 (N_19491,N_19248,N_19338);
or U19492 (N_19492,N_19268,N_19333);
or U19493 (N_19493,N_19279,N_19293);
nor U19494 (N_19494,N_19220,N_19319);
nand U19495 (N_19495,N_19337,N_19226);
nand U19496 (N_19496,N_19292,N_19209);
nand U19497 (N_19497,N_19285,N_19230);
or U19498 (N_19498,N_19316,N_19317);
xor U19499 (N_19499,N_19250,N_19287);
nor U19500 (N_19500,N_19220,N_19206);
xnor U19501 (N_19501,N_19268,N_19285);
nor U19502 (N_19502,N_19315,N_19247);
and U19503 (N_19503,N_19380,N_19343);
or U19504 (N_19504,N_19284,N_19339);
nor U19505 (N_19505,N_19208,N_19309);
and U19506 (N_19506,N_19300,N_19201);
or U19507 (N_19507,N_19388,N_19241);
xnor U19508 (N_19508,N_19354,N_19291);
nor U19509 (N_19509,N_19340,N_19295);
xnor U19510 (N_19510,N_19299,N_19249);
nand U19511 (N_19511,N_19261,N_19380);
and U19512 (N_19512,N_19347,N_19389);
and U19513 (N_19513,N_19378,N_19294);
nor U19514 (N_19514,N_19345,N_19246);
nand U19515 (N_19515,N_19381,N_19203);
xor U19516 (N_19516,N_19388,N_19281);
xnor U19517 (N_19517,N_19298,N_19350);
nand U19518 (N_19518,N_19357,N_19377);
and U19519 (N_19519,N_19384,N_19373);
xor U19520 (N_19520,N_19322,N_19257);
nor U19521 (N_19521,N_19359,N_19289);
or U19522 (N_19522,N_19223,N_19386);
nand U19523 (N_19523,N_19343,N_19272);
xnor U19524 (N_19524,N_19378,N_19375);
and U19525 (N_19525,N_19280,N_19248);
and U19526 (N_19526,N_19349,N_19319);
or U19527 (N_19527,N_19221,N_19399);
nand U19528 (N_19528,N_19319,N_19268);
nor U19529 (N_19529,N_19359,N_19389);
nand U19530 (N_19530,N_19260,N_19214);
nor U19531 (N_19531,N_19325,N_19243);
or U19532 (N_19532,N_19386,N_19337);
nand U19533 (N_19533,N_19255,N_19365);
or U19534 (N_19534,N_19220,N_19275);
or U19535 (N_19535,N_19236,N_19252);
nand U19536 (N_19536,N_19391,N_19278);
or U19537 (N_19537,N_19302,N_19221);
nor U19538 (N_19538,N_19281,N_19334);
and U19539 (N_19539,N_19261,N_19236);
nor U19540 (N_19540,N_19342,N_19328);
and U19541 (N_19541,N_19222,N_19289);
nand U19542 (N_19542,N_19327,N_19304);
or U19543 (N_19543,N_19254,N_19384);
or U19544 (N_19544,N_19298,N_19322);
nand U19545 (N_19545,N_19200,N_19343);
nor U19546 (N_19546,N_19241,N_19267);
xnor U19547 (N_19547,N_19324,N_19355);
or U19548 (N_19548,N_19313,N_19256);
nand U19549 (N_19549,N_19261,N_19213);
xor U19550 (N_19550,N_19301,N_19237);
nand U19551 (N_19551,N_19368,N_19345);
nor U19552 (N_19552,N_19258,N_19376);
nor U19553 (N_19553,N_19299,N_19272);
and U19554 (N_19554,N_19359,N_19201);
and U19555 (N_19555,N_19371,N_19390);
or U19556 (N_19556,N_19261,N_19277);
xnor U19557 (N_19557,N_19340,N_19325);
nand U19558 (N_19558,N_19242,N_19337);
or U19559 (N_19559,N_19368,N_19244);
xnor U19560 (N_19560,N_19396,N_19207);
and U19561 (N_19561,N_19316,N_19330);
nand U19562 (N_19562,N_19362,N_19279);
xor U19563 (N_19563,N_19207,N_19289);
and U19564 (N_19564,N_19214,N_19277);
and U19565 (N_19565,N_19305,N_19374);
nor U19566 (N_19566,N_19335,N_19244);
xor U19567 (N_19567,N_19211,N_19364);
nand U19568 (N_19568,N_19282,N_19272);
xor U19569 (N_19569,N_19227,N_19203);
and U19570 (N_19570,N_19258,N_19277);
and U19571 (N_19571,N_19265,N_19279);
and U19572 (N_19572,N_19361,N_19241);
or U19573 (N_19573,N_19272,N_19312);
nand U19574 (N_19574,N_19223,N_19369);
nand U19575 (N_19575,N_19337,N_19254);
nor U19576 (N_19576,N_19263,N_19275);
nor U19577 (N_19577,N_19387,N_19353);
nor U19578 (N_19578,N_19297,N_19353);
nor U19579 (N_19579,N_19228,N_19316);
nand U19580 (N_19580,N_19307,N_19214);
xnor U19581 (N_19581,N_19212,N_19230);
nor U19582 (N_19582,N_19265,N_19254);
nor U19583 (N_19583,N_19209,N_19362);
xnor U19584 (N_19584,N_19343,N_19248);
nor U19585 (N_19585,N_19274,N_19221);
nand U19586 (N_19586,N_19233,N_19379);
xor U19587 (N_19587,N_19255,N_19371);
xor U19588 (N_19588,N_19358,N_19267);
or U19589 (N_19589,N_19221,N_19213);
or U19590 (N_19590,N_19307,N_19255);
nand U19591 (N_19591,N_19382,N_19397);
nand U19592 (N_19592,N_19283,N_19328);
or U19593 (N_19593,N_19202,N_19257);
nand U19594 (N_19594,N_19236,N_19312);
xor U19595 (N_19595,N_19258,N_19238);
nand U19596 (N_19596,N_19212,N_19381);
and U19597 (N_19597,N_19366,N_19260);
xnor U19598 (N_19598,N_19215,N_19325);
xor U19599 (N_19599,N_19284,N_19399);
xnor U19600 (N_19600,N_19598,N_19499);
nor U19601 (N_19601,N_19543,N_19548);
or U19602 (N_19602,N_19433,N_19466);
nand U19603 (N_19603,N_19498,N_19444);
nand U19604 (N_19604,N_19468,N_19490);
nor U19605 (N_19605,N_19539,N_19436);
xor U19606 (N_19606,N_19537,N_19551);
or U19607 (N_19607,N_19536,N_19530);
xnor U19608 (N_19608,N_19420,N_19587);
or U19609 (N_19609,N_19467,N_19592);
nand U19610 (N_19610,N_19505,N_19478);
xnor U19611 (N_19611,N_19559,N_19406);
xor U19612 (N_19612,N_19589,N_19486);
nand U19613 (N_19613,N_19535,N_19462);
or U19614 (N_19614,N_19469,N_19400);
xnor U19615 (N_19615,N_19407,N_19540);
nor U19616 (N_19616,N_19402,N_19561);
xor U19617 (N_19617,N_19558,N_19541);
and U19618 (N_19618,N_19480,N_19445);
and U19619 (N_19619,N_19545,N_19446);
or U19620 (N_19620,N_19451,N_19557);
nand U19621 (N_19621,N_19572,N_19487);
nor U19622 (N_19622,N_19597,N_19524);
and U19623 (N_19623,N_19410,N_19426);
xor U19624 (N_19624,N_19404,N_19501);
or U19625 (N_19625,N_19447,N_19482);
and U19626 (N_19626,N_19519,N_19474);
or U19627 (N_19627,N_19494,N_19599);
and U19628 (N_19628,N_19416,N_19405);
xnor U19629 (N_19629,N_19595,N_19522);
or U19630 (N_19630,N_19514,N_19517);
or U19631 (N_19631,N_19431,N_19528);
nor U19632 (N_19632,N_19504,N_19588);
nand U19633 (N_19633,N_19434,N_19428);
or U19634 (N_19634,N_19585,N_19508);
nand U19635 (N_19635,N_19593,N_19497);
and U19636 (N_19636,N_19571,N_19526);
nand U19637 (N_19637,N_19429,N_19415);
xor U19638 (N_19638,N_19565,N_19430);
and U19639 (N_19639,N_19542,N_19584);
nor U19640 (N_19640,N_19529,N_19552);
and U19641 (N_19641,N_19596,N_19534);
xnor U19642 (N_19642,N_19417,N_19531);
and U19643 (N_19643,N_19579,N_19586);
nand U19644 (N_19644,N_19450,N_19456);
xnor U19645 (N_19645,N_19509,N_19567);
nor U19646 (N_19646,N_19566,N_19577);
nor U19647 (N_19647,N_19513,N_19488);
nor U19648 (N_19648,N_19570,N_19510);
or U19649 (N_19649,N_19581,N_19483);
xnor U19650 (N_19650,N_19470,N_19441);
or U19651 (N_19651,N_19560,N_19403);
and U19652 (N_19652,N_19465,N_19527);
and U19653 (N_19653,N_19550,N_19472);
nor U19654 (N_19654,N_19575,N_19496);
nand U19655 (N_19655,N_19547,N_19582);
xnor U19656 (N_19656,N_19518,N_19481);
and U19657 (N_19657,N_19573,N_19440);
nor U19658 (N_19658,N_19435,N_19553);
and U19659 (N_19659,N_19473,N_19515);
xor U19660 (N_19660,N_19424,N_19413);
nand U19661 (N_19661,N_19564,N_19562);
xnor U19662 (N_19662,N_19507,N_19459);
nor U19663 (N_19663,N_19448,N_19576);
nand U19664 (N_19664,N_19516,N_19411);
or U19665 (N_19665,N_19484,N_19432);
xor U19666 (N_19666,N_19418,N_19457);
nor U19667 (N_19667,N_19438,N_19549);
nand U19668 (N_19668,N_19476,N_19439);
or U19669 (N_19669,N_19533,N_19464);
nand U19670 (N_19670,N_19409,N_19555);
and U19671 (N_19671,N_19475,N_19554);
and U19672 (N_19672,N_19512,N_19563);
nor U19673 (N_19673,N_19492,N_19454);
or U19674 (N_19674,N_19412,N_19449);
nand U19675 (N_19675,N_19401,N_19463);
nor U19676 (N_19676,N_19422,N_19442);
nor U19677 (N_19677,N_19591,N_19511);
nand U19678 (N_19678,N_19455,N_19520);
and U19679 (N_19679,N_19479,N_19525);
nor U19680 (N_19680,N_19502,N_19521);
and U19681 (N_19681,N_19532,N_19461);
xnor U19682 (N_19682,N_19569,N_19568);
nand U19683 (N_19683,N_19538,N_19523);
and U19684 (N_19684,N_19590,N_19506);
nand U19685 (N_19685,N_19500,N_19594);
or U19686 (N_19686,N_19458,N_19556);
nand U19687 (N_19687,N_19421,N_19578);
or U19688 (N_19688,N_19460,N_19546);
xnor U19689 (N_19689,N_19437,N_19453);
and U19690 (N_19690,N_19423,N_19580);
xnor U19691 (N_19691,N_19503,N_19583);
and U19692 (N_19692,N_19574,N_19485);
and U19693 (N_19693,N_19452,N_19491);
nand U19694 (N_19694,N_19471,N_19493);
nand U19695 (N_19695,N_19414,N_19544);
and U19696 (N_19696,N_19489,N_19495);
nor U19697 (N_19697,N_19443,N_19408);
nand U19698 (N_19698,N_19427,N_19419);
xnor U19699 (N_19699,N_19425,N_19477);
nand U19700 (N_19700,N_19489,N_19548);
xor U19701 (N_19701,N_19487,N_19523);
xor U19702 (N_19702,N_19499,N_19454);
xor U19703 (N_19703,N_19590,N_19587);
nand U19704 (N_19704,N_19475,N_19435);
nand U19705 (N_19705,N_19467,N_19405);
xor U19706 (N_19706,N_19534,N_19517);
nand U19707 (N_19707,N_19515,N_19504);
nor U19708 (N_19708,N_19416,N_19553);
and U19709 (N_19709,N_19476,N_19494);
nand U19710 (N_19710,N_19491,N_19522);
nor U19711 (N_19711,N_19599,N_19581);
nand U19712 (N_19712,N_19438,N_19539);
or U19713 (N_19713,N_19563,N_19561);
or U19714 (N_19714,N_19453,N_19578);
xor U19715 (N_19715,N_19487,N_19597);
nand U19716 (N_19716,N_19566,N_19481);
and U19717 (N_19717,N_19584,N_19453);
nand U19718 (N_19718,N_19509,N_19570);
nand U19719 (N_19719,N_19573,N_19418);
nor U19720 (N_19720,N_19506,N_19584);
nor U19721 (N_19721,N_19420,N_19536);
xor U19722 (N_19722,N_19534,N_19536);
nand U19723 (N_19723,N_19583,N_19514);
nor U19724 (N_19724,N_19447,N_19545);
and U19725 (N_19725,N_19472,N_19455);
nor U19726 (N_19726,N_19401,N_19421);
and U19727 (N_19727,N_19548,N_19529);
xnor U19728 (N_19728,N_19598,N_19439);
nor U19729 (N_19729,N_19578,N_19482);
xnor U19730 (N_19730,N_19489,N_19424);
xnor U19731 (N_19731,N_19515,N_19583);
nand U19732 (N_19732,N_19558,N_19493);
or U19733 (N_19733,N_19526,N_19543);
and U19734 (N_19734,N_19511,N_19557);
xor U19735 (N_19735,N_19531,N_19544);
nand U19736 (N_19736,N_19527,N_19493);
nand U19737 (N_19737,N_19491,N_19424);
or U19738 (N_19738,N_19574,N_19436);
xor U19739 (N_19739,N_19576,N_19484);
nand U19740 (N_19740,N_19510,N_19425);
and U19741 (N_19741,N_19469,N_19545);
xnor U19742 (N_19742,N_19445,N_19444);
and U19743 (N_19743,N_19508,N_19509);
nor U19744 (N_19744,N_19519,N_19426);
or U19745 (N_19745,N_19434,N_19587);
or U19746 (N_19746,N_19447,N_19408);
xnor U19747 (N_19747,N_19574,N_19576);
nor U19748 (N_19748,N_19598,N_19599);
xnor U19749 (N_19749,N_19504,N_19556);
nor U19750 (N_19750,N_19586,N_19464);
nand U19751 (N_19751,N_19436,N_19408);
nor U19752 (N_19752,N_19475,N_19425);
and U19753 (N_19753,N_19465,N_19501);
nand U19754 (N_19754,N_19589,N_19543);
and U19755 (N_19755,N_19583,N_19529);
and U19756 (N_19756,N_19494,N_19536);
nor U19757 (N_19757,N_19573,N_19422);
nand U19758 (N_19758,N_19471,N_19485);
or U19759 (N_19759,N_19597,N_19491);
or U19760 (N_19760,N_19587,N_19453);
xnor U19761 (N_19761,N_19512,N_19459);
nor U19762 (N_19762,N_19502,N_19593);
nor U19763 (N_19763,N_19517,N_19593);
nand U19764 (N_19764,N_19508,N_19449);
nand U19765 (N_19765,N_19589,N_19467);
and U19766 (N_19766,N_19446,N_19523);
or U19767 (N_19767,N_19535,N_19599);
or U19768 (N_19768,N_19597,N_19579);
nand U19769 (N_19769,N_19489,N_19456);
nand U19770 (N_19770,N_19542,N_19582);
and U19771 (N_19771,N_19508,N_19534);
or U19772 (N_19772,N_19521,N_19583);
or U19773 (N_19773,N_19587,N_19526);
nand U19774 (N_19774,N_19576,N_19519);
nor U19775 (N_19775,N_19487,N_19563);
nand U19776 (N_19776,N_19444,N_19559);
xnor U19777 (N_19777,N_19534,N_19495);
nand U19778 (N_19778,N_19580,N_19447);
xor U19779 (N_19779,N_19437,N_19424);
or U19780 (N_19780,N_19462,N_19512);
nand U19781 (N_19781,N_19438,N_19565);
and U19782 (N_19782,N_19487,N_19440);
or U19783 (N_19783,N_19460,N_19556);
and U19784 (N_19784,N_19492,N_19450);
nand U19785 (N_19785,N_19464,N_19585);
and U19786 (N_19786,N_19549,N_19436);
nand U19787 (N_19787,N_19532,N_19458);
xnor U19788 (N_19788,N_19558,N_19484);
and U19789 (N_19789,N_19498,N_19404);
xnor U19790 (N_19790,N_19567,N_19487);
nor U19791 (N_19791,N_19515,N_19534);
nand U19792 (N_19792,N_19577,N_19428);
nor U19793 (N_19793,N_19402,N_19429);
nor U19794 (N_19794,N_19495,N_19562);
or U19795 (N_19795,N_19535,N_19470);
xnor U19796 (N_19796,N_19488,N_19546);
nand U19797 (N_19797,N_19515,N_19407);
nand U19798 (N_19798,N_19578,N_19535);
nand U19799 (N_19799,N_19584,N_19439);
or U19800 (N_19800,N_19752,N_19649);
nor U19801 (N_19801,N_19665,N_19782);
and U19802 (N_19802,N_19628,N_19681);
or U19803 (N_19803,N_19641,N_19619);
or U19804 (N_19804,N_19621,N_19609);
xor U19805 (N_19805,N_19695,N_19618);
xnor U19806 (N_19806,N_19678,N_19707);
or U19807 (N_19807,N_19722,N_19690);
nand U19808 (N_19808,N_19684,N_19749);
xnor U19809 (N_19809,N_19734,N_19640);
and U19810 (N_19810,N_19719,N_19625);
or U19811 (N_19811,N_19645,N_19666);
xor U19812 (N_19812,N_19655,N_19693);
nand U19813 (N_19813,N_19703,N_19731);
nand U19814 (N_19814,N_19688,N_19664);
and U19815 (N_19815,N_19616,N_19667);
and U19816 (N_19816,N_19783,N_19786);
or U19817 (N_19817,N_19697,N_19622);
and U19818 (N_19818,N_19714,N_19698);
xnor U19819 (N_19819,N_19632,N_19745);
nor U19820 (N_19820,N_19612,N_19699);
nor U19821 (N_19821,N_19751,N_19735);
or U19822 (N_19822,N_19663,N_19738);
or U19823 (N_19823,N_19636,N_19706);
or U19824 (N_19824,N_19670,N_19650);
nor U19825 (N_19825,N_19773,N_19737);
nand U19826 (N_19826,N_19654,N_19617);
nand U19827 (N_19827,N_19740,N_19794);
xor U19828 (N_19828,N_19653,N_19607);
or U19829 (N_19829,N_19652,N_19713);
nand U19830 (N_19830,N_19605,N_19717);
nand U19831 (N_19831,N_19730,N_19774);
nand U19832 (N_19832,N_19798,N_19762);
or U19833 (N_19833,N_19742,N_19658);
nand U19834 (N_19834,N_19767,N_19696);
and U19835 (N_19835,N_19610,N_19766);
nand U19836 (N_19836,N_19614,N_19765);
nand U19837 (N_19837,N_19729,N_19631);
or U19838 (N_19838,N_19602,N_19779);
or U19839 (N_19839,N_19680,N_19781);
and U19840 (N_19840,N_19686,N_19700);
nor U19841 (N_19841,N_19732,N_19685);
nand U19842 (N_19842,N_19637,N_19701);
xnor U19843 (N_19843,N_19676,N_19736);
or U19844 (N_19844,N_19630,N_19764);
nor U19845 (N_19845,N_19741,N_19760);
and U19846 (N_19846,N_19604,N_19721);
or U19847 (N_19847,N_19739,N_19600);
nor U19848 (N_19848,N_19727,N_19776);
xor U19849 (N_19849,N_19635,N_19708);
nand U19850 (N_19850,N_19788,N_19753);
nand U19851 (N_19851,N_19709,N_19763);
and U19852 (N_19852,N_19692,N_19629);
nand U19853 (N_19853,N_19675,N_19743);
xnor U19854 (N_19854,N_19711,N_19647);
xor U19855 (N_19855,N_19777,N_19646);
nor U19856 (N_19856,N_19672,N_19780);
or U19857 (N_19857,N_19784,N_19728);
or U19858 (N_19858,N_19657,N_19793);
nand U19859 (N_19859,N_19673,N_19620);
and U19860 (N_19860,N_19785,N_19603);
nor U19861 (N_19861,N_19613,N_19694);
nand U19862 (N_19862,N_19661,N_19660);
xor U19863 (N_19863,N_19789,N_19691);
and U19864 (N_19864,N_19687,N_19758);
or U19865 (N_19865,N_19725,N_19795);
and U19866 (N_19866,N_19626,N_19643);
and U19867 (N_19867,N_19677,N_19770);
or U19868 (N_19868,N_19796,N_19601);
and U19869 (N_19869,N_19651,N_19790);
xnor U19870 (N_19870,N_19791,N_19683);
nor U19871 (N_19871,N_19748,N_19799);
xor U19872 (N_19872,N_19689,N_19744);
nand U19873 (N_19873,N_19669,N_19775);
nand U19874 (N_19874,N_19797,N_19787);
or U19875 (N_19875,N_19750,N_19715);
and U19876 (N_19876,N_19756,N_19716);
nand U19877 (N_19877,N_19623,N_19724);
xor U19878 (N_19878,N_19634,N_19648);
and U19879 (N_19879,N_19772,N_19726);
nand U19880 (N_19880,N_19705,N_19682);
nand U19881 (N_19881,N_19778,N_19642);
nand U19882 (N_19882,N_19662,N_19768);
and U19883 (N_19883,N_19608,N_19712);
and U19884 (N_19884,N_19679,N_19761);
or U19885 (N_19885,N_19624,N_19615);
nand U19886 (N_19886,N_19723,N_19759);
xor U19887 (N_19887,N_19674,N_19668);
and U19888 (N_19888,N_19733,N_19792);
nand U19889 (N_19889,N_19639,N_19769);
nand U19890 (N_19890,N_19771,N_19718);
xor U19891 (N_19891,N_19656,N_19754);
nand U19892 (N_19892,N_19746,N_19720);
nand U19893 (N_19893,N_19638,N_19702);
nor U19894 (N_19894,N_19710,N_19755);
or U19895 (N_19895,N_19644,N_19747);
or U19896 (N_19896,N_19611,N_19704);
nor U19897 (N_19897,N_19627,N_19606);
and U19898 (N_19898,N_19671,N_19659);
or U19899 (N_19899,N_19633,N_19757);
xnor U19900 (N_19900,N_19775,N_19614);
and U19901 (N_19901,N_19791,N_19703);
or U19902 (N_19902,N_19627,N_19610);
and U19903 (N_19903,N_19723,N_19727);
nand U19904 (N_19904,N_19647,N_19694);
and U19905 (N_19905,N_19755,N_19745);
and U19906 (N_19906,N_19756,N_19661);
nor U19907 (N_19907,N_19649,N_19724);
and U19908 (N_19908,N_19794,N_19631);
or U19909 (N_19909,N_19706,N_19799);
or U19910 (N_19910,N_19749,N_19656);
or U19911 (N_19911,N_19790,N_19625);
or U19912 (N_19912,N_19685,N_19627);
nand U19913 (N_19913,N_19734,N_19799);
nor U19914 (N_19914,N_19613,N_19727);
and U19915 (N_19915,N_19668,N_19693);
or U19916 (N_19916,N_19616,N_19610);
and U19917 (N_19917,N_19763,N_19751);
or U19918 (N_19918,N_19797,N_19611);
nor U19919 (N_19919,N_19659,N_19763);
nor U19920 (N_19920,N_19634,N_19610);
xnor U19921 (N_19921,N_19670,N_19704);
nand U19922 (N_19922,N_19766,N_19616);
nand U19923 (N_19923,N_19704,N_19706);
nand U19924 (N_19924,N_19700,N_19767);
and U19925 (N_19925,N_19746,N_19747);
nand U19926 (N_19926,N_19647,N_19754);
and U19927 (N_19927,N_19631,N_19616);
nor U19928 (N_19928,N_19680,N_19724);
and U19929 (N_19929,N_19766,N_19647);
and U19930 (N_19930,N_19731,N_19791);
or U19931 (N_19931,N_19779,N_19653);
or U19932 (N_19932,N_19660,N_19799);
xor U19933 (N_19933,N_19625,N_19779);
nor U19934 (N_19934,N_19677,N_19742);
or U19935 (N_19935,N_19714,N_19635);
nand U19936 (N_19936,N_19656,N_19669);
and U19937 (N_19937,N_19610,N_19726);
nor U19938 (N_19938,N_19763,N_19621);
and U19939 (N_19939,N_19698,N_19700);
nand U19940 (N_19940,N_19659,N_19734);
and U19941 (N_19941,N_19713,N_19664);
or U19942 (N_19942,N_19676,N_19773);
nor U19943 (N_19943,N_19773,N_19770);
xor U19944 (N_19944,N_19617,N_19600);
nor U19945 (N_19945,N_19661,N_19766);
nor U19946 (N_19946,N_19694,N_19677);
nand U19947 (N_19947,N_19711,N_19666);
and U19948 (N_19948,N_19790,N_19742);
or U19949 (N_19949,N_19792,N_19773);
nor U19950 (N_19950,N_19658,N_19678);
nand U19951 (N_19951,N_19656,N_19621);
nor U19952 (N_19952,N_19682,N_19718);
and U19953 (N_19953,N_19773,N_19704);
nor U19954 (N_19954,N_19656,N_19775);
xnor U19955 (N_19955,N_19691,N_19676);
nand U19956 (N_19956,N_19683,N_19680);
nor U19957 (N_19957,N_19634,N_19689);
or U19958 (N_19958,N_19794,N_19713);
nand U19959 (N_19959,N_19714,N_19719);
and U19960 (N_19960,N_19678,N_19757);
nand U19961 (N_19961,N_19665,N_19755);
nor U19962 (N_19962,N_19771,N_19760);
nand U19963 (N_19963,N_19623,N_19688);
nor U19964 (N_19964,N_19600,N_19652);
and U19965 (N_19965,N_19638,N_19645);
or U19966 (N_19966,N_19769,N_19723);
nor U19967 (N_19967,N_19749,N_19730);
xnor U19968 (N_19968,N_19673,N_19665);
nor U19969 (N_19969,N_19704,N_19751);
nand U19970 (N_19970,N_19659,N_19648);
xnor U19971 (N_19971,N_19708,N_19752);
nand U19972 (N_19972,N_19787,N_19666);
nor U19973 (N_19973,N_19645,N_19664);
or U19974 (N_19974,N_19638,N_19720);
xnor U19975 (N_19975,N_19737,N_19742);
nand U19976 (N_19976,N_19670,N_19794);
xnor U19977 (N_19977,N_19724,N_19685);
xnor U19978 (N_19978,N_19762,N_19734);
nand U19979 (N_19979,N_19771,N_19794);
xor U19980 (N_19980,N_19664,N_19629);
and U19981 (N_19981,N_19760,N_19688);
nor U19982 (N_19982,N_19679,N_19672);
xor U19983 (N_19983,N_19785,N_19657);
xor U19984 (N_19984,N_19753,N_19791);
nand U19985 (N_19985,N_19687,N_19767);
and U19986 (N_19986,N_19610,N_19784);
nor U19987 (N_19987,N_19641,N_19656);
and U19988 (N_19988,N_19703,N_19629);
nand U19989 (N_19989,N_19739,N_19706);
nor U19990 (N_19990,N_19604,N_19600);
or U19991 (N_19991,N_19663,N_19725);
nand U19992 (N_19992,N_19776,N_19662);
nand U19993 (N_19993,N_19721,N_19767);
or U19994 (N_19994,N_19686,N_19735);
xor U19995 (N_19995,N_19752,N_19775);
or U19996 (N_19996,N_19661,N_19762);
nand U19997 (N_19997,N_19785,N_19668);
nor U19998 (N_19998,N_19636,N_19617);
nor U19999 (N_19999,N_19640,N_19777);
or UO_0 (O_0,N_19965,N_19899);
nor UO_1 (O_1,N_19968,N_19889);
and UO_2 (O_2,N_19905,N_19868);
and UO_3 (O_3,N_19919,N_19835);
nor UO_4 (O_4,N_19870,N_19819);
or UO_5 (O_5,N_19849,N_19853);
nand UO_6 (O_6,N_19814,N_19976);
xor UO_7 (O_7,N_19990,N_19854);
or UO_8 (O_8,N_19820,N_19979);
or UO_9 (O_9,N_19852,N_19871);
nand UO_10 (O_10,N_19892,N_19865);
xnor UO_11 (O_11,N_19827,N_19898);
and UO_12 (O_12,N_19881,N_19817);
nor UO_13 (O_13,N_19867,N_19974);
or UO_14 (O_14,N_19945,N_19913);
nor UO_15 (O_15,N_19863,N_19877);
or UO_16 (O_16,N_19900,N_19930);
nand UO_17 (O_17,N_19934,N_19918);
nor UO_18 (O_18,N_19925,N_19878);
or UO_19 (O_19,N_19922,N_19843);
nor UO_20 (O_20,N_19887,N_19997);
and UO_21 (O_21,N_19987,N_19837);
xor UO_22 (O_22,N_19811,N_19932);
and UO_23 (O_23,N_19917,N_19908);
nor UO_24 (O_24,N_19986,N_19864);
xor UO_25 (O_25,N_19935,N_19904);
nor UO_26 (O_26,N_19812,N_19903);
xnor UO_27 (O_27,N_19801,N_19906);
and UO_28 (O_28,N_19909,N_19857);
nor UO_29 (O_29,N_19882,N_19886);
nor UO_30 (O_30,N_19995,N_19933);
and UO_31 (O_31,N_19879,N_19858);
xor UO_32 (O_32,N_19959,N_19901);
and UO_33 (O_33,N_19893,N_19891);
or UO_34 (O_34,N_19821,N_19920);
nand UO_35 (O_35,N_19880,N_19941);
xor UO_36 (O_36,N_19961,N_19834);
nand UO_37 (O_37,N_19947,N_19824);
or UO_38 (O_38,N_19815,N_19938);
and UO_39 (O_39,N_19829,N_19943);
xnor UO_40 (O_40,N_19856,N_19890);
xnor UO_41 (O_41,N_19942,N_19805);
nand UO_42 (O_42,N_19855,N_19822);
nor UO_43 (O_43,N_19874,N_19931);
nand UO_44 (O_44,N_19842,N_19888);
nand UO_45 (O_45,N_19911,N_19948);
or UO_46 (O_46,N_19956,N_19989);
xnor UO_47 (O_47,N_19894,N_19924);
nand UO_48 (O_48,N_19912,N_19973);
nor UO_49 (O_49,N_19929,N_19847);
xor UO_50 (O_50,N_19826,N_19993);
nand UO_51 (O_51,N_19915,N_19872);
and UO_52 (O_52,N_19895,N_19982);
nand UO_53 (O_53,N_19960,N_19970);
xnor UO_54 (O_54,N_19830,N_19996);
nand UO_55 (O_55,N_19946,N_19839);
or UO_56 (O_56,N_19980,N_19955);
nand UO_57 (O_57,N_19952,N_19937);
nand UO_58 (O_58,N_19949,N_19806);
and UO_59 (O_59,N_19950,N_19985);
xor UO_60 (O_60,N_19988,N_19969);
or UO_61 (O_61,N_19992,N_19964);
or UO_62 (O_62,N_19954,N_19999);
or UO_63 (O_63,N_19963,N_19838);
and UO_64 (O_64,N_19923,N_19828);
nand UO_65 (O_65,N_19846,N_19841);
nor UO_66 (O_66,N_19875,N_19994);
nand UO_67 (O_67,N_19951,N_19831);
nand UO_68 (O_68,N_19818,N_19802);
and UO_69 (O_69,N_19896,N_19800);
and UO_70 (O_70,N_19957,N_19884);
nor UO_71 (O_71,N_19971,N_19803);
nand UO_72 (O_72,N_19809,N_19869);
nand UO_73 (O_73,N_19866,N_19914);
or UO_74 (O_74,N_19984,N_19958);
xor UO_75 (O_75,N_19808,N_19998);
nand UO_76 (O_76,N_19836,N_19833);
and UO_77 (O_77,N_19897,N_19907);
or UO_78 (O_78,N_19848,N_19940);
xor UO_79 (O_79,N_19804,N_19807);
or UO_80 (O_80,N_19936,N_19910);
or UO_81 (O_81,N_19859,N_19953);
or UO_82 (O_82,N_19977,N_19832);
nand UO_83 (O_83,N_19981,N_19816);
nand UO_84 (O_84,N_19823,N_19862);
or UO_85 (O_85,N_19972,N_19883);
xnor UO_86 (O_86,N_19885,N_19810);
or UO_87 (O_87,N_19966,N_19962);
and UO_88 (O_88,N_19840,N_19975);
or UO_89 (O_89,N_19928,N_19902);
xnor UO_90 (O_90,N_19944,N_19967);
nand UO_91 (O_91,N_19978,N_19860);
nand UO_92 (O_92,N_19844,N_19851);
nand UO_93 (O_93,N_19926,N_19873);
xnor UO_94 (O_94,N_19813,N_19991);
xnor UO_95 (O_95,N_19916,N_19861);
nand UO_96 (O_96,N_19825,N_19983);
or UO_97 (O_97,N_19921,N_19939);
and UO_98 (O_98,N_19927,N_19876);
nor UO_99 (O_99,N_19845,N_19850);
xnor UO_100 (O_100,N_19822,N_19940);
nand UO_101 (O_101,N_19817,N_19987);
nor UO_102 (O_102,N_19886,N_19951);
nor UO_103 (O_103,N_19942,N_19947);
xor UO_104 (O_104,N_19820,N_19983);
xor UO_105 (O_105,N_19852,N_19997);
xor UO_106 (O_106,N_19944,N_19875);
nor UO_107 (O_107,N_19862,N_19958);
nand UO_108 (O_108,N_19830,N_19813);
and UO_109 (O_109,N_19884,N_19909);
nand UO_110 (O_110,N_19846,N_19869);
nor UO_111 (O_111,N_19999,N_19946);
and UO_112 (O_112,N_19976,N_19807);
xnor UO_113 (O_113,N_19982,N_19939);
or UO_114 (O_114,N_19959,N_19955);
xnor UO_115 (O_115,N_19887,N_19964);
xor UO_116 (O_116,N_19904,N_19979);
nand UO_117 (O_117,N_19932,N_19926);
xnor UO_118 (O_118,N_19918,N_19972);
and UO_119 (O_119,N_19835,N_19972);
and UO_120 (O_120,N_19852,N_19944);
or UO_121 (O_121,N_19968,N_19960);
or UO_122 (O_122,N_19957,N_19922);
or UO_123 (O_123,N_19833,N_19925);
or UO_124 (O_124,N_19932,N_19896);
xnor UO_125 (O_125,N_19859,N_19911);
or UO_126 (O_126,N_19815,N_19911);
nor UO_127 (O_127,N_19990,N_19964);
nor UO_128 (O_128,N_19914,N_19861);
or UO_129 (O_129,N_19903,N_19883);
and UO_130 (O_130,N_19924,N_19952);
nand UO_131 (O_131,N_19845,N_19935);
and UO_132 (O_132,N_19945,N_19981);
or UO_133 (O_133,N_19835,N_19915);
and UO_134 (O_134,N_19956,N_19855);
xnor UO_135 (O_135,N_19988,N_19887);
and UO_136 (O_136,N_19817,N_19962);
xor UO_137 (O_137,N_19865,N_19942);
xnor UO_138 (O_138,N_19841,N_19938);
and UO_139 (O_139,N_19916,N_19935);
xnor UO_140 (O_140,N_19808,N_19890);
xor UO_141 (O_141,N_19835,N_19983);
and UO_142 (O_142,N_19866,N_19842);
or UO_143 (O_143,N_19809,N_19850);
and UO_144 (O_144,N_19873,N_19975);
nor UO_145 (O_145,N_19848,N_19903);
and UO_146 (O_146,N_19886,N_19958);
or UO_147 (O_147,N_19912,N_19891);
or UO_148 (O_148,N_19830,N_19995);
xor UO_149 (O_149,N_19943,N_19804);
or UO_150 (O_150,N_19963,N_19904);
nand UO_151 (O_151,N_19973,N_19827);
or UO_152 (O_152,N_19987,N_19916);
and UO_153 (O_153,N_19973,N_19895);
xnor UO_154 (O_154,N_19958,N_19957);
nand UO_155 (O_155,N_19850,N_19961);
and UO_156 (O_156,N_19908,N_19857);
nor UO_157 (O_157,N_19813,N_19955);
nand UO_158 (O_158,N_19866,N_19975);
nor UO_159 (O_159,N_19952,N_19814);
and UO_160 (O_160,N_19943,N_19888);
or UO_161 (O_161,N_19853,N_19936);
nor UO_162 (O_162,N_19817,N_19960);
nor UO_163 (O_163,N_19929,N_19933);
nand UO_164 (O_164,N_19864,N_19968);
xnor UO_165 (O_165,N_19819,N_19833);
and UO_166 (O_166,N_19824,N_19831);
nand UO_167 (O_167,N_19913,N_19853);
nor UO_168 (O_168,N_19868,N_19892);
nor UO_169 (O_169,N_19970,N_19815);
and UO_170 (O_170,N_19911,N_19917);
xnor UO_171 (O_171,N_19810,N_19804);
and UO_172 (O_172,N_19826,N_19959);
nor UO_173 (O_173,N_19945,N_19917);
and UO_174 (O_174,N_19949,N_19819);
or UO_175 (O_175,N_19889,N_19869);
nand UO_176 (O_176,N_19880,N_19979);
xnor UO_177 (O_177,N_19906,N_19985);
or UO_178 (O_178,N_19837,N_19887);
or UO_179 (O_179,N_19925,N_19840);
nand UO_180 (O_180,N_19902,N_19854);
and UO_181 (O_181,N_19859,N_19956);
and UO_182 (O_182,N_19822,N_19952);
nor UO_183 (O_183,N_19984,N_19901);
nor UO_184 (O_184,N_19959,N_19956);
nand UO_185 (O_185,N_19974,N_19894);
nand UO_186 (O_186,N_19824,N_19891);
or UO_187 (O_187,N_19815,N_19916);
xor UO_188 (O_188,N_19995,N_19993);
or UO_189 (O_189,N_19852,N_19981);
and UO_190 (O_190,N_19840,N_19801);
or UO_191 (O_191,N_19991,N_19823);
xnor UO_192 (O_192,N_19884,N_19890);
nor UO_193 (O_193,N_19906,N_19819);
nor UO_194 (O_194,N_19971,N_19840);
or UO_195 (O_195,N_19917,N_19948);
nand UO_196 (O_196,N_19935,N_19858);
nand UO_197 (O_197,N_19831,N_19990);
xnor UO_198 (O_198,N_19954,N_19961);
xnor UO_199 (O_199,N_19984,N_19871);
or UO_200 (O_200,N_19937,N_19894);
and UO_201 (O_201,N_19916,N_19936);
and UO_202 (O_202,N_19869,N_19978);
nor UO_203 (O_203,N_19822,N_19968);
nor UO_204 (O_204,N_19861,N_19929);
nand UO_205 (O_205,N_19873,N_19901);
or UO_206 (O_206,N_19843,N_19985);
nand UO_207 (O_207,N_19943,N_19833);
nand UO_208 (O_208,N_19810,N_19892);
and UO_209 (O_209,N_19989,N_19945);
xnor UO_210 (O_210,N_19971,N_19907);
nor UO_211 (O_211,N_19923,N_19829);
nor UO_212 (O_212,N_19852,N_19835);
or UO_213 (O_213,N_19937,N_19877);
or UO_214 (O_214,N_19966,N_19975);
and UO_215 (O_215,N_19897,N_19856);
xor UO_216 (O_216,N_19958,N_19817);
nor UO_217 (O_217,N_19939,N_19936);
nor UO_218 (O_218,N_19891,N_19809);
or UO_219 (O_219,N_19890,N_19813);
and UO_220 (O_220,N_19992,N_19892);
xnor UO_221 (O_221,N_19865,N_19946);
xnor UO_222 (O_222,N_19917,N_19806);
nor UO_223 (O_223,N_19933,N_19856);
xnor UO_224 (O_224,N_19843,N_19873);
and UO_225 (O_225,N_19849,N_19907);
and UO_226 (O_226,N_19823,N_19895);
xnor UO_227 (O_227,N_19831,N_19844);
nor UO_228 (O_228,N_19985,N_19932);
nand UO_229 (O_229,N_19846,N_19854);
or UO_230 (O_230,N_19856,N_19957);
nand UO_231 (O_231,N_19938,N_19985);
and UO_232 (O_232,N_19851,N_19826);
xor UO_233 (O_233,N_19885,N_19814);
and UO_234 (O_234,N_19890,N_19958);
xnor UO_235 (O_235,N_19848,N_19970);
xnor UO_236 (O_236,N_19902,N_19820);
xnor UO_237 (O_237,N_19833,N_19953);
or UO_238 (O_238,N_19888,N_19806);
and UO_239 (O_239,N_19805,N_19883);
nand UO_240 (O_240,N_19818,N_19834);
and UO_241 (O_241,N_19842,N_19910);
nand UO_242 (O_242,N_19924,N_19971);
and UO_243 (O_243,N_19885,N_19942);
nand UO_244 (O_244,N_19943,N_19878);
or UO_245 (O_245,N_19815,N_19885);
and UO_246 (O_246,N_19849,N_19942);
nand UO_247 (O_247,N_19872,N_19939);
xor UO_248 (O_248,N_19847,N_19943);
nor UO_249 (O_249,N_19935,N_19961);
nor UO_250 (O_250,N_19984,N_19935);
nand UO_251 (O_251,N_19966,N_19849);
and UO_252 (O_252,N_19841,N_19880);
nor UO_253 (O_253,N_19871,N_19966);
nand UO_254 (O_254,N_19939,N_19915);
nor UO_255 (O_255,N_19937,N_19822);
xnor UO_256 (O_256,N_19933,N_19809);
or UO_257 (O_257,N_19838,N_19920);
and UO_258 (O_258,N_19970,N_19817);
and UO_259 (O_259,N_19811,N_19921);
or UO_260 (O_260,N_19997,N_19857);
xnor UO_261 (O_261,N_19972,N_19955);
and UO_262 (O_262,N_19801,N_19871);
nand UO_263 (O_263,N_19924,N_19998);
and UO_264 (O_264,N_19936,N_19988);
or UO_265 (O_265,N_19996,N_19843);
or UO_266 (O_266,N_19924,N_19821);
or UO_267 (O_267,N_19833,N_19807);
nand UO_268 (O_268,N_19910,N_19808);
xor UO_269 (O_269,N_19867,N_19914);
or UO_270 (O_270,N_19940,N_19922);
and UO_271 (O_271,N_19975,N_19904);
xnor UO_272 (O_272,N_19936,N_19989);
and UO_273 (O_273,N_19868,N_19872);
or UO_274 (O_274,N_19998,N_19999);
nand UO_275 (O_275,N_19975,N_19836);
or UO_276 (O_276,N_19806,N_19941);
xor UO_277 (O_277,N_19903,N_19975);
nor UO_278 (O_278,N_19876,N_19922);
nand UO_279 (O_279,N_19984,N_19803);
xnor UO_280 (O_280,N_19868,N_19869);
nand UO_281 (O_281,N_19867,N_19917);
and UO_282 (O_282,N_19947,N_19896);
nand UO_283 (O_283,N_19950,N_19940);
and UO_284 (O_284,N_19973,N_19967);
xor UO_285 (O_285,N_19984,N_19995);
nand UO_286 (O_286,N_19838,N_19822);
xor UO_287 (O_287,N_19973,N_19892);
or UO_288 (O_288,N_19883,N_19899);
nor UO_289 (O_289,N_19938,N_19892);
or UO_290 (O_290,N_19834,N_19957);
nand UO_291 (O_291,N_19831,N_19920);
xor UO_292 (O_292,N_19824,N_19848);
or UO_293 (O_293,N_19953,N_19834);
and UO_294 (O_294,N_19811,N_19927);
nor UO_295 (O_295,N_19806,N_19910);
nor UO_296 (O_296,N_19977,N_19848);
nor UO_297 (O_297,N_19902,N_19922);
or UO_298 (O_298,N_19901,N_19852);
nor UO_299 (O_299,N_19917,N_19965);
nand UO_300 (O_300,N_19900,N_19816);
or UO_301 (O_301,N_19969,N_19884);
nor UO_302 (O_302,N_19830,N_19973);
or UO_303 (O_303,N_19884,N_19926);
nand UO_304 (O_304,N_19820,N_19987);
xnor UO_305 (O_305,N_19878,N_19928);
xor UO_306 (O_306,N_19964,N_19881);
xnor UO_307 (O_307,N_19965,N_19933);
nand UO_308 (O_308,N_19981,N_19925);
nor UO_309 (O_309,N_19809,N_19917);
xnor UO_310 (O_310,N_19839,N_19855);
xnor UO_311 (O_311,N_19874,N_19933);
nor UO_312 (O_312,N_19927,N_19994);
nand UO_313 (O_313,N_19821,N_19833);
and UO_314 (O_314,N_19844,N_19811);
or UO_315 (O_315,N_19886,N_19915);
xnor UO_316 (O_316,N_19800,N_19922);
or UO_317 (O_317,N_19832,N_19997);
and UO_318 (O_318,N_19973,N_19913);
xnor UO_319 (O_319,N_19989,N_19978);
xor UO_320 (O_320,N_19903,N_19835);
xor UO_321 (O_321,N_19848,N_19849);
nor UO_322 (O_322,N_19879,N_19930);
or UO_323 (O_323,N_19933,N_19864);
or UO_324 (O_324,N_19940,N_19883);
and UO_325 (O_325,N_19871,N_19842);
nor UO_326 (O_326,N_19988,N_19807);
and UO_327 (O_327,N_19831,N_19842);
and UO_328 (O_328,N_19825,N_19861);
or UO_329 (O_329,N_19886,N_19947);
xnor UO_330 (O_330,N_19940,N_19969);
nor UO_331 (O_331,N_19936,N_19997);
and UO_332 (O_332,N_19833,N_19969);
nor UO_333 (O_333,N_19823,N_19859);
nor UO_334 (O_334,N_19802,N_19987);
and UO_335 (O_335,N_19859,N_19828);
or UO_336 (O_336,N_19963,N_19890);
and UO_337 (O_337,N_19954,N_19910);
nand UO_338 (O_338,N_19852,N_19924);
nand UO_339 (O_339,N_19966,N_19997);
or UO_340 (O_340,N_19927,N_19989);
or UO_341 (O_341,N_19834,N_19832);
and UO_342 (O_342,N_19980,N_19919);
or UO_343 (O_343,N_19894,N_19820);
nor UO_344 (O_344,N_19940,N_19979);
or UO_345 (O_345,N_19888,N_19917);
or UO_346 (O_346,N_19958,N_19929);
xor UO_347 (O_347,N_19960,N_19867);
or UO_348 (O_348,N_19924,N_19988);
xnor UO_349 (O_349,N_19887,N_19897);
xor UO_350 (O_350,N_19831,N_19941);
nand UO_351 (O_351,N_19935,N_19941);
xor UO_352 (O_352,N_19865,N_19895);
or UO_353 (O_353,N_19901,N_19846);
xnor UO_354 (O_354,N_19943,N_19999);
and UO_355 (O_355,N_19895,N_19958);
nand UO_356 (O_356,N_19834,N_19948);
nand UO_357 (O_357,N_19895,N_19845);
or UO_358 (O_358,N_19818,N_19840);
xnor UO_359 (O_359,N_19890,N_19875);
nand UO_360 (O_360,N_19917,N_19846);
nor UO_361 (O_361,N_19839,N_19849);
or UO_362 (O_362,N_19939,N_19922);
and UO_363 (O_363,N_19986,N_19856);
and UO_364 (O_364,N_19826,N_19985);
nor UO_365 (O_365,N_19910,N_19856);
and UO_366 (O_366,N_19957,N_19847);
and UO_367 (O_367,N_19866,N_19938);
xor UO_368 (O_368,N_19862,N_19972);
and UO_369 (O_369,N_19972,N_19969);
and UO_370 (O_370,N_19854,N_19817);
nand UO_371 (O_371,N_19831,N_19895);
nor UO_372 (O_372,N_19932,N_19812);
nor UO_373 (O_373,N_19883,N_19965);
nand UO_374 (O_374,N_19818,N_19892);
or UO_375 (O_375,N_19986,N_19929);
and UO_376 (O_376,N_19873,N_19903);
or UO_377 (O_377,N_19870,N_19897);
nand UO_378 (O_378,N_19911,N_19907);
nor UO_379 (O_379,N_19980,N_19883);
nand UO_380 (O_380,N_19840,N_19961);
and UO_381 (O_381,N_19950,N_19986);
and UO_382 (O_382,N_19850,N_19832);
and UO_383 (O_383,N_19897,N_19923);
nor UO_384 (O_384,N_19959,N_19962);
and UO_385 (O_385,N_19903,N_19840);
and UO_386 (O_386,N_19912,N_19808);
or UO_387 (O_387,N_19973,N_19901);
or UO_388 (O_388,N_19897,N_19978);
nand UO_389 (O_389,N_19921,N_19930);
xor UO_390 (O_390,N_19919,N_19873);
xnor UO_391 (O_391,N_19847,N_19949);
nand UO_392 (O_392,N_19873,N_19834);
xnor UO_393 (O_393,N_19860,N_19903);
xor UO_394 (O_394,N_19976,N_19991);
nand UO_395 (O_395,N_19863,N_19948);
and UO_396 (O_396,N_19868,N_19882);
xor UO_397 (O_397,N_19896,N_19994);
or UO_398 (O_398,N_19869,N_19832);
xor UO_399 (O_399,N_19858,N_19800);
or UO_400 (O_400,N_19818,N_19950);
nand UO_401 (O_401,N_19887,N_19855);
nand UO_402 (O_402,N_19959,N_19856);
and UO_403 (O_403,N_19908,N_19961);
and UO_404 (O_404,N_19918,N_19910);
or UO_405 (O_405,N_19829,N_19866);
xnor UO_406 (O_406,N_19912,N_19898);
and UO_407 (O_407,N_19981,N_19889);
or UO_408 (O_408,N_19808,N_19975);
xor UO_409 (O_409,N_19820,N_19862);
nand UO_410 (O_410,N_19801,N_19981);
nor UO_411 (O_411,N_19935,N_19836);
nand UO_412 (O_412,N_19940,N_19801);
xor UO_413 (O_413,N_19974,N_19959);
nor UO_414 (O_414,N_19972,N_19976);
and UO_415 (O_415,N_19875,N_19840);
xor UO_416 (O_416,N_19840,N_19886);
nor UO_417 (O_417,N_19848,N_19836);
nand UO_418 (O_418,N_19976,N_19955);
nand UO_419 (O_419,N_19988,N_19973);
nor UO_420 (O_420,N_19826,N_19997);
nand UO_421 (O_421,N_19940,N_19956);
nand UO_422 (O_422,N_19980,N_19857);
nor UO_423 (O_423,N_19949,N_19801);
xor UO_424 (O_424,N_19850,N_19802);
nand UO_425 (O_425,N_19851,N_19817);
nand UO_426 (O_426,N_19985,N_19912);
nor UO_427 (O_427,N_19922,N_19825);
nor UO_428 (O_428,N_19896,N_19856);
and UO_429 (O_429,N_19892,N_19857);
xor UO_430 (O_430,N_19958,N_19928);
or UO_431 (O_431,N_19832,N_19985);
xor UO_432 (O_432,N_19861,N_19904);
and UO_433 (O_433,N_19841,N_19802);
or UO_434 (O_434,N_19987,N_19876);
nand UO_435 (O_435,N_19910,N_19919);
xnor UO_436 (O_436,N_19905,N_19855);
and UO_437 (O_437,N_19832,N_19948);
nand UO_438 (O_438,N_19968,N_19961);
and UO_439 (O_439,N_19851,N_19976);
xnor UO_440 (O_440,N_19956,N_19840);
or UO_441 (O_441,N_19800,N_19803);
and UO_442 (O_442,N_19966,N_19845);
and UO_443 (O_443,N_19866,N_19876);
or UO_444 (O_444,N_19955,N_19893);
xnor UO_445 (O_445,N_19844,N_19903);
nand UO_446 (O_446,N_19964,N_19809);
nand UO_447 (O_447,N_19970,N_19830);
or UO_448 (O_448,N_19913,N_19979);
and UO_449 (O_449,N_19836,N_19899);
nor UO_450 (O_450,N_19911,N_19853);
or UO_451 (O_451,N_19913,N_19942);
xnor UO_452 (O_452,N_19926,N_19998);
xnor UO_453 (O_453,N_19833,N_19981);
nand UO_454 (O_454,N_19882,N_19928);
and UO_455 (O_455,N_19975,N_19828);
or UO_456 (O_456,N_19988,N_19835);
xnor UO_457 (O_457,N_19836,N_19852);
xor UO_458 (O_458,N_19969,N_19958);
nand UO_459 (O_459,N_19862,N_19995);
xor UO_460 (O_460,N_19950,N_19991);
and UO_461 (O_461,N_19978,N_19914);
nor UO_462 (O_462,N_19878,N_19990);
nor UO_463 (O_463,N_19906,N_19921);
or UO_464 (O_464,N_19881,N_19836);
and UO_465 (O_465,N_19859,N_19991);
nand UO_466 (O_466,N_19811,N_19816);
or UO_467 (O_467,N_19894,N_19978);
nor UO_468 (O_468,N_19955,N_19989);
and UO_469 (O_469,N_19914,N_19838);
nor UO_470 (O_470,N_19944,N_19891);
or UO_471 (O_471,N_19873,N_19869);
and UO_472 (O_472,N_19854,N_19901);
or UO_473 (O_473,N_19801,N_19865);
or UO_474 (O_474,N_19855,N_19950);
or UO_475 (O_475,N_19812,N_19847);
nor UO_476 (O_476,N_19962,N_19828);
xnor UO_477 (O_477,N_19945,N_19901);
nor UO_478 (O_478,N_19864,N_19914);
xor UO_479 (O_479,N_19908,N_19888);
xor UO_480 (O_480,N_19967,N_19970);
or UO_481 (O_481,N_19916,N_19857);
or UO_482 (O_482,N_19901,N_19979);
nand UO_483 (O_483,N_19913,N_19907);
and UO_484 (O_484,N_19933,N_19865);
xor UO_485 (O_485,N_19909,N_19889);
nor UO_486 (O_486,N_19835,N_19843);
and UO_487 (O_487,N_19916,N_19973);
or UO_488 (O_488,N_19962,N_19941);
or UO_489 (O_489,N_19852,N_19838);
nor UO_490 (O_490,N_19823,N_19990);
nor UO_491 (O_491,N_19930,N_19904);
or UO_492 (O_492,N_19831,N_19918);
nor UO_493 (O_493,N_19982,N_19912);
nor UO_494 (O_494,N_19875,N_19895);
nand UO_495 (O_495,N_19996,N_19968);
and UO_496 (O_496,N_19961,N_19913);
xor UO_497 (O_497,N_19875,N_19947);
and UO_498 (O_498,N_19874,N_19924);
and UO_499 (O_499,N_19945,N_19855);
or UO_500 (O_500,N_19883,N_19929);
and UO_501 (O_501,N_19946,N_19967);
xor UO_502 (O_502,N_19815,N_19857);
and UO_503 (O_503,N_19921,N_19831);
and UO_504 (O_504,N_19991,N_19966);
nand UO_505 (O_505,N_19853,N_19841);
xor UO_506 (O_506,N_19808,N_19858);
nand UO_507 (O_507,N_19993,N_19859);
nand UO_508 (O_508,N_19887,N_19822);
nand UO_509 (O_509,N_19870,N_19985);
xor UO_510 (O_510,N_19944,N_19975);
xnor UO_511 (O_511,N_19932,N_19836);
xnor UO_512 (O_512,N_19936,N_19993);
and UO_513 (O_513,N_19995,N_19953);
nor UO_514 (O_514,N_19990,N_19988);
nand UO_515 (O_515,N_19995,N_19982);
xor UO_516 (O_516,N_19813,N_19980);
or UO_517 (O_517,N_19843,N_19850);
or UO_518 (O_518,N_19866,N_19816);
xor UO_519 (O_519,N_19872,N_19930);
nand UO_520 (O_520,N_19909,N_19874);
and UO_521 (O_521,N_19988,N_19849);
xor UO_522 (O_522,N_19958,N_19880);
or UO_523 (O_523,N_19873,N_19882);
xor UO_524 (O_524,N_19986,N_19988);
nand UO_525 (O_525,N_19920,N_19830);
xnor UO_526 (O_526,N_19923,N_19873);
xor UO_527 (O_527,N_19904,N_19860);
nand UO_528 (O_528,N_19868,N_19803);
and UO_529 (O_529,N_19878,N_19957);
xnor UO_530 (O_530,N_19838,N_19971);
nor UO_531 (O_531,N_19955,N_19977);
xnor UO_532 (O_532,N_19998,N_19815);
or UO_533 (O_533,N_19924,N_19808);
xor UO_534 (O_534,N_19906,N_19944);
xor UO_535 (O_535,N_19839,N_19831);
or UO_536 (O_536,N_19973,N_19908);
nand UO_537 (O_537,N_19999,N_19843);
xor UO_538 (O_538,N_19836,N_19802);
nor UO_539 (O_539,N_19870,N_19929);
xnor UO_540 (O_540,N_19871,N_19950);
nand UO_541 (O_541,N_19895,N_19826);
nor UO_542 (O_542,N_19818,N_19959);
or UO_543 (O_543,N_19822,N_19950);
xor UO_544 (O_544,N_19804,N_19883);
and UO_545 (O_545,N_19931,N_19849);
and UO_546 (O_546,N_19888,N_19913);
or UO_547 (O_547,N_19886,N_19890);
and UO_548 (O_548,N_19845,N_19889);
and UO_549 (O_549,N_19945,N_19888);
xnor UO_550 (O_550,N_19938,N_19853);
nand UO_551 (O_551,N_19830,N_19954);
nand UO_552 (O_552,N_19905,N_19822);
nand UO_553 (O_553,N_19824,N_19935);
or UO_554 (O_554,N_19922,N_19865);
xor UO_555 (O_555,N_19897,N_19899);
and UO_556 (O_556,N_19857,N_19965);
xor UO_557 (O_557,N_19981,N_19934);
nor UO_558 (O_558,N_19960,N_19964);
nor UO_559 (O_559,N_19998,N_19878);
nand UO_560 (O_560,N_19923,N_19854);
nor UO_561 (O_561,N_19940,N_19978);
or UO_562 (O_562,N_19951,N_19927);
nand UO_563 (O_563,N_19975,N_19856);
and UO_564 (O_564,N_19871,N_19971);
xor UO_565 (O_565,N_19861,N_19938);
xnor UO_566 (O_566,N_19874,N_19905);
nand UO_567 (O_567,N_19950,N_19923);
and UO_568 (O_568,N_19984,N_19967);
nor UO_569 (O_569,N_19961,N_19878);
nor UO_570 (O_570,N_19962,N_19815);
xor UO_571 (O_571,N_19952,N_19911);
xor UO_572 (O_572,N_19820,N_19907);
or UO_573 (O_573,N_19800,N_19912);
and UO_574 (O_574,N_19928,N_19997);
and UO_575 (O_575,N_19992,N_19903);
and UO_576 (O_576,N_19953,N_19840);
nor UO_577 (O_577,N_19980,N_19990);
and UO_578 (O_578,N_19871,N_19935);
or UO_579 (O_579,N_19898,N_19870);
nor UO_580 (O_580,N_19893,N_19841);
xor UO_581 (O_581,N_19942,N_19992);
xnor UO_582 (O_582,N_19849,N_19999);
nand UO_583 (O_583,N_19926,N_19948);
or UO_584 (O_584,N_19850,N_19955);
and UO_585 (O_585,N_19840,N_19998);
xor UO_586 (O_586,N_19950,N_19840);
or UO_587 (O_587,N_19975,N_19839);
nor UO_588 (O_588,N_19889,N_19839);
xor UO_589 (O_589,N_19840,N_19958);
and UO_590 (O_590,N_19968,N_19984);
nor UO_591 (O_591,N_19853,N_19950);
xnor UO_592 (O_592,N_19968,N_19833);
nor UO_593 (O_593,N_19878,N_19893);
and UO_594 (O_594,N_19841,N_19995);
nor UO_595 (O_595,N_19924,N_19944);
nor UO_596 (O_596,N_19892,N_19901);
and UO_597 (O_597,N_19935,N_19873);
or UO_598 (O_598,N_19900,N_19948);
nand UO_599 (O_599,N_19807,N_19904);
or UO_600 (O_600,N_19802,N_19832);
and UO_601 (O_601,N_19878,N_19987);
nor UO_602 (O_602,N_19828,N_19936);
nand UO_603 (O_603,N_19840,N_19879);
or UO_604 (O_604,N_19874,N_19937);
or UO_605 (O_605,N_19835,N_19838);
xnor UO_606 (O_606,N_19870,N_19835);
nand UO_607 (O_607,N_19922,N_19897);
nor UO_608 (O_608,N_19880,N_19948);
nand UO_609 (O_609,N_19897,N_19824);
xnor UO_610 (O_610,N_19869,N_19885);
and UO_611 (O_611,N_19882,N_19893);
nand UO_612 (O_612,N_19942,N_19879);
or UO_613 (O_613,N_19994,N_19835);
and UO_614 (O_614,N_19896,N_19919);
xor UO_615 (O_615,N_19938,N_19946);
nand UO_616 (O_616,N_19816,N_19977);
nor UO_617 (O_617,N_19995,N_19880);
or UO_618 (O_618,N_19890,N_19919);
nor UO_619 (O_619,N_19896,N_19971);
nand UO_620 (O_620,N_19867,N_19800);
and UO_621 (O_621,N_19807,N_19903);
xnor UO_622 (O_622,N_19869,N_19941);
or UO_623 (O_623,N_19953,N_19961);
and UO_624 (O_624,N_19822,N_19974);
or UO_625 (O_625,N_19940,N_19997);
and UO_626 (O_626,N_19901,N_19870);
xor UO_627 (O_627,N_19999,N_19887);
and UO_628 (O_628,N_19881,N_19833);
xnor UO_629 (O_629,N_19863,N_19824);
nor UO_630 (O_630,N_19980,N_19978);
and UO_631 (O_631,N_19925,N_19973);
and UO_632 (O_632,N_19958,N_19937);
nand UO_633 (O_633,N_19965,N_19943);
xor UO_634 (O_634,N_19914,N_19873);
nand UO_635 (O_635,N_19998,N_19964);
nor UO_636 (O_636,N_19974,N_19859);
xnor UO_637 (O_637,N_19825,N_19969);
nor UO_638 (O_638,N_19965,N_19867);
nor UO_639 (O_639,N_19914,N_19955);
nand UO_640 (O_640,N_19893,N_19935);
xnor UO_641 (O_641,N_19980,N_19817);
xnor UO_642 (O_642,N_19969,N_19815);
nor UO_643 (O_643,N_19828,N_19845);
xnor UO_644 (O_644,N_19996,N_19924);
nor UO_645 (O_645,N_19971,N_19928);
or UO_646 (O_646,N_19890,N_19834);
nand UO_647 (O_647,N_19948,N_19969);
and UO_648 (O_648,N_19944,N_19895);
xor UO_649 (O_649,N_19949,N_19992);
and UO_650 (O_650,N_19968,N_19821);
and UO_651 (O_651,N_19826,N_19883);
and UO_652 (O_652,N_19874,N_19830);
or UO_653 (O_653,N_19867,N_19877);
or UO_654 (O_654,N_19896,N_19920);
and UO_655 (O_655,N_19911,N_19897);
xor UO_656 (O_656,N_19973,N_19883);
and UO_657 (O_657,N_19909,N_19985);
xor UO_658 (O_658,N_19851,N_19821);
xnor UO_659 (O_659,N_19980,N_19885);
nand UO_660 (O_660,N_19895,N_19938);
xor UO_661 (O_661,N_19930,N_19949);
and UO_662 (O_662,N_19992,N_19982);
xnor UO_663 (O_663,N_19911,N_19857);
xor UO_664 (O_664,N_19854,N_19867);
nor UO_665 (O_665,N_19962,N_19834);
nor UO_666 (O_666,N_19829,N_19828);
and UO_667 (O_667,N_19985,N_19895);
nor UO_668 (O_668,N_19881,N_19902);
nand UO_669 (O_669,N_19832,N_19868);
xnor UO_670 (O_670,N_19899,N_19952);
xnor UO_671 (O_671,N_19810,N_19852);
xnor UO_672 (O_672,N_19980,N_19976);
nor UO_673 (O_673,N_19998,N_19880);
and UO_674 (O_674,N_19938,N_19837);
and UO_675 (O_675,N_19889,N_19902);
nor UO_676 (O_676,N_19837,N_19863);
xnor UO_677 (O_677,N_19869,N_19904);
or UO_678 (O_678,N_19881,N_19863);
and UO_679 (O_679,N_19861,N_19947);
xor UO_680 (O_680,N_19869,N_19977);
nor UO_681 (O_681,N_19888,N_19942);
nand UO_682 (O_682,N_19820,N_19823);
and UO_683 (O_683,N_19868,N_19883);
or UO_684 (O_684,N_19845,N_19926);
nand UO_685 (O_685,N_19915,N_19973);
nand UO_686 (O_686,N_19981,N_19996);
and UO_687 (O_687,N_19868,N_19805);
xor UO_688 (O_688,N_19952,N_19978);
nand UO_689 (O_689,N_19812,N_19964);
nor UO_690 (O_690,N_19885,N_19958);
or UO_691 (O_691,N_19800,N_19877);
and UO_692 (O_692,N_19941,N_19913);
nand UO_693 (O_693,N_19866,N_19963);
and UO_694 (O_694,N_19999,N_19857);
and UO_695 (O_695,N_19923,N_19869);
and UO_696 (O_696,N_19918,N_19903);
nand UO_697 (O_697,N_19915,N_19853);
and UO_698 (O_698,N_19911,N_19889);
or UO_699 (O_699,N_19922,N_19951);
and UO_700 (O_700,N_19842,N_19895);
or UO_701 (O_701,N_19804,N_19893);
nand UO_702 (O_702,N_19854,N_19992);
xnor UO_703 (O_703,N_19822,N_19877);
or UO_704 (O_704,N_19813,N_19898);
nor UO_705 (O_705,N_19908,N_19801);
and UO_706 (O_706,N_19825,N_19801);
nand UO_707 (O_707,N_19812,N_19864);
xor UO_708 (O_708,N_19986,N_19857);
or UO_709 (O_709,N_19832,N_19933);
nand UO_710 (O_710,N_19991,N_19887);
or UO_711 (O_711,N_19911,N_19835);
nand UO_712 (O_712,N_19859,N_19807);
nand UO_713 (O_713,N_19815,N_19981);
or UO_714 (O_714,N_19948,N_19840);
or UO_715 (O_715,N_19888,N_19941);
xor UO_716 (O_716,N_19920,N_19966);
or UO_717 (O_717,N_19907,N_19965);
and UO_718 (O_718,N_19864,N_19897);
nor UO_719 (O_719,N_19804,N_19838);
xor UO_720 (O_720,N_19907,N_19866);
or UO_721 (O_721,N_19994,N_19824);
or UO_722 (O_722,N_19811,N_19868);
and UO_723 (O_723,N_19942,N_19961);
or UO_724 (O_724,N_19889,N_19973);
and UO_725 (O_725,N_19821,N_19801);
or UO_726 (O_726,N_19849,N_19857);
nand UO_727 (O_727,N_19802,N_19914);
nand UO_728 (O_728,N_19956,N_19854);
nor UO_729 (O_729,N_19812,N_19933);
nor UO_730 (O_730,N_19964,N_19832);
or UO_731 (O_731,N_19904,N_19821);
nand UO_732 (O_732,N_19977,N_19934);
xnor UO_733 (O_733,N_19941,N_19915);
or UO_734 (O_734,N_19877,N_19883);
or UO_735 (O_735,N_19983,N_19993);
xnor UO_736 (O_736,N_19930,N_19824);
xnor UO_737 (O_737,N_19952,N_19832);
xnor UO_738 (O_738,N_19802,N_19986);
nand UO_739 (O_739,N_19800,N_19935);
nand UO_740 (O_740,N_19828,N_19822);
nand UO_741 (O_741,N_19880,N_19926);
or UO_742 (O_742,N_19816,N_19936);
or UO_743 (O_743,N_19896,N_19959);
and UO_744 (O_744,N_19802,N_19993);
xnor UO_745 (O_745,N_19849,N_19846);
or UO_746 (O_746,N_19867,N_19971);
nand UO_747 (O_747,N_19902,N_19822);
and UO_748 (O_748,N_19993,N_19894);
or UO_749 (O_749,N_19860,N_19995);
nor UO_750 (O_750,N_19826,N_19892);
or UO_751 (O_751,N_19944,N_19836);
and UO_752 (O_752,N_19855,N_19814);
xor UO_753 (O_753,N_19875,N_19901);
nand UO_754 (O_754,N_19862,N_19913);
and UO_755 (O_755,N_19892,N_19823);
or UO_756 (O_756,N_19937,N_19986);
and UO_757 (O_757,N_19826,N_19960);
or UO_758 (O_758,N_19802,N_19882);
and UO_759 (O_759,N_19985,N_19851);
nand UO_760 (O_760,N_19999,N_19939);
nand UO_761 (O_761,N_19927,N_19950);
xnor UO_762 (O_762,N_19856,N_19980);
nand UO_763 (O_763,N_19906,N_19911);
nand UO_764 (O_764,N_19998,N_19811);
xnor UO_765 (O_765,N_19838,N_19841);
and UO_766 (O_766,N_19892,N_19904);
and UO_767 (O_767,N_19920,N_19867);
and UO_768 (O_768,N_19824,N_19878);
or UO_769 (O_769,N_19857,N_19949);
and UO_770 (O_770,N_19863,N_19977);
or UO_771 (O_771,N_19875,N_19808);
or UO_772 (O_772,N_19889,N_19991);
or UO_773 (O_773,N_19973,N_19943);
and UO_774 (O_774,N_19967,N_19877);
nand UO_775 (O_775,N_19950,N_19806);
nand UO_776 (O_776,N_19961,N_19991);
nor UO_777 (O_777,N_19959,N_19879);
nor UO_778 (O_778,N_19875,N_19907);
nand UO_779 (O_779,N_19827,N_19931);
and UO_780 (O_780,N_19930,N_19896);
or UO_781 (O_781,N_19915,N_19807);
xor UO_782 (O_782,N_19838,N_19810);
nor UO_783 (O_783,N_19891,N_19883);
and UO_784 (O_784,N_19959,N_19840);
and UO_785 (O_785,N_19885,N_19985);
or UO_786 (O_786,N_19975,N_19810);
xor UO_787 (O_787,N_19934,N_19970);
and UO_788 (O_788,N_19942,N_19962);
or UO_789 (O_789,N_19912,N_19960);
and UO_790 (O_790,N_19841,N_19913);
or UO_791 (O_791,N_19860,N_19934);
and UO_792 (O_792,N_19922,N_19905);
or UO_793 (O_793,N_19812,N_19983);
or UO_794 (O_794,N_19814,N_19963);
nand UO_795 (O_795,N_19820,N_19900);
and UO_796 (O_796,N_19994,N_19953);
nand UO_797 (O_797,N_19936,N_19896);
nand UO_798 (O_798,N_19883,N_19854);
or UO_799 (O_799,N_19991,N_19874);
xor UO_800 (O_800,N_19841,N_19912);
or UO_801 (O_801,N_19942,N_19989);
or UO_802 (O_802,N_19865,N_19910);
xor UO_803 (O_803,N_19951,N_19936);
xnor UO_804 (O_804,N_19968,N_19963);
nand UO_805 (O_805,N_19983,N_19887);
or UO_806 (O_806,N_19957,N_19914);
nor UO_807 (O_807,N_19841,N_19946);
or UO_808 (O_808,N_19884,N_19911);
or UO_809 (O_809,N_19893,N_19900);
and UO_810 (O_810,N_19927,N_19843);
nand UO_811 (O_811,N_19879,N_19841);
xnor UO_812 (O_812,N_19933,N_19908);
nand UO_813 (O_813,N_19954,N_19865);
or UO_814 (O_814,N_19979,N_19934);
nand UO_815 (O_815,N_19856,N_19934);
nor UO_816 (O_816,N_19805,N_19812);
and UO_817 (O_817,N_19806,N_19998);
or UO_818 (O_818,N_19885,N_19875);
and UO_819 (O_819,N_19949,N_19975);
and UO_820 (O_820,N_19822,N_19817);
nor UO_821 (O_821,N_19946,N_19922);
nand UO_822 (O_822,N_19990,N_19813);
xnor UO_823 (O_823,N_19856,N_19842);
xor UO_824 (O_824,N_19982,N_19844);
or UO_825 (O_825,N_19900,N_19901);
nor UO_826 (O_826,N_19808,N_19882);
nor UO_827 (O_827,N_19818,N_19943);
nor UO_828 (O_828,N_19897,N_19985);
nand UO_829 (O_829,N_19907,N_19958);
nor UO_830 (O_830,N_19823,N_19952);
nor UO_831 (O_831,N_19987,N_19935);
and UO_832 (O_832,N_19813,N_19880);
and UO_833 (O_833,N_19878,N_19803);
nor UO_834 (O_834,N_19899,N_19926);
and UO_835 (O_835,N_19914,N_19924);
nand UO_836 (O_836,N_19981,N_19961);
and UO_837 (O_837,N_19968,N_19847);
nor UO_838 (O_838,N_19868,N_19890);
xnor UO_839 (O_839,N_19965,N_19906);
xor UO_840 (O_840,N_19959,N_19892);
nor UO_841 (O_841,N_19827,N_19825);
nor UO_842 (O_842,N_19831,N_19853);
or UO_843 (O_843,N_19987,N_19947);
xor UO_844 (O_844,N_19911,N_19898);
nor UO_845 (O_845,N_19811,N_19884);
xor UO_846 (O_846,N_19903,N_19936);
nand UO_847 (O_847,N_19841,N_19804);
nor UO_848 (O_848,N_19874,N_19949);
or UO_849 (O_849,N_19993,N_19851);
or UO_850 (O_850,N_19900,N_19831);
nand UO_851 (O_851,N_19901,N_19868);
or UO_852 (O_852,N_19816,N_19864);
or UO_853 (O_853,N_19906,N_19892);
xnor UO_854 (O_854,N_19971,N_19863);
xnor UO_855 (O_855,N_19944,N_19989);
nand UO_856 (O_856,N_19999,N_19908);
nand UO_857 (O_857,N_19807,N_19870);
nor UO_858 (O_858,N_19960,N_19954);
and UO_859 (O_859,N_19999,N_19888);
or UO_860 (O_860,N_19973,N_19979);
xnor UO_861 (O_861,N_19981,N_19860);
xor UO_862 (O_862,N_19932,N_19813);
nor UO_863 (O_863,N_19880,N_19909);
nor UO_864 (O_864,N_19838,N_19953);
or UO_865 (O_865,N_19961,N_19915);
and UO_866 (O_866,N_19805,N_19802);
xnor UO_867 (O_867,N_19926,N_19894);
nand UO_868 (O_868,N_19964,N_19892);
nand UO_869 (O_869,N_19856,N_19826);
and UO_870 (O_870,N_19841,N_19989);
or UO_871 (O_871,N_19871,N_19850);
nand UO_872 (O_872,N_19915,N_19873);
and UO_873 (O_873,N_19866,N_19832);
nor UO_874 (O_874,N_19827,N_19970);
nand UO_875 (O_875,N_19931,N_19976);
or UO_876 (O_876,N_19821,N_19934);
nand UO_877 (O_877,N_19978,N_19811);
nand UO_878 (O_878,N_19982,N_19868);
or UO_879 (O_879,N_19891,N_19945);
nor UO_880 (O_880,N_19930,N_19861);
or UO_881 (O_881,N_19905,N_19830);
xnor UO_882 (O_882,N_19993,N_19881);
nand UO_883 (O_883,N_19959,N_19825);
or UO_884 (O_884,N_19801,N_19997);
nand UO_885 (O_885,N_19910,N_19925);
xor UO_886 (O_886,N_19900,N_19993);
xnor UO_887 (O_887,N_19933,N_19915);
or UO_888 (O_888,N_19963,N_19856);
nand UO_889 (O_889,N_19809,N_19968);
nand UO_890 (O_890,N_19815,N_19864);
xnor UO_891 (O_891,N_19846,N_19985);
nand UO_892 (O_892,N_19817,N_19929);
nand UO_893 (O_893,N_19861,N_19983);
and UO_894 (O_894,N_19910,N_19860);
nand UO_895 (O_895,N_19868,N_19939);
xor UO_896 (O_896,N_19898,N_19985);
nand UO_897 (O_897,N_19958,N_19883);
or UO_898 (O_898,N_19801,N_19986);
or UO_899 (O_899,N_19961,N_19929);
and UO_900 (O_900,N_19889,N_19868);
nor UO_901 (O_901,N_19802,N_19899);
xnor UO_902 (O_902,N_19950,N_19942);
nor UO_903 (O_903,N_19907,N_19800);
xor UO_904 (O_904,N_19861,N_19844);
nand UO_905 (O_905,N_19908,N_19930);
and UO_906 (O_906,N_19904,N_19983);
nand UO_907 (O_907,N_19981,N_19986);
or UO_908 (O_908,N_19803,N_19889);
xnor UO_909 (O_909,N_19910,N_19834);
or UO_910 (O_910,N_19868,N_19955);
xnor UO_911 (O_911,N_19828,N_19985);
xor UO_912 (O_912,N_19943,N_19956);
and UO_913 (O_913,N_19844,N_19847);
and UO_914 (O_914,N_19888,N_19903);
and UO_915 (O_915,N_19997,N_19915);
or UO_916 (O_916,N_19974,N_19826);
nand UO_917 (O_917,N_19880,N_19855);
nor UO_918 (O_918,N_19821,N_19953);
nor UO_919 (O_919,N_19968,N_19839);
or UO_920 (O_920,N_19956,N_19845);
or UO_921 (O_921,N_19867,N_19813);
xor UO_922 (O_922,N_19842,N_19884);
and UO_923 (O_923,N_19803,N_19992);
nand UO_924 (O_924,N_19991,N_19984);
and UO_925 (O_925,N_19977,N_19896);
nor UO_926 (O_926,N_19960,N_19952);
nand UO_927 (O_927,N_19944,N_19870);
nand UO_928 (O_928,N_19949,N_19966);
and UO_929 (O_929,N_19866,N_19980);
xor UO_930 (O_930,N_19874,N_19930);
xor UO_931 (O_931,N_19832,N_19940);
nand UO_932 (O_932,N_19925,N_19808);
and UO_933 (O_933,N_19925,N_19842);
or UO_934 (O_934,N_19950,N_19947);
nand UO_935 (O_935,N_19977,N_19810);
and UO_936 (O_936,N_19961,N_19902);
or UO_937 (O_937,N_19842,N_19829);
and UO_938 (O_938,N_19882,N_19914);
and UO_939 (O_939,N_19902,N_19897);
nor UO_940 (O_940,N_19932,N_19933);
nor UO_941 (O_941,N_19892,N_19858);
and UO_942 (O_942,N_19959,N_19999);
nor UO_943 (O_943,N_19956,N_19869);
and UO_944 (O_944,N_19982,N_19969);
or UO_945 (O_945,N_19873,N_19927);
nand UO_946 (O_946,N_19889,N_19828);
and UO_947 (O_947,N_19982,N_19879);
xnor UO_948 (O_948,N_19926,N_19865);
and UO_949 (O_949,N_19904,N_19876);
nor UO_950 (O_950,N_19853,N_19852);
and UO_951 (O_951,N_19987,N_19845);
xor UO_952 (O_952,N_19820,N_19940);
and UO_953 (O_953,N_19895,N_19809);
xnor UO_954 (O_954,N_19917,N_19830);
xnor UO_955 (O_955,N_19815,N_19881);
xnor UO_956 (O_956,N_19890,N_19909);
or UO_957 (O_957,N_19812,N_19966);
and UO_958 (O_958,N_19822,N_19967);
nor UO_959 (O_959,N_19855,N_19828);
nand UO_960 (O_960,N_19918,N_19866);
nor UO_961 (O_961,N_19908,N_19880);
xor UO_962 (O_962,N_19882,N_19896);
and UO_963 (O_963,N_19838,N_19830);
nand UO_964 (O_964,N_19986,N_19926);
nand UO_965 (O_965,N_19866,N_19884);
nand UO_966 (O_966,N_19966,N_19884);
nor UO_967 (O_967,N_19848,N_19806);
or UO_968 (O_968,N_19824,N_19940);
or UO_969 (O_969,N_19885,N_19864);
nand UO_970 (O_970,N_19989,N_19958);
xnor UO_971 (O_971,N_19868,N_19814);
or UO_972 (O_972,N_19820,N_19919);
nand UO_973 (O_973,N_19833,N_19992);
nand UO_974 (O_974,N_19871,N_19800);
xnor UO_975 (O_975,N_19943,N_19819);
nand UO_976 (O_976,N_19985,N_19841);
nor UO_977 (O_977,N_19845,N_19811);
and UO_978 (O_978,N_19976,N_19850);
or UO_979 (O_979,N_19839,N_19914);
and UO_980 (O_980,N_19849,N_19881);
and UO_981 (O_981,N_19937,N_19982);
xnor UO_982 (O_982,N_19969,N_19883);
or UO_983 (O_983,N_19947,N_19984);
and UO_984 (O_984,N_19803,N_19902);
xnor UO_985 (O_985,N_19876,N_19882);
xnor UO_986 (O_986,N_19862,N_19865);
nor UO_987 (O_987,N_19836,N_19957);
or UO_988 (O_988,N_19835,N_19883);
nor UO_989 (O_989,N_19946,N_19890);
or UO_990 (O_990,N_19932,N_19930);
nor UO_991 (O_991,N_19847,N_19958);
nor UO_992 (O_992,N_19913,N_19910);
nand UO_993 (O_993,N_19839,N_19990);
and UO_994 (O_994,N_19870,N_19818);
or UO_995 (O_995,N_19907,N_19871);
nor UO_996 (O_996,N_19837,N_19965);
or UO_997 (O_997,N_19947,N_19819);
or UO_998 (O_998,N_19889,N_19950);
nor UO_999 (O_999,N_19884,N_19977);
and UO_1000 (O_1000,N_19871,N_19985);
and UO_1001 (O_1001,N_19899,N_19938);
xor UO_1002 (O_1002,N_19860,N_19814);
xor UO_1003 (O_1003,N_19954,N_19979);
nand UO_1004 (O_1004,N_19814,N_19895);
xor UO_1005 (O_1005,N_19929,N_19853);
or UO_1006 (O_1006,N_19911,N_19816);
or UO_1007 (O_1007,N_19858,N_19824);
or UO_1008 (O_1008,N_19902,N_19875);
nand UO_1009 (O_1009,N_19860,N_19808);
and UO_1010 (O_1010,N_19805,N_19849);
nand UO_1011 (O_1011,N_19988,N_19808);
or UO_1012 (O_1012,N_19984,N_19918);
or UO_1013 (O_1013,N_19849,N_19887);
nand UO_1014 (O_1014,N_19828,N_19825);
nor UO_1015 (O_1015,N_19847,N_19803);
and UO_1016 (O_1016,N_19922,N_19958);
and UO_1017 (O_1017,N_19960,N_19893);
nor UO_1018 (O_1018,N_19932,N_19858);
nor UO_1019 (O_1019,N_19838,N_19906);
or UO_1020 (O_1020,N_19959,N_19991);
xor UO_1021 (O_1021,N_19820,N_19854);
xor UO_1022 (O_1022,N_19813,N_19841);
or UO_1023 (O_1023,N_19861,N_19884);
nand UO_1024 (O_1024,N_19836,N_19825);
xnor UO_1025 (O_1025,N_19862,N_19938);
xor UO_1026 (O_1026,N_19849,N_19868);
xor UO_1027 (O_1027,N_19965,N_19992);
nand UO_1028 (O_1028,N_19966,N_19967);
xor UO_1029 (O_1029,N_19919,N_19938);
nor UO_1030 (O_1030,N_19948,N_19952);
nand UO_1031 (O_1031,N_19881,N_19910);
and UO_1032 (O_1032,N_19964,N_19991);
nand UO_1033 (O_1033,N_19946,N_19882);
and UO_1034 (O_1034,N_19897,N_19973);
nand UO_1035 (O_1035,N_19814,N_19876);
nor UO_1036 (O_1036,N_19973,N_19946);
or UO_1037 (O_1037,N_19825,N_19933);
xnor UO_1038 (O_1038,N_19908,N_19953);
nor UO_1039 (O_1039,N_19921,N_19905);
nor UO_1040 (O_1040,N_19964,N_19827);
nand UO_1041 (O_1041,N_19843,N_19838);
xnor UO_1042 (O_1042,N_19831,N_19810);
and UO_1043 (O_1043,N_19927,N_19930);
or UO_1044 (O_1044,N_19806,N_19896);
or UO_1045 (O_1045,N_19814,N_19806);
or UO_1046 (O_1046,N_19970,N_19847);
and UO_1047 (O_1047,N_19800,N_19834);
xor UO_1048 (O_1048,N_19918,N_19897);
nor UO_1049 (O_1049,N_19872,N_19810);
and UO_1050 (O_1050,N_19929,N_19951);
nand UO_1051 (O_1051,N_19817,N_19911);
or UO_1052 (O_1052,N_19850,N_19901);
nor UO_1053 (O_1053,N_19872,N_19859);
or UO_1054 (O_1054,N_19944,N_19974);
or UO_1055 (O_1055,N_19855,N_19949);
nand UO_1056 (O_1056,N_19852,N_19982);
or UO_1057 (O_1057,N_19843,N_19858);
nand UO_1058 (O_1058,N_19894,N_19938);
xnor UO_1059 (O_1059,N_19828,N_19818);
nand UO_1060 (O_1060,N_19985,N_19966);
or UO_1061 (O_1061,N_19859,N_19868);
nor UO_1062 (O_1062,N_19886,N_19860);
nand UO_1063 (O_1063,N_19892,N_19982);
nand UO_1064 (O_1064,N_19918,N_19821);
nor UO_1065 (O_1065,N_19923,N_19911);
and UO_1066 (O_1066,N_19831,N_19992);
or UO_1067 (O_1067,N_19816,N_19809);
nand UO_1068 (O_1068,N_19930,N_19995);
xnor UO_1069 (O_1069,N_19929,N_19925);
xor UO_1070 (O_1070,N_19968,N_19943);
and UO_1071 (O_1071,N_19876,N_19965);
or UO_1072 (O_1072,N_19818,N_19946);
nor UO_1073 (O_1073,N_19912,N_19874);
and UO_1074 (O_1074,N_19967,N_19963);
nor UO_1075 (O_1075,N_19882,N_19923);
and UO_1076 (O_1076,N_19805,N_19966);
xnor UO_1077 (O_1077,N_19921,N_19835);
nor UO_1078 (O_1078,N_19975,N_19863);
xnor UO_1079 (O_1079,N_19884,N_19973);
nand UO_1080 (O_1080,N_19851,N_19945);
and UO_1081 (O_1081,N_19813,N_19836);
nor UO_1082 (O_1082,N_19878,N_19902);
xnor UO_1083 (O_1083,N_19996,N_19813);
or UO_1084 (O_1084,N_19806,N_19849);
xor UO_1085 (O_1085,N_19828,N_19894);
nand UO_1086 (O_1086,N_19816,N_19883);
nor UO_1087 (O_1087,N_19978,N_19959);
nand UO_1088 (O_1088,N_19963,N_19947);
nand UO_1089 (O_1089,N_19879,N_19911);
xor UO_1090 (O_1090,N_19922,N_19807);
or UO_1091 (O_1091,N_19896,N_19916);
nor UO_1092 (O_1092,N_19875,N_19999);
xor UO_1093 (O_1093,N_19950,N_19882);
or UO_1094 (O_1094,N_19818,N_19935);
or UO_1095 (O_1095,N_19942,N_19883);
and UO_1096 (O_1096,N_19955,N_19875);
and UO_1097 (O_1097,N_19862,N_19838);
nor UO_1098 (O_1098,N_19967,N_19903);
xor UO_1099 (O_1099,N_19946,N_19867);
nor UO_1100 (O_1100,N_19849,N_19867);
nand UO_1101 (O_1101,N_19983,N_19970);
nor UO_1102 (O_1102,N_19887,N_19898);
and UO_1103 (O_1103,N_19969,N_19802);
nand UO_1104 (O_1104,N_19812,N_19875);
nand UO_1105 (O_1105,N_19843,N_19833);
nand UO_1106 (O_1106,N_19917,N_19914);
or UO_1107 (O_1107,N_19907,N_19955);
xor UO_1108 (O_1108,N_19828,N_19879);
xor UO_1109 (O_1109,N_19818,N_19817);
nand UO_1110 (O_1110,N_19832,N_19838);
nor UO_1111 (O_1111,N_19934,N_19963);
nor UO_1112 (O_1112,N_19976,N_19937);
nor UO_1113 (O_1113,N_19965,N_19820);
and UO_1114 (O_1114,N_19907,N_19879);
and UO_1115 (O_1115,N_19807,N_19889);
or UO_1116 (O_1116,N_19909,N_19965);
and UO_1117 (O_1117,N_19861,N_19859);
and UO_1118 (O_1118,N_19850,N_19946);
and UO_1119 (O_1119,N_19852,N_19918);
and UO_1120 (O_1120,N_19800,N_19925);
xnor UO_1121 (O_1121,N_19872,N_19800);
nand UO_1122 (O_1122,N_19865,N_19991);
nand UO_1123 (O_1123,N_19801,N_19860);
or UO_1124 (O_1124,N_19983,N_19930);
and UO_1125 (O_1125,N_19981,N_19878);
and UO_1126 (O_1126,N_19825,N_19831);
nand UO_1127 (O_1127,N_19971,N_19970);
and UO_1128 (O_1128,N_19853,N_19855);
and UO_1129 (O_1129,N_19827,N_19946);
nand UO_1130 (O_1130,N_19904,N_19921);
nand UO_1131 (O_1131,N_19957,N_19953);
and UO_1132 (O_1132,N_19884,N_19925);
nor UO_1133 (O_1133,N_19901,N_19860);
nor UO_1134 (O_1134,N_19864,N_19825);
xnor UO_1135 (O_1135,N_19964,N_19949);
nand UO_1136 (O_1136,N_19865,N_19952);
or UO_1137 (O_1137,N_19886,N_19880);
xor UO_1138 (O_1138,N_19945,N_19844);
xor UO_1139 (O_1139,N_19968,N_19923);
nor UO_1140 (O_1140,N_19846,N_19931);
nor UO_1141 (O_1141,N_19887,N_19958);
or UO_1142 (O_1142,N_19992,N_19870);
and UO_1143 (O_1143,N_19941,N_19927);
nand UO_1144 (O_1144,N_19910,N_19914);
xnor UO_1145 (O_1145,N_19970,N_19840);
nand UO_1146 (O_1146,N_19849,N_19976);
and UO_1147 (O_1147,N_19843,N_19815);
nand UO_1148 (O_1148,N_19828,N_19917);
xor UO_1149 (O_1149,N_19986,N_19854);
nor UO_1150 (O_1150,N_19886,N_19833);
or UO_1151 (O_1151,N_19855,N_19973);
nand UO_1152 (O_1152,N_19908,N_19811);
nor UO_1153 (O_1153,N_19927,N_19959);
nand UO_1154 (O_1154,N_19933,N_19900);
nor UO_1155 (O_1155,N_19845,N_19967);
nand UO_1156 (O_1156,N_19992,N_19856);
nor UO_1157 (O_1157,N_19833,N_19988);
and UO_1158 (O_1158,N_19944,N_19802);
nand UO_1159 (O_1159,N_19826,N_19864);
xor UO_1160 (O_1160,N_19932,N_19894);
and UO_1161 (O_1161,N_19822,N_19936);
nor UO_1162 (O_1162,N_19999,N_19973);
nand UO_1163 (O_1163,N_19857,N_19864);
nor UO_1164 (O_1164,N_19875,N_19891);
xor UO_1165 (O_1165,N_19857,N_19805);
nor UO_1166 (O_1166,N_19842,N_19852);
and UO_1167 (O_1167,N_19841,N_19945);
nand UO_1168 (O_1168,N_19924,N_19974);
nor UO_1169 (O_1169,N_19939,N_19902);
xor UO_1170 (O_1170,N_19992,N_19998);
or UO_1171 (O_1171,N_19995,N_19918);
nor UO_1172 (O_1172,N_19811,N_19899);
or UO_1173 (O_1173,N_19844,N_19935);
and UO_1174 (O_1174,N_19862,N_19974);
nand UO_1175 (O_1175,N_19998,N_19849);
nor UO_1176 (O_1176,N_19804,N_19834);
or UO_1177 (O_1177,N_19914,N_19950);
nor UO_1178 (O_1178,N_19819,N_19970);
nor UO_1179 (O_1179,N_19854,N_19929);
nor UO_1180 (O_1180,N_19838,N_19896);
nor UO_1181 (O_1181,N_19865,N_19958);
or UO_1182 (O_1182,N_19860,N_19916);
xnor UO_1183 (O_1183,N_19908,N_19951);
nand UO_1184 (O_1184,N_19989,N_19949);
or UO_1185 (O_1185,N_19968,N_19997);
nand UO_1186 (O_1186,N_19966,N_19950);
nand UO_1187 (O_1187,N_19906,N_19873);
xor UO_1188 (O_1188,N_19815,N_19838);
nor UO_1189 (O_1189,N_19896,N_19864);
and UO_1190 (O_1190,N_19912,N_19812);
or UO_1191 (O_1191,N_19986,N_19978);
or UO_1192 (O_1192,N_19820,N_19875);
xnor UO_1193 (O_1193,N_19834,N_19955);
nand UO_1194 (O_1194,N_19967,N_19905);
nand UO_1195 (O_1195,N_19987,N_19839);
and UO_1196 (O_1196,N_19990,N_19999);
or UO_1197 (O_1197,N_19817,N_19847);
and UO_1198 (O_1198,N_19829,N_19898);
nor UO_1199 (O_1199,N_19800,N_19863);
xnor UO_1200 (O_1200,N_19954,N_19888);
xor UO_1201 (O_1201,N_19926,N_19859);
or UO_1202 (O_1202,N_19849,N_19831);
xnor UO_1203 (O_1203,N_19965,N_19845);
nand UO_1204 (O_1204,N_19833,N_19985);
xor UO_1205 (O_1205,N_19980,N_19848);
xnor UO_1206 (O_1206,N_19806,N_19976);
nand UO_1207 (O_1207,N_19904,N_19988);
nor UO_1208 (O_1208,N_19845,N_19875);
and UO_1209 (O_1209,N_19906,N_19917);
nor UO_1210 (O_1210,N_19951,N_19830);
nor UO_1211 (O_1211,N_19868,N_19969);
and UO_1212 (O_1212,N_19819,N_19961);
nand UO_1213 (O_1213,N_19971,N_19850);
xor UO_1214 (O_1214,N_19911,N_19999);
or UO_1215 (O_1215,N_19900,N_19931);
xor UO_1216 (O_1216,N_19893,N_19982);
xnor UO_1217 (O_1217,N_19977,N_19956);
nand UO_1218 (O_1218,N_19820,N_19817);
or UO_1219 (O_1219,N_19999,N_19866);
and UO_1220 (O_1220,N_19882,N_19803);
or UO_1221 (O_1221,N_19865,N_19869);
xor UO_1222 (O_1222,N_19990,N_19962);
and UO_1223 (O_1223,N_19807,N_19952);
and UO_1224 (O_1224,N_19845,N_19855);
nor UO_1225 (O_1225,N_19948,N_19892);
nor UO_1226 (O_1226,N_19835,N_19976);
nand UO_1227 (O_1227,N_19981,N_19959);
nor UO_1228 (O_1228,N_19945,N_19918);
xor UO_1229 (O_1229,N_19943,N_19997);
and UO_1230 (O_1230,N_19813,N_19998);
xnor UO_1231 (O_1231,N_19839,N_19978);
or UO_1232 (O_1232,N_19849,N_19832);
xor UO_1233 (O_1233,N_19972,N_19920);
nor UO_1234 (O_1234,N_19993,N_19960);
and UO_1235 (O_1235,N_19977,N_19942);
or UO_1236 (O_1236,N_19987,N_19867);
and UO_1237 (O_1237,N_19894,N_19931);
nand UO_1238 (O_1238,N_19915,N_19891);
and UO_1239 (O_1239,N_19968,N_19876);
and UO_1240 (O_1240,N_19895,N_19962);
xnor UO_1241 (O_1241,N_19841,N_19933);
nor UO_1242 (O_1242,N_19923,N_19997);
nand UO_1243 (O_1243,N_19834,N_19925);
nand UO_1244 (O_1244,N_19817,N_19933);
nand UO_1245 (O_1245,N_19879,N_19801);
nand UO_1246 (O_1246,N_19972,N_19858);
and UO_1247 (O_1247,N_19994,N_19926);
nand UO_1248 (O_1248,N_19985,N_19916);
xor UO_1249 (O_1249,N_19876,N_19916);
xor UO_1250 (O_1250,N_19877,N_19843);
or UO_1251 (O_1251,N_19999,N_19951);
nand UO_1252 (O_1252,N_19856,N_19828);
nand UO_1253 (O_1253,N_19887,N_19955);
xor UO_1254 (O_1254,N_19986,N_19957);
nand UO_1255 (O_1255,N_19999,N_19916);
nand UO_1256 (O_1256,N_19860,N_19855);
or UO_1257 (O_1257,N_19860,N_19970);
nor UO_1258 (O_1258,N_19821,N_19837);
nor UO_1259 (O_1259,N_19916,N_19902);
xor UO_1260 (O_1260,N_19924,N_19831);
nor UO_1261 (O_1261,N_19801,N_19978);
nand UO_1262 (O_1262,N_19881,N_19844);
nand UO_1263 (O_1263,N_19987,N_19968);
and UO_1264 (O_1264,N_19871,N_19924);
nand UO_1265 (O_1265,N_19894,N_19896);
nand UO_1266 (O_1266,N_19908,N_19852);
nor UO_1267 (O_1267,N_19919,N_19932);
and UO_1268 (O_1268,N_19849,N_19927);
and UO_1269 (O_1269,N_19862,N_19868);
and UO_1270 (O_1270,N_19932,N_19889);
or UO_1271 (O_1271,N_19946,N_19981);
or UO_1272 (O_1272,N_19966,N_19921);
nor UO_1273 (O_1273,N_19951,N_19864);
or UO_1274 (O_1274,N_19819,N_19967);
and UO_1275 (O_1275,N_19923,N_19912);
nor UO_1276 (O_1276,N_19970,N_19936);
xnor UO_1277 (O_1277,N_19821,N_19986);
nand UO_1278 (O_1278,N_19917,N_19860);
and UO_1279 (O_1279,N_19984,N_19874);
and UO_1280 (O_1280,N_19844,N_19923);
or UO_1281 (O_1281,N_19918,N_19887);
nor UO_1282 (O_1282,N_19869,N_19934);
xnor UO_1283 (O_1283,N_19925,N_19967);
nor UO_1284 (O_1284,N_19821,N_19949);
nand UO_1285 (O_1285,N_19898,N_19905);
and UO_1286 (O_1286,N_19828,N_19880);
and UO_1287 (O_1287,N_19920,N_19969);
or UO_1288 (O_1288,N_19913,N_19943);
nor UO_1289 (O_1289,N_19805,N_19850);
or UO_1290 (O_1290,N_19822,N_19882);
nand UO_1291 (O_1291,N_19954,N_19977);
and UO_1292 (O_1292,N_19828,N_19841);
nand UO_1293 (O_1293,N_19959,N_19964);
or UO_1294 (O_1294,N_19944,N_19960);
nand UO_1295 (O_1295,N_19993,N_19897);
or UO_1296 (O_1296,N_19890,N_19933);
xor UO_1297 (O_1297,N_19929,N_19928);
nor UO_1298 (O_1298,N_19910,N_19928);
or UO_1299 (O_1299,N_19839,N_19846);
nand UO_1300 (O_1300,N_19985,N_19836);
xnor UO_1301 (O_1301,N_19985,N_19937);
nor UO_1302 (O_1302,N_19896,N_19981);
nor UO_1303 (O_1303,N_19943,N_19966);
nand UO_1304 (O_1304,N_19926,N_19846);
or UO_1305 (O_1305,N_19833,N_19860);
xnor UO_1306 (O_1306,N_19800,N_19856);
and UO_1307 (O_1307,N_19809,N_19913);
xor UO_1308 (O_1308,N_19835,N_19809);
or UO_1309 (O_1309,N_19809,N_19955);
nor UO_1310 (O_1310,N_19856,N_19883);
or UO_1311 (O_1311,N_19853,N_19899);
nor UO_1312 (O_1312,N_19821,N_19936);
and UO_1313 (O_1313,N_19933,N_19951);
nand UO_1314 (O_1314,N_19856,N_19914);
nand UO_1315 (O_1315,N_19997,N_19870);
nand UO_1316 (O_1316,N_19983,N_19985);
nor UO_1317 (O_1317,N_19900,N_19889);
or UO_1318 (O_1318,N_19945,N_19999);
nor UO_1319 (O_1319,N_19931,N_19927);
xnor UO_1320 (O_1320,N_19894,N_19816);
and UO_1321 (O_1321,N_19915,N_19986);
nor UO_1322 (O_1322,N_19988,N_19903);
or UO_1323 (O_1323,N_19865,N_19824);
and UO_1324 (O_1324,N_19905,N_19826);
and UO_1325 (O_1325,N_19924,N_19826);
xnor UO_1326 (O_1326,N_19941,N_19898);
nor UO_1327 (O_1327,N_19832,N_19912);
nand UO_1328 (O_1328,N_19820,N_19957);
xor UO_1329 (O_1329,N_19950,N_19838);
and UO_1330 (O_1330,N_19937,N_19904);
or UO_1331 (O_1331,N_19894,N_19991);
or UO_1332 (O_1332,N_19882,N_19859);
nand UO_1333 (O_1333,N_19814,N_19983);
and UO_1334 (O_1334,N_19909,N_19949);
or UO_1335 (O_1335,N_19808,N_19801);
xnor UO_1336 (O_1336,N_19937,N_19980);
nor UO_1337 (O_1337,N_19826,N_19890);
xor UO_1338 (O_1338,N_19925,N_19880);
and UO_1339 (O_1339,N_19907,N_19834);
and UO_1340 (O_1340,N_19872,N_19889);
or UO_1341 (O_1341,N_19855,N_19921);
nand UO_1342 (O_1342,N_19895,N_19922);
nand UO_1343 (O_1343,N_19901,N_19885);
nor UO_1344 (O_1344,N_19993,N_19956);
nand UO_1345 (O_1345,N_19971,N_19982);
xnor UO_1346 (O_1346,N_19857,N_19975);
or UO_1347 (O_1347,N_19993,N_19996);
nand UO_1348 (O_1348,N_19853,N_19910);
or UO_1349 (O_1349,N_19934,N_19880);
nand UO_1350 (O_1350,N_19844,N_19911);
xnor UO_1351 (O_1351,N_19963,N_19964);
or UO_1352 (O_1352,N_19900,N_19953);
nor UO_1353 (O_1353,N_19913,N_19864);
or UO_1354 (O_1354,N_19854,N_19897);
or UO_1355 (O_1355,N_19923,N_19933);
nand UO_1356 (O_1356,N_19919,N_19979);
and UO_1357 (O_1357,N_19804,N_19902);
nor UO_1358 (O_1358,N_19802,N_19910);
and UO_1359 (O_1359,N_19955,N_19820);
and UO_1360 (O_1360,N_19879,N_19927);
xor UO_1361 (O_1361,N_19872,N_19923);
and UO_1362 (O_1362,N_19906,N_19913);
and UO_1363 (O_1363,N_19931,N_19855);
nor UO_1364 (O_1364,N_19836,N_19879);
nand UO_1365 (O_1365,N_19850,N_19938);
nand UO_1366 (O_1366,N_19804,N_19954);
xnor UO_1367 (O_1367,N_19963,N_19852);
or UO_1368 (O_1368,N_19819,N_19875);
or UO_1369 (O_1369,N_19968,N_19806);
and UO_1370 (O_1370,N_19969,N_19849);
and UO_1371 (O_1371,N_19938,N_19979);
nor UO_1372 (O_1372,N_19956,N_19972);
or UO_1373 (O_1373,N_19965,N_19913);
and UO_1374 (O_1374,N_19894,N_19960);
and UO_1375 (O_1375,N_19989,N_19863);
and UO_1376 (O_1376,N_19986,N_19841);
nand UO_1377 (O_1377,N_19815,N_19896);
or UO_1378 (O_1378,N_19804,N_19912);
xor UO_1379 (O_1379,N_19906,N_19815);
or UO_1380 (O_1380,N_19850,N_19862);
nand UO_1381 (O_1381,N_19867,N_19918);
xnor UO_1382 (O_1382,N_19936,N_19819);
nor UO_1383 (O_1383,N_19881,N_19991);
xnor UO_1384 (O_1384,N_19829,N_19931);
or UO_1385 (O_1385,N_19938,N_19907);
and UO_1386 (O_1386,N_19825,N_19886);
xor UO_1387 (O_1387,N_19831,N_19808);
or UO_1388 (O_1388,N_19833,N_19800);
and UO_1389 (O_1389,N_19927,N_19917);
xor UO_1390 (O_1390,N_19882,N_19892);
and UO_1391 (O_1391,N_19881,N_19840);
nor UO_1392 (O_1392,N_19819,N_19878);
nor UO_1393 (O_1393,N_19887,N_19985);
nor UO_1394 (O_1394,N_19804,N_19953);
and UO_1395 (O_1395,N_19900,N_19944);
nand UO_1396 (O_1396,N_19816,N_19922);
nor UO_1397 (O_1397,N_19979,N_19937);
nand UO_1398 (O_1398,N_19823,N_19884);
and UO_1399 (O_1399,N_19852,N_19929);
or UO_1400 (O_1400,N_19927,N_19909);
nor UO_1401 (O_1401,N_19930,N_19910);
and UO_1402 (O_1402,N_19909,N_19912);
xor UO_1403 (O_1403,N_19833,N_19951);
or UO_1404 (O_1404,N_19854,N_19834);
nor UO_1405 (O_1405,N_19954,N_19969);
nand UO_1406 (O_1406,N_19989,N_19903);
xor UO_1407 (O_1407,N_19836,N_19901);
and UO_1408 (O_1408,N_19957,N_19943);
or UO_1409 (O_1409,N_19971,N_19846);
xor UO_1410 (O_1410,N_19808,N_19856);
nand UO_1411 (O_1411,N_19911,N_19937);
and UO_1412 (O_1412,N_19825,N_19979);
xnor UO_1413 (O_1413,N_19893,N_19992);
nor UO_1414 (O_1414,N_19807,N_19818);
or UO_1415 (O_1415,N_19887,N_19934);
xnor UO_1416 (O_1416,N_19877,N_19901);
nor UO_1417 (O_1417,N_19919,N_19937);
and UO_1418 (O_1418,N_19879,N_19867);
or UO_1419 (O_1419,N_19851,N_19932);
nand UO_1420 (O_1420,N_19902,N_19824);
and UO_1421 (O_1421,N_19860,N_19972);
nand UO_1422 (O_1422,N_19835,N_19987);
nand UO_1423 (O_1423,N_19998,N_19856);
and UO_1424 (O_1424,N_19902,N_19926);
xor UO_1425 (O_1425,N_19949,N_19915);
nor UO_1426 (O_1426,N_19842,N_19996);
or UO_1427 (O_1427,N_19898,N_19867);
xnor UO_1428 (O_1428,N_19838,N_19873);
nand UO_1429 (O_1429,N_19851,N_19963);
nand UO_1430 (O_1430,N_19980,N_19921);
nand UO_1431 (O_1431,N_19819,N_19948);
or UO_1432 (O_1432,N_19938,N_19804);
nand UO_1433 (O_1433,N_19913,N_19878);
xnor UO_1434 (O_1434,N_19812,N_19936);
nand UO_1435 (O_1435,N_19914,N_19846);
xor UO_1436 (O_1436,N_19911,N_19931);
and UO_1437 (O_1437,N_19945,N_19895);
nor UO_1438 (O_1438,N_19855,N_19903);
and UO_1439 (O_1439,N_19979,N_19803);
nor UO_1440 (O_1440,N_19854,N_19908);
nor UO_1441 (O_1441,N_19895,N_19833);
nor UO_1442 (O_1442,N_19815,N_19921);
nor UO_1443 (O_1443,N_19982,N_19904);
nor UO_1444 (O_1444,N_19870,N_19994);
nand UO_1445 (O_1445,N_19926,N_19987);
and UO_1446 (O_1446,N_19817,N_19961);
nand UO_1447 (O_1447,N_19865,N_19839);
or UO_1448 (O_1448,N_19976,N_19821);
nor UO_1449 (O_1449,N_19816,N_19828);
nor UO_1450 (O_1450,N_19987,N_19978);
and UO_1451 (O_1451,N_19934,N_19815);
nor UO_1452 (O_1452,N_19841,N_19832);
nand UO_1453 (O_1453,N_19806,N_19853);
and UO_1454 (O_1454,N_19817,N_19984);
nor UO_1455 (O_1455,N_19857,N_19891);
and UO_1456 (O_1456,N_19866,N_19806);
and UO_1457 (O_1457,N_19970,N_19921);
or UO_1458 (O_1458,N_19938,N_19838);
nor UO_1459 (O_1459,N_19972,N_19985);
nor UO_1460 (O_1460,N_19908,N_19823);
nand UO_1461 (O_1461,N_19900,N_19912);
nor UO_1462 (O_1462,N_19927,N_19890);
or UO_1463 (O_1463,N_19900,N_19807);
xnor UO_1464 (O_1464,N_19840,N_19909);
nor UO_1465 (O_1465,N_19918,N_19944);
xor UO_1466 (O_1466,N_19801,N_19923);
nand UO_1467 (O_1467,N_19844,N_19971);
nand UO_1468 (O_1468,N_19810,N_19947);
nand UO_1469 (O_1469,N_19862,N_19962);
nand UO_1470 (O_1470,N_19921,N_19972);
or UO_1471 (O_1471,N_19853,N_19994);
or UO_1472 (O_1472,N_19996,N_19988);
nand UO_1473 (O_1473,N_19945,N_19858);
and UO_1474 (O_1474,N_19944,N_19922);
nand UO_1475 (O_1475,N_19908,N_19816);
nand UO_1476 (O_1476,N_19965,N_19949);
xor UO_1477 (O_1477,N_19946,N_19988);
nor UO_1478 (O_1478,N_19928,N_19881);
and UO_1479 (O_1479,N_19995,N_19972);
nand UO_1480 (O_1480,N_19964,N_19907);
or UO_1481 (O_1481,N_19832,N_19809);
and UO_1482 (O_1482,N_19980,N_19991);
xnor UO_1483 (O_1483,N_19979,N_19992);
and UO_1484 (O_1484,N_19984,N_19904);
xnor UO_1485 (O_1485,N_19889,N_19862);
xor UO_1486 (O_1486,N_19949,N_19924);
and UO_1487 (O_1487,N_19899,N_19951);
or UO_1488 (O_1488,N_19972,N_19949);
or UO_1489 (O_1489,N_19902,N_19991);
xor UO_1490 (O_1490,N_19958,N_19869);
or UO_1491 (O_1491,N_19918,N_19979);
and UO_1492 (O_1492,N_19951,N_19938);
nand UO_1493 (O_1493,N_19856,N_19974);
nand UO_1494 (O_1494,N_19952,N_19973);
and UO_1495 (O_1495,N_19921,N_19800);
xor UO_1496 (O_1496,N_19820,N_19852);
and UO_1497 (O_1497,N_19951,N_19963);
nand UO_1498 (O_1498,N_19946,N_19960);
xnor UO_1499 (O_1499,N_19983,N_19987);
or UO_1500 (O_1500,N_19818,N_19983);
xor UO_1501 (O_1501,N_19862,N_19980);
nor UO_1502 (O_1502,N_19993,N_19985);
xor UO_1503 (O_1503,N_19977,N_19871);
nand UO_1504 (O_1504,N_19974,N_19922);
nand UO_1505 (O_1505,N_19828,N_19944);
nor UO_1506 (O_1506,N_19856,N_19804);
or UO_1507 (O_1507,N_19897,N_19910);
nor UO_1508 (O_1508,N_19989,N_19857);
nor UO_1509 (O_1509,N_19959,N_19982);
nand UO_1510 (O_1510,N_19998,N_19884);
xor UO_1511 (O_1511,N_19888,N_19846);
or UO_1512 (O_1512,N_19910,N_19984);
or UO_1513 (O_1513,N_19841,N_19927);
and UO_1514 (O_1514,N_19947,N_19928);
nand UO_1515 (O_1515,N_19865,N_19884);
nand UO_1516 (O_1516,N_19999,N_19871);
nor UO_1517 (O_1517,N_19900,N_19960);
nor UO_1518 (O_1518,N_19923,N_19956);
nand UO_1519 (O_1519,N_19851,N_19914);
and UO_1520 (O_1520,N_19844,N_19926);
or UO_1521 (O_1521,N_19870,N_19919);
or UO_1522 (O_1522,N_19871,N_19835);
xor UO_1523 (O_1523,N_19999,N_19848);
or UO_1524 (O_1524,N_19837,N_19913);
xor UO_1525 (O_1525,N_19902,N_19826);
nor UO_1526 (O_1526,N_19992,N_19921);
nand UO_1527 (O_1527,N_19969,N_19922);
nor UO_1528 (O_1528,N_19840,N_19939);
or UO_1529 (O_1529,N_19960,N_19918);
or UO_1530 (O_1530,N_19847,N_19982);
nand UO_1531 (O_1531,N_19886,N_19861);
and UO_1532 (O_1532,N_19951,N_19875);
nor UO_1533 (O_1533,N_19872,N_19938);
or UO_1534 (O_1534,N_19991,N_19896);
xor UO_1535 (O_1535,N_19949,N_19910);
nor UO_1536 (O_1536,N_19841,N_19937);
nand UO_1537 (O_1537,N_19876,N_19944);
and UO_1538 (O_1538,N_19840,N_19882);
and UO_1539 (O_1539,N_19832,N_19825);
nand UO_1540 (O_1540,N_19942,N_19800);
and UO_1541 (O_1541,N_19840,N_19816);
or UO_1542 (O_1542,N_19934,N_19975);
nand UO_1543 (O_1543,N_19992,N_19885);
xnor UO_1544 (O_1544,N_19940,N_19881);
and UO_1545 (O_1545,N_19959,N_19810);
nand UO_1546 (O_1546,N_19808,N_19810);
or UO_1547 (O_1547,N_19811,N_19847);
nor UO_1548 (O_1548,N_19902,N_19912);
nand UO_1549 (O_1549,N_19996,N_19987);
nor UO_1550 (O_1550,N_19809,N_19800);
nor UO_1551 (O_1551,N_19932,N_19948);
nor UO_1552 (O_1552,N_19823,N_19949);
or UO_1553 (O_1553,N_19840,N_19969);
or UO_1554 (O_1554,N_19913,N_19851);
nor UO_1555 (O_1555,N_19995,N_19888);
xnor UO_1556 (O_1556,N_19900,N_19844);
and UO_1557 (O_1557,N_19932,N_19846);
nor UO_1558 (O_1558,N_19844,N_19835);
or UO_1559 (O_1559,N_19828,N_19842);
and UO_1560 (O_1560,N_19802,N_19922);
and UO_1561 (O_1561,N_19873,N_19996);
nand UO_1562 (O_1562,N_19974,N_19872);
xnor UO_1563 (O_1563,N_19876,N_19902);
nand UO_1564 (O_1564,N_19939,N_19900);
nand UO_1565 (O_1565,N_19882,N_19890);
nand UO_1566 (O_1566,N_19912,N_19957);
and UO_1567 (O_1567,N_19805,N_19816);
and UO_1568 (O_1568,N_19858,N_19842);
xnor UO_1569 (O_1569,N_19967,N_19997);
or UO_1570 (O_1570,N_19990,N_19892);
nor UO_1571 (O_1571,N_19853,N_19902);
nor UO_1572 (O_1572,N_19985,N_19857);
or UO_1573 (O_1573,N_19924,N_19922);
or UO_1574 (O_1574,N_19897,N_19981);
nor UO_1575 (O_1575,N_19883,N_19857);
nor UO_1576 (O_1576,N_19892,N_19944);
xnor UO_1577 (O_1577,N_19926,N_19966);
and UO_1578 (O_1578,N_19923,N_19922);
nand UO_1579 (O_1579,N_19853,N_19932);
nor UO_1580 (O_1580,N_19870,N_19964);
nor UO_1581 (O_1581,N_19971,N_19882);
nand UO_1582 (O_1582,N_19859,N_19801);
or UO_1583 (O_1583,N_19972,N_19881);
nand UO_1584 (O_1584,N_19862,N_19814);
and UO_1585 (O_1585,N_19822,N_19891);
nor UO_1586 (O_1586,N_19845,N_19979);
or UO_1587 (O_1587,N_19820,N_19826);
nor UO_1588 (O_1588,N_19981,N_19831);
or UO_1589 (O_1589,N_19934,N_19819);
nand UO_1590 (O_1590,N_19949,N_19906);
nor UO_1591 (O_1591,N_19836,N_19837);
nand UO_1592 (O_1592,N_19966,N_19912);
nand UO_1593 (O_1593,N_19909,N_19863);
and UO_1594 (O_1594,N_19812,N_19979);
xnor UO_1595 (O_1595,N_19968,N_19850);
nor UO_1596 (O_1596,N_19985,N_19901);
xor UO_1597 (O_1597,N_19873,N_19802);
nor UO_1598 (O_1598,N_19944,N_19931);
nor UO_1599 (O_1599,N_19832,N_19820);
nor UO_1600 (O_1600,N_19857,N_19918);
and UO_1601 (O_1601,N_19973,N_19818);
and UO_1602 (O_1602,N_19938,N_19929);
nand UO_1603 (O_1603,N_19951,N_19942);
nand UO_1604 (O_1604,N_19984,N_19911);
and UO_1605 (O_1605,N_19811,N_19990);
or UO_1606 (O_1606,N_19822,N_19945);
nor UO_1607 (O_1607,N_19976,N_19857);
and UO_1608 (O_1608,N_19809,N_19929);
and UO_1609 (O_1609,N_19975,N_19907);
xnor UO_1610 (O_1610,N_19982,N_19811);
or UO_1611 (O_1611,N_19992,N_19970);
nand UO_1612 (O_1612,N_19844,N_19937);
and UO_1613 (O_1613,N_19815,N_19933);
or UO_1614 (O_1614,N_19839,N_19917);
and UO_1615 (O_1615,N_19883,N_19849);
xor UO_1616 (O_1616,N_19837,N_19882);
nor UO_1617 (O_1617,N_19867,N_19901);
nor UO_1618 (O_1618,N_19928,N_19937);
nor UO_1619 (O_1619,N_19811,N_19946);
and UO_1620 (O_1620,N_19895,N_19930);
or UO_1621 (O_1621,N_19961,N_19999);
nand UO_1622 (O_1622,N_19955,N_19811);
nand UO_1623 (O_1623,N_19945,N_19817);
xor UO_1624 (O_1624,N_19989,N_19926);
or UO_1625 (O_1625,N_19825,N_19877);
xnor UO_1626 (O_1626,N_19883,N_19948);
or UO_1627 (O_1627,N_19829,N_19954);
nor UO_1628 (O_1628,N_19974,N_19860);
nor UO_1629 (O_1629,N_19810,N_19881);
or UO_1630 (O_1630,N_19872,N_19860);
nor UO_1631 (O_1631,N_19871,N_19998);
xor UO_1632 (O_1632,N_19819,N_19938);
or UO_1633 (O_1633,N_19809,N_19971);
nor UO_1634 (O_1634,N_19857,N_19853);
or UO_1635 (O_1635,N_19984,N_19836);
or UO_1636 (O_1636,N_19845,N_19898);
and UO_1637 (O_1637,N_19888,N_19884);
nor UO_1638 (O_1638,N_19867,N_19975);
xor UO_1639 (O_1639,N_19810,N_19995);
nand UO_1640 (O_1640,N_19984,N_19818);
or UO_1641 (O_1641,N_19898,N_19833);
nand UO_1642 (O_1642,N_19882,N_19910);
nor UO_1643 (O_1643,N_19940,N_19876);
or UO_1644 (O_1644,N_19813,N_19850);
or UO_1645 (O_1645,N_19801,N_19932);
nand UO_1646 (O_1646,N_19943,N_19856);
nor UO_1647 (O_1647,N_19976,N_19878);
nor UO_1648 (O_1648,N_19939,N_19839);
nor UO_1649 (O_1649,N_19805,N_19903);
xor UO_1650 (O_1650,N_19852,N_19873);
and UO_1651 (O_1651,N_19964,N_19894);
or UO_1652 (O_1652,N_19866,N_19948);
nor UO_1653 (O_1653,N_19975,N_19918);
xor UO_1654 (O_1654,N_19961,N_19940);
xor UO_1655 (O_1655,N_19963,N_19833);
xor UO_1656 (O_1656,N_19856,N_19953);
or UO_1657 (O_1657,N_19942,N_19829);
xnor UO_1658 (O_1658,N_19981,N_19822);
or UO_1659 (O_1659,N_19916,N_19998);
and UO_1660 (O_1660,N_19961,N_19879);
xnor UO_1661 (O_1661,N_19999,N_19962);
nand UO_1662 (O_1662,N_19954,N_19948);
or UO_1663 (O_1663,N_19853,N_19882);
nor UO_1664 (O_1664,N_19813,N_19903);
xnor UO_1665 (O_1665,N_19806,N_19818);
xnor UO_1666 (O_1666,N_19911,N_19860);
xnor UO_1667 (O_1667,N_19843,N_19938);
xnor UO_1668 (O_1668,N_19826,N_19832);
nor UO_1669 (O_1669,N_19996,N_19925);
and UO_1670 (O_1670,N_19864,N_19970);
and UO_1671 (O_1671,N_19962,N_19804);
nand UO_1672 (O_1672,N_19921,N_19851);
or UO_1673 (O_1673,N_19818,N_19916);
xor UO_1674 (O_1674,N_19902,N_19975);
nand UO_1675 (O_1675,N_19927,N_19967);
nand UO_1676 (O_1676,N_19847,N_19932);
nor UO_1677 (O_1677,N_19978,N_19943);
or UO_1678 (O_1678,N_19872,N_19901);
nor UO_1679 (O_1679,N_19886,N_19900);
nand UO_1680 (O_1680,N_19817,N_19894);
nand UO_1681 (O_1681,N_19963,N_19831);
and UO_1682 (O_1682,N_19820,N_19899);
and UO_1683 (O_1683,N_19868,N_19867);
nor UO_1684 (O_1684,N_19903,N_19943);
and UO_1685 (O_1685,N_19998,N_19956);
and UO_1686 (O_1686,N_19966,N_19888);
nor UO_1687 (O_1687,N_19967,N_19959);
or UO_1688 (O_1688,N_19940,N_19868);
and UO_1689 (O_1689,N_19891,N_19958);
or UO_1690 (O_1690,N_19875,N_19803);
nor UO_1691 (O_1691,N_19871,N_19836);
or UO_1692 (O_1692,N_19862,N_19836);
and UO_1693 (O_1693,N_19892,N_19969);
or UO_1694 (O_1694,N_19966,N_19829);
or UO_1695 (O_1695,N_19802,N_19998);
and UO_1696 (O_1696,N_19949,N_19879);
nor UO_1697 (O_1697,N_19870,N_19980);
nand UO_1698 (O_1698,N_19857,N_19935);
and UO_1699 (O_1699,N_19919,N_19941);
xnor UO_1700 (O_1700,N_19859,N_19870);
nand UO_1701 (O_1701,N_19971,N_19904);
xor UO_1702 (O_1702,N_19930,N_19849);
nand UO_1703 (O_1703,N_19988,N_19898);
nand UO_1704 (O_1704,N_19953,N_19847);
or UO_1705 (O_1705,N_19866,N_19892);
xor UO_1706 (O_1706,N_19971,N_19910);
or UO_1707 (O_1707,N_19892,N_19935);
nand UO_1708 (O_1708,N_19879,N_19947);
or UO_1709 (O_1709,N_19819,N_19818);
or UO_1710 (O_1710,N_19971,N_19913);
and UO_1711 (O_1711,N_19863,N_19965);
nand UO_1712 (O_1712,N_19917,N_19810);
xor UO_1713 (O_1713,N_19979,N_19961);
xnor UO_1714 (O_1714,N_19940,N_19924);
and UO_1715 (O_1715,N_19853,N_19817);
nor UO_1716 (O_1716,N_19807,N_19971);
and UO_1717 (O_1717,N_19996,N_19904);
or UO_1718 (O_1718,N_19801,N_19870);
nand UO_1719 (O_1719,N_19847,N_19833);
and UO_1720 (O_1720,N_19920,N_19843);
xor UO_1721 (O_1721,N_19829,N_19912);
xnor UO_1722 (O_1722,N_19895,N_19917);
nand UO_1723 (O_1723,N_19901,N_19968);
xnor UO_1724 (O_1724,N_19873,N_19931);
nor UO_1725 (O_1725,N_19927,N_19942);
and UO_1726 (O_1726,N_19953,N_19996);
nand UO_1727 (O_1727,N_19815,N_19920);
and UO_1728 (O_1728,N_19947,N_19964);
or UO_1729 (O_1729,N_19968,N_19903);
nand UO_1730 (O_1730,N_19916,N_19855);
nor UO_1731 (O_1731,N_19975,N_19823);
and UO_1732 (O_1732,N_19849,N_19809);
and UO_1733 (O_1733,N_19942,N_19824);
and UO_1734 (O_1734,N_19843,N_19915);
and UO_1735 (O_1735,N_19847,N_19894);
or UO_1736 (O_1736,N_19951,N_19896);
nor UO_1737 (O_1737,N_19935,N_19872);
nand UO_1738 (O_1738,N_19822,N_19848);
or UO_1739 (O_1739,N_19909,N_19893);
nor UO_1740 (O_1740,N_19882,N_19827);
xnor UO_1741 (O_1741,N_19895,N_19819);
xnor UO_1742 (O_1742,N_19883,N_19924);
or UO_1743 (O_1743,N_19919,N_19876);
xnor UO_1744 (O_1744,N_19829,N_19895);
or UO_1745 (O_1745,N_19922,N_19993);
nand UO_1746 (O_1746,N_19932,N_19996);
nor UO_1747 (O_1747,N_19866,N_19862);
nand UO_1748 (O_1748,N_19970,N_19916);
nand UO_1749 (O_1749,N_19817,N_19829);
nand UO_1750 (O_1750,N_19945,N_19831);
or UO_1751 (O_1751,N_19994,N_19976);
nor UO_1752 (O_1752,N_19957,N_19842);
nand UO_1753 (O_1753,N_19955,N_19876);
nand UO_1754 (O_1754,N_19846,N_19832);
xnor UO_1755 (O_1755,N_19917,N_19994);
xor UO_1756 (O_1756,N_19818,N_19958);
nand UO_1757 (O_1757,N_19817,N_19844);
and UO_1758 (O_1758,N_19852,N_19950);
xor UO_1759 (O_1759,N_19849,N_19922);
or UO_1760 (O_1760,N_19994,N_19814);
xnor UO_1761 (O_1761,N_19919,N_19948);
xor UO_1762 (O_1762,N_19880,N_19960);
nor UO_1763 (O_1763,N_19965,N_19960);
and UO_1764 (O_1764,N_19804,N_19963);
nor UO_1765 (O_1765,N_19886,N_19897);
nand UO_1766 (O_1766,N_19891,N_19957);
xnor UO_1767 (O_1767,N_19860,N_19871);
xor UO_1768 (O_1768,N_19885,N_19934);
or UO_1769 (O_1769,N_19816,N_19819);
and UO_1770 (O_1770,N_19890,N_19899);
xor UO_1771 (O_1771,N_19951,N_19819);
or UO_1772 (O_1772,N_19813,N_19871);
xor UO_1773 (O_1773,N_19875,N_19827);
nor UO_1774 (O_1774,N_19823,N_19835);
nor UO_1775 (O_1775,N_19844,N_19895);
xor UO_1776 (O_1776,N_19949,N_19996);
nand UO_1777 (O_1777,N_19804,N_19925);
or UO_1778 (O_1778,N_19940,N_19889);
or UO_1779 (O_1779,N_19847,N_19882);
or UO_1780 (O_1780,N_19959,N_19985);
nor UO_1781 (O_1781,N_19902,N_19988);
xor UO_1782 (O_1782,N_19947,N_19940);
or UO_1783 (O_1783,N_19904,N_19968);
xnor UO_1784 (O_1784,N_19905,N_19955);
xnor UO_1785 (O_1785,N_19892,N_19922);
nor UO_1786 (O_1786,N_19941,N_19905);
nor UO_1787 (O_1787,N_19979,N_19924);
or UO_1788 (O_1788,N_19877,N_19914);
and UO_1789 (O_1789,N_19920,N_19955);
nand UO_1790 (O_1790,N_19871,N_19826);
nand UO_1791 (O_1791,N_19958,N_19872);
nor UO_1792 (O_1792,N_19941,N_19894);
and UO_1793 (O_1793,N_19868,N_19934);
nor UO_1794 (O_1794,N_19972,N_19808);
nor UO_1795 (O_1795,N_19983,N_19964);
and UO_1796 (O_1796,N_19883,N_19812);
and UO_1797 (O_1797,N_19858,N_19887);
nor UO_1798 (O_1798,N_19837,N_19877);
nand UO_1799 (O_1799,N_19897,N_19843);
nand UO_1800 (O_1800,N_19842,N_19854);
and UO_1801 (O_1801,N_19867,N_19928);
nand UO_1802 (O_1802,N_19896,N_19958);
or UO_1803 (O_1803,N_19985,N_19913);
and UO_1804 (O_1804,N_19896,N_19898);
or UO_1805 (O_1805,N_19886,N_19983);
nand UO_1806 (O_1806,N_19925,N_19896);
and UO_1807 (O_1807,N_19861,N_19933);
and UO_1808 (O_1808,N_19967,N_19832);
nand UO_1809 (O_1809,N_19866,N_19910);
nand UO_1810 (O_1810,N_19831,N_19961);
and UO_1811 (O_1811,N_19913,N_19950);
or UO_1812 (O_1812,N_19885,N_19951);
xor UO_1813 (O_1813,N_19985,N_19949);
or UO_1814 (O_1814,N_19967,N_19837);
nor UO_1815 (O_1815,N_19995,N_19861);
nand UO_1816 (O_1816,N_19826,N_19957);
nand UO_1817 (O_1817,N_19974,N_19906);
nor UO_1818 (O_1818,N_19939,N_19811);
nor UO_1819 (O_1819,N_19946,N_19835);
nand UO_1820 (O_1820,N_19960,N_19936);
xor UO_1821 (O_1821,N_19899,N_19991);
or UO_1822 (O_1822,N_19821,N_19807);
and UO_1823 (O_1823,N_19806,N_19852);
or UO_1824 (O_1824,N_19912,N_19826);
nor UO_1825 (O_1825,N_19961,N_19848);
and UO_1826 (O_1826,N_19811,N_19967);
or UO_1827 (O_1827,N_19955,N_19837);
or UO_1828 (O_1828,N_19981,N_19921);
xor UO_1829 (O_1829,N_19946,N_19998);
nand UO_1830 (O_1830,N_19802,N_19939);
nor UO_1831 (O_1831,N_19944,N_19889);
nand UO_1832 (O_1832,N_19839,N_19838);
or UO_1833 (O_1833,N_19954,N_19868);
xnor UO_1834 (O_1834,N_19933,N_19913);
xor UO_1835 (O_1835,N_19883,N_19823);
xor UO_1836 (O_1836,N_19819,N_19908);
nor UO_1837 (O_1837,N_19988,N_19974);
nor UO_1838 (O_1838,N_19930,N_19865);
and UO_1839 (O_1839,N_19950,N_19872);
xor UO_1840 (O_1840,N_19958,N_19962);
xnor UO_1841 (O_1841,N_19949,N_19947);
nor UO_1842 (O_1842,N_19893,N_19917);
xnor UO_1843 (O_1843,N_19813,N_19895);
nor UO_1844 (O_1844,N_19855,N_19857);
and UO_1845 (O_1845,N_19831,N_19929);
xnor UO_1846 (O_1846,N_19817,N_19899);
nand UO_1847 (O_1847,N_19818,N_19835);
or UO_1848 (O_1848,N_19866,N_19872);
nor UO_1849 (O_1849,N_19807,N_19901);
and UO_1850 (O_1850,N_19907,N_19922);
or UO_1851 (O_1851,N_19943,N_19843);
and UO_1852 (O_1852,N_19896,N_19845);
xor UO_1853 (O_1853,N_19824,N_19972);
nand UO_1854 (O_1854,N_19922,N_19962);
or UO_1855 (O_1855,N_19952,N_19955);
or UO_1856 (O_1856,N_19803,N_19962);
or UO_1857 (O_1857,N_19832,N_19980);
nand UO_1858 (O_1858,N_19928,N_19800);
nand UO_1859 (O_1859,N_19831,N_19907);
nand UO_1860 (O_1860,N_19895,N_19849);
and UO_1861 (O_1861,N_19839,N_19891);
and UO_1862 (O_1862,N_19959,N_19909);
nor UO_1863 (O_1863,N_19886,N_19935);
or UO_1864 (O_1864,N_19921,N_19979);
nand UO_1865 (O_1865,N_19884,N_19961);
and UO_1866 (O_1866,N_19954,N_19897);
xnor UO_1867 (O_1867,N_19892,N_19898);
and UO_1868 (O_1868,N_19978,N_19929);
and UO_1869 (O_1869,N_19841,N_19897);
xor UO_1870 (O_1870,N_19988,N_19883);
or UO_1871 (O_1871,N_19829,N_19909);
and UO_1872 (O_1872,N_19926,N_19912);
or UO_1873 (O_1873,N_19914,N_19962);
or UO_1874 (O_1874,N_19864,N_19963);
or UO_1875 (O_1875,N_19807,N_19850);
or UO_1876 (O_1876,N_19831,N_19984);
nor UO_1877 (O_1877,N_19902,N_19950);
or UO_1878 (O_1878,N_19866,N_19886);
and UO_1879 (O_1879,N_19913,N_19823);
or UO_1880 (O_1880,N_19876,N_19816);
nand UO_1881 (O_1881,N_19831,N_19852);
xor UO_1882 (O_1882,N_19952,N_19894);
or UO_1883 (O_1883,N_19847,N_19863);
nand UO_1884 (O_1884,N_19951,N_19890);
xor UO_1885 (O_1885,N_19963,N_19845);
and UO_1886 (O_1886,N_19909,N_19907);
nor UO_1887 (O_1887,N_19854,N_19894);
and UO_1888 (O_1888,N_19829,N_19995);
nor UO_1889 (O_1889,N_19809,N_19976);
nand UO_1890 (O_1890,N_19858,N_19992);
xor UO_1891 (O_1891,N_19891,N_19836);
or UO_1892 (O_1892,N_19886,N_19955);
or UO_1893 (O_1893,N_19897,N_19959);
xnor UO_1894 (O_1894,N_19980,N_19906);
xnor UO_1895 (O_1895,N_19862,N_19857);
nand UO_1896 (O_1896,N_19800,N_19888);
and UO_1897 (O_1897,N_19917,N_19905);
or UO_1898 (O_1898,N_19923,N_19901);
or UO_1899 (O_1899,N_19886,N_19883);
nand UO_1900 (O_1900,N_19833,N_19938);
xnor UO_1901 (O_1901,N_19863,N_19833);
and UO_1902 (O_1902,N_19844,N_19892);
and UO_1903 (O_1903,N_19834,N_19990);
nor UO_1904 (O_1904,N_19985,N_19847);
nand UO_1905 (O_1905,N_19808,N_19871);
and UO_1906 (O_1906,N_19903,N_19948);
and UO_1907 (O_1907,N_19880,N_19929);
xor UO_1908 (O_1908,N_19965,N_19944);
nor UO_1909 (O_1909,N_19907,N_19853);
nand UO_1910 (O_1910,N_19948,N_19864);
xnor UO_1911 (O_1911,N_19837,N_19806);
and UO_1912 (O_1912,N_19820,N_19961);
or UO_1913 (O_1913,N_19982,N_19958);
or UO_1914 (O_1914,N_19934,N_19804);
nand UO_1915 (O_1915,N_19898,N_19951);
and UO_1916 (O_1916,N_19991,N_19872);
nor UO_1917 (O_1917,N_19842,N_19977);
nand UO_1918 (O_1918,N_19894,N_19916);
nor UO_1919 (O_1919,N_19805,N_19859);
nor UO_1920 (O_1920,N_19967,N_19964);
and UO_1921 (O_1921,N_19856,N_19968);
nand UO_1922 (O_1922,N_19960,N_19858);
or UO_1923 (O_1923,N_19924,N_19860);
or UO_1924 (O_1924,N_19935,N_19972);
xnor UO_1925 (O_1925,N_19810,N_19817);
xnor UO_1926 (O_1926,N_19891,N_19811);
nor UO_1927 (O_1927,N_19910,N_19831);
and UO_1928 (O_1928,N_19872,N_19814);
nor UO_1929 (O_1929,N_19878,N_19810);
nand UO_1930 (O_1930,N_19804,N_19910);
or UO_1931 (O_1931,N_19995,N_19850);
nand UO_1932 (O_1932,N_19944,N_19882);
and UO_1933 (O_1933,N_19852,N_19870);
or UO_1934 (O_1934,N_19944,N_19983);
nand UO_1935 (O_1935,N_19800,N_19828);
xnor UO_1936 (O_1936,N_19981,N_19969);
nand UO_1937 (O_1937,N_19983,N_19928);
xnor UO_1938 (O_1938,N_19937,N_19853);
and UO_1939 (O_1939,N_19933,N_19937);
xnor UO_1940 (O_1940,N_19969,N_19844);
nor UO_1941 (O_1941,N_19802,N_19972);
and UO_1942 (O_1942,N_19948,N_19941);
xor UO_1943 (O_1943,N_19964,N_19885);
and UO_1944 (O_1944,N_19844,N_19968);
or UO_1945 (O_1945,N_19811,N_19866);
nand UO_1946 (O_1946,N_19825,N_19915);
xnor UO_1947 (O_1947,N_19995,N_19898);
and UO_1948 (O_1948,N_19949,N_19900);
xnor UO_1949 (O_1949,N_19906,N_19990);
xnor UO_1950 (O_1950,N_19847,N_19854);
or UO_1951 (O_1951,N_19852,N_19951);
and UO_1952 (O_1952,N_19817,N_19875);
nor UO_1953 (O_1953,N_19989,N_19950);
nand UO_1954 (O_1954,N_19918,N_19891);
or UO_1955 (O_1955,N_19834,N_19958);
and UO_1956 (O_1956,N_19813,N_19957);
nand UO_1957 (O_1957,N_19895,N_19915);
and UO_1958 (O_1958,N_19860,N_19876);
xnor UO_1959 (O_1959,N_19933,N_19999);
xor UO_1960 (O_1960,N_19981,N_19992);
or UO_1961 (O_1961,N_19846,N_19831);
nand UO_1962 (O_1962,N_19968,N_19875);
nand UO_1963 (O_1963,N_19980,N_19869);
nand UO_1964 (O_1964,N_19952,N_19891);
nor UO_1965 (O_1965,N_19964,N_19912);
xnor UO_1966 (O_1966,N_19975,N_19864);
and UO_1967 (O_1967,N_19975,N_19961);
and UO_1968 (O_1968,N_19929,N_19873);
nand UO_1969 (O_1969,N_19968,N_19969);
nand UO_1970 (O_1970,N_19950,N_19956);
xnor UO_1971 (O_1971,N_19839,N_19817);
xnor UO_1972 (O_1972,N_19915,N_19832);
or UO_1973 (O_1973,N_19819,N_19940);
nand UO_1974 (O_1974,N_19822,N_19927);
nor UO_1975 (O_1975,N_19932,N_19899);
xnor UO_1976 (O_1976,N_19876,N_19925);
nand UO_1977 (O_1977,N_19892,N_19970);
nor UO_1978 (O_1978,N_19869,N_19981);
or UO_1979 (O_1979,N_19852,N_19900);
nand UO_1980 (O_1980,N_19966,N_19819);
nor UO_1981 (O_1981,N_19815,N_19903);
nand UO_1982 (O_1982,N_19969,N_19919);
nor UO_1983 (O_1983,N_19836,N_19875);
xor UO_1984 (O_1984,N_19977,N_19933);
nand UO_1985 (O_1985,N_19949,N_19958);
nor UO_1986 (O_1986,N_19835,N_19869);
nand UO_1987 (O_1987,N_19868,N_19957);
and UO_1988 (O_1988,N_19804,N_19999);
and UO_1989 (O_1989,N_19834,N_19915);
or UO_1990 (O_1990,N_19922,N_19823);
and UO_1991 (O_1991,N_19960,N_19980);
nand UO_1992 (O_1992,N_19969,N_19814);
nor UO_1993 (O_1993,N_19865,N_19830);
xor UO_1994 (O_1994,N_19821,N_19856);
or UO_1995 (O_1995,N_19851,N_19900);
or UO_1996 (O_1996,N_19983,N_19929);
or UO_1997 (O_1997,N_19917,N_19998);
or UO_1998 (O_1998,N_19997,N_19803);
xnor UO_1999 (O_1999,N_19997,N_19837);
or UO_2000 (O_2000,N_19839,N_19981);
xnor UO_2001 (O_2001,N_19809,N_19896);
xnor UO_2002 (O_2002,N_19855,N_19834);
xnor UO_2003 (O_2003,N_19879,N_19878);
or UO_2004 (O_2004,N_19892,N_19997);
nand UO_2005 (O_2005,N_19886,N_19841);
or UO_2006 (O_2006,N_19978,N_19924);
and UO_2007 (O_2007,N_19809,N_19969);
and UO_2008 (O_2008,N_19838,N_19877);
xnor UO_2009 (O_2009,N_19861,N_19838);
and UO_2010 (O_2010,N_19933,N_19852);
xnor UO_2011 (O_2011,N_19914,N_19875);
and UO_2012 (O_2012,N_19956,N_19858);
xor UO_2013 (O_2013,N_19884,N_19940);
and UO_2014 (O_2014,N_19952,N_19994);
or UO_2015 (O_2015,N_19982,N_19994);
nor UO_2016 (O_2016,N_19812,N_19822);
nor UO_2017 (O_2017,N_19919,N_19899);
nand UO_2018 (O_2018,N_19860,N_19963);
and UO_2019 (O_2019,N_19864,N_19868);
nand UO_2020 (O_2020,N_19969,N_19893);
or UO_2021 (O_2021,N_19935,N_19998);
xnor UO_2022 (O_2022,N_19948,N_19801);
xnor UO_2023 (O_2023,N_19858,N_19840);
and UO_2024 (O_2024,N_19925,N_19831);
or UO_2025 (O_2025,N_19920,N_19958);
and UO_2026 (O_2026,N_19943,N_19983);
nand UO_2027 (O_2027,N_19819,N_19814);
or UO_2028 (O_2028,N_19873,N_19951);
and UO_2029 (O_2029,N_19987,N_19810);
nand UO_2030 (O_2030,N_19873,N_19801);
or UO_2031 (O_2031,N_19971,N_19887);
and UO_2032 (O_2032,N_19866,N_19919);
nand UO_2033 (O_2033,N_19829,N_19928);
or UO_2034 (O_2034,N_19986,N_19903);
xnor UO_2035 (O_2035,N_19903,N_19847);
nor UO_2036 (O_2036,N_19828,N_19810);
and UO_2037 (O_2037,N_19869,N_19943);
nor UO_2038 (O_2038,N_19900,N_19836);
nor UO_2039 (O_2039,N_19879,N_19809);
and UO_2040 (O_2040,N_19909,N_19924);
nor UO_2041 (O_2041,N_19808,N_19999);
or UO_2042 (O_2042,N_19802,N_19861);
and UO_2043 (O_2043,N_19838,N_19977);
xor UO_2044 (O_2044,N_19963,N_19942);
nand UO_2045 (O_2045,N_19996,N_19991);
nor UO_2046 (O_2046,N_19951,N_19857);
nor UO_2047 (O_2047,N_19961,N_19866);
nor UO_2048 (O_2048,N_19965,N_19986);
and UO_2049 (O_2049,N_19850,N_19855);
xnor UO_2050 (O_2050,N_19919,N_19881);
or UO_2051 (O_2051,N_19951,N_19914);
or UO_2052 (O_2052,N_19835,N_19930);
or UO_2053 (O_2053,N_19900,N_19880);
or UO_2054 (O_2054,N_19817,N_19823);
nand UO_2055 (O_2055,N_19871,N_19914);
nor UO_2056 (O_2056,N_19949,N_19803);
and UO_2057 (O_2057,N_19998,N_19883);
nand UO_2058 (O_2058,N_19993,N_19866);
and UO_2059 (O_2059,N_19910,N_19872);
and UO_2060 (O_2060,N_19807,N_19910);
or UO_2061 (O_2061,N_19953,N_19858);
and UO_2062 (O_2062,N_19912,N_19954);
or UO_2063 (O_2063,N_19925,N_19863);
xnor UO_2064 (O_2064,N_19991,N_19929);
xor UO_2065 (O_2065,N_19902,N_19841);
and UO_2066 (O_2066,N_19962,N_19924);
nor UO_2067 (O_2067,N_19991,N_19979);
nor UO_2068 (O_2068,N_19882,N_19816);
xnor UO_2069 (O_2069,N_19999,N_19915);
nor UO_2070 (O_2070,N_19956,N_19871);
nor UO_2071 (O_2071,N_19984,N_19890);
nor UO_2072 (O_2072,N_19867,N_19969);
nor UO_2073 (O_2073,N_19997,N_19903);
xor UO_2074 (O_2074,N_19921,N_19816);
xnor UO_2075 (O_2075,N_19999,N_19932);
nor UO_2076 (O_2076,N_19821,N_19885);
or UO_2077 (O_2077,N_19898,N_19937);
or UO_2078 (O_2078,N_19987,N_19974);
or UO_2079 (O_2079,N_19977,N_19853);
nand UO_2080 (O_2080,N_19875,N_19888);
nor UO_2081 (O_2081,N_19953,N_19808);
xor UO_2082 (O_2082,N_19803,N_19811);
nand UO_2083 (O_2083,N_19873,N_19833);
and UO_2084 (O_2084,N_19969,N_19997);
nand UO_2085 (O_2085,N_19967,N_19820);
and UO_2086 (O_2086,N_19874,N_19903);
nor UO_2087 (O_2087,N_19875,N_19847);
and UO_2088 (O_2088,N_19861,N_19854);
and UO_2089 (O_2089,N_19949,N_19848);
nand UO_2090 (O_2090,N_19845,N_19975);
xor UO_2091 (O_2091,N_19839,N_19937);
nor UO_2092 (O_2092,N_19873,N_19812);
or UO_2093 (O_2093,N_19991,N_19926);
xor UO_2094 (O_2094,N_19999,N_19953);
xnor UO_2095 (O_2095,N_19945,N_19979);
and UO_2096 (O_2096,N_19934,N_19894);
nand UO_2097 (O_2097,N_19942,N_19929);
xnor UO_2098 (O_2098,N_19975,N_19992);
nand UO_2099 (O_2099,N_19999,N_19942);
or UO_2100 (O_2100,N_19847,N_19987);
or UO_2101 (O_2101,N_19976,N_19917);
and UO_2102 (O_2102,N_19940,N_19890);
and UO_2103 (O_2103,N_19847,N_19938);
xnor UO_2104 (O_2104,N_19945,N_19873);
and UO_2105 (O_2105,N_19810,N_19836);
nor UO_2106 (O_2106,N_19981,N_19966);
nand UO_2107 (O_2107,N_19998,N_19938);
or UO_2108 (O_2108,N_19951,N_19910);
xnor UO_2109 (O_2109,N_19889,N_19980);
nand UO_2110 (O_2110,N_19996,N_19867);
and UO_2111 (O_2111,N_19823,N_19901);
nand UO_2112 (O_2112,N_19800,N_19808);
nor UO_2113 (O_2113,N_19892,N_19812);
xnor UO_2114 (O_2114,N_19839,N_19823);
and UO_2115 (O_2115,N_19868,N_19840);
and UO_2116 (O_2116,N_19827,N_19997);
nand UO_2117 (O_2117,N_19976,N_19839);
or UO_2118 (O_2118,N_19843,N_19890);
and UO_2119 (O_2119,N_19890,N_19977);
nand UO_2120 (O_2120,N_19946,N_19898);
xor UO_2121 (O_2121,N_19851,N_19861);
nand UO_2122 (O_2122,N_19993,N_19864);
xor UO_2123 (O_2123,N_19980,N_19838);
nand UO_2124 (O_2124,N_19830,N_19827);
and UO_2125 (O_2125,N_19810,N_19994);
nand UO_2126 (O_2126,N_19936,N_19913);
or UO_2127 (O_2127,N_19924,N_19919);
nand UO_2128 (O_2128,N_19961,N_19952);
nor UO_2129 (O_2129,N_19862,N_19811);
nand UO_2130 (O_2130,N_19830,N_19993);
and UO_2131 (O_2131,N_19890,N_19833);
nor UO_2132 (O_2132,N_19849,N_19871);
or UO_2133 (O_2133,N_19995,N_19886);
nand UO_2134 (O_2134,N_19906,N_19953);
nand UO_2135 (O_2135,N_19959,N_19881);
or UO_2136 (O_2136,N_19850,N_19940);
nand UO_2137 (O_2137,N_19859,N_19952);
or UO_2138 (O_2138,N_19813,N_19888);
nand UO_2139 (O_2139,N_19936,N_19987);
and UO_2140 (O_2140,N_19912,N_19939);
nand UO_2141 (O_2141,N_19966,N_19911);
and UO_2142 (O_2142,N_19851,N_19858);
and UO_2143 (O_2143,N_19971,N_19826);
nand UO_2144 (O_2144,N_19855,N_19897);
nand UO_2145 (O_2145,N_19975,N_19826);
xnor UO_2146 (O_2146,N_19807,N_19950);
and UO_2147 (O_2147,N_19985,N_19940);
or UO_2148 (O_2148,N_19986,N_19946);
xor UO_2149 (O_2149,N_19906,N_19946);
nor UO_2150 (O_2150,N_19806,N_19807);
nor UO_2151 (O_2151,N_19949,N_19941);
xor UO_2152 (O_2152,N_19960,N_19907);
nor UO_2153 (O_2153,N_19854,N_19891);
xnor UO_2154 (O_2154,N_19815,N_19900);
or UO_2155 (O_2155,N_19934,N_19989);
nor UO_2156 (O_2156,N_19828,N_19914);
or UO_2157 (O_2157,N_19833,N_19851);
xor UO_2158 (O_2158,N_19937,N_19989);
nand UO_2159 (O_2159,N_19953,N_19907);
nand UO_2160 (O_2160,N_19997,N_19981);
xor UO_2161 (O_2161,N_19973,N_19891);
or UO_2162 (O_2162,N_19943,N_19932);
xor UO_2163 (O_2163,N_19884,N_19879);
nand UO_2164 (O_2164,N_19892,N_19862);
nand UO_2165 (O_2165,N_19948,N_19925);
nand UO_2166 (O_2166,N_19981,N_19807);
or UO_2167 (O_2167,N_19898,N_19940);
or UO_2168 (O_2168,N_19868,N_19935);
and UO_2169 (O_2169,N_19819,N_19888);
nand UO_2170 (O_2170,N_19800,N_19855);
and UO_2171 (O_2171,N_19984,N_19842);
or UO_2172 (O_2172,N_19854,N_19852);
xnor UO_2173 (O_2173,N_19864,N_19961);
or UO_2174 (O_2174,N_19961,N_19861);
nand UO_2175 (O_2175,N_19896,N_19865);
and UO_2176 (O_2176,N_19826,N_19807);
nor UO_2177 (O_2177,N_19981,N_19857);
nor UO_2178 (O_2178,N_19864,N_19941);
or UO_2179 (O_2179,N_19995,N_19986);
nor UO_2180 (O_2180,N_19972,N_19836);
nand UO_2181 (O_2181,N_19846,N_19946);
and UO_2182 (O_2182,N_19908,N_19952);
nor UO_2183 (O_2183,N_19997,N_19983);
nand UO_2184 (O_2184,N_19981,N_19888);
nor UO_2185 (O_2185,N_19904,N_19915);
xnor UO_2186 (O_2186,N_19955,N_19942);
or UO_2187 (O_2187,N_19978,N_19981);
nand UO_2188 (O_2188,N_19903,N_19912);
and UO_2189 (O_2189,N_19892,N_19840);
and UO_2190 (O_2190,N_19918,N_19859);
nor UO_2191 (O_2191,N_19910,N_19964);
and UO_2192 (O_2192,N_19963,N_19858);
and UO_2193 (O_2193,N_19995,N_19853);
and UO_2194 (O_2194,N_19861,N_19963);
and UO_2195 (O_2195,N_19994,N_19858);
nor UO_2196 (O_2196,N_19900,N_19849);
nand UO_2197 (O_2197,N_19963,N_19817);
xnor UO_2198 (O_2198,N_19816,N_19963);
or UO_2199 (O_2199,N_19978,N_19898);
nand UO_2200 (O_2200,N_19836,N_19908);
xnor UO_2201 (O_2201,N_19970,N_19961);
nor UO_2202 (O_2202,N_19980,N_19834);
and UO_2203 (O_2203,N_19865,N_19888);
xnor UO_2204 (O_2204,N_19807,N_19866);
xnor UO_2205 (O_2205,N_19899,N_19815);
nand UO_2206 (O_2206,N_19993,N_19933);
nor UO_2207 (O_2207,N_19873,N_19868);
xnor UO_2208 (O_2208,N_19867,N_19900);
nand UO_2209 (O_2209,N_19920,N_19943);
or UO_2210 (O_2210,N_19944,N_19901);
or UO_2211 (O_2211,N_19856,N_19961);
or UO_2212 (O_2212,N_19849,N_19877);
nand UO_2213 (O_2213,N_19976,N_19900);
or UO_2214 (O_2214,N_19914,N_19860);
and UO_2215 (O_2215,N_19858,N_19973);
nand UO_2216 (O_2216,N_19889,N_19923);
and UO_2217 (O_2217,N_19848,N_19807);
nor UO_2218 (O_2218,N_19809,N_19965);
xnor UO_2219 (O_2219,N_19927,N_19995);
nand UO_2220 (O_2220,N_19827,N_19834);
and UO_2221 (O_2221,N_19902,N_19812);
nand UO_2222 (O_2222,N_19870,N_19823);
or UO_2223 (O_2223,N_19868,N_19902);
xor UO_2224 (O_2224,N_19917,N_19813);
nand UO_2225 (O_2225,N_19982,N_19980);
nand UO_2226 (O_2226,N_19966,N_19951);
xnor UO_2227 (O_2227,N_19861,N_19864);
nand UO_2228 (O_2228,N_19838,N_19802);
or UO_2229 (O_2229,N_19868,N_19886);
nand UO_2230 (O_2230,N_19944,N_19941);
nand UO_2231 (O_2231,N_19967,N_19806);
nor UO_2232 (O_2232,N_19827,N_19902);
nor UO_2233 (O_2233,N_19830,N_19868);
nand UO_2234 (O_2234,N_19905,N_19829);
xnor UO_2235 (O_2235,N_19829,N_19872);
or UO_2236 (O_2236,N_19921,N_19932);
nand UO_2237 (O_2237,N_19844,N_19930);
or UO_2238 (O_2238,N_19895,N_19952);
xor UO_2239 (O_2239,N_19955,N_19825);
xnor UO_2240 (O_2240,N_19987,N_19843);
nand UO_2241 (O_2241,N_19914,N_19814);
xnor UO_2242 (O_2242,N_19885,N_19858);
and UO_2243 (O_2243,N_19903,N_19845);
and UO_2244 (O_2244,N_19979,N_19922);
nand UO_2245 (O_2245,N_19856,N_19970);
xnor UO_2246 (O_2246,N_19847,N_19885);
nor UO_2247 (O_2247,N_19907,N_19946);
xor UO_2248 (O_2248,N_19814,N_19894);
and UO_2249 (O_2249,N_19917,N_19861);
or UO_2250 (O_2250,N_19815,N_19901);
nand UO_2251 (O_2251,N_19824,N_19830);
and UO_2252 (O_2252,N_19805,N_19842);
nand UO_2253 (O_2253,N_19860,N_19847);
xor UO_2254 (O_2254,N_19847,N_19870);
and UO_2255 (O_2255,N_19883,N_19820);
xnor UO_2256 (O_2256,N_19952,N_19902);
xnor UO_2257 (O_2257,N_19840,N_19935);
nand UO_2258 (O_2258,N_19896,N_19949);
nand UO_2259 (O_2259,N_19889,N_19964);
xnor UO_2260 (O_2260,N_19845,N_19846);
or UO_2261 (O_2261,N_19821,N_19822);
or UO_2262 (O_2262,N_19824,N_19874);
nor UO_2263 (O_2263,N_19939,N_19911);
or UO_2264 (O_2264,N_19974,N_19836);
and UO_2265 (O_2265,N_19924,N_19936);
nor UO_2266 (O_2266,N_19875,N_19971);
nand UO_2267 (O_2267,N_19915,N_19864);
xnor UO_2268 (O_2268,N_19963,N_19848);
nand UO_2269 (O_2269,N_19899,N_19961);
or UO_2270 (O_2270,N_19950,N_19958);
or UO_2271 (O_2271,N_19831,N_19954);
or UO_2272 (O_2272,N_19954,N_19891);
nand UO_2273 (O_2273,N_19981,N_19811);
and UO_2274 (O_2274,N_19994,N_19964);
nor UO_2275 (O_2275,N_19995,N_19996);
and UO_2276 (O_2276,N_19877,N_19859);
nand UO_2277 (O_2277,N_19858,N_19861);
nor UO_2278 (O_2278,N_19942,N_19946);
nor UO_2279 (O_2279,N_19841,N_19843);
nand UO_2280 (O_2280,N_19813,N_19834);
or UO_2281 (O_2281,N_19890,N_19870);
nor UO_2282 (O_2282,N_19929,N_19998);
nor UO_2283 (O_2283,N_19839,N_19996);
and UO_2284 (O_2284,N_19940,N_19835);
nand UO_2285 (O_2285,N_19885,N_19911);
xor UO_2286 (O_2286,N_19900,N_19803);
or UO_2287 (O_2287,N_19997,N_19878);
nand UO_2288 (O_2288,N_19854,N_19836);
xor UO_2289 (O_2289,N_19929,N_19947);
nor UO_2290 (O_2290,N_19808,N_19839);
nand UO_2291 (O_2291,N_19991,N_19888);
xor UO_2292 (O_2292,N_19968,N_19956);
nand UO_2293 (O_2293,N_19897,N_19884);
and UO_2294 (O_2294,N_19941,N_19981);
nor UO_2295 (O_2295,N_19981,N_19813);
xor UO_2296 (O_2296,N_19966,N_19842);
nand UO_2297 (O_2297,N_19999,N_19986);
or UO_2298 (O_2298,N_19954,N_19848);
xor UO_2299 (O_2299,N_19921,N_19912);
or UO_2300 (O_2300,N_19928,N_19897);
or UO_2301 (O_2301,N_19959,N_19815);
nor UO_2302 (O_2302,N_19836,N_19930);
or UO_2303 (O_2303,N_19872,N_19981);
and UO_2304 (O_2304,N_19908,N_19922);
xor UO_2305 (O_2305,N_19908,N_19875);
and UO_2306 (O_2306,N_19882,N_19888);
xor UO_2307 (O_2307,N_19806,N_19801);
xnor UO_2308 (O_2308,N_19979,N_19932);
xnor UO_2309 (O_2309,N_19893,N_19890);
nor UO_2310 (O_2310,N_19833,N_19841);
or UO_2311 (O_2311,N_19894,N_19942);
xor UO_2312 (O_2312,N_19999,N_19861);
nor UO_2313 (O_2313,N_19973,N_19837);
and UO_2314 (O_2314,N_19809,N_19925);
or UO_2315 (O_2315,N_19851,N_19803);
nand UO_2316 (O_2316,N_19888,N_19809);
xor UO_2317 (O_2317,N_19868,N_19973);
or UO_2318 (O_2318,N_19991,N_19987);
nand UO_2319 (O_2319,N_19875,N_19913);
xnor UO_2320 (O_2320,N_19858,N_19826);
nor UO_2321 (O_2321,N_19906,N_19950);
or UO_2322 (O_2322,N_19897,N_19800);
or UO_2323 (O_2323,N_19938,N_19994);
nor UO_2324 (O_2324,N_19863,N_19928);
or UO_2325 (O_2325,N_19946,N_19966);
and UO_2326 (O_2326,N_19978,N_19904);
nor UO_2327 (O_2327,N_19916,N_19824);
nand UO_2328 (O_2328,N_19828,N_19986);
nand UO_2329 (O_2329,N_19800,N_19978);
and UO_2330 (O_2330,N_19960,N_19958);
and UO_2331 (O_2331,N_19991,N_19923);
nor UO_2332 (O_2332,N_19877,N_19844);
xor UO_2333 (O_2333,N_19946,N_19880);
nand UO_2334 (O_2334,N_19895,N_19905);
nor UO_2335 (O_2335,N_19843,N_19808);
and UO_2336 (O_2336,N_19997,N_19835);
nor UO_2337 (O_2337,N_19933,N_19936);
or UO_2338 (O_2338,N_19920,N_19861);
xor UO_2339 (O_2339,N_19996,N_19966);
nor UO_2340 (O_2340,N_19872,N_19985);
nor UO_2341 (O_2341,N_19857,N_19881);
or UO_2342 (O_2342,N_19875,N_19898);
nand UO_2343 (O_2343,N_19987,N_19891);
nand UO_2344 (O_2344,N_19982,N_19997);
xnor UO_2345 (O_2345,N_19807,N_19867);
xnor UO_2346 (O_2346,N_19959,N_19875);
or UO_2347 (O_2347,N_19894,N_19819);
and UO_2348 (O_2348,N_19868,N_19981);
and UO_2349 (O_2349,N_19925,N_19987);
xor UO_2350 (O_2350,N_19842,N_19917);
xnor UO_2351 (O_2351,N_19801,N_19998);
nand UO_2352 (O_2352,N_19880,N_19997);
and UO_2353 (O_2353,N_19969,N_19875);
nand UO_2354 (O_2354,N_19814,N_19950);
and UO_2355 (O_2355,N_19854,N_19809);
or UO_2356 (O_2356,N_19889,N_19957);
nor UO_2357 (O_2357,N_19863,N_19944);
xor UO_2358 (O_2358,N_19913,N_19881);
or UO_2359 (O_2359,N_19961,N_19917);
nand UO_2360 (O_2360,N_19823,N_19940);
nor UO_2361 (O_2361,N_19952,N_19941);
nand UO_2362 (O_2362,N_19882,N_19820);
nand UO_2363 (O_2363,N_19832,N_19983);
nand UO_2364 (O_2364,N_19838,N_19962);
nor UO_2365 (O_2365,N_19830,N_19974);
xor UO_2366 (O_2366,N_19953,N_19828);
nand UO_2367 (O_2367,N_19874,N_19915);
or UO_2368 (O_2368,N_19856,N_19973);
nor UO_2369 (O_2369,N_19952,N_19820);
nand UO_2370 (O_2370,N_19911,N_19822);
and UO_2371 (O_2371,N_19822,N_19942);
nor UO_2372 (O_2372,N_19925,N_19944);
and UO_2373 (O_2373,N_19982,N_19898);
and UO_2374 (O_2374,N_19988,N_19997);
xnor UO_2375 (O_2375,N_19852,N_19823);
xor UO_2376 (O_2376,N_19883,N_19806);
nor UO_2377 (O_2377,N_19840,N_19896);
nor UO_2378 (O_2378,N_19844,N_19909);
nand UO_2379 (O_2379,N_19978,N_19903);
nand UO_2380 (O_2380,N_19867,N_19811);
and UO_2381 (O_2381,N_19800,N_19875);
nor UO_2382 (O_2382,N_19845,N_19835);
nor UO_2383 (O_2383,N_19812,N_19981);
and UO_2384 (O_2384,N_19981,N_19995);
xnor UO_2385 (O_2385,N_19878,N_19952);
nand UO_2386 (O_2386,N_19909,N_19869);
or UO_2387 (O_2387,N_19812,N_19865);
and UO_2388 (O_2388,N_19892,N_19802);
nor UO_2389 (O_2389,N_19936,N_19895);
or UO_2390 (O_2390,N_19980,N_19966);
xor UO_2391 (O_2391,N_19859,N_19917);
or UO_2392 (O_2392,N_19851,N_19862);
nor UO_2393 (O_2393,N_19952,N_19996);
nor UO_2394 (O_2394,N_19865,N_19881);
or UO_2395 (O_2395,N_19924,N_19986);
nand UO_2396 (O_2396,N_19839,N_19904);
xnor UO_2397 (O_2397,N_19858,N_19822);
nand UO_2398 (O_2398,N_19826,N_19930);
or UO_2399 (O_2399,N_19843,N_19906);
nor UO_2400 (O_2400,N_19857,N_19875);
xor UO_2401 (O_2401,N_19836,N_19892);
xor UO_2402 (O_2402,N_19939,N_19953);
or UO_2403 (O_2403,N_19809,N_19820);
or UO_2404 (O_2404,N_19994,N_19909);
or UO_2405 (O_2405,N_19880,N_19895);
xor UO_2406 (O_2406,N_19981,N_19953);
and UO_2407 (O_2407,N_19950,N_19901);
xnor UO_2408 (O_2408,N_19869,N_19942);
and UO_2409 (O_2409,N_19946,N_19958);
nand UO_2410 (O_2410,N_19989,N_19930);
nor UO_2411 (O_2411,N_19971,N_19888);
nor UO_2412 (O_2412,N_19913,N_19801);
or UO_2413 (O_2413,N_19892,N_19910);
nand UO_2414 (O_2414,N_19953,N_19968);
and UO_2415 (O_2415,N_19852,N_19914);
and UO_2416 (O_2416,N_19815,N_19908);
nand UO_2417 (O_2417,N_19808,N_19900);
nor UO_2418 (O_2418,N_19922,N_19854);
or UO_2419 (O_2419,N_19891,N_19979);
and UO_2420 (O_2420,N_19864,N_19870);
xor UO_2421 (O_2421,N_19942,N_19845);
nand UO_2422 (O_2422,N_19804,N_19982);
xnor UO_2423 (O_2423,N_19820,N_19991);
or UO_2424 (O_2424,N_19821,N_19857);
or UO_2425 (O_2425,N_19957,N_19926);
xnor UO_2426 (O_2426,N_19811,N_19958);
xor UO_2427 (O_2427,N_19820,N_19851);
nand UO_2428 (O_2428,N_19946,N_19866);
xnor UO_2429 (O_2429,N_19978,N_19819);
and UO_2430 (O_2430,N_19902,N_19857);
xor UO_2431 (O_2431,N_19955,N_19938);
nor UO_2432 (O_2432,N_19828,N_19907);
and UO_2433 (O_2433,N_19878,N_19844);
and UO_2434 (O_2434,N_19926,N_19830);
and UO_2435 (O_2435,N_19884,N_19870);
nor UO_2436 (O_2436,N_19870,N_19946);
nor UO_2437 (O_2437,N_19930,N_19893);
or UO_2438 (O_2438,N_19804,N_19882);
and UO_2439 (O_2439,N_19961,N_19947);
nor UO_2440 (O_2440,N_19818,N_19906);
and UO_2441 (O_2441,N_19987,N_19854);
nor UO_2442 (O_2442,N_19954,N_19800);
nand UO_2443 (O_2443,N_19883,N_19916);
nand UO_2444 (O_2444,N_19838,N_19879);
or UO_2445 (O_2445,N_19810,N_19956);
xor UO_2446 (O_2446,N_19949,N_19999);
nor UO_2447 (O_2447,N_19969,N_19931);
and UO_2448 (O_2448,N_19853,N_19819);
or UO_2449 (O_2449,N_19811,N_19997);
nand UO_2450 (O_2450,N_19973,N_19849);
nor UO_2451 (O_2451,N_19951,N_19805);
and UO_2452 (O_2452,N_19845,N_19910);
nand UO_2453 (O_2453,N_19982,N_19888);
and UO_2454 (O_2454,N_19963,N_19997);
and UO_2455 (O_2455,N_19961,N_19875);
and UO_2456 (O_2456,N_19861,N_19806);
nand UO_2457 (O_2457,N_19898,N_19899);
and UO_2458 (O_2458,N_19985,N_19884);
nor UO_2459 (O_2459,N_19853,N_19881);
nand UO_2460 (O_2460,N_19988,N_19856);
and UO_2461 (O_2461,N_19895,N_19879);
nor UO_2462 (O_2462,N_19954,N_19938);
nor UO_2463 (O_2463,N_19958,N_19876);
xor UO_2464 (O_2464,N_19878,N_19873);
or UO_2465 (O_2465,N_19921,N_19999);
xnor UO_2466 (O_2466,N_19831,N_19833);
or UO_2467 (O_2467,N_19900,N_19864);
xnor UO_2468 (O_2468,N_19997,N_19939);
or UO_2469 (O_2469,N_19939,N_19844);
nor UO_2470 (O_2470,N_19908,N_19916);
nand UO_2471 (O_2471,N_19851,N_19928);
xnor UO_2472 (O_2472,N_19981,N_19903);
nor UO_2473 (O_2473,N_19949,N_19844);
nor UO_2474 (O_2474,N_19969,N_19925);
or UO_2475 (O_2475,N_19887,N_19827);
nor UO_2476 (O_2476,N_19923,N_19943);
nor UO_2477 (O_2477,N_19862,N_19931);
xor UO_2478 (O_2478,N_19981,N_19920);
or UO_2479 (O_2479,N_19892,N_19813);
or UO_2480 (O_2480,N_19892,N_19917);
xnor UO_2481 (O_2481,N_19942,N_19970);
nand UO_2482 (O_2482,N_19831,N_19802);
and UO_2483 (O_2483,N_19916,N_19917);
or UO_2484 (O_2484,N_19948,N_19897);
xor UO_2485 (O_2485,N_19972,N_19874);
nand UO_2486 (O_2486,N_19883,N_19888);
xnor UO_2487 (O_2487,N_19833,N_19901);
and UO_2488 (O_2488,N_19938,N_19821);
and UO_2489 (O_2489,N_19992,N_19874);
nor UO_2490 (O_2490,N_19854,N_19802);
xor UO_2491 (O_2491,N_19884,N_19979);
xnor UO_2492 (O_2492,N_19984,N_19847);
nand UO_2493 (O_2493,N_19964,N_19962);
nand UO_2494 (O_2494,N_19889,N_19977);
and UO_2495 (O_2495,N_19969,N_19952);
nand UO_2496 (O_2496,N_19885,N_19923);
xor UO_2497 (O_2497,N_19988,N_19945);
and UO_2498 (O_2498,N_19830,N_19943);
xor UO_2499 (O_2499,N_19968,N_19928);
endmodule