module basic_3000_30000_3500_50_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1860,In_589);
nand U1 (N_1,In_1944,In_183);
or U2 (N_2,In_149,In_687);
nand U3 (N_3,In_2531,In_2748);
nand U4 (N_4,In_2632,In_838);
nand U5 (N_5,In_1466,In_2651);
and U6 (N_6,In_264,In_213);
nand U7 (N_7,In_1877,In_26);
and U8 (N_8,In_787,In_2679);
nor U9 (N_9,In_2298,In_2764);
nand U10 (N_10,In_1300,In_744);
nand U11 (N_11,In_1534,In_963);
or U12 (N_12,In_1372,In_386);
or U13 (N_13,In_1796,In_2424);
nand U14 (N_14,In_2201,In_2143);
nand U15 (N_15,In_221,In_627);
nand U16 (N_16,In_558,In_749);
and U17 (N_17,In_2714,In_2304);
nor U18 (N_18,In_2879,In_128);
and U19 (N_19,In_2561,In_1406);
nor U20 (N_20,In_2930,In_648);
and U21 (N_21,In_679,In_1618);
and U22 (N_22,In_174,In_62);
nand U23 (N_23,In_241,In_847);
nand U24 (N_24,In_1768,In_1553);
or U25 (N_25,In_311,In_1779);
nor U26 (N_26,In_2546,In_693);
and U27 (N_27,In_730,In_309);
nand U28 (N_28,In_1644,In_1211);
and U29 (N_29,In_813,In_307);
or U30 (N_30,In_2245,In_2408);
and U31 (N_31,In_1705,In_160);
nor U32 (N_32,In_224,In_2630);
nand U33 (N_33,In_837,In_1809);
or U34 (N_34,In_372,In_1351);
nand U35 (N_35,In_962,In_1836);
xor U36 (N_36,In_2653,In_1449);
nand U37 (N_37,In_1452,In_115);
nor U38 (N_38,In_315,In_907);
or U39 (N_39,In_2309,In_1682);
and U40 (N_40,In_529,In_185);
or U41 (N_41,In_1100,In_2157);
nand U42 (N_42,In_105,In_812);
nand U43 (N_43,In_1925,In_112);
or U44 (N_44,In_2988,In_1309);
nor U45 (N_45,In_1482,In_596);
and U46 (N_46,In_205,In_1681);
and U47 (N_47,In_1435,In_2732);
and U48 (N_48,In_1942,In_2367);
and U49 (N_49,In_2027,In_1379);
nor U50 (N_50,In_2968,In_740);
nand U51 (N_51,In_1824,In_1600);
or U52 (N_52,In_2737,In_1933);
and U53 (N_53,In_1993,In_152);
or U54 (N_54,In_2292,In_2490);
nor U55 (N_55,In_1310,In_755);
or U56 (N_56,In_464,In_1488);
or U57 (N_57,In_1914,In_2513);
or U58 (N_58,In_762,In_2856);
and U59 (N_59,In_1967,In_2606);
and U60 (N_60,In_2072,In_2729);
or U61 (N_61,In_1661,In_2962);
and U62 (N_62,In_564,In_91);
nand U63 (N_63,In_2542,In_1880);
nand U64 (N_64,In_2413,In_1072);
and U65 (N_65,In_108,In_2938);
or U66 (N_66,In_2358,In_652);
nor U67 (N_67,In_1783,In_1612);
nor U68 (N_68,In_2660,In_2277);
or U69 (N_69,In_1471,In_119);
nor U70 (N_70,In_236,In_737);
or U71 (N_71,In_1380,In_2381);
nor U72 (N_72,In_1569,In_598);
and U73 (N_73,In_2465,In_293);
nand U74 (N_74,In_2836,In_1142);
nor U75 (N_75,In_2011,In_2921);
nor U76 (N_76,In_342,In_2070);
and U77 (N_77,In_1749,In_535);
nand U78 (N_78,In_1823,In_1523);
nand U79 (N_79,In_828,In_1637);
and U80 (N_80,In_1075,In_921);
and U81 (N_81,In_654,In_2472);
and U82 (N_82,In_491,In_2004);
nor U83 (N_83,In_1619,In_1392);
nand U84 (N_84,In_69,In_42);
or U85 (N_85,In_839,In_2569);
or U86 (N_86,In_521,In_2347);
nor U87 (N_87,In_2956,In_417);
and U88 (N_88,In_1187,In_912);
nor U89 (N_89,In_1598,In_1725);
nand U90 (N_90,In_429,In_18);
or U91 (N_91,In_822,In_1089);
nand U92 (N_92,In_52,In_520);
nand U93 (N_93,In_951,In_93);
nand U94 (N_94,In_759,In_2012);
nand U95 (N_95,In_2395,In_436);
or U96 (N_96,In_312,In_2698);
nand U97 (N_97,In_2948,In_1795);
and U98 (N_98,In_180,In_1848);
or U99 (N_99,In_1256,In_30);
or U100 (N_100,In_1630,In_639);
or U101 (N_101,In_156,In_2843);
or U102 (N_102,In_2604,In_1722);
nand U103 (N_103,In_1601,In_2855);
nand U104 (N_104,In_1786,In_741);
nand U105 (N_105,In_78,In_1259);
and U106 (N_106,In_120,In_1891);
nand U107 (N_107,In_1108,In_2433);
or U108 (N_108,In_2686,In_1893);
nor U109 (N_109,In_339,In_2094);
nand U110 (N_110,In_2754,In_2863);
nor U111 (N_111,In_1053,In_1235);
nor U112 (N_112,In_1752,In_1260);
nor U113 (N_113,In_1456,In_1789);
nand U114 (N_114,In_1447,In_2107);
xnor U115 (N_115,In_2726,In_118);
or U116 (N_116,In_2873,In_384);
xnor U117 (N_117,In_1057,In_405);
nor U118 (N_118,In_1778,In_1551);
or U119 (N_119,In_1912,In_1158);
nand U120 (N_120,In_277,In_2017);
nor U121 (N_121,In_956,In_2940);
nor U122 (N_122,In_355,In_1923);
nand U123 (N_123,In_2915,In_397);
or U124 (N_124,In_1539,In_368);
nor U125 (N_125,In_198,In_2589);
xnor U126 (N_126,In_2755,In_2861);
or U127 (N_127,In_1638,In_1662);
or U128 (N_128,In_2551,In_575);
xor U129 (N_129,In_2766,In_28);
nor U130 (N_130,In_1321,In_1790);
and U131 (N_131,In_228,In_2419);
and U132 (N_132,In_431,In_1341);
and U133 (N_133,In_680,In_967);
and U134 (N_134,In_2285,In_876);
nand U135 (N_135,In_1385,In_68);
nand U136 (N_136,In_642,In_1154);
or U137 (N_137,In_733,In_2680);
and U138 (N_138,In_2573,In_2898);
nor U139 (N_139,In_2346,In_1011);
or U140 (N_140,In_1130,In_1263);
nor U141 (N_141,In_1908,In_5);
or U142 (N_142,In_432,In_1508);
and U143 (N_143,In_276,In_1839);
and U144 (N_144,In_2341,In_1355);
nor U145 (N_145,In_641,In_422);
xor U146 (N_146,In_2378,In_259);
nor U147 (N_147,In_1280,In_1969);
nor U148 (N_148,In_1027,In_712);
and U149 (N_149,In_1805,In_1909);
or U150 (N_150,In_636,In_1002);
nand U151 (N_151,In_2804,In_861);
nor U152 (N_152,In_1966,In_1878);
or U153 (N_153,In_1141,In_375);
nor U154 (N_154,In_176,In_2130);
and U155 (N_155,In_1067,In_2103);
nand U156 (N_156,In_752,In_389);
or U157 (N_157,In_2437,In_1915);
nand U158 (N_158,In_1066,In_1974);
nor U159 (N_159,In_2080,In_2671);
nor U160 (N_160,In_2506,In_1401);
xnor U161 (N_161,In_2601,In_2069);
or U162 (N_162,In_1439,In_480);
and U163 (N_163,In_433,In_2954);
nand U164 (N_164,In_2077,In_856);
nor U165 (N_165,In_155,In_2456);
nand U166 (N_166,In_288,In_193);
and U167 (N_167,In_1294,In_2743);
and U168 (N_168,In_2638,In_991);
or U169 (N_169,In_1718,In_2817);
and U170 (N_170,In_1090,In_466);
nand U171 (N_171,In_2498,In_892);
nand U172 (N_172,In_2010,In_2730);
xnor U173 (N_173,In_2301,In_1584);
or U174 (N_174,In_428,In_2108);
nor U175 (N_175,In_1436,In_434);
and U176 (N_176,In_1051,In_2065);
or U177 (N_177,In_2744,In_1388);
and U178 (N_178,In_483,In_2361);
nor U179 (N_179,In_2055,In_2090);
nand U180 (N_180,In_410,In_1833);
and U181 (N_181,In_1649,In_349);
and U182 (N_182,In_449,In_2648);
or U183 (N_183,In_1448,In_857);
nor U184 (N_184,In_545,In_2977);
or U185 (N_185,In_325,In_633);
and U186 (N_186,In_2134,In_1064);
or U187 (N_187,In_1180,In_2970);
and U188 (N_188,In_958,In_824);
and U189 (N_189,In_1943,In_544);
nand U190 (N_190,In_1652,In_2180);
or U191 (N_191,In_2228,In_2987);
nand U192 (N_192,In_2295,In_2198);
or U193 (N_193,In_1911,In_2100);
and U194 (N_194,In_2575,In_1314);
xnor U195 (N_195,In_371,In_909);
nor U196 (N_196,In_1015,In_143);
nand U197 (N_197,In_15,In_578);
nor U198 (N_198,In_206,In_2866);
nor U199 (N_199,In_399,In_2832);
or U200 (N_200,In_2181,In_765);
or U201 (N_201,In_1148,In_1641);
nand U202 (N_202,In_1973,In_1048);
nand U203 (N_203,In_2388,In_801);
nand U204 (N_204,In_688,In_2355);
nand U205 (N_205,In_1826,In_2600);
nor U206 (N_206,In_1927,In_889);
and U207 (N_207,In_490,In_248);
and U208 (N_208,In_1034,In_809);
xor U209 (N_209,In_474,In_407);
or U210 (N_210,In_82,In_2236);
or U211 (N_211,In_1825,In_1906);
nand U212 (N_212,In_1579,In_2955);
nor U213 (N_213,In_2602,In_1459);
or U214 (N_214,In_2677,In_2858);
and U215 (N_215,In_2024,In_561);
and U216 (N_216,In_711,In_1085);
xnor U217 (N_217,In_460,In_1399);
or U218 (N_218,In_2800,In_308);
xor U219 (N_219,In_2510,In_1895);
nand U220 (N_220,In_1196,In_1693);
or U221 (N_221,In_2944,In_1497);
and U222 (N_222,In_59,In_1024);
nor U223 (N_223,In_278,In_751);
nor U224 (N_224,In_478,In_2106);
or U225 (N_225,In_2318,In_2684);
nor U226 (N_226,In_1921,In_806);
and U227 (N_227,In_999,In_2663);
or U228 (N_228,In_2548,In_2981);
and U229 (N_229,In_646,In_1326);
or U230 (N_230,In_2274,In_1801);
and U231 (N_231,In_2078,In_2187);
nand U232 (N_232,In_1339,In_1496);
nand U233 (N_233,In_1615,In_247);
or U234 (N_234,In_2040,In_1279);
nand U235 (N_235,In_1093,In_88);
nand U236 (N_236,In_1156,In_2667);
nor U237 (N_237,In_1047,In_1020);
and U238 (N_238,In_379,In_896);
and U239 (N_239,In_2683,In_532);
nand U240 (N_240,In_2784,In_1567);
and U241 (N_241,In_548,In_1892);
nor U242 (N_242,In_2704,In_2316);
or U243 (N_243,In_2523,In_2877);
nand U244 (N_244,In_923,In_2362);
or U245 (N_245,In_775,In_1869);
and U246 (N_246,In_2001,In_1575);
nor U247 (N_247,In_2993,In_2820);
nand U248 (N_248,In_2919,In_2943);
nand U249 (N_249,In_166,In_2509);
or U250 (N_250,In_911,In_440);
nor U251 (N_251,In_510,In_1746);
nand U252 (N_252,In_2390,In_471);
or U253 (N_253,In_255,In_1342);
or U254 (N_254,In_2633,In_2847);
or U255 (N_255,In_707,In_650);
xnor U256 (N_256,In_2499,In_1139);
or U257 (N_257,In_1865,In_1357);
nor U258 (N_258,In_200,In_511);
or U259 (N_259,In_1188,In_1656);
or U260 (N_260,In_1126,In_2235);
nand U261 (N_261,In_1116,In_333);
and U262 (N_262,In_2294,In_719);
or U263 (N_263,In_2788,In_795);
or U264 (N_264,In_1177,In_1419);
nor U265 (N_265,In_2917,In_626);
nor U266 (N_266,In_265,In_159);
nand U267 (N_267,In_899,In_2190);
nor U268 (N_268,In_769,In_1843);
nor U269 (N_269,In_1952,In_237);
nand U270 (N_270,In_2992,In_287);
nor U271 (N_271,In_1604,In_779);
nand U272 (N_272,In_1084,In_1252);
xnor U273 (N_273,In_2963,In_900);
and U274 (N_274,In_1953,In_2066);
nor U275 (N_275,In_219,In_859);
and U276 (N_276,In_1757,In_702);
or U277 (N_277,In_2243,In_1480);
nand U278 (N_278,In_528,In_1948);
nand U279 (N_279,In_2918,In_2670);
and U280 (N_280,In_2517,In_1077);
and U281 (N_281,In_2312,In_605);
and U282 (N_282,In_218,In_2526);
nor U283 (N_283,In_2911,In_418);
nor U284 (N_284,In_2000,In_883);
and U285 (N_285,In_2062,In_481);
nor U286 (N_286,In_1687,In_2481);
nand U287 (N_287,In_36,In_2371);
or U288 (N_288,In_1688,In_1119);
nand U289 (N_289,In_2076,In_1098);
and U290 (N_290,In_2170,In_1498);
nand U291 (N_291,In_2960,In_2691);
nor U292 (N_292,In_2881,In_356);
nand U293 (N_293,In_1247,In_1956);
or U294 (N_294,In_2276,In_2984);
nor U295 (N_295,In_1335,In_138);
and U296 (N_296,In_222,In_1161);
nor U297 (N_297,In_2852,In_2192);
and U298 (N_298,In_1000,In_1520);
nor U299 (N_299,In_1103,In_1734);
nor U300 (N_300,In_136,In_1135);
nand U301 (N_301,In_1262,In_175);
and U302 (N_302,In_1989,In_1081);
or U303 (N_303,In_621,In_2706);
nor U304 (N_304,In_706,In_403);
and U305 (N_305,In_628,In_331);
or U306 (N_306,In_1963,In_757);
nor U307 (N_307,In_1542,In_1748);
nor U308 (N_308,In_1068,In_981);
or U309 (N_309,In_1492,In_1731);
nand U310 (N_310,In_2350,In_1174);
nor U311 (N_311,In_2782,In_1735);
and U312 (N_312,In_2745,In_2214);
and U313 (N_313,In_2910,In_671);
or U314 (N_314,In_83,In_1328);
nor U315 (N_315,In_1761,In_2615);
or U316 (N_316,In_2998,In_2030);
and U317 (N_317,In_2478,In_455);
nand U318 (N_318,In_2994,In_2177);
nand U319 (N_319,In_2893,In_571);
or U320 (N_320,In_1995,In_1217);
nand U321 (N_321,In_2191,In_2469);
or U322 (N_322,In_1950,In_2302);
nand U323 (N_323,In_1353,In_2525);
or U324 (N_324,In_1666,In_1102);
and U325 (N_325,In_209,In_1958);
and U326 (N_326,In_2226,In_691);
nand U327 (N_327,In_826,In_2032);
nand U328 (N_328,In_1494,In_1434);
and U329 (N_329,In_188,In_971);
nand U330 (N_330,In_1882,In_2717);
and U331 (N_331,In_1421,In_1487);
nand U332 (N_332,In_2247,In_1916);
and U333 (N_333,In_1663,In_2234);
or U334 (N_334,In_734,In_2623);
nor U335 (N_335,In_1964,In_2071);
and U336 (N_336,In_938,In_2185);
and U337 (N_337,In_447,In_2572);
nor U338 (N_338,In_1679,In_1531);
or U339 (N_339,In_1420,In_1629);
nor U340 (N_340,In_1347,In_1138);
or U341 (N_341,In_1955,In_318);
nand U342 (N_342,In_2657,In_51);
nor U343 (N_343,In_1056,In_1800);
and U344 (N_344,In_2532,In_1560);
or U345 (N_345,In_786,In_123);
nand U346 (N_346,In_866,In_354);
or U347 (N_347,In_969,In_1215);
and U348 (N_348,In_2713,In_2656);
or U349 (N_349,In_2278,In_1432);
or U350 (N_350,In_615,In_1896);
and U351 (N_351,In_1515,In_2013);
nand U352 (N_352,In_1798,In_1292);
and U353 (N_353,In_2727,In_2892);
nand U354 (N_354,In_1131,In_234);
nor U355 (N_355,In_2197,In_2369);
nor U356 (N_356,In_1842,In_348);
or U357 (N_357,In_1519,In_1369);
or U358 (N_358,In_1599,In_404);
nand U359 (N_359,In_2484,In_201);
nand U360 (N_360,In_2443,In_774);
nand U361 (N_361,In_2172,In_314);
xor U362 (N_362,In_96,In_2935);
or U363 (N_363,In_2979,In_2765);
or U364 (N_364,In_134,In_1623);
and U365 (N_365,In_101,In_260);
or U366 (N_366,In_1457,In_1782);
xor U367 (N_367,In_1636,In_360);
and U368 (N_368,In_65,In_376);
nand U369 (N_369,In_2854,In_412);
nor U370 (N_370,In_2756,In_461);
nand U371 (N_371,In_84,In_1437);
nor U372 (N_372,In_2352,In_1544);
or U373 (N_373,In_1017,In_1881);
nand U374 (N_374,In_1898,In_1558);
or U375 (N_375,In_835,In_506);
nor U376 (N_376,In_39,In_2406);
nand U377 (N_377,In_1835,In_1879);
nor U378 (N_378,In_1590,In_784);
nor U379 (N_379,In_761,In_2046);
and U380 (N_380,In_1132,In_2434);
and U381 (N_381,In_2398,In_933);
nor U382 (N_382,In_2015,In_2747);
and U383 (N_383,In_1849,In_1932);
nand U384 (N_384,In_2824,In_1461);
nand U385 (N_385,In_2439,In_2850);
nand U386 (N_386,In_1738,In_282);
nor U387 (N_387,In_332,In_1977);
nand U388 (N_388,In_2248,In_2636);
nand U389 (N_389,In_17,In_1087);
nand U390 (N_390,In_853,In_199);
and U391 (N_391,In_2289,In_2597);
and U392 (N_392,In_1143,In_2099);
and U393 (N_393,In_713,In_1403);
nor U394 (N_394,In_576,In_937);
and U395 (N_395,In_2223,In_106);
nand U396 (N_396,In_66,In_539);
nand U397 (N_397,In_854,In_1478);
and U398 (N_398,In_1041,In_2495);
nand U399 (N_399,In_413,In_799);
nand U400 (N_400,In_1134,In_402);
or U401 (N_401,In_1744,In_549);
and U402 (N_402,In_2722,In_2026);
nor U403 (N_403,In_767,In_459);
nand U404 (N_404,In_867,In_182);
and U405 (N_405,In_2121,In_989);
or U406 (N_406,In_2577,In_2061);
nor U407 (N_407,In_714,In_975);
and U408 (N_408,In_2089,In_557);
and U409 (N_409,In_1418,In_768);
nor U410 (N_410,In_541,In_1996);
or U411 (N_411,In_2401,In_1546);
or U412 (N_412,In_53,In_1268);
nor U413 (N_413,In_662,In_522);
xor U414 (N_414,In_2828,In_181);
nor U415 (N_415,In_2654,In_1643);
nand U416 (N_416,In_645,In_1828);
xnor U417 (N_417,In_2467,In_1223);
nor U418 (N_418,In_1762,In_1264);
or U419 (N_419,In_484,In_1094);
nor U420 (N_420,In_37,In_438);
nand U421 (N_421,In_1557,In_1648);
nor U422 (N_422,In_298,In_1166);
nand U423 (N_423,In_2942,In_170);
nand U424 (N_424,In_924,In_132);
and U425 (N_425,In_2105,In_2151);
and U426 (N_426,In_750,In_2758);
or U427 (N_427,In_689,In_4);
or U428 (N_428,In_1758,In_546);
and U429 (N_429,In_275,In_2771);
and U430 (N_430,In_2628,In_1712);
or U431 (N_431,In_2724,In_1697);
and U432 (N_432,In_1887,In_925);
or U433 (N_433,In_2932,In_1532);
nand U434 (N_434,In_238,In_773);
nor U435 (N_435,In_1120,In_2934);
or U436 (N_436,In_286,In_2239);
and U437 (N_437,In_202,In_1506);
or U438 (N_438,In_780,In_2562);
or U439 (N_439,In_1468,In_1529);
or U440 (N_440,In_2812,In_942);
or U441 (N_441,In_559,In_1552);
nor U442 (N_442,In_1282,In_210);
nand U443 (N_443,In_2451,In_416);
nor U444 (N_444,In_2871,In_2608);
nand U445 (N_445,In_2452,In_2);
nand U446 (N_446,In_726,In_168);
xor U447 (N_447,In_2497,In_2845);
nor U448 (N_448,In_2193,In_2022);
and U449 (N_449,In_1775,In_1269);
or U450 (N_450,In_1866,In_1767);
and U451 (N_451,In_2005,In_1222);
xnor U452 (N_452,In_1834,In_1293);
nor U453 (N_453,In_1295,In_638);
nand U454 (N_454,In_2521,In_841);
nor U455 (N_455,In_2313,In_1571);
or U456 (N_456,In_233,In_1191);
or U457 (N_457,In_2780,In_2682);
and U458 (N_458,In_1961,In_910);
and U459 (N_459,In_1713,In_1224);
and U460 (N_460,In_936,In_322);
or U461 (N_461,In_2545,In_2989);
xnor U462 (N_462,In_1417,In_1430);
nor U463 (N_463,In_2462,In_1807);
nand U464 (N_464,In_1988,In_1010);
and U465 (N_465,In_2777,In_1685);
nand U466 (N_466,In_1168,In_970);
and U467 (N_467,In_215,In_1595);
and U468 (N_468,In_1274,In_2407);
and U469 (N_469,In_1791,In_1062);
nand U470 (N_470,In_340,In_2926);
nand U471 (N_471,In_1278,In_1907);
nand U472 (N_472,In_2153,In_1237);
and U473 (N_473,In_2598,In_303);
nand U474 (N_474,In_1105,In_1137);
or U475 (N_475,In_935,In_789);
and U476 (N_476,In_2795,In_220);
xnor U477 (N_477,In_1483,In_2961);
nor U478 (N_478,In_1822,In_1129);
xnor U479 (N_479,In_731,In_1763);
or U480 (N_480,In_791,In_44);
nor U481 (N_481,In_2793,In_710);
nor U482 (N_482,In_135,In_2377);
or U483 (N_483,In_40,In_2950);
and U484 (N_484,In_940,In_718);
xor U485 (N_485,In_2924,In_187);
nor U486 (N_486,In_2659,In_2741);
or U487 (N_487,In_2326,In_274);
nor U488 (N_488,In_80,In_1639);
nand U489 (N_489,In_2339,In_2431);
and U490 (N_490,In_230,In_2646);
nor U491 (N_491,In_2502,In_1855);
nor U492 (N_492,In_519,In_2949);
nor U493 (N_493,In_2464,In_1346);
nor U494 (N_494,In_1781,In_2386);
nand U495 (N_495,In_302,In_994);
and U496 (N_496,In_406,In_1383);
nand U497 (N_497,In_2844,In_2665);
or U498 (N_498,In_1626,In_2254);
nor U499 (N_499,In_231,In_943);
xnor U500 (N_500,In_1751,In_2848);
and U501 (N_501,In_863,In_2035);
and U502 (N_502,In_1793,In_1549);
nand U503 (N_503,In_1979,In_56);
nor U504 (N_504,In_760,In_1362);
nand U505 (N_505,In_1913,In_2527);
and U506 (N_506,In_2880,In_1651);
nand U507 (N_507,In_1813,In_1250);
nand U508 (N_508,In_2188,In_831);
nand U509 (N_509,In_1303,In_1179);
and U510 (N_510,In_1946,In_1940);
nand U511 (N_511,In_1334,In_1573);
nor U512 (N_512,In_721,In_1200);
nand U513 (N_513,In_2129,In_2311);
nand U514 (N_514,In_1819,In_2503);
nor U515 (N_515,In_1711,In_805);
nand U516 (N_516,In_2564,In_1340);
or U517 (N_517,In_2635,In_1336);
nand U518 (N_518,In_1970,In_2626);
nor U519 (N_519,In_2101,In_313);
or U520 (N_520,In_75,In_2964);
or U521 (N_521,In_2815,In_1503);
nor U522 (N_522,In_2662,In_2849);
nor U523 (N_523,In_1467,In_1536);
nand U524 (N_524,In_2702,In_1667);
nor U525 (N_525,In_1861,In_1720);
and U526 (N_526,In_2028,In_1994);
or U527 (N_527,In_352,In_965);
or U528 (N_528,In_1484,In_2681);
nor U529 (N_529,In_1182,In_2846);
nand U530 (N_530,In_142,In_2508);
or U531 (N_531,In_1074,In_203);
nor U532 (N_532,In_137,In_2946);
nor U533 (N_533,In_1980,In_2480);
nand U534 (N_534,In_1811,In_454);
nor U535 (N_535,In_502,In_979);
or U536 (N_536,In_22,In_2222);
nor U537 (N_537,In_451,In_1117);
or U538 (N_538,In_1227,In_1899);
and U539 (N_539,In_1287,In_2178);
nand U540 (N_540,In_244,In_1838);
and U541 (N_541,In_895,In_1859);
and U542 (N_542,In_2271,In_903);
nor U543 (N_543,In_871,In_1710);
and U544 (N_544,In_2379,In_1935);
nor U545 (N_545,In_616,In_2068);
nand U546 (N_546,In_1845,In_1565);
or U547 (N_547,In_2430,In_1683);
nor U548 (N_548,In_2916,In_658);
nor U549 (N_549,In_2634,In_21);
and U550 (N_550,In_2265,In_848);
and U551 (N_551,In_2882,In_1990);
and U552 (N_552,In_2461,In_398);
nand U553 (N_553,In_2734,In_229);
nand U554 (N_554,In_1371,In_291);
nor U555 (N_555,In_1170,In_817);
nor U556 (N_556,In_151,In_977);
nor U557 (N_557,In_99,In_2057);
and U558 (N_558,In_2825,In_2438);
nor U559 (N_559,In_552,In_89);
nand U560 (N_560,In_2599,In_1157);
and U561 (N_561,In_507,In_1541);
nor U562 (N_562,In_2048,In_1209);
and U563 (N_563,In_1704,In_2558);
or U564 (N_564,In_1511,In_2233);
or U565 (N_565,In_830,In_2232);
xnor U566 (N_566,In_1570,In_211);
or U567 (N_567,In_1548,In_179);
and U568 (N_568,In_901,In_1118);
nand U569 (N_569,In_1065,In_2300);
and U570 (N_570,In_1937,In_2353);
nand U571 (N_571,In_885,In_1240);
nand U572 (N_572,In_2971,In_457);
or U573 (N_573,In_1453,In_1375);
nand U574 (N_574,In_2982,In_1184);
nand U575 (N_575,In_140,In_2092);
nor U576 (N_576,In_2221,In_336);
nor U577 (N_577,In_425,In_1427);
nor U578 (N_578,In_1082,In_2216);
or U579 (N_579,In_663,In_281);
nor U580 (N_580,In_1463,In_2567);
or U581 (N_581,In_2735,In_2230);
and U582 (N_582,In_2161,In_184);
nand U583 (N_583,In_2928,In_1680);
nor U584 (N_584,In_266,In_54);
and U585 (N_585,In_2445,In_1924);
nand U586 (N_586,In_1609,In_2041);
or U587 (N_587,In_2200,In_2966);
and U588 (N_588,In_2841,In_300);
nand U589 (N_589,In_2163,In_2603);
nand U590 (N_590,In_1073,In_2584);
nor U591 (N_591,In_2136,In_947);
and U592 (N_592,In_2450,In_2842);
nor U593 (N_593,In_708,In_1517);
or U594 (N_594,In_2019,In_1992);
nand U595 (N_595,In_1675,In_1533);
and U596 (N_596,In_849,In_2029);
and U597 (N_597,In_664,In_476);
nand U598 (N_598,In_591,In_2416);
and U599 (N_599,In_2189,In_683);
and U600 (N_600,In_534,In_2760);
and U601 (N_601,N_474,In_465);
and U602 (N_602,In_2283,In_2709);
and U603 (N_603,In_2025,In_631);
nor U604 (N_604,N_42,N_82);
nand U605 (N_605,N_284,In_1597);
and U606 (N_606,In_2827,In_19);
or U607 (N_607,N_255,In_2237);
or U608 (N_608,In_77,N_438);
nand U609 (N_609,In_2712,In_1766);
nor U610 (N_610,In_2280,In_2908);
nor U611 (N_611,In_2330,In_2417);
or U612 (N_612,N_447,In_1525);
nor U613 (N_613,In_430,In_14);
and U614 (N_614,In_1764,In_1079);
and U615 (N_615,In_1396,In_2468);
and U616 (N_616,In_2692,N_354);
nor U617 (N_617,In_2210,N_137);
and U618 (N_618,In_2299,In_976);
nor U619 (N_619,In_776,In_836);
or U620 (N_620,In_245,N_274);
or U621 (N_621,In_2923,In_1033);
or U622 (N_622,N_279,In_790);
nand U623 (N_623,In_249,In_392);
nor U624 (N_624,N_266,N_177);
or U625 (N_625,In_2056,N_254);
nand U626 (N_626,In_1830,In_1521);
nor U627 (N_627,In_2972,In_1331);
nand U628 (N_628,In_802,In_2500);
nor U629 (N_629,In_2536,In_2435);
or U630 (N_630,In_547,In_2394);
nor U631 (N_631,N_43,In_2110);
nor U632 (N_632,N_567,In_939);
nand U633 (N_633,N_392,N_355);
or U634 (N_634,In_369,In_1076);
or U635 (N_635,In_148,N_496);
or U636 (N_636,In_1389,In_2436);
nand U637 (N_637,In_523,In_462);
nand U638 (N_638,N_223,In_2391);
and U639 (N_639,N_133,In_1853);
nand U640 (N_640,In_1462,N_17);
nand U641 (N_641,N_588,In_1717);
nor U642 (N_642,In_2590,In_7);
nand U643 (N_643,In_1755,In_560);
nand U644 (N_644,N_262,In_1324);
or U645 (N_645,N_510,In_1178);
nand U646 (N_646,N_119,In_1045);
and U647 (N_647,In_337,In_498);
or U648 (N_648,In_2269,N_59);
nor U649 (N_649,In_2859,N_210);
and U650 (N_650,In_2673,In_85);
nand U651 (N_651,N_587,In_2279);
nor U652 (N_652,In_171,In_1984);
nor U653 (N_653,In_2494,In_1424);
and U654 (N_654,In_2409,In_778);
and U655 (N_655,N_63,In_395);
nand U656 (N_656,N_220,N_381);
xnor U657 (N_657,In_2904,In_2087);
nand U658 (N_658,N_408,In_1042);
and U659 (N_659,In_2329,In_1867);
nor U660 (N_660,In_147,In_196);
nor U661 (N_661,In_667,N_348);
or U662 (N_662,In_846,In_86);
or U663 (N_663,N_596,In_2516);
and U664 (N_664,N_484,N_538);
nor U665 (N_665,In_2128,In_2332);
nor U666 (N_666,In_258,N_418);
nand U667 (N_667,In_961,In_2305);
and U668 (N_668,In_1225,In_2447);
nor U669 (N_669,In_110,In_1678);
and U670 (N_670,In_2393,In_2797);
nor U671 (N_671,In_1344,In_2907);
nor U672 (N_672,N_136,In_2006);
and U673 (N_673,In_686,N_153);
and U674 (N_674,In_2772,N_345);
nand U675 (N_675,In_823,In_574);
and U676 (N_676,In_2574,In_1960);
or U677 (N_677,N_313,In_487);
and U678 (N_678,N_183,N_580);
nand U679 (N_679,N_5,In_1871);
or U680 (N_680,N_73,In_1312);
and U681 (N_681,In_1367,N_227);
or U682 (N_682,In_2619,In_1572);
and U683 (N_683,In_2496,In_1400);
nor U684 (N_684,N_541,In_1112);
nand U685 (N_685,N_163,In_1863);
nand U686 (N_686,N_467,In_715);
xor U687 (N_687,In_1425,In_1476);
and U688 (N_688,In_2723,In_1611);
nor U689 (N_689,In_1691,In_1220);
and U690 (N_690,In_2286,N_155);
or U691 (N_691,In_1320,In_2580);
nor U692 (N_692,In_643,In_393);
nor U693 (N_693,N_591,In_1397);
or U694 (N_694,In_783,In_2023);
nand U695 (N_695,In_2770,In_2186);
or U696 (N_696,In_2783,N_151);
nand U697 (N_697,In_2145,In_2838);
nand U698 (N_698,In_2038,N_6);
nor U699 (N_699,In_599,In_2995);
nand U700 (N_700,In_1201,In_1605);
and U701 (N_701,In_850,In_124);
nand U702 (N_702,In_1894,In_2518);
or U703 (N_703,In_2366,In_2168);
and U704 (N_704,In_870,In_1333);
nand U705 (N_705,In_1797,N_344);
nor U706 (N_706,In_2901,In_335);
or U707 (N_707,N_166,In_2306);
nand U708 (N_708,In_1715,N_522);
or U709 (N_709,N_339,In_1317);
nand U710 (N_710,In_2969,In_1627);
nand U711 (N_711,In_2351,In_2382);
nor U712 (N_712,In_1164,In_391);
or U713 (N_713,In_141,In_1245);
and U714 (N_714,In_2082,In_1640);
or U715 (N_715,N_500,In_2486);
xnor U716 (N_716,In_1657,In_197);
and U717 (N_717,N_307,N_211);
nand U718 (N_718,In_2297,N_39);
or U719 (N_719,In_60,In_1233);
or U720 (N_720,In_1837,N_531);
and U721 (N_721,In_214,In_2591);
nor U722 (N_722,In_2290,N_305);
nor U723 (N_723,In_2872,In_2194);
nor U724 (N_724,In_2582,N_368);
nor U725 (N_725,In_2678,In_1358);
xnor U726 (N_726,In_1469,N_413);
or U727 (N_727,N_280,N_555);
nor U728 (N_728,In_1423,In_682);
or U729 (N_729,N_142,N_129);
nand U730 (N_730,In_370,N_514);
and U731 (N_731,In_2579,In_2144);
or U732 (N_732,In_614,In_2166);
nand U733 (N_733,In_1677,In_486);
nor U734 (N_734,In_1155,N_189);
nand U735 (N_735,In_111,In_2256);
and U736 (N_736,In_1361,In_980);
and U737 (N_737,In_2328,N_337);
nor U738 (N_738,In_2073,In_2563);
or U739 (N_739,In_326,In_1799);
and U740 (N_740,In_608,N_525);
and U741 (N_741,In_411,In_1370);
or U742 (N_742,In_985,In_2156);
or U743 (N_743,In_242,In_1271);
nand U744 (N_744,N_135,N_564);
or U745 (N_745,In_1820,In_810);
nand U746 (N_746,In_2576,In_1086);
nand U747 (N_747,N_19,In_1050);
nand U748 (N_748,N_487,In_1472);
nand U749 (N_749,In_1070,In_1244);
and U750 (N_750,N_314,In_2571);
nand U751 (N_751,N_516,In_953);
and U752 (N_752,N_125,In_632);
nor U753 (N_753,In_2272,In_1586);
nor U754 (N_754,N_312,In_268);
or U755 (N_755,In_1277,In_530);
or U756 (N_756,N_462,In_1373);
nor U757 (N_757,In_2511,In_2675);
nand U758 (N_758,In_1936,In_1127);
or U759 (N_759,In_94,In_2334);
or U760 (N_760,In_656,In_2553);
nor U761 (N_761,In_357,In_782);
nand U762 (N_762,In_1206,N_472);
nor U763 (N_763,In_2141,In_2839);
and U764 (N_764,In_2348,N_93);
or U765 (N_765,N_287,In_2264);
nor U766 (N_766,In_1886,In_1847);
nand U767 (N_767,In_798,In_129);
and U768 (N_768,In_1337,N_170);
nor U769 (N_769,In_1987,In_1753);
or U770 (N_770,In_844,In_2740);
and U771 (N_771,N_507,In_1624);
nand U772 (N_772,In_479,In_1490);
and U773 (N_773,In_2142,In_2474);
and U774 (N_774,In_2586,In_1147);
nand U775 (N_775,In_2997,In_1165);
nand U776 (N_776,In_1858,In_2616);
or U777 (N_777,In_2514,In_1664);
and U778 (N_778,N_27,N_554);
or U779 (N_779,In_684,In_2903);
nor U780 (N_780,In_922,In_2454);
nor U781 (N_781,N_232,N_172);
xnor U782 (N_782,In_2036,N_235);
or U783 (N_783,In_1582,In_2115);
or U784 (N_784,In_1518,In_869);
and U785 (N_785,In_2725,In_1405);
xnor U786 (N_786,In_1776,In_1585);
or U787 (N_787,In_1202,N_387);
nor U788 (N_788,In_1700,In_95);
and U789 (N_789,In_20,In_1078);
nand U790 (N_790,In_609,In_1394);
nor U791 (N_791,In_232,In_50);
and U792 (N_792,N_482,In_74);
nand U793 (N_793,In_280,N_221);
nand U794 (N_794,In_2058,In_2868);
nand U795 (N_795,In_1673,In_2524);
and U796 (N_796,In_2083,In_64);
or U797 (N_797,In_208,In_635);
nand U798 (N_798,In_2937,In_1398);
and U799 (N_799,In_2152,In_1930);
nand U800 (N_800,In_1509,In_1742);
and U801 (N_801,N_468,In_2308);
nor U802 (N_802,N_53,In_1356);
nand U803 (N_803,In_1978,In_579);
nor U804 (N_804,N_530,In_660);
or U805 (N_805,In_1167,In_2957);
or U806 (N_806,In_728,In_2959);
nor U807 (N_807,In_164,N_296);
nand U808 (N_808,In_2045,In_1810);
nor U809 (N_809,N_409,In_1698);
nand U810 (N_810,In_875,In_1991);
nand U811 (N_811,N_459,In_864);
nand U812 (N_812,N_501,In_2540);
nand U813 (N_813,N_203,In_190);
and U814 (N_814,In_2126,In_2202);
xnor U815 (N_815,In_2176,In_705);
nor U816 (N_816,N_62,In_2707);
nor U817 (N_817,In_2552,In_2895);
and U818 (N_818,In_2323,In_1069);
nand U819 (N_819,In_1107,N_512);
or U820 (N_820,N_506,N_191);
and U821 (N_821,In_509,In_2043);
or U822 (N_822,In_2674,In_611);
or U823 (N_823,In_793,In_1475);
nand U824 (N_824,In_2535,In_515);
nor U825 (N_825,In_2753,In_1920);
nand U826 (N_826,In_1918,In_986);
nor U827 (N_827,In_2610,N_583);
or U828 (N_828,In_1026,In_2890);
and U829 (N_829,In_700,In_1818);
nor U830 (N_830,In_2593,In_1253);
and U831 (N_831,N_24,N_593);
nor U832 (N_832,In_73,In_157);
or U833 (N_833,In_2596,N_173);
xor U834 (N_834,In_1607,In_1298);
and U835 (N_835,In_1377,N_91);
nor U836 (N_836,N_149,In_169);
nor U837 (N_837,In_217,In_2985);
or U838 (N_838,In_504,In_653);
nand U839 (N_839,In_2491,In_2644);
nand U840 (N_840,In_2874,In_1889);
or U841 (N_841,In_1928,In_1621);
nor U842 (N_842,In_420,N_521);
nor U843 (N_843,In_76,In_2088);
and U844 (N_844,In_1444,In_254);
nor U845 (N_845,In_644,In_2373);
or U846 (N_846,In_1743,N_230);
nor U847 (N_847,In_851,In_586);
and U848 (N_848,In_623,N_394);
nor U849 (N_849,In_2869,N_281);
nand U850 (N_850,In_1150,In_104);
and U851 (N_851,N_569,In_1670);
or U852 (N_852,In_1945,N_66);
nor U853 (N_853,In_1063,In_0);
or U854 (N_854,N_115,In_383);
nor U855 (N_855,N_49,N_532);
xor U856 (N_856,In_1646,In_2209);
xnor U857 (N_857,In_1030,In_1628);
nand U858 (N_858,In_1566,In_2775);
nor U859 (N_859,In_2578,In_618);
nor U860 (N_860,N_595,In_891);
nor U861 (N_861,N_499,In_2262);
and U862 (N_862,In_821,N_15);
nor U863 (N_863,In_1266,In_1538);
or U864 (N_864,In_441,In_1305);
and U865 (N_865,In_328,N_439);
nand U866 (N_866,N_10,N_31);
xor U867 (N_867,N_396,N_423);
nor U868 (N_868,In_2183,In_2171);
or U869 (N_869,In_832,In_887);
and U870 (N_870,In_2976,N_425);
or U871 (N_871,In_1732,In_670);
nand U872 (N_872,In_2618,N_380);
nand U873 (N_873,In_178,In_820);
and U874 (N_874,N_74,In_1443);
nand U875 (N_875,N_575,N_465);
nand U876 (N_876,N_25,In_1578);
nor U877 (N_877,N_245,In_1721);
and U878 (N_878,In_1857,In_2652);
xnor U879 (N_879,In_668,In_978);
xnor U880 (N_880,N_405,In_554);
and U881 (N_881,N_156,N_326);
nand U882 (N_882,In_9,N_359);
nand U883 (N_883,In_2980,In_1773);
or U884 (N_884,In_43,N_34);
or U885 (N_885,N_469,In_1275);
and U886 (N_886,In_1160,In_1986);
or U887 (N_887,N_316,In_973);
nand U888 (N_888,In_2640,N_318);
nand U889 (N_889,In_2607,N_527);
nand U890 (N_890,In_122,N_70);
nand U891 (N_891,In_1832,In_1198);
nor U892 (N_892,In_764,In_2205);
nand U893 (N_893,In_1962,In_473);
nand U894 (N_894,In_2376,In_927);
or U895 (N_895,N_519,In_674);
nor U896 (N_896,In_1535,In_2778);
and U897 (N_897,N_357,In_893);
and U898 (N_898,In_884,In_1350);
and U899 (N_899,N_376,In_1486);
or U900 (N_900,N_520,In_2059);
nand U901 (N_901,In_577,N_363);
or U902 (N_902,N_292,In_619);
nand U903 (N_903,In_2044,In_2912);
xnor U904 (N_904,N_148,In_2703);
or U905 (N_905,N_406,In_2363);
nor U906 (N_906,In_1588,In_1109);
and U907 (N_907,In_373,In_1528);
and U908 (N_908,In_1674,In_2007);
nor U909 (N_909,In_2063,In_1516);
nand U910 (N_910,In_1589,In_212);
or U911 (N_911,In_957,In_2487);
or U912 (N_912,N_197,N_452);
or U913 (N_913,In_1736,In_1784);
nor U914 (N_914,In_567,In_1512);
or U915 (N_915,N_502,In_1199);
and U916 (N_916,In_1123,N_108);
or U917 (N_917,N_160,N_64);
or U918 (N_918,In_1603,In_472);
nand U919 (N_919,In_323,In_617);
nand U920 (N_920,In_2885,In_2444);
and U921 (N_921,In_2581,N_80);
nand U922 (N_922,N_278,N_293);
nor U923 (N_923,N_404,In_292);
or U924 (N_924,N_533,In_125);
or U925 (N_925,In_1386,In_735);
nor U926 (N_926,In_2453,In_1574);
nor U927 (N_927,N_257,In_2335);
nand U928 (N_928,N_3,N_68);
or U929 (N_929,In_2257,In_192);
nor U930 (N_930,In_496,N_22);
nor U931 (N_931,N_561,In_450);
nand U932 (N_932,N_71,In_1226);
and U933 (N_933,In_2840,In_882);
or U934 (N_934,In_1232,In_263);
nor U935 (N_935,In_2676,In_2164);
or U936 (N_936,In_2042,In_622);
nor U937 (N_937,In_2135,In_746);
and U938 (N_938,In_1110,In_1189);
nor U939 (N_939,In_1316,In_2967);
nor U940 (N_940,In_1393,In_1464);
nand U941 (N_941,In_343,N_167);
and U942 (N_942,In_2282,In_49);
and U943 (N_943,In_1501,In_1364);
or U944 (N_944,In_968,N_370);
or U945 (N_945,N_457,In_1481);
nor U946 (N_946,N_11,In_868);
nor U947 (N_947,In_2947,In_423);
and U948 (N_948,In_697,In_2383);
or U949 (N_949,In_2034,In_1745);
and U950 (N_950,In_1829,In_926);
nand U951 (N_951,In_1740,In_1897);
nand U952 (N_952,In_2519,In_1931);
and U953 (N_953,In_1770,N_273);
nor U954 (N_954,In_556,In_2412);
nand U955 (N_955,In_2054,N_85);
nand U956 (N_956,N_195,In_1537);
nand U957 (N_957,In_1780,In_299);
or U958 (N_958,In_1429,In_2718);
nor U959 (N_959,In_2085,In_329);
or U960 (N_960,N_548,In_2620);
or U961 (N_961,In_555,In_114);
xnor U962 (N_962,N_308,N_327);
or U963 (N_963,In_1151,In_898);
nor U964 (N_964,In_1929,In_2260);
or U965 (N_965,In_2009,N_386);
nor U966 (N_966,In_897,In_944);
or U967 (N_967,In_1959,N_529);
nor U968 (N_968,In_2556,In_2238);
nor U969 (N_969,In_1228,In_367);
xor U970 (N_970,N_295,In_1903);
nand U971 (N_971,In_2251,In_426);
nor U972 (N_972,In_995,In_2693);
and U973 (N_973,In_1125,In_597);
nand U974 (N_974,N_171,In_1760);
and U975 (N_975,In_1479,In_570);
or U976 (N_976,In_1404,N_414);
nor U977 (N_977,In_1686,N_196);
and U978 (N_978,N_347,In_1771);
xnor U979 (N_979,In_1097,In_2470);
nand U980 (N_980,N_182,In_1054);
or U981 (N_981,In_1046,N_219);
and U982 (N_982,In_1971,In_1267);
nand U983 (N_983,In_1888,In_974);
and U984 (N_984,In_2515,In_1212);
nand U985 (N_985,N_574,N_101);
or U986 (N_986,In_2655,In_2067);
nor U987 (N_987,In_1777,In_816);
nor U988 (N_988,In_1387,N_491);
and U989 (N_989,In_1,In_289);
nor U990 (N_990,N_536,In_2796);
or U991 (N_991,N_131,In_2485);
or U992 (N_992,In_1001,N_475);
nand U993 (N_993,In_2359,N_460);
nand U994 (N_994,In_2365,In_983);
or U995 (N_995,In_1106,In_1999);
nor U996 (N_996,In_624,In_2364);
or U997 (N_997,In_2442,N_571);
nand U998 (N_998,In_1241,In_1008);
nand U999 (N_999,In_11,N_388);
or U1000 (N_1000,In_1144,In_1904);
and U1001 (N_1001,In_2387,In_1175);
nor U1002 (N_1002,In_1190,In_825);
nand U1003 (N_1003,N_277,In_1169);
or U1004 (N_1004,N_100,In_2695);
nand U1005 (N_1005,In_2458,In_2592);
and U1006 (N_1006,In_996,In_113);
nor U1007 (N_1007,In_2696,In_722);
and U1008 (N_1008,N_239,In_409);
and U1009 (N_1009,In_1186,N_397);
nor U1010 (N_1010,In_2973,In_1634);
and U1011 (N_1011,In_2700,N_353);
or U1012 (N_1012,In_701,In_2184);
nor U1013 (N_1013,In_1625,In_435);
and U1014 (N_1014,In_666,N_226);
nand U1015 (N_1015,In_186,In_533);
or U1016 (N_1016,In_2336,In_2883);
and U1017 (N_1017,In_394,In_2549);
and U1018 (N_1018,In_1592,In_917);
nand U1019 (N_1019,In_673,In_743);
nand U1020 (N_1020,N_325,In_1510);
nand U1021 (N_1021,N_169,In_777);
nor U1022 (N_1022,N_497,In_2217);
or U1023 (N_1023,In_146,In_1171);
and U1024 (N_1024,In_456,In_107);
or U1025 (N_1025,N_420,In_493);
or U1026 (N_1026,In_2344,N_509);
or U1027 (N_1027,In_296,In_736);
nor U1028 (N_1028,In_877,In_1101);
or U1029 (N_1029,In_1128,N_237);
nor U1030 (N_1030,N_188,In_1957);
nor U1031 (N_1031,In_2482,In_2658);
or U1032 (N_1032,In_516,In_1019);
nor U1033 (N_1033,In_582,N_132);
or U1034 (N_1034,In_23,In_1219);
nand U1035 (N_1035,In_1204,In_2534);
nand U1036 (N_1036,In_1007,In_1140);
and U1037 (N_1037,In_665,In_1111);
nand U1038 (N_1038,In_2627,N_455);
nand U1039 (N_1039,N_464,N_350);
nor U1040 (N_1040,In_2244,In_2479);
xnor U1041 (N_1041,In_2093,In_1411);
or U1042 (N_1042,In_2520,N_495);
or U1043 (N_1043,In_651,In_1910);
and U1044 (N_1044,In_2267,N_60);
or U1045 (N_1045,In_2544,In_2206);
and U1046 (N_1046,In_1724,In_526);
and U1047 (N_1047,N_184,In_982);
and U1048 (N_1048,In_63,In_2522);
or U1049 (N_1049,In_503,In_1660);
and U1050 (N_1050,In_443,In_1307);
or U1051 (N_1051,In_2167,In_2809);
nand U1052 (N_1052,N_120,In_477);
nand U1053 (N_1053,N_116,In_2466);
nor U1054 (N_1054,In_2621,In_2806);
nor U1055 (N_1055,In_1655,In_1747);
and U1056 (N_1056,In_1672,In_2501);
or U1057 (N_1057,In_2736,N_92);
nand U1058 (N_1058,In_448,In_1122);
nor U1059 (N_1059,In_1868,In_834);
nand U1060 (N_1060,N_20,N_57);
nand U1061 (N_1061,In_1230,N_585);
nor U1062 (N_1062,In_2936,N_374);
nor U1063 (N_1063,In_1061,In_766);
nand U1064 (N_1064,In_1029,In_2690);
nor U1065 (N_1065,In_1037,In_1451);
and U1066 (N_1066,N_503,In_223);
nand U1067 (N_1067,N_402,N_598);
xor U1068 (N_1068,In_81,In_284);
or U1069 (N_1069,In_2112,In_261);
nor U1070 (N_1070,N_550,N_168);
and U1071 (N_1071,In_1049,In_993);
xor U1072 (N_1072,N_48,In_2384);
and U1073 (N_1073,In_1258,In_808);
nor U1074 (N_1074,In_304,In_2504);
and U1075 (N_1075,In_239,In_878);
nor U1076 (N_1076,N_222,N_546);
or U1077 (N_1077,In_45,In_536);
nand U1078 (N_1078,In_1949,N_297);
and U1079 (N_1079,In_419,In_1794);
nand U1080 (N_1080,In_2225,In_694);
and U1081 (N_1081,In_1485,In_2195);
and U1082 (N_1082,In_1635,In_2021);
nand U1083 (N_1083,In_2263,N_21);
nand U1084 (N_1084,N_185,In_2776);
nand U1085 (N_1085,N_403,In_879);
nor U1086 (N_1086,In_934,In_1694);
nand U1087 (N_1087,In_1493,In_1197);
or U1088 (N_1088,N_269,N_46);
and U1089 (N_1089,In_1642,In_2774);
or U1090 (N_1090,N_105,In_240);
or U1091 (N_1091,N_551,In_2876);
nand U1092 (N_1092,In_1378,In_2242);
nor U1093 (N_1093,In_489,In_2708);
or U1094 (N_1094,In_2091,In_468);
nand U1095 (N_1095,N_539,In_2931);
nor U1096 (N_1096,In_1060,In_1159);
and U1097 (N_1097,In_739,In_2829);
nor U1098 (N_1098,In_525,In_1450);
or U1099 (N_1099,N_41,In_2802);
nor U1100 (N_1100,In_2647,In_344);
xnor U1101 (N_1101,In_992,In_990);
or U1102 (N_1102,In_640,N_597);
nand U1103 (N_1103,In_1596,N_289);
and U1104 (N_1104,In_524,N_246);
nor U1105 (N_1105,N_400,In_2629);
nand U1106 (N_1106,N_586,In_2104);
or U1107 (N_1107,In_669,In_1540);
nor U1108 (N_1108,In_321,N_523);
nor U1109 (N_1109,N_332,In_2685);
or U1110 (N_1110,In_2159,In_1096);
nand U1111 (N_1111,In_2568,In_2457);
or U1112 (N_1112,In_195,N_300);
or U1113 (N_1113,In_250,In_1526);
or U1114 (N_1114,N_473,In_246);
or U1115 (N_1115,N_419,In_1543);
or U1116 (N_1116,N_454,N_338);
or U1117 (N_1117,In_1701,In_2902);
nor U1118 (N_1118,In_794,In_1706);
nor U1119 (N_1119,In_2052,In_747);
nand U1120 (N_1120,In_1500,In_913);
or U1121 (N_1121,N_123,N_389);
or U1122 (N_1122,N_78,In_2441);
or U1123 (N_1123,In_1014,In_1727);
nand U1124 (N_1124,N_385,In_2400);
nor U1125 (N_1125,In_2291,In_191);
nand U1126 (N_1126,In_1458,N_592);
nand U1127 (N_1127,N_52,In_1313);
nor U1128 (N_1128,N_304,N_407);
and U1129 (N_1129,N_140,In_1555);
nand U1130 (N_1130,N_243,In_482);
or U1131 (N_1131,N_102,N_549);
nand U1132 (N_1132,N_88,N_30);
or U1133 (N_1133,N_9,In_2821);
nand U1134 (N_1134,In_948,In_1149);
nand U1135 (N_1135,In_492,In_2392);
and U1136 (N_1136,In_109,N_67);
or U1137 (N_1137,In_310,N_431);
nand U1138 (N_1138,In_2273,In_2146);
or U1139 (N_1139,N_29,In_1692);
and U1140 (N_1140,N_72,In_1231);
or U1141 (N_1141,In_2705,In_1080);
nand U1142 (N_1142,In_1851,N_461);
or U1143 (N_1143,In_1728,In_1545);
nor U1144 (N_1144,In_600,In_2865);
nor U1145 (N_1145,In_2697,In_1919);
and U1146 (N_1146,N_253,In_2420);
and U1147 (N_1147,In_565,In_319);
or U1148 (N_1148,In_2064,In_71);
nand U1149 (N_1149,In_2990,In_2721);
nor U1150 (N_1150,In_2886,In_2650);
nor U1151 (N_1151,N_236,In_984);
and U1152 (N_1152,In_1561,In_2429);
or U1153 (N_1153,In_347,In_1276);
nor U1154 (N_1154,In_33,In_1152);
nand U1155 (N_1155,In_950,In_1922);
or U1156 (N_1156,N_384,In_601);
and U1157 (N_1157,In_2375,In_590);
and U1158 (N_1158,N_18,In_2560);
nand U1159 (N_1159,In_756,N_428);
and U1160 (N_1160,In_2996,In_862);
xor U1161 (N_1161,In_858,In_1018);
or U1162 (N_1162,In_1213,In_2039);
nand U1163 (N_1163,N_175,N_590);
nor U1164 (N_1164,N_12,In_1306);
nand U1165 (N_1165,N_393,In_2941);
or U1166 (N_1166,In_1788,In_1329);
nand U1167 (N_1167,In_807,In_2864);
nor U1168 (N_1168,In_2528,In_1055);
nor U1169 (N_1169,In_2140,N_433);
and U1170 (N_1170,In_1815,In_2255);
nor U1171 (N_1171,N_282,In_2728);
and U1172 (N_1172,In_2816,In_2594);
nor U1173 (N_1173,N_47,In_1058);
or U1174 (N_1174,In_1917,N_121);
or U1175 (N_1175,In_1133,In_2303);
and U1176 (N_1176,In_139,In_272);
nand U1177 (N_1177,N_391,In_1248);
or U1178 (N_1178,N_352,In_2120);
nand U1179 (N_1179,In_872,In_2530);
nor U1180 (N_1180,In_2953,In_1214);
nand U1181 (N_1181,In_2125,In_1441);
nor U1182 (N_1182,In_301,N_56);
or U1183 (N_1183,In_678,In_1901);
or U1184 (N_1184,In_2818,In_2097);
xor U1185 (N_1185,In_377,In_2787);
nand U1186 (N_1186,In_1504,N_329);
nor U1187 (N_1187,In_1363,In_2288);
and U1188 (N_1188,In_2933,In_366);
and U1189 (N_1189,In_537,In_1951);
or U1190 (N_1190,In_2492,In_72);
nor U1191 (N_1191,In_1547,N_552);
and U1192 (N_1192,In_1554,In_1146);
nor U1193 (N_1193,In_543,In_2293);
and U1194 (N_1194,In_551,N_158);
nor U1195 (N_1195,In_216,In_987);
nand U1196 (N_1196,N_331,In_1614);
nor U1197 (N_1197,N_79,In_117);
nand U1198 (N_1198,In_902,In_1454);
nor U1199 (N_1199,N_261,In_1003);
nand U1200 (N_1200,In_2798,In_1322);
nand U1201 (N_1201,In_1239,N_799);
nor U1202 (N_1202,N_434,In_359);
or U1203 (N_1203,N_867,N_940);
and U1204 (N_1204,N_779,N_1034);
nor U1205 (N_1205,In_1709,N_634);
or U1206 (N_1206,N_451,In_2287);
nor U1207 (N_1207,In_797,In_1283);
nor U1208 (N_1208,In_2079,In_363);
nor U1209 (N_1209,In_1965,N_966);
xnor U1210 (N_1210,In_2611,N_793);
nand U1211 (N_1211,N_720,N_373);
xor U1212 (N_1212,In_945,In_550);
nor U1213 (N_1213,In_748,In_2333);
nor U1214 (N_1214,N_1101,In_2811);
nor U1215 (N_1215,In_681,N_809);
nor U1216 (N_1216,In_1366,In_1972);
nor U1217 (N_1217,In_2418,N_463);
or U1218 (N_1218,In_133,In_2694);
and U1219 (N_1219,In_1844,In_1733);
nand U1220 (N_1220,N_792,In_1390);
or U1221 (N_1221,In_3,N_919);
or U1222 (N_1222,N_272,N_959);
and U1223 (N_1223,N_696,N_340);
nand U1224 (N_1224,N_466,N_204);
and U1225 (N_1225,In_1031,In_31);
nand U1226 (N_1226,N_703,In_1238);
nand U1227 (N_1227,In_2925,In_672);
nand U1228 (N_1228,N_217,In_2446);
nor U1229 (N_1229,N_214,N_1026);
and U1230 (N_1230,In_97,In_2207);
nand U1231 (N_1231,In_424,In_629);
xnor U1232 (N_1232,In_1285,N_1159);
nor U1233 (N_1233,In_27,In_2098);
nor U1234 (N_1234,In_2037,In_771);
and U1235 (N_1235,In_2169,In_1759);
nand U1236 (N_1236,N_178,N_765);
nor U1237 (N_1237,In_2733,In_2891);
xor U1238 (N_1238,N_1168,N_984);
nor U1239 (N_1239,In_1301,In_1840);
nor U1240 (N_1240,In_758,In_649);
nand U1241 (N_1241,In_1564,N_488);
nand U1242 (N_1242,N_106,In_500);
nor U1243 (N_1243,N_234,In_2476);
or U1244 (N_1244,N_743,N_320);
and U1245 (N_1245,In_204,In_2426);
or U1246 (N_1246,N_1123,In_2643);
nand U1247 (N_1247,N_625,N_553);
or U1248 (N_1248,N_1188,N_946);
nand U1249 (N_1249,In_2905,N_366);
or U1250 (N_1250,In_1059,In_469);
and U1251 (N_1251,In_470,In_955);
and U1252 (N_1252,N_700,In_676);
and U1253 (N_1253,N_1019,N_1040);
and U1254 (N_1254,N_826,In_2833);
nand U1255 (N_1255,In_2182,N_37);
nor U1256 (N_1256,In_495,In_2196);
and U1257 (N_1257,N_437,N_850);
nor U1258 (N_1258,N_1066,In_1502);
and U1259 (N_1259,N_736,N_855);
and U1260 (N_1260,In_2945,In_2889);
nand U1261 (N_1261,In_2147,N_1008);
and U1262 (N_1262,In_1507,In_16);
nor U1263 (N_1263,N_727,N_306);
nand U1264 (N_1264,N_77,In_865);
nand U1265 (N_1265,In_2661,In_442);
nor U1266 (N_1266,In_2231,In_87);
and U1267 (N_1267,In_1446,N_89);
or U1268 (N_1268,N_377,N_1005);
and U1269 (N_1269,In_1669,In_1676);
and U1270 (N_1270,N_65,In_1249);
and U1271 (N_1271,N_717,N_761);
nand U1272 (N_1272,In_772,N_927);
nor U1273 (N_1273,In_172,In_1559);
nor U1274 (N_1274,N_1174,In_364);
or U1275 (N_1275,In_709,N_224);
nand U1276 (N_1276,N_738,N_895);
and U1277 (N_1277,In_1194,N_1058);
nand U1278 (N_1278,In_1726,In_1689);
and U1279 (N_1279,In_1513,In_603);
or U1280 (N_1280,N_528,In_2687);
and U1281 (N_1281,N_44,N_915);
and U1282 (N_1282,N_1028,N_576);
nand U1283 (N_1283,N_1055,N_1172);
nand U1284 (N_1284,N_849,N_1179);
nor U1285 (N_1285,N_476,N_1139);
and U1286 (N_1286,N_752,N_942);
xnor U1287 (N_1287,In_130,N_971);
and U1288 (N_1288,In_915,In_1254);
xor U1289 (N_1289,N_974,In_1831);
and U1290 (N_1290,N_268,N_283);
and U1291 (N_1291,N_113,N_1082);
nand U1292 (N_1292,N_914,In_1702);
xor U1293 (N_1293,In_2204,In_840);
and U1294 (N_1294,In_569,In_1739);
or U1295 (N_1295,N_260,In_390);
or U1296 (N_1296,N_609,N_782);
nor U1297 (N_1297,N_1166,In_1905);
or U1298 (N_1298,In_1653,In_595);
and U1299 (N_1299,N_714,In_70);
nand U1300 (N_1300,N_252,N_1083);
and U1301 (N_1301,In_2875,In_1229);
or U1302 (N_1302,In_2116,N_362);
nor U1303 (N_1303,N_726,N_118);
nor U1304 (N_1304,N_104,N_864);
or U1305 (N_1305,N_747,N_1175);
nor U1306 (N_1306,N_122,N_298);
and U1307 (N_1307,In_2605,N_1018);
or U1308 (N_1308,N_824,N_734);
and U1309 (N_1309,In_458,In_501);
nor U1310 (N_1310,In_1113,In_1716);
or U1311 (N_1311,In_2122,N_909);
nor U1312 (N_1312,N_524,In_2014);
and U1313 (N_1313,N_901,In_173);
nor U1314 (N_1314,In_1696,In_2173);
and U1315 (N_1315,N_650,N_920);
xor U1316 (N_1316,N_957,In_2894);
and U1317 (N_1317,N_1129,N_859);
nor U1318 (N_1318,In_2805,In_2867);
nand U1319 (N_1319,N_545,In_770);
or U1320 (N_1320,In_1856,In_2053);
nor U1321 (N_1321,In_2554,In_508);
nand U1322 (N_1322,N_745,In_1281);
and U1323 (N_1323,N_916,N_1130);
nor U1324 (N_1324,In_1088,N_929);
nor U1325 (N_1325,N_328,N_719);
nand U1326 (N_1326,N_669,In_2668);
or U1327 (N_1327,N_663,In_2762);
nor U1328 (N_1328,N_1105,In_283);
nand U1329 (N_1329,N_95,N_694);
nand U1330 (N_1330,N_55,N_505);
and U1331 (N_1331,N_813,In_2215);
or U1332 (N_1332,In_154,N_1045);
and U1333 (N_1333,In_2710,N_860);
or U1334 (N_1334,N_1044,N_334);
xnor U1335 (N_1335,In_845,In_612);
nand U1336 (N_1336,In_717,N_623);
and U1337 (N_1337,In_960,N_775);
or U1338 (N_1338,In_1708,In_581);
or U1339 (N_1339,In_1005,In_243);
nand U1340 (N_1340,In_2719,N_490);
nand U1341 (N_1341,N_756,In_1428);
nor U1342 (N_1342,In_1785,In_657);
nand U1343 (N_1343,N_1192,N_679);
or U1344 (N_1344,N_432,In_763);
nor U1345 (N_1345,N_684,In_792);
and U1346 (N_1346,In_754,In_1040);
nor U1347 (N_1347,In_1947,N_250);
xnor U1348 (N_1348,In_35,N_953);
or U1349 (N_1349,In_1613,N_448);
nand U1350 (N_1350,In_527,N_429);
nor U1351 (N_1351,In_1104,N_1090);
or U1352 (N_1352,In_518,In_1315);
nor U1353 (N_1353,In_1821,In_2631);
or U1354 (N_1354,N_721,In_928);
xnor U1355 (N_1355,N_1038,N_846);
nand U1356 (N_1356,In_568,N_751);
or U1357 (N_1357,N_213,N_993);
and U1358 (N_1358,N_1199,In_2555);
nand U1359 (N_1359,N_1095,N_996);
or U1360 (N_1360,In_1021,In_2471);
xnor U1361 (N_1361,In_2327,In_2410);
and U1362 (N_1362,N_130,In_998);
and U1363 (N_1363,N_422,In_860);
or U1364 (N_1364,In_467,N_150);
nor U1365 (N_1365,In_1580,N_897);
nor U1366 (N_1366,N_805,In_2792);
or U1367 (N_1367,In_2897,N_930);
or U1368 (N_1368,In_2081,In_2888);
and U1369 (N_1369,In_1382,N_286);
nor U1370 (N_1370,In_12,In_61);
xnor U1371 (N_1371,N_441,N_358);
and U1372 (N_1372,N_299,N_903);
and U1373 (N_1373,In_585,In_2372);
and U1374 (N_1374,In_2133,In_2952);
nand U1375 (N_1375,N_666,In_1591);
xor U1376 (N_1376,In_2249,N_1069);
or U1377 (N_1377,N_1029,N_445);
nor U1378 (N_1378,In_563,In_2779);
or U1379 (N_1379,N_670,In_695);
or U1380 (N_1380,N_656,In_1265);
xnor U1381 (N_1381,In_290,In_2345);
nand U1382 (N_1382,In_2810,In_729);
and U1383 (N_1383,N_1127,In_592);
and U1384 (N_1384,N_157,In_997);
nand U1385 (N_1385,In_1013,N_547);
or U1386 (N_1386,In_1941,N_477);
nor U1387 (N_1387,In_2033,N_1003);
nand U1388 (N_1388,In_1022,N_435);
nor U1389 (N_1389,In_1210,N_817);
nand U1390 (N_1390,N_212,N_86);
or U1391 (N_1391,N_1102,In_1192);
nor U1392 (N_1392,N_653,N_685);
nand U1393 (N_1393,In_1527,In_1442);
nand U1394 (N_1394,In_163,In_1052);
nor U1395 (N_1395,In_505,In_2768);
or U1396 (N_1396,N_992,In_842);
nor U1397 (N_1397,In_625,N_302);
or U1398 (N_1398,N_1096,In_1602);
and U1399 (N_1399,In_2649,N_768);
and U1400 (N_1400,N_341,In_1556);
nor U1401 (N_1401,In_1981,N_847);
nand U1402 (N_1402,N_954,In_330);
or U1403 (N_1403,N_839,In_2731);
and U1404 (N_1404,N_1064,In_1354);
and U1405 (N_1405,N_1042,N_998);
and U1406 (N_1406,In_2751,In_2175);
nand U1407 (N_1407,N_493,In_150);
nand U1408 (N_1408,In_573,N_424);
or U1409 (N_1409,In_890,N_557);
or U1410 (N_1410,In_855,N_1037);
and U1411 (N_1411,In_444,In_67);
nor U1412 (N_1412,N_117,N_1153);
or U1413 (N_1413,N_1189,In_2986);
and U1414 (N_1414,N_710,In_538);
or U1415 (N_1415,In_2588,N_563);
nor U1416 (N_1416,N_111,N_568);
or U1417 (N_1417,In_1243,N_871);
and U1418 (N_1418,In_2317,In_345);
nor U1419 (N_1419,N_40,In_1873);
nor U1420 (N_1420,In_1440,N_218);
and U1421 (N_1421,In_880,N_771);
or U1422 (N_1422,N_361,N_784);
or U1423 (N_1423,N_1009,In_1684);
and U1424 (N_1424,N_542,In_415);
and U1425 (N_1425,In_1349,In_2160);
nand U1426 (N_1426,In_2752,In_1345);
and U1427 (N_1427,N_683,N_619);
or U1428 (N_1428,In_2138,N_975);
or U1429 (N_1429,N_410,N_815);
or U1430 (N_1430,N_248,N_383);
nand U1431 (N_1431,In_1875,N_822);
nor U1432 (N_1432,In_2913,N_599);
nand U1433 (N_1433,In_803,In_2060);
and U1434 (N_1434,N_395,In_2857);
nor U1435 (N_1435,In_1414,In_2315);
nor U1436 (N_1436,N_534,In_1163);
nand U1437 (N_1437,N_785,In_144);
and U1438 (N_1438,N_1094,N_1191);
nor U1439 (N_1439,In_2179,N_1165);
and U1440 (N_1440,In_2349,N_937);
nor U1441 (N_1441,N_321,In_2162);
and U1442 (N_1442,In_1695,N_637);
nor U1443 (N_1443,N_945,In_2750);
or U1444 (N_1444,N_661,In_2823);
and U1445 (N_1445,In_2565,In_79);
and U1446 (N_1446,In_1255,N_1075);
nor U1447 (N_1447,In_6,N_881);
nor U1448 (N_1448,N_1006,N_84);
nand U1449 (N_1449,In_2261,In_796);
and U1450 (N_1450,In_2208,N_336);
and U1451 (N_1451,N_865,N_825);
nand U1452 (N_1452,N_205,N_187);
or U1453 (N_1453,N_1049,N_489);
nor U1454 (N_1454,In_2624,In_2307);
or U1455 (N_1455,In_2137,N_127);
and U1456 (N_1456,N_288,N_4);
and U1457 (N_1457,N_225,In_2834);
nand U1458 (N_1458,N_910,N_570);
nand U1459 (N_1459,In_271,In_2220);
and U1460 (N_1460,N_654,N_811);
or U1461 (N_1461,In_1038,In_2111);
or U1462 (N_1462,N_426,N_731);
or U1463 (N_1463,N_1167,N_797);
nand U1464 (N_1464,N_513,In_2199);
and U1465 (N_1465,N_778,In_2284);
and U1466 (N_1466,In_2711,N_256);
nor U1467 (N_1467,In_2124,In_2117);
nand U1468 (N_1468,N_436,N_1022);
or U1469 (N_1469,In_2370,N_1110);
or U1470 (N_1470,In_881,In_2794);
or U1471 (N_1471,N_950,N_1081);
or U1472 (N_1472,In_894,N_1183);
and U1473 (N_1473,N_594,In_723);
xnor U1474 (N_1474,N_535,N_600);
nand U1475 (N_1475,In_699,In_2154);
xor U1476 (N_1476,N_76,N_614);
nor U1477 (N_1477,In_1668,N_816);
or U1478 (N_1478,N_1187,N_842);
nor U1479 (N_1479,N_1,N_1148);
and U1480 (N_1480,In_24,N_275);
and U1481 (N_1481,N_124,In_1032);
nand U1482 (N_1482,N_50,N_691);
nor U1483 (N_1483,In_324,In_452);
xnor U1484 (N_1484,In_972,N_964);
or U1485 (N_1485,In_2331,In_2625);
or U1486 (N_1486,N_828,N_617);
nor U1487 (N_1487,N_1061,In_1359);
nor U1488 (N_1488,In_1954,In_2505);
or U1489 (N_1489,N_851,N_152);
or U1490 (N_1490,N_643,In_194);
nor U1491 (N_1491,In_1323,In_2449);
nand U1492 (N_1492,N_1052,In_2860);
nand U1493 (N_1493,In_127,In_2738);
nor U1494 (N_1494,In_873,In_2884);
nor U1495 (N_1495,N_757,N_1020);
nor U1496 (N_1496,In_1153,N_258);
or U1497 (N_1497,In_2270,In_2448);
xor U1498 (N_1498,In_488,In_815);
and U1499 (N_1499,In_358,N_660);
nand U1500 (N_1500,In_2113,N_1078);
nand U1501 (N_1501,In_2324,In_2999);
nand U1502 (N_1502,In_1563,In_162);
or U1503 (N_1503,In_1426,N_680);
and U1504 (N_1504,N_838,N_952);
and U1505 (N_1505,In_745,N_777);
and U1506 (N_1506,N_581,N_961);
nor U1507 (N_1507,N_922,In_2084);
nand U1508 (N_1508,N_633,N_810);
and U1509 (N_1509,In_1343,In_2259);
nor U1510 (N_1510,N_498,N_837);
or U1511 (N_1511,In_2789,In_2896);
or U1512 (N_1512,N_578,In_2761);
nand U1513 (N_1513,In_606,In_513);
nand U1514 (N_1514,N_605,In_613);
nor U1515 (N_1515,In_2354,In_916);
nor U1516 (N_1516,N_1031,N_1046);
nor U1517 (N_1517,In_2587,In_2158);
or U1518 (N_1518,N_54,N_644);
and U1519 (N_1519,N_1162,In_297);
nand U1520 (N_1520,In_158,N_365);
or U1521 (N_1521,N_707,N_773);
xor U1522 (N_1522,In_2460,N_896);
and U1523 (N_1523,N_632,In_1645);
and U1524 (N_1524,In_361,N_658);
and U1525 (N_1525,N_819,N_75);
nor U1526 (N_1526,N_589,N_943);
or U1527 (N_1527,In_1926,In_92);
nand U1528 (N_1528,N_613,N_958);
or U1529 (N_1529,In_1284,In_295);
and U1530 (N_1530,N_968,In_954);
nand U1531 (N_1531,In_1162,In_2477);
nor U1532 (N_1532,N_651,N_845);
nand U1533 (N_1533,N_967,N_2);
and U1534 (N_1534,In_439,N_990);
and U1535 (N_1535,N_812,N_238);
and U1536 (N_1536,N_1133,N_631);
or U1537 (N_1537,N_1053,N_655);
nand U1538 (N_1538,N_960,In_1207);
or U1539 (N_1539,In_2016,N_323);
nand U1540 (N_1540,In_1327,N_16);
nand U1541 (N_1541,In_738,In_400);
nand U1542 (N_1542,N_907,In_427);
xor U1543 (N_1543,In_584,In_2118);
nor U1544 (N_1544,N_759,N_126);
nor U1545 (N_1545,In_1530,N_1104);
nand U1546 (N_1546,N_1157,In_2321);
or U1547 (N_1547,N_1051,N_814);
nor U1548 (N_1548,In_225,N_1196);
or U1549 (N_1549,N_401,In_2314);
or U1550 (N_1550,N_889,In_320);
or U1551 (N_1551,In_499,In_1550);
and U1552 (N_1552,In_2432,In_262);
nor U1553 (N_1553,N_83,In_2853);
nor U1554 (N_1554,In_351,N_832);
or U1555 (N_1555,In_685,In_381);
nor U1556 (N_1556,N_161,In_1384);
and U1557 (N_1557,N_956,In_387);
and U1558 (N_1558,In_1985,N_818);
and U1559 (N_1559,In_445,N_1085);
or U1560 (N_1560,In_1145,N_1138);
or U1561 (N_1561,In_2781,N_862);
and U1562 (N_1562,In_58,N_1086);
nand U1563 (N_1563,In_580,N_877);
and U1564 (N_1564,N_1039,In_2922);
nor U1565 (N_1565,In_2319,In_788);
nor U1566 (N_1566,N_701,In_1438);
nand U1567 (N_1567,In_655,N_7);
or U1568 (N_1568,In_2415,N_231);
and U1569 (N_1569,In_1741,N_543);
or U1570 (N_1570,N_343,N_718);
nand U1571 (N_1571,N_141,N_1079);
or U1572 (N_1572,N_955,In_341);
nand U1573 (N_1573,In_1308,N_638);
or U1574 (N_1574,In_1583,In_1671);
or U1575 (N_1575,In_1311,N_1001);
nor U1576 (N_1576,N_450,In_843);
and U1577 (N_1577,N_562,In_988);
and U1578 (N_1578,N_369,N_112);
nor U1579 (N_1579,In_1203,N_620);
or U1580 (N_1580,N_540,In_1124);
nand U1581 (N_1581,In_1524,N_1124);
or U1582 (N_1582,In_38,In_1804);
or U1583 (N_1583,In_29,N_878);
and U1584 (N_1584,In_25,In_362);
and U1585 (N_1585,N_1142,In_2666);
nor U1586 (N_1586,In_10,N_1158);
or U1587 (N_1587,In_41,In_2958);
and U1588 (N_1588,In_2399,N_572);
nor U1589 (N_1589,N_291,N_442);
nor U1590 (N_1590,In_874,N_724);
nand U1591 (N_1591,In_1703,In_388);
and U1592 (N_1592,N_1017,N_1035);
nor U1593 (N_1593,N_608,N_1152);
nor U1594 (N_1594,In_553,N_444);
and U1595 (N_1595,N_976,N_723);
and U1596 (N_1596,In_279,In_253);
and U1597 (N_1597,In_1765,In_2622);
nand U1598 (N_1598,In_2746,N_1092);
nor U1599 (N_1599,In_1365,N_904);
or U1600 (N_1600,N_518,N_271);
or U1601 (N_1601,N_780,N_1036);
or U1602 (N_1602,In_1173,N_38);
and U1603 (N_1603,N_1120,N_1062);
nor U1604 (N_1604,N_251,In_1976);
nand U1605 (N_1605,N_485,In_1009);
nand U1606 (N_1606,N_789,In_1470);
nand U1607 (N_1607,In_2533,N_657);
or U1608 (N_1608,In_1998,N_621);
nor U1609 (N_1609,In_2900,N_686);
nor U1610 (N_1610,N_367,In_1193);
xor U1611 (N_1611,N_769,N_925);
and U1612 (N_1612,N_893,N_1121);
nand U1613 (N_1613,In_2742,N_806);
and U1614 (N_1614,In_48,N_430);
or U1615 (N_1615,N_1067,In_2380);
nand U1616 (N_1616,N_1107,N_1194);
nor U1617 (N_1617,N_999,N_823);
nor U1618 (N_1618,N_1030,In_833);
nor U1619 (N_1619,In_1286,N_873);
nand U1620 (N_1620,N_1007,In_47);
nor U1621 (N_1621,N_739,In_2475);
nor U1622 (N_1622,N_962,N_883);
or U1623 (N_1623,In_1391,In_1610);
nand U1624 (N_1624,In_2002,N_667);
nand U1625 (N_1625,N_1011,In_1631);
or U1626 (N_1626,N_681,N_645);
and U1627 (N_1627,N_900,N_866);
or U1628 (N_1628,In_1289,In_165);
or U1629 (N_1629,In_2149,N_270);
nor U1630 (N_1630,N_81,N_852);
or U1631 (N_1631,In_804,N_885);
nor U1632 (N_1632,In_1841,N_894);
or U1633 (N_1633,In_732,In_2114);
and U1634 (N_1634,In_1690,In_966);
nor U1635 (N_1635,In_2203,In_1756);
and U1636 (N_1636,N_1132,In_583);
nand U1637 (N_1637,In_2241,N_1076);
xnor U1638 (N_1638,N_821,In_269);
and U1639 (N_1639,N_841,N_240);
nand U1640 (N_1640,N_988,In_602);
and U1641 (N_1641,N_558,In_2411);
and U1642 (N_1642,In_2224,N_1068);
nor U1643 (N_1643,N_868,N_921);
nor U1644 (N_1644,N_786,N_880);
or U1645 (N_1645,In_514,In_1257);
nand U1646 (N_1646,In_2340,In_1622);
nand U1647 (N_1647,N_582,In_365);
xnor U1648 (N_1648,N_456,In_2008);
and U1649 (N_1649,In_121,N_1016);
nand U1650 (N_1650,N_884,N_0);
nand U1651 (N_1651,N_228,In_1827);
or U1652 (N_1652,N_844,In_90);
nor U1653 (N_1653,N_699,N_1150);
nand U1654 (N_1654,N_242,N_938);
and U1655 (N_1655,N_1146,In_2906);
nor U1656 (N_1656,In_116,N_1106);
and U1657 (N_1657,N_664,N_1025);
and U1658 (N_1658,In_1043,N_690);
and U1659 (N_1659,N_705,N_1084);
xor U1660 (N_1660,N_762,In_818);
nor U1661 (N_1661,N_453,In_2550);
nor U1662 (N_1662,N_928,In_1872);
and U1663 (N_1663,N_486,In_2404);
and U1664 (N_1664,N_804,In_2455);
or U1665 (N_1665,In_2018,N_764);
or U1666 (N_1666,In_1968,In_1288);
nor U1667 (N_1667,In_1983,In_2049);
nand U1668 (N_1668,N_899,N_994);
nor U1669 (N_1669,In_1095,In_1035);
and U1670 (N_1670,In_2031,N_1070);
nand U1671 (N_1671,In_2557,N_647);
nor U1672 (N_1672,In_2899,In_497);
nand U1673 (N_1673,N_887,N_1155);
nand U1674 (N_1674,N_965,In_1416);
nor U1675 (N_1675,In_2813,In_374);
or U1676 (N_1676,In_904,In_1750);
nand U1677 (N_1677,N_763,N_421);
or U1678 (N_1678,In_350,N_672);
nor U1679 (N_1679,N_159,In_1594);
or U1680 (N_1680,N_1013,In_2102);
nor U1681 (N_1681,N_1144,N_1197);
or U1682 (N_1682,In_594,In_396);
nand U1683 (N_1683,In_2837,In_334);
nand U1684 (N_1684,In_1884,N_265);
nor U1685 (N_1685,In_446,In_1723);
nand U1686 (N_1686,In_2614,N_711);
nor U1687 (N_1687,N_411,N_674);
nand U1688 (N_1688,N_932,In_2227);
nand U1689 (N_1689,In_2131,In_1568);
nor U1690 (N_1690,N_1171,In_2974);
or U1691 (N_1691,In_2229,In_2150);
nor U1692 (N_1692,In_1707,N_615);
nor U1693 (N_1693,N_1043,N_788);
nor U1694 (N_1694,In_949,In_675);
nor U1695 (N_1695,N_616,In_2688);
nor U1696 (N_1696,In_2268,N_682);
nand U1697 (N_1697,N_767,N_835);
nor U1698 (N_1698,N_23,In_453);
and U1699 (N_1699,In_1272,N_697);
nor U1700 (N_1700,N_712,In_256);
nor U1701 (N_1701,In_2543,In_1221);
nand U1702 (N_1702,N_61,N_479);
nor U1703 (N_1703,In_2769,N_544);
or U1704 (N_1704,In_1412,In_2275);
nand U1705 (N_1705,N_772,N_646);
nor U1706 (N_1706,N_1088,In_1092);
nand U1707 (N_1707,N_735,In_13);
or U1708 (N_1708,In_2050,In_562);
or U1709 (N_1709,N_934,In_103);
or U1710 (N_1710,N_565,In_1714);
nand U1711 (N_1711,N_186,N_872);
and U1712 (N_1712,In_2851,N_511);
nor U1713 (N_1713,N_1178,N_1193);
nor U1714 (N_1714,N_1047,N_390);
and U1715 (N_1715,N_795,N_1048);
and U1716 (N_1716,In_2749,N_399);
and U1717 (N_1717,N_515,N_107);
and U1718 (N_1718,N_1180,In_2266);
nand U1719 (N_1719,In_1407,In_2473);
and U1720 (N_1720,N_740,In_886);
and U1721 (N_1721,N_875,In_2831);
nor U1722 (N_1722,N_87,N_315);
and U1723 (N_1723,N_259,N_741);
nand U1724 (N_1724,In_2322,In_919);
or U1725 (N_1725,N_1181,N_709);
nor U1726 (N_1726,N_1184,N_360);
nand U1727 (N_1727,N_801,N_263);
nor U1728 (N_1728,N_192,In_475);
and U1729 (N_1729,N_933,In_1814);
nor U1730 (N_1730,In_1862,In_1514);
nand U1731 (N_1731,N_869,N_1054);
nor U1732 (N_1732,In_1185,In_1665);
and U1733 (N_1733,In_1410,In_2975);
nor U1734 (N_1734,In_1870,In_126);
and U1735 (N_1735,In_1997,N_774);
and U1736 (N_1736,In_1273,N_902);
nor U1737 (N_1737,N_716,In_2139);
nand U1738 (N_1738,N_1080,In_294);
nand U1739 (N_1739,In_306,N_1087);
xnor U1740 (N_1740,N_1169,N_1145);
or U1741 (N_1741,N_449,N_1041);
nand U1742 (N_1742,N_673,N_986);
nor U1743 (N_1743,In_1025,In_414);
or U1744 (N_1744,N_886,In_1846);
or U1745 (N_1745,In_1505,In_2790);
or U1746 (N_1746,N_537,In_1348);
nor U1747 (N_1747,N_1093,N_829);
nor U1748 (N_1748,N_1147,N_923);
or U1749 (N_1749,N_179,In_207);
nand U1750 (N_1750,In_1325,N_969);
nor U1751 (N_1751,In_1900,In_2132);
nand U1752 (N_1752,In_2281,In_2325);
and U1753 (N_1753,N_695,In_1360);
or U1754 (N_1754,N_629,In_1395);
nand U1755 (N_1755,N_164,In_1216);
nor U1756 (N_1756,N_99,N_69);
nor U1757 (N_1757,In_2320,In_2095);
or U1758 (N_1758,N_706,In_906);
nand U1759 (N_1759,In_2385,In_2559);
nand U1760 (N_1760,N_624,N_622);
or U1761 (N_1761,N_303,In_98);
and U1762 (N_1762,N_128,In_1270);
or U1763 (N_1763,In_2483,N_97);
nand U1764 (N_1764,In_2808,In_1205);
and U1765 (N_1765,In_1489,N_194);
or U1766 (N_1766,In_2664,In_1319);
nand U1767 (N_1767,In_1938,In_2862);
nor U1768 (N_1768,In_2127,N_1073);
nand U1769 (N_1769,In_1338,N_753);
and U1770 (N_1770,In_946,N_285);
and U1771 (N_1771,In_2757,N_912);
and U1772 (N_1772,N_754,In_167);
and U1773 (N_1773,N_1000,N_443);
nand U1774 (N_1774,N_181,N_1137);
nand U1775 (N_1775,In_720,N_642);
and U1776 (N_1776,In_2689,N_1100);
or U1777 (N_1777,N_1140,In_1012);
nand U1778 (N_1778,N_96,In_637);
nand U1779 (N_1779,N_1113,In_1465);
or U1780 (N_1780,N_103,N_198);
and U1781 (N_1781,N_848,N_671);
nor U1782 (N_1782,N_668,In_1071);
or U1783 (N_1783,In_2613,N_480);
and U1784 (N_1784,In_1587,In_2096);
xnor U1785 (N_1785,In_2716,In_2414);
and U1786 (N_1786,In_285,In_2402);
nor U1787 (N_1787,N_351,In_2423);
and U1788 (N_1788,N_863,N_989);
or U1789 (N_1789,N_606,In_1299);
nand U1790 (N_1790,In_1296,N_708);
nor U1791 (N_1791,In_1374,In_270);
and U1792 (N_1792,In_918,In_2310);
and U1793 (N_1793,In_1606,In_2785);
and U1794 (N_1794,N_836,N_931);
nand U1795 (N_1795,In_696,In_1982);
or U1796 (N_1796,In_100,N_8);
nor U1797 (N_1797,N_244,In_698);
nand U1798 (N_1798,N_58,N_458);
and U1799 (N_1799,In_1617,In_1803);
and U1800 (N_1800,In_2927,In_1136);
nor U1801 (N_1801,In_1633,N_1108);
and U1802 (N_1802,In_1806,N_807);
nor U1803 (N_1803,N_1286,In_2212);
or U1804 (N_1804,N_1253,N_1465);
or U1805 (N_1805,N_997,N_1467);
nor U1806 (N_1806,N_1348,N_1208);
nand U1807 (N_1807,N_1674,In_2342);
nor U1808 (N_1808,In_2165,N_1700);
nor U1809 (N_1809,N_1769,N_440);
nor U1810 (N_1810,N_611,N_1210);
or U1811 (N_1811,N_1709,In_2074);
nand U1812 (N_1812,N_319,N_1214);
nand U1813 (N_1813,N_1670,N_618);
and U1814 (N_1814,N_1767,In_2541);
or U1815 (N_1815,In_2991,In_2830);
and U1816 (N_1816,In_235,N_732);
and U1817 (N_1817,In_252,In_572);
xnor U1818 (N_1818,N_796,N_1689);
or U1819 (N_1819,N_556,In_1413);
and U1820 (N_1820,N_1527,In_2914);
or U1821 (N_1821,N_648,N_834);
and U1822 (N_1822,In_1934,N_936);
and U1823 (N_1823,N_1282,N_1632);
and U1824 (N_1824,N_1365,N_794);
nor U1825 (N_1825,In_1455,N_627);
or U1826 (N_1826,N_1114,N_1346);
nor U1827 (N_1827,N_1622,N_1378);
nor U1828 (N_1828,N_1203,N_1401);
and U1829 (N_1829,N_1446,N_267);
or U1830 (N_1830,In_2759,N_905);
and U1831 (N_1831,In_2739,In_2463);
nand U1832 (N_1832,N_604,N_1305);
nor U1833 (N_1833,N_1718,N_1326);
nor U1834 (N_1834,N_1560,N_1620);
nand U1835 (N_1835,N_1466,N_1233);
xnor U1836 (N_1836,N_1422,N_1349);
nor U1837 (N_1837,N_1059,N_665);
and U1838 (N_1838,In_2155,N_659);
or U1839 (N_1839,In_1172,In_145);
or U1840 (N_1840,N_913,In_588);
and U1841 (N_1841,In_385,N_1134);
nand U1842 (N_1842,N_1212,N_1524);
or U1843 (N_1843,N_1491,In_2374);
nor U1844 (N_1844,N_517,In_2357);
or U1845 (N_1845,N_1631,In_1802);
nand U1846 (N_1846,In_2396,In_257);
or U1847 (N_1847,N_790,In_630);
and U1848 (N_1848,N_333,N_1673);
nor U1849 (N_1849,In_2701,In_1433);
nor U1850 (N_1850,N_346,N_924);
nor U1851 (N_1851,N_1010,N_1458);
nand U1852 (N_1852,N_1473,In_703);
xnor U1853 (N_1853,In_2252,In_1850);
nor U1854 (N_1854,In_2343,N_1414);
nor U1855 (N_1855,In_485,N_1575);
nor U1856 (N_1856,N_1695,N_1245);
nor U1857 (N_1857,N_601,N_1512);
nor U1858 (N_1858,N_1333,N_13);
or U1859 (N_1859,N_1482,N_1211);
nor U1860 (N_1860,In_620,N_470);
xnor U1861 (N_1861,N_1545,N_1161);
and U1862 (N_1862,N_1431,N_1584);
and U1863 (N_1863,In_1939,N_770);
or U1864 (N_1864,N_1321,N_1724);
and U1865 (N_1865,In_177,N_755);
nor U1866 (N_1866,N_1418,N_983);
or U1867 (N_1867,In_2595,N_944);
and U1868 (N_1868,N_1307,N_1633);
and U1869 (N_1869,N_1763,N_1383);
nor U1870 (N_1870,N_1582,N_1509);
and U1871 (N_1871,N_1705,In_131);
nand U1872 (N_1872,N_1372,N_1683);
nand U1873 (N_1873,N_1565,In_1699);
nor U1874 (N_1874,N_1439,In_2003);
and U1875 (N_1875,N_290,N_1639);
or U1876 (N_1876,In_1318,In_690);
or U1877 (N_1877,N_199,In_1028);
nand U1878 (N_1878,In_1808,N_146);
or U1879 (N_1879,N_1313,N_1519);
nor U1880 (N_1880,N_1755,N_1520);
nand U1881 (N_1881,N_1135,N_1630);
xor U1882 (N_1882,N_1597,N_1487);
nand U1883 (N_1883,In_607,In_378);
or U1884 (N_1884,In_2799,N_1347);
nand U1885 (N_1885,N_1112,N_1736);
nor U1886 (N_1886,In_1608,N_1738);
and U1887 (N_1887,N_843,N_1250);
nand U1888 (N_1888,N_174,N_688);
nor U1889 (N_1889,N_1259,N_504);
nand U1890 (N_1890,N_1793,N_1766);
and U1891 (N_1891,In_2246,In_1368);
nand U1892 (N_1892,In_1902,In_2920);
and U1893 (N_1893,N_1266,N_1412);
nand U1894 (N_1894,N_1646,N_1280);
nand U1895 (N_1895,N_202,N_1296);
or U1896 (N_1896,N_1213,In_1659);
and U1897 (N_1897,N_1562,N_330);
or U1898 (N_1898,N_1580,N_1765);
nor U1899 (N_1899,N_26,N_335);
nor U1900 (N_1900,N_1660,In_929);
nand U1901 (N_1901,N_1363,In_2786);
nor U1902 (N_1902,N_1251,In_2493);
and U1903 (N_1903,N_1662,In_1874);
nand U1904 (N_1904,N_1623,N_1111);
or U1905 (N_1905,N_1289,N_1770);
and U1906 (N_1906,N_1514,N_1248);
nand U1907 (N_1907,N_1706,N_1627);
nor U1908 (N_1908,N_110,N_1375);
nor U1909 (N_1909,N_675,N_1456);
or U1910 (N_1910,In_2909,N_134);
nor U1911 (N_1911,N_1621,N_1475);
xor U1912 (N_1912,N_1547,N_579);
nand U1913 (N_1913,N_1074,N_1471);
nand U1914 (N_1914,N_1315,N_1484);
nor U1915 (N_1915,N_1409,N_1419);
nand U1916 (N_1916,N_1595,N_1201);
and U1917 (N_1917,N_90,In_1632);
or U1918 (N_1918,In_1251,N_208);
nand U1919 (N_1919,N_702,N_1583);
or U1920 (N_1920,In_1004,In_1769);
and U1921 (N_1921,In_1195,N_1534);
nor U1922 (N_1922,In_852,In_1332);
or U1923 (N_1923,N_949,N_1402);
or U1924 (N_1924,N_1436,N_1243);
nor U1925 (N_1925,In_1864,N_1200);
nor U1926 (N_1926,N_1264,N_139);
nand U1927 (N_1927,N_193,N_1273);
and U1928 (N_1928,N_1703,In_1304);
and U1929 (N_1929,N_1274,N_854);
nor U1930 (N_1930,N_1198,N_398);
nand U1931 (N_1931,In_2119,N_1672);
or U1932 (N_1932,N_1784,N_636);
or U1933 (N_1933,In_161,N_1607);
nor U1934 (N_1934,In_1616,N_1693);
or U1935 (N_1935,N_1617,N_1782);
xor U1936 (N_1936,N_1285,N_1711);
and U1937 (N_1937,N_1218,N_1712);
or U1938 (N_1938,N_1408,N_1608);
nand U1939 (N_1939,N_1265,N_1556);
nor U1940 (N_1940,N_1024,N_918);
nor U1941 (N_1941,N_1302,N_1576);
and U1942 (N_1942,In_753,N_1272);
nor U1943 (N_1943,N_1379,N_1792);
and U1944 (N_1944,N_1344,N_630);
nor U1945 (N_1945,N_1551,N_973);
nand U1946 (N_1946,In_1817,N_1410);
or U1947 (N_1947,In_1302,N_602);
nand U1948 (N_1948,N_1444,N_1154);
nor U1949 (N_1949,In_964,In_1376);
nand U1950 (N_1950,N_1327,N_1303);
and U1951 (N_1951,N_311,In_785);
nor U1952 (N_1952,In_401,N_980);
xnor U1953 (N_1953,N_1744,N_143);
or U1954 (N_1954,N_1681,N_417);
or U1955 (N_1955,N_1521,N_1548);
nand U1956 (N_1956,N_1587,N_730);
or U1957 (N_1957,In_1006,N_1677);
or U1958 (N_1958,In_1812,In_273);
or U1959 (N_1959,N_1748,In_1246);
nor U1960 (N_1960,N_1495,N_948);
xnor U1961 (N_1961,N_1745,N_1377);
nor U1962 (N_1962,In_1477,N_1564);
and U1963 (N_1963,N_1710,N_1641);
or U1964 (N_1964,N_1715,In_2699);
or U1965 (N_1965,N_577,N_1329);
nor U1966 (N_1966,In_267,In_1883);
or U1967 (N_1967,N_1612,N_1666);
nand U1968 (N_1968,N_1470,N_1702);
and U1969 (N_1969,N_207,N_478);
or U1970 (N_1970,N_1295,In_1381);
nor U1971 (N_1971,N_888,N_1225);
nor U1972 (N_1972,N_1653,N_1581);
or U1973 (N_1973,N_1109,In_1620);
xnor U1974 (N_1974,N_856,N_803);
and U1975 (N_1975,In_542,In_1261);
nor U1976 (N_1976,In_2250,In_1562);
nor U1977 (N_1977,N_831,N_781);
or U1978 (N_1978,In_1234,In_1352);
nor U1979 (N_1979,N_748,N_1382);
nand U1980 (N_1980,N_1506,N_987);
or U1981 (N_1981,N_1242,In_1121);
or U1982 (N_1982,N_1014,N_1386);
nor U1983 (N_1983,N_1341,N_898);
or U1984 (N_1984,In_1114,In_1091);
nor U1985 (N_1985,N_1215,N_1649);
or U1986 (N_1986,N_827,N_1668);
xor U1987 (N_1987,N_1256,N_1433);
nand U1988 (N_1988,N_1513,N_1448);
or U1989 (N_1989,N_1246,In_437);
and U1990 (N_1990,N_206,N_249);
and U1991 (N_1991,N_1552,In_1473);
and U1992 (N_1992,N_1063,N_722);
nand U1993 (N_1993,N_1361,In_1408);
or U1994 (N_1994,In_2803,N_1761);
nand U1995 (N_1995,N_412,N_635);
nand U1996 (N_1996,N_1515,N_1542);
nor U1997 (N_1997,N_1671,N_1421);
and U1998 (N_1998,N_342,In_2617);
nor U1999 (N_1999,N_1789,In_1409);
and U2000 (N_2000,N_1247,N_378);
or U2001 (N_2001,N_1783,N_1790);
and U2002 (N_2002,N_1526,N_1091);
or U2003 (N_2003,In_2213,N_1616);
and U2004 (N_2004,N_1481,N_1566);
nand U2005 (N_2005,In_827,In_2512);
and U2006 (N_2006,N_1538,In_540);
and U2007 (N_2007,N_1701,In_2051);
and U2008 (N_2008,N_963,N_1260);
and U2009 (N_2009,In_1297,N_1486);
or U2010 (N_2010,N_1376,N_1311);
nor U2011 (N_2011,In_317,N_1717);
nand U2012 (N_2012,In_2356,N_639);
xnor U2013 (N_2013,N_991,N_1730);
nor U2014 (N_2014,N_560,N_1636);
or U2015 (N_2015,N_1126,N_746);
or U2016 (N_2016,In_2669,N_874);
nor U2017 (N_2017,In_494,N_1304);
nor U2018 (N_2018,N_995,N_1480);
and U2019 (N_2019,N_766,N_1293);
or U2020 (N_2020,In_8,N_371);
or U2021 (N_2021,N_981,N_1428);
nor U2022 (N_2022,In_932,N_1032);
or U2023 (N_2023,In_2389,In_2219);
nand U2024 (N_2024,In_2428,In_2878);
and U2025 (N_2025,N_1772,In_2020);
nand U2026 (N_2026,In_380,N_1268);
or U2027 (N_2027,In_34,In_1039);
and U2028 (N_2028,N_1751,N_1535);
and U2029 (N_2029,N_1544,N_1479);
or U2030 (N_2030,N_1734,N_1033);
nand U2031 (N_2031,N_1604,N_1397);
nand U2032 (N_2032,In_930,N_165);
nor U2033 (N_2033,N_1232,N_882);
or U2034 (N_2034,N_481,In_2488);
nor U2035 (N_2035,In_2253,In_704);
and U2036 (N_2036,N_1308,N_1523);
nand U2037 (N_2037,In_819,N_1452);
and U2038 (N_2038,N_1600,N_1432);
or U2039 (N_2039,N_677,N_1721);
or U2040 (N_2040,N_1787,N_1531);
nor U2041 (N_2041,N_729,In_604);
nand U2042 (N_2042,In_2641,In_2258);
nand U2043 (N_2043,N_610,N_1577);
or U2044 (N_2044,N_1469,N_1442);
nor U2045 (N_2045,N_1640,In_2547);
or U2046 (N_2046,N_1395,N_1425);
and U2047 (N_2047,N_1223,N_833);
and U2048 (N_2048,N_1072,N_1186);
nor U2049 (N_2049,In_1792,N_1796);
nor U2050 (N_2050,N_1360,N_1490);
nand U2051 (N_2051,N_1602,In_2405);
nand U2052 (N_2052,N_870,N_1065);
or U2053 (N_2053,N_1656,N_1380);
nand U2054 (N_2054,In_353,In_647);
nand U2055 (N_2055,N_1316,N_1429);
and U2056 (N_2056,N_1511,N_1244);
or U2057 (N_2057,N_1461,N_324);
nor U2058 (N_2058,N_264,N_1405);
nor U2059 (N_2059,N_698,N_1550);
and U2060 (N_2060,N_1638,N_176);
or U2061 (N_2061,In_189,N_215);
and U2062 (N_2062,N_1510,N_1619);
and U2063 (N_2063,N_1393,In_2403);
nand U2064 (N_2064,In_2639,N_1559);
nand U2065 (N_2065,N_1392,N_109);
nand U2066 (N_2066,N_1438,N_917);
or U2067 (N_2067,In_2951,In_2672);
xor U2068 (N_2068,In_952,N_526);
nand U2069 (N_2069,N_749,N_51);
and U2070 (N_2070,N_209,N_808);
nand U2071 (N_2071,N_1650,In_659);
or U2072 (N_2072,N_1235,N_1325);
nand U2073 (N_2073,N_1328,N_1799);
or U2074 (N_2074,N_1455,N_1635);
nor U2075 (N_2075,In_724,In_2529);
nor U2076 (N_2076,In_914,N_1269);
nor U2077 (N_2077,N_1571,N_1685);
and U2078 (N_2078,N_1306,In_716);
or U2079 (N_2079,N_1603,N_1271);
or U2080 (N_2080,N_1779,N_1477);
nand U2081 (N_2081,In_1330,In_227);
or U2082 (N_2082,N_28,N_1555);
nand U2083 (N_2083,N_1493,N_1217);
nor U2084 (N_2084,N_1119,N_1719);
nor U2085 (N_2085,In_2337,N_1504);
and U2086 (N_2086,N_1502,N_1454);
or U2087 (N_2087,N_32,N_233);
and U2088 (N_2088,N_1609,N_1658);
and U2089 (N_2089,In_1474,N_941);
nor U2090 (N_2090,N_972,N_1774);
and U2091 (N_2091,N_364,N_1115);
nor U2092 (N_2092,N_1240,N_1435);
and U2093 (N_2093,In_2720,In_1183);
xnor U2094 (N_2094,N_1732,N_728);
or U2095 (N_2095,N_649,In_2801);
or U2096 (N_2096,In_1730,In_2822);
nor U2097 (N_2097,N_982,N_1680);
nand U2098 (N_2098,N_1747,In_2539);
and U2099 (N_2099,N_1398,N_317);
nor U2100 (N_2100,In_1083,N_1457);
nand U2101 (N_2101,N_1497,N_1390);
or U2102 (N_2102,N_1056,In_2939);
and U2103 (N_2103,N_1601,N_641);
and U2104 (N_2104,In_2123,N_154);
or U2105 (N_2105,N_1292,N_1518);
and U2106 (N_2106,N_687,N_1567);
nor U2107 (N_2107,In_338,N_1340);
and U2108 (N_2108,N_1537,N_162);
and U2109 (N_2109,N_1310,N_607);
or U2110 (N_2110,N_1498,In_46);
nor U2111 (N_2111,N_309,In_421);
nand U2112 (N_2112,N_1427,N_1420);
nand U2113 (N_2113,N_1794,In_2537);
or U2114 (N_2114,N_1207,N_1536);
and U2115 (N_2115,N_1777,N_1553);
or U2116 (N_2116,N_1532,N_890);
nand U2117 (N_2117,N_1221,In_2767);
nor U2118 (N_2118,N_1355,In_1816);
or U2119 (N_2119,In_153,N_1643);
nand U2120 (N_2120,N_349,N_1543);
nor U2121 (N_2121,N_1021,N_1483);
nand U2122 (N_2122,N_820,N_1023);
nand U2123 (N_2123,N_676,N_1591);
and U2124 (N_2124,N_1499,In_2240);
or U2125 (N_2125,N_1399,In_2075);
nand U2126 (N_2126,In_2835,In_905);
nand U2127 (N_2127,N_1728,N_147);
nor U2128 (N_2128,N_382,N_322);
nand U2129 (N_2129,N_1222,N_1319);
nand U2130 (N_2130,N_1356,N_1262);
nand U2131 (N_2131,In_2870,N_584);
nand U2132 (N_2132,In_327,N_138);
nor U2133 (N_2133,N_1417,N_301);
or U2134 (N_2134,In_2148,N_1163);
nor U2135 (N_2135,N_1505,N_1659);
nor U2136 (N_2136,N_1239,N_1764);
or U2137 (N_2137,N_1366,N_1219);
and U2138 (N_2138,N_692,In_888);
and U2139 (N_2139,N_1746,N_1160);
and U2140 (N_2140,N_1585,N_1644);
nor U2141 (N_2141,N_427,N_725);
or U2142 (N_2142,In_2507,N_1230);
and U2143 (N_2143,N_1270,N_704);
nor U2144 (N_2144,N_1374,In_727);
and U2145 (N_2145,N_446,N_1367);
xnor U2146 (N_2146,N_1324,N_1387);
nor U2147 (N_2147,N_1596,N_857);
or U2148 (N_2148,N_1593,N_1426);
or U2149 (N_2149,In_677,N_1057);
nand U2150 (N_2150,N_626,N_947);
and U2151 (N_2151,N_1275,N_1578);
nor U2152 (N_2152,N_1151,N_1731);
and U2153 (N_2153,N_1234,N_1637);
nor U2154 (N_2154,N_1508,In_2109);
nand U2155 (N_2155,In_1099,N_1798);
nor U2156 (N_2156,N_1384,N_1773);
and U2157 (N_2157,N_1572,In_2645);
nand U2158 (N_2158,N_1750,N_1231);
nor U2159 (N_2159,N_1753,In_2211);
or U2160 (N_2160,N_802,N_1141);
nand U2161 (N_2161,N_1574,In_781);
nor U2162 (N_2162,In_692,In_1290);
nand U2163 (N_2163,N_1615,N_1205);
or U2164 (N_2164,N_1533,N_1411);
nor U2165 (N_2165,N_1173,N_951);
and U2166 (N_2166,N_94,N_1723);
or U2167 (N_2167,N_1688,N_1451);
xor U2168 (N_2168,In_661,N_241);
and U2169 (N_2169,N_1441,N_375);
nand U2170 (N_2170,N_1778,N_1729);
nor U2171 (N_2171,N_652,N_1118);
nand U2172 (N_2172,N_1279,In_2421);
and U2173 (N_2173,N_1759,N_1733);
or U2174 (N_2174,N_1450,N_1391);
nor U2175 (N_2175,N_1592,N_1665);
or U2176 (N_2176,N_1117,N_1737);
and U2177 (N_2177,In_2047,In_1036);
or U2178 (N_2178,N_180,N_1561);
and U2179 (N_2179,N_879,N_1704);
nor U2180 (N_2180,N_1447,N_1460);
and U2181 (N_2181,N_1237,N_1558);
and U2182 (N_2182,In_1402,N_45);
nor U2183 (N_2183,In_1242,N_1071);
or U2184 (N_2184,N_1227,In_2929);
nor U2185 (N_2185,N_1464,In_2360);
nand U2186 (N_2186,N_415,N_1624);
and U2187 (N_2187,In_2583,N_1202);
or U2188 (N_2188,In_305,N_294);
nand U2189 (N_2189,N_977,In_55);
and U2190 (N_2190,N_1618,In_931);
or U2191 (N_2191,N_1338,In_1729);
or U2192 (N_2192,N_876,N_798);
and U2193 (N_2193,In_1650,In_1044);
and U2194 (N_2194,N_1336,N_1281);
and U2195 (N_2195,N_1357,N_145);
or U2196 (N_2196,N_1756,N_1209);
and U2197 (N_2197,N_1795,N_892);
or U2198 (N_2198,In_1737,N_1517);
nand U2199 (N_2199,N_1220,N_1170);
nor U2200 (N_2200,N_1176,N_970);
or U2201 (N_2201,In_2566,N_1320);
nand U2202 (N_2202,N_1351,In_2791);
nor U2203 (N_2203,N_1786,In_2642);
nor U2204 (N_2204,N_1406,N_1507);
or U2205 (N_2205,In_800,N_1687);
nor U2206 (N_2206,N_612,N_1546);
nor U2207 (N_2207,N_1468,N_1768);
and U2208 (N_2208,N_1478,In_102);
nand U2209 (N_2209,In_1654,N_1678);
and U2210 (N_2210,N_1463,N_1740);
nor U2211 (N_2211,N_1686,In_1176);
and U2212 (N_2212,In_2612,N_1089);
nand U2213 (N_2213,N_1727,N_1522);
or U2214 (N_2214,N_200,In_346);
and U2215 (N_2215,N_640,N_1573);
and U2216 (N_2216,In_2807,N_1400);
and U2217 (N_2217,In_829,N_858);
or U2218 (N_2218,N_1015,N_758);
and U2219 (N_2219,N_1754,In_566);
or U2220 (N_2220,N_1277,N_1453);
and U2221 (N_2221,N_1699,N_1654);
and U2222 (N_2222,N_787,In_2609);
and U2223 (N_2223,N_1300,N_310);
and U2224 (N_2224,N_1492,N_1404);
and U2225 (N_2225,N_1528,In_2814);
and U2226 (N_2226,N_1050,N_979);
nor U2227 (N_2227,In_1754,N_1791);
nand U2228 (N_2228,N_1647,N_1667);
nor U2229 (N_2229,N_1350,N_1388);
or U2230 (N_2230,In_908,N_98);
nand U2231 (N_2231,In_587,N_1330);
nand U2232 (N_2232,N_1570,In_2978);
and U2233 (N_2233,N_1489,N_1440);
and U2234 (N_2234,N_1651,N_1675);
nand U2235 (N_2235,N_372,In_2086);
nand U2236 (N_2236,N_1309,In_1218);
and U2237 (N_2237,In_2338,N_190);
and U2238 (N_2238,N_1634,In_408);
nand U2239 (N_2239,N_1339,N_1381);
nor U2240 (N_2240,N_1625,N_1394);
or U2241 (N_2241,N_1004,N_1642);
and U2242 (N_2242,N_1669,N_1216);
or U2243 (N_2243,N_1136,N_1288);
or U2244 (N_2244,N_1462,N_742);
or U2245 (N_2245,In_1581,N_1317);
and U2246 (N_2246,N_1599,N_1541);
nand U2247 (N_2247,N_662,N_1598);
or U2248 (N_2248,N_1735,N_1629);
and U2249 (N_2249,In_1852,N_1278);
nor U2250 (N_2250,In_742,In_2368);
nand U2251 (N_2251,N_471,N_1396);
nand U2252 (N_2252,N_1226,N_1252);
nand U2253 (N_2253,N_1720,N_1771);
nand U2254 (N_2254,N_483,In_1460);
nor U2255 (N_2255,N_1716,N_1263);
nand U2256 (N_2256,N_1708,N_1722);
nand U2257 (N_2257,In_1890,N_1563);
and U2258 (N_2258,N_1757,N_1149);
nor U2259 (N_2259,N_1116,In_1208);
or U2260 (N_2260,N_1415,N_1525);
nor U2261 (N_2261,N_1371,In_2826);
nand U2262 (N_2262,N_1776,N_908);
and U2263 (N_2263,N_713,N_1496);
nand U2264 (N_2264,N_1362,In_1787);
nand U2265 (N_2265,In_1431,N_733);
and U2266 (N_2266,N_1474,N_1472);
and U2267 (N_2267,N_1077,N_566);
nor U2268 (N_2268,N_1322,N_1423);
or U2269 (N_2269,N_1254,N_1314);
or U2270 (N_2270,N_1788,N_1443);
and U2271 (N_2271,N_1610,N_1131);
and U2272 (N_2272,N_1529,N_1368);
or U2273 (N_2273,N_1060,In_1774);
or U2274 (N_2274,In_814,N_1290);
nor U2275 (N_2275,N_1694,In_1115);
nor U2276 (N_2276,N_1605,In_463);
or U2277 (N_2277,N_1103,N_1258);
and U2278 (N_2278,N_1488,N_1449);
or U2279 (N_2279,N_356,N_1554);
or U2280 (N_2280,N_1679,In_226);
nor U2281 (N_2281,N_276,In_251);
nand U2282 (N_2282,In_1016,N_1590);
and U2283 (N_2283,N_1501,N_1445);
nand U2284 (N_2284,In_811,N_1283);
and U2285 (N_2285,N_1516,N_678);
nor U2286 (N_2286,N_1569,N_1298);
or U2287 (N_2287,N_1204,N_1684);
and U2288 (N_2288,N_1318,N_1332);
and U2289 (N_2289,In_57,N_35);
or U2290 (N_2290,N_1284,In_1522);
nor U2291 (N_2291,In_2459,In_1491);
or U2292 (N_2292,N_1267,N_1682);
and U2293 (N_2293,N_1334,In_941);
nor U2294 (N_2294,N_1190,N_1287);
nor U2295 (N_2295,N_737,N_1628);
or U2296 (N_2296,In_32,N_1714);
and U2297 (N_2297,In_610,N_1255);
xnor U2298 (N_2298,N_1698,In_1576);
and U2299 (N_2299,N_776,In_1975);
and U2300 (N_2300,In_1876,N_1437);
nand U2301 (N_2301,In_1499,N_1760);
and U2302 (N_2302,N_201,N_760);
nand U2303 (N_2303,N_891,N_830);
nor U2304 (N_2304,N_1343,N_1323);
nor U2305 (N_2305,N_1206,N_1780);
or U2306 (N_2306,N_791,N_1540);
nand U2307 (N_2307,N_1241,N_1485);
or U2308 (N_2308,In_725,N_1385);
nor U2309 (N_2309,N_1416,N_1785);
nor U2310 (N_2310,N_1589,N_1261);
xnor U2311 (N_2311,N_935,N_1312);
nand U2312 (N_2312,N_559,In_2218);
or U2313 (N_2313,N_1353,N_1781);
and U2314 (N_2314,In_2715,N_1707);
nand U2315 (N_2315,N_1749,N_1228);
nand U2316 (N_2316,N_1294,In_2819);
xnor U2317 (N_2317,N_628,N_508);
or U2318 (N_2318,In_2427,N_1726);
nor U2319 (N_2319,N_1664,In_634);
nor U2320 (N_2320,N_1122,N_1594);
and U2321 (N_2321,N_1549,N_1331);
nor U2322 (N_2322,N_1249,N_1557);
nand U2323 (N_2323,N_247,N_36);
and U2324 (N_2324,N_1797,N_1500);
nor U2325 (N_2325,N_603,In_2422);
nand U2326 (N_2326,N_1645,In_2489);
or U2327 (N_2327,N_33,N_1713);
or U2328 (N_2328,In_1577,In_1719);
and U2329 (N_2329,In_2425,In_531);
and U2330 (N_2330,In_920,N_1345);
or U2331 (N_2331,N_494,N_1335);
and U2332 (N_2332,In_593,N_750);
nor U2333 (N_2333,N_1337,In_2538);
and U2334 (N_2334,N_1185,N_1655);
nand U2335 (N_2335,In_1885,N_985);
and U2336 (N_2336,N_1182,N_1098);
or U2337 (N_2337,N_1156,In_2965);
nor U2338 (N_2338,N_1661,N_840);
or U2339 (N_2339,N_1359,N_853);
and U2340 (N_2340,N_1012,In_1415);
or U2341 (N_2341,N_861,N_1236);
and U2342 (N_2342,In_2887,N_1692);
nor U2343 (N_2343,N_1648,N_1606);
or U2344 (N_2344,N_1291,N_1352);
and U2345 (N_2345,N_1301,N_1775);
or U2346 (N_2346,N_715,N_1229);
nand U2347 (N_2347,N_216,In_2296);
xor U2348 (N_2348,N_1125,N_911);
or U2349 (N_2349,N_1027,N_573);
or U2350 (N_2350,N_744,In_2983);
xnor U2351 (N_2351,In_2440,N_1407);
and U2352 (N_2352,N_1224,In_1593);
nor U2353 (N_2353,N_783,N_1434);
or U2354 (N_2354,In_2570,In_2637);
and U2355 (N_2355,N_1373,N_1276);
nand U2356 (N_2356,N_1568,In_2773);
nand U2357 (N_2357,N_1413,N_1690);
nor U2358 (N_2358,N_1752,N_689);
or U2359 (N_2359,In_1291,N_1530);
nand U2360 (N_2360,N_1403,N_1579);
and U2361 (N_2361,N_1725,N_926);
xor U2362 (N_2362,N_1257,N_1143);
and U2363 (N_2363,In_2397,N_14);
nor U2364 (N_2364,N_1424,In_2585);
nor U2365 (N_2365,N_1195,N_379);
and U2366 (N_2366,In_512,In_1422);
nand U2367 (N_2367,N_1696,N_144);
and U2368 (N_2368,N_1613,N_1364);
and U2369 (N_2369,In_1023,N_1494);
or U2370 (N_2370,N_1758,N_1238);
or U2371 (N_2371,In_1647,N_1297);
or U2372 (N_2372,N_1503,N_1743);
nor U2373 (N_2373,N_800,N_1370);
nand U2374 (N_2374,N_1342,N_1586);
and U2375 (N_2375,N_1002,In_2174);
nor U2376 (N_2376,N_1742,N_939);
nand U2377 (N_2377,N_1177,In_959);
and U2378 (N_2378,N_1676,In_382);
and U2379 (N_2379,N_1697,In_1236);
nor U2380 (N_2380,N_1626,N_492);
nor U2381 (N_2381,N_1691,N_1164);
or U2382 (N_2382,N_1369,N_1741);
or U2383 (N_2383,In_1445,In_1658);
nand U2384 (N_2384,In_1854,N_1476);
nor U2385 (N_2385,N_229,N_1539);
nand U2386 (N_2386,N_416,N_1099);
or U2387 (N_2387,N_1588,In_517);
or U2388 (N_2388,N_693,N_1299);
nand U2389 (N_2389,N_1657,N_1459);
and U2390 (N_2390,N_1614,In_1495);
or U2391 (N_2391,N_978,N_1354);
nor U2392 (N_2392,N_1389,In_316);
and U2393 (N_2393,In_2763,In_1181);
nor U2394 (N_2394,N_1739,N_906);
or U2395 (N_2395,N_1652,N_1358);
nand U2396 (N_2396,N_114,In_1772);
nor U2397 (N_2397,N_1762,N_1097);
and U2398 (N_2398,N_1663,N_1128);
and U2399 (N_2399,N_1611,N_1430);
or U2400 (N_2400,N_2141,N_2119);
nor U2401 (N_2401,N_1962,N_2376);
and U2402 (N_2402,N_2146,N_2007);
and U2403 (N_2403,N_2044,N_1954);
or U2404 (N_2404,N_1963,N_2140);
nor U2405 (N_2405,N_1897,N_1807);
nand U2406 (N_2406,N_1924,N_1970);
nand U2407 (N_2407,N_1923,N_2287);
or U2408 (N_2408,N_2344,N_1916);
or U2409 (N_2409,N_1889,N_2348);
and U2410 (N_2410,N_2265,N_2294);
or U2411 (N_2411,N_1899,N_1898);
and U2412 (N_2412,N_2027,N_2128);
and U2413 (N_2413,N_2256,N_1876);
or U2414 (N_2414,N_2058,N_2154);
or U2415 (N_2415,N_2037,N_2258);
or U2416 (N_2416,N_1888,N_2399);
nand U2417 (N_2417,N_1943,N_1951);
nand U2418 (N_2418,N_2109,N_2185);
or U2419 (N_2419,N_2130,N_2239);
and U2420 (N_2420,N_2317,N_2270);
nand U2421 (N_2421,N_1944,N_2355);
or U2422 (N_2422,N_2215,N_2072);
or U2423 (N_2423,N_2240,N_1956);
and U2424 (N_2424,N_2031,N_2024);
or U2425 (N_2425,N_1937,N_2023);
xnor U2426 (N_2426,N_1860,N_2257);
and U2427 (N_2427,N_1905,N_1826);
nand U2428 (N_2428,N_2006,N_2049);
nor U2429 (N_2429,N_2387,N_2361);
nand U2430 (N_2430,N_1988,N_1903);
nor U2431 (N_2431,N_2319,N_2112);
nand U2432 (N_2432,N_2295,N_2009);
nand U2433 (N_2433,N_2184,N_1985);
or U2434 (N_2434,N_2307,N_1852);
nand U2435 (N_2435,N_2202,N_2192);
nor U2436 (N_2436,N_1875,N_2016);
or U2437 (N_2437,N_2209,N_2190);
nor U2438 (N_2438,N_2153,N_2151);
or U2439 (N_2439,N_1839,N_2032);
nor U2440 (N_2440,N_2237,N_2325);
nand U2441 (N_2441,N_2137,N_2218);
nand U2442 (N_2442,N_2250,N_2326);
nand U2443 (N_2443,N_2067,N_2338);
nand U2444 (N_2444,N_1958,N_2288);
nand U2445 (N_2445,N_1982,N_1893);
and U2446 (N_2446,N_1906,N_2332);
nor U2447 (N_2447,N_1999,N_2122);
or U2448 (N_2448,N_2042,N_2198);
xor U2449 (N_2449,N_1877,N_1856);
and U2450 (N_2450,N_2167,N_1993);
nor U2451 (N_2451,N_2331,N_2269);
and U2452 (N_2452,N_1997,N_1827);
and U2453 (N_2453,N_2330,N_2262);
nand U2454 (N_2454,N_2203,N_1849);
or U2455 (N_2455,N_2121,N_2231);
nor U2456 (N_2456,N_2089,N_2242);
and U2457 (N_2457,N_1966,N_2139);
or U2458 (N_2458,N_2360,N_2208);
nand U2459 (N_2459,N_1821,N_1820);
or U2460 (N_2460,N_2368,N_2345);
nor U2461 (N_2461,N_2371,N_2278);
or U2462 (N_2462,N_1977,N_1878);
nand U2463 (N_2463,N_2356,N_2074);
and U2464 (N_2464,N_1834,N_2124);
or U2465 (N_2465,N_1832,N_2245);
or U2466 (N_2466,N_2100,N_1929);
nor U2467 (N_2467,N_2068,N_1902);
nand U2468 (N_2468,N_1862,N_2187);
nor U2469 (N_2469,N_2059,N_2020);
nor U2470 (N_2470,N_1994,N_1915);
and U2471 (N_2471,N_2160,N_1907);
or U2472 (N_2472,N_1829,N_2388);
nor U2473 (N_2473,N_1911,N_2143);
nand U2474 (N_2474,N_2116,N_2358);
nor U2475 (N_2475,N_2088,N_2291);
nand U2476 (N_2476,N_2354,N_2200);
or U2477 (N_2477,N_2254,N_1851);
nor U2478 (N_2478,N_1959,N_2102);
nand U2479 (N_2479,N_2373,N_2080);
or U2480 (N_2480,N_1838,N_2195);
nor U2481 (N_2481,N_1935,N_2244);
nor U2482 (N_2482,N_1955,N_2318);
and U2483 (N_2483,N_1974,N_2105);
and U2484 (N_2484,N_2223,N_2324);
nand U2485 (N_2485,N_2255,N_1855);
or U2486 (N_2486,N_2021,N_2114);
nand U2487 (N_2487,N_2306,N_2308);
and U2488 (N_2488,N_1953,N_1918);
nor U2489 (N_2489,N_1921,N_2043);
nand U2490 (N_2490,N_2147,N_2339);
or U2491 (N_2491,N_1976,N_1801);
nor U2492 (N_2492,N_2149,N_1947);
nand U2493 (N_2493,N_2086,N_1882);
nand U2494 (N_2494,N_1968,N_2191);
nor U2495 (N_2495,N_2064,N_2272);
and U2496 (N_2496,N_2186,N_2372);
or U2497 (N_2497,N_2108,N_2001);
or U2498 (N_2498,N_1967,N_1814);
nand U2499 (N_2499,N_2211,N_2230);
or U2500 (N_2500,N_1831,N_1922);
or U2501 (N_2501,N_1835,N_2129);
or U2502 (N_2502,N_1914,N_2103);
nor U2503 (N_2503,N_1981,N_2221);
or U2504 (N_2504,N_2040,N_2238);
nand U2505 (N_2505,N_2393,N_2219);
or U2506 (N_2506,N_2382,N_2075);
nand U2507 (N_2507,N_1913,N_1850);
nor U2508 (N_2508,N_2188,N_1984);
nor U2509 (N_2509,N_2333,N_2003);
nor U2510 (N_2510,N_2166,N_2159);
nand U2511 (N_2511,N_2273,N_2011);
nor U2512 (N_2512,N_2359,N_1995);
and U2513 (N_2513,N_2028,N_1992);
nor U2514 (N_2514,N_2321,N_2390);
and U2515 (N_2515,N_2304,N_2093);
and U2516 (N_2516,N_2314,N_1926);
or U2517 (N_2517,N_2030,N_2289);
or U2518 (N_2518,N_2070,N_1854);
nand U2519 (N_2519,N_2377,N_2174);
and U2520 (N_2520,N_2334,N_2161);
nor U2521 (N_2521,N_1950,N_1900);
or U2522 (N_2522,N_2320,N_1910);
or U2523 (N_2523,N_2353,N_2045);
or U2524 (N_2524,N_2090,N_1806);
and U2525 (N_2525,N_2169,N_2236);
nor U2526 (N_2526,N_2213,N_1810);
and U2527 (N_2527,N_2041,N_2181);
or U2528 (N_2528,N_2298,N_2302);
nor U2529 (N_2529,N_1932,N_1872);
or U2530 (N_2530,N_2248,N_1863);
nor U2531 (N_2531,N_2350,N_1837);
xnor U2532 (N_2532,N_2087,N_2386);
and U2533 (N_2533,N_1980,N_1987);
nand U2534 (N_2534,N_1973,N_2066);
nor U2535 (N_2535,N_2366,N_1931);
and U2536 (N_2536,N_2381,N_2183);
nand U2537 (N_2537,N_2046,N_1919);
nand U2538 (N_2538,N_2310,N_2347);
nand U2539 (N_2539,N_1983,N_1842);
nor U2540 (N_2540,N_1887,N_1942);
nor U2541 (N_2541,N_2225,N_2038);
and U2542 (N_2542,N_1928,N_2229);
nand U2543 (N_2543,N_2327,N_1841);
and U2544 (N_2544,N_2276,N_2017);
and U2545 (N_2545,N_2290,N_1930);
nand U2546 (N_2546,N_2235,N_2374);
nor U2547 (N_2547,N_1812,N_2336);
and U2548 (N_2548,N_2301,N_2152);
or U2549 (N_2549,N_1949,N_2014);
nand U2550 (N_2550,N_2123,N_2165);
nor U2551 (N_2551,N_2106,N_2252);
nor U2552 (N_2552,N_2134,N_1886);
or U2553 (N_2553,N_1848,N_1961);
nand U2554 (N_2554,N_2085,N_2227);
or U2555 (N_2555,N_2002,N_2052);
or U2556 (N_2556,N_2398,N_1901);
nor U2557 (N_2557,N_1836,N_2107);
xor U2558 (N_2558,N_2117,N_2069);
or U2559 (N_2559,N_2172,N_2267);
and U2560 (N_2560,N_1803,N_2284);
nand U2561 (N_2561,N_1991,N_2328);
and U2562 (N_2562,N_2279,N_2133);
nand U2563 (N_2563,N_2145,N_1811);
xor U2564 (N_2564,N_2010,N_1964);
nor U2565 (N_2565,N_1945,N_1904);
or U2566 (N_2566,N_2115,N_2025);
nand U2567 (N_2567,N_2363,N_2197);
nand U2568 (N_2568,N_2061,N_2005);
or U2569 (N_2569,N_1894,N_2234);
nor U2570 (N_2570,N_1873,N_2083);
or U2571 (N_2571,N_1866,N_2228);
nand U2572 (N_2572,N_1975,N_2346);
and U2573 (N_2573,N_1927,N_1885);
or U2574 (N_2574,N_2018,N_2383);
nor U2575 (N_2575,N_2311,N_2065);
or U2576 (N_2576,N_2182,N_2035);
nor U2577 (N_2577,N_1845,N_2176);
nor U2578 (N_2578,N_2341,N_1952);
nor U2579 (N_2579,N_1925,N_2034);
nand U2580 (N_2580,N_1892,N_2050);
nand U2581 (N_2581,N_2253,N_2053);
nand U2582 (N_2582,N_2029,N_2051);
nor U2583 (N_2583,N_2084,N_2394);
nor U2584 (N_2584,N_2156,N_2274);
nor U2585 (N_2585,N_2039,N_1971);
or U2586 (N_2586,N_2177,N_1909);
nand U2587 (N_2587,N_2155,N_2362);
nor U2588 (N_2588,N_2364,N_2077);
or U2589 (N_2589,N_2092,N_2391);
nor U2590 (N_2590,N_2232,N_1978);
or U2591 (N_2591,N_2392,N_2268);
and U2592 (N_2592,N_1867,N_1822);
nand U2593 (N_2593,N_1868,N_2312);
nand U2594 (N_2594,N_2125,N_2144);
nor U2595 (N_2595,N_2081,N_2063);
or U2596 (N_2596,N_1933,N_1920);
nand U2597 (N_2597,N_1881,N_2060);
and U2598 (N_2598,N_2299,N_2309);
nand U2599 (N_2599,N_1809,N_2206);
nand U2600 (N_2600,N_2286,N_2384);
nand U2601 (N_2601,N_2196,N_2012);
nand U2602 (N_2602,N_2099,N_1864);
and U2603 (N_2603,N_2389,N_2241);
or U2604 (N_2604,N_2094,N_2054);
and U2605 (N_2605,N_2170,N_1986);
nand U2606 (N_2606,N_2277,N_2095);
and U2607 (N_2607,N_2164,N_2179);
and U2608 (N_2608,N_2322,N_2135);
or U2609 (N_2609,N_1979,N_1936);
nand U2610 (N_2610,N_2297,N_2013);
nand U2611 (N_2611,N_1865,N_2217);
nand U2612 (N_2612,N_2148,N_2266);
or U2613 (N_2613,N_1883,N_2222);
nor U2614 (N_2614,N_2205,N_2096);
and U2615 (N_2615,N_2204,N_1828);
nand U2616 (N_2616,N_2048,N_2282);
nand U2617 (N_2617,N_1990,N_2104);
nor U2618 (N_2618,N_1940,N_2150);
nand U2619 (N_2619,N_1896,N_1939);
and U2620 (N_2620,N_2340,N_2079);
and U2621 (N_2621,N_2136,N_1857);
and U2622 (N_2622,N_1825,N_2375);
nor U2623 (N_2623,N_2380,N_1890);
or U2624 (N_2624,N_2026,N_1869);
and U2625 (N_2625,N_2249,N_2396);
or U2626 (N_2626,N_2178,N_2131);
nor U2627 (N_2627,N_1853,N_1846);
nor U2628 (N_2628,N_1884,N_1946);
and U2629 (N_2629,N_1805,N_2163);
and U2630 (N_2630,N_2226,N_1996);
and U2631 (N_2631,N_2263,N_2057);
and U2632 (N_2632,N_2110,N_2243);
nand U2633 (N_2633,N_2292,N_1816);
and U2634 (N_2634,N_1912,N_2303);
or U2635 (N_2635,N_1819,N_2015);
or U2636 (N_2636,N_1934,N_1972);
nand U2637 (N_2637,N_2329,N_2210);
nor U2638 (N_2638,N_1813,N_2264);
nor U2639 (N_2639,N_1823,N_1965);
or U2640 (N_2640,N_1891,N_1960);
and U2641 (N_2641,N_2033,N_2293);
nor U2642 (N_2642,N_2082,N_2158);
nor U2643 (N_2643,N_1871,N_2315);
nand U2644 (N_2644,N_1989,N_2091);
or U2645 (N_2645,N_2078,N_2138);
nand U2646 (N_2646,N_2126,N_2300);
and U2647 (N_2647,N_2370,N_2071);
or U2648 (N_2648,N_1874,N_1800);
nand U2649 (N_2649,N_2120,N_2313);
or U2650 (N_2650,N_1840,N_1861);
and U2651 (N_2651,N_2357,N_2275);
and U2652 (N_2652,N_1815,N_2212);
or U2653 (N_2653,N_2285,N_2118);
and U2654 (N_2654,N_2162,N_2207);
nand U2655 (N_2655,N_1858,N_1802);
nor U2656 (N_2656,N_1818,N_2283);
nand U2657 (N_2657,N_1847,N_2261);
nor U2658 (N_2658,N_2216,N_2220);
nand U2659 (N_2659,N_2113,N_2352);
nand U2660 (N_2660,N_2189,N_2316);
or U2661 (N_2661,N_2022,N_1843);
and U2662 (N_2662,N_2365,N_2351);
or U2663 (N_2663,N_2224,N_1817);
or U2664 (N_2664,N_2323,N_2173);
nor U2665 (N_2665,N_1917,N_2047);
or U2666 (N_2666,N_2342,N_1830);
nor U2667 (N_2667,N_1957,N_2214);
nor U2668 (N_2668,N_2175,N_2101);
nand U2669 (N_2669,N_1859,N_2142);
nor U2670 (N_2670,N_2397,N_1844);
and U2671 (N_2671,N_2251,N_2367);
nand U2672 (N_2672,N_1948,N_2296);
or U2673 (N_2673,N_2004,N_2008);
nand U2674 (N_2674,N_2271,N_1998);
or U2675 (N_2675,N_2343,N_2194);
or U2676 (N_2676,N_2260,N_2111);
nor U2677 (N_2677,N_2395,N_1880);
or U2678 (N_2678,N_2379,N_2233);
and U2679 (N_2679,N_2076,N_2201);
or U2680 (N_2680,N_1879,N_2062);
nand U2681 (N_2681,N_2168,N_2335);
or U2682 (N_2682,N_1908,N_2259);
nor U2683 (N_2683,N_2378,N_1808);
and U2684 (N_2684,N_1969,N_2349);
and U2685 (N_2685,N_2171,N_2281);
and U2686 (N_2686,N_1833,N_2193);
nor U2687 (N_2687,N_2056,N_2280);
nand U2688 (N_2688,N_1895,N_1938);
nand U2689 (N_2689,N_2036,N_2199);
or U2690 (N_2690,N_2000,N_2247);
nand U2691 (N_2691,N_2055,N_1824);
and U2692 (N_2692,N_2098,N_2385);
nand U2693 (N_2693,N_2097,N_2127);
nor U2694 (N_2694,N_1870,N_2157);
nand U2695 (N_2695,N_2369,N_1804);
and U2696 (N_2696,N_2019,N_2180);
and U2697 (N_2697,N_2246,N_2132);
nor U2698 (N_2698,N_2073,N_1941);
or U2699 (N_2699,N_2337,N_2305);
nand U2700 (N_2700,N_2192,N_2282);
nand U2701 (N_2701,N_1855,N_1896);
nand U2702 (N_2702,N_2077,N_2164);
nand U2703 (N_2703,N_2080,N_2003);
or U2704 (N_2704,N_1830,N_2367);
nor U2705 (N_2705,N_1991,N_1887);
nand U2706 (N_2706,N_2346,N_1881);
and U2707 (N_2707,N_2391,N_2339);
or U2708 (N_2708,N_2207,N_2002);
and U2709 (N_2709,N_2195,N_1929);
nand U2710 (N_2710,N_2183,N_2308);
and U2711 (N_2711,N_2096,N_2170);
nor U2712 (N_2712,N_2259,N_2029);
nand U2713 (N_2713,N_2339,N_2258);
nand U2714 (N_2714,N_2216,N_1917);
and U2715 (N_2715,N_1966,N_1919);
and U2716 (N_2716,N_1932,N_2191);
or U2717 (N_2717,N_2006,N_2034);
nor U2718 (N_2718,N_2021,N_2239);
nor U2719 (N_2719,N_2272,N_2026);
or U2720 (N_2720,N_2253,N_1954);
or U2721 (N_2721,N_1840,N_1912);
or U2722 (N_2722,N_2173,N_1884);
and U2723 (N_2723,N_1934,N_2306);
nor U2724 (N_2724,N_2189,N_1948);
or U2725 (N_2725,N_2128,N_1929);
xor U2726 (N_2726,N_2163,N_2177);
nand U2727 (N_2727,N_2133,N_2106);
nand U2728 (N_2728,N_2255,N_1882);
or U2729 (N_2729,N_1851,N_1863);
nand U2730 (N_2730,N_1917,N_2008);
nor U2731 (N_2731,N_2179,N_2138);
nand U2732 (N_2732,N_2082,N_2287);
nand U2733 (N_2733,N_2219,N_1966);
nand U2734 (N_2734,N_2246,N_2129);
nand U2735 (N_2735,N_2003,N_1852);
nor U2736 (N_2736,N_2000,N_2062);
or U2737 (N_2737,N_2045,N_2176);
and U2738 (N_2738,N_1971,N_2262);
nor U2739 (N_2739,N_2224,N_1948);
nor U2740 (N_2740,N_2328,N_2043);
or U2741 (N_2741,N_1948,N_2016);
nand U2742 (N_2742,N_2162,N_1968);
nor U2743 (N_2743,N_2377,N_1902);
nand U2744 (N_2744,N_2119,N_1885);
and U2745 (N_2745,N_2185,N_2346);
nand U2746 (N_2746,N_2033,N_2221);
nand U2747 (N_2747,N_2303,N_2214);
or U2748 (N_2748,N_2291,N_1842);
or U2749 (N_2749,N_1967,N_2389);
nor U2750 (N_2750,N_1805,N_1937);
nand U2751 (N_2751,N_2320,N_1810);
nand U2752 (N_2752,N_2207,N_1803);
nand U2753 (N_2753,N_2137,N_2192);
nor U2754 (N_2754,N_1957,N_2307);
or U2755 (N_2755,N_2235,N_2263);
or U2756 (N_2756,N_2163,N_1890);
or U2757 (N_2757,N_2128,N_2279);
or U2758 (N_2758,N_2372,N_2275);
nand U2759 (N_2759,N_1946,N_1800);
nor U2760 (N_2760,N_1866,N_2086);
nand U2761 (N_2761,N_2217,N_1975);
or U2762 (N_2762,N_1812,N_2350);
or U2763 (N_2763,N_2074,N_2312);
or U2764 (N_2764,N_2259,N_2287);
and U2765 (N_2765,N_2243,N_2233);
nand U2766 (N_2766,N_2274,N_2222);
and U2767 (N_2767,N_1926,N_2098);
or U2768 (N_2768,N_2226,N_2064);
nor U2769 (N_2769,N_2141,N_2201);
or U2770 (N_2770,N_2080,N_1823);
nor U2771 (N_2771,N_1918,N_1843);
and U2772 (N_2772,N_2110,N_2354);
and U2773 (N_2773,N_2080,N_1848);
and U2774 (N_2774,N_2138,N_1879);
nand U2775 (N_2775,N_2284,N_2361);
nand U2776 (N_2776,N_2169,N_2202);
nand U2777 (N_2777,N_2015,N_1832);
nand U2778 (N_2778,N_2184,N_2191);
or U2779 (N_2779,N_2206,N_2311);
nor U2780 (N_2780,N_2358,N_1993);
nor U2781 (N_2781,N_1943,N_1989);
nand U2782 (N_2782,N_2091,N_1946);
and U2783 (N_2783,N_2057,N_2281);
and U2784 (N_2784,N_2070,N_2035);
nand U2785 (N_2785,N_2361,N_2373);
nand U2786 (N_2786,N_2090,N_1978);
nor U2787 (N_2787,N_2322,N_2376);
or U2788 (N_2788,N_1880,N_1864);
or U2789 (N_2789,N_2084,N_2364);
and U2790 (N_2790,N_2150,N_2115);
nor U2791 (N_2791,N_1936,N_2100);
nand U2792 (N_2792,N_1919,N_1818);
or U2793 (N_2793,N_1995,N_1851);
nand U2794 (N_2794,N_2017,N_2021);
nand U2795 (N_2795,N_2373,N_2292);
or U2796 (N_2796,N_2030,N_2155);
nand U2797 (N_2797,N_2025,N_2302);
nor U2798 (N_2798,N_1950,N_2050);
or U2799 (N_2799,N_2349,N_1905);
or U2800 (N_2800,N_2382,N_1999);
and U2801 (N_2801,N_2037,N_2040);
nor U2802 (N_2802,N_2398,N_2397);
nand U2803 (N_2803,N_1897,N_2175);
nor U2804 (N_2804,N_1936,N_2178);
nand U2805 (N_2805,N_1988,N_1929);
nor U2806 (N_2806,N_2224,N_2321);
and U2807 (N_2807,N_1845,N_2271);
or U2808 (N_2808,N_1949,N_2334);
and U2809 (N_2809,N_1850,N_1968);
or U2810 (N_2810,N_2199,N_1870);
and U2811 (N_2811,N_1848,N_1985);
or U2812 (N_2812,N_2103,N_2097);
or U2813 (N_2813,N_2128,N_2377);
nor U2814 (N_2814,N_1961,N_2300);
nor U2815 (N_2815,N_2197,N_1999);
nor U2816 (N_2816,N_2081,N_1804);
or U2817 (N_2817,N_1964,N_1860);
or U2818 (N_2818,N_2234,N_2137);
and U2819 (N_2819,N_2285,N_2253);
nor U2820 (N_2820,N_1807,N_1920);
and U2821 (N_2821,N_1873,N_1915);
nor U2822 (N_2822,N_2293,N_2040);
nor U2823 (N_2823,N_1894,N_1933);
and U2824 (N_2824,N_2036,N_2145);
or U2825 (N_2825,N_1827,N_1987);
or U2826 (N_2826,N_2055,N_2177);
or U2827 (N_2827,N_1983,N_2257);
or U2828 (N_2828,N_1882,N_2075);
nor U2829 (N_2829,N_2099,N_2068);
or U2830 (N_2830,N_2192,N_1880);
nor U2831 (N_2831,N_2036,N_2224);
or U2832 (N_2832,N_2335,N_2315);
nand U2833 (N_2833,N_2162,N_2246);
nand U2834 (N_2834,N_2246,N_1909);
or U2835 (N_2835,N_2362,N_2148);
and U2836 (N_2836,N_2197,N_2099);
nor U2837 (N_2837,N_2203,N_1909);
and U2838 (N_2838,N_1995,N_1811);
or U2839 (N_2839,N_1948,N_2117);
nor U2840 (N_2840,N_2199,N_1800);
or U2841 (N_2841,N_1808,N_1965);
and U2842 (N_2842,N_2020,N_2312);
nand U2843 (N_2843,N_2355,N_1855);
and U2844 (N_2844,N_1890,N_2188);
nor U2845 (N_2845,N_2015,N_2385);
and U2846 (N_2846,N_1998,N_2127);
or U2847 (N_2847,N_2105,N_2284);
nand U2848 (N_2848,N_2305,N_2325);
or U2849 (N_2849,N_2070,N_2050);
xnor U2850 (N_2850,N_2350,N_1997);
nor U2851 (N_2851,N_2247,N_1846);
and U2852 (N_2852,N_2159,N_2394);
or U2853 (N_2853,N_2343,N_1820);
and U2854 (N_2854,N_1803,N_2164);
or U2855 (N_2855,N_2362,N_2263);
nor U2856 (N_2856,N_1988,N_2290);
or U2857 (N_2857,N_1997,N_1809);
xor U2858 (N_2858,N_2094,N_2305);
nand U2859 (N_2859,N_2221,N_2034);
or U2860 (N_2860,N_2348,N_2007);
nor U2861 (N_2861,N_1904,N_2243);
and U2862 (N_2862,N_2397,N_2311);
nor U2863 (N_2863,N_2040,N_2301);
nand U2864 (N_2864,N_2356,N_1957);
or U2865 (N_2865,N_2223,N_2285);
nor U2866 (N_2866,N_2236,N_2110);
and U2867 (N_2867,N_1864,N_1964);
and U2868 (N_2868,N_2000,N_1856);
nand U2869 (N_2869,N_1914,N_2218);
or U2870 (N_2870,N_2118,N_2085);
nor U2871 (N_2871,N_1861,N_1918);
nand U2872 (N_2872,N_2047,N_2342);
nand U2873 (N_2873,N_1969,N_2359);
or U2874 (N_2874,N_2226,N_2056);
or U2875 (N_2875,N_2365,N_2104);
nor U2876 (N_2876,N_2107,N_2370);
or U2877 (N_2877,N_2361,N_1869);
nand U2878 (N_2878,N_2202,N_1972);
nor U2879 (N_2879,N_1812,N_2150);
nor U2880 (N_2880,N_2154,N_2117);
and U2881 (N_2881,N_2329,N_1831);
nand U2882 (N_2882,N_2220,N_1800);
and U2883 (N_2883,N_2291,N_2275);
and U2884 (N_2884,N_1978,N_2218);
xor U2885 (N_2885,N_2347,N_1951);
and U2886 (N_2886,N_2221,N_2374);
nand U2887 (N_2887,N_2092,N_2019);
and U2888 (N_2888,N_1876,N_2059);
nand U2889 (N_2889,N_2187,N_2314);
nand U2890 (N_2890,N_2331,N_1964);
and U2891 (N_2891,N_2100,N_2215);
and U2892 (N_2892,N_2278,N_2359);
and U2893 (N_2893,N_2290,N_1877);
nand U2894 (N_2894,N_1898,N_1946);
or U2895 (N_2895,N_1872,N_1828);
and U2896 (N_2896,N_2384,N_1885);
nand U2897 (N_2897,N_1802,N_2228);
and U2898 (N_2898,N_2025,N_1857);
and U2899 (N_2899,N_1912,N_1998);
xnor U2900 (N_2900,N_2251,N_2074);
nand U2901 (N_2901,N_2072,N_2337);
nor U2902 (N_2902,N_2023,N_2194);
nand U2903 (N_2903,N_1861,N_2063);
nor U2904 (N_2904,N_2037,N_2296);
nand U2905 (N_2905,N_2373,N_1887);
and U2906 (N_2906,N_2030,N_2016);
and U2907 (N_2907,N_1853,N_2217);
and U2908 (N_2908,N_2349,N_1808);
nor U2909 (N_2909,N_1946,N_2223);
xnor U2910 (N_2910,N_1872,N_2352);
nor U2911 (N_2911,N_2191,N_2132);
and U2912 (N_2912,N_2249,N_2222);
and U2913 (N_2913,N_2166,N_2316);
or U2914 (N_2914,N_1873,N_2155);
or U2915 (N_2915,N_2340,N_2140);
or U2916 (N_2916,N_2175,N_1811);
nand U2917 (N_2917,N_2250,N_1844);
nand U2918 (N_2918,N_1929,N_2267);
nor U2919 (N_2919,N_1840,N_1954);
nor U2920 (N_2920,N_2258,N_2271);
nand U2921 (N_2921,N_2007,N_2190);
and U2922 (N_2922,N_1978,N_2028);
and U2923 (N_2923,N_1891,N_2372);
xnor U2924 (N_2924,N_1954,N_2351);
or U2925 (N_2925,N_2395,N_2096);
and U2926 (N_2926,N_2343,N_2144);
nand U2927 (N_2927,N_2134,N_1849);
nor U2928 (N_2928,N_1871,N_1814);
or U2929 (N_2929,N_2207,N_2046);
xnor U2930 (N_2930,N_2220,N_2057);
nand U2931 (N_2931,N_2033,N_2234);
nor U2932 (N_2932,N_2225,N_2251);
and U2933 (N_2933,N_1808,N_2179);
nor U2934 (N_2934,N_1878,N_2048);
and U2935 (N_2935,N_1851,N_2395);
and U2936 (N_2936,N_2279,N_1800);
nor U2937 (N_2937,N_1906,N_2043);
and U2938 (N_2938,N_2104,N_2199);
or U2939 (N_2939,N_2064,N_2254);
or U2940 (N_2940,N_2306,N_1986);
or U2941 (N_2941,N_1816,N_2027);
nor U2942 (N_2942,N_2101,N_1932);
nor U2943 (N_2943,N_1805,N_2129);
xnor U2944 (N_2944,N_2198,N_1969);
nand U2945 (N_2945,N_2306,N_2099);
nor U2946 (N_2946,N_2274,N_2234);
or U2947 (N_2947,N_2246,N_1911);
and U2948 (N_2948,N_1827,N_2082);
nand U2949 (N_2949,N_1868,N_2131);
nand U2950 (N_2950,N_2082,N_1956);
or U2951 (N_2951,N_1932,N_2053);
nand U2952 (N_2952,N_1957,N_2064);
or U2953 (N_2953,N_2361,N_2262);
or U2954 (N_2954,N_2287,N_2067);
or U2955 (N_2955,N_2062,N_2099);
or U2956 (N_2956,N_2027,N_2093);
or U2957 (N_2957,N_2054,N_2052);
nor U2958 (N_2958,N_1849,N_2154);
or U2959 (N_2959,N_2030,N_1845);
and U2960 (N_2960,N_1821,N_2111);
and U2961 (N_2961,N_2133,N_1912);
or U2962 (N_2962,N_1883,N_2035);
or U2963 (N_2963,N_2363,N_1910);
nand U2964 (N_2964,N_2202,N_2231);
and U2965 (N_2965,N_1931,N_1829);
nand U2966 (N_2966,N_1959,N_1831);
nor U2967 (N_2967,N_1983,N_2208);
and U2968 (N_2968,N_2023,N_1995);
or U2969 (N_2969,N_2277,N_2024);
and U2970 (N_2970,N_2107,N_2090);
or U2971 (N_2971,N_2250,N_1986);
and U2972 (N_2972,N_1963,N_2166);
nor U2973 (N_2973,N_2171,N_1888);
and U2974 (N_2974,N_2152,N_1802);
or U2975 (N_2975,N_2019,N_1831);
and U2976 (N_2976,N_2097,N_2125);
and U2977 (N_2977,N_2162,N_1947);
and U2978 (N_2978,N_2057,N_1978);
nand U2979 (N_2979,N_1817,N_2241);
or U2980 (N_2980,N_2241,N_2394);
and U2981 (N_2981,N_2056,N_2010);
or U2982 (N_2982,N_1863,N_1924);
or U2983 (N_2983,N_2288,N_2157);
and U2984 (N_2984,N_2365,N_2391);
or U2985 (N_2985,N_1920,N_1821);
and U2986 (N_2986,N_2094,N_2004);
nor U2987 (N_2987,N_2238,N_2131);
or U2988 (N_2988,N_2005,N_2172);
or U2989 (N_2989,N_2142,N_1946);
nand U2990 (N_2990,N_2175,N_2255);
nor U2991 (N_2991,N_2022,N_2161);
nor U2992 (N_2992,N_2177,N_1928);
and U2993 (N_2993,N_2350,N_2065);
nor U2994 (N_2994,N_2307,N_2074);
and U2995 (N_2995,N_2308,N_1985);
nor U2996 (N_2996,N_1933,N_2112);
nand U2997 (N_2997,N_2116,N_2396);
or U2998 (N_2998,N_2073,N_2373);
and U2999 (N_2999,N_2041,N_2173);
nor U3000 (N_3000,N_2607,N_2935);
nand U3001 (N_3001,N_2863,N_2884);
nand U3002 (N_3002,N_2593,N_2846);
nand U3003 (N_3003,N_2597,N_2862);
nand U3004 (N_3004,N_2524,N_2584);
and U3005 (N_3005,N_2818,N_2923);
nand U3006 (N_3006,N_2528,N_2518);
xor U3007 (N_3007,N_2747,N_2745);
nor U3008 (N_3008,N_2474,N_2601);
or U3009 (N_3009,N_2605,N_2835);
or U3010 (N_3010,N_2682,N_2979);
or U3011 (N_3011,N_2987,N_2968);
nand U3012 (N_3012,N_2566,N_2770);
nand U3013 (N_3013,N_2877,N_2422);
nor U3014 (N_3014,N_2702,N_2828);
or U3015 (N_3015,N_2841,N_2675);
nor U3016 (N_3016,N_2455,N_2814);
or U3017 (N_3017,N_2880,N_2727);
and U3018 (N_3018,N_2598,N_2875);
and U3019 (N_3019,N_2905,N_2509);
and U3020 (N_3020,N_2452,N_2696);
nor U3021 (N_3021,N_2471,N_2646);
nor U3022 (N_3022,N_2918,N_2517);
nor U3023 (N_3023,N_2891,N_2894);
and U3024 (N_3024,N_2466,N_2774);
nand U3025 (N_3025,N_2937,N_2401);
and U3026 (N_3026,N_2489,N_2465);
xnor U3027 (N_3027,N_2402,N_2430);
and U3028 (N_3028,N_2826,N_2640);
and U3029 (N_3029,N_2473,N_2982);
and U3030 (N_3030,N_2903,N_2544);
or U3031 (N_3031,N_2656,N_2490);
or U3032 (N_3032,N_2619,N_2676);
and U3033 (N_3033,N_2998,N_2406);
nor U3034 (N_3034,N_2678,N_2761);
and U3035 (N_3035,N_2912,N_2723);
nor U3036 (N_3036,N_2834,N_2762);
and U3037 (N_3037,N_2824,N_2683);
nand U3038 (N_3038,N_2867,N_2458);
nor U3039 (N_3039,N_2405,N_2749);
nand U3040 (N_3040,N_2815,N_2913);
or U3041 (N_3041,N_2421,N_2966);
or U3042 (N_3042,N_2861,N_2716);
nor U3043 (N_3043,N_2999,N_2725);
nor U3044 (N_3044,N_2632,N_2641);
nand U3045 (N_3045,N_2475,N_2781);
nor U3046 (N_3046,N_2708,N_2782);
nor U3047 (N_3047,N_2794,N_2462);
nor U3048 (N_3048,N_2609,N_2901);
nor U3049 (N_3049,N_2472,N_2844);
or U3050 (N_3050,N_2695,N_2576);
nand U3051 (N_3051,N_2570,N_2796);
or U3052 (N_3052,N_2984,N_2831);
or U3053 (N_3053,N_2843,N_2572);
and U3054 (N_3054,N_2647,N_2625);
nand U3055 (N_3055,N_2525,N_2574);
and U3056 (N_3056,N_2849,N_2952);
xnor U3057 (N_3057,N_2942,N_2526);
and U3058 (N_3058,N_2541,N_2537);
and U3059 (N_3059,N_2642,N_2898);
nand U3060 (N_3060,N_2718,N_2470);
nand U3061 (N_3061,N_2461,N_2701);
nand U3062 (N_3062,N_2811,N_2460);
nand U3063 (N_3063,N_2519,N_2516);
and U3064 (N_3064,N_2934,N_2773);
nor U3065 (N_3065,N_2674,N_2569);
nand U3066 (N_3066,N_2902,N_2639);
or U3067 (N_3067,N_2945,N_2542);
nor U3068 (N_3068,N_2553,N_2986);
or U3069 (N_3069,N_2667,N_2737);
nor U3070 (N_3070,N_2748,N_2783);
nor U3071 (N_3071,N_2950,N_2715);
and U3072 (N_3072,N_2755,N_2658);
nand U3073 (N_3073,N_2825,N_2514);
and U3074 (N_3074,N_2837,N_2970);
nor U3075 (N_3075,N_2494,N_2842);
and U3076 (N_3076,N_2659,N_2507);
nand U3077 (N_3077,N_2531,N_2839);
and U3078 (N_3078,N_2586,N_2550);
and U3079 (N_3079,N_2477,N_2627);
and U3080 (N_3080,N_2753,N_2580);
and U3081 (N_3081,N_2820,N_2568);
and U3082 (N_3082,N_2582,N_2792);
or U3083 (N_3083,N_2956,N_2651);
and U3084 (N_3084,N_2751,N_2413);
nand U3085 (N_3085,N_2546,N_2561);
nor U3086 (N_3086,N_2744,N_2628);
or U3087 (N_3087,N_2415,N_2963);
nand U3088 (N_3088,N_2855,N_2878);
xnor U3089 (N_3089,N_2448,N_2686);
nand U3090 (N_3090,N_2946,N_2851);
and U3091 (N_3091,N_2545,N_2453);
nand U3092 (N_3092,N_2734,N_2850);
nor U3093 (N_3093,N_2602,N_2527);
and U3094 (N_3094,N_2685,N_2692);
nand U3095 (N_3095,N_2480,N_2868);
and U3096 (N_3096,N_2975,N_2510);
and U3097 (N_3097,N_2739,N_2743);
and U3098 (N_3098,N_2864,N_2504);
nand U3099 (N_3099,N_2872,N_2596);
and U3100 (N_3100,N_2463,N_2491);
or U3101 (N_3101,N_2575,N_2439);
nand U3102 (N_3102,N_2957,N_2909);
or U3103 (N_3103,N_2555,N_2931);
nand U3104 (N_3104,N_2941,N_2819);
and U3105 (N_3105,N_2548,N_2859);
and U3106 (N_3106,N_2503,N_2662);
nand U3107 (N_3107,N_2694,N_2485);
nor U3108 (N_3108,N_2629,N_2626);
nand U3109 (N_3109,N_2446,N_2958);
nor U3110 (N_3110,N_2983,N_2562);
nand U3111 (N_3111,N_2775,N_2938);
nor U3112 (N_3112,N_2432,N_2621);
and U3113 (N_3113,N_2776,N_2496);
nor U3114 (N_3114,N_2436,N_2717);
nand U3115 (N_3115,N_2549,N_2994);
or U3116 (N_3116,N_2922,N_2429);
or U3117 (N_3117,N_2735,N_2577);
nand U3118 (N_3118,N_2634,N_2411);
and U3119 (N_3119,N_2869,N_2652);
or U3120 (N_3120,N_2672,N_2660);
or U3121 (N_3121,N_2408,N_2721);
xor U3122 (N_3122,N_2758,N_2400);
nand U3123 (N_3123,N_2728,N_2705);
nor U3124 (N_3124,N_2889,N_2693);
or U3125 (N_3125,N_2876,N_2883);
nor U3126 (N_3126,N_2492,N_2926);
nand U3127 (N_3127,N_2690,N_2417);
nand U3128 (N_3128,N_2483,N_2425);
and U3129 (N_3129,N_2707,N_2440);
xnor U3130 (N_3130,N_2713,N_2499);
and U3131 (N_3131,N_2539,N_2590);
nand U3132 (N_3132,N_2559,N_2681);
or U3133 (N_3133,N_2766,N_2495);
or U3134 (N_3134,N_2791,N_2447);
nand U3135 (N_3135,N_2523,N_2976);
and U3136 (N_3136,N_2907,N_2554);
nor U3137 (N_3137,N_2767,N_2779);
or U3138 (N_3138,N_2534,N_2680);
and U3139 (N_3139,N_2997,N_2959);
nand U3140 (N_3140,N_2925,N_2616);
nor U3141 (N_3141,N_2738,N_2585);
nor U3142 (N_3142,N_2454,N_2915);
and U3143 (N_3143,N_2412,N_2671);
nand U3144 (N_3144,N_2801,N_2600);
nor U3145 (N_3145,N_2887,N_2533);
nand U3146 (N_3146,N_2592,N_2414);
or U3147 (N_3147,N_2654,N_2615);
or U3148 (N_3148,N_2505,N_2564);
or U3149 (N_3149,N_2858,N_2557);
nor U3150 (N_3150,N_2960,N_2906);
or U3151 (N_3151,N_2468,N_2703);
nor U3152 (N_3152,N_2740,N_2896);
or U3153 (N_3153,N_2778,N_2606);
and U3154 (N_3154,N_2636,N_2729);
nor U3155 (N_3155,N_2944,N_2435);
nor U3156 (N_3156,N_2985,N_2469);
and U3157 (N_3157,N_2481,N_2764);
or U3158 (N_3158,N_2486,N_2464);
or U3159 (N_3159,N_2589,N_2637);
nand U3160 (N_3160,N_2742,N_2866);
nand U3161 (N_3161,N_2445,N_2578);
or U3162 (N_3162,N_2790,N_2431);
nor U3163 (N_3163,N_2512,N_2892);
nand U3164 (N_3164,N_2964,N_2724);
and U3165 (N_3165,N_2949,N_2746);
nor U3166 (N_3166,N_2911,N_2513);
nor U3167 (N_3167,N_2832,N_2990);
and U3168 (N_3168,N_2404,N_2547);
nand U3169 (N_3169,N_2860,N_2930);
nor U3170 (N_3170,N_2812,N_2441);
and U3171 (N_3171,N_2522,N_2433);
nor U3172 (N_3172,N_2643,N_2910);
and U3173 (N_3173,N_2684,N_2560);
or U3174 (N_3174,N_2874,N_2992);
xnor U3175 (N_3175,N_2438,N_2799);
nor U3176 (N_3176,N_2928,N_2612);
nor U3177 (N_3177,N_2501,N_2852);
nand U3178 (N_3178,N_2420,N_2802);
nor U3179 (N_3179,N_2787,N_2423);
and U3180 (N_3180,N_2810,N_2857);
nor U3181 (N_3181,N_2805,N_2977);
or U3182 (N_3182,N_2836,N_2426);
nor U3183 (N_3183,N_2854,N_2583);
nand U3184 (N_3184,N_2763,N_2511);
and U3185 (N_3185,N_2587,N_2954);
nor U3186 (N_3186,N_2476,N_2943);
nand U3187 (N_3187,N_2653,N_2649);
nor U3188 (N_3188,N_2720,N_2710);
nand U3189 (N_3189,N_2888,N_2921);
xnor U3190 (N_3190,N_2962,N_2914);
or U3191 (N_3191,N_2697,N_2899);
nand U3192 (N_3192,N_2974,N_2870);
nor U3193 (N_3193,N_2416,N_2885);
or U3194 (N_3194,N_2532,N_2881);
or U3195 (N_3195,N_2594,N_2630);
nor U3196 (N_3196,N_2515,N_2830);
or U3197 (N_3197,N_2784,N_2599);
or U3198 (N_3198,N_2845,N_2648);
nor U3199 (N_3199,N_2822,N_2916);
nand U3200 (N_3200,N_2882,N_2437);
nand U3201 (N_3201,N_2558,N_2788);
or U3202 (N_3202,N_2506,N_2904);
nor U3203 (N_3203,N_2551,N_2443);
and U3204 (N_3204,N_2969,N_2478);
and U3205 (N_3205,N_2579,N_2603);
nand U3206 (N_3206,N_2700,N_2664);
nor U3207 (N_3207,N_2563,N_2591);
nand U3208 (N_3208,N_2687,N_2719);
or U3209 (N_3209,N_2530,N_2709);
or U3210 (N_3210,N_2456,N_2493);
nand U3211 (N_3211,N_2712,N_2487);
and U3212 (N_3212,N_2879,N_2795);
or U3213 (N_3213,N_2711,N_2691);
and U3214 (N_3214,N_2847,N_2807);
and U3215 (N_3215,N_2768,N_2611);
nand U3216 (N_3216,N_2813,N_2677);
or U3217 (N_3217,N_2919,N_2565);
nor U3218 (N_3218,N_2613,N_2571);
nor U3219 (N_3219,N_2622,N_2673);
nor U3220 (N_3220,N_2924,N_2552);
or U3221 (N_3221,N_2529,N_2635);
and U3222 (N_3222,N_2936,N_2953);
nor U3223 (N_3223,N_2661,N_2848);
nor U3224 (N_3224,N_2502,N_2618);
and U3225 (N_3225,N_2679,N_2624);
nor U3226 (N_3226,N_2409,N_2610);
nand U3227 (N_3227,N_2933,N_2663);
nand U3228 (N_3228,N_2459,N_2971);
or U3229 (N_3229,N_2699,N_2484);
nand U3230 (N_3230,N_2670,N_2500);
and U3231 (N_3231,N_2722,N_2543);
and U3232 (N_3232,N_2731,N_2581);
nor U3233 (N_3233,N_2772,N_2760);
and U3234 (N_3234,N_2809,N_2967);
or U3235 (N_3235,N_2827,N_2714);
nand U3236 (N_3236,N_2821,N_2991);
nand U3237 (N_3237,N_2457,N_2488);
and U3238 (N_3238,N_2785,N_2951);
and U3239 (N_3239,N_2920,N_2939);
nand U3240 (N_3240,N_2604,N_2873);
nand U3241 (N_3241,N_2595,N_2965);
nand U3242 (N_3242,N_2427,N_2623);
or U3243 (N_3243,N_2765,N_2442);
nor U3244 (N_3244,N_2840,N_2620);
and U3245 (N_3245,N_2741,N_2978);
or U3246 (N_3246,N_2786,N_2424);
or U3247 (N_3247,N_2816,N_2482);
nand U3248 (N_3248,N_2726,N_2567);
or U3249 (N_3249,N_2932,N_2657);
and U3250 (N_3250,N_2961,N_2608);
or U3251 (N_3251,N_2665,N_2980);
or U3252 (N_3252,N_2886,N_2871);
nand U3253 (N_3253,N_2508,N_2467);
and U3254 (N_3254,N_2757,N_2434);
xnor U3255 (N_3255,N_2535,N_2451);
nor U3256 (N_3256,N_2940,N_2759);
and U3257 (N_3257,N_2736,N_2806);
and U3258 (N_3258,N_2981,N_2633);
or U3259 (N_3259,N_2897,N_2947);
or U3260 (N_3260,N_2895,N_2993);
nand U3261 (N_3261,N_2730,N_2955);
nor U3262 (N_3262,N_2520,N_2804);
nor U3263 (N_3263,N_2800,N_2780);
nor U3264 (N_3264,N_2829,N_2444);
or U3265 (N_3265,N_2777,N_2750);
or U3266 (N_3266,N_2893,N_2521);
and U3267 (N_3267,N_2972,N_2838);
and U3268 (N_3268,N_2890,N_2428);
nor U3269 (N_3269,N_2973,N_2669);
nor U3270 (N_3270,N_2650,N_2908);
nand U3271 (N_3271,N_2927,N_2449);
and U3272 (N_3272,N_2732,N_2645);
and U3273 (N_3273,N_2865,N_2948);
and U3274 (N_3274,N_2900,N_2733);
and U3275 (N_3275,N_2418,N_2498);
and U3276 (N_3276,N_2988,N_2803);
and U3277 (N_3277,N_2479,N_2419);
xor U3278 (N_3278,N_2536,N_2996);
or U3279 (N_3279,N_2644,N_2617);
nand U3280 (N_3280,N_2752,N_2823);
nor U3281 (N_3281,N_2995,N_2756);
nand U3282 (N_3282,N_2407,N_2698);
nor U3283 (N_3283,N_2817,N_2688);
nor U3284 (N_3284,N_2403,N_2573);
nand U3285 (N_3285,N_2989,N_2450);
nor U3286 (N_3286,N_2410,N_2917);
or U3287 (N_3287,N_2638,N_2704);
nor U3288 (N_3288,N_2540,N_2666);
nand U3289 (N_3289,N_2614,N_2929);
nand U3290 (N_3290,N_2769,N_2833);
xnor U3291 (N_3291,N_2538,N_2556);
or U3292 (N_3292,N_2853,N_2798);
nor U3293 (N_3293,N_2655,N_2856);
and U3294 (N_3294,N_2797,N_2631);
and U3295 (N_3295,N_2808,N_2754);
nand U3296 (N_3296,N_2689,N_2497);
and U3297 (N_3297,N_2668,N_2789);
and U3298 (N_3298,N_2706,N_2793);
nor U3299 (N_3299,N_2771,N_2588);
nand U3300 (N_3300,N_2728,N_2997);
or U3301 (N_3301,N_2572,N_2680);
nand U3302 (N_3302,N_2459,N_2847);
or U3303 (N_3303,N_2666,N_2432);
nand U3304 (N_3304,N_2917,N_2955);
nand U3305 (N_3305,N_2777,N_2789);
nand U3306 (N_3306,N_2528,N_2609);
or U3307 (N_3307,N_2810,N_2577);
or U3308 (N_3308,N_2597,N_2943);
or U3309 (N_3309,N_2587,N_2710);
or U3310 (N_3310,N_2968,N_2469);
nand U3311 (N_3311,N_2754,N_2994);
nand U3312 (N_3312,N_2460,N_2887);
and U3313 (N_3313,N_2963,N_2642);
and U3314 (N_3314,N_2550,N_2483);
and U3315 (N_3315,N_2404,N_2668);
and U3316 (N_3316,N_2754,N_2998);
or U3317 (N_3317,N_2628,N_2833);
nor U3318 (N_3318,N_2534,N_2513);
or U3319 (N_3319,N_2864,N_2578);
or U3320 (N_3320,N_2773,N_2784);
or U3321 (N_3321,N_2620,N_2802);
nor U3322 (N_3322,N_2484,N_2846);
and U3323 (N_3323,N_2834,N_2510);
and U3324 (N_3324,N_2885,N_2553);
or U3325 (N_3325,N_2596,N_2939);
nand U3326 (N_3326,N_2851,N_2546);
nand U3327 (N_3327,N_2974,N_2574);
nand U3328 (N_3328,N_2674,N_2408);
nand U3329 (N_3329,N_2901,N_2795);
nand U3330 (N_3330,N_2434,N_2807);
nand U3331 (N_3331,N_2816,N_2422);
and U3332 (N_3332,N_2569,N_2632);
nor U3333 (N_3333,N_2610,N_2542);
nor U3334 (N_3334,N_2922,N_2509);
and U3335 (N_3335,N_2868,N_2714);
or U3336 (N_3336,N_2981,N_2778);
or U3337 (N_3337,N_2821,N_2495);
nor U3338 (N_3338,N_2747,N_2740);
or U3339 (N_3339,N_2893,N_2920);
nor U3340 (N_3340,N_2770,N_2835);
or U3341 (N_3341,N_2947,N_2619);
nand U3342 (N_3342,N_2595,N_2436);
and U3343 (N_3343,N_2962,N_2975);
nor U3344 (N_3344,N_2598,N_2740);
nand U3345 (N_3345,N_2493,N_2742);
and U3346 (N_3346,N_2556,N_2692);
nand U3347 (N_3347,N_2519,N_2417);
nor U3348 (N_3348,N_2749,N_2875);
nand U3349 (N_3349,N_2527,N_2756);
or U3350 (N_3350,N_2815,N_2628);
and U3351 (N_3351,N_2403,N_2802);
nand U3352 (N_3352,N_2454,N_2711);
nand U3353 (N_3353,N_2779,N_2439);
nor U3354 (N_3354,N_2776,N_2685);
nand U3355 (N_3355,N_2829,N_2643);
nand U3356 (N_3356,N_2723,N_2459);
nand U3357 (N_3357,N_2687,N_2879);
and U3358 (N_3358,N_2849,N_2696);
nand U3359 (N_3359,N_2934,N_2677);
nor U3360 (N_3360,N_2872,N_2787);
nand U3361 (N_3361,N_2482,N_2694);
xnor U3362 (N_3362,N_2893,N_2740);
or U3363 (N_3363,N_2596,N_2611);
and U3364 (N_3364,N_2623,N_2478);
nand U3365 (N_3365,N_2524,N_2768);
or U3366 (N_3366,N_2473,N_2948);
nand U3367 (N_3367,N_2498,N_2435);
and U3368 (N_3368,N_2742,N_2774);
and U3369 (N_3369,N_2915,N_2993);
or U3370 (N_3370,N_2750,N_2441);
nor U3371 (N_3371,N_2528,N_2612);
nand U3372 (N_3372,N_2905,N_2750);
and U3373 (N_3373,N_2795,N_2485);
or U3374 (N_3374,N_2972,N_2520);
nand U3375 (N_3375,N_2717,N_2875);
nor U3376 (N_3376,N_2842,N_2667);
or U3377 (N_3377,N_2867,N_2980);
nor U3378 (N_3378,N_2528,N_2895);
and U3379 (N_3379,N_2465,N_2454);
nand U3380 (N_3380,N_2953,N_2425);
nor U3381 (N_3381,N_2687,N_2421);
and U3382 (N_3382,N_2721,N_2971);
or U3383 (N_3383,N_2491,N_2934);
nor U3384 (N_3384,N_2663,N_2443);
nor U3385 (N_3385,N_2753,N_2449);
nand U3386 (N_3386,N_2671,N_2893);
or U3387 (N_3387,N_2921,N_2754);
nand U3388 (N_3388,N_2978,N_2502);
nand U3389 (N_3389,N_2405,N_2940);
and U3390 (N_3390,N_2587,N_2815);
or U3391 (N_3391,N_2770,N_2500);
nand U3392 (N_3392,N_2892,N_2525);
nand U3393 (N_3393,N_2925,N_2820);
and U3394 (N_3394,N_2595,N_2582);
nand U3395 (N_3395,N_2590,N_2781);
nand U3396 (N_3396,N_2491,N_2751);
and U3397 (N_3397,N_2942,N_2973);
nor U3398 (N_3398,N_2529,N_2535);
nand U3399 (N_3399,N_2952,N_2848);
or U3400 (N_3400,N_2841,N_2941);
nor U3401 (N_3401,N_2707,N_2844);
and U3402 (N_3402,N_2837,N_2999);
nand U3403 (N_3403,N_2845,N_2472);
or U3404 (N_3404,N_2922,N_2952);
nand U3405 (N_3405,N_2706,N_2658);
nand U3406 (N_3406,N_2462,N_2700);
nor U3407 (N_3407,N_2997,N_2720);
or U3408 (N_3408,N_2726,N_2624);
or U3409 (N_3409,N_2904,N_2995);
and U3410 (N_3410,N_2524,N_2599);
nor U3411 (N_3411,N_2664,N_2710);
nor U3412 (N_3412,N_2496,N_2464);
nor U3413 (N_3413,N_2436,N_2424);
and U3414 (N_3414,N_2961,N_2643);
nand U3415 (N_3415,N_2915,N_2797);
nor U3416 (N_3416,N_2805,N_2953);
or U3417 (N_3417,N_2983,N_2814);
and U3418 (N_3418,N_2836,N_2601);
and U3419 (N_3419,N_2911,N_2866);
and U3420 (N_3420,N_2671,N_2746);
and U3421 (N_3421,N_2411,N_2682);
or U3422 (N_3422,N_2755,N_2429);
or U3423 (N_3423,N_2730,N_2783);
xnor U3424 (N_3424,N_2495,N_2739);
xnor U3425 (N_3425,N_2833,N_2559);
or U3426 (N_3426,N_2642,N_2888);
nand U3427 (N_3427,N_2986,N_2976);
nand U3428 (N_3428,N_2491,N_2839);
or U3429 (N_3429,N_2529,N_2814);
or U3430 (N_3430,N_2712,N_2517);
nor U3431 (N_3431,N_2622,N_2615);
nand U3432 (N_3432,N_2436,N_2764);
nand U3433 (N_3433,N_2998,N_2450);
and U3434 (N_3434,N_2888,N_2609);
and U3435 (N_3435,N_2414,N_2621);
nor U3436 (N_3436,N_2848,N_2476);
nand U3437 (N_3437,N_2578,N_2941);
and U3438 (N_3438,N_2913,N_2616);
or U3439 (N_3439,N_2677,N_2970);
xnor U3440 (N_3440,N_2882,N_2516);
nand U3441 (N_3441,N_2605,N_2547);
nor U3442 (N_3442,N_2644,N_2862);
and U3443 (N_3443,N_2471,N_2742);
or U3444 (N_3444,N_2672,N_2531);
and U3445 (N_3445,N_2914,N_2609);
or U3446 (N_3446,N_2686,N_2944);
nor U3447 (N_3447,N_2725,N_2800);
and U3448 (N_3448,N_2475,N_2498);
and U3449 (N_3449,N_2776,N_2756);
or U3450 (N_3450,N_2938,N_2694);
nand U3451 (N_3451,N_2638,N_2505);
nor U3452 (N_3452,N_2747,N_2754);
nor U3453 (N_3453,N_2413,N_2492);
or U3454 (N_3454,N_2497,N_2787);
and U3455 (N_3455,N_2959,N_2530);
nor U3456 (N_3456,N_2649,N_2463);
xnor U3457 (N_3457,N_2755,N_2502);
or U3458 (N_3458,N_2682,N_2787);
and U3459 (N_3459,N_2456,N_2905);
or U3460 (N_3460,N_2825,N_2900);
and U3461 (N_3461,N_2412,N_2804);
nand U3462 (N_3462,N_2852,N_2553);
nor U3463 (N_3463,N_2740,N_2675);
nor U3464 (N_3464,N_2654,N_2922);
nand U3465 (N_3465,N_2570,N_2988);
or U3466 (N_3466,N_2931,N_2653);
nor U3467 (N_3467,N_2473,N_2813);
nand U3468 (N_3468,N_2534,N_2896);
or U3469 (N_3469,N_2961,N_2585);
nand U3470 (N_3470,N_2617,N_2700);
and U3471 (N_3471,N_2990,N_2807);
and U3472 (N_3472,N_2476,N_2593);
nor U3473 (N_3473,N_2647,N_2437);
and U3474 (N_3474,N_2519,N_2764);
and U3475 (N_3475,N_2816,N_2873);
or U3476 (N_3476,N_2544,N_2838);
or U3477 (N_3477,N_2726,N_2463);
nor U3478 (N_3478,N_2877,N_2887);
nor U3479 (N_3479,N_2941,N_2874);
and U3480 (N_3480,N_2916,N_2809);
nor U3481 (N_3481,N_2822,N_2509);
nor U3482 (N_3482,N_2449,N_2774);
nand U3483 (N_3483,N_2501,N_2889);
nor U3484 (N_3484,N_2614,N_2810);
and U3485 (N_3485,N_2556,N_2625);
nor U3486 (N_3486,N_2757,N_2740);
nor U3487 (N_3487,N_2843,N_2969);
or U3488 (N_3488,N_2861,N_2687);
nor U3489 (N_3489,N_2697,N_2781);
or U3490 (N_3490,N_2402,N_2882);
and U3491 (N_3491,N_2928,N_2849);
and U3492 (N_3492,N_2939,N_2494);
and U3493 (N_3493,N_2799,N_2560);
nand U3494 (N_3494,N_2952,N_2472);
and U3495 (N_3495,N_2776,N_2701);
and U3496 (N_3496,N_2821,N_2579);
nand U3497 (N_3497,N_2512,N_2779);
and U3498 (N_3498,N_2402,N_2486);
xnor U3499 (N_3499,N_2405,N_2928);
nand U3500 (N_3500,N_2744,N_2492);
and U3501 (N_3501,N_2592,N_2511);
xor U3502 (N_3502,N_2454,N_2881);
and U3503 (N_3503,N_2719,N_2577);
nand U3504 (N_3504,N_2640,N_2889);
nor U3505 (N_3505,N_2664,N_2472);
nand U3506 (N_3506,N_2531,N_2720);
nand U3507 (N_3507,N_2796,N_2728);
nor U3508 (N_3508,N_2742,N_2482);
or U3509 (N_3509,N_2500,N_2466);
or U3510 (N_3510,N_2790,N_2641);
or U3511 (N_3511,N_2575,N_2642);
and U3512 (N_3512,N_2557,N_2524);
or U3513 (N_3513,N_2988,N_2535);
and U3514 (N_3514,N_2547,N_2857);
and U3515 (N_3515,N_2922,N_2939);
nor U3516 (N_3516,N_2712,N_2496);
nor U3517 (N_3517,N_2580,N_2897);
and U3518 (N_3518,N_2737,N_2695);
and U3519 (N_3519,N_2668,N_2956);
or U3520 (N_3520,N_2824,N_2761);
or U3521 (N_3521,N_2694,N_2780);
or U3522 (N_3522,N_2692,N_2803);
or U3523 (N_3523,N_2800,N_2824);
or U3524 (N_3524,N_2600,N_2953);
or U3525 (N_3525,N_2527,N_2833);
or U3526 (N_3526,N_2555,N_2467);
and U3527 (N_3527,N_2764,N_2752);
or U3528 (N_3528,N_2438,N_2595);
nand U3529 (N_3529,N_2654,N_2624);
and U3530 (N_3530,N_2652,N_2613);
nand U3531 (N_3531,N_2579,N_2783);
and U3532 (N_3532,N_2444,N_2660);
and U3533 (N_3533,N_2783,N_2506);
and U3534 (N_3534,N_2471,N_2562);
and U3535 (N_3535,N_2867,N_2756);
nor U3536 (N_3536,N_2902,N_2913);
nor U3537 (N_3537,N_2448,N_2944);
and U3538 (N_3538,N_2563,N_2731);
nand U3539 (N_3539,N_2872,N_2439);
and U3540 (N_3540,N_2922,N_2431);
or U3541 (N_3541,N_2805,N_2421);
nand U3542 (N_3542,N_2439,N_2527);
nor U3543 (N_3543,N_2794,N_2967);
and U3544 (N_3544,N_2895,N_2986);
and U3545 (N_3545,N_2912,N_2883);
or U3546 (N_3546,N_2516,N_2465);
nor U3547 (N_3547,N_2843,N_2977);
or U3548 (N_3548,N_2775,N_2594);
and U3549 (N_3549,N_2589,N_2535);
or U3550 (N_3550,N_2909,N_2585);
and U3551 (N_3551,N_2786,N_2961);
and U3552 (N_3552,N_2855,N_2765);
and U3553 (N_3553,N_2620,N_2413);
nand U3554 (N_3554,N_2518,N_2805);
nand U3555 (N_3555,N_2786,N_2466);
or U3556 (N_3556,N_2482,N_2673);
and U3557 (N_3557,N_2657,N_2970);
and U3558 (N_3558,N_2646,N_2526);
nand U3559 (N_3559,N_2729,N_2649);
nor U3560 (N_3560,N_2642,N_2700);
nand U3561 (N_3561,N_2619,N_2406);
or U3562 (N_3562,N_2763,N_2530);
and U3563 (N_3563,N_2969,N_2949);
nor U3564 (N_3564,N_2920,N_2475);
and U3565 (N_3565,N_2565,N_2724);
and U3566 (N_3566,N_2530,N_2404);
nand U3567 (N_3567,N_2990,N_2796);
or U3568 (N_3568,N_2569,N_2654);
nor U3569 (N_3569,N_2652,N_2914);
nand U3570 (N_3570,N_2569,N_2635);
nor U3571 (N_3571,N_2747,N_2630);
and U3572 (N_3572,N_2939,N_2858);
and U3573 (N_3573,N_2479,N_2676);
and U3574 (N_3574,N_2716,N_2805);
nand U3575 (N_3575,N_2793,N_2758);
nor U3576 (N_3576,N_2525,N_2672);
nor U3577 (N_3577,N_2930,N_2418);
nor U3578 (N_3578,N_2756,N_2412);
or U3579 (N_3579,N_2899,N_2813);
nor U3580 (N_3580,N_2559,N_2721);
nand U3581 (N_3581,N_2857,N_2470);
and U3582 (N_3582,N_2715,N_2461);
or U3583 (N_3583,N_2596,N_2512);
nor U3584 (N_3584,N_2811,N_2714);
or U3585 (N_3585,N_2537,N_2415);
nor U3586 (N_3586,N_2552,N_2699);
and U3587 (N_3587,N_2989,N_2433);
or U3588 (N_3588,N_2755,N_2438);
nor U3589 (N_3589,N_2638,N_2675);
and U3590 (N_3590,N_2505,N_2409);
and U3591 (N_3591,N_2476,N_2531);
or U3592 (N_3592,N_2900,N_2449);
and U3593 (N_3593,N_2912,N_2611);
or U3594 (N_3594,N_2556,N_2797);
and U3595 (N_3595,N_2928,N_2743);
or U3596 (N_3596,N_2464,N_2998);
and U3597 (N_3597,N_2636,N_2755);
and U3598 (N_3598,N_2673,N_2587);
nand U3599 (N_3599,N_2870,N_2761);
nor U3600 (N_3600,N_3120,N_3525);
and U3601 (N_3601,N_3534,N_3175);
and U3602 (N_3602,N_3055,N_3369);
nor U3603 (N_3603,N_3455,N_3370);
or U3604 (N_3604,N_3279,N_3003);
nor U3605 (N_3605,N_3000,N_3133);
or U3606 (N_3606,N_3156,N_3523);
nand U3607 (N_3607,N_3463,N_3173);
or U3608 (N_3608,N_3046,N_3255);
nand U3609 (N_3609,N_3430,N_3547);
and U3610 (N_3610,N_3365,N_3020);
nor U3611 (N_3611,N_3163,N_3065);
or U3612 (N_3612,N_3006,N_3162);
xnor U3613 (N_3613,N_3249,N_3294);
and U3614 (N_3614,N_3037,N_3233);
or U3615 (N_3615,N_3590,N_3242);
or U3616 (N_3616,N_3122,N_3366);
and U3617 (N_3617,N_3351,N_3337);
or U3618 (N_3618,N_3565,N_3446);
and U3619 (N_3619,N_3361,N_3059);
xnor U3620 (N_3620,N_3155,N_3514);
or U3621 (N_3621,N_3416,N_3537);
nand U3622 (N_3622,N_3021,N_3033);
nand U3623 (N_3623,N_3450,N_3253);
nor U3624 (N_3624,N_3114,N_3013);
or U3625 (N_3625,N_3218,N_3034);
nand U3626 (N_3626,N_3464,N_3154);
or U3627 (N_3627,N_3007,N_3573);
or U3628 (N_3628,N_3354,N_3581);
and U3629 (N_3629,N_3499,N_3344);
xnor U3630 (N_3630,N_3519,N_3123);
nand U3631 (N_3631,N_3228,N_3124);
nand U3632 (N_3632,N_3554,N_3305);
nand U3633 (N_3633,N_3584,N_3313);
and U3634 (N_3634,N_3527,N_3580);
xor U3635 (N_3635,N_3243,N_3176);
and U3636 (N_3636,N_3392,N_3489);
nor U3637 (N_3637,N_3004,N_3202);
or U3638 (N_3638,N_3387,N_3212);
nand U3639 (N_3639,N_3404,N_3393);
and U3640 (N_3640,N_3290,N_3141);
and U3641 (N_3641,N_3467,N_3030);
and U3642 (N_3642,N_3582,N_3032);
nor U3643 (N_3643,N_3300,N_3427);
nand U3644 (N_3644,N_3472,N_3011);
xnor U3645 (N_3645,N_3078,N_3074);
or U3646 (N_3646,N_3509,N_3390);
or U3647 (N_3647,N_3139,N_3147);
nor U3648 (N_3648,N_3482,N_3397);
and U3649 (N_3649,N_3056,N_3268);
or U3650 (N_3650,N_3599,N_3116);
nand U3651 (N_3651,N_3301,N_3371);
and U3652 (N_3652,N_3342,N_3411);
or U3653 (N_3653,N_3359,N_3597);
or U3654 (N_3654,N_3496,N_3015);
nand U3655 (N_3655,N_3367,N_3112);
or U3656 (N_3656,N_3262,N_3346);
nor U3657 (N_3657,N_3225,N_3358);
or U3658 (N_3658,N_3500,N_3447);
nand U3659 (N_3659,N_3186,N_3398);
nand U3660 (N_3660,N_3049,N_3246);
or U3661 (N_3661,N_3363,N_3552);
nor U3662 (N_3662,N_3240,N_3276);
nor U3663 (N_3663,N_3014,N_3296);
and U3664 (N_3664,N_3043,N_3483);
and U3665 (N_3665,N_3183,N_3364);
nor U3666 (N_3666,N_3044,N_3019);
nor U3667 (N_3667,N_3577,N_3488);
xnor U3668 (N_3668,N_3150,N_3579);
nand U3669 (N_3669,N_3136,N_3281);
and U3670 (N_3670,N_3199,N_3062);
nand U3671 (N_3671,N_3017,N_3381);
or U3672 (N_3672,N_3435,N_3185);
or U3673 (N_3673,N_3480,N_3553);
nand U3674 (N_3674,N_3475,N_3031);
or U3675 (N_3675,N_3576,N_3314);
nand U3676 (N_3676,N_3545,N_3506);
nand U3677 (N_3677,N_3385,N_3018);
nor U3678 (N_3678,N_3336,N_3091);
and U3679 (N_3679,N_3302,N_3257);
nor U3680 (N_3680,N_3293,N_3317);
nand U3681 (N_3681,N_3087,N_3140);
and U3682 (N_3682,N_3515,N_3022);
or U3683 (N_3683,N_3159,N_3110);
nand U3684 (N_3684,N_3066,N_3591);
nand U3685 (N_3685,N_3415,N_3278);
or U3686 (N_3686,N_3226,N_3431);
or U3687 (N_3687,N_3588,N_3170);
nand U3688 (N_3688,N_3035,N_3318);
nor U3689 (N_3689,N_3291,N_3439);
or U3690 (N_3690,N_3008,N_3556);
and U3691 (N_3691,N_3395,N_3571);
nand U3692 (N_3692,N_3187,N_3511);
or U3693 (N_3693,N_3047,N_3461);
or U3694 (N_3694,N_3520,N_3075);
nand U3695 (N_3695,N_3459,N_3321);
nand U3696 (N_3696,N_3048,N_3205);
nand U3697 (N_3697,N_3535,N_3105);
nor U3698 (N_3698,N_3221,N_3169);
nand U3699 (N_3699,N_3138,N_3109);
nor U3700 (N_3700,N_3260,N_3077);
and U3701 (N_3701,N_3039,N_3328);
nor U3702 (N_3702,N_3270,N_3117);
or U3703 (N_3703,N_3272,N_3266);
nor U3704 (N_3704,N_3587,N_3191);
or U3705 (N_3705,N_3287,N_3490);
and U3706 (N_3706,N_3115,N_3143);
nand U3707 (N_3707,N_3353,N_3448);
or U3708 (N_3708,N_3211,N_3379);
nand U3709 (N_3709,N_3219,N_3437);
and U3710 (N_3710,N_3569,N_3438);
or U3711 (N_3711,N_3544,N_3360);
nor U3712 (N_3712,N_3441,N_3100);
nor U3713 (N_3713,N_3132,N_3513);
nor U3714 (N_3714,N_3247,N_3286);
nand U3715 (N_3715,N_3418,N_3241);
nor U3716 (N_3716,N_3434,N_3009);
or U3717 (N_3717,N_3086,N_3469);
nand U3718 (N_3718,N_3494,N_3103);
nand U3719 (N_3719,N_3274,N_3531);
nand U3720 (N_3720,N_3174,N_3196);
and U3721 (N_3721,N_3200,N_3144);
nand U3722 (N_3722,N_3195,N_3157);
nand U3723 (N_3723,N_3094,N_3258);
nand U3724 (N_3724,N_3306,N_3473);
or U3725 (N_3725,N_3181,N_3401);
and U3726 (N_3726,N_3516,N_3252);
nand U3727 (N_3727,N_3512,N_3182);
nor U3728 (N_3728,N_3320,N_3327);
nand U3729 (N_3729,N_3478,N_3023);
nor U3730 (N_3730,N_3410,N_3555);
nor U3731 (N_3731,N_3568,N_3010);
or U3732 (N_3732,N_3244,N_3166);
or U3733 (N_3733,N_3384,N_3421);
or U3734 (N_3734,N_3507,N_3025);
nor U3735 (N_3735,N_3217,N_3304);
and U3736 (N_3736,N_3308,N_3505);
or U3737 (N_3737,N_3498,N_3206);
and U3738 (N_3738,N_3510,N_3468);
and U3739 (N_3739,N_3179,N_3562);
nand U3740 (N_3740,N_3493,N_3106);
nor U3741 (N_3741,N_3350,N_3101);
nand U3742 (N_3742,N_3551,N_3029);
nor U3743 (N_3743,N_3129,N_3058);
and U3744 (N_3744,N_3542,N_3085);
or U3745 (N_3745,N_3236,N_3130);
and U3746 (N_3746,N_3315,N_3566);
nor U3747 (N_3747,N_3097,N_3288);
and U3748 (N_3748,N_3343,N_3053);
nor U3749 (N_3749,N_3425,N_3319);
or U3750 (N_3750,N_3082,N_3456);
nand U3751 (N_3751,N_3177,N_3477);
nor U3752 (N_3752,N_3457,N_3083);
or U3753 (N_3753,N_3026,N_3099);
or U3754 (N_3754,N_3214,N_3382);
or U3755 (N_3755,N_3423,N_3341);
nand U3756 (N_3756,N_3502,N_3549);
and U3757 (N_3757,N_3378,N_3491);
or U3758 (N_3758,N_3238,N_3424);
nor U3759 (N_3759,N_3526,N_3178);
or U3760 (N_3760,N_3089,N_3108);
and U3761 (N_3761,N_3299,N_3376);
nand U3762 (N_3762,N_3528,N_3307);
nand U3763 (N_3763,N_3297,N_3107);
xnor U3764 (N_3764,N_3192,N_3152);
and U3765 (N_3765,N_3201,N_3068);
and U3766 (N_3766,N_3119,N_3149);
or U3767 (N_3767,N_3040,N_3209);
or U3768 (N_3768,N_3076,N_3203);
nor U3769 (N_3769,N_3422,N_3072);
xnor U3770 (N_3770,N_3060,N_3374);
nor U3771 (N_3771,N_3237,N_3208);
or U3772 (N_3772,N_3198,N_3057);
and U3773 (N_3773,N_3067,N_3230);
or U3774 (N_3774,N_3229,N_3349);
nor U3775 (N_3775,N_3578,N_3271);
nor U3776 (N_3776,N_3593,N_3567);
or U3777 (N_3777,N_3102,N_3180);
nand U3778 (N_3778,N_3284,N_3050);
and U3779 (N_3779,N_3380,N_3460);
or U3780 (N_3780,N_3090,N_3184);
and U3781 (N_3781,N_3570,N_3292);
nor U3782 (N_3782,N_3557,N_3042);
and U3783 (N_3783,N_3322,N_3227);
or U3784 (N_3784,N_3399,N_3412);
or U3785 (N_3785,N_3064,N_3171);
nand U3786 (N_3786,N_3540,N_3484);
nor U3787 (N_3787,N_3440,N_3476);
nor U3788 (N_3788,N_3407,N_3355);
nor U3789 (N_3789,N_3234,N_3080);
nor U3790 (N_3790,N_3362,N_3536);
and U3791 (N_3791,N_3197,N_3093);
and U3792 (N_3792,N_3054,N_3027);
nand U3793 (N_3793,N_3128,N_3148);
nor U3794 (N_3794,N_3347,N_3561);
or U3795 (N_3795,N_3081,N_3405);
nor U3796 (N_3796,N_3492,N_3215);
or U3797 (N_3797,N_3316,N_3312);
nand U3798 (N_3798,N_3550,N_3095);
and U3799 (N_3799,N_3503,N_3583);
nand U3800 (N_3800,N_3388,N_3486);
and U3801 (N_3801,N_3168,N_3465);
or U3802 (N_3802,N_3332,N_3310);
nand U3803 (N_3803,N_3220,N_3045);
or U3804 (N_3804,N_3331,N_3239);
nand U3805 (N_3805,N_3016,N_3267);
and U3806 (N_3806,N_3433,N_3134);
or U3807 (N_3807,N_3071,N_3028);
nor U3808 (N_3808,N_3487,N_3224);
nor U3809 (N_3809,N_3232,N_3245);
nand U3810 (N_3810,N_3559,N_3326);
nand U3811 (N_3811,N_3289,N_3449);
and U3812 (N_3812,N_3403,N_3298);
or U3813 (N_3813,N_3036,N_3546);
nand U3814 (N_3814,N_3495,N_3146);
and U3815 (N_3815,N_3428,N_3231);
and U3816 (N_3816,N_3400,N_3548);
or U3817 (N_3817,N_3466,N_3564);
or U3818 (N_3818,N_3479,N_3521);
nand U3819 (N_3819,N_3596,N_3160);
nand U3820 (N_3820,N_3452,N_3436);
or U3821 (N_3821,N_3222,N_3558);
and U3822 (N_3822,N_3137,N_3283);
or U3823 (N_3823,N_3470,N_3394);
and U3824 (N_3824,N_3204,N_3586);
nand U3825 (N_3825,N_3073,N_3210);
nor U3826 (N_3826,N_3481,N_3126);
nor U3827 (N_3827,N_3575,N_3330);
nand U3828 (N_3828,N_3420,N_3442);
or U3829 (N_3829,N_3275,N_3061);
nand U3830 (N_3830,N_3453,N_3541);
nor U3831 (N_3831,N_3263,N_3508);
nor U3832 (N_3832,N_3118,N_3190);
and U3833 (N_3833,N_3277,N_3193);
nand U3834 (N_3834,N_3522,N_3098);
nand U3835 (N_3835,N_3264,N_3529);
or U3836 (N_3836,N_3352,N_3069);
and U3837 (N_3837,N_3084,N_3386);
nand U3838 (N_3838,N_3265,N_3532);
nand U3839 (N_3839,N_3572,N_3063);
or U3840 (N_3840,N_3145,N_3164);
nand U3841 (N_3841,N_3356,N_3339);
nor U3842 (N_3842,N_3323,N_3485);
or U3843 (N_3843,N_3530,N_3251);
or U3844 (N_3844,N_3375,N_3213);
nand U3845 (N_3845,N_3443,N_3135);
nor U3846 (N_3846,N_3092,N_3161);
nand U3847 (N_3847,N_3172,N_3396);
nor U3848 (N_3848,N_3088,N_3372);
nand U3849 (N_3849,N_3165,N_3402);
and U3850 (N_3850,N_3451,N_3269);
or U3851 (N_3851,N_3104,N_3595);
or U3852 (N_3852,N_3216,N_3038);
nor U3853 (N_3853,N_3261,N_3345);
and U3854 (N_3854,N_3563,N_3311);
and U3855 (N_3855,N_3167,N_3254);
and U3856 (N_3856,N_3194,N_3121);
or U3857 (N_3857,N_3189,N_3002);
or U3858 (N_3858,N_3429,N_3524);
nand U3859 (N_3859,N_3052,N_3417);
nand U3860 (N_3860,N_3406,N_3585);
nor U3861 (N_3861,N_3334,N_3444);
nand U3862 (N_3862,N_3079,N_3333);
nor U3863 (N_3863,N_3113,N_3153);
nand U3864 (N_3864,N_3426,N_3504);
nand U3865 (N_3865,N_3329,N_3325);
nand U3866 (N_3866,N_3096,N_3501);
nand U3867 (N_3867,N_3051,N_3391);
nand U3868 (N_3868,N_3273,N_3598);
and U3869 (N_3869,N_3001,N_3419);
or U3870 (N_3870,N_3259,N_3533);
nor U3871 (N_3871,N_3131,N_3070);
nor U3872 (N_3872,N_3235,N_3539);
nor U3873 (N_3873,N_3207,N_3471);
and U3874 (N_3874,N_3041,N_3151);
nor U3875 (N_3875,N_3324,N_3368);
nor U3876 (N_3876,N_3432,N_3295);
nand U3877 (N_3877,N_3285,N_3589);
nand U3878 (N_3878,N_3282,N_3409);
or U3879 (N_3879,N_3024,N_3223);
or U3880 (N_3880,N_3335,N_3250);
nor U3881 (N_3881,N_3338,N_3309);
nand U3882 (N_3882,N_3594,N_3408);
nor U3883 (N_3883,N_3454,N_3256);
nand U3884 (N_3884,N_3538,N_3560);
or U3885 (N_3885,N_3413,N_3142);
or U3886 (N_3886,N_3383,N_3373);
or U3887 (N_3887,N_3497,N_3389);
or U3888 (N_3888,N_3303,N_3592);
nor U3889 (N_3889,N_3518,N_3517);
and U3890 (N_3890,N_3357,N_3012);
nand U3891 (N_3891,N_3474,N_3280);
nor U3892 (N_3892,N_3127,N_3158);
nor U3893 (N_3893,N_3462,N_3340);
nand U3894 (N_3894,N_3574,N_3111);
or U3895 (N_3895,N_3348,N_3248);
or U3896 (N_3896,N_3445,N_3125);
nand U3897 (N_3897,N_3414,N_3005);
or U3898 (N_3898,N_3543,N_3188);
or U3899 (N_3899,N_3458,N_3377);
nand U3900 (N_3900,N_3218,N_3372);
nand U3901 (N_3901,N_3497,N_3582);
and U3902 (N_3902,N_3493,N_3581);
and U3903 (N_3903,N_3072,N_3091);
nand U3904 (N_3904,N_3059,N_3589);
nand U3905 (N_3905,N_3147,N_3234);
xnor U3906 (N_3906,N_3550,N_3112);
and U3907 (N_3907,N_3562,N_3503);
nand U3908 (N_3908,N_3018,N_3548);
nand U3909 (N_3909,N_3040,N_3151);
or U3910 (N_3910,N_3577,N_3403);
or U3911 (N_3911,N_3199,N_3578);
nor U3912 (N_3912,N_3077,N_3039);
nor U3913 (N_3913,N_3032,N_3187);
xnor U3914 (N_3914,N_3096,N_3468);
or U3915 (N_3915,N_3121,N_3136);
nor U3916 (N_3916,N_3089,N_3514);
or U3917 (N_3917,N_3136,N_3233);
and U3918 (N_3918,N_3476,N_3083);
or U3919 (N_3919,N_3365,N_3423);
xnor U3920 (N_3920,N_3053,N_3107);
and U3921 (N_3921,N_3228,N_3549);
and U3922 (N_3922,N_3509,N_3458);
nand U3923 (N_3923,N_3182,N_3378);
nor U3924 (N_3924,N_3191,N_3419);
nor U3925 (N_3925,N_3083,N_3568);
or U3926 (N_3926,N_3099,N_3083);
nand U3927 (N_3927,N_3043,N_3585);
or U3928 (N_3928,N_3213,N_3285);
or U3929 (N_3929,N_3245,N_3443);
nor U3930 (N_3930,N_3448,N_3581);
or U3931 (N_3931,N_3375,N_3141);
nand U3932 (N_3932,N_3082,N_3208);
nor U3933 (N_3933,N_3465,N_3485);
nor U3934 (N_3934,N_3291,N_3481);
nor U3935 (N_3935,N_3599,N_3566);
nor U3936 (N_3936,N_3248,N_3445);
or U3937 (N_3937,N_3331,N_3268);
or U3938 (N_3938,N_3345,N_3516);
and U3939 (N_3939,N_3239,N_3052);
nor U3940 (N_3940,N_3488,N_3359);
nor U3941 (N_3941,N_3526,N_3568);
or U3942 (N_3942,N_3562,N_3037);
or U3943 (N_3943,N_3525,N_3402);
or U3944 (N_3944,N_3252,N_3423);
and U3945 (N_3945,N_3419,N_3379);
or U3946 (N_3946,N_3542,N_3366);
nand U3947 (N_3947,N_3511,N_3465);
nor U3948 (N_3948,N_3015,N_3059);
nand U3949 (N_3949,N_3555,N_3275);
nor U3950 (N_3950,N_3554,N_3306);
nor U3951 (N_3951,N_3043,N_3037);
or U3952 (N_3952,N_3387,N_3156);
nor U3953 (N_3953,N_3457,N_3321);
nand U3954 (N_3954,N_3544,N_3193);
and U3955 (N_3955,N_3123,N_3080);
and U3956 (N_3956,N_3417,N_3548);
or U3957 (N_3957,N_3094,N_3336);
nand U3958 (N_3958,N_3172,N_3500);
or U3959 (N_3959,N_3017,N_3304);
and U3960 (N_3960,N_3206,N_3429);
or U3961 (N_3961,N_3343,N_3490);
and U3962 (N_3962,N_3227,N_3483);
and U3963 (N_3963,N_3260,N_3132);
or U3964 (N_3964,N_3084,N_3111);
nor U3965 (N_3965,N_3471,N_3510);
or U3966 (N_3966,N_3343,N_3150);
nand U3967 (N_3967,N_3190,N_3459);
or U3968 (N_3968,N_3530,N_3339);
xnor U3969 (N_3969,N_3331,N_3300);
or U3970 (N_3970,N_3063,N_3504);
and U3971 (N_3971,N_3206,N_3087);
xor U3972 (N_3972,N_3352,N_3597);
or U3973 (N_3973,N_3478,N_3039);
and U3974 (N_3974,N_3383,N_3258);
and U3975 (N_3975,N_3424,N_3005);
and U3976 (N_3976,N_3077,N_3182);
xor U3977 (N_3977,N_3528,N_3449);
or U3978 (N_3978,N_3218,N_3572);
or U3979 (N_3979,N_3412,N_3348);
or U3980 (N_3980,N_3357,N_3541);
or U3981 (N_3981,N_3121,N_3140);
and U3982 (N_3982,N_3499,N_3145);
and U3983 (N_3983,N_3044,N_3218);
and U3984 (N_3984,N_3082,N_3414);
nand U3985 (N_3985,N_3595,N_3140);
or U3986 (N_3986,N_3309,N_3331);
and U3987 (N_3987,N_3428,N_3353);
nand U3988 (N_3988,N_3039,N_3258);
and U3989 (N_3989,N_3355,N_3265);
or U3990 (N_3990,N_3102,N_3161);
nor U3991 (N_3991,N_3439,N_3096);
xor U3992 (N_3992,N_3517,N_3553);
nor U3993 (N_3993,N_3285,N_3591);
nor U3994 (N_3994,N_3179,N_3560);
and U3995 (N_3995,N_3380,N_3570);
nand U3996 (N_3996,N_3497,N_3218);
nand U3997 (N_3997,N_3099,N_3327);
or U3998 (N_3998,N_3504,N_3414);
and U3999 (N_3999,N_3491,N_3181);
and U4000 (N_4000,N_3457,N_3268);
nand U4001 (N_4001,N_3524,N_3152);
and U4002 (N_4002,N_3367,N_3569);
or U4003 (N_4003,N_3155,N_3401);
and U4004 (N_4004,N_3011,N_3286);
xnor U4005 (N_4005,N_3441,N_3190);
nor U4006 (N_4006,N_3108,N_3349);
xnor U4007 (N_4007,N_3479,N_3173);
and U4008 (N_4008,N_3492,N_3033);
nor U4009 (N_4009,N_3064,N_3046);
nor U4010 (N_4010,N_3573,N_3333);
and U4011 (N_4011,N_3035,N_3163);
nor U4012 (N_4012,N_3469,N_3444);
nor U4013 (N_4013,N_3166,N_3193);
or U4014 (N_4014,N_3177,N_3077);
nor U4015 (N_4015,N_3498,N_3445);
nand U4016 (N_4016,N_3010,N_3477);
and U4017 (N_4017,N_3342,N_3596);
xor U4018 (N_4018,N_3197,N_3391);
nor U4019 (N_4019,N_3135,N_3417);
nor U4020 (N_4020,N_3310,N_3344);
or U4021 (N_4021,N_3353,N_3571);
nand U4022 (N_4022,N_3386,N_3340);
nor U4023 (N_4023,N_3127,N_3251);
and U4024 (N_4024,N_3387,N_3114);
or U4025 (N_4025,N_3165,N_3172);
or U4026 (N_4026,N_3528,N_3036);
or U4027 (N_4027,N_3279,N_3017);
nor U4028 (N_4028,N_3287,N_3453);
or U4029 (N_4029,N_3103,N_3070);
nand U4030 (N_4030,N_3005,N_3588);
nor U4031 (N_4031,N_3078,N_3150);
nand U4032 (N_4032,N_3137,N_3112);
xnor U4033 (N_4033,N_3537,N_3289);
or U4034 (N_4034,N_3127,N_3382);
or U4035 (N_4035,N_3542,N_3349);
nand U4036 (N_4036,N_3547,N_3260);
and U4037 (N_4037,N_3207,N_3336);
nand U4038 (N_4038,N_3535,N_3188);
and U4039 (N_4039,N_3375,N_3469);
and U4040 (N_4040,N_3355,N_3400);
or U4041 (N_4041,N_3580,N_3099);
nand U4042 (N_4042,N_3290,N_3047);
or U4043 (N_4043,N_3057,N_3395);
or U4044 (N_4044,N_3068,N_3389);
and U4045 (N_4045,N_3513,N_3595);
or U4046 (N_4046,N_3273,N_3548);
and U4047 (N_4047,N_3163,N_3169);
nand U4048 (N_4048,N_3360,N_3552);
nand U4049 (N_4049,N_3542,N_3179);
nor U4050 (N_4050,N_3006,N_3473);
or U4051 (N_4051,N_3391,N_3150);
nand U4052 (N_4052,N_3391,N_3336);
nor U4053 (N_4053,N_3115,N_3125);
and U4054 (N_4054,N_3057,N_3516);
nor U4055 (N_4055,N_3594,N_3062);
nand U4056 (N_4056,N_3074,N_3077);
or U4057 (N_4057,N_3312,N_3329);
and U4058 (N_4058,N_3574,N_3057);
nor U4059 (N_4059,N_3385,N_3451);
and U4060 (N_4060,N_3490,N_3383);
and U4061 (N_4061,N_3179,N_3033);
nor U4062 (N_4062,N_3472,N_3403);
and U4063 (N_4063,N_3357,N_3535);
nor U4064 (N_4064,N_3289,N_3044);
or U4065 (N_4065,N_3363,N_3038);
xnor U4066 (N_4066,N_3498,N_3508);
and U4067 (N_4067,N_3092,N_3275);
nand U4068 (N_4068,N_3119,N_3331);
or U4069 (N_4069,N_3018,N_3169);
nor U4070 (N_4070,N_3148,N_3439);
nor U4071 (N_4071,N_3018,N_3309);
nand U4072 (N_4072,N_3277,N_3549);
nand U4073 (N_4073,N_3246,N_3551);
nand U4074 (N_4074,N_3059,N_3374);
or U4075 (N_4075,N_3459,N_3246);
nand U4076 (N_4076,N_3086,N_3058);
nand U4077 (N_4077,N_3081,N_3027);
nor U4078 (N_4078,N_3000,N_3254);
and U4079 (N_4079,N_3561,N_3237);
or U4080 (N_4080,N_3558,N_3271);
or U4081 (N_4081,N_3136,N_3157);
nor U4082 (N_4082,N_3530,N_3519);
xor U4083 (N_4083,N_3434,N_3566);
nor U4084 (N_4084,N_3292,N_3308);
or U4085 (N_4085,N_3576,N_3593);
nand U4086 (N_4086,N_3099,N_3261);
nand U4087 (N_4087,N_3037,N_3381);
nand U4088 (N_4088,N_3219,N_3231);
or U4089 (N_4089,N_3234,N_3250);
and U4090 (N_4090,N_3444,N_3524);
xnor U4091 (N_4091,N_3260,N_3264);
or U4092 (N_4092,N_3194,N_3319);
or U4093 (N_4093,N_3192,N_3486);
nand U4094 (N_4094,N_3078,N_3505);
nor U4095 (N_4095,N_3113,N_3198);
or U4096 (N_4096,N_3385,N_3376);
and U4097 (N_4097,N_3315,N_3529);
and U4098 (N_4098,N_3228,N_3107);
and U4099 (N_4099,N_3380,N_3217);
nor U4100 (N_4100,N_3347,N_3328);
and U4101 (N_4101,N_3247,N_3023);
nor U4102 (N_4102,N_3568,N_3020);
nor U4103 (N_4103,N_3436,N_3062);
or U4104 (N_4104,N_3542,N_3505);
nor U4105 (N_4105,N_3562,N_3059);
nor U4106 (N_4106,N_3248,N_3398);
nor U4107 (N_4107,N_3345,N_3499);
or U4108 (N_4108,N_3287,N_3060);
nand U4109 (N_4109,N_3108,N_3263);
nand U4110 (N_4110,N_3266,N_3177);
or U4111 (N_4111,N_3098,N_3265);
nand U4112 (N_4112,N_3479,N_3566);
or U4113 (N_4113,N_3005,N_3586);
and U4114 (N_4114,N_3090,N_3052);
nand U4115 (N_4115,N_3389,N_3421);
or U4116 (N_4116,N_3364,N_3324);
nor U4117 (N_4117,N_3544,N_3442);
nand U4118 (N_4118,N_3515,N_3108);
and U4119 (N_4119,N_3451,N_3228);
or U4120 (N_4120,N_3186,N_3180);
nor U4121 (N_4121,N_3028,N_3020);
and U4122 (N_4122,N_3347,N_3093);
nand U4123 (N_4123,N_3068,N_3122);
and U4124 (N_4124,N_3592,N_3449);
or U4125 (N_4125,N_3041,N_3072);
or U4126 (N_4126,N_3235,N_3321);
nor U4127 (N_4127,N_3239,N_3542);
and U4128 (N_4128,N_3083,N_3587);
nand U4129 (N_4129,N_3045,N_3469);
or U4130 (N_4130,N_3349,N_3280);
or U4131 (N_4131,N_3268,N_3098);
nand U4132 (N_4132,N_3457,N_3110);
nor U4133 (N_4133,N_3383,N_3194);
or U4134 (N_4134,N_3085,N_3572);
nor U4135 (N_4135,N_3484,N_3557);
nor U4136 (N_4136,N_3276,N_3466);
nor U4137 (N_4137,N_3553,N_3280);
nor U4138 (N_4138,N_3536,N_3357);
nor U4139 (N_4139,N_3353,N_3371);
xnor U4140 (N_4140,N_3375,N_3240);
nor U4141 (N_4141,N_3358,N_3347);
nand U4142 (N_4142,N_3129,N_3407);
nor U4143 (N_4143,N_3463,N_3258);
or U4144 (N_4144,N_3278,N_3419);
xor U4145 (N_4145,N_3156,N_3312);
and U4146 (N_4146,N_3044,N_3454);
nor U4147 (N_4147,N_3515,N_3036);
and U4148 (N_4148,N_3323,N_3293);
or U4149 (N_4149,N_3531,N_3145);
nand U4150 (N_4150,N_3003,N_3506);
nor U4151 (N_4151,N_3415,N_3506);
or U4152 (N_4152,N_3089,N_3000);
nor U4153 (N_4153,N_3316,N_3186);
nand U4154 (N_4154,N_3053,N_3044);
xor U4155 (N_4155,N_3586,N_3473);
or U4156 (N_4156,N_3032,N_3553);
nor U4157 (N_4157,N_3203,N_3404);
nor U4158 (N_4158,N_3143,N_3031);
nor U4159 (N_4159,N_3125,N_3438);
or U4160 (N_4160,N_3443,N_3371);
and U4161 (N_4161,N_3136,N_3272);
nand U4162 (N_4162,N_3025,N_3387);
nor U4163 (N_4163,N_3378,N_3249);
nand U4164 (N_4164,N_3009,N_3498);
xor U4165 (N_4165,N_3551,N_3057);
nand U4166 (N_4166,N_3330,N_3577);
and U4167 (N_4167,N_3083,N_3492);
or U4168 (N_4168,N_3202,N_3313);
or U4169 (N_4169,N_3403,N_3557);
nand U4170 (N_4170,N_3565,N_3592);
or U4171 (N_4171,N_3364,N_3256);
nor U4172 (N_4172,N_3081,N_3135);
xnor U4173 (N_4173,N_3487,N_3366);
nand U4174 (N_4174,N_3598,N_3466);
or U4175 (N_4175,N_3070,N_3372);
nand U4176 (N_4176,N_3414,N_3441);
or U4177 (N_4177,N_3217,N_3331);
and U4178 (N_4178,N_3316,N_3480);
or U4179 (N_4179,N_3026,N_3524);
and U4180 (N_4180,N_3594,N_3036);
nor U4181 (N_4181,N_3426,N_3142);
nand U4182 (N_4182,N_3038,N_3412);
and U4183 (N_4183,N_3552,N_3149);
and U4184 (N_4184,N_3077,N_3426);
nor U4185 (N_4185,N_3148,N_3343);
and U4186 (N_4186,N_3383,N_3334);
or U4187 (N_4187,N_3163,N_3400);
and U4188 (N_4188,N_3472,N_3188);
xor U4189 (N_4189,N_3006,N_3164);
or U4190 (N_4190,N_3003,N_3409);
and U4191 (N_4191,N_3512,N_3491);
nor U4192 (N_4192,N_3214,N_3499);
nand U4193 (N_4193,N_3332,N_3144);
and U4194 (N_4194,N_3363,N_3034);
nor U4195 (N_4195,N_3090,N_3412);
and U4196 (N_4196,N_3045,N_3505);
xor U4197 (N_4197,N_3330,N_3272);
nor U4198 (N_4198,N_3341,N_3292);
nor U4199 (N_4199,N_3031,N_3067);
or U4200 (N_4200,N_3966,N_3717);
or U4201 (N_4201,N_3666,N_3801);
and U4202 (N_4202,N_3947,N_4134);
or U4203 (N_4203,N_3982,N_3798);
xnor U4204 (N_4204,N_3827,N_4067);
or U4205 (N_4205,N_3687,N_4135);
nor U4206 (N_4206,N_3726,N_3670);
nor U4207 (N_4207,N_4113,N_3774);
nand U4208 (N_4208,N_3880,N_3925);
or U4209 (N_4209,N_4138,N_3794);
nand U4210 (N_4210,N_3816,N_3958);
or U4211 (N_4211,N_3749,N_4165);
nor U4212 (N_4212,N_3693,N_3828);
and U4213 (N_4213,N_3865,N_4055);
nor U4214 (N_4214,N_3845,N_4192);
nor U4215 (N_4215,N_3876,N_3973);
nand U4216 (N_4216,N_3983,N_4058);
xor U4217 (N_4217,N_4176,N_3721);
and U4218 (N_4218,N_4167,N_3911);
nand U4219 (N_4219,N_3955,N_4140);
nand U4220 (N_4220,N_3644,N_3921);
xnor U4221 (N_4221,N_4129,N_4150);
or U4222 (N_4222,N_3641,N_3817);
or U4223 (N_4223,N_4152,N_4006);
and U4224 (N_4224,N_3919,N_3961);
and U4225 (N_4225,N_3942,N_3667);
nor U4226 (N_4226,N_3884,N_4062);
or U4227 (N_4227,N_4195,N_3682);
or U4228 (N_4228,N_4181,N_3710);
nand U4229 (N_4229,N_4002,N_4158);
and U4230 (N_4230,N_3993,N_4108);
or U4231 (N_4231,N_3661,N_3821);
nand U4232 (N_4232,N_3640,N_3875);
or U4233 (N_4233,N_3879,N_3643);
nand U4234 (N_4234,N_3986,N_3872);
nand U4235 (N_4235,N_3791,N_4091);
nand U4236 (N_4236,N_3658,N_3924);
and U4237 (N_4237,N_3752,N_3680);
nand U4238 (N_4238,N_4180,N_3810);
or U4239 (N_4239,N_3665,N_4066);
xnor U4240 (N_4240,N_4013,N_4096);
nor U4241 (N_4241,N_3807,N_4070);
and U4242 (N_4242,N_4123,N_4142);
xor U4243 (N_4243,N_3743,N_4056);
nor U4244 (N_4244,N_4071,N_4052);
and U4245 (N_4245,N_3606,N_4196);
nor U4246 (N_4246,N_4026,N_3716);
nand U4247 (N_4247,N_3762,N_4157);
and U4248 (N_4248,N_4080,N_3722);
nor U4249 (N_4249,N_3771,N_3824);
nor U4250 (N_4250,N_4049,N_3988);
nand U4251 (N_4251,N_3776,N_3852);
nor U4252 (N_4252,N_4128,N_3608);
nand U4253 (N_4253,N_3652,N_3873);
or U4254 (N_4254,N_3916,N_4190);
nand U4255 (N_4255,N_3618,N_4147);
and U4256 (N_4256,N_3938,N_3709);
or U4257 (N_4257,N_3883,N_3688);
and U4258 (N_4258,N_3907,N_4073);
nand U4259 (N_4259,N_3655,N_4044);
nand U4260 (N_4260,N_3702,N_3783);
nand U4261 (N_4261,N_4008,N_3874);
or U4262 (N_4262,N_3963,N_3900);
or U4263 (N_4263,N_3920,N_3839);
nand U4264 (N_4264,N_3788,N_4105);
or U4265 (N_4265,N_3645,N_3663);
nor U4266 (N_4266,N_3744,N_4098);
or U4267 (N_4267,N_3719,N_3782);
or U4268 (N_4268,N_3631,N_3893);
or U4269 (N_4269,N_3602,N_3601);
and U4270 (N_4270,N_3795,N_3979);
or U4271 (N_4271,N_4061,N_3648);
or U4272 (N_4272,N_4185,N_3755);
and U4273 (N_4273,N_4077,N_4125);
and U4274 (N_4274,N_3843,N_4145);
nand U4275 (N_4275,N_3844,N_3994);
and U4276 (N_4276,N_3818,N_4041);
and U4277 (N_4277,N_3895,N_4189);
and U4278 (N_4278,N_3838,N_3781);
nand U4279 (N_4279,N_4175,N_3713);
nor U4280 (N_4280,N_3909,N_4164);
or U4281 (N_4281,N_3703,N_3835);
nand U4282 (N_4282,N_3630,N_3615);
nor U4283 (N_4283,N_4017,N_4072);
or U4284 (N_4284,N_3625,N_4101);
and U4285 (N_4285,N_4115,N_3917);
nor U4286 (N_4286,N_4161,N_4160);
and U4287 (N_4287,N_4110,N_4036);
and U4288 (N_4288,N_3992,N_3674);
nor U4289 (N_4289,N_4112,N_3864);
and U4290 (N_4290,N_4075,N_3633);
and U4291 (N_4291,N_4102,N_3767);
and U4292 (N_4292,N_3662,N_4000);
nand U4293 (N_4293,N_4148,N_3940);
nand U4294 (N_4294,N_4114,N_3738);
and U4295 (N_4295,N_3996,N_3639);
or U4296 (N_4296,N_3811,N_3696);
nand U4297 (N_4297,N_4035,N_3737);
or U4298 (N_4298,N_3941,N_3734);
or U4299 (N_4299,N_3770,N_3851);
nand U4300 (N_4300,N_3636,N_3853);
nand U4301 (N_4301,N_4095,N_4116);
or U4302 (N_4302,N_3632,N_3977);
nand U4303 (N_4303,N_4172,N_4089);
or U4304 (N_4304,N_4100,N_4159);
and U4305 (N_4305,N_3678,N_3860);
and U4306 (N_4306,N_3745,N_4018);
nor U4307 (N_4307,N_3691,N_4076);
nor U4308 (N_4308,N_3624,N_3748);
nand U4309 (N_4309,N_3954,N_3899);
nor U4310 (N_4310,N_3764,N_3918);
and U4311 (N_4311,N_3929,N_3683);
or U4312 (N_4312,N_4069,N_3803);
nand U4313 (N_4313,N_3672,N_3820);
or U4314 (N_4314,N_4153,N_4126);
nand U4315 (N_4315,N_3765,N_3854);
or U4316 (N_4316,N_3711,N_3849);
nand U4317 (N_4317,N_3787,N_3987);
xor U4318 (N_4318,N_4179,N_3967);
nor U4319 (N_4319,N_3712,N_3891);
nor U4320 (N_4320,N_4020,N_4198);
and U4321 (N_4321,N_3769,N_4149);
nor U4322 (N_4322,N_3614,N_3877);
nand U4323 (N_4323,N_4107,N_3888);
or U4324 (N_4324,N_3964,N_3705);
nand U4325 (N_4325,N_3825,N_3904);
nand U4326 (N_4326,N_3786,N_3647);
or U4327 (N_4327,N_3778,N_4120);
or U4328 (N_4328,N_4169,N_3978);
nand U4329 (N_4329,N_3664,N_3905);
xor U4330 (N_4330,N_3708,N_3796);
nand U4331 (N_4331,N_3952,N_3815);
or U4332 (N_4332,N_4117,N_3707);
nor U4333 (N_4333,N_3960,N_4156);
and U4334 (N_4334,N_3841,N_4063);
nand U4335 (N_4335,N_3732,N_4038);
nor U4336 (N_4336,N_3866,N_3723);
or U4337 (N_4337,N_4048,N_3837);
nand U4338 (N_4338,N_4019,N_4182);
or U4339 (N_4339,N_4005,N_3830);
or U4340 (N_4340,N_3690,N_3740);
and U4341 (N_4341,N_3944,N_4022);
or U4342 (N_4342,N_3634,N_3646);
nor U4343 (N_4343,N_4121,N_3932);
and U4344 (N_4344,N_3689,N_3991);
nand U4345 (N_4345,N_3892,N_3981);
or U4346 (N_4346,N_3780,N_4193);
nor U4347 (N_4347,N_3651,N_3867);
or U4348 (N_4348,N_3603,N_4016);
or U4349 (N_4349,N_4111,N_3962);
or U4350 (N_4350,N_4074,N_4030);
and U4351 (N_4351,N_3701,N_4068);
and U4352 (N_4352,N_3971,N_3936);
nor U4353 (N_4353,N_3903,N_3735);
nor U4354 (N_4354,N_4003,N_3605);
nand U4355 (N_4355,N_3657,N_3659);
nor U4356 (N_4356,N_3746,N_3863);
nand U4357 (N_4357,N_3889,N_4133);
and U4358 (N_4358,N_4137,N_3747);
nand U4359 (N_4359,N_3751,N_4131);
nor U4360 (N_4360,N_3990,N_3935);
nand U4361 (N_4361,N_3676,N_3698);
or U4362 (N_4362,N_4104,N_4039);
or U4363 (N_4363,N_3914,N_4092);
nor U4364 (N_4364,N_4132,N_3706);
nor U4365 (N_4365,N_3937,N_4184);
or U4366 (N_4366,N_3896,N_3975);
nor U4367 (N_4367,N_3997,N_3612);
nand U4368 (N_4368,N_3730,N_4060);
nand U4369 (N_4369,N_3819,N_4014);
nor U4370 (N_4370,N_4094,N_3834);
xnor U4371 (N_4371,N_3831,N_3980);
nor U4372 (N_4372,N_3616,N_3793);
or U4373 (N_4373,N_3934,N_3842);
nand U4374 (N_4374,N_3861,N_4144);
nand U4375 (N_4375,N_3699,N_3802);
or U4376 (N_4376,N_3809,N_3731);
nor U4377 (N_4377,N_3733,N_3621);
nor U4378 (N_4378,N_4082,N_4043);
nand U4379 (N_4379,N_3859,N_3758);
nand U4380 (N_4380,N_3933,N_3804);
nand U4381 (N_4381,N_4032,N_3692);
and U4382 (N_4382,N_4154,N_3619);
and U4383 (N_4383,N_3926,N_4024);
nand U4384 (N_4384,N_3768,N_4177);
nor U4385 (N_4385,N_3972,N_4199);
and U4386 (N_4386,N_4197,N_4168);
nand U4387 (N_4387,N_4139,N_3650);
and U4388 (N_4388,N_3753,N_4188);
or U4389 (N_4389,N_3908,N_3976);
nor U4390 (N_4390,N_3974,N_4103);
nor U4391 (N_4391,N_3686,N_3846);
or U4392 (N_4392,N_3739,N_3999);
nand U4393 (N_4393,N_3777,N_3923);
nand U4394 (N_4394,N_3995,N_3829);
or U4395 (N_4395,N_3638,N_3789);
and U4396 (N_4396,N_4086,N_3985);
and U4397 (N_4397,N_3671,N_3617);
or U4398 (N_4398,N_3913,N_3669);
nor U4399 (N_4399,N_4045,N_3620);
and U4400 (N_4400,N_3953,N_3928);
nand U4401 (N_4401,N_4021,N_4109);
and U4402 (N_4402,N_3881,N_4033);
and U4403 (N_4403,N_3850,N_3931);
nand U4404 (N_4404,N_3681,N_4015);
nand U4405 (N_4405,N_3727,N_3922);
or U4406 (N_4406,N_3894,N_3906);
nand U4407 (N_4407,N_3660,N_3729);
nor U4408 (N_4408,N_3898,N_4143);
and U4409 (N_4409,N_3679,N_3998);
and U4410 (N_4410,N_3943,N_4023);
or U4411 (N_4411,N_4141,N_4031);
nor U4412 (N_4412,N_3642,N_3949);
nor U4413 (N_4413,N_4025,N_3628);
nor U4414 (N_4414,N_4053,N_3784);
or U4415 (N_4415,N_3622,N_3808);
xor U4416 (N_4416,N_3948,N_4059);
nand U4417 (N_4417,N_3959,N_3956);
nand U4418 (N_4418,N_3772,N_3653);
or U4419 (N_4419,N_3790,N_3609);
or U4420 (N_4420,N_4118,N_3763);
nand U4421 (N_4421,N_4124,N_3868);
xor U4422 (N_4422,N_3623,N_4012);
and U4423 (N_4423,N_4088,N_4064);
or U4424 (N_4424,N_4065,N_4079);
or U4425 (N_4425,N_4083,N_3946);
and U4426 (N_4426,N_4054,N_3945);
and U4427 (N_4427,N_4084,N_3607);
or U4428 (N_4428,N_4011,N_3950);
and U4429 (N_4429,N_3858,N_3969);
nand U4430 (N_4430,N_3741,N_4163);
nand U4431 (N_4431,N_3797,N_3910);
and U4432 (N_4432,N_3742,N_3890);
or U4433 (N_4433,N_4001,N_3814);
nor U4434 (N_4434,N_4042,N_4155);
nor U4435 (N_4435,N_3965,N_3856);
and U4436 (N_4436,N_3759,N_4047);
or U4437 (N_4437,N_3968,N_3757);
nor U4438 (N_4438,N_3887,N_3761);
nand U4439 (N_4439,N_4183,N_4146);
nand U4440 (N_4440,N_3600,N_3832);
nand U4441 (N_4441,N_3870,N_3800);
nand U4442 (N_4442,N_3626,N_3927);
and U4443 (N_4443,N_4170,N_4097);
or U4444 (N_4444,N_4093,N_3792);
and U4445 (N_4445,N_3754,N_4166);
and U4446 (N_4446,N_3613,N_3812);
and U4447 (N_4447,N_4004,N_4040);
and U4448 (N_4448,N_4037,N_3848);
nor U4449 (N_4449,N_4171,N_4162);
nor U4450 (N_4450,N_4173,N_4085);
or U4451 (N_4451,N_3649,N_3885);
nor U4452 (N_4452,N_4187,N_4151);
and U4453 (N_4453,N_3654,N_3715);
nor U4454 (N_4454,N_4078,N_3840);
nand U4455 (N_4455,N_3984,N_3951);
nor U4456 (N_4456,N_3704,N_4127);
nand U4457 (N_4457,N_3823,N_3799);
nor U4458 (N_4458,N_3882,N_3750);
nand U4459 (N_4459,N_3813,N_3656);
nand U4460 (N_4460,N_4090,N_4130);
nor U4461 (N_4461,N_4106,N_3836);
nand U4462 (N_4462,N_4051,N_3912);
nand U4463 (N_4463,N_3668,N_4050);
nor U4464 (N_4464,N_3635,N_3610);
and U4465 (N_4465,N_3637,N_3939);
or U4466 (N_4466,N_3902,N_4119);
nand U4467 (N_4467,N_3736,N_4029);
nor U4468 (N_4468,N_3833,N_3694);
nand U4469 (N_4469,N_4057,N_3970);
nor U4470 (N_4470,N_4178,N_3847);
and U4471 (N_4471,N_3611,N_4009);
or U4472 (N_4472,N_3766,N_3857);
xor U4473 (N_4473,N_3930,N_4046);
or U4474 (N_4474,N_3673,N_3855);
nor U4475 (N_4475,N_3806,N_4081);
and U4476 (N_4476,N_4136,N_4194);
or U4477 (N_4477,N_4122,N_4027);
and U4478 (N_4478,N_3728,N_3901);
and U4479 (N_4479,N_3862,N_3714);
nand U4480 (N_4480,N_4099,N_3675);
or U4481 (N_4481,N_3700,N_3957);
and U4482 (N_4482,N_3760,N_3886);
and U4483 (N_4483,N_3878,N_3718);
and U4484 (N_4484,N_4007,N_3604);
nor U4485 (N_4485,N_4034,N_3779);
or U4486 (N_4486,N_3871,N_3915);
nor U4487 (N_4487,N_3695,N_3627);
nor U4488 (N_4488,N_3826,N_3775);
nand U4489 (N_4489,N_3684,N_3773);
nor U4490 (N_4490,N_3822,N_3720);
or U4491 (N_4491,N_3989,N_4186);
nand U4492 (N_4492,N_4010,N_4191);
or U4493 (N_4493,N_3869,N_3629);
or U4494 (N_4494,N_3785,N_3685);
or U4495 (N_4495,N_3756,N_3897);
nand U4496 (N_4496,N_4028,N_3724);
nand U4497 (N_4497,N_3725,N_3805);
or U4498 (N_4498,N_3677,N_4174);
and U4499 (N_4499,N_3697,N_4087);
or U4500 (N_4500,N_3759,N_3610);
and U4501 (N_4501,N_4150,N_3889);
nor U4502 (N_4502,N_3739,N_3890);
nor U4503 (N_4503,N_3963,N_3679);
or U4504 (N_4504,N_3814,N_3669);
and U4505 (N_4505,N_3705,N_3860);
or U4506 (N_4506,N_3922,N_3822);
or U4507 (N_4507,N_3605,N_4180);
and U4508 (N_4508,N_3746,N_4054);
nand U4509 (N_4509,N_4081,N_3913);
and U4510 (N_4510,N_4029,N_3847);
nor U4511 (N_4511,N_4066,N_4042);
nand U4512 (N_4512,N_3637,N_4146);
or U4513 (N_4513,N_4101,N_4032);
and U4514 (N_4514,N_4048,N_3905);
and U4515 (N_4515,N_4139,N_3987);
and U4516 (N_4516,N_3604,N_4140);
or U4517 (N_4517,N_4088,N_3618);
nor U4518 (N_4518,N_3638,N_3628);
and U4519 (N_4519,N_3619,N_4043);
xor U4520 (N_4520,N_3850,N_3797);
and U4521 (N_4521,N_3732,N_4065);
nand U4522 (N_4522,N_3829,N_3840);
nor U4523 (N_4523,N_3906,N_3860);
nand U4524 (N_4524,N_3702,N_3630);
and U4525 (N_4525,N_3928,N_3635);
nand U4526 (N_4526,N_4075,N_3774);
and U4527 (N_4527,N_3622,N_3926);
and U4528 (N_4528,N_3876,N_3807);
nand U4529 (N_4529,N_4147,N_4084);
nor U4530 (N_4530,N_3890,N_3897);
nor U4531 (N_4531,N_3665,N_3980);
and U4532 (N_4532,N_3804,N_3838);
or U4533 (N_4533,N_3901,N_4078);
nor U4534 (N_4534,N_3624,N_3815);
nor U4535 (N_4535,N_4125,N_3842);
nand U4536 (N_4536,N_3866,N_4025);
nor U4537 (N_4537,N_3945,N_3811);
nor U4538 (N_4538,N_3723,N_4195);
nand U4539 (N_4539,N_3704,N_3953);
nand U4540 (N_4540,N_4185,N_4003);
or U4541 (N_4541,N_3677,N_4183);
nand U4542 (N_4542,N_4037,N_3741);
nand U4543 (N_4543,N_3647,N_4078);
nand U4544 (N_4544,N_3749,N_3725);
nand U4545 (N_4545,N_3750,N_3619);
or U4546 (N_4546,N_3883,N_3651);
nand U4547 (N_4547,N_4007,N_3936);
nand U4548 (N_4548,N_4171,N_3866);
or U4549 (N_4549,N_3612,N_3802);
nor U4550 (N_4550,N_3767,N_3825);
nand U4551 (N_4551,N_4082,N_4121);
nand U4552 (N_4552,N_3866,N_3971);
or U4553 (N_4553,N_3848,N_4057);
xor U4554 (N_4554,N_3705,N_4074);
and U4555 (N_4555,N_3956,N_3756);
nand U4556 (N_4556,N_3717,N_3879);
and U4557 (N_4557,N_3888,N_3703);
and U4558 (N_4558,N_4090,N_4135);
nor U4559 (N_4559,N_3855,N_4024);
nand U4560 (N_4560,N_3615,N_3921);
or U4561 (N_4561,N_4051,N_3610);
and U4562 (N_4562,N_4110,N_3713);
nor U4563 (N_4563,N_3759,N_3639);
nor U4564 (N_4564,N_3672,N_3661);
nor U4565 (N_4565,N_3927,N_3669);
nor U4566 (N_4566,N_4129,N_3629);
and U4567 (N_4567,N_3651,N_3881);
or U4568 (N_4568,N_4181,N_3971);
and U4569 (N_4569,N_3705,N_3770);
nand U4570 (N_4570,N_4050,N_3984);
or U4571 (N_4571,N_4147,N_3625);
nand U4572 (N_4572,N_4075,N_3870);
and U4573 (N_4573,N_3829,N_4091);
and U4574 (N_4574,N_3925,N_3998);
or U4575 (N_4575,N_3820,N_4159);
nor U4576 (N_4576,N_3910,N_4120);
nand U4577 (N_4577,N_4066,N_3789);
nand U4578 (N_4578,N_4060,N_4199);
nand U4579 (N_4579,N_3950,N_4041);
nor U4580 (N_4580,N_3639,N_3683);
nor U4581 (N_4581,N_3779,N_3930);
and U4582 (N_4582,N_3684,N_4035);
nand U4583 (N_4583,N_4010,N_4058);
or U4584 (N_4584,N_3687,N_4157);
nand U4585 (N_4585,N_3937,N_4171);
nor U4586 (N_4586,N_4176,N_4083);
or U4587 (N_4587,N_3620,N_3960);
nor U4588 (N_4588,N_3840,N_4026);
or U4589 (N_4589,N_4030,N_4111);
or U4590 (N_4590,N_3731,N_4035);
nand U4591 (N_4591,N_3729,N_3972);
nand U4592 (N_4592,N_3806,N_3714);
nor U4593 (N_4593,N_3949,N_4096);
and U4594 (N_4594,N_3683,N_3630);
nand U4595 (N_4595,N_3941,N_3738);
nor U4596 (N_4596,N_3809,N_4113);
nand U4597 (N_4597,N_3682,N_4109);
and U4598 (N_4598,N_3618,N_4139);
or U4599 (N_4599,N_4041,N_4072);
xnor U4600 (N_4600,N_3602,N_3938);
xor U4601 (N_4601,N_3720,N_3661);
and U4602 (N_4602,N_3894,N_3849);
nand U4603 (N_4603,N_3652,N_3865);
nand U4604 (N_4604,N_3769,N_3767);
or U4605 (N_4605,N_4064,N_3694);
or U4606 (N_4606,N_3622,N_3798);
or U4607 (N_4607,N_3613,N_3708);
and U4608 (N_4608,N_4159,N_3821);
or U4609 (N_4609,N_3737,N_3704);
and U4610 (N_4610,N_3972,N_3933);
or U4611 (N_4611,N_3981,N_3961);
nor U4612 (N_4612,N_3919,N_3766);
or U4613 (N_4613,N_3862,N_3742);
nor U4614 (N_4614,N_4009,N_4044);
and U4615 (N_4615,N_3896,N_4155);
nor U4616 (N_4616,N_3751,N_3722);
nor U4617 (N_4617,N_3964,N_3627);
or U4618 (N_4618,N_3824,N_3710);
xor U4619 (N_4619,N_4164,N_3787);
nand U4620 (N_4620,N_4111,N_3991);
nand U4621 (N_4621,N_4102,N_4172);
or U4622 (N_4622,N_3840,N_3965);
or U4623 (N_4623,N_4064,N_4040);
or U4624 (N_4624,N_3977,N_4008);
nor U4625 (N_4625,N_3961,N_4066);
and U4626 (N_4626,N_4131,N_4038);
nand U4627 (N_4627,N_3700,N_3940);
nand U4628 (N_4628,N_4105,N_4141);
and U4629 (N_4629,N_3851,N_3679);
or U4630 (N_4630,N_4168,N_4049);
nor U4631 (N_4631,N_4045,N_4145);
or U4632 (N_4632,N_3931,N_4116);
nor U4633 (N_4633,N_3690,N_4143);
nand U4634 (N_4634,N_3669,N_4106);
and U4635 (N_4635,N_3808,N_3654);
nor U4636 (N_4636,N_3725,N_3947);
or U4637 (N_4637,N_3922,N_4011);
and U4638 (N_4638,N_3711,N_4105);
and U4639 (N_4639,N_3953,N_3613);
and U4640 (N_4640,N_4092,N_3673);
nor U4641 (N_4641,N_3961,N_4097);
or U4642 (N_4642,N_3952,N_3606);
nor U4643 (N_4643,N_4070,N_3667);
and U4644 (N_4644,N_3654,N_4013);
nor U4645 (N_4645,N_3918,N_3844);
or U4646 (N_4646,N_3704,N_4069);
or U4647 (N_4647,N_4040,N_4054);
and U4648 (N_4648,N_3817,N_3802);
nand U4649 (N_4649,N_4058,N_3831);
nand U4650 (N_4650,N_4005,N_4031);
or U4651 (N_4651,N_3688,N_3797);
nor U4652 (N_4652,N_4085,N_4167);
nand U4653 (N_4653,N_3711,N_3725);
or U4654 (N_4654,N_4126,N_4124);
nand U4655 (N_4655,N_3798,N_3659);
nor U4656 (N_4656,N_3710,N_4160);
and U4657 (N_4657,N_4180,N_3890);
and U4658 (N_4658,N_4106,N_3703);
or U4659 (N_4659,N_4119,N_4031);
and U4660 (N_4660,N_3728,N_3788);
xnor U4661 (N_4661,N_3779,N_3859);
and U4662 (N_4662,N_3891,N_3829);
and U4663 (N_4663,N_3749,N_3964);
nand U4664 (N_4664,N_3884,N_3659);
or U4665 (N_4665,N_4106,N_4112);
nor U4666 (N_4666,N_4088,N_4083);
nor U4667 (N_4667,N_4111,N_4001);
nand U4668 (N_4668,N_3934,N_3837);
or U4669 (N_4669,N_4180,N_3842);
nand U4670 (N_4670,N_4034,N_3656);
and U4671 (N_4671,N_4066,N_3855);
or U4672 (N_4672,N_3948,N_4027);
and U4673 (N_4673,N_3934,N_3960);
nand U4674 (N_4674,N_4132,N_3858);
nor U4675 (N_4675,N_3820,N_3808);
and U4676 (N_4676,N_4129,N_3813);
nand U4677 (N_4677,N_3973,N_3777);
nor U4678 (N_4678,N_4082,N_3925);
nand U4679 (N_4679,N_3699,N_4140);
nand U4680 (N_4680,N_4134,N_3747);
nor U4681 (N_4681,N_3983,N_3719);
or U4682 (N_4682,N_3762,N_3745);
nand U4683 (N_4683,N_3800,N_3926);
or U4684 (N_4684,N_4053,N_3601);
nand U4685 (N_4685,N_3990,N_3974);
nand U4686 (N_4686,N_3991,N_3723);
nor U4687 (N_4687,N_3626,N_4106);
or U4688 (N_4688,N_3997,N_4083);
or U4689 (N_4689,N_3659,N_3743);
nor U4690 (N_4690,N_3668,N_4198);
and U4691 (N_4691,N_3733,N_3941);
nor U4692 (N_4692,N_4147,N_4024);
or U4693 (N_4693,N_4159,N_3830);
nor U4694 (N_4694,N_4098,N_3955);
xnor U4695 (N_4695,N_3874,N_3669);
nand U4696 (N_4696,N_3695,N_4145);
nor U4697 (N_4697,N_3844,N_4109);
xor U4698 (N_4698,N_4041,N_3639);
or U4699 (N_4699,N_3786,N_3695);
and U4700 (N_4700,N_3875,N_3735);
nand U4701 (N_4701,N_3875,N_3883);
nand U4702 (N_4702,N_3954,N_3787);
nand U4703 (N_4703,N_3769,N_3751);
nor U4704 (N_4704,N_4044,N_4094);
nor U4705 (N_4705,N_4100,N_3936);
nand U4706 (N_4706,N_3620,N_4057);
and U4707 (N_4707,N_3939,N_3815);
nor U4708 (N_4708,N_4095,N_3877);
and U4709 (N_4709,N_4070,N_4106);
and U4710 (N_4710,N_3671,N_4027);
and U4711 (N_4711,N_3734,N_4064);
nand U4712 (N_4712,N_4064,N_3865);
or U4713 (N_4713,N_4057,N_3925);
nand U4714 (N_4714,N_3977,N_3931);
or U4715 (N_4715,N_3669,N_3763);
or U4716 (N_4716,N_3964,N_4028);
and U4717 (N_4717,N_4128,N_3935);
or U4718 (N_4718,N_3843,N_3801);
or U4719 (N_4719,N_3612,N_3664);
or U4720 (N_4720,N_3696,N_3820);
and U4721 (N_4721,N_3902,N_4122);
nor U4722 (N_4722,N_3974,N_4188);
nor U4723 (N_4723,N_3688,N_4034);
nand U4724 (N_4724,N_3628,N_4171);
or U4725 (N_4725,N_4152,N_3617);
nand U4726 (N_4726,N_3792,N_3907);
or U4727 (N_4727,N_3624,N_4044);
and U4728 (N_4728,N_4078,N_4157);
or U4729 (N_4729,N_3790,N_3765);
nor U4730 (N_4730,N_3833,N_3934);
and U4731 (N_4731,N_3814,N_4119);
nand U4732 (N_4732,N_3620,N_3612);
nand U4733 (N_4733,N_3679,N_3958);
and U4734 (N_4734,N_3602,N_3611);
nor U4735 (N_4735,N_4002,N_4159);
nand U4736 (N_4736,N_3839,N_4042);
nand U4737 (N_4737,N_4149,N_3699);
or U4738 (N_4738,N_3853,N_4194);
nor U4739 (N_4739,N_3777,N_4021);
nand U4740 (N_4740,N_4140,N_3770);
nand U4741 (N_4741,N_3729,N_3620);
nand U4742 (N_4742,N_4066,N_4024);
or U4743 (N_4743,N_4033,N_4101);
nand U4744 (N_4744,N_4016,N_3763);
nor U4745 (N_4745,N_3679,N_3896);
nand U4746 (N_4746,N_4193,N_4025);
and U4747 (N_4747,N_3963,N_3930);
or U4748 (N_4748,N_4080,N_3725);
and U4749 (N_4749,N_3751,N_3681);
nor U4750 (N_4750,N_4107,N_4114);
nand U4751 (N_4751,N_3945,N_4050);
nor U4752 (N_4752,N_4090,N_3948);
and U4753 (N_4753,N_3737,N_3968);
nand U4754 (N_4754,N_3803,N_3836);
and U4755 (N_4755,N_3816,N_4110);
nand U4756 (N_4756,N_3602,N_3867);
nand U4757 (N_4757,N_4044,N_3869);
nor U4758 (N_4758,N_4140,N_4150);
or U4759 (N_4759,N_4134,N_3849);
and U4760 (N_4760,N_3746,N_4195);
and U4761 (N_4761,N_3789,N_3954);
nand U4762 (N_4762,N_4007,N_3803);
or U4763 (N_4763,N_3824,N_4194);
and U4764 (N_4764,N_4170,N_3929);
or U4765 (N_4765,N_3953,N_3973);
nand U4766 (N_4766,N_4019,N_3948);
or U4767 (N_4767,N_3639,N_3625);
and U4768 (N_4768,N_3792,N_4000);
or U4769 (N_4769,N_4108,N_3714);
nor U4770 (N_4770,N_4043,N_3940);
and U4771 (N_4771,N_3744,N_4069);
and U4772 (N_4772,N_3956,N_3796);
or U4773 (N_4773,N_4057,N_4179);
xnor U4774 (N_4774,N_3887,N_3657);
nand U4775 (N_4775,N_4072,N_3950);
or U4776 (N_4776,N_3801,N_4185);
and U4777 (N_4777,N_3635,N_4036);
nor U4778 (N_4778,N_3922,N_4088);
or U4779 (N_4779,N_3873,N_4109);
nor U4780 (N_4780,N_4015,N_4039);
and U4781 (N_4781,N_3792,N_3761);
nor U4782 (N_4782,N_3997,N_4086);
or U4783 (N_4783,N_4173,N_3970);
and U4784 (N_4784,N_3659,N_3964);
and U4785 (N_4785,N_3649,N_3655);
or U4786 (N_4786,N_4113,N_3968);
nand U4787 (N_4787,N_3769,N_3962);
nor U4788 (N_4788,N_3956,N_3640);
nand U4789 (N_4789,N_3770,N_4114);
and U4790 (N_4790,N_4196,N_3943);
or U4791 (N_4791,N_3904,N_3636);
nand U4792 (N_4792,N_3716,N_3835);
nand U4793 (N_4793,N_3672,N_3861);
nand U4794 (N_4794,N_3828,N_3696);
or U4795 (N_4795,N_4114,N_3674);
or U4796 (N_4796,N_3972,N_4023);
or U4797 (N_4797,N_4089,N_3624);
or U4798 (N_4798,N_3795,N_4000);
nand U4799 (N_4799,N_3626,N_3756);
and U4800 (N_4800,N_4245,N_4602);
and U4801 (N_4801,N_4678,N_4405);
or U4802 (N_4802,N_4365,N_4780);
or U4803 (N_4803,N_4616,N_4227);
and U4804 (N_4804,N_4325,N_4549);
nor U4805 (N_4805,N_4640,N_4622);
and U4806 (N_4806,N_4217,N_4387);
nor U4807 (N_4807,N_4313,N_4503);
or U4808 (N_4808,N_4257,N_4258);
and U4809 (N_4809,N_4322,N_4215);
nor U4810 (N_4810,N_4551,N_4564);
or U4811 (N_4811,N_4440,N_4455);
nand U4812 (N_4812,N_4472,N_4766);
or U4813 (N_4813,N_4438,N_4691);
nor U4814 (N_4814,N_4483,N_4441);
or U4815 (N_4815,N_4666,N_4637);
and U4816 (N_4816,N_4231,N_4315);
nand U4817 (N_4817,N_4728,N_4534);
nand U4818 (N_4818,N_4388,N_4461);
xor U4819 (N_4819,N_4497,N_4372);
nand U4820 (N_4820,N_4307,N_4779);
or U4821 (N_4821,N_4479,N_4722);
or U4822 (N_4822,N_4758,N_4341);
nand U4823 (N_4823,N_4799,N_4788);
nand U4824 (N_4824,N_4792,N_4273);
nand U4825 (N_4825,N_4287,N_4264);
and U4826 (N_4826,N_4267,N_4517);
nor U4827 (N_4827,N_4422,N_4467);
nor U4828 (N_4828,N_4255,N_4567);
nand U4829 (N_4829,N_4796,N_4425);
nand U4830 (N_4830,N_4574,N_4716);
or U4831 (N_4831,N_4228,N_4401);
nor U4832 (N_4832,N_4571,N_4458);
and U4833 (N_4833,N_4777,N_4703);
nand U4834 (N_4834,N_4765,N_4488);
nor U4835 (N_4835,N_4558,N_4721);
nand U4836 (N_4836,N_4394,N_4414);
nand U4837 (N_4837,N_4545,N_4668);
and U4838 (N_4838,N_4331,N_4709);
and U4839 (N_4839,N_4452,N_4300);
and U4840 (N_4840,N_4206,N_4630);
or U4841 (N_4841,N_4573,N_4533);
or U4842 (N_4842,N_4363,N_4595);
nand U4843 (N_4843,N_4278,N_4229);
nor U4844 (N_4844,N_4554,N_4544);
nand U4845 (N_4845,N_4220,N_4644);
nor U4846 (N_4846,N_4239,N_4606);
and U4847 (N_4847,N_4738,N_4795);
or U4848 (N_4848,N_4759,N_4403);
and U4849 (N_4849,N_4762,N_4456);
nor U4850 (N_4850,N_4211,N_4499);
nor U4851 (N_4851,N_4661,N_4782);
nand U4852 (N_4852,N_4601,N_4240);
and U4853 (N_4853,N_4619,N_4726);
or U4854 (N_4854,N_4581,N_4326);
nor U4855 (N_4855,N_4706,N_4731);
or U4856 (N_4856,N_4495,N_4282);
or U4857 (N_4857,N_4344,N_4279);
or U4858 (N_4858,N_4340,N_4643);
or U4859 (N_4859,N_4646,N_4633);
nor U4860 (N_4860,N_4310,N_4512);
xor U4861 (N_4861,N_4547,N_4419);
nor U4862 (N_4862,N_4358,N_4289);
nand U4863 (N_4863,N_4757,N_4711);
nand U4864 (N_4864,N_4409,N_4397);
nor U4865 (N_4865,N_4755,N_4271);
or U4866 (N_4866,N_4244,N_4481);
or U4867 (N_4867,N_4689,N_4348);
or U4868 (N_4868,N_4254,N_4510);
or U4869 (N_4869,N_4433,N_4507);
or U4870 (N_4870,N_4587,N_4210);
xor U4871 (N_4871,N_4505,N_4690);
nor U4872 (N_4872,N_4377,N_4687);
nand U4873 (N_4873,N_4626,N_4418);
or U4874 (N_4874,N_4724,N_4489);
nand U4875 (N_4875,N_4203,N_4527);
nor U4876 (N_4876,N_4209,N_4761);
nand U4877 (N_4877,N_4454,N_4775);
nor U4878 (N_4878,N_4566,N_4311);
nor U4879 (N_4879,N_4304,N_4241);
or U4880 (N_4880,N_4540,N_4599);
xnor U4881 (N_4881,N_4374,N_4727);
nor U4882 (N_4882,N_4539,N_4280);
or U4883 (N_4883,N_4371,N_4362);
nand U4884 (N_4884,N_4265,N_4589);
nor U4885 (N_4885,N_4500,N_4338);
and U4886 (N_4886,N_4443,N_4222);
or U4887 (N_4887,N_4747,N_4491);
or U4888 (N_4888,N_4426,N_4615);
nor U4889 (N_4889,N_4445,N_4671);
nand U4890 (N_4890,N_4327,N_4786);
or U4891 (N_4891,N_4218,N_4552);
or U4892 (N_4892,N_4612,N_4314);
or U4893 (N_4893,N_4553,N_4675);
nand U4894 (N_4894,N_4350,N_4238);
or U4895 (N_4895,N_4578,N_4369);
nand U4896 (N_4896,N_4763,N_4519);
nand U4897 (N_4897,N_4743,N_4502);
nor U4898 (N_4898,N_4442,N_4476);
and U4899 (N_4899,N_4748,N_4657);
or U4900 (N_4900,N_4773,N_4337);
nand U4901 (N_4901,N_4734,N_4555);
nor U4902 (N_4902,N_4754,N_4610);
nor U4903 (N_4903,N_4439,N_4592);
nor U4904 (N_4904,N_4404,N_4660);
nor U4905 (N_4905,N_4434,N_4576);
and U4906 (N_4906,N_4309,N_4712);
or U4907 (N_4907,N_4291,N_4431);
and U4908 (N_4908,N_4583,N_4334);
nand U4909 (N_4909,N_4778,N_4694);
nand U4910 (N_4910,N_4375,N_4333);
nand U4911 (N_4911,N_4276,N_4723);
nand U4912 (N_4912,N_4312,N_4353);
nor U4913 (N_4913,N_4641,N_4355);
and U4914 (N_4914,N_4597,N_4432);
nand U4915 (N_4915,N_4477,N_4319);
nor U4916 (N_4916,N_4275,N_4525);
and U4917 (N_4917,N_4474,N_4624);
and U4918 (N_4918,N_4396,N_4769);
nor U4919 (N_4919,N_4774,N_4223);
nor U4920 (N_4920,N_4294,N_4707);
or U4921 (N_4921,N_4794,N_4647);
nand U4922 (N_4922,N_4412,N_4580);
and U4923 (N_4923,N_4532,N_4277);
and U4924 (N_4924,N_4357,N_4650);
nor U4925 (N_4925,N_4680,N_4339);
or U4926 (N_4926,N_4760,N_4674);
nor U4927 (N_4927,N_4494,N_4705);
or U4928 (N_4928,N_4586,N_4613);
and U4929 (N_4929,N_4746,N_4214);
xnor U4930 (N_4930,N_4569,N_4410);
and U4931 (N_4931,N_4430,N_4618);
and U4932 (N_4932,N_4306,N_4336);
nand U4933 (N_4933,N_4603,N_4305);
nor U4934 (N_4934,N_4234,N_4684);
or U4935 (N_4935,N_4537,N_4465);
or U4936 (N_4936,N_4484,N_4744);
nor U4937 (N_4937,N_4635,N_4560);
or U4938 (N_4938,N_4283,N_4688);
nor U4939 (N_4939,N_4368,N_4207);
and U4940 (N_4940,N_4463,N_4253);
and U4941 (N_4941,N_4400,N_4714);
and U4942 (N_4942,N_4208,N_4632);
or U4943 (N_4943,N_4679,N_4642);
nor U4944 (N_4944,N_4729,N_4598);
and U4945 (N_4945,N_4732,N_4563);
and U4946 (N_4946,N_4511,N_4478);
nor U4947 (N_4947,N_4570,N_4296);
nor U4948 (N_4948,N_4733,N_4740);
nor U4949 (N_4949,N_4367,N_4685);
nor U4950 (N_4950,N_4346,N_4324);
nor U4951 (N_4951,N_4770,N_4379);
nand U4952 (N_4952,N_4509,N_4683);
and U4953 (N_4953,N_4390,N_4793);
nor U4954 (N_4954,N_4750,N_4493);
or U4955 (N_4955,N_4235,N_4708);
nor U4956 (N_4956,N_4428,N_4295);
nor U4957 (N_4957,N_4411,N_4669);
nor U4958 (N_4958,N_4261,N_4415);
nor U4959 (N_4959,N_4392,N_4787);
nor U4960 (N_4960,N_4652,N_4219);
and U4961 (N_4961,N_4715,N_4359);
and U4962 (N_4962,N_4204,N_4764);
nor U4963 (N_4963,N_4343,N_4631);
and U4964 (N_4964,N_4444,N_4473);
nand U4965 (N_4965,N_4676,N_4656);
nand U4966 (N_4966,N_4704,N_4538);
or U4967 (N_4967,N_4698,N_4789);
or U4968 (N_4968,N_4243,N_4528);
and U4969 (N_4969,N_4742,N_4262);
nor U4970 (N_4970,N_4585,N_4356);
or U4971 (N_4971,N_4516,N_4249);
xnor U4972 (N_4972,N_4301,N_4471);
or U4973 (N_4973,N_4508,N_4591);
or U4974 (N_4974,N_4201,N_4424);
and U4975 (N_4975,N_4783,N_4651);
and U4976 (N_4976,N_4741,N_4448);
and U4977 (N_4977,N_4216,N_4720);
or U4978 (N_4978,N_4634,N_4446);
nand U4979 (N_4979,N_4590,N_4237);
nand U4980 (N_4980,N_4614,N_4274);
and U4981 (N_4981,N_4272,N_4791);
nand U4982 (N_4982,N_4475,N_4224);
and U4983 (N_4983,N_4332,N_4308);
and U4984 (N_4984,N_4559,N_4482);
nor U4985 (N_4985,N_4719,N_4772);
nand U4986 (N_4986,N_4385,N_4342);
nor U4987 (N_4987,N_4462,N_4609);
nand U4988 (N_4988,N_4451,N_4468);
nor U4989 (N_4989,N_4692,N_4370);
nand U4990 (N_4990,N_4546,N_4399);
and U4991 (N_4991,N_4556,N_4548);
and U4992 (N_4992,N_4349,N_4212);
nor U4993 (N_4993,N_4436,N_4663);
and U4994 (N_4994,N_4501,N_4594);
nor U4995 (N_4995,N_4513,N_4607);
or U4996 (N_4996,N_4485,N_4629);
or U4997 (N_4997,N_4250,N_4298);
or U4998 (N_4998,N_4604,N_4466);
nand U4999 (N_4999,N_4449,N_4579);
nand U5000 (N_5000,N_4284,N_4395);
xor U5001 (N_5001,N_4328,N_4389);
nand U5002 (N_5002,N_4246,N_4596);
and U5003 (N_5003,N_4673,N_4302);
nor U5004 (N_5004,N_4316,N_4251);
and U5005 (N_5005,N_4515,N_4730);
nor U5006 (N_5006,N_4520,N_4423);
nand U5007 (N_5007,N_4628,N_4713);
nor U5008 (N_5008,N_4259,N_4470);
or U5009 (N_5009,N_4506,N_4330);
nor U5010 (N_5010,N_4384,N_4320);
or U5011 (N_5011,N_4364,N_4699);
nor U5012 (N_5012,N_4236,N_4286);
nand U5013 (N_5013,N_4736,N_4450);
nor U5014 (N_5014,N_4568,N_4625);
or U5015 (N_5015,N_4266,N_4526);
nand U5016 (N_5016,N_4268,N_4248);
nor U5017 (N_5017,N_4664,N_4753);
nor U5018 (N_5018,N_4514,N_4351);
nor U5019 (N_5019,N_4781,N_4784);
nand U5020 (N_5020,N_4751,N_4281);
and U5021 (N_5021,N_4407,N_4393);
and U5022 (N_5022,N_4670,N_4608);
nand U5023 (N_5023,N_4260,N_4297);
or U5024 (N_5024,N_4557,N_4427);
or U5025 (N_5025,N_4398,N_4459);
or U5026 (N_5026,N_4605,N_4521);
nand U5027 (N_5027,N_4636,N_4498);
or U5028 (N_5028,N_4232,N_4575);
or U5029 (N_5029,N_4290,N_4453);
and U5030 (N_5030,N_4293,N_4230);
nor U5031 (N_5031,N_4288,N_4682);
nand U5032 (N_5032,N_4256,N_4417);
nor U5033 (N_5033,N_4535,N_4402);
or U5034 (N_5034,N_4797,N_4323);
or U5035 (N_5035,N_4464,N_4413);
nor U5036 (N_5036,N_4492,N_4562);
nand U5037 (N_5037,N_4460,N_4785);
and U5038 (N_5038,N_4518,N_4299);
and U5039 (N_5039,N_4378,N_4696);
or U5040 (N_5040,N_4524,N_4490);
and U5041 (N_5041,N_4620,N_4386);
nor U5042 (N_5042,N_4700,N_4225);
or U5043 (N_5043,N_4318,N_4718);
or U5044 (N_5044,N_4529,N_4376);
and U5045 (N_5045,N_4202,N_4522);
nor U5046 (N_5046,N_4242,N_4550);
or U5047 (N_5047,N_4710,N_4270);
and U5048 (N_5048,N_4536,N_4221);
nand U5049 (N_5049,N_4381,N_4292);
nand U5050 (N_5050,N_4285,N_4701);
xor U5051 (N_5051,N_4623,N_4542);
and U5052 (N_5052,N_4469,N_4480);
nor U5053 (N_5053,N_4735,N_4649);
nand U5054 (N_5054,N_4686,N_4543);
and U5055 (N_5055,N_4667,N_4588);
or U5056 (N_5056,N_4653,N_4408);
or U5057 (N_5057,N_4321,N_4739);
and U5058 (N_5058,N_4659,N_4329);
nand U5059 (N_5059,N_4317,N_4345);
nor U5060 (N_5060,N_4303,N_4383);
and U5061 (N_5061,N_4205,N_4745);
nor U5062 (N_5062,N_4382,N_4798);
nor U5063 (N_5063,N_4749,N_4627);
and U5064 (N_5064,N_4697,N_4681);
or U5065 (N_5065,N_4366,N_4654);
nor U5066 (N_5066,N_4226,N_4665);
and U5067 (N_5067,N_4658,N_4702);
and U5068 (N_5068,N_4361,N_4638);
nand U5069 (N_5069,N_4639,N_4600);
nand U5070 (N_5070,N_4756,N_4335);
nor U5071 (N_5071,N_4677,N_4582);
or U5072 (N_5072,N_4771,N_4247);
nand U5073 (N_5073,N_4725,N_4437);
nor U5074 (N_5074,N_4655,N_4406);
nor U5075 (N_5075,N_4737,N_4416);
nor U5076 (N_5076,N_4695,N_4269);
or U5077 (N_5077,N_4420,N_4572);
or U5078 (N_5078,N_4447,N_4200);
and U5079 (N_5079,N_4611,N_4790);
nor U5080 (N_5080,N_4693,N_4233);
or U5081 (N_5081,N_4496,N_4523);
and U5082 (N_5082,N_4252,N_4435);
nor U5083 (N_5083,N_4486,N_4648);
or U5084 (N_5084,N_4768,N_4429);
nor U5085 (N_5085,N_4530,N_4752);
nand U5086 (N_5086,N_4347,N_4621);
nand U5087 (N_5087,N_4504,N_4263);
nand U5088 (N_5088,N_4380,N_4487);
and U5089 (N_5089,N_4354,N_4561);
and U5090 (N_5090,N_4213,N_4577);
or U5091 (N_5091,N_4717,N_4645);
nand U5092 (N_5092,N_4531,N_4617);
nor U5093 (N_5093,N_4672,N_4391);
or U5094 (N_5094,N_4565,N_4767);
and U5095 (N_5095,N_4373,N_4541);
nor U5096 (N_5096,N_4352,N_4360);
nand U5097 (N_5097,N_4421,N_4662);
nor U5098 (N_5098,N_4776,N_4457);
or U5099 (N_5099,N_4593,N_4584);
and U5100 (N_5100,N_4417,N_4462);
and U5101 (N_5101,N_4648,N_4389);
and U5102 (N_5102,N_4365,N_4653);
or U5103 (N_5103,N_4546,N_4562);
or U5104 (N_5104,N_4584,N_4766);
nor U5105 (N_5105,N_4548,N_4741);
nor U5106 (N_5106,N_4378,N_4353);
xnor U5107 (N_5107,N_4295,N_4548);
nand U5108 (N_5108,N_4429,N_4612);
nor U5109 (N_5109,N_4713,N_4753);
nand U5110 (N_5110,N_4596,N_4298);
nand U5111 (N_5111,N_4734,N_4396);
or U5112 (N_5112,N_4760,N_4379);
and U5113 (N_5113,N_4243,N_4315);
or U5114 (N_5114,N_4505,N_4231);
or U5115 (N_5115,N_4281,N_4477);
or U5116 (N_5116,N_4444,N_4333);
nor U5117 (N_5117,N_4743,N_4241);
nand U5118 (N_5118,N_4757,N_4469);
and U5119 (N_5119,N_4311,N_4572);
nor U5120 (N_5120,N_4560,N_4201);
or U5121 (N_5121,N_4491,N_4773);
or U5122 (N_5122,N_4572,N_4283);
xor U5123 (N_5123,N_4429,N_4322);
nor U5124 (N_5124,N_4603,N_4292);
or U5125 (N_5125,N_4217,N_4279);
nand U5126 (N_5126,N_4649,N_4357);
and U5127 (N_5127,N_4405,N_4278);
xor U5128 (N_5128,N_4430,N_4541);
nor U5129 (N_5129,N_4406,N_4390);
or U5130 (N_5130,N_4429,N_4532);
nor U5131 (N_5131,N_4230,N_4534);
and U5132 (N_5132,N_4447,N_4280);
nand U5133 (N_5133,N_4528,N_4429);
or U5134 (N_5134,N_4499,N_4235);
and U5135 (N_5135,N_4245,N_4548);
nor U5136 (N_5136,N_4676,N_4383);
nor U5137 (N_5137,N_4696,N_4307);
or U5138 (N_5138,N_4500,N_4350);
xor U5139 (N_5139,N_4763,N_4359);
nand U5140 (N_5140,N_4397,N_4520);
nor U5141 (N_5141,N_4517,N_4632);
nor U5142 (N_5142,N_4308,N_4226);
nand U5143 (N_5143,N_4346,N_4362);
nand U5144 (N_5144,N_4569,N_4334);
nor U5145 (N_5145,N_4376,N_4325);
nand U5146 (N_5146,N_4723,N_4271);
nand U5147 (N_5147,N_4206,N_4205);
or U5148 (N_5148,N_4687,N_4741);
nor U5149 (N_5149,N_4388,N_4596);
or U5150 (N_5150,N_4356,N_4627);
nand U5151 (N_5151,N_4688,N_4474);
nor U5152 (N_5152,N_4691,N_4505);
or U5153 (N_5153,N_4426,N_4484);
and U5154 (N_5154,N_4419,N_4329);
or U5155 (N_5155,N_4745,N_4357);
nor U5156 (N_5156,N_4518,N_4615);
nor U5157 (N_5157,N_4604,N_4349);
or U5158 (N_5158,N_4334,N_4286);
or U5159 (N_5159,N_4464,N_4624);
nor U5160 (N_5160,N_4483,N_4738);
nand U5161 (N_5161,N_4747,N_4640);
nor U5162 (N_5162,N_4293,N_4718);
and U5163 (N_5163,N_4452,N_4297);
and U5164 (N_5164,N_4698,N_4353);
and U5165 (N_5165,N_4429,N_4468);
nand U5166 (N_5166,N_4634,N_4462);
nand U5167 (N_5167,N_4371,N_4484);
nor U5168 (N_5168,N_4549,N_4441);
or U5169 (N_5169,N_4686,N_4584);
nand U5170 (N_5170,N_4438,N_4431);
xor U5171 (N_5171,N_4406,N_4374);
and U5172 (N_5172,N_4518,N_4430);
or U5173 (N_5173,N_4643,N_4488);
or U5174 (N_5174,N_4653,N_4236);
nand U5175 (N_5175,N_4569,N_4749);
nand U5176 (N_5176,N_4404,N_4712);
nand U5177 (N_5177,N_4369,N_4430);
nor U5178 (N_5178,N_4338,N_4436);
or U5179 (N_5179,N_4323,N_4556);
nor U5180 (N_5180,N_4388,N_4707);
and U5181 (N_5181,N_4377,N_4624);
or U5182 (N_5182,N_4590,N_4760);
and U5183 (N_5183,N_4273,N_4360);
and U5184 (N_5184,N_4309,N_4232);
nor U5185 (N_5185,N_4213,N_4431);
nor U5186 (N_5186,N_4600,N_4251);
nand U5187 (N_5187,N_4543,N_4548);
nor U5188 (N_5188,N_4349,N_4295);
xor U5189 (N_5189,N_4367,N_4228);
or U5190 (N_5190,N_4250,N_4318);
nand U5191 (N_5191,N_4551,N_4379);
and U5192 (N_5192,N_4675,N_4382);
nor U5193 (N_5193,N_4466,N_4430);
nor U5194 (N_5194,N_4508,N_4635);
or U5195 (N_5195,N_4389,N_4548);
or U5196 (N_5196,N_4425,N_4353);
nand U5197 (N_5197,N_4592,N_4239);
or U5198 (N_5198,N_4226,N_4384);
nand U5199 (N_5199,N_4399,N_4349);
nand U5200 (N_5200,N_4568,N_4274);
and U5201 (N_5201,N_4548,N_4667);
and U5202 (N_5202,N_4729,N_4307);
nand U5203 (N_5203,N_4448,N_4585);
and U5204 (N_5204,N_4473,N_4304);
and U5205 (N_5205,N_4604,N_4251);
nand U5206 (N_5206,N_4513,N_4289);
and U5207 (N_5207,N_4406,N_4278);
and U5208 (N_5208,N_4606,N_4493);
nor U5209 (N_5209,N_4552,N_4429);
or U5210 (N_5210,N_4385,N_4383);
nor U5211 (N_5211,N_4429,N_4562);
and U5212 (N_5212,N_4303,N_4298);
nand U5213 (N_5213,N_4330,N_4660);
xor U5214 (N_5214,N_4623,N_4265);
or U5215 (N_5215,N_4757,N_4781);
and U5216 (N_5216,N_4657,N_4374);
nor U5217 (N_5217,N_4473,N_4412);
nor U5218 (N_5218,N_4454,N_4551);
nand U5219 (N_5219,N_4635,N_4700);
xnor U5220 (N_5220,N_4521,N_4281);
or U5221 (N_5221,N_4276,N_4222);
or U5222 (N_5222,N_4435,N_4230);
nand U5223 (N_5223,N_4680,N_4645);
nor U5224 (N_5224,N_4354,N_4636);
nand U5225 (N_5225,N_4697,N_4223);
nand U5226 (N_5226,N_4385,N_4791);
nor U5227 (N_5227,N_4629,N_4606);
and U5228 (N_5228,N_4435,N_4740);
or U5229 (N_5229,N_4794,N_4399);
nor U5230 (N_5230,N_4281,N_4577);
nand U5231 (N_5231,N_4620,N_4402);
nand U5232 (N_5232,N_4647,N_4624);
nor U5233 (N_5233,N_4588,N_4628);
and U5234 (N_5234,N_4507,N_4230);
or U5235 (N_5235,N_4505,N_4656);
and U5236 (N_5236,N_4673,N_4634);
or U5237 (N_5237,N_4581,N_4586);
or U5238 (N_5238,N_4712,N_4435);
nor U5239 (N_5239,N_4647,N_4388);
and U5240 (N_5240,N_4281,N_4479);
nor U5241 (N_5241,N_4210,N_4507);
nor U5242 (N_5242,N_4226,N_4792);
and U5243 (N_5243,N_4207,N_4222);
and U5244 (N_5244,N_4716,N_4665);
nand U5245 (N_5245,N_4307,N_4497);
nand U5246 (N_5246,N_4386,N_4303);
or U5247 (N_5247,N_4389,N_4561);
and U5248 (N_5248,N_4775,N_4721);
or U5249 (N_5249,N_4249,N_4384);
or U5250 (N_5250,N_4763,N_4634);
nor U5251 (N_5251,N_4323,N_4699);
or U5252 (N_5252,N_4243,N_4695);
nor U5253 (N_5253,N_4300,N_4739);
or U5254 (N_5254,N_4754,N_4376);
nor U5255 (N_5255,N_4321,N_4645);
nor U5256 (N_5256,N_4450,N_4288);
nand U5257 (N_5257,N_4492,N_4236);
and U5258 (N_5258,N_4209,N_4374);
xor U5259 (N_5259,N_4408,N_4318);
and U5260 (N_5260,N_4291,N_4287);
nand U5261 (N_5261,N_4629,N_4344);
or U5262 (N_5262,N_4729,N_4613);
nand U5263 (N_5263,N_4363,N_4768);
and U5264 (N_5264,N_4495,N_4363);
and U5265 (N_5265,N_4310,N_4231);
and U5266 (N_5266,N_4692,N_4675);
and U5267 (N_5267,N_4226,N_4687);
or U5268 (N_5268,N_4428,N_4640);
nand U5269 (N_5269,N_4695,N_4484);
and U5270 (N_5270,N_4213,N_4525);
or U5271 (N_5271,N_4774,N_4234);
and U5272 (N_5272,N_4616,N_4798);
nand U5273 (N_5273,N_4648,N_4371);
nor U5274 (N_5274,N_4514,N_4767);
and U5275 (N_5275,N_4720,N_4201);
or U5276 (N_5276,N_4597,N_4484);
or U5277 (N_5277,N_4499,N_4202);
or U5278 (N_5278,N_4717,N_4348);
nor U5279 (N_5279,N_4668,N_4247);
nor U5280 (N_5280,N_4261,N_4421);
nand U5281 (N_5281,N_4468,N_4641);
nor U5282 (N_5282,N_4343,N_4200);
nand U5283 (N_5283,N_4422,N_4374);
nor U5284 (N_5284,N_4419,N_4368);
nand U5285 (N_5285,N_4727,N_4686);
nor U5286 (N_5286,N_4469,N_4587);
nor U5287 (N_5287,N_4752,N_4469);
nand U5288 (N_5288,N_4418,N_4485);
nor U5289 (N_5289,N_4245,N_4459);
nor U5290 (N_5290,N_4752,N_4683);
and U5291 (N_5291,N_4767,N_4770);
xor U5292 (N_5292,N_4308,N_4657);
or U5293 (N_5293,N_4630,N_4217);
or U5294 (N_5294,N_4362,N_4245);
or U5295 (N_5295,N_4522,N_4316);
and U5296 (N_5296,N_4606,N_4377);
xor U5297 (N_5297,N_4379,N_4292);
or U5298 (N_5298,N_4217,N_4738);
and U5299 (N_5299,N_4619,N_4224);
and U5300 (N_5300,N_4745,N_4635);
xnor U5301 (N_5301,N_4599,N_4771);
nor U5302 (N_5302,N_4522,N_4490);
and U5303 (N_5303,N_4422,N_4435);
and U5304 (N_5304,N_4248,N_4362);
nor U5305 (N_5305,N_4618,N_4426);
and U5306 (N_5306,N_4735,N_4276);
xnor U5307 (N_5307,N_4513,N_4536);
nand U5308 (N_5308,N_4497,N_4701);
nor U5309 (N_5309,N_4572,N_4711);
and U5310 (N_5310,N_4306,N_4598);
nor U5311 (N_5311,N_4699,N_4264);
and U5312 (N_5312,N_4737,N_4376);
xnor U5313 (N_5313,N_4375,N_4230);
nor U5314 (N_5314,N_4247,N_4334);
or U5315 (N_5315,N_4649,N_4724);
nand U5316 (N_5316,N_4673,N_4358);
nand U5317 (N_5317,N_4465,N_4721);
nor U5318 (N_5318,N_4797,N_4625);
or U5319 (N_5319,N_4478,N_4234);
nand U5320 (N_5320,N_4344,N_4265);
and U5321 (N_5321,N_4399,N_4751);
or U5322 (N_5322,N_4537,N_4320);
or U5323 (N_5323,N_4779,N_4777);
nor U5324 (N_5324,N_4681,N_4400);
nor U5325 (N_5325,N_4533,N_4417);
or U5326 (N_5326,N_4635,N_4676);
and U5327 (N_5327,N_4702,N_4606);
and U5328 (N_5328,N_4580,N_4385);
nor U5329 (N_5329,N_4281,N_4742);
nand U5330 (N_5330,N_4693,N_4527);
and U5331 (N_5331,N_4310,N_4396);
or U5332 (N_5332,N_4695,N_4687);
xor U5333 (N_5333,N_4729,N_4620);
nand U5334 (N_5334,N_4504,N_4257);
and U5335 (N_5335,N_4616,N_4302);
and U5336 (N_5336,N_4448,N_4618);
or U5337 (N_5337,N_4677,N_4200);
nand U5338 (N_5338,N_4519,N_4441);
xnor U5339 (N_5339,N_4311,N_4766);
nor U5340 (N_5340,N_4779,N_4278);
nand U5341 (N_5341,N_4429,N_4218);
nor U5342 (N_5342,N_4759,N_4263);
or U5343 (N_5343,N_4581,N_4332);
nor U5344 (N_5344,N_4740,N_4476);
or U5345 (N_5345,N_4253,N_4625);
and U5346 (N_5346,N_4256,N_4562);
nand U5347 (N_5347,N_4471,N_4525);
nand U5348 (N_5348,N_4585,N_4674);
xnor U5349 (N_5349,N_4470,N_4776);
xor U5350 (N_5350,N_4799,N_4467);
nor U5351 (N_5351,N_4684,N_4289);
nor U5352 (N_5352,N_4755,N_4308);
nand U5353 (N_5353,N_4248,N_4431);
and U5354 (N_5354,N_4498,N_4778);
nand U5355 (N_5355,N_4489,N_4693);
nand U5356 (N_5356,N_4549,N_4426);
and U5357 (N_5357,N_4555,N_4417);
nand U5358 (N_5358,N_4255,N_4261);
nor U5359 (N_5359,N_4619,N_4574);
and U5360 (N_5360,N_4237,N_4532);
or U5361 (N_5361,N_4762,N_4635);
and U5362 (N_5362,N_4691,N_4381);
and U5363 (N_5363,N_4562,N_4761);
nor U5364 (N_5364,N_4586,N_4388);
xnor U5365 (N_5365,N_4230,N_4235);
or U5366 (N_5366,N_4492,N_4209);
or U5367 (N_5367,N_4468,N_4558);
nor U5368 (N_5368,N_4487,N_4595);
or U5369 (N_5369,N_4311,N_4684);
xnor U5370 (N_5370,N_4540,N_4478);
nand U5371 (N_5371,N_4424,N_4782);
nand U5372 (N_5372,N_4731,N_4265);
and U5373 (N_5373,N_4752,N_4277);
and U5374 (N_5374,N_4671,N_4245);
or U5375 (N_5375,N_4310,N_4463);
or U5376 (N_5376,N_4659,N_4569);
nand U5377 (N_5377,N_4320,N_4761);
and U5378 (N_5378,N_4438,N_4738);
nand U5379 (N_5379,N_4295,N_4688);
nand U5380 (N_5380,N_4248,N_4417);
nor U5381 (N_5381,N_4709,N_4691);
or U5382 (N_5382,N_4504,N_4675);
nor U5383 (N_5383,N_4429,N_4207);
or U5384 (N_5384,N_4404,N_4425);
nand U5385 (N_5385,N_4361,N_4202);
nand U5386 (N_5386,N_4285,N_4498);
or U5387 (N_5387,N_4510,N_4280);
nand U5388 (N_5388,N_4320,N_4324);
and U5389 (N_5389,N_4526,N_4384);
and U5390 (N_5390,N_4475,N_4283);
nor U5391 (N_5391,N_4387,N_4358);
nand U5392 (N_5392,N_4493,N_4559);
or U5393 (N_5393,N_4527,N_4524);
nor U5394 (N_5394,N_4769,N_4667);
nor U5395 (N_5395,N_4420,N_4577);
nor U5396 (N_5396,N_4739,N_4371);
or U5397 (N_5397,N_4488,N_4660);
or U5398 (N_5398,N_4384,N_4777);
and U5399 (N_5399,N_4243,N_4616);
and U5400 (N_5400,N_5062,N_5027);
or U5401 (N_5401,N_5327,N_4998);
nor U5402 (N_5402,N_4840,N_5377);
and U5403 (N_5403,N_5365,N_5375);
xnor U5404 (N_5404,N_5104,N_5015);
and U5405 (N_5405,N_4860,N_5356);
nor U5406 (N_5406,N_4847,N_4886);
nand U5407 (N_5407,N_4825,N_5235);
nor U5408 (N_5408,N_5001,N_5218);
and U5409 (N_5409,N_5086,N_5190);
nor U5410 (N_5410,N_5009,N_5342);
nor U5411 (N_5411,N_5227,N_4979);
nor U5412 (N_5412,N_5204,N_4974);
nor U5413 (N_5413,N_5025,N_4902);
or U5414 (N_5414,N_5233,N_5150);
or U5415 (N_5415,N_5386,N_5095);
or U5416 (N_5416,N_4896,N_5284);
and U5417 (N_5417,N_5128,N_5296);
or U5418 (N_5418,N_4955,N_5048);
and U5419 (N_5419,N_5311,N_5213);
nor U5420 (N_5420,N_5011,N_4967);
and U5421 (N_5421,N_5304,N_4940);
and U5422 (N_5422,N_4897,N_5347);
and U5423 (N_5423,N_5023,N_4879);
and U5424 (N_5424,N_5170,N_5394);
nor U5425 (N_5425,N_4822,N_4813);
nor U5426 (N_5426,N_5329,N_4993);
nor U5427 (N_5427,N_5334,N_5200);
and U5428 (N_5428,N_5199,N_4853);
and U5429 (N_5429,N_4842,N_5266);
nand U5430 (N_5430,N_5156,N_4984);
or U5431 (N_5431,N_5254,N_5191);
and U5432 (N_5432,N_4829,N_4841);
and U5433 (N_5433,N_5181,N_5106);
nor U5434 (N_5434,N_4924,N_5357);
and U5435 (N_5435,N_5203,N_5073);
nor U5436 (N_5436,N_5164,N_4827);
and U5437 (N_5437,N_5026,N_5019);
nand U5438 (N_5438,N_5237,N_4923);
and U5439 (N_5439,N_5238,N_4812);
and U5440 (N_5440,N_5344,N_5306);
xnor U5441 (N_5441,N_5182,N_5189);
nor U5442 (N_5442,N_5331,N_4921);
and U5443 (N_5443,N_5391,N_5163);
and U5444 (N_5444,N_4958,N_5042);
nand U5445 (N_5445,N_4850,N_5349);
nor U5446 (N_5446,N_5064,N_5038);
or U5447 (N_5447,N_5148,N_5206);
and U5448 (N_5448,N_5116,N_5393);
nor U5449 (N_5449,N_4999,N_5360);
or U5450 (N_5450,N_5217,N_5096);
nor U5451 (N_5451,N_5288,N_5007);
xor U5452 (N_5452,N_5010,N_5390);
or U5453 (N_5453,N_5176,N_5255);
and U5454 (N_5454,N_5399,N_5320);
and U5455 (N_5455,N_5083,N_5300);
nor U5456 (N_5456,N_5022,N_5376);
or U5457 (N_5457,N_4845,N_5052);
nand U5458 (N_5458,N_4875,N_5325);
or U5459 (N_5459,N_4884,N_4820);
or U5460 (N_5460,N_5302,N_4932);
nand U5461 (N_5461,N_5228,N_5321);
or U5462 (N_5462,N_4959,N_5184);
nor U5463 (N_5463,N_5216,N_5058);
or U5464 (N_5464,N_5317,N_4803);
nor U5465 (N_5465,N_5014,N_5242);
or U5466 (N_5466,N_4887,N_5326);
nor U5467 (N_5467,N_5281,N_5241);
nor U5468 (N_5468,N_5250,N_5142);
nor U5469 (N_5469,N_5274,N_5054);
nand U5470 (N_5470,N_5291,N_5348);
and U5471 (N_5471,N_5352,N_5308);
nand U5472 (N_5472,N_4913,N_4851);
nor U5473 (N_5473,N_5107,N_5060);
nor U5474 (N_5474,N_5397,N_5032);
nor U5475 (N_5475,N_4944,N_4818);
or U5476 (N_5476,N_4995,N_4945);
or U5477 (N_5477,N_5364,N_5382);
and U5478 (N_5478,N_5120,N_4912);
xnor U5479 (N_5479,N_5367,N_5127);
or U5480 (N_5480,N_4872,N_5279);
nand U5481 (N_5481,N_5290,N_5339);
nand U5482 (N_5482,N_5336,N_5172);
nor U5483 (N_5483,N_5369,N_4889);
nor U5484 (N_5484,N_4929,N_4927);
or U5485 (N_5485,N_5387,N_5310);
xor U5486 (N_5486,N_4905,N_4870);
xor U5487 (N_5487,N_4997,N_4833);
or U5488 (N_5488,N_5253,N_5040);
and U5489 (N_5489,N_5309,N_4966);
nor U5490 (N_5490,N_4868,N_4961);
or U5491 (N_5491,N_4809,N_4920);
nor U5492 (N_5492,N_5074,N_4973);
and U5493 (N_5493,N_5185,N_5381);
and U5494 (N_5494,N_4881,N_4843);
nor U5495 (N_5495,N_5335,N_5175);
nor U5496 (N_5496,N_5282,N_5353);
or U5497 (N_5497,N_5202,N_5395);
nand U5498 (N_5498,N_4819,N_5097);
nand U5499 (N_5499,N_5051,N_4989);
or U5500 (N_5500,N_5146,N_5151);
and U5501 (N_5501,N_4919,N_5117);
nor U5502 (N_5502,N_5141,N_5268);
or U5503 (N_5503,N_4888,N_5065);
or U5504 (N_5504,N_5355,N_5041);
nor U5505 (N_5505,N_4900,N_5211);
nor U5506 (N_5506,N_5078,N_5122);
nor U5507 (N_5507,N_4970,N_5134);
and U5508 (N_5508,N_5214,N_5215);
and U5509 (N_5509,N_4891,N_5366);
or U5510 (N_5510,N_4909,N_5244);
or U5511 (N_5511,N_5071,N_5257);
nand U5512 (N_5512,N_4988,N_4865);
nor U5513 (N_5513,N_5084,N_5021);
nand U5514 (N_5514,N_4895,N_4869);
nand U5515 (N_5515,N_4941,N_5076);
nand U5516 (N_5516,N_4992,N_4807);
nor U5517 (N_5517,N_4908,N_4834);
nand U5518 (N_5518,N_4986,N_4878);
or U5519 (N_5519,N_5131,N_4949);
nand U5520 (N_5520,N_5144,N_4934);
or U5521 (N_5521,N_4882,N_5225);
and U5522 (N_5522,N_4983,N_4951);
and U5523 (N_5523,N_5186,N_5138);
and U5524 (N_5524,N_4950,N_5256);
and U5525 (N_5525,N_4873,N_5043);
and U5526 (N_5526,N_5082,N_5036);
nand U5527 (N_5527,N_4880,N_5292);
and U5528 (N_5528,N_5105,N_5035);
and U5529 (N_5529,N_4823,N_5016);
and U5530 (N_5530,N_5318,N_5059);
xor U5531 (N_5531,N_5396,N_4866);
or U5532 (N_5532,N_5037,N_5363);
and U5533 (N_5533,N_5119,N_5247);
or U5534 (N_5534,N_5069,N_5187);
nand U5535 (N_5535,N_5207,N_4801);
nor U5536 (N_5536,N_5209,N_5328);
and U5537 (N_5537,N_5314,N_5162);
and U5538 (N_5538,N_4901,N_5240);
nand U5539 (N_5539,N_5384,N_5029);
and U5540 (N_5540,N_5262,N_5020);
nor U5541 (N_5541,N_4964,N_5323);
and U5542 (N_5542,N_5273,N_4991);
and U5543 (N_5543,N_5285,N_5103);
nand U5544 (N_5544,N_5208,N_5003);
nor U5545 (N_5545,N_5220,N_5350);
and U5546 (N_5546,N_4933,N_4987);
nand U5547 (N_5547,N_4971,N_4938);
nor U5548 (N_5548,N_5383,N_4925);
and U5549 (N_5549,N_5109,N_5155);
or U5550 (N_5550,N_4968,N_5180);
nor U5551 (N_5551,N_4990,N_5088);
nor U5552 (N_5552,N_5392,N_4864);
and U5553 (N_5553,N_4969,N_5046);
or U5554 (N_5554,N_5210,N_5110);
nand U5555 (N_5555,N_4874,N_5201);
nor U5556 (N_5556,N_5275,N_4982);
nor U5557 (N_5557,N_4857,N_5243);
or U5558 (N_5558,N_5072,N_4837);
or U5559 (N_5559,N_5371,N_5287);
and U5560 (N_5560,N_5188,N_5299);
or U5561 (N_5561,N_4815,N_5159);
nor U5562 (N_5562,N_4838,N_5121);
xnor U5563 (N_5563,N_4848,N_5280);
and U5564 (N_5564,N_5388,N_5231);
nand U5565 (N_5565,N_5263,N_5087);
nor U5566 (N_5566,N_5113,N_4885);
xnor U5567 (N_5567,N_4942,N_5112);
nor U5568 (N_5568,N_4814,N_4839);
and U5569 (N_5569,N_5005,N_5012);
and U5570 (N_5570,N_5099,N_5283);
nor U5571 (N_5571,N_5293,N_4802);
or U5572 (N_5572,N_5070,N_4894);
nor U5573 (N_5573,N_5123,N_5219);
nor U5574 (N_5574,N_5313,N_5006);
nand U5575 (N_5575,N_5153,N_4917);
nand U5576 (N_5576,N_5398,N_5135);
nand U5577 (N_5577,N_5261,N_5091);
nand U5578 (N_5578,N_4935,N_5179);
and U5579 (N_5579,N_5248,N_5340);
and U5580 (N_5580,N_5270,N_5232);
and U5581 (N_5581,N_5130,N_4861);
nand U5582 (N_5582,N_5034,N_5315);
nor U5583 (N_5583,N_4899,N_5165);
nand U5584 (N_5584,N_4844,N_5298);
nor U5585 (N_5585,N_5358,N_5081);
or U5586 (N_5586,N_5249,N_5139);
and U5587 (N_5587,N_5177,N_4846);
and U5588 (N_5588,N_4832,N_4922);
or U5589 (N_5589,N_4821,N_5264);
nand U5590 (N_5590,N_5137,N_4811);
or U5591 (N_5591,N_5251,N_4858);
nand U5592 (N_5592,N_5000,N_5033);
nor U5593 (N_5593,N_5324,N_5024);
nand U5594 (N_5594,N_5140,N_5212);
nand U5595 (N_5595,N_5111,N_5197);
and U5596 (N_5596,N_5147,N_5183);
nor U5597 (N_5597,N_5239,N_5226);
or U5598 (N_5598,N_5126,N_4963);
and U5599 (N_5599,N_5359,N_4862);
nand U5600 (N_5600,N_4810,N_4867);
and U5601 (N_5601,N_5169,N_5312);
or U5602 (N_5602,N_4911,N_5267);
or U5603 (N_5603,N_4856,N_5008);
or U5604 (N_5604,N_5013,N_5192);
or U5605 (N_5605,N_5161,N_4852);
nand U5606 (N_5606,N_4863,N_5278);
nand U5607 (N_5607,N_4904,N_5337);
nor U5608 (N_5608,N_4859,N_5223);
or U5609 (N_5609,N_5018,N_5098);
nor U5610 (N_5610,N_5193,N_4871);
nor U5611 (N_5611,N_4806,N_4828);
or U5612 (N_5612,N_5380,N_5289);
nand U5613 (N_5613,N_4883,N_5085);
and U5614 (N_5614,N_5379,N_5224);
nor U5615 (N_5615,N_5271,N_5090);
nor U5616 (N_5616,N_5368,N_5143);
and U5617 (N_5617,N_4928,N_5236);
and U5618 (N_5618,N_5166,N_5333);
or U5619 (N_5619,N_4965,N_4947);
nand U5620 (N_5620,N_4826,N_5294);
nand U5621 (N_5621,N_5272,N_5067);
or U5622 (N_5622,N_5258,N_4980);
nand U5623 (N_5623,N_5171,N_5322);
nand U5624 (N_5624,N_5246,N_5075);
nor U5625 (N_5625,N_4910,N_5080);
nand U5626 (N_5626,N_5125,N_4835);
or U5627 (N_5627,N_5370,N_5361);
nor U5628 (N_5628,N_5049,N_4824);
and U5629 (N_5629,N_5265,N_4985);
nor U5630 (N_5630,N_4915,N_5174);
or U5631 (N_5631,N_5030,N_5297);
nor U5632 (N_5632,N_4918,N_5385);
and U5633 (N_5633,N_4943,N_5222);
nand U5634 (N_5634,N_5221,N_4893);
or U5635 (N_5635,N_4890,N_5145);
nand U5636 (N_5636,N_5295,N_4855);
and U5637 (N_5637,N_4831,N_4960);
or U5638 (N_5638,N_5044,N_5028);
nand U5639 (N_5639,N_5152,N_5305);
and U5640 (N_5640,N_5031,N_5346);
nand U5641 (N_5641,N_5286,N_4916);
and U5642 (N_5642,N_5343,N_5167);
nand U5643 (N_5643,N_5102,N_5341);
nor U5644 (N_5644,N_5089,N_5269);
and U5645 (N_5645,N_4817,N_5124);
nand U5646 (N_5646,N_5056,N_5157);
nand U5647 (N_5647,N_5351,N_4805);
nand U5648 (N_5648,N_4906,N_4953);
nand U5649 (N_5649,N_5061,N_5063);
and U5650 (N_5650,N_5002,N_5354);
nand U5651 (N_5651,N_5158,N_5093);
or U5652 (N_5652,N_5205,N_4962);
or U5653 (N_5653,N_4876,N_4804);
or U5654 (N_5654,N_4898,N_5316);
and U5655 (N_5655,N_5050,N_4954);
nand U5656 (N_5656,N_5389,N_5259);
nor U5657 (N_5657,N_4914,N_4849);
or U5658 (N_5658,N_5362,N_4836);
and U5659 (N_5659,N_4903,N_5168);
and U5660 (N_5660,N_5234,N_4956);
and U5661 (N_5661,N_5319,N_4981);
or U5662 (N_5662,N_5332,N_5195);
nor U5663 (N_5663,N_4957,N_5154);
nor U5664 (N_5664,N_5115,N_5330);
xnor U5665 (N_5665,N_5303,N_4816);
nor U5666 (N_5666,N_5194,N_5307);
nand U5667 (N_5667,N_4948,N_5230);
and U5668 (N_5668,N_4930,N_5057);
or U5669 (N_5669,N_5132,N_4830);
xnor U5670 (N_5670,N_5100,N_4977);
or U5671 (N_5671,N_5066,N_4808);
nor U5672 (N_5672,N_5277,N_4877);
nor U5673 (N_5673,N_4972,N_5045);
nand U5674 (N_5674,N_5077,N_4937);
nand U5675 (N_5675,N_5149,N_5047);
and U5676 (N_5676,N_5374,N_4931);
or U5677 (N_5677,N_5068,N_4907);
and U5678 (N_5678,N_5101,N_4996);
and U5679 (N_5679,N_4975,N_5133);
nand U5680 (N_5680,N_5178,N_4994);
nor U5681 (N_5681,N_5094,N_5372);
nand U5682 (N_5682,N_5055,N_5092);
nor U5683 (N_5683,N_4854,N_5173);
nand U5684 (N_5684,N_4946,N_4939);
nor U5685 (N_5685,N_5229,N_5245);
or U5686 (N_5686,N_4976,N_5198);
nor U5687 (N_5687,N_5017,N_4936);
nand U5688 (N_5688,N_5039,N_5053);
nand U5689 (N_5689,N_5129,N_5252);
or U5690 (N_5690,N_4800,N_5260);
and U5691 (N_5691,N_5276,N_5196);
and U5692 (N_5692,N_5301,N_5108);
nor U5693 (N_5693,N_5118,N_5079);
nor U5694 (N_5694,N_5373,N_4926);
nor U5695 (N_5695,N_4952,N_4978);
nor U5696 (N_5696,N_5378,N_5114);
and U5697 (N_5697,N_5338,N_5345);
and U5698 (N_5698,N_5004,N_4892);
and U5699 (N_5699,N_5136,N_5160);
or U5700 (N_5700,N_4827,N_5169);
nand U5701 (N_5701,N_4924,N_5285);
nand U5702 (N_5702,N_5168,N_5107);
nor U5703 (N_5703,N_5002,N_5201);
nor U5704 (N_5704,N_5073,N_4940);
nand U5705 (N_5705,N_5099,N_5211);
or U5706 (N_5706,N_5089,N_5004);
or U5707 (N_5707,N_5230,N_5167);
or U5708 (N_5708,N_5013,N_5030);
and U5709 (N_5709,N_4956,N_4847);
and U5710 (N_5710,N_5152,N_5272);
and U5711 (N_5711,N_4902,N_4832);
or U5712 (N_5712,N_5088,N_5037);
and U5713 (N_5713,N_5053,N_5226);
and U5714 (N_5714,N_5348,N_4834);
or U5715 (N_5715,N_5084,N_5085);
nor U5716 (N_5716,N_5228,N_5060);
and U5717 (N_5717,N_4924,N_4847);
or U5718 (N_5718,N_4862,N_4961);
nor U5719 (N_5719,N_5231,N_5377);
xnor U5720 (N_5720,N_5258,N_4818);
xnor U5721 (N_5721,N_4863,N_5319);
nor U5722 (N_5722,N_5320,N_5397);
nand U5723 (N_5723,N_5319,N_4874);
nand U5724 (N_5724,N_5153,N_5237);
nand U5725 (N_5725,N_5144,N_5262);
nor U5726 (N_5726,N_5213,N_5319);
nand U5727 (N_5727,N_5315,N_5278);
or U5728 (N_5728,N_5093,N_5310);
nand U5729 (N_5729,N_4931,N_4921);
and U5730 (N_5730,N_4815,N_5300);
nand U5731 (N_5731,N_4891,N_4929);
and U5732 (N_5732,N_5086,N_4879);
nor U5733 (N_5733,N_4822,N_5124);
nor U5734 (N_5734,N_5065,N_4993);
nor U5735 (N_5735,N_5372,N_5187);
and U5736 (N_5736,N_5069,N_5272);
nor U5737 (N_5737,N_5322,N_5103);
and U5738 (N_5738,N_5246,N_5361);
and U5739 (N_5739,N_5324,N_4813);
and U5740 (N_5740,N_5098,N_4916);
or U5741 (N_5741,N_5314,N_4871);
or U5742 (N_5742,N_5043,N_5133);
nand U5743 (N_5743,N_5289,N_4972);
nand U5744 (N_5744,N_5135,N_5187);
or U5745 (N_5745,N_5339,N_5115);
nand U5746 (N_5746,N_4907,N_5049);
nand U5747 (N_5747,N_5104,N_5124);
and U5748 (N_5748,N_5217,N_4803);
and U5749 (N_5749,N_4963,N_5353);
or U5750 (N_5750,N_4838,N_4995);
and U5751 (N_5751,N_5165,N_4872);
nor U5752 (N_5752,N_4934,N_5170);
or U5753 (N_5753,N_4900,N_5065);
or U5754 (N_5754,N_5290,N_5164);
nor U5755 (N_5755,N_4979,N_5028);
or U5756 (N_5756,N_5399,N_5365);
nor U5757 (N_5757,N_4895,N_5050);
nand U5758 (N_5758,N_5261,N_4982);
nand U5759 (N_5759,N_4923,N_5358);
or U5760 (N_5760,N_4956,N_5042);
nand U5761 (N_5761,N_4819,N_5152);
or U5762 (N_5762,N_5339,N_5191);
and U5763 (N_5763,N_5198,N_4850);
or U5764 (N_5764,N_4949,N_5277);
nor U5765 (N_5765,N_5223,N_5334);
or U5766 (N_5766,N_5326,N_5011);
or U5767 (N_5767,N_4954,N_4936);
and U5768 (N_5768,N_4849,N_4856);
nand U5769 (N_5769,N_5252,N_5073);
or U5770 (N_5770,N_5374,N_5024);
nand U5771 (N_5771,N_5122,N_4839);
and U5772 (N_5772,N_5393,N_5274);
nor U5773 (N_5773,N_5347,N_5345);
nor U5774 (N_5774,N_5085,N_5211);
or U5775 (N_5775,N_5353,N_5387);
nand U5776 (N_5776,N_4960,N_5321);
nand U5777 (N_5777,N_4965,N_5394);
or U5778 (N_5778,N_5109,N_5040);
or U5779 (N_5779,N_5084,N_5298);
nor U5780 (N_5780,N_4957,N_4881);
nand U5781 (N_5781,N_4813,N_5121);
nor U5782 (N_5782,N_5088,N_5376);
nor U5783 (N_5783,N_5189,N_4979);
nand U5784 (N_5784,N_4923,N_5002);
nor U5785 (N_5785,N_5366,N_4865);
xor U5786 (N_5786,N_5058,N_5292);
nand U5787 (N_5787,N_4810,N_5133);
nand U5788 (N_5788,N_5164,N_5394);
nor U5789 (N_5789,N_4980,N_4821);
nand U5790 (N_5790,N_4949,N_5137);
and U5791 (N_5791,N_5058,N_4915);
nand U5792 (N_5792,N_4875,N_4983);
or U5793 (N_5793,N_5301,N_5369);
or U5794 (N_5794,N_5167,N_4899);
or U5795 (N_5795,N_5093,N_4937);
or U5796 (N_5796,N_5269,N_5144);
nand U5797 (N_5797,N_4813,N_5294);
or U5798 (N_5798,N_4953,N_5228);
nor U5799 (N_5799,N_5068,N_5094);
nor U5800 (N_5800,N_5279,N_5172);
nand U5801 (N_5801,N_5193,N_5283);
nand U5802 (N_5802,N_4963,N_5120);
or U5803 (N_5803,N_4834,N_4863);
nand U5804 (N_5804,N_4957,N_5255);
nand U5805 (N_5805,N_5001,N_5093);
and U5806 (N_5806,N_5382,N_5114);
nand U5807 (N_5807,N_4816,N_5244);
nand U5808 (N_5808,N_5169,N_5391);
nor U5809 (N_5809,N_5263,N_4876);
and U5810 (N_5810,N_5074,N_4946);
or U5811 (N_5811,N_5332,N_4880);
or U5812 (N_5812,N_5107,N_4838);
nor U5813 (N_5813,N_4822,N_4928);
nor U5814 (N_5814,N_5007,N_4951);
nand U5815 (N_5815,N_5159,N_4970);
xnor U5816 (N_5816,N_4878,N_5368);
nor U5817 (N_5817,N_4882,N_5127);
or U5818 (N_5818,N_5038,N_4887);
nand U5819 (N_5819,N_5228,N_5049);
and U5820 (N_5820,N_4820,N_5121);
or U5821 (N_5821,N_4952,N_5003);
and U5822 (N_5822,N_5056,N_5260);
and U5823 (N_5823,N_4887,N_4877);
or U5824 (N_5824,N_4838,N_5200);
and U5825 (N_5825,N_5253,N_5255);
or U5826 (N_5826,N_4975,N_4813);
or U5827 (N_5827,N_5217,N_5194);
nor U5828 (N_5828,N_5120,N_5228);
nand U5829 (N_5829,N_5115,N_5258);
or U5830 (N_5830,N_4892,N_4863);
or U5831 (N_5831,N_4999,N_4906);
and U5832 (N_5832,N_5141,N_4941);
or U5833 (N_5833,N_4986,N_5130);
nor U5834 (N_5834,N_5073,N_5371);
nand U5835 (N_5835,N_5226,N_5153);
or U5836 (N_5836,N_4821,N_4954);
or U5837 (N_5837,N_5040,N_5387);
nor U5838 (N_5838,N_5320,N_4921);
nand U5839 (N_5839,N_4918,N_5095);
and U5840 (N_5840,N_5144,N_5177);
and U5841 (N_5841,N_5151,N_4973);
or U5842 (N_5842,N_5211,N_5385);
nor U5843 (N_5843,N_5318,N_5004);
and U5844 (N_5844,N_5159,N_4964);
or U5845 (N_5845,N_5122,N_5002);
and U5846 (N_5846,N_4904,N_4837);
nand U5847 (N_5847,N_5044,N_5217);
or U5848 (N_5848,N_4984,N_5070);
and U5849 (N_5849,N_4836,N_4920);
nor U5850 (N_5850,N_5208,N_5226);
nor U5851 (N_5851,N_5103,N_5061);
nand U5852 (N_5852,N_5021,N_5241);
nor U5853 (N_5853,N_5237,N_5184);
or U5854 (N_5854,N_4838,N_5334);
and U5855 (N_5855,N_4908,N_5314);
nor U5856 (N_5856,N_5299,N_4917);
nand U5857 (N_5857,N_5134,N_5233);
and U5858 (N_5858,N_4922,N_5222);
or U5859 (N_5859,N_4974,N_5324);
nor U5860 (N_5860,N_4896,N_5083);
nand U5861 (N_5861,N_4885,N_5161);
nor U5862 (N_5862,N_5189,N_5150);
and U5863 (N_5863,N_5033,N_4847);
and U5864 (N_5864,N_4992,N_5215);
and U5865 (N_5865,N_5140,N_5219);
and U5866 (N_5866,N_5243,N_5267);
nand U5867 (N_5867,N_5064,N_5197);
and U5868 (N_5868,N_5244,N_5175);
and U5869 (N_5869,N_5079,N_4811);
nand U5870 (N_5870,N_5190,N_5032);
and U5871 (N_5871,N_5368,N_5198);
nand U5872 (N_5872,N_4868,N_5223);
or U5873 (N_5873,N_5366,N_5204);
nor U5874 (N_5874,N_5075,N_5207);
and U5875 (N_5875,N_5373,N_5362);
xor U5876 (N_5876,N_4879,N_5080);
and U5877 (N_5877,N_5000,N_5054);
or U5878 (N_5878,N_5131,N_5233);
nor U5879 (N_5879,N_5174,N_5182);
or U5880 (N_5880,N_4954,N_5178);
nor U5881 (N_5881,N_4990,N_4888);
or U5882 (N_5882,N_5204,N_4827);
and U5883 (N_5883,N_5297,N_5019);
and U5884 (N_5884,N_4954,N_5124);
nand U5885 (N_5885,N_5197,N_5154);
or U5886 (N_5886,N_4968,N_5230);
and U5887 (N_5887,N_4843,N_4893);
or U5888 (N_5888,N_5378,N_5053);
nand U5889 (N_5889,N_5183,N_4982);
nor U5890 (N_5890,N_5048,N_5325);
nor U5891 (N_5891,N_5290,N_4824);
nand U5892 (N_5892,N_5166,N_5257);
nor U5893 (N_5893,N_4940,N_5393);
or U5894 (N_5894,N_4904,N_5322);
and U5895 (N_5895,N_4806,N_4937);
nand U5896 (N_5896,N_5335,N_5133);
and U5897 (N_5897,N_5284,N_4868);
nand U5898 (N_5898,N_5326,N_5174);
nand U5899 (N_5899,N_5062,N_5310);
and U5900 (N_5900,N_5385,N_5153);
nand U5901 (N_5901,N_5332,N_5213);
and U5902 (N_5902,N_4896,N_4999);
or U5903 (N_5903,N_5366,N_5143);
or U5904 (N_5904,N_5337,N_5002);
or U5905 (N_5905,N_4851,N_4936);
nand U5906 (N_5906,N_4855,N_4833);
xnor U5907 (N_5907,N_5074,N_5230);
or U5908 (N_5908,N_4966,N_5334);
nor U5909 (N_5909,N_5332,N_5064);
nor U5910 (N_5910,N_5121,N_5148);
or U5911 (N_5911,N_4867,N_5396);
and U5912 (N_5912,N_5390,N_4860);
and U5913 (N_5913,N_5374,N_5084);
nor U5914 (N_5914,N_5391,N_5238);
nor U5915 (N_5915,N_5131,N_5336);
nand U5916 (N_5916,N_5020,N_4895);
nand U5917 (N_5917,N_5267,N_5262);
nor U5918 (N_5918,N_5065,N_4802);
nor U5919 (N_5919,N_4932,N_5174);
and U5920 (N_5920,N_4805,N_4892);
or U5921 (N_5921,N_4938,N_4866);
or U5922 (N_5922,N_5030,N_5011);
nor U5923 (N_5923,N_4966,N_4946);
or U5924 (N_5924,N_4978,N_4925);
xor U5925 (N_5925,N_5132,N_4997);
and U5926 (N_5926,N_5083,N_5142);
or U5927 (N_5927,N_5029,N_5068);
nand U5928 (N_5928,N_5390,N_4822);
xor U5929 (N_5929,N_4874,N_4972);
or U5930 (N_5930,N_5019,N_4877);
nand U5931 (N_5931,N_5380,N_5368);
and U5932 (N_5932,N_5307,N_4879);
and U5933 (N_5933,N_5291,N_5350);
and U5934 (N_5934,N_5259,N_4873);
or U5935 (N_5935,N_4837,N_4832);
nor U5936 (N_5936,N_4927,N_5238);
nor U5937 (N_5937,N_5384,N_5030);
or U5938 (N_5938,N_5291,N_4874);
xnor U5939 (N_5939,N_4907,N_5043);
nand U5940 (N_5940,N_5176,N_5254);
nor U5941 (N_5941,N_4991,N_5136);
and U5942 (N_5942,N_4817,N_5147);
xnor U5943 (N_5943,N_5363,N_4803);
nand U5944 (N_5944,N_5196,N_5000);
and U5945 (N_5945,N_5248,N_4904);
nor U5946 (N_5946,N_5187,N_5133);
and U5947 (N_5947,N_4997,N_5191);
nand U5948 (N_5948,N_4965,N_5349);
or U5949 (N_5949,N_4808,N_5154);
xor U5950 (N_5950,N_5214,N_5068);
or U5951 (N_5951,N_4821,N_5287);
or U5952 (N_5952,N_5313,N_4836);
or U5953 (N_5953,N_4985,N_5111);
nand U5954 (N_5954,N_4864,N_5033);
and U5955 (N_5955,N_4905,N_5189);
and U5956 (N_5956,N_5355,N_5237);
and U5957 (N_5957,N_5364,N_5007);
nand U5958 (N_5958,N_5069,N_5381);
or U5959 (N_5959,N_5198,N_4885);
nor U5960 (N_5960,N_5356,N_5370);
or U5961 (N_5961,N_5296,N_5211);
nand U5962 (N_5962,N_5011,N_4973);
nand U5963 (N_5963,N_5052,N_5161);
or U5964 (N_5964,N_5178,N_5186);
xnor U5965 (N_5965,N_4973,N_5023);
or U5966 (N_5966,N_4823,N_4935);
and U5967 (N_5967,N_5003,N_5083);
and U5968 (N_5968,N_5282,N_5080);
nor U5969 (N_5969,N_4917,N_4818);
and U5970 (N_5970,N_5395,N_4886);
nor U5971 (N_5971,N_5204,N_5083);
nand U5972 (N_5972,N_4804,N_5144);
nand U5973 (N_5973,N_4849,N_5047);
nand U5974 (N_5974,N_5158,N_5088);
nor U5975 (N_5975,N_5185,N_5146);
and U5976 (N_5976,N_5238,N_4985);
nand U5977 (N_5977,N_4840,N_5366);
nor U5978 (N_5978,N_5068,N_5371);
nand U5979 (N_5979,N_5068,N_5370);
and U5980 (N_5980,N_5180,N_5366);
and U5981 (N_5981,N_5288,N_5211);
or U5982 (N_5982,N_5200,N_4816);
and U5983 (N_5983,N_5383,N_4904);
and U5984 (N_5984,N_5020,N_4904);
and U5985 (N_5985,N_5029,N_4827);
or U5986 (N_5986,N_5101,N_5300);
nor U5987 (N_5987,N_5210,N_5041);
nand U5988 (N_5988,N_4866,N_4830);
and U5989 (N_5989,N_4984,N_5192);
nor U5990 (N_5990,N_5023,N_4812);
and U5991 (N_5991,N_4931,N_4825);
and U5992 (N_5992,N_4987,N_4957);
and U5993 (N_5993,N_4890,N_5024);
and U5994 (N_5994,N_4814,N_5103);
nor U5995 (N_5995,N_5373,N_5307);
nor U5996 (N_5996,N_5228,N_5385);
nand U5997 (N_5997,N_4803,N_4945);
and U5998 (N_5998,N_4819,N_4916);
and U5999 (N_5999,N_4893,N_4829);
nand U6000 (N_6000,N_5432,N_5663);
and U6001 (N_6001,N_5622,N_5721);
or U6002 (N_6002,N_5894,N_5883);
or U6003 (N_6003,N_5672,N_5475);
nand U6004 (N_6004,N_5732,N_5849);
nor U6005 (N_6005,N_5743,N_5494);
nand U6006 (N_6006,N_5470,N_5697);
nor U6007 (N_6007,N_5918,N_5689);
nand U6008 (N_6008,N_5940,N_5811);
nand U6009 (N_6009,N_5921,N_5565);
nand U6010 (N_6010,N_5691,N_5758);
nor U6011 (N_6011,N_5944,N_5499);
nor U6012 (N_6012,N_5704,N_5945);
nor U6013 (N_6013,N_5932,N_5805);
and U6014 (N_6014,N_5870,N_5576);
nor U6015 (N_6015,N_5681,N_5603);
and U6016 (N_6016,N_5460,N_5679);
nand U6017 (N_6017,N_5562,N_5736);
nand U6018 (N_6018,N_5986,N_5403);
or U6019 (N_6019,N_5560,N_5786);
nor U6020 (N_6020,N_5517,N_5873);
nand U6021 (N_6021,N_5995,N_5591);
nor U6022 (N_6022,N_5901,N_5429);
xor U6023 (N_6023,N_5557,N_5774);
xnor U6024 (N_6024,N_5535,N_5968);
nor U6025 (N_6025,N_5485,N_5893);
nor U6026 (N_6026,N_5520,N_5440);
or U6027 (N_6027,N_5451,N_5652);
nor U6028 (N_6028,N_5884,N_5513);
nor U6029 (N_6029,N_5990,N_5818);
or U6030 (N_6030,N_5419,N_5843);
nand U6031 (N_6031,N_5505,N_5874);
or U6032 (N_6032,N_5827,N_5751);
or U6033 (N_6033,N_5804,N_5480);
nand U6034 (N_6034,N_5790,N_5872);
and U6035 (N_6035,N_5706,N_5972);
nand U6036 (N_6036,N_5580,N_5406);
and U6037 (N_6037,N_5842,N_5973);
nor U6038 (N_6038,N_5956,N_5529);
or U6039 (N_6039,N_5501,N_5960);
nor U6040 (N_6040,N_5518,N_5851);
and U6041 (N_6041,N_5596,N_5924);
and U6042 (N_6042,N_5631,N_5522);
nand U6043 (N_6043,N_5542,N_5490);
nor U6044 (N_6044,N_5625,N_5477);
and U6045 (N_6045,N_5779,N_5421);
or U6046 (N_6046,N_5910,N_5674);
nand U6047 (N_6047,N_5869,N_5571);
nand U6048 (N_6048,N_5889,N_5902);
or U6049 (N_6049,N_5712,N_5434);
and U6050 (N_6050,N_5589,N_5738);
nand U6051 (N_6051,N_5913,N_5838);
and U6052 (N_6052,N_5664,N_5569);
nor U6053 (N_6053,N_5868,N_5821);
nand U6054 (N_6054,N_5546,N_5961);
nand U6055 (N_6055,N_5802,N_5464);
xor U6056 (N_6056,N_5585,N_5629);
xor U6057 (N_6057,N_5987,N_5498);
nand U6058 (N_6058,N_5436,N_5680);
nand U6059 (N_6059,N_5831,N_5466);
and U6060 (N_6060,N_5447,N_5947);
nand U6061 (N_6061,N_5621,N_5639);
nand U6062 (N_6062,N_5796,N_5531);
or U6063 (N_6063,N_5781,N_5558);
and U6064 (N_6064,N_5538,N_5446);
xor U6065 (N_6065,N_5896,N_5942);
or U6066 (N_6066,N_5782,N_5441);
nand U6067 (N_6067,N_5416,N_5864);
and U6068 (N_6068,N_5525,N_5483);
nand U6069 (N_6069,N_5633,N_5906);
nor U6070 (N_6070,N_5590,N_5530);
nor U6071 (N_6071,N_5524,N_5601);
and U6072 (N_6072,N_5424,N_5948);
xor U6073 (N_6073,N_5701,N_5605);
and U6074 (N_6074,N_5931,N_5439);
and U6075 (N_6075,N_5867,N_5813);
nand U6076 (N_6076,N_5801,N_5482);
or U6077 (N_6077,N_5858,N_5807);
or U6078 (N_6078,N_5481,N_5887);
nand U6079 (N_6079,N_5547,N_5764);
nor U6080 (N_6080,N_5405,N_5928);
or U6081 (N_6081,N_5800,N_5503);
and U6082 (N_6082,N_5404,N_5934);
and U6083 (N_6083,N_5552,N_5541);
nor U6084 (N_6084,N_5567,N_5830);
and U6085 (N_6085,N_5668,N_5991);
and U6086 (N_6086,N_5472,N_5527);
or U6087 (N_6087,N_5904,N_5471);
and U6088 (N_6088,N_5402,N_5555);
nor U6089 (N_6089,N_5602,N_5716);
and U6090 (N_6090,N_5820,N_5719);
and U6091 (N_6091,N_5950,N_5788);
or U6092 (N_6092,N_5620,N_5479);
and U6093 (N_6093,N_5671,N_5880);
and U6094 (N_6094,N_5410,N_5741);
nand U6095 (N_6095,N_5753,N_5614);
or U6096 (N_6096,N_5519,N_5853);
nand U6097 (N_6097,N_5635,N_5778);
nand U6098 (N_6098,N_5927,N_5898);
and U6099 (N_6099,N_5957,N_5919);
and U6100 (N_6100,N_5428,N_5792);
nor U6101 (N_6101,N_5694,N_5638);
or U6102 (N_6102,N_5768,N_5551);
or U6103 (N_6103,N_5840,N_5866);
nor U6104 (N_6104,N_5512,N_5545);
and U6105 (N_6105,N_5992,N_5985);
and U6106 (N_6106,N_5597,N_5666);
nand U6107 (N_6107,N_5740,N_5826);
and U6108 (N_6108,N_5444,N_5568);
and U6109 (N_6109,N_5757,N_5443);
nor U6110 (N_6110,N_5999,N_5715);
or U6111 (N_6111,N_5920,N_5845);
nor U6112 (N_6112,N_5650,N_5452);
nand U6113 (N_6113,N_5900,N_5413);
or U6114 (N_6114,N_5795,N_5577);
or U6115 (N_6115,N_5534,N_5657);
and U6116 (N_6116,N_5967,N_5581);
nor U6117 (N_6117,N_5455,N_5431);
and U6118 (N_6118,N_5963,N_5859);
and U6119 (N_6119,N_5645,N_5854);
nor U6120 (N_6120,N_5579,N_5791);
xnor U6121 (N_6121,N_5862,N_5970);
and U6122 (N_6122,N_5578,N_5739);
and U6123 (N_6123,N_5699,N_5848);
or U6124 (N_6124,N_5613,N_5766);
and U6125 (N_6125,N_5623,N_5426);
and U6126 (N_6126,N_5595,N_5537);
nand U6127 (N_6127,N_5488,N_5946);
and U6128 (N_6128,N_5677,N_5685);
nor U6129 (N_6129,N_5952,N_5911);
xnor U6130 (N_6130,N_5510,N_5616);
or U6131 (N_6131,N_5915,N_5533);
nor U6132 (N_6132,N_5773,N_5411);
nor U6133 (N_6133,N_5574,N_5882);
or U6134 (N_6134,N_5607,N_5815);
nor U6135 (N_6135,N_5700,N_5438);
or U6136 (N_6136,N_5765,N_5762);
nand U6137 (N_6137,N_5926,N_5745);
or U6138 (N_6138,N_5610,N_5702);
or U6139 (N_6139,N_5653,N_5628);
nor U6140 (N_6140,N_5420,N_5606);
nand U6141 (N_6141,N_5632,N_5974);
and U6142 (N_6142,N_5624,N_5717);
nand U6143 (N_6143,N_5852,N_5856);
or U6144 (N_6144,N_5885,N_5727);
or U6145 (N_6145,N_5785,N_5909);
and U6146 (N_6146,N_5756,N_5713);
nand U6147 (N_6147,N_5718,N_5598);
or U6148 (N_6148,N_5509,N_5857);
and U6149 (N_6149,N_5760,N_5618);
and U6150 (N_6150,N_5878,N_5561);
nand U6151 (N_6151,N_5548,N_5695);
and U6152 (N_6152,N_5892,N_5592);
nor U6153 (N_6153,N_5504,N_5759);
nand U6154 (N_6154,N_5746,N_5720);
nand U6155 (N_6155,N_5539,N_5835);
nand U6156 (N_6156,N_5489,N_5834);
nand U6157 (N_6157,N_5445,N_5993);
and U6158 (N_6158,N_5937,N_5556);
nor U6159 (N_6159,N_5980,N_5566);
nor U6160 (N_6160,N_5982,N_5855);
nand U6161 (N_6161,N_5832,N_5954);
nor U6162 (N_6162,N_5500,N_5793);
nand U6163 (N_6163,N_5506,N_5769);
nand U6164 (N_6164,N_5881,N_5922);
xor U6165 (N_6165,N_5861,N_5914);
nand U6166 (N_6166,N_5450,N_5905);
nand U6167 (N_6167,N_5794,N_5863);
or U6168 (N_6168,N_5737,N_5492);
and U6169 (N_6169,N_5593,N_5675);
nor U6170 (N_6170,N_5507,N_5467);
xnor U6171 (N_6171,N_5516,N_5819);
or U6172 (N_6172,N_5449,N_5797);
nor U6173 (N_6173,N_5808,N_5875);
nor U6174 (N_6174,N_5423,N_5977);
or U6175 (N_6175,N_5409,N_5828);
and U6176 (N_6176,N_5733,N_5705);
and U6177 (N_6177,N_5461,N_5619);
and U6178 (N_6178,N_5678,N_5726);
and U6179 (N_6179,N_5860,N_5493);
nor U6180 (N_6180,N_5617,N_5684);
nand U6181 (N_6181,N_5656,N_5630);
and U6182 (N_6182,N_5640,N_5908);
nand U6183 (N_6183,N_5731,N_5983);
nand U6184 (N_6184,N_5708,N_5748);
nor U6185 (N_6185,N_5654,N_5511);
and U6186 (N_6186,N_5953,N_5435);
nand U6187 (N_6187,N_5888,N_5703);
and U6188 (N_6188,N_5770,N_5536);
nor U6189 (N_6189,N_5611,N_5798);
xor U6190 (N_6190,N_5427,N_5641);
xnor U6191 (N_6191,N_5682,N_5814);
nand U6192 (N_6192,N_5456,N_5457);
nor U6193 (N_6193,N_5612,N_5964);
and U6194 (N_6194,N_5923,N_5707);
nor U6195 (N_6195,N_5780,N_5673);
nand U6196 (N_6196,N_5925,N_5809);
and U6197 (N_6197,N_5825,N_5586);
or U6198 (N_6198,N_5609,N_5899);
xor U6199 (N_6199,N_5951,N_5514);
nand U6200 (N_6200,N_5943,N_5763);
or U6201 (N_6201,N_5891,N_5687);
nor U6202 (N_6202,N_5777,N_5554);
and U6203 (N_6203,N_5787,N_5709);
or U6204 (N_6204,N_5588,N_5698);
and U6205 (N_6205,N_5938,N_5949);
nor U6206 (N_6206,N_5474,N_5829);
nor U6207 (N_6207,N_5989,N_5729);
or U6208 (N_6208,N_5600,N_5462);
nand U6209 (N_6209,N_5415,N_5676);
or U6210 (N_6210,N_5941,N_5651);
nor U6211 (N_6211,N_5844,N_5407);
nand U6212 (N_6212,N_5890,N_5803);
and U6213 (N_6213,N_5563,N_5749);
and U6214 (N_6214,N_5484,N_5667);
or U6215 (N_6215,N_5478,N_5917);
or U6216 (N_6216,N_5463,N_5903);
and U6217 (N_6217,N_5907,N_5604);
xor U6218 (N_6218,N_5540,N_5553);
or U6219 (N_6219,N_5839,N_5559);
nand U6220 (N_6220,N_5570,N_5532);
nand U6221 (N_6221,N_5816,N_5508);
nor U6222 (N_6222,N_5955,N_5626);
or U6223 (N_6223,N_5487,N_5933);
or U6224 (N_6224,N_5425,N_5543);
nor U6225 (N_6225,N_5476,N_5752);
or U6226 (N_6226,N_5669,N_5573);
and U6227 (N_6227,N_5806,N_5996);
and U6228 (N_6228,N_5710,N_5637);
and U6229 (N_6229,N_5526,N_5448);
nand U6230 (N_6230,N_5627,N_5496);
nor U6231 (N_6231,N_5877,N_5725);
and U6232 (N_6232,N_5929,N_5583);
nor U6233 (N_6233,N_5935,N_5523);
or U6234 (N_6234,N_5784,N_5418);
nor U6235 (N_6235,N_5783,N_5660);
nand U6236 (N_6236,N_5817,N_5572);
nand U6237 (N_6237,N_5984,N_5966);
or U6238 (N_6238,N_5958,N_5771);
nor U6239 (N_6239,N_5730,N_5458);
nand U6240 (N_6240,N_5822,N_5648);
or U6241 (N_6241,N_5670,N_5647);
nor U6242 (N_6242,N_5750,N_5454);
or U6243 (N_6243,N_5722,N_5442);
or U6244 (N_6244,N_5491,N_5688);
nor U6245 (N_6245,N_5594,N_5912);
nor U6246 (N_6246,N_5564,N_5812);
nor U6247 (N_6247,N_5636,N_5417);
and U6248 (N_6248,N_5661,N_5599);
nand U6249 (N_6249,N_5495,N_5886);
xor U6250 (N_6250,N_5936,N_5846);
or U6251 (N_6251,N_5502,N_5734);
nand U6252 (N_6252,N_5930,N_5401);
nand U6253 (N_6253,N_5690,N_5742);
xor U6254 (N_6254,N_5549,N_5841);
nor U6255 (N_6255,N_5665,N_5473);
and U6256 (N_6256,N_5582,N_5400);
and U6257 (N_6257,N_5959,N_5521);
and U6258 (N_6258,N_5772,N_5998);
xnor U6259 (N_6259,N_5865,N_5544);
and U6260 (N_6260,N_5714,N_5711);
xnor U6261 (N_6261,N_5823,N_5789);
nor U6262 (N_6262,N_5997,N_5646);
and U6263 (N_6263,N_5497,N_5761);
and U6264 (N_6264,N_5895,N_5939);
nor U6265 (N_6265,N_5584,N_5897);
nor U6266 (N_6266,N_5683,N_5747);
nor U6267 (N_6267,N_5981,N_5755);
and U6268 (N_6268,N_5969,N_5836);
and U6269 (N_6269,N_5468,N_5469);
nor U6270 (N_6270,N_5976,N_5988);
nand U6271 (N_6271,N_5414,N_5528);
or U6272 (N_6272,N_5459,N_5412);
and U6273 (N_6273,N_5587,N_5515);
and U6274 (N_6274,N_5810,N_5486);
or U6275 (N_6275,N_5430,N_5658);
or U6276 (N_6276,N_5971,N_5962);
nand U6277 (N_6277,N_5696,N_5837);
nor U6278 (N_6278,N_5979,N_5644);
and U6279 (N_6279,N_5965,N_5408);
nor U6280 (N_6280,N_5833,N_5550);
nand U6281 (N_6281,N_5634,N_5916);
and U6282 (N_6282,N_5754,N_5876);
and U6283 (N_6283,N_5615,N_5799);
or U6284 (N_6284,N_5728,N_5693);
and U6285 (N_6285,N_5994,N_5453);
and U6286 (N_6286,N_5850,N_5692);
nand U6287 (N_6287,N_5649,N_5775);
or U6288 (N_6288,N_5978,N_5824);
nand U6289 (N_6289,N_5723,N_5767);
and U6290 (N_6290,N_5662,N_5465);
nor U6291 (N_6291,N_5975,N_5437);
or U6292 (N_6292,N_5879,N_5659);
or U6293 (N_6293,N_5847,N_5776);
and U6294 (N_6294,N_5643,N_5871);
nor U6295 (N_6295,N_5433,N_5686);
nor U6296 (N_6296,N_5744,N_5422);
nor U6297 (N_6297,N_5608,N_5655);
or U6298 (N_6298,N_5642,N_5724);
or U6299 (N_6299,N_5575,N_5735);
or U6300 (N_6300,N_5965,N_5800);
and U6301 (N_6301,N_5571,N_5447);
and U6302 (N_6302,N_5928,N_5509);
or U6303 (N_6303,N_5907,N_5441);
or U6304 (N_6304,N_5483,N_5836);
nand U6305 (N_6305,N_5580,N_5737);
xor U6306 (N_6306,N_5657,N_5741);
and U6307 (N_6307,N_5535,N_5940);
nand U6308 (N_6308,N_5411,N_5639);
and U6309 (N_6309,N_5982,N_5937);
or U6310 (N_6310,N_5899,N_5525);
or U6311 (N_6311,N_5985,N_5504);
or U6312 (N_6312,N_5619,N_5800);
or U6313 (N_6313,N_5682,N_5965);
nor U6314 (N_6314,N_5484,N_5858);
nor U6315 (N_6315,N_5762,N_5464);
xnor U6316 (N_6316,N_5624,N_5637);
nor U6317 (N_6317,N_5418,N_5875);
nor U6318 (N_6318,N_5664,N_5862);
nand U6319 (N_6319,N_5741,N_5739);
nand U6320 (N_6320,N_5449,N_5739);
nand U6321 (N_6321,N_5786,N_5641);
nor U6322 (N_6322,N_5646,N_5754);
nor U6323 (N_6323,N_5806,N_5974);
nand U6324 (N_6324,N_5501,N_5680);
nor U6325 (N_6325,N_5833,N_5941);
nand U6326 (N_6326,N_5806,N_5887);
or U6327 (N_6327,N_5965,N_5659);
nor U6328 (N_6328,N_5656,N_5585);
or U6329 (N_6329,N_5797,N_5799);
nand U6330 (N_6330,N_5591,N_5563);
nor U6331 (N_6331,N_5863,N_5460);
nor U6332 (N_6332,N_5514,N_5905);
nand U6333 (N_6333,N_5807,N_5663);
nand U6334 (N_6334,N_5792,N_5418);
and U6335 (N_6335,N_5916,N_5714);
nor U6336 (N_6336,N_5691,N_5752);
and U6337 (N_6337,N_5915,N_5976);
or U6338 (N_6338,N_5823,N_5617);
and U6339 (N_6339,N_5604,N_5573);
or U6340 (N_6340,N_5888,N_5543);
and U6341 (N_6341,N_5869,N_5404);
or U6342 (N_6342,N_5676,N_5642);
nand U6343 (N_6343,N_5727,N_5863);
or U6344 (N_6344,N_5442,N_5792);
or U6345 (N_6345,N_5966,N_5522);
nor U6346 (N_6346,N_5647,N_5784);
or U6347 (N_6347,N_5517,N_5545);
nand U6348 (N_6348,N_5925,N_5986);
or U6349 (N_6349,N_5914,N_5889);
and U6350 (N_6350,N_5693,N_5823);
and U6351 (N_6351,N_5983,N_5991);
nor U6352 (N_6352,N_5961,N_5424);
xor U6353 (N_6353,N_5421,N_5508);
or U6354 (N_6354,N_5856,N_5987);
and U6355 (N_6355,N_5554,N_5711);
nand U6356 (N_6356,N_5568,N_5633);
nor U6357 (N_6357,N_5894,N_5819);
and U6358 (N_6358,N_5696,N_5744);
or U6359 (N_6359,N_5897,N_5451);
and U6360 (N_6360,N_5709,N_5778);
nor U6361 (N_6361,N_5923,N_5928);
and U6362 (N_6362,N_5886,N_5665);
nand U6363 (N_6363,N_5962,N_5867);
xor U6364 (N_6364,N_5418,N_5776);
nand U6365 (N_6365,N_5751,N_5447);
and U6366 (N_6366,N_5720,N_5947);
nand U6367 (N_6367,N_5603,N_5530);
nand U6368 (N_6368,N_5873,N_5826);
or U6369 (N_6369,N_5720,N_5803);
nor U6370 (N_6370,N_5591,N_5630);
nand U6371 (N_6371,N_5474,N_5467);
nand U6372 (N_6372,N_5850,N_5571);
and U6373 (N_6373,N_5917,N_5922);
and U6374 (N_6374,N_5490,N_5872);
nor U6375 (N_6375,N_5554,N_5835);
nand U6376 (N_6376,N_5729,N_5448);
xnor U6377 (N_6377,N_5808,N_5764);
nor U6378 (N_6378,N_5812,N_5464);
nor U6379 (N_6379,N_5996,N_5514);
nor U6380 (N_6380,N_5403,N_5836);
nand U6381 (N_6381,N_5711,N_5530);
and U6382 (N_6382,N_5543,N_5968);
or U6383 (N_6383,N_5532,N_5530);
and U6384 (N_6384,N_5680,N_5662);
or U6385 (N_6385,N_5561,N_5779);
or U6386 (N_6386,N_5733,N_5485);
or U6387 (N_6387,N_5944,N_5757);
nor U6388 (N_6388,N_5996,N_5759);
nand U6389 (N_6389,N_5643,N_5915);
nand U6390 (N_6390,N_5845,N_5727);
or U6391 (N_6391,N_5708,N_5579);
nand U6392 (N_6392,N_5603,N_5777);
nand U6393 (N_6393,N_5559,N_5912);
nand U6394 (N_6394,N_5671,N_5490);
or U6395 (N_6395,N_5536,N_5895);
or U6396 (N_6396,N_5679,N_5443);
or U6397 (N_6397,N_5637,N_5400);
nand U6398 (N_6398,N_5596,N_5419);
nand U6399 (N_6399,N_5627,N_5990);
nor U6400 (N_6400,N_5576,N_5527);
and U6401 (N_6401,N_5828,N_5487);
nor U6402 (N_6402,N_5712,N_5940);
or U6403 (N_6403,N_5785,N_5908);
nand U6404 (N_6404,N_5848,N_5859);
nand U6405 (N_6405,N_5752,N_5450);
and U6406 (N_6406,N_5928,N_5796);
nand U6407 (N_6407,N_5607,N_5854);
nand U6408 (N_6408,N_5536,N_5905);
or U6409 (N_6409,N_5588,N_5581);
nor U6410 (N_6410,N_5915,N_5722);
and U6411 (N_6411,N_5797,N_5519);
nor U6412 (N_6412,N_5576,N_5726);
or U6413 (N_6413,N_5608,N_5723);
nor U6414 (N_6414,N_5798,N_5532);
and U6415 (N_6415,N_5560,N_5696);
and U6416 (N_6416,N_5617,N_5422);
xnor U6417 (N_6417,N_5965,N_5825);
nand U6418 (N_6418,N_5446,N_5923);
and U6419 (N_6419,N_5891,N_5960);
nor U6420 (N_6420,N_5756,N_5488);
nor U6421 (N_6421,N_5472,N_5777);
and U6422 (N_6422,N_5622,N_5912);
and U6423 (N_6423,N_5610,N_5405);
nor U6424 (N_6424,N_5661,N_5500);
and U6425 (N_6425,N_5610,N_5513);
nand U6426 (N_6426,N_5706,N_5415);
and U6427 (N_6427,N_5829,N_5418);
or U6428 (N_6428,N_5955,N_5993);
and U6429 (N_6429,N_5680,N_5957);
nand U6430 (N_6430,N_5450,N_5633);
nand U6431 (N_6431,N_5630,N_5675);
nand U6432 (N_6432,N_5524,N_5493);
and U6433 (N_6433,N_5656,N_5738);
nand U6434 (N_6434,N_5486,N_5918);
or U6435 (N_6435,N_5971,N_5534);
or U6436 (N_6436,N_5604,N_5727);
and U6437 (N_6437,N_5757,N_5433);
and U6438 (N_6438,N_5727,N_5805);
nand U6439 (N_6439,N_5460,N_5729);
or U6440 (N_6440,N_5471,N_5790);
nor U6441 (N_6441,N_5527,N_5598);
or U6442 (N_6442,N_5569,N_5575);
and U6443 (N_6443,N_5510,N_5694);
and U6444 (N_6444,N_5459,N_5841);
or U6445 (N_6445,N_5582,N_5861);
nor U6446 (N_6446,N_5686,N_5757);
or U6447 (N_6447,N_5982,N_5439);
or U6448 (N_6448,N_5673,N_5698);
nand U6449 (N_6449,N_5769,N_5807);
or U6450 (N_6450,N_5833,N_5558);
nand U6451 (N_6451,N_5624,N_5933);
xnor U6452 (N_6452,N_5437,N_5655);
nand U6453 (N_6453,N_5761,N_5637);
and U6454 (N_6454,N_5619,N_5632);
or U6455 (N_6455,N_5612,N_5716);
nand U6456 (N_6456,N_5443,N_5781);
nand U6457 (N_6457,N_5653,N_5953);
nand U6458 (N_6458,N_5831,N_5813);
nor U6459 (N_6459,N_5904,N_5881);
or U6460 (N_6460,N_5571,N_5916);
nor U6461 (N_6461,N_5514,N_5537);
nand U6462 (N_6462,N_5709,N_5741);
and U6463 (N_6463,N_5832,N_5674);
and U6464 (N_6464,N_5789,N_5615);
and U6465 (N_6465,N_5982,N_5592);
or U6466 (N_6466,N_5770,N_5599);
and U6467 (N_6467,N_5597,N_5621);
or U6468 (N_6468,N_5457,N_5437);
nor U6469 (N_6469,N_5898,N_5418);
and U6470 (N_6470,N_5401,N_5546);
or U6471 (N_6471,N_5453,N_5715);
or U6472 (N_6472,N_5553,N_5642);
nor U6473 (N_6473,N_5757,N_5430);
and U6474 (N_6474,N_5626,N_5647);
or U6475 (N_6475,N_5895,N_5862);
nor U6476 (N_6476,N_5848,N_5463);
and U6477 (N_6477,N_5620,N_5658);
and U6478 (N_6478,N_5408,N_5793);
nor U6479 (N_6479,N_5424,N_5583);
or U6480 (N_6480,N_5961,N_5913);
xnor U6481 (N_6481,N_5866,N_5752);
nor U6482 (N_6482,N_5612,N_5915);
or U6483 (N_6483,N_5511,N_5625);
nand U6484 (N_6484,N_5779,N_5677);
or U6485 (N_6485,N_5498,N_5679);
and U6486 (N_6486,N_5698,N_5998);
and U6487 (N_6487,N_5488,N_5670);
and U6488 (N_6488,N_5409,N_5459);
and U6489 (N_6489,N_5587,N_5608);
nor U6490 (N_6490,N_5851,N_5964);
nor U6491 (N_6491,N_5618,N_5799);
and U6492 (N_6492,N_5915,N_5833);
xnor U6493 (N_6493,N_5427,N_5788);
nand U6494 (N_6494,N_5598,N_5906);
and U6495 (N_6495,N_5861,N_5611);
and U6496 (N_6496,N_5522,N_5850);
nor U6497 (N_6497,N_5887,N_5696);
xnor U6498 (N_6498,N_5620,N_5697);
nor U6499 (N_6499,N_5802,N_5859);
or U6500 (N_6500,N_5628,N_5849);
nand U6501 (N_6501,N_5871,N_5515);
nand U6502 (N_6502,N_5799,N_5832);
nor U6503 (N_6503,N_5638,N_5790);
and U6504 (N_6504,N_5925,N_5961);
or U6505 (N_6505,N_5474,N_5957);
and U6506 (N_6506,N_5407,N_5937);
nand U6507 (N_6507,N_5940,N_5959);
nor U6508 (N_6508,N_5455,N_5568);
nor U6509 (N_6509,N_5579,N_5422);
or U6510 (N_6510,N_5420,N_5903);
nand U6511 (N_6511,N_5977,N_5605);
or U6512 (N_6512,N_5683,N_5986);
nand U6513 (N_6513,N_5553,N_5439);
nand U6514 (N_6514,N_5983,N_5838);
nor U6515 (N_6515,N_5450,N_5599);
nand U6516 (N_6516,N_5750,N_5772);
and U6517 (N_6517,N_5523,N_5970);
nand U6518 (N_6518,N_5463,N_5870);
and U6519 (N_6519,N_5653,N_5861);
nand U6520 (N_6520,N_5666,N_5830);
nor U6521 (N_6521,N_5972,N_5550);
nand U6522 (N_6522,N_5704,N_5862);
and U6523 (N_6523,N_5517,N_5643);
nor U6524 (N_6524,N_5462,N_5665);
or U6525 (N_6525,N_5882,N_5466);
nor U6526 (N_6526,N_5619,N_5477);
or U6527 (N_6527,N_5643,N_5576);
nor U6528 (N_6528,N_5655,N_5509);
and U6529 (N_6529,N_5995,N_5916);
nor U6530 (N_6530,N_5416,N_5548);
nand U6531 (N_6531,N_5981,N_5400);
nor U6532 (N_6532,N_5695,N_5700);
nor U6533 (N_6533,N_5673,N_5645);
nand U6534 (N_6534,N_5986,N_5513);
nand U6535 (N_6535,N_5511,N_5823);
nand U6536 (N_6536,N_5419,N_5446);
and U6537 (N_6537,N_5943,N_5561);
or U6538 (N_6538,N_5578,N_5623);
or U6539 (N_6539,N_5584,N_5488);
nor U6540 (N_6540,N_5720,N_5683);
xor U6541 (N_6541,N_5916,N_5788);
nand U6542 (N_6542,N_5425,N_5811);
or U6543 (N_6543,N_5810,N_5602);
nand U6544 (N_6544,N_5642,N_5997);
nand U6545 (N_6545,N_5995,N_5983);
or U6546 (N_6546,N_5492,N_5673);
nor U6547 (N_6547,N_5533,N_5880);
or U6548 (N_6548,N_5410,N_5655);
or U6549 (N_6549,N_5514,N_5556);
nor U6550 (N_6550,N_5494,N_5448);
nand U6551 (N_6551,N_5940,N_5955);
nand U6552 (N_6552,N_5642,N_5751);
nor U6553 (N_6553,N_5624,N_5568);
and U6554 (N_6554,N_5840,N_5772);
nand U6555 (N_6555,N_5487,N_5495);
nor U6556 (N_6556,N_5471,N_5555);
and U6557 (N_6557,N_5520,N_5789);
nor U6558 (N_6558,N_5526,N_5484);
and U6559 (N_6559,N_5545,N_5840);
or U6560 (N_6560,N_5584,N_5614);
or U6561 (N_6561,N_5418,N_5949);
or U6562 (N_6562,N_5815,N_5891);
nand U6563 (N_6563,N_5973,N_5892);
and U6564 (N_6564,N_5810,N_5589);
and U6565 (N_6565,N_5732,N_5519);
or U6566 (N_6566,N_5961,N_5780);
nand U6567 (N_6567,N_5814,N_5577);
and U6568 (N_6568,N_5609,N_5552);
nand U6569 (N_6569,N_5958,N_5445);
or U6570 (N_6570,N_5960,N_5782);
or U6571 (N_6571,N_5953,N_5951);
and U6572 (N_6572,N_5662,N_5698);
or U6573 (N_6573,N_5985,N_5625);
and U6574 (N_6574,N_5617,N_5421);
or U6575 (N_6575,N_5461,N_5850);
nand U6576 (N_6576,N_5939,N_5849);
nand U6577 (N_6577,N_5998,N_5512);
or U6578 (N_6578,N_5507,N_5567);
nor U6579 (N_6579,N_5450,N_5755);
nand U6580 (N_6580,N_5527,N_5631);
nor U6581 (N_6581,N_5875,N_5572);
nor U6582 (N_6582,N_5674,N_5913);
or U6583 (N_6583,N_5614,N_5906);
nand U6584 (N_6584,N_5820,N_5850);
nand U6585 (N_6585,N_5660,N_5816);
or U6586 (N_6586,N_5809,N_5930);
or U6587 (N_6587,N_5482,N_5931);
or U6588 (N_6588,N_5925,N_5767);
and U6589 (N_6589,N_5965,N_5994);
nor U6590 (N_6590,N_5662,N_5577);
and U6591 (N_6591,N_5621,N_5470);
nand U6592 (N_6592,N_5884,N_5623);
and U6593 (N_6593,N_5874,N_5591);
or U6594 (N_6594,N_5936,N_5490);
or U6595 (N_6595,N_5962,N_5947);
nand U6596 (N_6596,N_5562,N_5626);
nor U6597 (N_6597,N_5716,N_5523);
nor U6598 (N_6598,N_5647,N_5522);
nand U6599 (N_6599,N_5671,N_5720);
or U6600 (N_6600,N_6553,N_6211);
and U6601 (N_6601,N_6357,N_6468);
nor U6602 (N_6602,N_6419,N_6339);
nor U6603 (N_6603,N_6016,N_6459);
nand U6604 (N_6604,N_6060,N_6243);
and U6605 (N_6605,N_6286,N_6565);
nand U6606 (N_6606,N_6163,N_6203);
and U6607 (N_6607,N_6237,N_6366);
nand U6608 (N_6608,N_6253,N_6088);
nand U6609 (N_6609,N_6241,N_6020);
nor U6610 (N_6610,N_6127,N_6529);
and U6611 (N_6611,N_6336,N_6255);
nor U6612 (N_6612,N_6526,N_6348);
or U6613 (N_6613,N_6099,N_6170);
or U6614 (N_6614,N_6591,N_6145);
nor U6615 (N_6615,N_6083,N_6316);
nand U6616 (N_6616,N_6311,N_6065);
or U6617 (N_6617,N_6374,N_6261);
nor U6618 (N_6618,N_6475,N_6530);
nor U6619 (N_6619,N_6157,N_6148);
nand U6620 (N_6620,N_6054,N_6318);
nor U6621 (N_6621,N_6461,N_6572);
and U6622 (N_6622,N_6308,N_6111);
or U6623 (N_6623,N_6595,N_6043);
or U6624 (N_6624,N_6588,N_6413);
or U6625 (N_6625,N_6491,N_6452);
nand U6626 (N_6626,N_6039,N_6110);
nor U6627 (N_6627,N_6564,N_6106);
nand U6628 (N_6628,N_6257,N_6375);
and U6629 (N_6629,N_6151,N_6301);
nor U6630 (N_6630,N_6554,N_6424);
or U6631 (N_6631,N_6382,N_6482);
nand U6632 (N_6632,N_6469,N_6297);
nor U6633 (N_6633,N_6403,N_6354);
and U6634 (N_6634,N_6173,N_6159);
and U6635 (N_6635,N_6149,N_6304);
xor U6636 (N_6636,N_6046,N_6494);
nand U6637 (N_6637,N_6119,N_6195);
or U6638 (N_6638,N_6386,N_6266);
or U6639 (N_6639,N_6463,N_6271);
nor U6640 (N_6640,N_6277,N_6324);
and U6641 (N_6641,N_6184,N_6226);
or U6642 (N_6642,N_6189,N_6567);
and U6643 (N_6643,N_6175,N_6546);
nand U6644 (N_6644,N_6185,N_6209);
and U6645 (N_6645,N_6230,N_6381);
or U6646 (N_6646,N_6109,N_6490);
nor U6647 (N_6647,N_6280,N_6344);
nand U6648 (N_6648,N_6136,N_6421);
and U6649 (N_6649,N_6462,N_6331);
and U6650 (N_6650,N_6125,N_6275);
nand U6651 (N_6651,N_6001,N_6259);
or U6652 (N_6652,N_6502,N_6333);
and U6653 (N_6653,N_6343,N_6368);
and U6654 (N_6654,N_6483,N_6210);
nand U6655 (N_6655,N_6228,N_6037);
nand U6656 (N_6656,N_6577,N_6300);
nor U6657 (N_6657,N_6496,N_6342);
and U6658 (N_6658,N_6295,N_6090);
or U6659 (N_6659,N_6123,N_6080);
nand U6660 (N_6660,N_6035,N_6156);
and U6661 (N_6661,N_6009,N_6448);
nand U6662 (N_6662,N_6356,N_6247);
and U6663 (N_6663,N_6434,N_6476);
and U6664 (N_6664,N_6076,N_6274);
or U6665 (N_6665,N_6555,N_6458);
nor U6666 (N_6666,N_6194,N_6025);
and U6667 (N_6667,N_6484,N_6442);
or U6668 (N_6668,N_6500,N_6117);
nand U6669 (N_6669,N_6390,N_6049);
and U6670 (N_6670,N_6281,N_6227);
or U6671 (N_6671,N_6066,N_6470);
and U6672 (N_6672,N_6004,N_6124);
or U6673 (N_6673,N_6018,N_6244);
nor U6674 (N_6674,N_6044,N_6391);
nor U6675 (N_6675,N_6379,N_6341);
nand U6676 (N_6676,N_6140,N_6177);
nand U6677 (N_6677,N_6078,N_6235);
or U6678 (N_6678,N_6457,N_6309);
and U6679 (N_6679,N_6139,N_6003);
and U6680 (N_6680,N_6351,N_6538);
nand U6681 (N_6681,N_6191,N_6095);
nor U6682 (N_6682,N_6401,N_6207);
nor U6683 (N_6683,N_6371,N_6063);
and U6684 (N_6684,N_6179,N_6539);
and U6685 (N_6685,N_6188,N_6542);
nor U6686 (N_6686,N_6597,N_6332);
nand U6687 (N_6687,N_6528,N_6430);
nand U6688 (N_6688,N_6330,N_6570);
and U6689 (N_6689,N_6079,N_6014);
xnor U6690 (N_6690,N_6019,N_6052);
and U6691 (N_6691,N_6422,N_6556);
and U6692 (N_6692,N_6094,N_6328);
nor U6693 (N_6693,N_6254,N_6130);
and U6694 (N_6694,N_6472,N_6074);
nor U6695 (N_6695,N_6396,N_6165);
nor U6696 (N_6696,N_6326,N_6447);
or U6697 (N_6697,N_6267,N_6134);
and U6698 (N_6698,N_6536,N_6091);
nor U6699 (N_6699,N_6384,N_6239);
nor U6700 (N_6700,N_6006,N_6238);
nor U6701 (N_6701,N_6439,N_6560);
nand U6702 (N_6702,N_6017,N_6135);
nand U6703 (N_6703,N_6105,N_6425);
or U6704 (N_6704,N_6535,N_6305);
and U6705 (N_6705,N_6455,N_6503);
nand U6706 (N_6706,N_6005,N_6206);
or U6707 (N_6707,N_6093,N_6168);
xor U6708 (N_6708,N_6389,N_6081);
and U6709 (N_6709,N_6508,N_6432);
or U6710 (N_6710,N_6543,N_6373);
nor U6711 (N_6711,N_6224,N_6214);
nor U6712 (N_6712,N_6319,N_6306);
or U6713 (N_6713,N_6249,N_6196);
nand U6714 (N_6714,N_6427,N_6531);
or U6715 (N_6715,N_6062,N_6186);
nor U6716 (N_6716,N_6493,N_6086);
or U6717 (N_6717,N_6598,N_6272);
or U6718 (N_6718,N_6585,N_6176);
nand U6719 (N_6719,N_6164,N_6467);
or U6720 (N_6720,N_6370,N_6576);
and U6721 (N_6721,N_6315,N_6358);
and U6722 (N_6722,N_6116,N_6312);
or U6723 (N_6723,N_6166,N_6096);
and U6724 (N_6724,N_6563,N_6103);
or U6725 (N_6725,N_6141,N_6441);
nand U6726 (N_6726,N_6040,N_6032);
nand U6727 (N_6727,N_6547,N_6417);
nand U6728 (N_6728,N_6561,N_6497);
and U6729 (N_6729,N_6558,N_6488);
or U6730 (N_6730,N_6222,N_6256);
and U6731 (N_6731,N_6152,N_6030);
nand U6732 (N_6732,N_6002,N_6592);
nor U6733 (N_6733,N_6479,N_6337);
or U6734 (N_6734,N_6213,N_6012);
or U6735 (N_6735,N_6340,N_6192);
nand U6736 (N_6736,N_6541,N_6571);
nand U6737 (N_6737,N_6533,N_6101);
nand U6738 (N_6738,N_6397,N_6445);
nand U6739 (N_6739,N_6008,N_6169);
xnor U6740 (N_6740,N_6137,N_6360);
nand U6741 (N_6741,N_6033,N_6248);
and U6742 (N_6742,N_6583,N_6011);
or U6743 (N_6743,N_6321,N_6231);
and U6744 (N_6744,N_6551,N_6378);
and U6745 (N_6745,N_6399,N_6132);
or U6746 (N_6746,N_6143,N_6223);
nand U6747 (N_6747,N_6376,N_6519);
nor U6748 (N_6748,N_6505,N_6064);
nor U6749 (N_6749,N_6015,N_6501);
nand U6750 (N_6750,N_6013,N_6404);
nand U6751 (N_6751,N_6084,N_6205);
nand U6752 (N_6752,N_6512,N_6120);
nand U6753 (N_6753,N_6473,N_6456);
nand U6754 (N_6754,N_6147,N_6359);
or U6755 (N_6755,N_6590,N_6045);
nand U6756 (N_6756,N_6245,N_6022);
xor U6757 (N_6757,N_6051,N_6294);
and U6758 (N_6758,N_6029,N_6055);
and U6759 (N_6759,N_6580,N_6112);
nand U6760 (N_6760,N_6050,N_6414);
nor U6761 (N_6761,N_6515,N_6487);
and U6762 (N_6762,N_6593,N_6158);
nand U6763 (N_6763,N_6562,N_6114);
or U6764 (N_6764,N_6265,N_6068);
and U6765 (N_6765,N_6446,N_6278);
and U6766 (N_6766,N_6586,N_6292);
nor U6767 (N_6767,N_6128,N_6489);
nor U6768 (N_6768,N_6537,N_6516);
nor U6769 (N_6769,N_6041,N_6513);
or U6770 (N_6770,N_6465,N_6104);
or U6771 (N_6771,N_6569,N_6178);
or U6772 (N_6772,N_6418,N_6024);
and U6773 (N_6773,N_6216,N_6365);
and U6774 (N_6774,N_6161,N_6581);
xnor U6775 (N_6775,N_6545,N_6480);
xor U6776 (N_6776,N_6440,N_6320);
nand U6777 (N_6777,N_6036,N_6225);
nand U6778 (N_6778,N_6303,N_6100);
and U6779 (N_6779,N_6221,N_6477);
or U6780 (N_6780,N_6089,N_6408);
or U6781 (N_6781,N_6108,N_6388);
nor U6782 (N_6782,N_6346,N_6097);
and U6783 (N_6783,N_6171,N_6270);
nor U6784 (N_6784,N_6474,N_6183);
nor U6785 (N_6785,N_6436,N_6352);
and U6786 (N_6786,N_6293,N_6220);
nand U6787 (N_6787,N_6387,N_6288);
or U6788 (N_6788,N_6058,N_6260);
and U6789 (N_6789,N_6144,N_6098);
nor U6790 (N_6790,N_6416,N_6420);
and U6791 (N_6791,N_6240,N_6402);
and U6792 (N_6792,N_6521,N_6251);
xnor U6793 (N_6793,N_6287,N_6478);
nor U6794 (N_6794,N_6252,N_6550);
nor U6795 (N_6795,N_6372,N_6217);
nand U6796 (N_6796,N_6575,N_6566);
nor U6797 (N_6797,N_6510,N_6444);
nand U6798 (N_6798,N_6527,N_6578);
nor U6799 (N_6799,N_6559,N_6518);
nor U6800 (N_6800,N_6453,N_6367);
or U6801 (N_6801,N_6437,N_6540);
nor U6802 (N_6802,N_6023,N_6353);
or U6803 (N_6803,N_6509,N_6138);
and U6804 (N_6804,N_6302,N_6317);
or U6805 (N_6805,N_6038,N_6589);
nor U6806 (N_6806,N_6236,N_6506);
nor U6807 (N_6807,N_6407,N_6197);
nor U6808 (N_6808,N_6454,N_6485);
nand U6809 (N_6809,N_6394,N_6071);
nand U6810 (N_6810,N_6059,N_6579);
and U6811 (N_6811,N_6073,N_6406);
xnor U6812 (N_6812,N_6327,N_6299);
xor U6813 (N_6813,N_6587,N_6481);
nor U6814 (N_6814,N_6273,N_6524);
and U6815 (N_6815,N_6498,N_6131);
nor U6816 (N_6816,N_6258,N_6544);
nor U6817 (N_6817,N_6268,N_6582);
or U6818 (N_6818,N_6363,N_6048);
and U6819 (N_6819,N_6426,N_6409);
nand U6820 (N_6820,N_6229,N_6338);
nand U6821 (N_6821,N_6599,N_6435);
nand U6822 (N_6822,N_6193,N_6466);
and U6823 (N_6823,N_6107,N_6057);
or U6824 (N_6824,N_6122,N_6250);
nor U6825 (N_6825,N_6167,N_6329);
nand U6826 (N_6826,N_6190,N_6150);
nand U6827 (N_6827,N_6180,N_6443);
nor U6828 (N_6828,N_6548,N_6198);
nand U6829 (N_6829,N_6082,N_6429);
or U6830 (N_6830,N_6400,N_6153);
xnor U6831 (N_6831,N_6115,N_6282);
or U6832 (N_6832,N_6160,N_6072);
or U6833 (N_6833,N_6200,N_6395);
nand U6834 (N_6834,N_6307,N_6233);
nor U6835 (N_6835,N_6405,N_6507);
nor U6836 (N_6836,N_6042,N_6380);
nor U6837 (N_6837,N_6323,N_6557);
nand U6838 (N_6838,N_6596,N_6199);
nand U6839 (N_6839,N_6313,N_6517);
nor U6840 (N_6840,N_6263,N_6383);
and U6841 (N_6841,N_6129,N_6034);
or U6842 (N_6842,N_6504,N_6298);
nor U6843 (N_6843,N_6499,N_6289);
or U6844 (N_6844,N_6495,N_6511);
nor U6845 (N_6845,N_6269,N_6285);
or U6846 (N_6846,N_6262,N_6102);
and U6847 (N_6847,N_6242,N_6549);
nor U6848 (N_6848,N_6296,N_6234);
nor U6849 (N_6849,N_6449,N_6181);
and U6850 (N_6850,N_6075,N_6172);
and U6851 (N_6851,N_6087,N_6412);
and U6852 (N_6852,N_6438,N_6369);
nor U6853 (N_6853,N_6431,N_6182);
or U6854 (N_6854,N_6520,N_6215);
nand U6855 (N_6855,N_6146,N_6028);
or U6856 (N_6856,N_6026,N_6314);
nor U6857 (N_6857,N_6212,N_6347);
nor U6858 (N_6858,N_6154,N_6364);
nand U6859 (N_6859,N_6155,N_6232);
and U6860 (N_6860,N_6433,N_6492);
nor U6861 (N_6861,N_6471,N_6010);
and U6862 (N_6862,N_6202,N_6392);
and U6863 (N_6863,N_6218,N_6522);
nor U6864 (N_6864,N_6070,N_6007);
or U6865 (N_6865,N_6092,N_6126);
nor U6866 (N_6866,N_6335,N_6279);
nand U6867 (N_6867,N_6514,N_6423);
and U6868 (N_6868,N_6061,N_6276);
or U6869 (N_6869,N_6573,N_6047);
or U6870 (N_6870,N_6568,N_6322);
or U6871 (N_6871,N_6532,N_6053);
nand U6872 (N_6872,N_6345,N_6118);
nor U6873 (N_6873,N_6486,N_6113);
nand U6874 (N_6874,N_6460,N_6219);
and U6875 (N_6875,N_6398,N_6162);
and U6876 (N_6876,N_6334,N_6450);
and U6877 (N_6877,N_6362,N_6584);
nor U6878 (N_6878,N_6208,N_6534);
or U6879 (N_6879,N_6451,N_6085);
and U6880 (N_6880,N_6246,N_6415);
and U6881 (N_6881,N_6464,N_6290);
or U6882 (N_6882,N_6411,N_6349);
nor U6883 (N_6883,N_6574,N_6201);
and U6884 (N_6884,N_6355,N_6031);
nor U6885 (N_6885,N_6552,N_6067);
nand U6886 (N_6886,N_6264,N_6077);
nand U6887 (N_6887,N_6133,N_6377);
and U6888 (N_6888,N_6594,N_6350);
and U6889 (N_6889,N_6283,N_6056);
and U6890 (N_6890,N_6121,N_6000);
nor U6891 (N_6891,N_6291,N_6204);
or U6892 (N_6892,N_6393,N_6027);
and U6893 (N_6893,N_6361,N_6310);
nand U6894 (N_6894,N_6284,N_6523);
nor U6895 (N_6895,N_6142,N_6187);
or U6896 (N_6896,N_6021,N_6325);
and U6897 (N_6897,N_6069,N_6525);
and U6898 (N_6898,N_6428,N_6385);
nand U6899 (N_6899,N_6174,N_6410);
and U6900 (N_6900,N_6476,N_6202);
nand U6901 (N_6901,N_6014,N_6083);
xnor U6902 (N_6902,N_6301,N_6444);
or U6903 (N_6903,N_6097,N_6167);
nand U6904 (N_6904,N_6353,N_6213);
nand U6905 (N_6905,N_6134,N_6538);
and U6906 (N_6906,N_6459,N_6303);
nand U6907 (N_6907,N_6232,N_6367);
nand U6908 (N_6908,N_6039,N_6192);
nand U6909 (N_6909,N_6162,N_6167);
or U6910 (N_6910,N_6552,N_6336);
nor U6911 (N_6911,N_6594,N_6257);
and U6912 (N_6912,N_6501,N_6598);
nor U6913 (N_6913,N_6273,N_6101);
or U6914 (N_6914,N_6346,N_6366);
or U6915 (N_6915,N_6208,N_6112);
nor U6916 (N_6916,N_6382,N_6007);
or U6917 (N_6917,N_6056,N_6027);
and U6918 (N_6918,N_6177,N_6217);
and U6919 (N_6919,N_6113,N_6212);
xnor U6920 (N_6920,N_6428,N_6284);
nor U6921 (N_6921,N_6418,N_6563);
xnor U6922 (N_6922,N_6229,N_6192);
or U6923 (N_6923,N_6588,N_6355);
nand U6924 (N_6924,N_6593,N_6010);
nor U6925 (N_6925,N_6158,N_6378);
xor U6926 (N_6926,N_6166,N_6052);
or U6927 (N_6927,N_6038,N_6522);
nor U6928 (N_6928,N_6402,N_6215);
and U6929 (N_6929,N_6282,N_6064);
or U6930 (N_6930,N_6027,N_6142);
or U6931 (N_6931,N_6262,N_6043);
or U6932 (N_6932,N_6037,N_6578);
and U6933 (N_6933,N_6505,N_6426);
or U6934 (N_6934,N_6400,N_6227);
and U6935 (N_6935,N_6332,N_6273);
nor U6936 (N_6936,N_6200,N_6389);
and U6937 (N_6937,N_6320,N_6410);
and U6938 (N_6938,N_6487,N_6061);
nand U6939 (N_6939,N_6035,N_6297);
nor U6940 (N_6940,N_6203,N_6522);
and U6941 (N_6941,N_6046,N_6549);
or U6942 (N_6942,N_6398,N_6254);
nand U6943 (N_6943,N_6165,N_6480);
or U6944 (N_6944,N_6337,N_6206);
and U6945 (N_6945,N_6559,N_6308);
nor U6946 (N_6946,N_6478,N_6535);
or U6947 (N_6947,N_6562,N_6345);
nor U6948 (N_6948,N_6506,N_6021);
and U6949 (N_6949,N_6475,N_6122);
or U6950 (N_6950,N_6167,N_6213);
xor U6951 (N_6951,N_6179,N_6192);
and U6952 (N_6952,N_6138,N_6166);
or U6953 (N_6953,N_6024,N_6431);
nand U6954 (N_6954,N_6320,N_6229);
or U6955 (N_6955,N_6001,N_6170);
or U6956 (N_6956,N_6538,N_6263);
nor U6957 (N_6957,N_6265,N_6355);
nor U6958 (N_6958,N_6071,N_6248);
nor U6959 (N_6959,N_6555,N_6585);
nand U6960 (N_6960,N_6353,N_6383);
nor U6961 (N_6961,N_6014,N_6506);
nand U6962 (N_6962,N_6502,N_6080);
nor U6963 (N_6963,N_6044,N_6490);
and U6964 (N_6964,N_6003,N_6478);
nand U6965 (N_6965,N_6480,N_6483);
and U6966 (N_6966,N_6337,N_6349);
or U6967 (N_6967,N_6548,N_6086);
or U6968 (N_6968,N_6034,N_6073);
nor U6969 (N_6969,N_6011,N_6236);
nand U6970 (N_6970,N_6415,N_6397);
nand U6971 (N_6971,N_6079,N_6294);
or U6972 (N_6972,N_6087,N_6080);
or U6973 (N_6973,N_6093,N_6120);
nand U6974 (N_6974,N_6268,N_6051);
or U6975 (N_6975,N_6077,N_6456);
and U6976 (N_6976,N_6202,N_6021);
or U6977 (N_6977,N_6599,N_6493);
nand U6978 (N_6978,N_6108,N_6520);
and U6979 (N_6979,N_6076,N_6410);
and U6980 (N_6980,N_6315,N_6212);
or U6981 (N_6981,N_6197,N_6598);
and U6982 (N_6982,N_6585,N_6146);
nand U6983 (N_6983,N_6047,N_6478);
or U6984 (N_6984,N_6216,N_6504);
nand U6985 (N_6985,N_6241,N_6387);
or U6986 (N_6986,N_6181,N_6527);
or U6987 (N_6987,N_6028,N_6599);
nor U6988 (N_6988,N_6376,N_6142);
or U6989 (N_6989,N_6195,N_6571);
and U6990 (N_6990,N_6226,N_6194);
and U6991 (N_6991,N_6354,N_6293);
and U6992 (N_6992,N_6324,N_6076);
nand U6993 (N_6993,N_6561,N_6567);
nand U6994 (N_6994,N_6486,N_6183);
or U6995 (N_6995,N_6077,N_6093);
and U6996 (N_6996,N_6244,N_6334);
nand U6997 (N_6997,N_6491,N_6581);
or U6998 (N_6998,N_6085,N_6253);
or U6999 (N_6999,N_6506,N_6093);
nor U7000 (N_7000,N_6355,N_6137);
xnor U7001 (N_7001,N_6504,N_6381);
nor U7002 (N_7002,N_6269,N_6433);
or U7003 (N_7003,N_6131,N_6588);
nor U7004 (N_7004,N_6293,N_6483);
or U7005 (N_7005,N_6401,N_6073);
and U7006 (N_7006,N_6544,N_6031);
and U7007 (N_7007,N_6378,N_6369);
and U7008 (N_7008,N_6147,N_6229);
nand U7009 (N_7009,N_6040,N_6489);
and U7010 (N_7010,N_6037,N_6115);
nor U7011 (N_7011,N_6161,N_6263);
nor U7012 (N_7012,N_6196,N_6162);
nand U7013 (N_7013,N_6196,N_6403);
nand U7014 (N_7014,N_6300,N_6214);
nor U7015 (N_7015,N_6039,N_6246);
nor U7016 (N_7016,N_6281,N_6067);
nor U7017 (N_7017,N_6001,N_6081);
nor U7018 (N_7018,N_6054,N_6119);
nor U7019 (N_7019,N_6476,N_6449);
and U7020 (N_7020,N_6047,N_6564);
and U7021 (N_7021,N_6243,N_6162);
nand U7022 (N_7022,N_6307,N_6464);
nand U7023 (N_7023,N_6459,N_6438);
and U7024 (N_7024,N_6476,N_6419);
nand U7025 (N_7025,N_6494,N_6589);
nand U7026 (N_7026,N_6269,N_6530);
nor U7027 (N_7027,N_6541,N_6500);
and U7028 (N_7028,N_6148,N_6323);
or U7029 (N_7029,N_6186,N_6031);
xor U7030 (N_7030,N_6008,N_6360);
nor U7031 (N_7031,N_6053,N_6387);
xor U7032 (N_7032,N_6446,N_6489);
nand U7033 (N_7033,N_6363,N_6288);
or U7034 (N_7034,N_6335,N_6065);
and U7035 (N_7035,N_6365,N_6572);
or U7036 (N_7036,N_6416,N_6288);
or U7037 (N_7037,N_6581,N_6179);
or U7038 (N_7038,N_6366,N_6386);
nor U7039 (N_7039,N_6077,N_6454);
and U7040 (N_7040,N_6445,N_6039);
xnor U7041 (N_7041,N_6561,N_6137);
or U7042 (N_7042,N_6240,N_6330);
nor U7043 (N_7043,N_6568,N_6485);
and U7044 (N_7044,N_6217,N_6399);
nand U7045 (N_7045,N_6408,N_6522);
and U7046 (N_7046,N_6332,N_6027);
or U7047 (N_7047,N_6224,N_6036);
nor U7048 (N_7048,N_6423,N_6375);
nand U7049 (N_7049,N_6426,N_6071);
and U7050 (N_7050,N_6400,N_6500);
nand U7051 (N_7051,N_6370,N_6103);
nand U7052 (N_7052,N_6065,N_6014);
or U7053 (N_7053,N_6117,N_6021);
and U7054 (N_7054,N_6495,N_6552);
and U7055 (N_7055,N_6287,N_6288);
or U7056 (N_7056,N_6043,N_6315);
nand U7057 (N_7057,N_6157,N_6541);
or U7058 (N_7058,N_6249,N_6533);
nand U7059 (N_7059,N_6474,N_6322);
xnor U7060 (N_7060,N_6138,N_6062);
or U7061 (N_7061,N_6022,N_6465);
or U7062 (N_7062,N_6294,N_6426);
and U7063 (N_7063,N_6555,N_6228);
or U7064 (N_7064,N_6137,N_6521);
nor U7065 (N_7065,N_6469,N_6153);
and U7066 (N_7066,N_6105,N_6296);
or U7067 (N_7067,N_6533,N_6299);
nor U7068 (N_7068,N_6559,N_6169);
xnor U7069 (N_7069,N_6554,N_6291);
or U7070 (N_7070,N_6598,N_6268);
nand U7071 (N_7071,N_6319,N_6102);
and U7072 (N_7072,N_6340,N_6420);
or U7073 (N_7073,N_6150,N_6448);
and U7074 (N_7074,N_6564,N_6242);
or U7075 (N_7075,N_6066,N_6254);
nor U7076 (N_7076,N_6150,N_6450);
nor U7077 (N_7077,N_6133,N_6149);
and U7078 (N_7078,N_6129,N_6485);
nor U7079 (N_7079,N_6490,N_6013);
nand U7080 (N_7080,N_6358,N_6262);
nand U7081 (N_7081,N_6267,N_6331);
nand U7082 (N_7082,N_6241,N_6092);
or U7083 (N_7083,N_6074,N_6253);
nand U7084 (N_7084,N_6557,N_6405);
or U7085 (N_7085,N_6214,N_6000);
or U7086 (N_7086,N_6368,N_6362);
nor U7087 (N_7087,N_6258,N_6237);
nand U7088 (N_7088,N_6316,N_6526);
nor U7089 (N_7089,N_6583,N_6445);
and U7090 (N_7090,N_6383,N_6107);
and U7091 (N_7091,N_6048,N_6167);
or U7092 (N_7092,N_6217,N_6471);
nand U7093 (N_7093,N_6207,N_6173);
and U7094 (N_7094,N_6590,N_6326);
nand U7095 (N_7095,N_6186,N_6493);
and U7096 (N_7096,N_6421,N_6143);
or U7097 (N_7097,N_6545,N_6030);
nand U7098 (N_7098,N_6105,N_6091);
or U7099 (N_7099,N_6359,N_6164);
nor U7100 (N_7100,N_6122,N_6204);
and U7101 (N_7101,N_6346,N_6426);
and U7102 (N_7102,N_6267,N_6217);
nor U7103 (N_7103,N_6142,N_6352);
nor U7104 (N_7104,N_6267,N_6453);
nand U7105 (N_7105,N_6123,N_6419);
or U7106 (N_7106,N_6237,N_6436);
nor U7107 (N_7107,N_6246,N_6598);
and U7108 (N_7108,N_6335,N_6492);
nand U7109 (N_7109,N_6509,N_6168);
nand U7110 (N_7110,N_6264,N_6318);
and U7111 (N_7111,N_6337,N_6550);
nor U7112 (N_7112,N_6428,N_6031);
nor U7113 (N_7113,N_6401,N_6505);
or U7114 (N_7114,N_6592,N_6014);
and U7115 (N_7115,N_6334,N_6320);
or U7116 (N_7116,N_6476,N_6111);
and U7117 (N_7117,N_6094,N_6487);
and U7118 (N_7118,N_6273,N_6275);
nor U7119 (N_7119,N_6208,N_6206);
and U7120 (N_7120,N_6212,N_6151);
nor U7121 (N_7121,N_6286,N_6005);
or U7122 (N_7122,N_6107,N_6237);
nor U7123 (N_7123,N_6272,N_6388);
nor U7124 (N_7124,N_6434,N_6586);
or U7125 (N_7125,N_6027,N_6227);
xor U7126 (N_7126,N_6144,N_6039);
nor U7127 (N_7127,N_6533,N_6280);
nand U7128 (N_7128,N_6352,N_6591);
and U7129 (N_7129,N_6350,N_6513);
nor U7130 (N_7130,N_6256,N_6454);
nor U7131 (N_7131,N_6449,N_6074);
xnor U7132 (N_7132,N_6093,N_6271);
nor U7133 (N_7133,N_6032,N_6217);
nand U7134 (N_7134,N_6376,N_6206);
nand U7135 (N_7135,N_6183,N_6360);
and U7136 (N_7136,N_6214,N_6475);
nor U7137 (N_7137,N_6180,N_6220);
nand U7138 (N_7138,N_6427,N_6263);
or U7139 (N_7139,N_6079,N_6363);
and U7140 (N_7140,N_6025,N_6251);
nand U7141 (N_7141,N_6408,N_6314);
and U7142 (N_7142,N_6084,N_6348);
nand U7143 (N_7143,N_6288,N_6140);
nor U7144 (N_7144,N_6163,N_6135);
nand U7145 (N_7145,N_6089,N_6117);
or U7146 (N_7146,N_6217,N_6578);
xnor U7147 (N_7147,N_6470,N_6330);
nand U7148 (N_7148,N_6422,N_6027);
nor U7149 (N_7149,N_6173,N_6455);
nand U7150 (N_7150,N_6492,N_6326);
or U7151 (N_7151,N_6222,N_6043);
nor U7152 (N_7152,N_6211,N_6319);
or U7153 (N_7153,N_6065,N_6040);
and U7154 (N_7154,N_6388,N_6595);
nor U7155 (N_7155,N_6481,N_6453);
or U7156 (N_7156,N_6345,N_6021);
and U7157 (N_7157,N_6579,N_6339);
or U7158 (N_7158,N_6573,N_6100);
xnor U7159 (N_7159,N_6356,N_6426);
or U7160 (N_7160,N_6314,N_6224);
nand U7161 (N_7161,N_6590,N_6129);
and U7162 (N_7162,N_6189,N_6287);
nand U7163 (N_7163,N_6404,N_6411);
and U7164 (N_7164,N_6476,N_6573);
and U7165 (N_7165,N_6410,N_6510);
or U7166 (N_7166,N_6194,N_6078);
nand U7167 (N_7167,N_6298,N_6497);
nand U7168 (N_7168,N_6239,N_6364);
nor U7169 (N_7169,N_6495,N_6037);
or U7170 (N_7170,N_6114,N_6285);
xnor U7171 (N_7171,N_6504,N_6174);
nor U7172 (N_7172,N_6504,N_6318);
or U7173 (N_7173,N_6315,N_6345);
nand U7174 (N_7174,N_6017,N_6100);
and U7175 (N_7175,N_6481,N_6308);
or U7176 (N_7176,N_6560,N_6129);
or U7177 (N_7177,N_6153,N_6371);
and U7178 (N_7178,N_6455,N_6494);
nand U7179 (N_7179,N_6496,N_6294);
or U7180 (N_7180,N_6424,N_6379);
nand U7181 (N_7181,N_6463,N_6081);
or U7182 (N_7182,N_6330,N_6581);
nand U7183 (N_7183,N_6249,N_6433);
nand U7184 (N_7184,N_6428,N_6596);
nor U7185 (N_7185,N_6419,N_6457);
and U7186 (N_7186,N_6399,N_6529);
or U7187 (N_7187,N_6352,N_6508);
and U7188 (N_7188,N_6338,N_6333);
nand U7189 (N_7189,N_6042,N_6350);
or U7190 (N_7190,N_6519,N_6564);
and U7191 (N_7191,N_6229,N_6028);
and U7192 (N_7192,N_6261,N_6142);
nand U7193 (N_7193,N_6355,N_6523);
or U7194 (N_7194,N_6221,N_6342);
nand U7195 (N_7195,N_6111,N_6003);
or U7196 (N_7196,N_6311,N_6331);
nand U7197 (N_7197,N_6556,N_6239);
and U7198 (N_7198,N_6143,N_6580);
and U7199 (N_7199,N_6511,N_6106);
and U7200 (N_7200,N_6717,N_6891);
nor U7201 (N_7201,N_7000,N_6852);
or U7202 (N_7202,N_6924,N_6793);
nor U7203 (N_7203,N_6901,N_6912);
nor U7204 (N_7204,N_6834,N_6607);
and U7205 (N_7205,N_7078,N_6678);
nor U7206 (N_7206,N_6613,N_7082);
and U7207 (N_7207,N_7074,N_7091);
or U7208 (N_7208,N_6655,N_6638);
nor U7209 (N_7209,N_6601,N_6919);
and U7210 (N_7210,N_6780,N_7127);
or U7211 (N_7211,N_7022,N_7173);
nor U7212 (N_7212,N_6832,N_6963);
and U7213 (N_7213,N_6746,N_6970);
and U7214 (N_7214,N_6624,N_6884);
or U7215 (N_7215,N_6931,N_7148);
or U7216 (N_7216,N_7062,N_6665);
nand U7217 (N_7217,N_7047,N_6606);
xnor U7218 (N_7218,N_6609,N_7165);
or U7219 (N_7219,N_7068,N_7032);
or U7220 (N_7220,N_6993,N_6979);
and U7221 (N_7221,N_7128,N_7070);
and U7222 (N_7222,N_6894,N_6913);
or U7223 (N_7223,N_7110,N_7051);
nand U7224 (N_7224,N_6889,N_7103);
and U7225 (N_7225,N_6971,N_6915);
or U7226 (N_7226,N_7066,N_6787);
nor U7227 (N_7227,N_7027,N_7015);
nand U7228 (N_7228,N_6698,N_7045);
nand U7229 (N_7229,N_6757,N_7021);
and U7230 (N_7230,N_6860,N_6959);
and U7231 (N_7231,N_6868,N_6741);
nor U7232 (N_7232,N_6699,N_6997);
and U7233 (N_7233,N_6998,N_6727);
nand U7234 (N_7234,N_6865,N_6791);
nor U7235 (N_7235,N_6898,N_6955);
nand U7236 (N_7236,N_6799,N_6822);
nor U7237 (N_7237,N_7094,N_6949);
or U7238 (N_7238,N_6694,N_7033);
nand U7239 (N_7239,N_6830,N_6795);
and U7240 (N_7240,N_6906,N_7132);
or U7241 (N_7241,N_6619,N_7176);
or U7242 (N_7242,N_6713,N_6776);
nand U7243 (N_7243,N_7156,N_6845);
nand U7244 (N_7244,N_7113,N_7063);
nand U7245 (N_7245,N_7170,N_7072);
or U7246 (N_7246,N_7149,N_7086);
xor U7247 (N_7247,N_6688,N_6841);
nor U7248 (N_7248,N_7152,N_6867);
nor U7249 (N_7249,N_6947,N_7046);
or U7250 (N_7250,N_6905,N_7126);
or U7251 (N_7251,N_7018,N_6680);
and U7252 (N_7252,N_7058,N_7161);
nor U7253 (N_7253,N_6728,N_6961);
or U7254 (N_7254,N_6662,N_6988);
nand U7255 (N_7255,N_7175,N_6895);
nand U7256 (N_7256,N_7038,N_7095);
or U7257 (N_7257,N_6668,N_6855);
nand U7258 (N_7258,N_6978,N_6771);
nand U7259 (N_7259,N_6944,N_6820);
or U7260 (N_7260,N_6805,N_6628);
nand U7261 (N_7261,N_6663,N_6985);
and U7262 (N_7262,N_6604,N_6632);
nor U7263 (N_7263,N_6740,N_6916);
or U7264 (N_7264,N_7183,N_7090);
nor U7265 (N_7265,N_6726,N_6842);
or U7266 (N_7266,N_6914,N_6785);
or U7267 (N_7267,N_6652,N_7197);
or U7268 (N_7268,N_6702,N_6853);
and U7269 (N_7269,N_6796,N_6752);
and U7270 (N_7270,N_6938,N_6811);
or U7271 (N_7271,N_6792,N_6951);
nand U7272 (N_7272,N_6801,N_6885);
and U7273 (N_7273,N_6747,N_6857);
nand U7274 (N_7274,N_7160,N_6756);
nand U7275 (N_7275,N_6870,N_6608);
and U7276 (N_7276,N_6958,N_6710);
or U7277 (N_7277,N_7042,N_6656);
and U7278 (N_7278,N_6763,N_7039);
or U7279 (N_7279,N_7092,N_7050);
or U7280 (N_7280,N_7104,N_6815);
nor U7281 (N_7281,N_6809,N_6614);
nand U7282 (N_7282,N_7168,N_6990);
nor U7283 (N_7283,N_7109,N_7006);
nor U7284 (N_7284,N_6715,N_6721);
nor U7285 (N_7285,N_6761,N_6783);
nand U7286 (N_7286,N_6966,N_6967);
and U7287 (N_7287,N_7158,N_6892);
or U7288 (N_7288,N_6847,N_6673);
and U7289 (N_7289,N_7135,N_6824);
nand U7290 (N_7290,N_7099,N_7081);
and U7291 (N_7291,N_7083,N_7191);
and U7292 (N_7292,N_6975,N_6875);
nand U7293 (N_7293,N_7107,N_7157);
and U7294 (N_7294,N_7096,N_6819);
nor U7295 (N_7295,N_6732,N_7196);
and U7296 (N_7296,N_6704,N_6769);
and U7297 (N_7297,N_7111,N_6882);
and U7298 (N_7298,N_6642,N_6786);
and U7299 (N_7299,N_7137,N_6935);
nor U7300 (N_7300,N_7116,N_6754);
nand U7301 (N_7301,N_6685,N_7134);
nand U7302 (N_7302,N_6888,N_6965);
nor U7303 (N_7303,N_7108,N_7024);
and U7304 (N_7304,N_6973,N_7112);
or U7305 (N_7305,N_6920,N_6605);
or U7306 (N_7306,N_7184,N_6735);
or U7307 (N_7307,N_6923,N_6952);
nor U7308 (N_7308,N_6765,N_7029);
nand U7309 (N_7309,N_6907,N_6705);
nor U7310 (N_7310,N_6810,N_6759);
nor U7311 (N_7311,N_6987,N_6734);
nor U7312 (N_7312,N_6880,N_6669);
nor U7313 (N_7313,N_6995,N_6616);
nand U7314 (N_7314,N_7118,N_7079);
and U7315 (N_7315,N_6731,N_6849);
nor U7316 (N_7316,N_7178,N_6829);
and U7317 (N_7317,N_6720,N_6660);
and U7318 (N_7318,N_6627,N_6730);
and U7319 (N_7319,N_6933,N_6869);
or U7320 (N_7320,N_6862,N_6804);
and U7321 (N_7321,N_7065,N_7169);
and U7322 (N_7322,N_6661,N_7187);
nor U7323 (N_7323,N_7001,N_6881);
nor U7324 (N_7324,N_7030,N_6911);
nand U7325 (N_7325,N_6758,N_6693);
and U7326 (N_7326,N_6921,N_6953);
or U7327 (N_7327,N_6784,N_6939);
nor U7328 (N_7328,N_7089,N_6802);
nor U7329 (N_7329,N_6719,N_6760);
nand U7330 (N_7330,N_6623,N_6817);
nor U7331 (N_7331,N_6788,N_7150);
nor U7332 (N_7332,N_6873,N_6942);
nand U7333 (N_7333,N_6976,N_6928);
and U7334 (N_7334,N_7023,N_7014);
nor U7335 (N_7335,N_6744,N_6789);
nor U7336 (N_7336,N_7131,N_7130);
nor U7337 (N_7337,N_6675,N_6812);
and U7338 (N_7338,N_6711,N_7177);
nor U7339 (N_7339,N_6682,N_6766);
and U7340 (N_7340,N_7106,N_6648);
nor U7341 (N_7341,N_6621,N_7025);
and U7342 (N_7342,N_7179,N_7142);
nand U7343 (N_7343,N_6737,N_6618);
and U7344 (N_7344,N_7093,N_7143);
and U7345 (N_7345,N_6634,N_6883);
and U7346 (N_7346,N_6695,N_7009);
nand U7347 (N_7347,N_6743,N_6779);
and U7348 (N_7348,N_6781,N_6777);
and U7349 (N_7349,N_6863,N_6982);
nor U7350 (N_7350,N_6999,N_6681);
nor U7351 (N_7351,N_7010,N_7028);
nand U7352 (N_7352,N_6918,N_6940);
nand U7353 (N_7353,N_6631,N_6878);
and U7354 (N_7354,N_6818,N_6709);
nor U7355 (N_7355,N_6635,N_6856);
and U7356 (N_7356,N_6934,N_6962);
nand U7357 (N_7357,N_6986,N_7192);
or U7358 (N_7358,N_7026,N_7139);
nor U7359 (N_7359,N_6981,N_6773);
nand U7360 (N_7360,N_6687,N_7147);
or U7361 (N_7361,N_6836,N_6644);
or U7362 (N_7362,N_7174,N_6808);
and U7363 (N_7363,N_6649,N_6877);
nor U7364 (N_7364,N_7097,N_7171);
nor U7365 (N_7365,N_7190,N_7146);
and U7366 (N_7366,N_7012,N_6859);
and U7367 (N_7367,N_6844,N_7061);
nor U7368 (N_7368,N_6750,N_6922);
nand U7369 (N_7369,N_6725,N_6722);
and U7370 (N_7370,N_6831,N_7044);
and U7371 (N_7371,N_6840,N_6748);
or U7372 (N_7372,N_7073,N_6828);
and U7373 (N_7373,N_6996,N_7145);
nand U7374 (N_7374,N_6697,N_6886);
nor U7375 (N_7375,N_7057,N_7181);
nor U7376 (N_7376,N_6909,N_7049);
nand U7377 (N_7377,N_7060,N_7163);
nor U7378 (N_7378,N_6816,N_6866);
nor U7379 (N_7379,N_6992,N_7071);
or U7380 (N_7380,N_6691,N_6643);
nor U7381 (N_7381,N_6778,N_6653);
and U7382 (N_7382,N_6689,N_7098);
and U7383 (N_7383,N_7136,N_6647);
and U7384 (N_7384,N_6637,N_6936);
nand U7385 (N_7385,N_6893,N_6874);
or U7386 (N_7386,N_7080,N_7055);
nor U7387 (N_7387,N_6739,N_6639);
and U7388 (N_7388,N_6879,N_6658);
nor U7389 (N_7389,N_6972,N_7188);
nor U7390 (N_7390,N_6736,N_7041);
nor U7391 (N_7391,N_7121,N_6708);
nand U7392 (N_7392,N_6626,N_6904);
nor U7393 (N_7393,N_6843,N_6686);
and U7394 (N_7394,N_6800,N_6943);
nand U7395 (N_7395,N_7043,N_6733);
or U7396 (N_7396,N_6782,N_6968);
nor U7397 (N_7397,N_6983,N_6646);
or U7398 (N_7398,N_6900,N_7129);
and U7399 (N_7399,N_6629,N_6602);
and U7400 (N_7400,N_7151,N_6823);
and U7401 (N_7401,N_6679,N_6672);
nand U7402 (N_7402,N_6960,N_7013);
and U7403 (N_7403,N_7198,N_7155);
and U7404 (N_7404,N_6927,N_6716);
or U7405 (N_7405,N_7002,N_6664);
and U7406 (N_7406,N_6600,N_7194);
and U7407 (N_7407,N_7115,N_6723);
nor U7408 (N_7408,N_6657,N_7138);
or U7409 (N_7409,N_7004,N_7017);
or U7410 (N_7410,N_7164,N_7064);
or U7411 (N_7411,N_6764,N_7124);
nand U7412 (N_7412,N_7053,N_7084);
nand U7413 (N_7413,N_6814,N_6745);
nand U7414 (N_7414,N_6692,N_6917);
and U7415 (N_7415,N_7154,N_6837);
and U7416 (N_7416,N_6899,N_6807);
nand U7417 (N_7417,N_6871,N_6729);
nand U7418 (N_7418,N_6848,N_7031);
nor U7419 (N_7419,N_6667,N_6714);
nand U7420 (N_7420,N_6790,N_6615);
nand U7421 (N_7421,N_6755,N_6794);
and U7422 (N_7422,N_6864,N_7189);
and U7423 (N_7423,N_6851,N_6703);
and U7424 (N_7424,N_6676,N_6775);
or U7425 (N_7425,N_6826,N_6645);
nor U7426 (N_7426,N_7166,N_7007);
nor U7427 (N_7427,N_7069,N_6650);
nand U7428 (N_7428,N_7185,N_7122);
or U7429 (N_7429,N_6762,N_6742);
nor U7430 (N_7430,N_7167,N_6611);
nor U7431 (N_7431,N_7114,N_6854);
or U7432 (N_7432,N_6897,N_6620);
and U7433 (N_7433,N_6994,N_7153);
or U7434 (N_7434,N_7162,N_6671);
nor U7435 (N_7435,N_7100,N_7008);
and U7436 (N_7436,N_6633,N_6835);
nor U7437 (N_7437,N_6945,N_6718);
and U7438 (N_7438,N_6930,N_7172);
or U7439 (N_7439,N_7193,N_6838);
and U7440 (N_7440,N_6896,N_7067);
nor U7441 (N_7441,N_6980,N_7052);
or U7442 (N_7442,N_6872,N_7182);
or U7443 (N_7443,N_7159,N_6846);
nand U7444 (N_7444,N_6630,N_6666);
nand U7445 (N_7445,N_6767,N_7101);
or U7446 (N_7446,N_6701,N_7133);
nor U7447 (N_7447,N_6707,N_6946);
nor U7448 (N_7448,N_6926,N_6768);
and U7449 (N_7449,N_6984,N_6850);
and U7450 (N_7450,N_6902,N_6977);
nor U7451 (N_7451,N_7059,N_6948);
nand U7452 (N_7452,N_7036,N_6929);
or U7453 (N_7453,N_6612,N_7085);
or U7454 (N_7454,N_6603,N_6887);
nand U7455 (N_7455,N_6770,N_6622);
or U7456 (N_7456,N_6925,N_7034);
and U7457 (N_7457,N_6683,N_6640);
or U7458 (N_7458,N_7056,N_7048);
nand U7459 (N_7459,N_6827,N_6833);
or U7460 (N_7460,N_6641,N_6651);
or U7461 (N_7461,N_6706,N_6890);
and U7462 (N_7462,N_6974,N_7186);
and U7463 (N_7463,N_6956,N_6903);
or U7464 (N_7464,N_7125,N_7102);
nand U7465 (N_7465,N_6751,N_7037);
or U7466 (N_7466,N_7117,N_7105);
or U7467 (N_7467,N_7020,N_6774);
nor U7468 (N_7468,N_6659,N_6749);
nand U7469 (N_7469,N_7141,N_7119);
nand U7470 (N_7470,N_6696,N_7016);
nand U7471 (N_7471,N_6636,N_7120);
or U7472 (N_7472,N_6684,N_6738);
and U7473 (N_7473,N_6724,N_7144);
and U7474 (N_7474,N_6969,N_7180);
and U7475 (N_7475,N_6910,N_7019);
nor U7476 (N_7476,N_6803,N_6813);
nand U7477 (N_7477,N_6797,N_6989);
nor U7478 (N_7478,N_6941,N_6839);
nand U7479 (N_7479,N_7199,N_6674);
or U7480 (N_7480,N_7123,N_7035);
nor U7481 (N_7481,N_7195,N_7077);
nand U7482 (N_7482,N_6677,N_7005);
nand U7483 (N_7483,N_6908,N_6821);
or U7484 (N_7484,N_6806,N_7087);
and U7485 (N_7485,N_6954,N_6876);
nand U7486 (N_7486,N_6858,N_6772);
nand U7487 (N_7487,N_6625,N_7076);
or U7488 (N_7488,N_6753,N_6690);
or U7489 (N_7489,N_6617,N_6670);
nand U7490 (N_7490,N_6991,N_7140);
or U7491 (N_7491,N_6825,N_6798);
and U7492 (N_7492,N_7088,N_6700);
or U7493 (N_7493,N_7040,N_6610);
or U7494 (N_7494,N_6950,N_6932);
or U7495 (N_7495,N_6861,N_7075);
nor U7496 (N_7496,N_6957,N_6654);
or U7497 (N_7497,N_7011,N_6964);
or U7498 (N_7498,N_7054,N_6937);
and U7499 (N_7499,N_7003,N_6712);
nand U7500 (N_7500,N_6780,N_6718);
nand U7501 (N_7501,N_7064,N_6799);
and U7502 (N_7502,N_6718,N_7120);
nor U7503 (N_7503,N_7012,N_6855);
nand U7504 (N_7504,N_6917,N_7037);
nand U7505 (N_7505,N_6934,N_6643);
nand U7506 (N_7506,N_7073,N_6921);
or U7507 (N_7507,N_6743,N_7123);
nand U7508 (N_7508,N_7055,N_7103);
nand U7509 (N_7509,N_6711,N_6722);
nor U7510 (N_7510,N_6880,N_7195);
and U7511 (N_7511,N_6911,N_7194);
and U7512 (N_7512,N_7098,N_7020);
nand U7513 (N_7513,N_6704,N_6657);
nor U7514 (N_7514,N_7113,N_6854);
and U7515 (N_7515,N_6628,N_6895);
xnor U7516 (N_7516,N_6621,N_6627);
and U7517 (N_7517,N_7186,N_7169);
or U7518 (N_7518,N_6967,N_6808);
nor U7519 (N_7519,N_6734,N_7114);
nor U7520 (N_7520,N_6643,N_6995);
nand U7521 (N_7521,N_6699,N_6869);
or U7522 (N_7522,N_6678,N_6784);
nand U7523 (N_7523,N_6964,N_6902);
and U7524 (N_7524,N_6894,N_6884);
nand U7525 (N_7525,N_6829,N_6940);
or U7526 (N_7526,N_6624,N_7112);
nor U7527 (N_7527,N_7016,N_6763);
xnor U7528 (N_7528,N_7135,N_6747);
nand U7529 (N_7529,N_6684,N_7148);
xor U7530 (N_7530,N_6918,N_6605);
nand U7531 (N_7531,N_6891,N_7096);
nor U7532 (N_7532,N_6672,N_6898);
or U7533 (N_7533,N_6723,N_6650);
or U7534 (N_7534,N_6948,N_6658);
nor U7535 (N_7535,N_6991,N_7059);
and U7536 (N_7536,N_6764,N_6899);
nor U7537 (N_7537,N_6759,N_6712);
nor U7538 (N_7538,N_6770,N_7041);
and U7539 (N_7539,N_6641,N_6763);
nor U7540 (N_7540,N_6725,N_6842);
nand U7541 (N_7541,N_7059,N_6815);
nand U7542 (N_7542,N_7147,N_7105);
nor U7543 (N_7543,N_7165,N_6607);
nor U7544 (N_7544,N_6895,N_7083);
and U7545 (N_7545,N_6981,N_6646);
nor U7546 (N_7546,N_6913,N_6835);
nor U7547 (N_7547,N_6649,N_7176);
nor U7548 (N_7548,N_6696,N_6875);
or U7549 (N_7549,N_7187,N_6693);
nor U7550 (N_7550,N_6914,N_6912);
nand U7551 (N_7551,N_6937,N_6965);
and U7552 (N_7552,N_6761,N_6653);
and U7553 (N_7553,N_6682,N_6903);
or U7554 (N_7554,N_6991,N_6960);
and U7555 (N_7555,N_6912,N_6850);
nor U7556 (N_7556,N_7002,N_6650);
and U7557 (N_7557,N_6969,N_7120);
nand U7558 (N_7558,N_6659,N_6806);
and U7559 (N_7559,N_6764,N_6801);
nor U7560 (N_7560,N_6909,N_6617);
nor U7561 (N_7561,N_6958,N_6650);
nand U7562 (N_7562,N_7197,N_6933);
nor U7563 (N_7563,N_6772,N_6916);
nor U7564 (N_7564,N_6889,N_6671);
xor U7565 (N_7565,N_6958,N_7166);
nand U7566 (N_7566,N_6700,N_6790);
and U7567 (N_7567,N_6690,N_7097);
nor U7568 (N_7568,N_6665,N_6767);
nor U7569 (N_7569,N_6869,N_6792);
nand U7570 (N_7570,N_7031,N_6931);
xnor U7571 (N_7571,N_6994,N_6794);
nor U7572 (N_7572,N_6951,N_6677);
nand U7573 (N_7573,N_7057,N_7186);
nand U7574 (N_7574,N_7164,N_6854);
nand U7575 (N_7575,N_6713,N_6707);
or U7576 (N_7576,N_7054,N_6897);
nor U7577 (N_7577,N_7113,N_7056);
or U7578 (N_7578,N_7094,N_6787);
or U7579 (N_7579,N_7159,N_6814);
xor U7580 (N_7580,N_7088,N_7081);
and U7581 (N_7581,N_6791,N_6904);
or U7582 (N_7582,N_6873,N_6754);
nand U7583 (N_7583,N_6730,N_6968);
nand U7584 (N_7584,N_7146,N_6794);
nor U7585 (N_7585,N_6796,N_6669);
nor U7586 (N_7586,N_6959,N_6620);
nor U7587 (N_7587,N_6953,N_6717);
or U7588 (N_7588,N_7152,N_6962);
nor U7589 (N_7589,N_6955,N_6763);
and U7590 (N_7590,N_6935,N_6956);
nand U7591 (N_7591,N_6662,N_6786);
and U7592 (N_7592,N_6959,N_6603);
or U7593 (N_7593,N_7058,N_6913);
nand U7594 (N_7594,N_6690,N_6966);
xor U7595 (N_7595,N_6693,N_6879);
nand U7596 (N_7596,N_7158,N_6774);
nor U7597 (N_7597,N_6878,N_6802);
or U7598 (N_7598,N_7141,N_6601);
nand U7599 (N_7599,N_7184,N_6612);
and U7600 (N_7600,N_7017,N_7155);
nand U7601 (N_7601,N_6736,N_6761);
and U7602 (N_7602,N_6861,N_6747);
nand U7603 (N_7603,N_7135,N_6806);
nor U7604 (N_7604,N_6610,N_6763);
or U7605 (N_7605,N_6668,N_6717);
or U7606 (N_7606,N_6725,N_7030);
and U7607 (N_7607,N_6809,N_7143);
or U7608 (N_7608,N_6813,N_7048);
nor U7609 (N_7609,N_7110,N_6970);
and U7610 (N_7610,N_7016,N_6954);
nand U7611 (N_7611,N_6775,N_7055);
or U7612 (N_7612,N_6786,N_7184);
and U7613 (N_7613,N_6705,N_6629);
nand U7614 (N_7614,N_6620,N_6860);
xor U7615 (N_7615,N_6718,N_7042);
or U7616 (N_7616,N_7119,N_6671);
and U7617 (N_7617,N_6651,N_7171);
and U7618 (N_7618,N_6827,N_6863);
nand U7619 (N_7619,N_6838,N_6984);
or U7620 (N_7620,N_6773,N_7057);
and U7621 (N_7621,N_6753,N_6749);
nand U7622 (N_7622,N_6843,N_6800);
or U7623 (N_7623,N_7164,N_6769);
and U7624 (N_7624,N_6875,N_6775);
xnor U7625 (N_7625,N_7038,N_7013);
or U7626 (N_7626,N_6892,N_7178);
and U7627 (N_7627,N_6944,N_6776);
nor U7628 (N_7628,N_7026,N_6708);
or U7629 (N_7629,N_7199,N_7086);
or U7630 (N_7630,N_7055,N_6642);
nor U7631 (N_7631,N_7156,N_6984);
or U7632 (N_7632,N_6845,N_6716);
nand U7633 (N_7633,N_7044,N_7176);
nand U7634 (N_7634,N_7185,N_6947);
or U7635 (N_7635,N_7125,N_6994);
or U7636 (N_7636,N_7050,N_7033);
or U7637 (N_7637,N_6941,N_6715);
nand U7638 (N_7638,N_7041,N_6873);
nor U7639 (N_7639,N_6914,N_6955);
and U7640 (N_7640,N_6606,N_6849);
nand U7641 (N_7641,N_6961,N_7105);
nand U7642 (N_7642,N_6779,N_6854);
nand U7643 (N_7643,N_6806,N_7192);
and U7644 (N_7644,N_7140,N_7112);
nand U7645 (N_7645,N_6607,N_6643);
nor U7646 (N_7646,N_6920,N_6908);
nor U7647 (N_7647,N_6961,N_6705);
or U7648 (N_7648,N_6611,N_6803);
or U7649 (N_7649,N_6602,N_6971);
and U7650 (N_7650,N_6989,N_6652);
nand U7651 (N_7651,N_6616,N_6979);
or U7652 (N_7652,N_6677,N_6856);
nand U7653 (N_7653,N_6814,N_6639);
nand U7654 (N_7654,N_6940,N_6903);
or U7655 (N_7655,N_6984,N_7021);
or U7656 (N_7656,N_6750,N_7179);
or U7657 (N_7657,N_6629,N_6667);
or U7658 (N_7658,N_6914,N_6918);
nor U7659 (N_7659,N_6778,N_7113);
and U7660 (N_7660,N_7067,N_6823);
or U7661 (N_7661,N_6795,N_6826);
and U7662 (N_7662,N_7044,N_6753);
nor U7663 (N_7663,N_6898,N_7145);
nor U7664 (N_7664,N_6709,N_6632);
xnor U7665 (N_7665,N_6706,N_7037);
nand U7666 (N_7666,N_7146,N_6631);
and U7667 (N_7667,N_6710,N_6982);
nor U7668 (N_7668,N_7053,N_6968);
nand U7669 (N_7669,N_6820,N_6830);
and U7670 (N_7670,N_6829,N_6966);
or U7671 (N_7671,N_6620,N_7111);
xor U7672 (N_7672,N_6888,N_6915);
or U7673 (N_7673,N_7157,N_6718);
or U7674 (N_7674,N_6784,N_6801);
or U7675 (N_7675,N_6826,N_6955);
nand U7676 (N_7676,N_7039,N_7170);
or U7677 (N_7677,N_7179,N_6934);
nand U7678 (N_7678,N_6946,N_6635);
nand U7679 (N_7679,N_6629,N_6604);
or U7680 (N_7680,N_7028,N_7122);
or U7681 (N_7681,N_6668,N_6983);
nand U7682 (N_7682,N_6656,N_6824);
nor U7683 (N_7683,N_7137,N_6985);
or U7684 (N_7684,N_6788,N_7170);
nand U7685 (N_7685,N_6914,N_7182);
xor U7686 (N_7686,N_6824,N_6950);
nor U7687 (N_7687,N_6948,N_7187);
and U7688 (N_7688,N_7047,N_6890);
nand U7689 (N_7689,N_6899,N_6886);
and U7690 (N_7690,N_6860,N_6744);
or U7691 (N_7691,N_6709,N_6919);
nor U7692 (N_7692,N_6698,N_6804);
or U7693 (N_7693,N_7113,N_7049);
nand U7694 (N_7694,N_7187,N_7122);
and U7695 (N_7695,N_7183,N_7038);
nor U7696 (N_7696,N_6766,N_7148);
nor U7697 (N_7697,N_7194,N_6839);
nor U7698 (N_7698,N_6665,N_7100);
nand U7699 (N_7699,N_6919,N_6791);
nand U7700 (N_7700,N_6801,N_6660);
or U7701 (N_7701,N_6912,N_7115);
xnor U7702 (N_7702,N_7079,N_6862);
or U7703 (N_7703,N_7013,N_6973);
nand U7704 (N_7704,N_6615,N_6826);
and U7705 (N_7705,N_6716,N_6762);
and U7706 (N_7706,N_6639,N_6966);
nor U7707 (N_7707,N_7033,N_7155);
and U7708 (N_7708,N_7066,N_7164);
nand U7709 (N_7709,N_7195,N_6916);
and U7710 (N_7710,N_6836,N_6982);
and U7711 (N_7711,N_6996,N_6736);
nand U7712 (N_7712,N_6972,N_7109);
nand U7713 (N_7713,N_6695,N_7162);
and U7714 (N_7714,N_7136,N_7132);
nor U7715 (N_7715,N_6760,N_6958);
or U7716 (N_7716,N_7025,N_6803);
nor U7717 (N_7717,N_6817,N_6861);
nand U7718 (N_7718,N_6790,N_6657);
nor U7719 (N_7719,N_7158,N_7169);
nand U7720 (N_7720,N_7080,N_7039);
and U7721 (N_7721,N_6802,N_7175);
nand U7722 (N_7722,N_6757,N_7073);
and U7723 (N_7723,N_6942,N_6836);
or U7724 (N_7724,N_6963,N_7182);
nor U7725 (N_7725,N_6651,N_6871);
and U7726 (N_7726,N_7144,N_6919);
nand U7727 (N_7727,N_7051,N_6627);
nor U7728 (N_7728,N_6789,N_6962);
or U7729 (N_7729,N_6642,N_6865);
and U7730 (N_7730,N_7146,N_6727);
nand U7731 (N_7731,N_7010,N_6862);
nor U7732 (N_7732,N_7026,N_6685);
and U7733 (N_7733,N_6665,N_7051);
nand U7734 (N_7734,N_6604,N_7011);
nand U7735 (N_7735,N_6808,N_7175);
nand U7736 (N_7736,N_6847,N_6751);
and U7737 (N_7737,N_6976,N_6734);
or U7738 (N_7738,N_7115,N_6815);
and U7739 (N_7739,N_7113,N_6878);
nor U7740 (N_7740,N_6895,N_7019);
or U7741 (N_7741,N_6895,N_7118);
or U7742 (N_7742,N_6827,N_7051);
nor U7743 (N_7743,N_7023,N_7005);
and U7744 (N_7744,N_6812,N_7095);
nor U7745 (N_7745,N_6860,N_6642);
and U7746 (N_7746,N_7008,N_6855);
nor U7747 (N_7747,N_6689,N_6627);
nor U7748 (N_7748,N_6723,N_7072);
nand U7749 (N_7749,N_6676,N_6649);
nand U7750 (N_7750,N_6915,N_6655);
or U7751 (N_7751,N_6874,N_7145);
and U7752 (N_7752,N_6850,N_6860);
nand U7753 (N_7753,N_7171,N_6803);
nor U7754 (N_7754,N_6823,N_6623);
or U7755 (N_7755,N_6766,N_7042);
nand U7756 (N_7756,N_7056,N_6954);
nand U7757 (N_7757,N_6774,N_6967);
nor U7758 (N_7758,N_6608,N_6718);
nand U7759 (N_7759,N_6676,N_7174);
nand U7760 (N_7760,N_6823,N_7136);
nand U7761 (N_7761,N_7149,N_6729);
and U7762 (N_7762,N_6965,N_6913);
and U7763 (N_7763,N_7034,N_7046);
or U7764 (N_7764,N_6937,N_6980);
and U7765 (N_7765,N_6856,N_6789);
nor U7766 (N_7766,N_6903,N_7118);
nor U7767 (N_7767,N_6659,N_7156);
and U7768 (N_7768,N_7162,N_6915);
nor U7769 (N_7769,N_6886,N_7048);
and U7770 (N_7770,N_6644,N_7098);
and U7771 (N_7771,N_7005,N_6895);
and U7772 (N_7772,N_6682,N_6723);
nor U7773 (N_7773,N_6972,N_6663);
or U7774 (N_7774,N_6881,N_6935);
nor U7775 (N_7775,N_6684,N_7093);
or U7776 (N_7776,N_7198,N_7143);
and U7777 (N_7777,N_7085,N_6668);
and U7778 (N_7778,N_7082,N_6881);
nand U7779 (N_7779,N_6942,N_6868);
or U7780 (N_7780,N_7111,N_6821);
nand U7781 (N_7781,N_6935,N_7128);
and U7782 (N_7782,N_6794,N_7157);
or U7783 (N_7783,N_6982,N_7033);
nand U7784 (N_7784,N_6813,N_7056);
nor U7785 (N_7785,N_6618,N_7157);
nor U7786 (N_7786,N_7107,N_6655);
and U7787 (N_7787,N_6828,N_6796);
and U7788 (N_7788,N_6655,N_7069);
nor U7789 (N_7789,N_6644,N_6940);
nand U7790 (N_7790,N_7033,N_7188);
nand U7791 (N_7791,N_6725,N_6644);
and U7792 (N_7792,N_7037,N_6989);
or U7793 (N_7793,N_6921,N_6773);
and U7794 (N_7794,N_6987,N_6858);
or U7795 (N_7795,N_7187,N_7072);
nor U7796 (N_7796,N_7199,N_6755);
nor U7797 (N_7797,N_7132,N_6869);
or U7798 (N_7798,N_6689,N_7062);
nor U7799 (N_7799,N_7120,N_6847);
nor U7800 (N_7800,N_7259,N_7201);
and U7801 (N_7801,N_7791,N_7226);
or U7802 (N_7802,N_7422,N_7405);
nand U7803 (N_7803,N_7735,N_7691);
or U7804 (N_7804,N_7440,N_7714);
and U7805 (N_7805,N_7231,N_7519);
or U7806 (N_7806,N_7426,N_7581);
nand U7807 (N_7807,N_7718,N_7565);
nor U7808 (N_7808,N_7493,N_7477);
nand U7809 (N_7809,N_7710,N_7577);
or U7810 (N_7810,N_7391,N_7766);
nand U7811 (N_7811,N_7678,N_7389);
or U7812 (N_7812,N_7212,N_7392);
nand U7813 (N_7813,N_7550,N_7795);
and U7814 (N_7814,N_7689,N_7309);
nor U7815 (N_7815,N_7723,N_7421);
or U7816 (N_7816,N_7758,N_7643);
nand U7817 (N_7817,N_7525,N_7749);
nand U7818 (N_7818,N_7645,N_7637);
or U7819 (N_7819,N_7311,N_7594);
nor U7820 (N_7820,N_7402,N_7656);
and U7821 (N_7821,N_7485,N_7273);
xnor U7822 (N_7822,N_7649,N_7324);
nor U7823 (N_7823,N_7788,N_7607);
or U7824 (N_7824,N_7303,N_7377);
and U7825 (N_7825,N_7692,N_7432);
nand U7826 (N_7826,N_7455,N_7228);
or U7827 (N_7827,N_7403,N_7564);
or U7828 (N_7828,N_7598,N_7599);
xor U7829 (N_7829,N_7468,N_7603);
and U7830 (N_7830,N_7543,N_7734);
nor U7831 (N_7831,N_7237,N_7667);
nor U7832 (N_7832,N_7478,N_7457);
nor U7833 (N_7833,N_7224,N_7773);
nand U7834 (N_7834,N_7664,N_7410);
or U7835 (N_7835,N_7339,N_7680);
nand U7836 (N_7836,N_7573,N_7359);
and U7837 (N_7837,N_7386,N_7220);
xnor U7838 (N_7838,N_7558,N_7612);
and U7839 (N_7839,N_7695,N_7699);
or U7840 (N_7840,N_7225,N_7778);
and U7841 (N_7841,N_7537,N_7469);
nor U7842 (N_7842,N_7286,N_7247);
or U7843 (N_7843,N_7401,N_7299);
nor U7844 (N_7844,N_7474,N_7613);
or U7845 (N_7845,N_7282,N_7772);
and U7846 (N_7846,N_7601,N_7650);
nor U7847 (N_7847,N_7738,N_7344);
and U7848 (N_7848,N_7527,N_7685);
or U7849 (N_7849,N_7730,N_7345);
and U7850 (N_7850,N_7502,N_7798);
and U7851 (N_7851,N_7541,N_7644);
or U7852 (N_7852,N_7743,N_7246);
or U7853 (N_7853,N_7317,N_7314);
or U7854 (N_7854,N_7713,N_7399);
nor U7855 (N_7855,N_7308,N_7358);
nand U7856 (N_7856,N_7780,N_7707);
and U7857 (N_7857,N_7559,N_7676);
and U7858 (N_7858,N_7630,N_7400);
xor U7859 (N_7859,N_7362,N_7239);
nand U7860 (N_7860,N_7210,N_7529);
or U7861 (N_7861,N_7510,N_7238);
nor U7862 (N_7862,N_7322,N_7412);
nor U7863 (N_7863,N_7762,N_7554);
xor U7864 (N_7864,N_7648,N_7204);
xnor U7865 (N_7865,N_7496,N_7736);
and U7866 (N_7866,N_7626,N_7448);
xnor U7867 (N_7867,N_7538,N_7351);
nor U7868 (N_7868,N_7215,N_7267);
and U7869 (N_7869,N_7655,N_7625);
nand U7870 (N_7870,N_7750,N_7495);
or U7871 (N_7871,N_7281,N_7356);
nor U7872 (N_7872,N_7438,N_7371);
and U7873 (N_7873,N_7652,N_7756);
or U7874 (N_7874,N_7770,N_7727);
or U7875 (N_7875,N_7482,N_7205);
and U7876 (N_7876,N_7361,N_7489);
or U7877 (N_7877,N_7294,N_7765);
and U7878 (N_7878,N_7546,N_7213);
nor U7879 (N_7879,N_7669,N_7506);
and U7880 (N_7880,N_7694,N_7511);
nand U7881 (N_7881,N_7753,N_7681);
nand U7882 (N_7882,N_7700,N_7744);
and U7883 (N_7883,N_7264,N_7670);
or U7884 (N_7884,N_7256,N_7471);
or U7885 (N_7885,N_7235,N_7290);
nor U7886 (N_7886,N_7447,N_7556);
or U7887 (N_7887,N_7557,N_7793);
nor U7888 (N_7888,N_7445,N_7549);
and U7889 (N_7889,N_7221,N_7217);
nand U7890 (N_7890,N_7370,N_7323);
and U7891 (N_7891,N_7512,N_7236);
and U7892 (N_7892,N_7250,N_7679);
nor U7893 (N_7893,N_7674,N_7590);
and U7894 (N_7894,N_7328,N_7330);
and U7895 (N_7895,N_7631,N_7767);
nor U7896 (N_7896,N_7384,N_7715);
nor U7897 (N_7897,N_7397,N_7492);
and U7898 (N_7898,N_7407,N_7484);
nor U7899 (N_7899,N_7796,N_7642);
nor U7900 (N_7900,N_7301,N_7435);
nand U7901 (N_7901,N_7582,N_7223);
and U7902 (N_7902,N_7575,N_7252);
nand U7903 (N_7903,N_7249,N_7320);
and U7904 (N_7904,N_7771,N_7731);
or U7905 (N_7905,N_7242,N_7305);
nor U7906 (N_7906,N_7646,N_7721);
nor U7907 (N_7907,N_7526,N_7385);
nor U7908 (N_7908,N_7499,N_7441);
or U7909 (N_7909,N_7464,N_7604);
nor U7910 (N_7910,N_7367,N_7618);
and U7911 (N_7911,N_7516,N_7373);
and U7912 (N_7912,N_7443,N_7675);
nand U7913 (N_7913,N_7243,N_7327);
xor U7914 (N_7914,N_7234,N_7697);
and U7915 (N_7915,N_7792,N_7374);
or U7916 (N_7916,N_7764,N_7504);
nand U7917 (N_7917,N_7218,N_7528);
or U7918 (N_7918,N_7611,N_7761);
and U7919 (N_7919,N_7254,N_7449);
or U7920 (N_7920,N_7433,N_7404);
and U7921 (N_7921,N_7206,N_7790);
or U7922 (N_7922,N_7544,N_7661);
nor U7923 (N_7923,N_7390,N_7561);
nor U7924 (N_7924,N_7548,N_7253);
and U7925 (N_7925,N_7708,N_7262);
nand U7926 (N_7926,N_7354,N_7589);
nor U7927 (N_7927,N_7462,N_7276);
nand U7928 (N_7928,N_7673,N_7291);
nand U7929 (N_7929,N_7737,N_7310);
and U7930 (N_7930,N_7423,N_7270);
nor U7931 (N_7931,N_7726,N_7783);
or U7932 (N_7932,N_7619,N_7568);
nand U7933 (N_7933,N_7536,N_7337);
or U7934 (N_7934,N_7346,N_7360);
and U7935 (N_7935,N_7746,N_7797);
nor U7936 (N_7936,N_7318,N_7313);
and U7937 (N_7937,N_7470,N_7636);
or U7938 (N_7938,N_7417,N_7515);
and U7939 (N_7939,N_7364,N_7307);
or U7940 (N_7940,N_7439,N_7409);
nand U7941 (N_7941,N_7216,N_7785);
nand U7942 (N_7942,N_7241,N_7583);
or U7943 (N_7943,N_7245,N_7271);
and U7944 (N_7944,N_7641,N_7263);
xor U7945 (N_7945,N_7269,N_7261);
and U7946 (N_7946,N_7752,N_7570);
nor U7947 (N_7947,N_7520,N_7639);
or U7948 (N_7948,N_7704,N_7660);
and U7949 (N_7949,N_7289,N_7497);
and U7950 (N_7950,N_7552,N_7450);
nor U7951 (N_7951,N_7709,N_7272);
nor U7952 (N_7952,N_7382,N_7574);
or U7953 (N_7953,N_7321,N_7295);
nand U7954 (N_7954,N_7739,N_7705);
and U7955 (N_7955,N_7296,N_7712);
or U7956 (N_7956,N_7429,N_7782);
nor U7957 (N_7957,N_7733,N_7326);
or U7958 (N_7958,N_7420,N_7789);
nand U7959 (N_7959,N_7534,N_7300);
and U7960 (N_7960,N_7352,N_7616);
nor U7961 (N_7961,N_7632,N_7488);
nand U7962 (N_7962,N_7306,N_7454);
or U7963 (N_7963,N_7283,N_7682);
nand U7964 (N_7964,N_7562,N_7722);
nand U7965 (N_7965,N_7640,N_7465);
or U7966 (N_7966,N_7312,N_7298);
and U7967 (N_7967,N_7463,N_7334);
and U7968 (N_7968,N_7395,N_7486);
and U7969 (N_7969,N_7248,N_7227);
and U7970 (N_7970,N_7702,N_7200);
nor U7971 (N_7971,N_7600,N_7687);
nand U7972 (N_7972,N_7503,N_7285);
nand U7973 (N_7973,N_7266,N_7341);
and U7974 (N_7974,N_7586,N_7686);
nand U7975 (N_7975,N_7533,N_7617);
nand U7976 (N_7976,N_7763,N_7287);
nand U7977 (N_7977,N_7621,N_7532);
nand U7978 (N_7978,N_7693,N_7366);
nor U7979 (N_7979,N_7605,N_7343);
nand U7980 (N_7980,N_7591,N_7703);
and U7981 (N_7981,N_7319,N_7268);
and U7982 (N_7982,N_7376,N_7514);
nand U7983 (N_7983,N_7501,N_7779);
nor U7984 (N_7984,N_7665,N_7348);
nand U7985 (N_7985,N_7336,N_7509);
nor U7986 (N_7986,N_7466,N_7428);
nor U7987 (N_7987,N_7535,N_7381);
and U7988 (N_7988,N_7755,N_7545);
and U7989 (N_7989,N_7325,N_7424);
and U7990 (N_7990,N_7375,N_7593);
xnor U7991 (N_7991,N_7458,N_7280);
nor U7992 (N_7992,N_7431,N_7659);
or U7993 (N_7993,N_7203,N_7350);
or U7994 (N_7994,N_7698,N_7732);
nand U7995 (N_7995,N_7569,N_7467);
nor U7996 (N_7996,N_7585,N_7316);
nor U7997 (N_7997,N_7209,N_7690);
nand U7998 (N_7998,N_7329,N_7208);
nor U7999 (N_7999,N_7518,N_7513);
nand U8000 (N_8000,N_7668,N_7427);
nor U8001 (N_8001,N_7768,N_7658);
or U8002 (N_8002,N_7398,N_7393);
nor U8003 (N_8003,N_7553,N_7233);
nand U8004 (N_8004,N_7717,N_7777);
or U8005 (N_8005,N_7774,N_7288);
or U8006 (N_8006,N_7741,N_7523);
and U8007 (N_8007,N_7629,N_7340);
nor U8008 (N_8008,N_7436,N_7335);
nand U8009 (N_8009,N_7539,N_7684);
nand U8010 (N_8010,N_7222,N_7365);
and U8011 (N_8011,N_7666,N_7425);
and U8012 (N_8012,N_7284,N_7662);
and U8013 (N_8013,N_7606,N_7292);
nor U8014 (N_8014,N_7711,N_7623);
nand U8015 (N_8015,N_7483,N_7657);
nand U8016 (N_8016,N_7794,N_7475);
or U8017 (N_8017,N_7608,N_7784);
and U8018 (N_8018,N_7754,N_7522);
or U8019 (N_8019,N_7653,N_7635);
nand U8020 (N_8020,N_7595,N_7274);
nand U8021 (N_8021,N_7609,N_7357);
nor U8022 (N_8022,N_7567,N_7260);
nor U8023 (N_8023,N_7540,N_7542);
or U8024 (N_8024,N_7418,N_7406);
and U8025 (N_8025,N_7597,N_7747);
and U8026 (N_8026,N_7232,N_7355);
nor U8027 (N_8027,N_7338,N_7654);
nor U8028 (N_8028,N_7278,N_7277);
nand U8029 (N_8029,N_7304,N_7628);
or U8030 (N_8030,N_7413,N_7560);
nand U8031 (N_8031,N_7740,N_7596);
nand U8032 (N_8032,N_7615,N_7219);
and U8033 (N_8033,N_7202,N_7214);
and U8034 (N_8034,N_7388,N_7588);
nor U8035 (N_8035,N_7776,N_7434);
nand U8036 (N_8036,N_7460,N_7473);
nand U8037 (N_8037,N_7452,N_7372);
and U8038 (N_8038,N_7672,N_7748);
nand U8039 (N_8039,N_7517,N_7799);
or U8040 (N_8040,N_7728,N_7745);
nor U8041 (N_8041,N_7229,N_7479);
nor U8042 (N_8042,N_7592,N_7786);
nand U8043 (N_8043,N_7579,N_7408);
nor U8044 (N_8044,N_7387,N_7487);
nand U8045 (N_8045,N_7729,N_7627);
and U8046 (N_8046,N_7781,N_7459);
or U8047 (N_8047,N_7461,N_7368);
nor U8048 (N_8048,N_7442,N_7576);
nor U8049 (N_8049,N_7494,N_7332);
nor U8050 (N_8050,N_7578,N_7349);
or U8051 (N_8051,N_7414,N_7363);
nor U8052 (N_8052,N_7416,N_7251);
and U8053 (N_8053,N_7584,N_7530);
or U8054 (N_8054,N_7456,N_7480);
or U8055 (N_8055,N_7725,N_7481);
and U8056 (N_8056,N_7258,N_7508);
nand U8057 (N_8057,N_7476,N_7378);
and U8058 (N_8058,N_7331,N_7555);
and U8059 (N_8059,N_7634,N_7571);
or U8060 (N_8060,N_7419,N_7706);
nand U8061 (N_8061,N_7531,N_7769);
and U8062 (N_8062,N_7620,N_7369);
or U8063 (N_8063,N_7724,N_7683);
or U8064 (N_8064,N_7411,N_7207);
nand U8065 (N_8065,N_7430,N_7490);
or U8066 (N_8066,N_7757,N_7587);
nor U8067 (N_8067,N_7505,N_7651);
and U8068 (N_8068,N_7446,N_7633);
and U8069 (N_8069,N_7647,N_7701);
nor U8070 (N_8070,N_7742,N_7302);
and U8071 (N_8071,N_7297,N_7719);
and U8072 (N_8072,N_7614,N_7663);
nand U8073 (N_8073,N_7572,N_7696);
nand U8074 (N_8074,N_7437,N_7265);
nand U8075 (N_8075,N_7622,N_7498);
nand U8076 (N_8076,N_7379,N_7257);
and U8077 (N_8077,N_7688,N_7353);
and U8078 (N_8078,N_7760,N_7602);
nand U8079 (N_8079,N_7342,N_7563);
nor U8080 (N_8080,N_7677,N_7507);
nor U8081 (N_8081,N_7279,N_7275);
nor U8082 (N_8082,N_7347,N_7333);
or U8083 (N_8083,N_7315,N_7293);
or U8084 (N_8084,N_7671,N_7500);
nor U8085 (N_8085,N_7415,N_7551);
and U8086 (N_8086,N_7491,N_7720);
and U8087 (N_8087,N_7230,N_7244);
and U8088 (N_8088,N_7716,N_7383);
nand U8089 (N_8089,N_7472,N_7240);
nor U8090 (N_8090,N_7787,N_7580);
or U8091 (N_8091,N_7211,N_7759);
nor U8092 (N_8092,N_7444,N_7624);
and U8093 (N_8093,N_7521,N_7638);
nand U8094 (N_8094,N_7380,N_7524);
or U8095 (N_8095,N_7255,N_7451);
nand U8096 (N_8096,N_7396,N_7751);
and U8097 (N_8097,N_7566,N_7453);
or U8098 (N_8098,N_7610,N_7547);
nand U8099 (N_8099,N_7775,N_7394);
xnor U8100 (N_8100,N_7720,N_7628);
and U8101 (N_8101,N_7207,N_7435);
and U8102 (N_8102,N_7203,N_7606);
nand U8103 (N_8103,N_7788,N_7623);
nand U8104 (N_8104,N_7319,N_7200);
nor U8105 (N_8105,N_7511,N_7353);
nor U8106 (N_8106,N_7491,N_7239);
nor U8107 (N_8107,N_7366,N_7686);
or U8108 (N_8108,N_7627,N_7360);
and U8109 (N_8109,N_7781,N_7454);
nand U8110 (N_8110,N_7245,N_7773);
nor U8111 (N_8111,N_7798,N_7729);
nand U8112 (N_8112,N_7298,N_7347);
nand U8113 (N_8113,N_7333,N_7589);
nand U8114 (N_8114,N_7586,N_7318);
nor U8115 (N_8115,N_7307,N_7779);
nor U8116 (N_8116,N_7687,N_7614);
nor U8117 (N_8117,N_7739,N_7761);
and U8118 (N_8118,N_7416,N_7525);
nor U8119 (N_8119,N_7490,N_7737);
nor U8120 (N_8120,N_7323,N_7364);
or U8121 (N_8121,N_7204,N_7305);
or U8122 (N_8122,N_7563,N_7562);
and U8123 (N_8123,N_7776,N_7499);
and U8124 (N_8124,N_7515,N_7525);
nand U8125 (N_8125,N_7783,N_7423);
or U8126 (N_8126,N_7673,N_7395);
and U8127 (N_8127,N_7355,N_7508);
nand U8128 (N_8128,N_7356,N_7508);
nor U8129 (N_8129,N_7757,N_7396);
or U8130 (N_8130,N_7455,N_7702);
nor U8131 (N_8131,N_7445,N_7627);
nand U8132 (N_8132,N_7476,N_7219);
nand U8133 (N_8133,N_7764,N_7255);
nor U8134 (N_8134,N_7205,N_7495);
and U8135 (N_8135,N_7686,N_7580);
or U8136 (N_8136,N_7565,N_7430);
or U8137 (N_8137,N_7455,N_7607);
or U8138 (N_8138,N_7237,N_7606);
nand U8139 (N_8139,N_7462,N_7511);
or U8140 (N_8140,N_7325,N_7640);
or U8141 (N_8141,N_7540,N_7310);
nand U8142 (N_8142,N_7254,N_7473);
or U8143 (N_8143,N_7302,N_7671);
xor U8144 (N_8144,N_7354,N_7782);
or U8145 (N_8145,N_7577,N_7237);
or U8146 (N_8146,N_7781,N_7403);
xor U8147 (N_8147,N_7264,N_7266);
nor U8148 (N_8148,N_7236,N_7708);
nand U8149 (N_8149,N_7691,N_7303);
nor U8150 (N_8150,N_7674,N_7652);
nand U8151 (N_8151,N_7491,N_7445);
nor U8152 (N_8152,N_7762,N_7627);
nor U8153 (N_8153,N_7600,N_7760);
nand U8154 (N_8154,N_7796,N_7271);
nand U8155 (N_8155,N_7321,N_7312);
nand U8156 (N_8156,N_7540,N_7779);
and U8157 (N_8157,N_7290,N_7351);
and U8158 (N_8158,N_7403,N_7433);
or U8159 (N_8159,N_7638,N_7445);
nand U8160 (N_8160,N_7250,N_7733);
nor U8161 (N_8161,N_7268,N_7522);
nor U8162 (N_8162,N_7207,N_7350);
and U8163 (N_8163,N_7201,N_7429);
or U8164 (N_8164,N_7253,N_7206);
nand U8165 (N_8165,N_7232,N_7477);
nand U8166 (N_8166,N_7774,N_7613);
nand U8167 (N_8167,N_7220,N_7372);
and U8168 (N_8168,N_7400,N_7495);
xor U8169 (N_8169,N_7305,N_7487);
and U8170 (N_8170,N_7712,N_7516);
nand U8171 (N_8171,N_7362,N_7430);
nor U8172 (N_8172,N_7699,N_7434);
or U8173 (N_8173,N_7408,N_7231);
and U8174 (N_8174,N_7442,N_7528);
nand U8175 (N_8175,N_7277,N_7289);
or U8176 (N_8176,N_7745,N_7247);
nand U8177 (N_8177,N_7407,N_7504);
and U8178 (N_8178,N_7785,N_7226);
and U8179 (N_8179,N_7720,N_7529);
nand U8180 (N_8180,N_7764,N_7215);
nand U8181 (N_8181,N_7617,N_7710);
nor U8182 (N_8182,N_7762,N_7304);
and U8183 (N_8183,N_7642,N_7464);
nor U8184 (N_8184,N_7276,N_7232);
nor U8185 (N_8185,N_7664,N_7680);
nand U8186 (N_8186,N_7727,N_7742);
nand U8187 (N_8187,N_7682,N_7381);
or U8188 (N_8188,N_7226,N_7254);
nor U8189 (N_8189,N_7684,N_7579);
nand U8190 (N_8190,N_7403,N_7698);
or U8191 (N_8191,N_7797,N_7332);
or U8192 (N_8192,N_7359,N_7665);
nor U8193 (N_8193,N_7433,N_7311);
nand U8194 (N_8194,N_7357,N_7647);
and U8195 (N_8195,N_7700,N_7670);
nor U8196 (N_8196,N_7599,N_7371);
or U8197 (N_8197,N_7572,N_7609);
and U8198 (N_8198,N_7663,N_7206);
or U8199 (N_8199,N_7716,N_7389);
nand U8200 (N_8200,N_7529,N_7387);
and U8201 (N_8201,N_7216,N_7287);
or U8202 (N_8202,N_7409,N_7250);
or U8203 (N_8203,N_7422,N_7452);
and U8204 (N_8204,N_7622,N_7241);
and U8205 (N_8205,N_7438,N_7666);
nor U8206 (N_8206,N_7676,N_7313);
nand U8207 (N_8207,N_7414,N_7640);
and U8208 (N_8208,N_7580,N_7689);
nand U8209 (N_8209,N_7369,N_7722);
xnor U8210 (N_8210,N_7652,N_7339);
or U8211 (N_8211,N_7298,N_7377);
and U8212 (N_8212,N_7610,N_7473);
nand U8213 (N_8213,N_7417,N_7764);
nand U8214 (N_8214,N_7499,N_7732);
and U8215 (N_8215,N_7396,N_7784);
or U8216 (N_8216,N_7232,N_7315);
nand U8217 (N_8217,N_7672,N_7597);
or U8218 (N_8218,N_7674,N_7563);
nor U8219 (N_8219,N_7311,N_7401);
and U8220 (N_8220,N_7747,N_7307);
nor U8221 (N_8221,N_7728,N_7746);
or U8222 (N_8222,N_7614,N_7211);
and U8223 (N_8223,N_7379,N_7250);
and U8224 (N_8224,N_7242,N_7610);
or U8225 (N_8225,N_7484,N_7611);
or U8226 (N_8226,N_7604,N_7665);
nand U8227 (N_8227,N_7267,N_7266);
xnor U8228 (N_8228,N_7483,N_7463);
and U8229 (N_8229,N_7347,N_7662);
and U8230 (N_8230,N_7326,N_7489);
and U8231 (N_8231,N_7552,N_7389);
nor U8232 (N_8232,N_7549,N_7403);
nand U8233 (N_8233,N_7412,N_7362);
or U8234 (N_8234,N_7673,N_7643);
nor U8235 (N_8235,N_7614,N_7514);
or U8236 (N_8236,N_7784,N_7690);
xor U8237 (N_8237,N_7538,N_7379);
and U8238 (N_8238,N_7334,N_7222);
nor U8239 (N_8239,N_7512,N_7629);
or U8240 (N_8240,N_7699,N_7411);
or U8241 (N_8241,N_7560,N_7742);
and U8242 (N_8242,N_7513,N_7670);
nor U8243 (N_8243,N_7593,N_7349);
nor U8244 (N_8244,N_7527,N_7720);
or U8245 (N_8245,N_7489,N_7383);
or U8246 (N_8246,N_7654,N_7593);
nand U8247 (N_8247,N_7697,N_7622);
nor U8248 (N_8248,N_7323,N_7677);
or U8249 (N_8249,N_7631,N_7771);
or U8250 (N_8250,N_7779,N_7698);
nor U8251 (N_8251,N_7668,N_7632);
or U8252 (N_8252,N_7615,N_7364);
and U8253 (N_8253,N_7583,N_7384);
and U8254 (N_8254,N_7435,N_7752);
or U8255 (N_8255,N_7390,N_7662);
and U8256 (N_8256,N_7492,N_7552);
nor U8257 (N_8257,N_7527,N_7715);
or U8258 (N_8258,N_7639,N_7359);
or U8259 (N_8259,N_7755,N_7283);
and U8260 (N_8260,N_7335,N_7213);
nand U8261 (N_8261,N_7496,N_7661);
nor U8262 (N_8262,N_7549,N_7628);
or U8263 (N_8263,N_7662,N_7659);
nor U8264 (N_8264,N_7453,N_7492);
or U8265 (N_8265,N_7618,N_7485);
nor U8266 (N_8266,N_7201,N_7211);
or U8267 (N_8267,N_7464,N_7606);
and U8268 (N_8268,N_7211,N_7772);
nand U8269 (N_8269,N_7637,N_7747);
nor U8270 (N_8270,N_7319,N_7470);
or U8271 (N_8271,N_7678,N_7271);
nand U8272 (N_8272,N_7689,N_7376);
and U8273 (N_8273,N_7691,N_7578);
or U8274 (N_8274,N_7427,N_7429);
or U8275 (N_8275,N_7571,N_7498);
and U8276 (N_8276,N_7471,N_7464);
and U8277 (N_8277,N_7328,N_7706);
nor U8278 (N_8278,N_7586,N_7487);
or U8279 (N_8279,N_7266,N_7627);
nand U8280 (N_8280,N_7515,N_7493);
nand U8281 (N_8281,N_7247,N_7315);
and U8282 (N_8282,N_7310,N_7439);
and U8283 (N_8283,N_7606,N_7622);
nor U8284 (N_8284,N_7202,N_7617);
and U8285 (N_8285,N_7366,N_7537);
nand U8286 (N_8286,N_7724,N_7423);
or U8287 (N_8287,N_7653,N_7284);
nor U8288 (N_8288,N_7650,N_7276);
nand U8289 (N_8289,N_7279,N_7235);
nand U8290 (N_8290,N_7553,N_7312);
and U8291 (N_8291,N_7490,N_7314);
and U8292 (N_8292,N_7288,N_7689);
and U8293 (N_8293,N_7239,N_7596);
nand U8294 (N_8294,N_7397,N_7274);
nor U8295 (N_8295,N_7678,N_7530);
nor U8296 (N_8296,N_7317,N_7405);
nand U8297 (N_8297,N_7437,N_7585);
or U8298 (N_8298,N_7385,N_7735);
nor U8299 (N_8299,N_7759,N_7504);
nor U8300 (N_8300,N_7501,N_7290);
nand U8301 (N_8301,N_7491,N_7762);
and U8302 (N_8302,N_7595,N_7415);
nor U8303 (N_8303,N_7334,N_7399);
nor U8304 (N_8304,N_7616,N_7600);
nor U8305 (N_8305,N_7712,N_7284);
nor U8306 (N_8306,N_7685,N_7467);
nand U8307 (N_8307,N_7214,N_7539);
nor U8308 (N_8308,N_7441,N_7338);
and U8309 (N_8309,N_7767,N_7551);
or U8310 (N_8310,N_7625,N_7720);
and U8311 (N_8311,N_7428,N_7657);
nor U8312 (N_8312,N_7410,N_7562);
nand U8313 (N_8313,N_7344,N_7726);
and U8314 (N_8314,N_7630,N_7339);
and U8315 (N_8315,N_7605,N_7530);
nand U8316 (N_8316,N_7294,N_7582);
nand U8317 (N_8317,N_7204,N_7628);
or U8318 (N_8318,N_7487,N_7270);
nor U8319 (N_8319,N_7246,N_7715);
and U8320 (N_8320,N_7631,N_7693);
and U8321 (N_8321,N_7503,N_7398);
or U8322 (N_8322,N_7247,N_7206);
and U8323 (N_8323,N_7246,N_7746);
nor U8324 (N_8324,N_7689,N_7220);
or U8325 (N_8325,N_7585,N_7627);
nand U8326 (N_8326,N_7700,N_7746);
nor U8327 (N_8327,N_7518,N_7450);
and U8328 (N_8328,N_7435,N_7643);
or U8329 (N_8329,N_7488,N_7256);
nor U8330 (N_8330,N_7707,N_7781);
nor U8331 (N_8331,N_7633,N_7459);
nor U8332 (N_8332,N_7765,N_7532);
nor U8333 (N_8333,N_7732,N_7424);
nor U8334 (N_8334,N_7492,N_7353);
nor U8335 (N_8335,N_7757,N_7276);
and U8336 (N_8336,N_7606,N_7731);
nor U8337 (N_8337,N_7711,N_7607);
or U8338 (N_8338,N_7235,N_7746);
nor U8339 (N_8339,N_7531,N_7553);
nand U8340 (N_8340,N_7374,N_7284);
and U8341 (N_8341,N_7518,N_7479);
or U8342 (N_8342,N_7365,N_7516);
or U8343 (N_8343,N_7746,N_7669);
or U8344 (N_8344,N_7282,N_7294);
nor U8345 (N_8345,N_7724,N_7343);
or U8346 (N_8346,N_7602,N_7724);
and U8347 (N_8347,N_7559,N_7369);
nand U8348 (N_8348,N_7638,N_7600);
nand U8349 (N_8349,N_7710,N_7443);
and U8350 (N_8350,N_7680,N_7757);
nand U8351 (N_8351,N_7761,N_7582);
or U8352 (N_8352,N_7309,N_7449);
nand U8353 (N_8353,N_7314,N_7667);
or U8354 (N_8354,N_7549,N_7590);
nor U8355 (N_8355,N_7325,N_7402);
and U8356 (N_8356,N_7598,N_7218);
nand U8357 (N_8357,N_7484,N_7314);
and U8358 (N_8358,N_7523,N_7715);
nand U8359 (N_8359,N_7414,N_7326);
nor U8360 (N_8360,N_7449,N_7558);
nor U8361 (N_8361,N_7477,N_7497);
or U8362 (N_8362,N_7496,N_7553);
or U8363 (N_8363,N_7493,N_7357);
nand U8364 (N_8364,N_7262,N_7792);
nor U8365 (N_8365,N_7472,N_7372);
nand U8366 (N_8366,N_7223,N_7259);
nor U8367 (N_8367,N_7507,N_7551);
nor U8368 (N_8368,N_7287,N_7793);
nand U8369 (N_8369,N_7288,N_7397);
or U8370 (N_8370,N_7763,N_7543);
nand U8371 (N_8371,N_7220,N_7530);
or U8372 (N_8372,N_7744,N_7380);
and U8373 (N_8373,N_7713,N_7350);
and U8374 (N_8374,N_7585,N_7425);
and U8375 (N_8375,N_7293,N_7634);
or U8376 (N_8376,N_7414,N_7469);
xor U8377 (N_8377,N_7257,N_7566);
or U8378 (N_8378,N_7376,N_7763);
and U8379 (N_8379,N_7799,N_7548);
nand U8380 (N_8380,N_7666,N_7498);
and U8381 (N_8381,N_7622,N_7268);
and U8382 (N_8382,N_7646,N_7486);
and U8383 (N_8383,N_7334,N_7212);
nor U8384 (N_8384,N_7290,N_7562);
nand U8385 (N_8385,N_7204,N_7298);
nor U8386 (N_8386,N_7498,N_7269);
nand U8387 (N_8387,N_7252,N_7345);
or U8388 (N_8388,N_7443,N_7471);
nor U8389 (N_8389,N_7628,N_7677);
or U8390 (N_8390,N_7417,N_7224);
and U8391 (N_8391,N_7700,N_7209);
and U8392 (N_8392,N_7712,N_7367);
nor U8393 (N_8393,N_7364,N_7563);
nand U8394 (N_8394,N_7776,N_7365);
and U8395 (N_8395,N_7359,N_7248);
nand U8396 (N_8396,N_7733,N_7638);
nor U8397 (N_8397,N_7466,N_7777);
or U8398 (N_8398,N_7344,N_7324);
nand U8399 (N_8399,N_7375,N_7572);
nand U8400 (N_8400,N_8077,N_8196);
and U8401 (N_8401,N_8261,N_8152);
and U8402 (N_8402,N_7935,N_8262);
nor U8403 (N_8403,N_8234,N_8211);
and U8404 (N_8404,N_7941,N_7930);
and U8405 (N_8405,N_8361,N_7910);
or U8406 (N_8406,N_8248,N_8022);
or U8407 (N_8407,N_7868,N_7883);
nor U8408 (N_8408,N_8214,N_7878);
nand U8409 (N_8409,N_7990,N_7816);
nor U8410 (N_8410,N_7885,N_8087);
nand U8411 (N_8411,N_8319,N_8111);
nand U8412 (N_8412,N_8073,N_8386);
or U8413 (N_8413,N_7921,N_8182);
nand U8414 (N_8414,N_8284,N_7914);
nor U8415 (N_8415,N_8300,N_8035);
nor U8416 (N_8416,N_8217,N_8024);
and U8417 (N_8417,N_7993,N_8044);
nor U8418 (N_8418,N_8114,N_8018);
and U8419 (N_8419,N_8320,N_8219);
nand U8420 (N_8420,N_8137,N_8083);
and U8421 (N_8421,N_8351,N_8068);
or U8422 (N_8422,N_7928,N_8384);
or U8423 (N_8423,N_8075,N_8021);
nand U8424 (N_8424,N_8358,N_8168);
nor U8425 (N_8425,N_8247,N_8078);
or U8426 (N_8426,N_8370,N_8173);
nand U8427 (N_8427,N_7875,N_7934);
and U8428 (N_8428,N_8306,N_8134);
nor U8429 (N_8429,N_8239,N_8100);
and U8430 (N_8430,N_8290,N_8079);
and U8431 (N_8431,N_7911,N_8368);
and U8432 (N_8432,N_7819,N_8353);
xor U8433 (N_8433,N_8051,N_8169);
nand U8434 (N_8434,N_8039,N_8054);
nand U8435 (N_8435,N_8145,N_8286);
nand U8436 (N_8436,N_8162,N_8123);
and U8437 (N_8437,N_8252,N_8237);
nand U8438 (N_8438,N_8226,N_8198);
or U8439 (N_8439,N_8050,N_7812);
xnor U8440 (N_8440,N_7938,N_8380);
and U8441 (N_8441,N_8121,N_7969);
and U8442 (N_8442,N_8258,N_7842);
and U8443 (N_8443,N_8243,N_8263);
and U8444 (N_8444,N_8388,N_8143);
and U8445 (N_8445,N_8174,N_8255);
nand U8446 (N_8446,N_8276,N_8185);
and U8447 (N_8447,N_8098,N_8313);
and U8448 (N_8448,N_8155,N_8141);
or U8449 (N_8449,N_8249,N_8325);
nand U8450 (N_8450,N_8347,N_8277);
or U8451 (N_8451,N_7858,N_8144);
or U8452 (N_8452,N_7957,N_7915);
or U8453 (N_8453,N_8374,N_8045);
nand U8454 (N_8454,N_8067,N_7877);
and U8455 (N_8455,N_8378,N_8326);
nand U8456 (N_8456,N_8375,N_7949);
xnor U8457 (N_8457,N_8164,N_8101);
nor U8458 (N_8458,N_8146,N_8203);
and U8459 (N_8459,N_8395,N_8007);
nor U8460 (N_8460,N_8228,N_8046);
and U8461 (N_8461,N_7817,N_7988);
nor U8462 (N_8462,N_8202,N_8092);
nor U8463 (N_8463,N_8357,N_8222);
nand U8464 (N_8464,N_7971,N_8321);
nand U8465 (N_8465,N_7968,N_8089);
and U8466 (N_8466,N_8016,N_7813);
or U8467 (N_8467,N_8015,N_7897);
nor U8468 (N_8468,N_8371,N_8342);
and U8469 (N_8469,N_8195,N_8317);
nor U8470 (N_8470,N_8085,N_7952);
and U8471 (N_8471,N_7963,N_8107);
nand U8472 (N_8472,N_7978,N_8186);
nand U8473 (N_8473,N_8148,N_7997);
nand U8474 (N_8474,N_7999,N_8381);
nor U8475 (N_8475,N_7942,N_8221);
nand U8476 (N_8476,N_7805,N_7815);
nor U8477 (N_8477,N_7986,N_7857);
nand U8478 (N_8478,N_8027,N_7840);
nand U8479 (N_8479,N_7996,N_8294);
nand U8480 (N_8480,N_7987,N_8009);
or U8481 (N_8481,N_8204,N_7814);
and U8482 (N_8482,N_8333,N_7848);
nand U8483 (N_8483,N_8028,N_8244);
or U8484 (N_8484,N_8270,N_8398);
nand U8485 (N_8485,N_8130,N_8177);
nand U8486 (N_8486,N_8070,N_7965);
and U8487 (N_8487,N_8029,N_8346);
xor U8488 (N_8488,N_7977,N_7959);
and U8489 (N_8489,N_8090,N_7822);
xor U8490 (N_8490,N_8036,N_8205);
and U8491 (N_8491,N_8298,N_8056);
nand U8492 (N_8492,N_8264,N_8212);
nor U8493 (N_8493,N_8133,N_7860);
nor U8494 (N_8494,N_8088,N_7943);
and U8495 (N_8495,N_8391,N_8136);
nand U8496 (N_8496,N_7899,N_7931);
and U8497 (N_8497,N_8251,N_8335);
xnor U8498 (N_8498,N_8181,N_7871);
and U8499 (N_8499,N_8063,N_8175);
or U8500 (N_8500,N_7803,N_7884);
nor U8501 (N_8501,N_8176,N_8309);
or U8502 (N_8502,N_8058,N_8301);
nor U8503 (N_8503,N_7922,N_8376);
nand U8504 (N_8504,N_8151,N_7887);
and U8505 (N_8505,N_8245,N_8280);
and U8506 (N_8506,N_8236,N_7892);
nor U8507 (N_8507,N_8207,N_8097);
nand U8508 (N_8508,N_8149,N_7886);
nand U8509 (N_8509,N_7843,N_7827);
nand U8510 (N_8510,N_7889,N_7820);
and U8511 (N_8511,N_8010,N_8129);
and U8512 (N_8512,N_8392,N_8102);
nand U8513 (N_8513,N_8030,N_8360);
nand U8514 (N_8514,N_8139,N_7958);
and U8515 (N_8515,N_7852,N_8257);
or U8516 (N_8516,N_8275,N_8308);
nand U8517 (N_8517,N_8316,N_8383);
nand U8518 (N_8518,N_8055,N_8315);
and U8519 (N_8519,N_8288,N_8311);
and U8520 (N_8520,N_7953,N_8084);
nor U8521 (N_8521,N_8364,N_8314);
nor U8522 (N_8522,N_7847,N_7984);
nor U8523 (N_8523,N_7900,N_7998);
nor U8524 (N_8524,N_7912,N_7845);
or U8525 (N_8525,N_8206,N_8118);
or U8526 (N_8526,N_8112,N_7893);
nand U8527 (N_8527,N_8233,N_7923);
nor U8528 (N_8528,N_7936,N_7947);
and U8529 (N_8529,N_7909,N_7927);
and U8530 (N_8530,N_8366,N_7916);
nor U8531 (N_8531,N_8158,N_8281);
or U8532 (N_8532,N_7826,N_8242);
or U8533 (N_8533,N_8385,N_8256);
nand U8534 (N_8534,N_8047,N_7823);
nand U8535 (N_8535,N_7995,N_7946);
nor U8536 (N_8536,N_8095,N_8193);
nor U8537 (N_8537,N_7834,N_7907);
nand U8538 (N_8538,N_8017,N_8283);
or U8539 (N_8539,N_7821,N_8240);
xnor U8540 (N_8540,N_8362,N_8059);
nand U8541 (N_8541,N_7979,N_7970);
nand U8542 (N_8542,N_8006,N_8119);
and U8543 (N_8543,N_7981,N_8235);
nand U8544 (N_8544,N_8379,N_7891);
nor U8545 (N_8545,N_8069,N_8393);
and U8546 (N_8546,N_8200,N_7985);
and U8547 (N_8547,N_8225,N_7994);
or U8548 (N_8548,N_7967,N_8166);
and U8549 (N_8549,N_8387,N_8218);
nor U8550 (N_8550,N_7865,N_7841);
or U8551 (N_8551,N_8272,N_7926);
and U8552 (N_8552,N_8216,N_8305);
xor U8553 (N_8553,N_8334,N_8231);
nand U8554 (N_8554,N_8170,N_8259);
or U8555 (N_8555,N_8302,N_7824);
or U8556 (N_8556,N_7908,N_8003);
nand U8557 (N_8557,N_8183,N_8147);
or U8558 (N_8558,N_8061,N_7830);
or U8559 (N_8559,N_8020,N_7945);
nor U8560 (N_8560,N_8012,N_7854);
or U8561 (N_8561,N_8105,N_8285);
or U8562 (N_8562,N_7825,N_8188);
and U8563 (N_8563,N_8132,N_7901);
nor U8564 (N_8564,N_8241,N_7870);
or U8565 (N_8565,N_7828,N_8382);
and U8566 (N_8566,N_8184,N_8328);
nor U8567 (N_8567,N_8064,N_8008);
and U8568 (N_8568,N_7818,N_8080);
or U8569 (N_8569,N_8341,N_7955);
nor U8570 (N_8570,N_7913,N_8113);
nand U8571 (N_8571,N_7807,N_7937);
and U8572 (N_8572,N_8343,N_8135);
xor U8573 (N_8573,N_8140,N_8254);
or U8574 (N_8574,N_7831,N_8033);
nand U8575 (N_8575,N_8373,N_8116);
nor U8576 (N_8576,N_7944,N_7804);
or U8577 (N_8577,N_8229,N_7983);
nor U8578 (N_8578,N_8348,N_7829);
nor U8579 (N_8579,N_8253,N_8295);
or U8580 (N_8580,N_8224,N_7940);
nand U8581 (N_8581,N_8138,N_8032);
nor U8582 (N_8582,N_8238,N_7849);
nand U8583 (N_8583,N_8363,N_8215);
nand U8584 (N_8584,N_8165,N_8001);
nand U8585 (N_8585,N_8345,N_8005);
or U8586 (N_8586,N_8025,N_8266);
nand U8587 (N_8587,N_8394,N_7801);
and U8588 (N_8588,N_8344,N_8318);
and U8589 (N_8589,N_7919,N_8299);
nor U8590 (N_8590,N_8093,N_7880);
nand U8591 (N_8591,N_8250,N_8023);
and U8592 (N_8592,N_8389,N_8273);
or U8593 (N_8593,N_8332,N_7898);
or U8594 (N_8594,N_8082,N_7962);
nand U8595 (N_8595,N_8156,N_8043);
and U8596 (N_8596,N_8356,N_8372);
nor U8597 (N_8597,N_8367,N_8338);
and U8598 (N_8598,N_7972,N_8310);
or U8599 (N_8599,N_7976,N_8287);
and U8600 (N_8600,N_8209,N_8349);
or U8601 (N_8601,N_8180,N_8397);
or U8602 (N_8602,N_7837,N_8062);
nand U8603 (N_8603,N_7961,N_8339);
nand U8604 (N_8604,N_7933,N_7881);
or U8605 (N_8605,N_8167,N_7973);
xor U8606 (N_8606,N_8279,N_7835);
nand U8607 (N_8607,N_7832,N_8327);
or U8608 (N_8608,N_7974,N_8293);
nand U8609 (N_8609,N_7863,N_8034);
nor U8610 (N_8610,N_8142,N_8312);
and U8611 (N_8611,N_8004,N_8072);
nor U8612 (N_8612,N_7917,N_8267);
nor U8613 (N_8613,N_8191,N_8260);
nand U8614 (N_8614,N_8013,N_8268);
nor U8615 (N_8615,N_8128,N_7850);
or U8616 (N_8616,N_8197,N_8049);
nor U8617 (N_8617,N_8103,N_8187);
nor U8618 (N_8618,N_8127,N_8038);
or U8619 (N_8619,N_8037,N_8227);
or U8620 (N_8620,N_7802,N_8269);
and U8621 (N_8621,N_7920,N_8359);
or U8622 (N_8622,N_8230,N_8099);
nand U8623 (N_8623,N_7809,N_8126);
nor U8624 (N_8624,N_8091,N_8369);
and U8625 (N_8625,N_7896,N_7800);
and U8626 (N_8626,N_8124,N_8131);
and U8627 (N_8627,N_7888,N_8019);
or U8628 (N_8628,N_8172,N_8210);
nand U8629 (N_8629,N_7879,N_7806);
nand U8630 (N_8630,N_7864,N_7991);
or U8631 (N_8631,N_7866,N_7833);
and U8632 (N_8632,N_8014,N_8048);
and U8633 (N_8633,N_8041,N_8086);
and U8634 (N_8634,N_8150,N_7929);
nor U8635 (N_8635,N_8213,N_7956);
nor U8636 (N_8636,N_8076,N_8324);
or U8637 (N_8637,N_8192,N_8071);
and U8638 (N_8638,N_7905,N_7918);
and U8639 (N_8639,N_7904,N_7939);
or U8640 (N_8640,N_7960,N_8104);
nor U8641 (N_8641,N_8352,N_7844);
xor U8642 (N_8642,N_7876,N_8220);
or U8643 (N_8643,N_8122,N_8026);
and U8644 (N_8644,N_7855,N_8065);
and U8645 (N_8645,N_8081,N_7836);
or U8646 (N_8646,N_7954,N_8154);
nor U8647 (N_8647,N_7894,N_7882);
nand U8648 (N_8648,N_8110,N_8000);
or U8649 (N_8649,N_7964,N_7902);
nand U8650 (N_8650,N_8291,N_8208);
or U8651 (N_8651,N_7989,N_8060);
nor U8652 (N_8652,N_7869,N_8271);
xor U8653 (N_8653,N_8296,N_8053);
nor U8654 (N_8654,N_8117,N_8282);
and U8655 (N_8655,N_8329,N_8115);
or U8656 (N_8656,N_8125,N_7851);
or U8657 (N_8657,N_7890,N_8365);
nand U8658 (N_8658,N_8163,N_8171);
nand U8659 (N_8659,N_7808,N_7859);
xnor U8660 (N_8660,N_8120,N_8190);
or U8661 (N_8661,N_7874,N_8002);
nand U8662 (N_8662,N_8108,N_8396);
and U8663 (N_8663,N_8323,N_8307);
or U8664 (N_8664,N_8246,N_8297);
or U8665 (N_8665,N_8223,N_8232);
or U8666 (N_8666,N_8074,N_7861);
and U8667 (N_8667,N_8303,N_7932);
nand U8668 (N_8668,N_8331,N_8199);
nand U8669 (N_8669,N_8330,N_7838);
nor U8670 (N_8670,N_7975,N_8178);
nor U8671 (N_8671,N_8201,N_8354);
and U8672 (N_8672,N_8194,N_8337);
nor U8673 (N_8673,N_7811,N_7810);
and U8674 (N_8674,N_8109,N_8066);
and U8675 (N_8675,N_7925,N_8159);
and U8676 (N_8676,N_8336,N_8265);
nor U8677 (N_8677,N_8042,N_8355);
nand U8678 (N_8678,N_7856,N_8094);
nand U8679 (N_8679,N_8189,N_7862);
nor U8680 (N_8680,N_8153,N_8040);
nand U8681 (N_8681,N_8161,N_8106);
nor U8682 (N_8682,N_7867,N_7895);
xnor U8683 (N_8683,N_8052,N_8322);
or U8684 (N_8684,N_8399,N_8292);
or U8685 (N_8685,N_8031,N_7980);
and U8686 (N_8686,N_7992,N_8278);
nand U8687 (N_8687,N_7906,N_8390);
nor U8688 (N_8688,N_7839,N_7951);
nand U8689 (N_8689,N_8011,N_8289);
or U8690 (N_8690,N_7982,N_7948);
nor U8691 (N_8691,N_8179,N_7853);
and U8692 (N_8692,N_7903,N_8096);
nand U8693 (N_8693,N_8340,N_7966);
and U8694 (N_8694,N_7924,N_7846);
nor U8695 (N_8695,N_8304,N_8274);
and U8696 (N_8696,N_8157,N_8057);
or U8697 (N_8697,N_7873,N_7950);
nor U8698 (N_8698,N_8350,N_8160);
nor U8699 (N_8699,N_7872,N_8377);
and U8700 (N_8700,N_7931,N_7935);
nor U8701 (N_8701,N_8353,N_8278);
nand U8702 (N_8702,N_8210,N_8301);
nor U8703 (N_8703,N_8161,N_8192);
nand U8704 (N_8704,N_8100,N_8107);
or U8705 (N_8705,N_7805,N_8352);
xnor U8706 (N_8706,N_8144,N_7878);
nor U8707 (N_8707,N_7841,N_7962);
nand U8708 (N_8708,N_7821,N_8145);
nand U8709 (N_8709,N_8002,N_7896);
or U8710 (N_8710,N_8289,N_7882);
xor U8711 (N_8711,N_8265,N_8275);
nor U8712 (N_8712,N_8095,N_7973);
or U8713 (N_8713,N_8262,N_7894);
nor U8714 (N_8714,N_8006,N_8368);
nand U8715 (N_8715,N_7992,N_8183);
or U8716 (N_8716,N_8208,N_7899);
nor U8717 (N_8717,N_8247,N_8294);
and U8718 (N_8718,N_8167,N_8216);
nand U8719 (N_8719,N_7933,N_8394);
and U8720 (N_8720,N_8152,N_8183);
nor U8721 (N_8721,N_7974,N_8062);
nor U8722 (N_8722,N_8087,N_8130);
nand U8723 (N_8723,N_8071,N_7828);
or U8724 (N_8724,N_8372,N_8235);
or U8725 (N_8725,N_7987,N_7914);
nor U8726 (N_8726,N_8188,N_7844);
nand U8727 (N_8727,N_8299,N_8133);
or U8728 (N_8728,N_8325,N_8135);
nor U8729 (N_8729,N_8190,N_8394);
or U8730 (N_8730,N_8216,N_8178);
and U8731 (N_8731,N_8391,N_8058);
or U8732 (N_8732,N_8384,N_8217);
and U8733 (N_8733,N_8273,N_7962);
or U8734 (N_8734,N_8005,N_8218);
or U8735 (N_8735,N_7898,N_7883);
xor U8736 (N_8736,N_8388,N_7891);
nor U8737 (N_8737,N_8122,N_8189);
or U8738 (N_8738,N_8323,N_8351);
and U8739 (N_8739,N_8323,N_8061);
nor U8740 (N_8740,N_8345,N_7909);
or U8741 (N_8741,N_7839,N_8332);
nor U8742 (N_8742,N_7964,N_8228);
and U8743 (N_8743,N_8058,N_8168);
nor U8744 (N_8744,N_8130,N_8076);
or U8745 (N_8745,N_8127,N_8255);
or U8746 (N_8746,N_8248,N_8206);
nor U8747 (N_8747,N_7933,N_7920);
nand U8748 (N_8748,N_8273,N_8246);
and U8749 (N_8749,N_8064,N_7898);
or U8750 (N_8750,N_8092,N_8026);
nor U8751 (N_8751,N_7894,N_8182);
nor U8752 (N_8752,N_7975,N_8065);
nand U8753 (N_8753,N_8291,N_8194);
nor U8754 (N_8754,N_8234,N_8024);
nand U8755 (N_8755,N_8059,N_8230);
nand U8756 (N_8756,N_7962,N_8040);
nor U8757 (N_8757,N_7804,N_7837);
and U8758 (N_8758,N_8364,N_7907);
nand U8759 (N_8759,N_8277,N_7853);
or U8760 (N_8760,N_7984,N_8068);
nor U8761 (N_8761,N_7910,N_8144);
or U8762 (N_8762,N_8053,N_8034);
or U8763 (N_8763,N_7845,N_8263);
nor U8764 (N_8764,N_7832,N_7999);
nand U8765 (N_8765,N_7901,N_7840);
and U8766 (N_8766,N_8141,N_8398);
and U8767 (N_8767,N_8141,N_8234);
or U8768 (N_8768,N_7852,N_8067);
nor U8769 (N_8769,N_8287,N_7856);
or U8770 (N_8770,N_7835,N_8217);
or U8771 (N_8771,N_8288,N_8179);
nor U8772 (N_8772,N_7995,N_8040);
and U8773 (N_8773,N_8054,N_8370);
xnor U8774 (N_8774,N_7905,N_8126);
or U8775 (N_8775,N_8310,N_8308);
or U8776 (N_8776,N_7896,N_8368);
nand U8777 (N_8777,N_8309,N_7925);
or U8778 (N_8778,N_8263,N_7936);
or U8779 (N_8779,N_7910,N_8116);
nor U8780 (N_8780,N_7911,N_8243);
and U8781 (N_8781,N_8164,N_8365);
nand U8782 (N_8782,N_8065,N_8096);
nand U8783 (N_8783,N_8348,N_8084);
or U8784 (N_8784,N_7818,N_8317);
nand U8785 (N_8785,N_8261,N_8349);
nand U8786 (N_8786,N_7912,N_7871);
or U8787 (N_8787,N_7957,N_8281);
nand U8788 (N_8788,N_8312,N_7837);
and U8789 (N_8789,N_8085,N_8311);
and U8790 (N_8790,N_8376,N_7925);
nor U8791 (N_8791,N_8237,N_7806);
nand U8792 (N_8792,N_8183,N_8096);
or U8793 (N_8793,N_8046,N_7829);
nand U8794 (N_8794,N_8162,N_8100);
nand U8795 (N_8795,N_8315,N_8002);
and U8796 (N_8796,N_8306,N_8192);
and U8797 (N_8797,N_7857,N_8153);
nor U8798 (N_8798,N_7896,N_7804);
or U8799 (N_8799,N_7999,N_7905);
nand U8800 (N_8800,N_8258,N_7956);
or U8801 (N_8801,N_7891,N_7877);
nand U8802 (N_8802,N_7982,N_8189);
and U8803 (N_8803,N_8209,N_8260);
and U8804 (N_8804,N_8093,N_8116);
or U8805 (N_8805,N_8106,N_8087);
nand U8806 (N_8806,N_7951,N_8258);
and U8807 (N_8807,N_7907,N_8076);
and U8808 (N_8808,N_7997,N_8271);
or U8809 (N_8809,N_8243,N_8185);
or U8810 (N_8810,N_7938,N_7957);
or U8811 (N_8811,N_8094,N_8148);
nor U8812 (N_8812,N_8132,N_7827);
and U8813 (N_8813,N_7929,N_8200);
nor U8814 (N_8814,N_7823,N_8003);
and U8815 (N_8815,N_7942,N_8076);
nand U8816 (N_8816,N_8329,N_8275);
or U8817 (N_8817,N_8393,N_7900);
or U8818 (N_8818,N_8243,N_8236);
and U8819 (N_8819,N_7998,N_7842);
or U8820 (N_8820,N_8163,N_8188);
nor U8821 (N_8821,N_8017,N_7907);
nand U8822 (N_8822,N_8134,N_8070);
and U8823 (N_8823,N_8386,N_8315);
nand U8824 (N_8824,N_8316,N_8301);
and U8825 (N_8825,N_7828,N_7883);
nor U8826 (N_8826,N_8332,N_8002);
or U8827 (N_8827,N_8094,N_8005);
or U8828 (N_8828,N_7802,N_8216);
nand U8829 (N_8829,N_8068,N_8319);
nor U8830 (N_8830,N_8366,N_7942);
or U8831 (N_8831,N_7990,N_8370);
or U8832 (N_8832,N_8224,N_8221);
nor U8833 (N_8833,N_8167,N_7918);
nor U8834 (N_8834,N_8236,N_8248);
or U8835 (N_8835,N_8152,N_8093);
nor U8836 (N_8836,N_8299,N_7907);
and U8837 (N_8837,N_8187,N_8013);
and U8838 (N_8838,N_8285,N_8077);
or U8839 (N_8839,N_7803,N_8248);
or U8840 (N_8840,N_7852,N_8183);
or U8841 (N_8841,N_8258,N_7859);
or U8842 (N_8842,N_7819,N_8184);
nand U8843 (N_8843,N_8006,N_7928);
or U8844 (N_8844,N_8310,N_7805);
or U8845 (N_8845,N_8007,N_8050);
or U8846 (N_8846,N_8277,N_8106);
xnor U8847 (N_8847,N_8173,N_8256);
nor U8848 (N_8848,N_8160,N_7975);
and U8849 (N_8849,N_8056,N_8379);
nor U8850 (N_8850,N_8006,N_8144);
nor U8851 (N_8851,N_7970,N_8391);
or U8852 (N_8852,N_8219,N_7839);
or U8853 (N_8853,N_8143,N_7885);
or U8854 (N_8854,N_7959,N_8357);
or U8855 (N_8855,N_8209,N_7892);
xnor U8856 (N_8856,N_8213,N_8269);
nor U8857 (N_8857,N_8044,N_8287);
or U8858 (N_8858,N_7816,N_7883);
and U8859 (N_8859,N_7908,N_8397);
or U8860 (N_8860,N_7819,N_8108);
nor U8861 (N_8861,N_8236,N_8245);
or U8862 (N_8862,N_8027,N_8343);
or U8863 (N_8863,N_7941,N_7842);
nand U8864 (N_8864,N_8166,N_8243);
and U8865 (N_8865,N_7985,N_8278);
nand U8866 (N_8866,N_8072,N_7854);
or U8867 (N_8867,N_7944,N_8187);
or U8868 (N_8868,N_8313,N_8013);
xnor U8869 (N_8869,N_8074,N_8284);
nand U8870 (N_8870,N_8333,N_8336);
and U8871 (N_8871,N_8181,N_8239);
nor U8872 (N_8872,N_7953,N_8036);
nor U8873 (N_8873,N_8040,N_8352);
and U8874 (N_8874,N_8251,N_8279);
or U8875 (N_8875,N_8332,N_8108);
or U8876 (N_8876,N_8254,N_8303);
or U8877 (N_8877,N_8322,N_8192);
and U8878 (N_8878,N_8106,N_8344);
nand U8879 (N_8879,N_8382,N_8247);
or U8880 (N_8880,N_8098,N_8094);
nor U8881 (N_8881,N_8245,N_7830);
or U8882 (N_8882,N_7827,N_8119);
nand U8883 (N_8883,N_8026,N_8019);
and U8884 (N_8884,N_8214,N_7822);
or U8885 (N_8885,N_8145,N_8085);
and U8886 (N_8886,N_8298,N_8085);
nand U8887 (N_8887,N_8073,N_8360);
nor U8888 (N_8888,N_8296,N_8307);
or U8889 (N_8889,N_7987,N_8311);
and U8890 (N_8890,N_8074,N_7874);
nor U8891 (N_8891,N_8175,N_7810);
nand U8892 (N_8892,N_8259,N_7802);
nand U8893 (N_8893,N_8210,N_7856);
or U8894 (N_8894,N_8083,N_8322);
or U8895 (N_8895,N_8062,N_7939);
and U8896 (N_8896,N_8034,N_7840);
nand U8897 (N_8897,N_8042,N_7938);
and U8898 (N_8898,N_7942,N_8359);
nand U8899 (N_8899,N_7842,N_8263);
nor U8900 (N_8900,N_8172,N_8396);
and U8901 (N_8901,N_8337,N_8366);
and U8902 (N_8902,N_8252,N_8359);
or U8903 (N_8903,N_8203,N_7991);
nor U8904 (N_8904,N_8238,N_8298);
nor U8905 (N_8905,N_7924,N_7963);
xor U8906 (N_8906,N_8256,N_7947);
nand U8907 (N_8907,N_7843,N_7802);
nor U8908 (N_8908,N_8109,N_7993);
or U8909 (N_8909,N_8122,N_8024);
nor U8910 (N_8910,N_8231,N_7897);
or U8911 (N_8911,N_8121,N_7995);
and U8912 (N_8912,N_8384,N_7812);
or U8913 (N_8913,N_8386,N_8276);
and U8914 (N_8914,N_7870,N_8077);
nor U8915 (N_8915,N_8032,N_8251);
nor U8916 (N_8916,N_8051,N_7968);
nor U8917 (N_8917,N_8074,N_8118);
or U8918 (N_8918,N_8111,N_7852);
or U8919 (N_8919,N_8067,N_8371);
or U8920 (N_8920,N_8126,N_8121);
nor U8921 (N_8921,N_7983,N_8308);
nand U8922 (N_8922,N_7909,N_8100);
nor U8923 (N_8923,N_7848,N_8352);
or U8924 (N_8924,N_8325,N_8092);
or U8925 (N_8925,N_7991,N_8241);
or U8926 (N_8926,N_8211,N_8015);
nand U8927 (N_8927,N_8048,N_8119);
nor U8928 (N_8928,N_8068,N_8185);
nor U8929 (N_8929,N_8170,N_8249);
nor U8930 (N_8930,N_7845,N_7962);
nor U8931 (N_8931,N_7942,N_7863);
and U8932 (N_8932,N_8234,N_7872);
and U8933 (N_8933,N_8380,N_7853);
and U8934 (N_8934,N_8096,N_8112);
or U8935 (N_8935,N_7925,N_8095);
nand U8936 (N_8936,N_8310,N_8288);
or U8937 (N_8937,N_8368,N_8062);
xor U8938 (N_8938,N_7879,N_8243);
nor U8939 (N_8939,N_8153,N_8115);
and U8940 (N_8940,N_7903,N_7941);
nor U8941 (N_8941,N_8261,N_7842);
or U8942 (N_8942,N_7955,N_8069);
and U8943 (N_8943,N_8266,N_7980);
or U8944 (N_8944,N_8026,N_8070);
nor U8945 (N_8945,N_7918,N_8238);
or U8946 (N_8946,N_7828,N_8280);
xnor U8947 (N_8947,N_7949,N_7960);
or U8948 (N_8948,N_8351,N_8121);
or U8949 (N_8949,N_8303,N_8050);
or U8950 (N_8950,N_8053,N_7848);
and U8951 (N_8951,N_8034,N_8121);
nand U8952 (N_8952,N_8378,N_8180);
nand U8953 (N_8953,N_8344,N_8373);
and U8954 (N_8954,N_8160,N_8386);
nor U8955 (N_8955,N_7971,N_7803);
nor U8956 (N_8956,N_8104,N_8064);
nand U8957 (N_8957,N_7851,N_8176);
xnor U8958 (N_8958,N_8165,N_8188);
nand U8959 (N_8959,N_8275,N_8356);
and U8960 (N_8960,N_8135,N_8170);
or U8961 (N_8961,N_8155,N_8184);
and U8962 (N_8962,N_8108,N_8193);
nor U8963 (N_8963,N_8144,N_8240);
or U8964 (N_8964,N_7883,N_8223);
and U8965 (N_8965,N_8095,N_8061);
or U8966 (N_8966,N_7813,N_8073);
or U8967 (N_8967,N_8020,N_8218);
and U8968 (N_8968,N_7928,N_8257);
or U8969 (N_8969,N_8399,N_8060);
xor U8970 (N_8970,N_8016,N_8083);
and U8971 (N_8971,N_8097,N_8292);
or U8972 (N_8972,N_8398,N_8273);
nor U8973 (N_8973,N_8142,N_7806);
nor U8974 (N_8974,N_8123,N_8190);
nor U8975 (N_8975,N_8285,N_7980);
or U8976 (N_8976,N_8222,N_7934);
or U8977 (N_8977,N_7933,N_7931);
or U8978 (N_8978,N_8379,N_7867);
nand U8979 (N_8979,N_8060,N_8393);
and U8980 (N_8980,N_7811,N_7875);
nor U8981 (N_8981,N_8359,N_8250);
or U8982 (N_8982,N_8098,N_7949);
and U8983 (N_8983,N_8397,N_7865);
xor U8984 (N_8984,N_8371,N_8130);
and U8985 (N_8985,N_7938,N_8157);
and U8986 (N_8986,N_8338,N_8329);
or U8987 (N_8987,N_8152,N_8105);
and U8988 (N_8988,N_8342,N_7916);
nor U8989 (N_8989,N_7960,N_8268);
or U8990 (N_8990,N_8178,N_7985);
nor U8991 (N_8991,N_8084,N_7908);
or U8992 (N_8992,N_8208,N_7923);
xor U8993 (N_8993,N_8167,N_7992);
and U8994 (N_8994,N_8181,N_8000);
nor U8995 (N_8995,N_8368,N_8255);
nand U8996 (N_8996,N_7873,N_8146);
nand U8997 (N_8997,N_8378,N_8088);
or U8998 (N_8998,N_7903,N_7878);
or U8999 (N_8999,N_8392,N_7803);
and U9000 (N_9000,N_8964,N_8777);
or U9001 (N_9001,N_8966,N_8547);
nand U9002 (N_9002,N_8879,N_8438);
nand U9003 (N_9003,N_8685,N_8554);
and U9004 (N_9004,N_8718,N_8949);
or U9005 (N_9005,N_8682,N_8735);
or U9006 (N_9006,N_8586,N_8443);
or U9007 (N_9007,N_8546,N_8490);
or U9008 (N_9008,N_8894,N_8409);
xnor U9009 (N_9009,N_8415,N_8472);
or U9010 (N_9010,N_8992,N_8551);
and U9011 (N_9011,N_8560,N_8857);
nor U9012 (N_9012,N_8874,N_8549);
or U9013 (N_9013,N_8976,N_8734);
nand U9014 (N_9014,N_8641,N_8462);
nor U9015 (N_9015,N_8829,N_8492);
nor U9016 (N_9016,N_8770,N_8656);
and U9017 (N_9017,N_8494,N_8557);
nor U9018 (N_9018,N_8985,N_8615);
and U9019 (N_9019,N_8723,N_8968);
nand U9020 (N_9020,N_8830,N_8499);
and U9021 (N_9021,N_8452,N_8540);
and U9022 (N_9022,N_8878,N_8833);
nand U9023 (N_9023,N_8428,N_8513);
nand U9024 (N_9024,N_8593,N_8463);
nand U9025 (N_9025,N_8402,N_8819);
nor U9026 (N_9026,N_8902,N_8827);
xor U9027 (N_9027,N_8792,N_8401);
nor U9028 (N_9028,N_8496,N_8784);
nand U9029 (N_9029,N_8901,N_8487);
and U9030 (N_9030,N_8449,N_8793);
and U9031 (N_9031,N_8788,N_8629);
nand U9032 (N_9032,N_8437,N_8934);
and U9033 (N_9033,N_8954,N_8654);
and U9034 (N_9034,N_8893,N_8464);
and U9035 (N_9035,N_8647,N_8600);
nand U9036 (N_9036,N_8681,N_8757);
and U9037 (N_9037,N_8884,N_8798);
or U9038 (N_9038,N_8691,N_8753);
or U9039 (N_9039,N_8710,N_8899);
nand U9040 (N_9040,N_8679,N_8425);
and U9041 (N_9041,N_8765,N_8939);
nor U9042 (N_9042,N_8674,N_8942);
nand U9043 (N_9043,N_8477,N_8671);
nor U9044 (N_9044,N_8693,N_8446);
nor U9045 (N_9045,N_8683,N_8643);
nand U9046 (N_9046,N_8731,N_8680);
and U9047 (N_9047,N_8516,N_8673);
nor U9048 (N_9048,N_8801,N_8931);
nand U9049 (N_9049,N_8522,N_8905);
and U9050 (N_9050,N_8950,N_8532);
or U9051 (N_9051,N_8977,N_8910);
or U9052 (N_9052,N_8775,N_8995);
or U9053 (N_9053,N_8736,N_8810);
and U9054 (N_9054,N_8818,N_8839);
nor U9055 (N_9055,N_8527,N_8483);
and U9056 (N_9056,N_8805,N_8800);
and U9057 (N_9057,N_8589,N_8442);
and U9058 (N_9058,N_8928,N_8536);
nand U9059 (N_9059,N_8658,N_8825);
nor U9060 (N_9060,N_8448,N_8947);
or U9061 (N_9061,N_8523,N_8826);
nand U9062 (N_9062,N_8561,N_8815);
or U9063 (N_9063,N_8553,N_8970);
or U9064 (N_9064,N_8426,N_8537);
nand U9065 (N_9065,N_8650,N_8435);
and U9066 (N_9066,N_8828,N_8760);
and U9067 (N_9067,N_8555,N_8860);
nor U9068 (N_9068,N_8628,N_8503);
nor U9069 (N_9069,N_8748,N_8745);
or U9070 (N_9070,N_8993,N_8576);
and U9071 (N_9071,N_8602,N_8927);
and U9072 (N_9072,N_8943,N_8669);
and U9073 (N_9073,N_8807,N_8972);
and U9074 (N_9074,N_8648,N_8720);
nor U9075 (N_9075,N_8459,N_8870);
or U9076 (N_9076,N_8512,N_8456);
or U9077 (N_9077,N_8771,N_8953);
and U9078 (N_9078,N_8678,N_8724);
nand U9079 (N_9079,N_8668,N_8809);
nor U9080 (N_9080,N_8454,N_8541);
and U9081 (N_9081,N_8940,N_8861);
xor U9082 (N_9082,N_8661,N_8984);
nand U9083 (N_9083,N_8406,N_8530);
nor U9084 (N_9084,N_8704,N_8416);
nor U9085 (N_9085,N_8872,N_8424);
nand U9086 (N_9086,N_8746,N_8762);
nand U9087 (N_9087,N_8982,N_8812);
and U9088 (N_9088,N_8609,N_8996);
nand U9089 (N_9089,N_8559,N_8920);
and U9090 (N_9090,N_8690,N_8582);
nor U9091 (N_9091,N_8751,N_8447);
nand U9092 (N_9092,N_8623,N_8856);
nor U9093 (N_9093,N_8543,N_8687);
nand U9094 (N_9094,N_8946,N_8677);
nor U9095 (N_9095,N_8596,N_8877);
or U9096 (N_9096,N_8969,N_8725);
or U9097 (N_9097,N_8686,N_8956);
and U9098 (N_9098,N_8484,N_8880);
nand U9099 (N_9099,N_8733,N_8853);
nand U9100 (N_9100,N_8816,N_8486);
nand U9101 (N_9101,N_8469,N_8836);
or U9102 (N_9102,N_8515,N_8676);
and U9103 (N_9103,N_8610,N_8419);
nor U9104 (N_9104,N_8842,N_8700);
nor U9105 (N_9105,N_8823,N_8444);
or U9106 (N_9106,N_8420,N_8544);
or U9107 (N_9107,N_8550,N_8892);
or U9108 (N_9108,N_8886,N_8922);
nor U9109 (N_9109,N_8919,N_8958);
and U9110 (N_9110,N_8854,N_8450);
nor U9111 (N_9111,N_8479,N_8948);
or U9112 (N_9112,N_8403,N_8408);
nor U9113 (N_9113,N_8843,N_8505);
nor U9114 (N_9114,N_8897,N_8497);
nor U9115 (N_9115,N_8611,N_8867);
and U9116 (N_9116,N_8646,N_8714);
or U9117 (N_9117,N_8534,N_8707);
or U9118 (N_9118,N_8627,N_8821);
nor U9119 (N_9119,N_8875,N_8410);
and U9120 (N_9120,N_8808,N_8458);
and U9121 (N_9121,N_8434,N_8730);
nand U9122 (N_9122,N_8577,N_8657);
nand U9123 (N_9123,N_8885,N_8852);
nor U9124 (N_9124,N_8614,N_8844);
or U9125 (N_9125,N_8994,N_8439);
nor U9126 (N_9126,N_8903,N_8865);
or U9127 (N_9127,N_8590,N_8445);
and U9128 (N_9128,N_8502,N_8684);
and U9129 (N_9129,N_8432,N_8620);
xnor U9130 (N_9130,N_8598,N_8869);
and U9131 (N_9131,N_8743,N_8621);
and U9132 (N_9132,N_8727,N_8849);
nor U9133 (N_9133,N_8405,N_8906);
nor U9134 (N_9134,N_8506,N_8457);
nor U9135 (N_9135,N_8606,N_8491);
nand U9136 (N_9136,N_8747,N_8585);
nor U9137 (N_9137,N_8759,N_8630);
or U9138 (N_9138,N_8573,N_8847);
nand U9139 (N_9139,N_8649,N_8990);
and U9140 (N_9140,N_8433,N_8514);
or U9141 (N_9141,N_8619,N_8599);
nand U9142 (N_9142,N_8890,N_8570);
nor U9143 (N_9143,N_8915,N_8695);
and U9144 (N_9144,N_8556,N_8539);
and U9145 (N_9145,N_8473,N_8900);
nor U9146 (N_9146,N_8697,N_8813);
nor U9147 (N_9147,N_8507,N_8740);
and U9148 (N_9148,N_8659,N_8850);
or U9149 (N_9149,N_8711,N_8701);
nand U9150 (N_9150,N_8631,N_8485);
or U9151 (N_9151,N_8912,N_8768);
or U9152 (N_9152,N_8575,N_8838);
nor U9153 (N_9153,N_8988,N_8755);
or U9154 (N_9154,N_8719,N_8592);
or U9155 (N_9155,N_8841,N_8617);
nor U9156 (N_9156,N_8862,N_8519);
xnor U9157 (N_9157,N_8563,N_8859);
or U9158 (N_9158,N_8422,N_8607);
and U9159 (N_9159,N_8761,N_8907);
nand U9160 (N_9160,N_8766,N_8480);
nand U9161 (N_9161,N_8520,N_8778);
nor U9162 (N_9162,N_8495,N_8764);
and U9163 (N_9163,N_8717,N_8722);
nor U9164 (N_9164,N_8476,N_8639);
nor U9165 (N_9165,N_8430,N_8637);
and U9166 (N_9166,N_8866,N_8471);
or U9167 (N_9167,N_8705,N_8509);
and U9168 (N_9168,N_8873,N_8455);
and U9169 (N_9169,N_8750,N_8981);
nor U9170 (N_9170,N_8664,N_8655);
and U9171 (N_9171,N_8538,N_8989);
or U9172 (N_9172,N_8584,N_8451);
nor U9173 (N_9173,N_8797,N_8467);
nand U9174 (N_9174,N_8489,N_8971);
nand U9175 (N_9175,N_8672,N_8804);
nor U9176 (N_9176,N_8732,N_8583);
or U9177 (N_9177,N_8665,N_8998);
and U9178 (N_9178,N_8511,N_8604);
nand U9179 (N_9179,N_8587,N_8698);
nor U9180 (N_9180,N_8882,N_8634);
nor U9181 (N_9181,N_8817,N_8528);
or U9182 (N_9182,N_8752,N_8979);
nand U9183 (N_9183,N_8913,N_8688);
or U9184 (N_9184,N_8889,N_8887);
nand U9185 (N_9185,N_8820,N_8997);
nor U9186 (N_9186,N_8973,N_8962);
or U9187 (N_9187,N_8914,N_8712);
and U9188 (N_9188,N_8742,N_8531);
and U9189 (N_9189,N_8715,N_8500);
nor U9190 (N_9190,N_8675,N_8796);
or U9191 (N_9191,N_8930,N_8831);
or U9192 (N_9192,N_8653,N_8400);
nand U9193 (N_9193,N_8651,N_8945);
nand U9194 (N_9194,N_8963,N_8666);
and U9195 (N_9195,N_8917,N_8524);
or U9196 (N_9196,N_8786,N_8822);
and U9197 (N_9197,N_8959,N_8951);
xnor U9198 (N_9198,N_8662,N_8780);
nand U9199 (N_9199,N_8542,N_8474);
nand U9200 (N_9200,N_8638,N_8888);
nand U9201 (N_9201,N_8978,N_8987);
xnor U9202 (N_9202,N_8909,N_8744);
and U9203 (N_9203,N_8967,N_8645);
or U9204 (N_9204,N_8789,N_8633);
or U9205 (N_9205,N_8421,N_8773);
nor U9206 (N_9206,N_8578,N_8957);
or U9207 (N_9207,N_8453,N_8595);
and U9208 (N_9208,N_8787,N_8588);
and U9209 (N_9209,N_8411,N_8824);
nor U9210 (N_9210,N_8726,N_8689);
nand U9211 (N_9211,N_8883,N_8591);
or U9212 (N_9212,N_8518,N_8418);
nor U9213 (N_9213,N_8925,N_8840);
xnor U9214 (N_9214,N_8568,N_8703);
nand U9215 (N_9215,N_8613,N_8465);
xor U9216 (N_9216,N_8908,N_8709);
nor U9217 (N_9217,N_8916,N_8565);
and U9218 (N_9218,N_8652,N_8708);
nor U9219 (N_9219,N_8904,N_8802);
nor U9220 (N_9220,N_8414,N_8635);
and U9221 (N_9221,N_8558,N_8407);
xnor U9222 (N_9222,N_8427,N_8644);
and U9223 (N_9223,N_8603,N_8848);
and U9224 (N_9224,N_8937,N_8498);
and U9225 (N_9225,N_8837,N_8605);
or U9226 (N_9226,N_8846,N_8626);
nor U9227 (N_9227,N_8468,N_8552);
nor U9228 (N_9228,N_8622,N_8508);
nor U9229 (N_9229,N_8533,N_8895);
nand U9230 (N_9230,N_8814,N_8794);
and U9231 (N_9231,N_8481,N_8470);
nor U9232 (N_9232,N_8737,N_8699);
nand U9233 (N_9233,N_8834,N_8923);
or U9234 (N_9234,N_8924,N_8845);
nand U9235 (N_9235,N_8574,N_8571);
nor U9236 (N_9236,N_8423,N_8504);
nor U9237 (N_9237,N_8772,N_8624);
or U9238 (N_9238,N_8535,N_8436);
and U9239 (N_9239,N_8640,N_8567);
xor U9240 (N_9240,N_8694,N_8713);
or U9241 (N_9241,N_8756,N_8932);
nor U9242 (N_9242,N_8729,N_8803);
nor U9243 (N_9243,N_8811,N_8980);
and U9244 (N_9244,N_8785,N_8965);
and U9245 (N_9245,N_8851,N_8868);
and U9246 (N_9246,N_8521,N_8612);
or U9247 (N_9247,N_8991,N_8616);
and U9248 (N_9248,N_8955,N_8413);
or U9249 (N_9249,N_8918,N_8855);
nand U9250 (N_9250,N_8417,N_8608);
and U9251 (N_9251,N_8758,N_8754);
nand U9252 (N_9252,N_8832,N_8774);
nor U9253 (N_9253,N_8728,N_8983);
or U9254 (N_9254,N_8493,N_8941);
nand U9255 (N_9255,N_8716,N_8896);
and U9256 (N_9256,N_8929,N_8625);
and U9257 (N_9257,N_8935,N_8763);
or U9258 (N_9258,N_8858,N_8545);
xnor U9259 (N_9259,N_8580,N_8579);
nor U9260 (N_9260,N_8938,N_8881);
or U9261 (N_9261,N_8767,N_8569);
nand U9262 (N_9262,N_8779,N_8952);
or U9263 (N_9263,N_8431,N_8660);
or U9264 (N_9264,N_8526,N_8933);
or U9265 (N_9265,N_8741,N_8936);
nand U9266 (N_9266,N_8696,N_8466);
or U9267 (N_9267,N_8961,N_8806);
nand U9268 (N_9268,N_8670,N_8986);
nor U9269 (N_9269,N_8636,N_8488);
and U9270 (N_9270,N_8769,N_8782);
and U9271 (N_9271,N_8926,N_8921);
or U9272 (N_9272,N_8475,N_8482);
nor U9273 (N_9273,N_8642,N_8864);
nor U9274 (N_9274,N_8974,N_8429);
and U9275 (N_9275,N_8548,N_8478);
and U9276 (N_9276,N_8799,N_8440);
and U9277 (N_9277,N_8597,N_8790);
and U9278 (N_9278,N_8562,N_8461);
nor U9279 (N_9279,N_8501,N_8566);
or U9280 (N_9280,N_8667,N_8795);
nand U9281 (N_9281,N_8572,N_8891);
or U9282 (N_9282,N_8706,N_8632);
nor U9283 (N_9283,N_8911,N_8663);
and U9284 (N_9284,N_8702,N_8776);
and U9285 (N_9285,N_8975,N_8835);
nand U9286 (N_9286,N_8692,N_8404);
nand U9287 (N_9287,N_8999,N_8749);
xor U9288 (N_9288,N_8525,N_8783);
or U9289 (N_9289,N_8517,N_8460);
nor U9290 (N_9290,N_8529,N_8960);
and U9291 (N_9291,N_8581,N_8863);
nand U9292 (N_9292,N_8944,N_8601);
nand U9293 (N_9293,N_8739,N_8412);
nand U9294 (N_9294,N_8510,N_8721);
or U9295 (N_9295,N_8871,N_8618);
nor U9296 (N_9296,N_8876,N_8898);
nor U9297 (N_9297,N_8564,N_8781);
nand U9298 (N_9298,N_8791,N_8594);
nor U9299 (N_9299,N_8738,N_8441);
or U9300 (N_9300,N_8706,N_8850);
nand U9301 (N_9301,N_8563,N_8934);
nor U9302 (N_9302,N_8688,N_8719);
nand U9303 (N_9303,N_8465,N_8639);
and U9304 (N_9304,N_8842,N_8479);
and U9305 (N_9305,N_8950,N_8723);
and U9306 (N_9306,N_8578,N_8532);
nand U9307 (N_9307,N_8816,N_8449);
nand U9308 (N_9308,N_8697,N_8664);
or U9309 (N_9309,N_8557,N_8805);
nor U9310 (N_9310,N_8668,N_8854);
nor U9311 (N_9311,N_8570,N_8927);
nand U9312 (N_9312,N_8842,N_8570);
nand U9313 (N_9313,N_8774,N_8574);
or U9314 (N_9314,N_8840,N_8802);
and U9315 (N_9315,N_8623,N_8630);
or U9316 (N_9316,N_8733,N_8753);
or U9317 (N_9317,N_8657,N_8741);
xor U9318 (N_9318,N_8672,N_8998);
nand U9319 (N_9319,N_8591,N_8829);
nor U9320 (N_9320,N_8588,N_8968);
nor U9321 (N_9321,N_8756,N_8834);
nor U9322 (N_9322,N_8792,N_8414);
or U9323 (N_9323,N_8581,N_8729);
or U9324 (N_9324,N_8800,N_8701);
and U9325 (N_9325,N_8773,N_8662);
and U9326 (N_9326,N_8577,N_8562);
nor U9327 (N_9327,N_8717,N_8885);
nor U9328 (N_9328,N_8901,N_8806);
nor U9329 (N_9329,N_8815,N_8468);
nor U9330 (N_9330,N_8501,N_8589);
or U9331 (N_9331,N_8944,N_8524);
or U9332 (N_9332,N_8540,N_8768);
and U9333 (N_9333,N_8958,N_8889);
or U9334 (N_9334,N_8579,N_8758);
and U9335 (N_9335,N_8723,N_8544);
xor U9336 (N_9336,N_8818,N_8912);
nand U9337 (N_9337,N_8759,N_8433);
nand U9338 (N_9338,N_8411,N_8716);
or U9339 (N_9339,N_8872,N_8997);
and U9340 (N_9340,N_8425,N_8445);
nor U9341 (N_9341,N_8801,N_8427);
nand U9342 (N_9342,N_8402,N_8516);
nor U9343 (N_9343,N_8670,N_8904);
or U9344 (N_9344,N_8752,N_8763);
or U9345 (N_9345,N_8730,N_8492);
nand U9346 (N_9346,N_8842,N_8995);
nand U9347 (N_9347,N_8565,N_8679);
and U9348 (N_9348,N_8659,N_8746);
or U9349 (N_9349,N_8566,N_8481);
nor U9350 (N_9350,N_8708,N_8408);
or U9351 (N_9351,N_8471,N_8832);
nor U9352 (N_9352,N_8833,N_8795);
nand U9353 (N_9353,N_8528,N_8875);
or U9354 (N_9354,N_8772,N_8580);
nor U9355 (N_9355,N_8588,N_8823);
nor U9356 (N_9356,N_8924,N_8462);
nor U9357 (N_9357,N_8952,N_8747);
and U9358 (N_9358,N_8755,N_8474);
nand U9359 (N_9359,N_8548,N_8882);
and U9360 (N_9360,N_8572,N_8475);
nor U9361 (N_9361,N_8904,N_8664);
nand U9362 (N_9362,N_8598,N_8559);
or U9363 (N_9363,N_8568,N_8416);
and U9364 (N_9364,N_8780,N_8872);
nor U9365 (N_9365,N_8775,N_8428);
or U9366 (N_9366,N_8805,N_8785);
and U9367 (N_9367,N_8609,N_8887);
or U9368 (N_9368,N_8611,N_8526);
and U9369 (N_9369,N_8949,N_8650);
or U9370 (N_9370,N_8622,N_8640);
or U9371 (N_9371,N_8886,N_8661);
or U9372 (N_9372,N_8562,N_8893);
nand U9373 (N_9373,N_8771,N_8963);
and U9374 (N_9374,N_8559,N_8451);
and U9375 (N_9375,N_8497,N_8717);
nand U9376 (N_9376,N_8706,N_8495);
or U9377 (N_9377,N_8674,N_8987);
nand U9378 (N_9378,N_8891,N_8940);
or U9379 (N_9379,N_8950,N_8986);
nor U9380 (N_9380,N_8612,N_8466);
or U9381 (N_9381,N_8540,N_8740);
nand U9382 (N_9382,N_8593,N_8610);
nand U9383 (N_9383,N_8887,N_8855);
nand U9384 (N_9384,N_8702,N_8904);
nor U9385 (N_9385,N_8661,N_8421);
nand U9386 (N_9386,N_8957,N_8494);
and U9387 (N_9387,N_8616,N_8979);
and U9388 (N_9388,N_8767,N_8552);
or U9389 (N_9389,N_8606,N_8611);
and U9390 (N_9390,N_8700,N_8878);
nand U9391 (N_9391,N_8737,N_8958);
and U9392 (N_9392,N_8461,N_8546);
or U9393 (N_9393,N_8648,N_8699);
or U9394 (N_9394,N_8927,N_8539);
nand U9395 (N_9395,N_8546,N_8532);
or U9396 (N_9396,N_8540,N_8651);
and U9397 (N_9397,N_8470,N_8638);
and U9398 (N_9398,N_8516,N_8491);
nor U9399 (N_9399,N_8883,N_8669);
nor U9400 (N_9400,N_8861,N_8678);
or U9401 (N_9401,N_8747,N_8577);
and U9402 (N_9402,N_8467,N_8786);
and U9403 (N_9403,N_8710,N_8614);
or U9404 (N_9404,N_8634,N_8573);
nor U9405 (N_9405,N_8843,N_8491);
or U9406 (N_9406,N_8807,N_8822);
and U9407 (N_9407,N_8866,N_8992);
or U9408 (N_9408,N_8457,N_8807);
nor U9409 (N_9409,N_8639,N_8577);
or U9410 (N_9410,N_8826,N_8414);
nor U9411 (N_9411,N_8558,N_8804);
xnor U9412 (N_9412,N_8963,N_8748);
nor U9413 (N_9413,N_8700,N_8781);
nand U9414 (N_9414,N_8591,N_8471);
nand U9415 (N_9415,N_8811,N_8774);
nor U9416 (N_9416,N_8705,N_8717);
and U9417 (N_9417,N_8657,N_8696);
nand U9418 (N_9418,N_8519,N_8668);
or U9419 (N_9419,N_8761,N_8691);
and U9420 (N_9420,N_8540,N_8480);
nor U9421 (N_9421,N_8889,N_8758);
nor U9422 (N_9422,N_8903,N_8646);
nor U9423 (N_9423,N_8506,N_8507);
nand U9424 (N_9424,N_8544,N_8611);
nor U9425 (N_9425,N_8656,N_8950);
nand U9426 (N_9426,N_8729,N_8518);
and U9427 (N_9427,N_8675,N_8585);
nor U9428 (N_9428,N_8469,N_8550);
nor U9429 (N_9429,N_8412,N_8993);
nor U9430 (N_9430,N_8699,N_8490);
and U9431 (N_9431,N_8935,N_8942);
or U9432 (N_9432,N_8995,N_8498);
and U9433 (N_9433,N_8965,N_8778);
or U9434 (N_9434,N_8852,N_8492);
nand U9435 (N_9435,N_8555,N_8479);
or U9436 (N_9436,N_8437,N_8928);
or U9437 (N_9437,N_8733,N_8668);
nor U9438 (N_9438,N_8425,N_8853);
or U9439 (N_9439,N_8431,N_8496);
nand U9440 (N_9440,N_8873,N_8780);
nand U9441 (N_9441,N_8614,N_8484);
and U9442 (N_9442,N_8985,N_8523);
nand U9443 (N_9443,N_8774,N_8751);
and U9444 (N_9444,N_8732,N_8958);
nor U9445 (N_9445,N_8796,N_8845);
and U9446 (N_9446,N_8450,N_8630);
nand U9447 (N_9447,N_8978,N_8895);
or U9448 (N_9448,N_8554,N_8463);
nand U9449 (N_9449,N_8736,N_8679);
or U9450 (N_9450,N_8509,N_8512);
nor U9451 (N_9451,N_8423,N_8986);
nor U9452 (N_9452,N_8634,N_8823);
nor U9453 (N_9453,N_8937,N_8407);
and U9454 (N_9454,N_8491,N_8595);
and U9455 (N_9455,N_8979,N_8669);
or U9456 (N_9456,N_8951,N_8886);
nand U9457 (N_9457,N_8962,N_8803);
nand U9458 (N_9458,N_8671,N_8972);
nor U9459 (N_9459,N_8519,N_8416);
or U9460 (N_9460,N_8672,N_8970);
and U9461 (N_9461,N_8557,N_8966);
or U9462 (N_9462,N_8713,N_8854);
or U9463 (N_9463,N_8668,N_8801);
or U9464 (N_9464,N_8653,N_8812);
or U9465 (N_9465,N_8576,N_8779);
nor U9466 (N_9466,N_8966,N_8992);
nor U9467 (N_9467,N_8971,N_8881);
nor U9468 (N_9468,N_8906,N_8857);
nor U9469 (N_9469,N_8525,N_8431);
and U9470 (N_9470,N_8714,N_8618);
nand U9471 (N_9471,N_8718,N_8932);
nor U9472 (N_9472,N_8628,N_8789);
xnor U9473 (N_9473,N_8707,N_8867);
and U9474 (N_9474,N_8619,N_8958);
nand U9475 (N_9475,N_8556,N_8813);
or U9476 (N_9476,N_8669,N_8581);
nor U9477 (N_9477,N_8829,N_8879);
nand U9478 (N_9478,N_8980,N_8837);
and U9479 (N_9479,N_8659,N_8495);
or U9480 (N_9480,N_8400,N_8729);
nand U9481 (N_9481,N_8490,N_8452);
nor U9482 (N_9482,N_8540,N_8907);
nor U9483 (N_9483,N_8467,N_8780);
nor U9484 (N_9484,N_8662,N_8963);
or U9485 (N_9485,N_8911,N_8402);
nor U9486 (N_9486,N_8999,N_8783);
nor U9487 (N_9487,N_8668,N_8456);
nand U9488 (N_9488,N_8606,N_8450);
nor U9489 (N_9489,N_8742,N_8645);
nand U9490 (N_9490,N_8481,N_8681);
nor U9491 (N_9491,N_8844,N_8987);
or U9492 (N_9492,N_8542,N_8587);
nand U9493 (N_9493,N_8924,N_8487);
nand U9494 (N_9494,N_8444,N_8597);
or U9495 (N_9495,N_8812,N_8828);
and U9496 (N_9496,N_8483,N_8682);
and U9497 (N_9497,N_8784,N_8993);
nor U9498 (N_9498,N_8779,N_8774);
or U9499 (N_9499,N_8438,N_8561);
nor U9500 (N_9500,N_8422,N_8983);
and U9501 (N_9501,N_8795,N_8759);
nand U9502 (N_9502,N_8669,N_8992);
nor U9503 (N_9503,N_8747,N_8525);
or U9504 (N_9504,N_8728,N_8950);
nor U9505 (N_9505,N_8509,N_8673);
or U9506 (N_9506,N_8583,N_8611);
or U9507 (N_9507,N_8648,N_8491);
or U9508 (N_9508,N_8899,N_8910);
nand U9509 (N_9509,N_8652,N_8845);
or U9510 (N_9510,N_8694,N_8679);
and U9511 (N_9511,N_8483,N_8463);
nand U9512 (N_9512,N_8435,N_8527);
nand U9513 (N_9513,N_8843,N_8765);
nor U9514 (N_9514,N_8892,N_8419);
or U9515 (N_9515,N_8880,N_8944);
nor U9516 (N_9516,N_8454,N_8962);
nand U9517 (N_9517,N_8858,N_8792);
nor U9518 (N_9518,N_8845,N_8976);
nand U9519 (N_9519,N_8812,N_8444);
nor U9520 (N_9520,N_8544,N_8526);
or U9521 (N_9521,N_8571,N_8872);
nor U9522 (N_9522,N_8630,N_8654);
or U9523 (N_9523,N_8818,N_8710);
or U9524 (N_9524,N_8568,N_8715);
nor U9525 (N_9525,N_8999,N_8499);
and U9526 (N_9526,N_8491,N_8475);
nand U9527 (N_9527,N_8933,N_8657);
or U9528 (N_9528,N_8684,N_8422);
nor U9529 (N_9529,N_8895,N_8906);
nand U9530 (N_9530,N_8447,N_8927);
and U9531 (N_9531,N_8702,N_8741);
nand U9532 (N_9532,N_8535,N_8444);
and U9533 (N_9533,N_8927,N_8732);
and U9534 (N_9534,N_8762,N_8520);
and U9535 (N_9535,N_8433,N_8559);
nor U9536 (N_9536,N_8730,N_8952);
or U9537 (N_9537,N_8774,N_8693);
or U9538 (N_9538,N_8430,N_8836);
nand U9539 (N_9539,N_8881,N_8525);
nor U9540 (N_9540,N_8921,N_8688);
or U9541 (N_9541,N_8942,N_8727);
or U9542 (N_9542,N_8575,N_8474);
or U9543 (N_9543,N_8767,N_8886);
or U9544 (N_9544,N_8981,N_8551);
and U9545 (N_9545,N_8538,N_8974);
nand U9546 (N_9546,N_8775,N_8937);
nand U9547 (N_9547,N_8518,N_8547);
or U9548 (N_9548,N_8737,N_8769);
and U9549 (N_9549,N_8530,N_8434);
nor U9550 (N_9550,N_8886,N_8818);
nor U9551 (N_9551,N_8680,N_8887);
nor U9552 (N_9552,N_8618,N_8507);
nor U9553 (N_9553,N_8892,N_8593);
nor U9554 (N_9554,N_8924,N_8436);
nand U9555 (N_9555,N_8783,N_8728);
and U9556 (N_9556,N_8621,N_8683);
nand U9557 (N_9557,N_8569,N_8972);
nor U9558 (N_9558,N_8558,N_8429);
xor U9559 (N_9559,N_8521,N_8720);
nand U9560 (N_9560,N_8514,N_8495);
nand U9561 (N_9561,N_8426,N_8725);
nand U9562 (N_9562,N_8759,N_8472);
or U9563 (N_9563,N_8727,N_8534);
and U9564 (N_9564,N_8519,N_8947);
nand U9565 (N_9565,N_8902,N_8524);
nor U9566 (N_9566,N_8964,N_8744);
and U9567 (N_9567,N_8454,N_8510);
nand U9568 (N_9568,N_8506,N_8932);
nand U9569 (N_9569,N_8830,N_8745);
nand U9570 (N_9570,N_8685,N_8690);
or U9571 (N_9571,N_8851,N_8941);
nand U9572 (N_9572,N_8683,N_8980);
or U9573 (N_9573,N_8784,N_8426);
and U9574 (N_9574,N_8439,N_8549);
nand U9575 (N_9575,N_8592,N_8643);
nor U9576 (N_9576,N_8774,N_8400);
xor U9577 (N_9577,N_8738,N_8710);
or U9578 (N_9578,N_8636,N_8926);
nand U9579 (N_9579,N_8663,N_8777);
nand U9580 (N_9580,N_8649,N_8652);
and U9581 (N_9581,N_8904,N_8809);
or U9582 (N_9582,N_8592,N_8660);
and U9583 (N_9583,N_8462,N_8956);
nand U9584 (N_9584,N_8466,N_8606);
nand U9585 (N_9585,N_8767,N_8900);
or U9586 (N_9586,N_8723,N_8782);
nand U9587 (N_9587,N_8928,N_8791);
nand U9588 (N_9588,N_8460,N_8925);
or U9589 (N_9589,N_8426,N_8791);
nand U9590 (N_9590,N_8996,N_8549);
and U9591 (N_9591,N_8908,N_8622);
or U9592 (N_9592,N_8623,N_8528);
and U9593 (N_9593,N_8600,N_8621);
nor U9594 (N_9594,N_8480,N_8425);
or U9595 (N_9595,N_8467,N_8720);
or U9596 (N_9596,N_8827,N_8423);
and U9597 (N_9597,N_8784,N_8941);
nand U9598 (N_9598,N_8433,N_8595);
nand U9599 (N_9599,N_8881,N_8705);
and U9600 (N_9600,N_9224,N_9203);
or U9601 (N_9601,N_9500,N_9196);
nand U9602 (N_9602,N_9443,N_9345);
and U9603 (N_9603,N_9068,N_9321);
or U9604 (N_9604,N_9061,N_9503);
nor U9605 (N_9605,N_9009,N_9377);
nor U9606 (N_9606,N_9384,N_9066);
or U9607 (N_9607,N_9506,N_9168);
and U9608 (N_9608,N_9366,N_9323);
and U9609 (N_9609,N_9257,N_9198);
nand U9610 (N_9610,N_9012,N_9405);
nand U9611 (N_9611,N_9391,N_9581);
and U9612 (N_9612,N_9056,N_9263);
and U9613 (N_9613,N_9327,N_9139);
or U9614 (N_9614,N_9325,N_9097);
or U9615 (N_9615,N_9385,N_9507);
nor U9616 (N_9616,N_9580,N_9406);
and U9617 (N_9617,N_9311,N_9572);
nor U9618 (N_9618,N_9359,N_9451);
nor U9619 (N_9619,N_9045,N_9047);
nor U9620 (N_9620,N_9111,N_9424);
nor U9621 (N_9621,N_9130,N_9192);
nand U9622 (N_9622,N_9392,N_9560);
nand U9623 (N_9623,N_9396,N_9439);
or U9624 (N_9624,N_9032,N_9081);
nand U9625 (N_9625,N_9389,N_9169);
nor U9626 (N_9626,N_9307,N_9156);
and U9627 (N_9627,N_9352,N_9563);
or U9628 (N_9628,N_9233,N_9453);
nand U9629 (N_9629,N_9176,N_9513);
nor U9630 (N_9630,N_9252,N_9310);
nor U9631 (N_9631,N_9238,N_9208);
nor U9632 (N_9632,N_9062,N_9495);
or U9633 (N_9633,N_9467,N_9449);
xor U9634 (N_9634,N_9255,N_9144);
xor U9635 (N_9635,N_9379,N_9488);
nand U9636 (N_9636,N_9473,N_9524);
and U9637 (N_9637,N_9283,N_9386);
nor U9638 (N_9638,N_9393,N_9445);
nor U9639 (N_9639,N_9207,N_9067);
and U9640 (N_9640,N_9021,N_9035);
and U9641 (N_9641,N_9149,N_9555);
and U9642 (N_9642,N_9214,N_9416);
nor U9643 (N_9643,N_9545,N_9222);
nand U9644 (N_9644,N_9582,N_9587);
and U9645 (N_9645,N_9378,N_9512);
or U9646 (N_9646,N_9167,N_9348);
nor U9647 (N_9647,N_9145,N_9562);
or U9648 (N_9648,N_9189,N_9529);
and U9649 (N_9649,N_9541,N_9499);
or U9650 (N_9650,N_9339,N_9330);
or U9651 (N_9651,N_9063,N_9150);
xor U9652 (N_9652,N_9369,N_9094);
nor U9653 (N_9653,N_9103,N_9522);
nand U9654 (N_9654,N_9256,N_9326);
nor U9655 (N_9655,N_9202,N_9458);
and U9656 (N_9656,N_9101,N_9082);
xnor U9657 (N_9657,N_9382,N_9195);
nand U9658 (N_9658,N_9277,N_9362);
nor U9659 (N_9659,N_9553,N_9209);
and U9660 (N_9660,N_9370,N_9480);
nand U9661 (N_9661,N_9459,N_9008);
nand U9662 (N_9662,N_9533,N_9053);
nor U9663 (N_9663,N_9590,N_9304);
xor U9664 (N_9664,N_9175,N_9430);
or U9665 (N_9665,N_9586,N_9285);
or U9666 (N_9666,N_9349,N_9039);
nor U9667 (N_9667,N_9092,N_9332);
nand U9668 (N_9668,N_9328,N_9388);
or U9669 (N_9669,N_9171,N_9452);
and U9670 (N_9670,N_9113,N_9177);
or U9671 (N_9671,N_9034,N_9598);
nand U9672 (N_9672,N_9197,N_9201);
or U9673 (N_9673,N_9414,N_9143);
or U9674 (N_9674,N_9276,N_9187);
or U9675 (N_9675,N_9407,N_9099);
or U9676 (N_9676,N_9069,N_9523);
and U9677 (N_9677,N_9341,N_9042);
nand U9678 (N_9678,N_9482,N_9337);
or U9679 (N_9679,N_9454,N_9278);
and U9680 (N_9680,N_9544,N_9002);
and U9681 (N_9681,N_9243,N_9227);
or U9682 (N_9682,N_9073,N_9474);
nor U9683 (N_9683,N_9287,N_9000);
or U9684 (N_9684,N_9051,N_9212);
nand U9685 (N_9685,N_9060,N_9329);
nor U9686 (N_9686,N_9122,N_9258);
nand U9687 (N_9687,N_9447,N_9153);
nand U9688 (N_9688,N_9525,N_9155);
or U9689 (N_9689,N_9134,N_9216);
and U9690 (N_9690,N_9185,N_9123);
nand U9691 (N_9691,N_9374,N_9096);
xor U9692 (N_9692,N_9270,N_9147);
and U9693 (N_9693,N_9041,N_9272);
nand U9694 (N_9694,N_9316,N_9429);
nand U9695 (N_9695,N_9117,N_9302);
xnor U9696 (N_9696,N_9336,N_9342);
nor U9697 (N_9697,N_9050,N_9478);
nor U9698 (N_9698,N_9074,N_9088);
nand U9699 (N_9699,N_9440,N_9353);
nor U9700 (N_9700,N_9136,N_9457);
nand U9701 (N_9701,N_9229,N_9210);
xor U9702 (N_9702,N_9223,N_9335);
and U9703 (N_9703,N_9496,N_9508);
or U9704 (N_9704,N_9059,N_9260);
or U9705 (N_9705,N_9427,N_9161);
nand U9706 (N_9706,N_9567,N_9006);
and U9707 (N_9707,N_9292,N_9133);
or U9708 (N_9708,N_9232,N_9599);
and U9709 (N_9709,N_9425,N_9048);
or U9710 (N_9710,N_9466,N_9104);
nand U9711 (N_9711,N_9400,N_9105);
nor U9712 (N_9712,N_9444,N_9291);
or U9713 (N_9713,N_9493,N_9472);
or U9714 (N_9714,N_9191,N_9084);
xnor U9715 (N_9715,N_9471,N_9286);
nand U9716 (N_9716,N_9593,N_9098);
nand U9717 (N_9717,N_9160,N_9317);
nor U9718 (N_9718,N_9019,N_9477);
nand U9719 (N_9719,N_9213,N_9079);
nor U9720 (N_9720,N_9519,N_9266);
nor U9721 (N_9721,N_9583,N_9417);
or U9722 (N_9722,N_9234,N_9220);
nand U9723 (N_9723,N_9170,N_9356);
nor U9724 (N_9724,N_9281,N_9078);
and U9725 (N_9725,N_9164,N_9237);
nand U9726 (N_9726,N_9033,N_9426);
nor U9727 (N_9727,N_9254,N_9262);
or U9728 (N_9728,N_9575,N_9455);
nand U9729 (N_9729,N_9020,N_9040);
or U9730 (N_9730,N_9148,N_9183);
nor U9731 (N_9731,N_9494,N_9433);
or U9732 (N_9732,N_9100,N_9072);
or U9733 (N_9733,N_9556,N_9180);
or U9734 (N_9734,N_9346,N_9456);
nor U9735 (N_9735,N_9413,N_9279);
nor U9736 (N_9736,N_9125,N_9569);
and U9737 (N_9737,N_9421,N_9225);
nand U9738 (N_9738,N_9131,N_9398);
and U9739 (N_9739,N_9244,N_9536);
and U9740 (N_9740,N_9158,N_9001);
nand U9741 (N_9741,N_9184,N_9594);
and U9742 (N_9742,N_9132,N_9230);
and U9743 (N_9743,N_9166,N_9313);
or U9744 (N_9744,N_9355,N_9547);
or U9745 (N_9745,N_9505,N_9319);
and U9746 (N_9746,N_9137,N_9010);
nor U9747 (N_9747,N_9247,N_9340);
and U9748 (N_9748,N_9200,N_9592);
nor U9749 (N_9749,N_9085,N_9057);
or U9750 (N_9750,N_9030,N_9299);
nor U9751 (N_9751,N_9566,N_9199);
nor U9752 (N_9752,N_9306,N_9242);
or U9753 (N_9753,N_9475,N_9595);
and U9754 (N_9754,N_9383,N_9024);
nor U9755 (N_9755,N_9294,N_9361);
nor U9756 (N_9756,N_9596,N_9463);
nor U9757 (N_9757,N_9215,N_9441);
nand U9758 (N_9758,N_9561,N_9365);
and U9759 (N_9759,N_9481,N_9129);
nor U9760 (N_9760,N_9106,N_9432);
nor U9761 (N_9761,N_9469,N_9570);
nand U9762 (N_9762,N_9387,N_9343);
or U9763 (N_9763,N_9080,N_9141);
nand U9764 (N_9764,N_9087,N_9597);
nand U9765 (N_9765,N_9004,N_9363);
or U9766 (N_9766,N_9465,N_9364);
nand U9767 (N_9767,N_9064,N_9403);
and U9768 (N_9768,N_9284,N_9376);
and U9769 (N_9769,N_9511,N_9288);
or U9770 (N_9770,N_9314,N_9504);
nand U9771 (N_9771,N_9322,N_9211);
nor U9772 (N_9772,N_9193,N_9172);
or U9773 (N_9773,N_9509,N_9435);
and U9774 (N_9774,N_9576,N_9240);
and U9775 (N_9775,N_9498,N_9239);
nor U9776 (N_9776,N_9483,N_9380);
and U9777 (N_9777,N_9253,N_9394);
or U9778 (N_9778,N_9521,N_9589);
or U9779 (N_9779,N_9401,N_9579);
nand U9780 (N_9780,N_9018,N_9071);
nand U9781 (N_9781,N_9282,N_9357);
and U9782 (N_9782,N_9036,N_9527);
nand U9783 (N_9783,N_9205,N_9419);
xnor U9784 (N_9784,N_9162,N_9151);
nand U9785 (N_9785,N_9520,N_9486);
nand U9786 (N_9786,N_9516,N_9194);
nand U9787 (N_9787,N_9052,N_9138);
nand U9788 (N_9788,N_9537,N_9017);
or U9789 (N_9789,N_9289,N_9502);
or U9790 (N_9790,N_9535,N_9146);
nor U9791 (N_9791,N_9182,N_9054);
nor U9792 (N_9792,N_9091,N_9577);
nor U9793 (N_9793,N_9275,N_9076);
and U9794 (N_9794,N_9565,N_9470);
or U9795 (N_9795,N_9462,N_9489);
and U9796 (N_9796,N_9464,N_9007);
and U9797 (N_9797,N_9070,N_9165);
and U9798 (N_9798,N_9381,N_9038);
and U9799 (N_9799,N_9043,N_9178);
and U9800 (N_9800,N_9204,N_9461);
and U9801 (N_9801,N_9028,N_9298);
or U9802 (N_9802,N_9246,N_9373);
nand U9803 (N_9803,N_9026,N_9551);
and U9804 (N_9804,N_9320,N_9485);
and U9805 (N_9805,N_9395,N_9118);
nand U9806 (N_9806,N_9308,N_9399);
nor U9807 (N_9807,N_9245,N_9557);
or U9808 (N_9808,N_9573,N_9190);
and U9809 (N_9809,N_9515,N_9089);
nand U9810 (N_9810,N_9174,N_9046);
and U9811 (N_9811,N_9497,N_9491);
and U9812 (N_9812,N_9154,N_9108);
and U9813 (N_9813,N_9179,N_9415);
nand U9814 (N_9814,N_9251,N_9492);
xnor U9815 (N_9815,N_9115,N_9114);
or U9816 (N_9816,N_9517,N_9448);
and U9817 (N_9817,N_9186,N_9152);
or U9818 (N_9818,N_9305,N_9003);
and U9819 (N_9819,N_9259,N_9542);
nor U9820 (N_9820,N_9241,N_9249);
and U9821 (N_9821,N_9109,N_9442);
nor U9822 (N_9822,N_9181,N_9031);
or U9823 (N_9823,N_9044,N_9083);
or U9824 (N_9824,N_9127,N_9418);
or U9825 (N_9825,N_9271,N_9501);
or U9826 (N_9826,N_9236,N_9264);
or U9827 (N_9827,N_9588,N_9368);
nor U9828 (N_9828,N_9410,N_9324);
nand U9829 (N_9829,N_9546,N_9090);
and U9830 (N_9830,N_9409,N_9333);
nor U9831 (N_9831,N_9102,N_9163);
nor U9832 (N_9832,N_9450,N_9273);
nor U9833 (N_9833,N_9408,N_9173);
nor U9834 (N_9834,N_9268,N_9309);
or U9835 (N_9835,N_9110,N_9011);
nand U9836 (N_9836,N_9086,N_9358);
and U9837 (N_9837,N_9530,N_9121);
or U9838 (N_9838,N_9584,N_9029);
and U9839 (N_9839,N_9434,N_9534);
and U9840 (N_9840,N_9295,N_9297);
xor U9841 (N_9841,N_9027,N_9518);
and U9842 (N_9842,N_9371,N_9124);
or U9843 (N_9843,N_9140,N_9428);
and U9844 (N_9844,N_9331,N_9228);
or U9845 (N_9845,N_9261,N_9206);
nand U9846 (N_9846,N_9157,N_9300);
and U9847 (N_9847,N_9350,N_9490);
or U9848 (N_9848,N_9301,N_9119);
or U9849 (N_9849,N_9221,N_9476);
nand U9850 (N_9850,N_9487,N_9159);
and U9851 (N_9851,N_9564,N_9438);
or U9852 (N_9852,N_9568,N_9005);
and U9853 (N_9853,N_9142,N_9531);
nor U9854 (N_9854,N_9397,N_9390);
and U9855 (N_9855,N_9338,N_9460);
or U9856 (N_9856,N_9218,N_9540);
nor U9857 (N_9857,N_9559,N_9549);
or U9858 (N_9858,N_9367,N_9274);
or U9859 (N_9859,N_9312,N_9112);
nor U9860 (N_9860,N_9436,N_9422);
or U9861 (N_9861,N_9558,N_9023);
and U9862 (N_9862,N_9049,N_9404);
or U9863 (N_9863,N_9280,N_9265);
and U9864 (N_9864,N_9226,N_9510);
or U9865 (N_9865,N_9075,N_9437);
nor U9866 (N_9866,N_9347,N_9095);
or U9867 (N_9867,N_9543,N_9296);
nand U9868 (N_9868,N_9116,N_9571);
nor U9869 (N_9869,N_9269,N_9318);
nor U9870 (N_9870,N_9248,N_9412);
and U9871 (N_9871,N_9446,N_9375);
and U9872 (N_9872,N_9231,N_9107);
nor U9873 (N_9873,N_9423,N_9484);
and U9874 (N_9874,N_9065,N_9217);
or U9875 (N_9875,N_9188,N_9514);
nand U9876 (N_9876,N_9013,N_9235);
or U9877 (N_9877,N_9548,N_9093);
nand U9878 (N_9878,N_9344,N_9574);
nor U9879 (N_9879,N_9552,N_9135);
and U9880 (N_9880,N_9267,N_9016);
or U9881 (N_9881,N_9351,N_9120);
and U9882 (N_9882,N_9058,N_9128);
nand U9883 (N_9883,N_9411,N_9126);
nor U9884 (N_9884,N_9354,N_9578);
nand U9885 (N_9885,N_9468,N_9290);
nand U9886 (N_9886,N_9402,N_9219);
nor U9887 (N_9887,N_9554,N_9532);
and U9888 (N_9888,N_9479,N_9015);
and U9889 (N_9889,N_9372,N_9539);
nor U9890 (N_9890,N_9431,N_9591);
nor U9891 (N_9891,N_9037,N_9528);
nand U9892 (N_9892,N_9250,N_9022);
xor U9893 (N_9893,N_9293,N_9526);
and U9894 (N_9894,N_9360,N_9585);
nor U9895 (N_9895,N_9025,N_9334);
nand U9896 (N_9896,N_9055,N_9538);
and U9897 (N_9897,N_9315,N_9077);
and U9898 (N_9898,N_9014,N_9420);
nor U9899 (N_9899,N_9550,N_9303);
and U9900 (N_9900,N_9016,N_9468);
nor U9901 (N_9901,N_9334,N_9543);
and U9902 (N_9902,N_9519,N_9440);
xnor U9903 (N_9903,N_9448,N_9301);
or U9904 (N_9904,N_9539,N_9307);
nand U9905 (N_9905,N_9004,N_9320);
nor U9906 (N_9906,N_9153,N_9543);
or U9907 (N_9907,N_9442,N_9577);
or U9908 (N_9908,N_9184,N_9449);
and U9909 (N_9909,N_9401,N_9260);
and U9910 (N_9910,N_9459,N_9437);
nand U9911 (N_9911,N_9220,N_9131);
nor U9912 (N_9912,N_9022,N_9206);
and U9913 (N_9913,N_9378,N_9224);
nor U9914 (N_9914,N_9074,N_9322);
nand U9915 (N_9915,N_9154,N_9451);
or U9916 (N_9916,N_9103,N_9052);
nand U9917 (N_9917,N_9280,N_9548);
nand U9918 (N_9918,N_9330,N_9522);
xor U9919 (N_9919,N_9479,N_9456);
nand U9920 (N_9920,N_9375,N_9037);
nor U9921 (N_9921,N_9030,N_9364);
nor U9922 (N_9922,N_9213,N_9013);
nor U9923 (N_9923,N_9109,N_9595);
or U9924 (N_9924,N_9239,N_9406);
xnor U9925 (N_9925,N_9189,N_9384);
nand U9926 (N_9926,N_9211,N_9294);
nand U9927 (N_9927,N_9370,N_9113);
nand U9928 (N_9928,N_9562,N_9418);
and U9929 (N_9929,N_9092,N_9493);
xor U9930 (N_9930,N_9574,N_9294);
or U9931 (N_9931,N_9058,N_9262);
and U9932 (N_9932,N_9447,N_9114);
nand U9933 (N_9933,N_9549,N_9379);
or U9934 (N_9934,N_9194,N_9138);
nand U9935 (N_9935,N_9496,N_9018);
nor U9936 (N_9936,N_9430,N_9045);
nor U9937 (N_9937,N_9164,N_9530);
nand U9938 (N_9938,N_9439,N_9243);
nand U9939 (N_9939,N_9309,N_9190);
nor U9940 (N_9940,N_9436,N_9245);
or U9941 (N_9941,N_9485,N_9026);
and U9942 (N_9942,N_9321,N_9144);
nor U9943 (N_9943,N_9096,N_9105);
nor U9944 (N_9944,N_9289,N_9546);
and U9945 (N_9945,N_9327,N_9575);
and U9946 (N_9946,N_9006,N_9370);
and U9947 (N_9947,N_9184,N_9222);
and U9948 (N_9948,N_9157,N_9520);
nor U9949 (N_9949,N_9156,N_9434);
nand U9950 (N_9950,N_9109,N_9072);
nor U9951 (N_9951,N_9236,N_9474);
or U9952 (N_9952,N_9463,N_9598);
and U9953 (N_9953,N_9186,N_9522);
nand U9954 (N_9954,N_9206,N_9353);
nand U9955 (N_9955,N_9144,N_9469);
or U9956 (N_9956,N_9235,N_9474);
and U9957 (N_9957,N_9435,N_9564);
nor U9958 (N_9958,N_9328,N_9561);
nand U9959 (N_9959,N_9000,N_9246);
and U9960 (N_9960,N_9379,N_9113);
nor U9961 (N_9961,N_9231,N_9406);
or U9962 (N_9962,N_9241,N_9554);
and U9963 (N_9963,N_9156,N_9523);
and U9964 (N_9964,N_9547,N_9046);
nand U9965 (N_9965,N_9387,N_9468);
or U9966 (N_9966,N_9280,N_9224);
and U9967 (N_9967,N_9304,N_9239);
and U9968 (N_9968,N_9251,N_9514);
or U9969 (N_9969,N_9360,N_9467);
or U9970 (N_9970,N_9127,N_9381);
or U9971 (N_9971,N_9393,N_9474);
nand U9972 (N_9972,N_9364,N_9131);
and U9973 (N_9973,N_9470,N_9355);
nor U9974 (N_9974,N_9298,N_9445);
and U9975 (N_9975,N_9495,N_9466);
nor U9976 (N_9976,N_9550,N_9397);
nand U9977 (N_9977,N_9138,N_9214);
nand U9978 (N_9978,N_9074,N_9057);
and U9979 (N_9979,N_9568,N_9598);
nand U9980 (N_9980,N_9557,N_9163);
and U9981 (N_9981,N_9485,N_9175);
nor U9982 (N_9982,N_9530,N_9234);
and U9983 (N_9983,N_9525,N_9589);
nand U9984 (N_9984,N_9556,N_9360);
nand U9985 (N_9985,N_9572,N_9204);
or U9986 (N_9986,N_9276,N_9192);
nand U9987 (N_9987,N_9532,N_9180);
and U9988 (N_9988,N_9045,N_9507);
nand U9989 (N_9989,N_9111,N_9207);
nand U9990 (N_9990,N_9120,N_9138);
nand U9991 (N_9991,N_9067,N_9325);
or U9992 (N_9992,N_9014,N_9403);
nor U9993 (N_9993,N_9572,N_9486);
nor U9994 (N_9994,N_9098,N_9205);
and U9995 (N_9995,N_9262,N_9232);
or U9996 (N_9996,N_9249,N_9133);
nor U9997 (N_9997,N_9194,N_9452);
and U9998 (N_9998,N_9565,N_9195);
nand U9999 (N_9999,N_9329,N_9241);
xnor U10000 (N_10000,N_9062,N_9203);
nand U10001 (N_10001,N_9442,N_9352);
nand U10002 (N_10002,N_9352,N_9484);
or U10003 (N_10003,N_9399,N_9339);
and U10004 (N_10004,N_9007,N_9164);
and U10005 (N_10005,N_9340,N_9035);
and U10006 (N_10006,N_9071,N_9281);
and U10007 (N_10007,N_9037,N_9093);
or U10008 (N_10008,N_9313,N_9119);
or U10009 (N_10009,N_9144,N_9429);
and U10010 (N_10010,N_9436,N_9234);
xnor U10011 (N_10011,N_9560,N_9074);
nor U10012 (N_10012,N_9437,N_9338);
or U10013 (N_10013,N_9266,N_9162);
nor U10014 (N_10014,N_9464,N_9246);
xor U10015 (N_10015,N_9250,N_9152);
nand U10016 (N_10016,N_9327,N_9563);
and U10017 (N_10017,N_9123,N_9434);
and U10018 (N_10018,N_9449,N_9198);
xor U10019 (N_10019,N_9079,N_9010);
nand U10020 (N_10020,N_9460,N_9381);
or U10021 (N_10021,N_9573,N_9055);
nand U10022 (N_10022,N_9558,N_9412);
or U10023 (N_10023,N_9023,N_9030);
and U10024 (N_10024,N_9372,N_9023);
or U10025 (N_10025,N_9176,N_9279);
or U10026 (N_10026,N_9496,N_9205);
nand U10027 (N_10027,N_9377,N_9584);
nor U10028 (N_10028,N_9202,N_9484);
nor U10029 (N_10029,N_9062,N_9261);
or U10030 (N_10030,N_9347,N_9233);
nor U10031 (N_10031,N_9518,N_9469);
nor U10032 (N_10032,N_9080,N_9496);
nor U10033 (N_10033,N_9585,N_9543);
nand U10034 (N_10034,N_9452,N_9252);
nor U10035 (N_10035,N_9471,N_9070);
nor U10036 (N_10036,N_9276,N_9471);
and U10037 (N_10037,N_9152,N_9597);
and U10038 (N_10038,N_9504,N_9246);
xnor U10039 (N_10039,N_9572,N_9046);
nor U10040 (N_10040,N_9028,N_9187);
nor U10041 (N_10041,N_9413,N_9457);
and U10042 (N_10042,N_9475,N_9096);
nand U10043 (N_10043,N_9429,N_9381);
nand U10044 (N_10044,N_9558,N_9144);
xor U10045 (N_10045,N_9438,N_9097);
nor U10046 (N_10046,N_9026,N_9125);
nand U10047 (N_10047,N_9518,N_9403);
and U10048 (N_10048,N_9477,N_9470);
nand U10049 (N_10049,N_9315,N_9551);
and U10050 (N_10050,N_9446,N_9425);
nor U10051 (N_10051,N_9479,N_9227);
or U10052 (N_10052,N_9061,N_9223);
nor U10053 (N_10053,N_9595,N_9042);
or U10054 (N_10054,N_9288,N_9314);
or U10055 (N_10055,N_9493,N_9555);
and U10056 (N_10056,N_9024,N_9330);
nor U10057 (N_10057,N_9162,N_9063);
xnor U10058 (N_10058,N_9061,N_9100);
or U10059 (N_10059,N_9239,N_9519);
or U10060 (N_10060,N_9250,N_9477);
nand U10061 (N_10061,N_9274,N_9407);
xnor U10062 (N_10062,N_9384,N_9322);
nor U10063 (N_10063,N_9280,N_9523);
nor U10064 (N_10064,N_9109,N_9087);
nand U10065 (N_10065,N_9064,N_9314);
xor U10066 (N_10066,N_9140,N_9211);
or U10067 (N_10067,N_9187,N_9371);
and U10068 (N_10068,N_9514,N_9265);
nor U10069 (N_10069,N_9196,N_9596);
and U10070 (N_10070,N_9001,N_9576);
or U10071 (N_10071,N_9403,N_9093);
nor U10072 (N_10072,N_9490,N_9387);
and U10073 (N_10073,N_9172,N_9313);
nor U10074 (N_10074,N_9296,N_9312);
nor U10075 (N_10075,N_9186,N_9586);
or U10076 (N_10076,N_9098,N_9223);
and U10077 (N_10077,N_9175,N_9060);
and U10078 (N_10078,N_9245,N_9002);
or U10079 (N_10079,N_9476,N_9274);
or U10080 (N_10080,N_9217,N_9326);
nand U10081 (N_10081,N_9546,N_9561);
and U10082 (N_10082,N_9266,N_9121);
and U10083 (N_10083,N_9393,N_9121);
and U10084 (N_10084,N_9503,N_9337);
nor U10085 (N_10085,N_9299,N_9455);
nand U10086 (N_10086,N_9525,N_9322);
and U10087 (N_10087,N_9286,N_9298);
nand U10088 (N_10088,N_9357,N_9511);
and U10089 (N_10089,N_9103,N_9001);
or U10090 (N_10090,N_9453,N_9401);
and U10091 (N_10091,N_9536,N_9522);
or U10092 (N_10092,N_9474,N_9509);
and U10093 (N_10093,N_9070,N_9251);
nand U10094 (N_10094,N_9560,N_9309);
nand U10095 (N_10095,N_9101,N_9234);
nor U10096 (N_10096,N_9378,N_9128);
nor U10097 (N_10097,N_9486,N_9443);
or U10098 (N_10098,N_9039,N_9453);
nand U10099 (N_10099,N_9284,N_9572);
and U10100 (N_10100,N_9180,N_9485);
nor U10101 (N_10101,N_9534,N_9077);
or U10102 (N_10102,N_9137,N_9310);
nor U10103 (N_10103,N_9025,N_9055);
nor U10104 (N_10104,N_9157,N_9485);
nand U10105 (N_10105,N_9184,N_9593);
nor U10106 (N_10106,N_9264,N_9528);
or U10107 (N_10107,N_9208,N_9094);
and U10108 (N_10108,N_9116,N_9201);
or U10109 (N_10109,N_9461,N_9219);
and U10110 (N_10110,N_9056,N_9322);
nand U10111 (N_10111,N_9145,N_9484);
nor U10112 (N_10112,N_9530,N_9037);
nand U10113 (N_10113,N_9445,N_9344);
and U10114 (N_10114,N_9191,N_9152);
and U10115 (N_10115,N_9205,N_9232);
or U10116 (N_10116,N_9444,N_9147);
nand U10117 (N_10117,N_9439,N_9055);
nor U10118 (N_10118,N_9226,N_9370);
nand U10119 (N_10119,N_9315,N_9308);
nand U10120 (N_10120,N_9481,N_9261);
nor U10121 (N_10121,N_9321,N_9008);
or U10122 (N_10122,N_9347,N_9507);
and U10123 (N_10123,N_9495,N_9268);
and U10124 (N_10124,N_9527,N_9157);
xor U10125 (N_10125,N_9107,N_9166);
nand U10126 (N_10126,N_9378,N_9235);
or U10127 (N_10127,N_9043,N_9432);
nand U10128 (N_10128,N_9002,N_9191);
or U10129 (N_10129,N_9396,N_9569);
nor U10130 (N_10130,N_9455,N_9366);
nor U10131 (N_10131,N_9116,N_9590);
nand U10132 (N_10132,N_9146,N_9255);
or U10133 (N_10133,N_9428,N_9332);
nand U10134 (N_10134,N_9337,N_9468);
xor U10135 (N_10135,N_9176,N_9410);
nand U10136 (N_10136,N_9454,N_9033);
nor U10137 (N_10137,N_9072,N_9409);
or U10138 (N_10138,N_9421,N_9531);
nor U10139 (N_10139,N_9206,N_9464);
or U10140 (N_10140,N_9450,N_9519);
and U10141 (N_10141,N_9018,N_9480);
and U10142 (N_10142,N_9090,N_9164);
nand U10143 (N_10143,N_9532,N_9490);
or U10144 (N_10144,N_9454,N_9017);
nor U10145 (N_10145,N_9425,N_9526);
and U10146 (N_10146,N_9140,N_9478);
and U10147 (N_10147,N_9259,N_9376);
nand U10148 (N_10148,N_9021,N_9360);
nor U10149 (N_10149,N_9298,N_9267);
nor U10150 (N_10150,N_9529,N_9567);
nor U10151 (N_10151,N_9592,N_9037);
xnor U10152 (N_10152,N_9095,N_9205);
nor U10153 (N_10153,N_9003,N_9195);
nor U10154 (N_10154,N_9038,N_9279);
or U10155 (N_10155,N_9172,N_9116);
nand U10156 (N_10156,N_9102,N_9059);
xnor U10157 (N_10157,N_9136,N_9382);
and U10158 (N_10158,N_9024,N_9193);
nor U10159 (N_10159,N_9306,N_9299);
or U10160 (N_10160,N_9575,N_9100);
xor U10161 (N_10161,N_9002,N_9065);
nor U10162 (N_10162,N_9049,N_9072);
or U10163 (N_10163,N_9367,N_9590);
nor U10164 (N_10164,N_9578,N_9182);
and U10165 (N_10165,N_9123,N_9292);
and U10166 (N_10166,N_9118,N_9183);
nor U10167 (N_10167,N_9046,N_9522);
or U10168 (N_10168,N_9438,N_9345);
nand U10169 (N_10169,N_9311,N_9419);
or U10170 (N_10170,N_9126,N_9211);
and U10171 (N_10171,N_9391,N_9494);
nor U10172 (N_10172,N_9070,N_9456);
or U10173 (N_10173,N_9442,N_9506);
and U10174 (N_10174,N_9228,N_9354);
nor U10175 (N_10175,N_9449,N_9579);
nand U10176 (N_10176,N_9413,N_9412);
nor U10177 (N_10177,N_9028,N_9220);
or U10178 (N_10178,N_9092,N_9127);
or U10179 (N_10179,N_9580,N_9288);
or U10180 (N_10180,N_9573,N_9540);
or U10181 (N_10181,N_9299,N_9531);
nand U10182 (N_10182,N_9366,N_9311);
nand U10183 (N_10183,N_9102,N_9397);
or U10184 (N_10184,N_9550,N_9445);
and U10185 (N_10185,N_9594,N_9560);
nand U10186 (N_10186,N_9061,N_9167);
or U10187 (N_10187,N_9324,N_9027);
nor U10188 (N_10188,N_9474,N_9407);
and U10189 (N_10189,N_9030,N_9418);
nand U10190 (N_10190,N_9298,N_9528);
or U10191 (N_10191,N_9233,N_9020);
nor U10192 (N_10192,N_9204,N_9241);
nor U10193 (N_10193,N_9251,N_9196);
nor U10194 (N_10194,N_9174,N_9413);
nand U10195 (N_10195,N_9159,N_9109);
nor U10196 (N_10196,N_9390,N_9164);
and U10197 (N_10197,N_9364,N_9139);
nor U10198 (N_10198,N_9195,N_9521);
or U10199 (N_10199,N_9146,N_9187);
and U10200 (N_10200,N_10168,N_9793);
nor U10201 (N_10201,N_9818,N_10071);
nand U10202 (N_10202,N_9707,N_10132);
or U10203 (N_10203,N_10166,N_9980);
nand U10204 (N_10204,N_10064,N_9758);
and U10205 (N_10205,N_10159,N_9735);
nand U10206 (N_10206,N_9892,N_9757);
and U10207 (N_10207,N_9846,N_9831);
or U10208 (N_10208,N_9690,N_9950);
nand U10209 (N_10209,N_9619,N_9745);
nand U10210 (N_10210,N_9863,N_9645);
nand U10211 (N_10211,N_9905,N_9605);
nor U10212 (N_10212,N_9736,N_10076);
and U10213 (N_10213,N_10155,N_9672);
nor U10214 (N_10214,N_9934,N_9855);
nand U10215 (N_10215,N_10023,N_9897);
nor U10216 (N_10216,N_9938,N_9865);
nand U10217 (N_10217,N_9716,N_9877);
and U10218 (N_10218,N_9723,N_10034);
or U10219 (N_10219,N_10014,N_10192);
and U10220 (N_10220,N_9643,N_10114);
nor U10221 (N_10221,N_9812,N_9906);
xor U10222 (N_10222,N_9623,N_10086);
and U10223 (N_10223,N_9648,N_9658);
or U10224 (N_10224,N_10189,N_9652);
xor U10225 (N_10225,N_9967,N_9894);
nand U10226 (N_10226,N_9771,N_9767);
and U10227 (N_10227,N_9978,N_9805);
or U10228 (N_10228,N_10121,N_10025);
or U10229 (N_10229,N_10158,N_9965);
nor U10230 (N_10230,N_10108,N_9669);
nand U10231 (N_10231,N_9610,N_9824);
nor U10232 (N_10232,N_10089,N_9974);
and U10233 (N_10233,N_9816,N_9659);
or U10234 (N_10234,N_9917,N_9712);
or U10235 (N_10235,N_9751,N_9976);
and U10236 (N_10236,N_9910,N_10184);
or U10237 (N_10237,N_9715,N_9692);
and U10238 (N_10238,N_9674,N_10117);
or U10239 (N_10239,N_9786,N_9656);
and U10240 (N_10240,N_10091,N_9624);
and U10241 (N_10241,N_9809,N_10165);
nor U10242 (N_10242,N_10107,N_9999);
nand U10243 (N_10243,N_10163,N_10171);
or U10244 (N_10244,N_9807,N_9673);
nand U10245 (N_10245,N_9922,N_10077);
and U10246 (N_10246,N_9891,N_9979);
nand U10247 (N_10247,N_10126,N_10142);
and U10248 (N_10248,N_10120,N_9682);
and U10249 (N_10249,N_9823,N_10161);
and U10250 (N_10250,N_10138,N_10179);
or U10251 (N_10251,N_10004,N_9700);
and U10252 (N_10252,N_10026,N_10090);
nand U10253 (N_10253,N_10024,N_9691);
or U10254 (N_10254,N_9677,N_9622);
nand U10255 (N_10255,N_9798,N_9861);
nor U10256 (N_10256,N_10147,N_9954);
nand U10257 (N_10257,N_9731,N_9803);
nand U10258 (N_10258,N_9890,N_9729);
nand U10259 (N_10259,N_10104,N_10035);
nand U10260 (N_10260,N_10151,N_9653);
nand U10261 (N_10261,N_10122,N_9627);
or U10262 (N_10262,N_10083,N_10154);
nor U10263 (N_10263,N_10055,N_10041);
nor U10264 (N_10264,N_9969,N_9843);
nand U10265 (N_10265,N_10016,N_10139);
nand U10266 (N_10266,N_9740,N_10169);
nor U10267 (N_10267,N_9832,N_9882);
or U10268 (N_10268,N_9949,N_9693);
nor U10269 (N_10269,N_9956,N_10020);
nand U10270 (N_10270,N_10198,N_9960);
nand U10271 (N_10271,N_9998,N_10186);
nor U10272 (N_10272,N_9900,N_9788);
nor U10273 (N_10273,N_9744,N_9935);
or U10274 (N_10274,N_9628,N_10075);
nor U10275 (N_10275,N_9721,N_10141);
nand U10276 (N_10276,N_10029,N_10058);
or U10277 (N_10277,N_10042,N_10000);
nor U10278 (N_10278,N_10053,N_9981);
or U10279 (N_10279,N_10196,N_10033);
nand U10280 (N_10280,N_9872,N_9738);
or U10281 (N_10281,N_9601,N_9792);
or U10282 (N_10282,N_9837,N_10017);
nand U10283 (N_10283,N_9940,N_9631);
nand U10284 (N_10284,N_10173,N_9613);
nand U10285 (N_10285,N_9774,N_9884);
nand U10286 (N_10286,N_9849,N_9930);
and U10287 (N_10287,N_10005,N_10145);
or U10288 (N_10288,N_9985,N_10148);
xnor U10289 (N_10289,N_10194,N_9853);
nand U10290 (N_10290,N_10109,N_10134);
and U10291 (N_10291,N_9703,N_9748);
nand U10292 (N_10292,N_10123,N_9795);
and U10293 (N_10293,N_9991,N_9914);
nor U10294 (N_10294,N_9880,N_9963);
nor U10295 (N_10295,N_9814,N_9983);
and U10296 (N_10296,N_9747,N_10150);
nor U10297 (N_10297,N_9870,N_10199);
nor U10298 (N_10298,N_9654,N_9944);
nor U10299 (N_10299,N_9763,N_10193);
or U10300 (N_10300,N_9862,N_9955);
or U10301 (N_10301,N_10146,N_9676);
xor U10302 (N_10302,N_9923,N_9995);
nor U10303 (N_10303,N_9663,N_9859);
and U10304 (N_10304,N_9777,N_9724);
or U10305 (N_10305,N_9603,N_10183);
and U10306 (N_10306,N_9947,N_9706);
nor U10307 (N_10307,N_10197,N_9615);
nor U10308 (N_10308,N_10097,N_9951);
nor U10309 (N_10309,N_9925,N_10054);
and U10310 (N_10310,N_9835,N_9994);
or U10311 (N_10311,N_9667,N_9699);
nor U10312 (N_10312,N_10012,N_9889);
and U10313 (N_10313,N_9679,N_10111);
or U10314 (N_10314,N_9684,N_9946);
or U10315 (N_10315,N_10060,N_9651);
nor U10316 (N_10316,N_9698,N_10007);
nand U10317 (N_10317,N_9928,N_10073);
and U10318 (N_10318,N_10069,N_9604);
nor U10319 (N_10319,N_9752,N_9796);
xnor U10320 (N_10320,N_9866,N_10156);
nor U10321 (N_10321,N_9683,N_9834);
or U10322 (N_10322,N_9661,N_9687);
nor U10323 (N_10323,N_9778,N_10178);
nand U10324 (N_10324,N_9675,N_9813);
nand U10325 (N_10325,N_10018,N_10131);
and U10326 (N_10326,N_9990,N_9689);
and U10327 (N_10327,N_10043,N_10181);
or U10328 (N_10328,N_9638,N_9856);
and U10329 (N_10329,N_9694,N_9921);
nand U10330 (N_10330,N_10125,N_10099);
and U10331 (N_10331,N_9657,N_10038);
nor U10332 (N_10332,N_9907,N_9727);
or U10333 (N_10333,N_10037,N_9898);
and U10334 (N_10334,N_9948,N_9895);
or U10335 (N_10335,N_9739,N_9953);
and U10336 (N_10336,N_9769,N_9919);
and U10337 (N_10337,N_10092,N_9733);
nand U10338 (N_10338,N_10070,N_10068);
and U10339 (N_10339,N_9701,N_9918);
nand U10340 (N_10340,N_9819,N_9825);
or U10341 (N_10341,N_9810,N_9828);
and U10342 (N_10342,N_9732,N_10105);
or U10343 (N_10343,N_10157,N_9722);
or U10344 (N_10344,N_9696,N_9761);
nand U10345 (N_10345,N_10103,N_9743);
and U10346 (N_10346,N_9997,N_10002);
nand U10347 (N_10347,N_9867,N_9913);
nor U10348 (N_10348,N_10098,N_9992);
nand U10349 (N_10349,N_9620,N_9868);
and U10350 (N_10350,N_9650,N_10003);
nand U10351 (N_10351,N_9695,N_9776);
or U10352 (N_10352,N_9606,N_9876);
and U10353 (N_10353,N_9854,N_9886);
nor U10354 (N_10354,N_9647,N_9959);
nor U10355 (N_10355,N_9901,N_9878);
nor U10356 (N_10356,N_10074,N_10110);
or U10357 (N_10357,N_9885,N_9833);
nand U10358 (N_10358,N_10087,N_9726);
nor U10359 (N_10359,N_9713,N_9896);
and U10360 (N_10360,N_9931,N_9970);
nand U10361 (N_10361,N_9904,N_10160);
or U10362 (N_10362,N_10096,N_9857);
or U10363 (N_10363,N_9799,N_9830);
and U10364 (N_10364,N_9714,N_9759);
xor U10365 (N_10365,N_9639,N_9734);
nor U10366 (N_10366,N_9986,N_10119);
nor U10367 (N_10367,N_9626,N_9755);
and U10368 (N_10368,N_10032,N_9836);
nor U10369 (N_10369,N_9760,N_9847);
nand U10370 (N_10370,N_9987,N_9908);
and U10371 (N_10371,N_9742,N_9621);
nand U10372 (N_10372,N_9797,N_9660);
nor U10373 (N_10373,N_9893,N_9842);
nand U10374 (N_10374,N_9655,N_9929);
or U10375 (N_10375,N_10065,N_10066);
and U10376 (N_10376,N_9802,N_9887);
nand U10377 (N_10377,N_9617,N_10019);
and U10378 (N_10378,N_9800,N_10036);
and U10379 (N_10379,N_9822,N_9609);
and U10380 (N_10380,N_9753,N_9780);
nand U10381 (N_10381,N_10191,N_9789);
or U10382 (N_10382,N_10124,N_9964);
or U10383 (N_10383,N_10082,N_10028);
nand U10384 (N_10384,N_10078,N_10133);
nand U10385 (N_10385,N_9697,N_10116);
or U10386 (N_10386,N_9633,N_10009);
and U10387 (N_10387,N_10057,N_9750);
or U10388 (N_10388,N_10063,N_9879);
or U10389 (N_10389,N_9903,N_9844);
nand U10390 (N_10390,N_10011,N_9629);
or U10391 (N_10391,N_9971,N_9720);
and U10392 (N_10392,N_9746,N_9719);
nand U10393 (N_10393,N_9966,N_9612);
nor U10394 (N_10394,N_10048,N_10047);
nand U10395 (N_10395,N_10188,N_9749);
and U10396 (N_10396,N_9664,N_9791);
nor U10397 (N_10397,N_10031,N_9784);
nor U10398 (N_10398,N_9977,N_9984);
and U10399 (N_10399,N_9635,N_9730);
or U10400 (N_10400,N_10062,N_10079);
nand U10401 (N_10401,N_10006,N_10072);
or U10402 (N_10402,N_9709,N_10180);
and U10403 (N_10403,N_9634,N_9794);
or U10404 (N_10404,N_9899,N_9932);
nor U10405 (N_10405,N_10052,N_9718);
nor U10406 (N_10406,N_10044,N_9945);
nor U10407 (N_10407,N_9916,N_10021);
nand U10408 (N_10408,N_9768,N_10080);
nand U10409 (N_10409,N_9717,N_9827);
nor U10410 (N_10410,N_9937,N_10137);
and U10411 (N_10411,N_9787,N_9765);
nor U10412 (N_10412,N_9864,N_9616);
or U10413 (N_10413,N_9641,N_10101);
and U10414 (N_10414,N_9851,N_9808);
nand U10415 (N_10415,N_9871,N_9644);
xnor U10416 (N_10416,N_9972,N_10115);
xor U10417 (N_10417,N_9725,N_10050);
nand U10418 (N_10418,N_10176,N_10051);
nor U10419 (N_10419,N_9671,N_10084);
or U10420 (N_10420,N_10127,N_9640);
nor U10421 (N_10421,N_10001,N_9611);
nor U10422 (N_10422,N_10010,N_9936);
and U10423 (N_10423,N_9666,N_9820);
nand U10424 (N_10424,N_9702,N_9845);
or U10425 (N_10425,N_9630,N_9852);
nor U10426 (N_10426,N_9600,N_10022);
and U10427 (N_10427,N_9728,N_9873);
nor U10428 (N_10428,N_9710,N_10095);
nor U10429 (N_10429,N_9783,N_9762);
nor U10430 (N_10430,N_9614,N_9608);
nor U10431 (N_10431,N_10027,N_10175);
nand U10432 (N_10432,N_9662,N_9670);
and U10433 (N_10433,N_10135,N_9680);
or U10434 (N_10434,N_10046,N_10056);
and U10435 (N_10435,N_9607,N_9804);
nand U10436 (N_10436,N_9902,N_9962);
nand U10437 (N_10437,N_10102,N_10113);
nand U10438 (N_10438,N_10015,N_10094);
nor U10439 (N_10439,N_9642,N_9711);
and U10440 (N_10440,N_9915,N_9688);
nor U10441 (N_10441,N_9770,N_9975);
nand U10442 (N_10442,N_10130,N_9775);
nand U10443 (N_10443,N_10185,N_9961);
nand U10444 (N_10444,N_9829,N_9850);
or U10445 (N_10445,N_10177,N_9602);
or U10446 (N_10446,N_10149,N_9958);
nand U10447 (N_10447,N_9632,N_9826);
nand U10448 (N_10448,N_10182,N_9737);
or U10449 (N_10449,N_10195,N_9754);
nor U10450 (N_10450,N_9681,N_9705);
or U10451 (N_10451,N_9858,N_9649);
nand U10452 (N_10452,N_9646,N_9766);
and U10453 (N_10453,N_10030,N_9926);
nor U10454 (N_10454,N_10013,N_9665);
nand U10455 (N_10455,N_10153,N_10008);
nand U10456 (N_10456,N_9801,N_9912);
and U10457 (N_10457,N_9618,N_9772);
nand U10458 (N_10458,N_10136,N_10061);
and U10459 (N_10459,N_9957,N_10088);
or U10460 (N_10460,N_9848,N_9708);
nand U10461 (N_10461,N_10100,N_9941);
and U10462 (N_10462,N_10039,N_9785);
nand U10463 (N_10463,N_9875,N_10190);
and U10464 (N_10464,N_9909,N_9993);
and U10465 (N_10465,N_9815,N_9636);
nor U10466 (N_10466,N_10170,N_9790);
nand U10467 (N_10467,N_10085,N_9841);
nand U10468 (N_10468,N_10174,N_9781);
or U10469 (N_10469,N_9686,N_9773);
and U10470 (N_10470,N_9668,N_9939);
nor U10471 (N_10471,N_9704,N_9943);
nand U10472 (N_10472,N_9996,N_10093);
nand U10473 (N_10473,N_9911,N_9952);
or U10474 (N_10474,N_10167,N_10128);
nor U10475 (N_10475,N_9881,N_10106);
nor U10476 (N_10476,N_10164,N_9779);
nor U10477 (N_10477,N_10049,N_9883);
or U10478 (N_10478,N_10162,N_9927);
and U10479 (N_10479,N_10187,N_9888);
nand U10480 (N_10480,N_9988,N_9860);
or U10481 (N_10481,N_9973,N_10140);
nor U10482 (N_10482,N_10129,N_9989);
nor U10483 (N_10483,N_9840,N_10144);
nor U10484 (N_10484,N_10143,N_9685);
and U10485 (N_10485,N_9968,N_9806);
or U10486 (N_10486,N_9782,N_9924);
and U10487 (N_10487,N_10081,N_9869);
nand U10488 (N_10488,N_10067,N_10040);
nor U10489 (N_10489,N_9838,N_9625);
nand U10490 (N_10490,N_9756,N_9817);
or U10491 (N_10491,N_9678,N_10112);
nand U10492 (N_10492,N_9839,N_9821);
or U10493 (N_10493,N_10172,N_9637);
nor U10494 (N_10494,N_9920,N_9811);
nand U10495 (N_10495,N_9942,N_10059);
or U10496 (N_10496,N_9764,N_10118);
nor U10497 (N_10497,N_9982,N_9874);
xnor U10498 (N_10498,N_10045,N_9741);
nor U10499 (N_10499,N_10152,N_9933);
or U10500 (N_10500,N_10105,N_9958);
nor U10501 (N_10501,N_10176,N_9885);
nand U10502 (N_10502,N_9903,N_10129);
nand U10503 (N_10503,N_9986,N_9862);
and U10504 (N_10504,N_10137,N_9917);
nor U10505 (N_10505,N_10067,N_9628);
and U10506 (N_10506,N_10156,N_10067);
nor U10507 (N_10507,N_9801,N_10090);
nand U10508 (N_10508,N_10092,N_10143);
nor U10509 (N_10509,N_10190,N_10067);
and U10510 (N_10510,N_10095,N_10009);
and U10511 (N_10511,N_9713,N_9922);
nor U10512 (N_10512,N_10011,N_10157);
or U10513 (N_10513,N_9759,N_9633);
and U10514 (N_10514,N_10092,N_10173);
nand U10515 (N_10515,N_10068,N_10133);
and U10516 (N_10516,N_10052,N_9859);
nand U10517 (N_10517,N_9644,N_9853);
and U10518 (N_10518,N_9756,N_9889);
and U10519 (N_10519,N_9749,N_9878);
and U10520 (N_10520,N_10149,N_9890);
nand U10521 (N_10521,N_10040,N_9792);
and U10522 (N_10522,N_9855,N_9741);
nor U10523 (N_10523,N_9737,N_9958);
nor U10524 (N_10524,N_9879,N_10104);
nand U10525 (N_10525,N_9951,N_9995);
nand U10526 (N_10526,N_9623,N_9791);
and U10527 (N_10527,N_9669,N_9668);
nor U10528 (N_10528,N_10198,N_9931);
or U10529 (N_10529,N_9613,N_9849);
nor U10530 (N_10530,N_10051,N_9945);
nand U10531 (N_10531,N_9661,N_10149);
and U10532 (N_10532,N_10163,N_9667);
xor U10533 (N_10533,N_10130,N_9638);
or U10534 (N_10534,N_9837,N_9920);
nand U10535 (N_10535,N_9945,N_9848);
and U10536 (N_10536,N_10053,N_9653);
nand U10537 (N_10537,N_9720,N_10124);
xor U10538 (N_10538,N_10143,N_10097);
nor U10539 (N_10539,N_9905,N_10159);
and U10540 (N_10540,N_9985,N_10048);
or U10541 (N_10541,N_9765,N_10185);
nor U10542 (N_10542,N_10103,N_9863);
nand U10543 (N_10543,N_10142,N_9735);
and U10544 (N_10544,N_9830,N_9695);
nand U10545 (N_10545,N_9603,N_10017);
and U10546 (N_10546,N_9717,N_10085);
and U10547 (N_10547,N_9827,N_9766);
or U10548 (N_10548,N_9644,N_10179);
and U10549 (N_10549,N_9933,N_9957);
or U10550 (N_10550,N_10194,N_9990);
nor U10551 (N_10551,N_10172,N_9749);
nor U10552 (N_10552,N_9975,N_9651);
or U10553 (N_10553,N_9855,N_10060);
nor U10554 (N_10554,N_10083,N_10009);
and U10555 (N_10555,N_9962,N_10036);
and U10556 (N_10556,N_9623,N_9717);
nand U10557 (N_10557,N_10199,N_9617);
and U10558 (N_10558,N_9654,N_9914);
nand U10559 (N_10559,N_10045,N_9824);
nor U10560 (N_10560,N_9824,N_9640);
and U10561 (N_10561,N_9901,N_9602);
xnor U10562 (N_10562,N_10131,N_9744);
or U10563 (N_10563,N_9604,N_9676);
and U10564 (N_10564,N_9862,N_9664);
and U10565 (N_10565,N_10122,N_9766);
nand U10566 (N_10566,N_9794,N_9658);
nor U10567 (N_10567,N_10193,N_9660);
or U10568 (N_10568,N_9796,N_9942);
xnor U10569 (N_10569,N_9659,N_9670);
and U10570 (N_10570,N_10129,N_9610);
and U10571 (N_10571,N_9845,N_10074);
nor U10572 (N_10572,N_9826,N_10112);
or U10573 (N_10573,N_9964,N_10048);
nand U10574 (N_10574,N_10195,N_9617);
nor U10575 (N_10575,N_9602,N_9663);
and U10576 (N_10576,N_10052,N_9778);
and U10577 (N_10577,N_10060,N_9897);
nand U10578 (N_10578,N_9768,N_10031);
nand U10579 (N_10579,N_9986,N_10121);
or U10580 (N_10580,N_9715,N_9928);
nor U10581 (N_10581,N_9880,N_10160);
and U10582 (N_10582,N_9642,N_9805);
and U10583 (N_10583,N_9951,N_10129);
nor U10584 (N_10584,N_10145,N_9622);
or U10585 (N_10585,N_10152,N_9935);
xor U10586 (N_10586,N_9780,N_9602);
nand U10587 (N_10587,N_10175,N_9915);
nor U10588 (N_10588,N_9837,N_10178);
nor U10589 (N_10589,N_9992,N_9958);
and U10590 (N_10590,N_10163,N_9807);
nand U10591 (N_10591,N_10111,N_10123);
and U10592 (N_10592,N_9941,N_10172);
nand U10593 (N_10593,N_10168,N_10120);
nand U10594 (N_10594,N_10036,N_9760);
nand U10595 (N_10595,N_9827,N_10085);
or U10596 (N_10596,N_10087,N_9762);
nand U10597 (N_10597,N_9980,N_10065);
nor U10598 (N_10598,N_9739,N_9606);
nor U10599 (N_10599,N_10179,N_9900);
and U10600 (N_10600,N_9700,N_9849);
and U10601 (N_10601,N_9748,N_9989);
or U10602 (N_10602,N_9770,N_9898);
and U10603 (N_10603,N_9744,N_9746);
nand U10604 (N_10604,N_9728,N_9624);
and U10605 (N_10605,N_10093,N_9722);
nand U10606 (N_10606,N_9719,N_9944);
nor U10607 (N_10607,N_9830,N_9818);
or U10608 (N_10608,N_10010,N_9903);
nand U10609 (N_10609,N_10148,N_9953);
nand U10610 (N_10610,N_9780,N_9836);
nand U10611 (N_10611,N_9926,N_10191);
and U10612 (N_10612,N_9672,N_9620);
nand U10613 (N_10613,N_9844,N_10038);
nand U10614 (N_10614,N_9914,N_9973);
or U10615 (N_10615,N_9638,N_9603);
nand U10616 (N_10616,N_10188,N_9787);
or U10617 (N_10617,N_9634,N_10100);
nor U10618 (N_10618,N_9735,N_9930);
nor U10619 (N_10619,N_9614,N_9960);
nor U10620 (N_10620,N_9986,N_9738);
nor U10621 (N_10621,N_10112,N_10104);
nor U10622 (N_10622,N_9712,N_9976);
or U10623 (N_10623,N_9964,N_10043);
nor U10624 (N_10624,N_9665,N_9779);
nor U10625 (N_10625,N_10010,N_10132);
nor U10626 (N_10626,N_9824,N_9936);
nor U10627 (N_10627,N_10119,N_10107);
nand U10628 (N_10628,N_9895,N_9900);
nor U10629 (N_10629,N_9691,N_9850);
or U10630 (N_10630,N_9676,N_10142);
and U10631 (N_10631,N_9849,N_10060);
or U10632 (N_10632,N_10191,N_9901);
nand U10633 (N_10633,N_9717,N_9837);
and U10634 (N_10634,N_9940,N_9704);
xor U10635 (N_10635,N_9608,N_9931);
nand U10636 (N_10636,N_10025,N_9694);
or U10637 (N_10637,N_10098,N_9942);
and U10638 (N_10638,N_10182,N_9800);
nand U10639 (N_10639,N_9761,N_9669);
or U10640 (N_10640,N_9647,N_10089);
nor U10641 (N_10641,N_9632,N_10041);
nand U10642 (N_10642,N_9873,N_10095);
and U10643 (N_10643,N_10004,N_9765);
and U10644 (N_10644,N_9734,N_9874);
and U10645 (N_10645,N_9833,N_9664);
nand U10646 (N_10646,N_9828,N_10170);
nand U10647 (N_10647,N_9659,N_10037);
xor U10648 (N_10648,N_9691,N_10056);
and U10649 (N_10649,N_9861,N_10187);
nand U10650 (N_10650,N_9926,N_10015);
or U10651 (N_10651,N_9862,N_10139);
nor U10652 (N_10652,N_10051,N_9685);
nand U10653 (N_10653,N_9824,N_9809);
or U10654 (N_10654,N_10094,N_9766);
or U10655 (N_10655,N_10080,N_9927);
nand U10656 (N_10656,N_9622,N_9887);
nor U10657 (N_10657,N_9861,N_9719);
and U10658 (N_10658,N_9854,N_9736);
nor U10659 (N_10659,N_10130,N_9795);
or U10660 (N_10660,N_9625,N_10117);
nor U10661 (N_10661,N_9856,N_9824);
or U10662 (N_10662,N_9771,N_10107);
nor U10663 (N_10663,N_9610,N_9625);
or U10664 (N_10664,N_9949,N_10010);
nand U10665 (N_10665,N_9895,N_10053);
nand U10666 (N_10666,N_9832,N_9947);
nand U10667 (N_10667,N_10075,N_9877);
nand U10668 (N_10668,N_9898,N_10186);
nor U10669 (N_10669,N_9915,N_9993);
nand U10670 (N_10670,N_9607,N_10131);
nand U10671 (N_10671,N_10188,N_9923);
nand U10672 (N_10672,N_10034,N_9860);
or U10673 (N_10673,N_10178,N_9735);
and U10674 (N_10674,N_9995,N_9963);
and U10675 (N_10675,N_9664,N_9728);
and U10676 (N_10676,N_10185,N_9919);
nand U10677 (N_10677,N_9646,N_9885);
nor U10678 (N_10678,N_9667,N_9605);
or U10679 (N_10679,N_10165,N_9840);
nand U10680 (N_10680,N_9618,N_9820);
or U10681 (N_10681,N_10142,N_9670);
and U10682 (N_10682,N_9798,N_9605);
nand U10683 (N_10683,N_9699,N_9794);
and U10684 (N_10684,N_9709,N_9745);
nor U10685 (N_10685,N_9947,N_10005);
or U10686 (N_10686,N_9646,N_9914);
nor U10687 (N_10687,N_9738,N_10102);
and U10688 (N_10688,N_9998,N_9688);
nand U10689 (N_10689,N_9858,N_10183);
nor U10690 (N_10690,N_9863,N_9859);
or U10691 (N_10691,N_9965,N_9821);
nand U10692 (N_10692,N_9946,N_9604);
and U10693 (N_10693,N_9796,N_9681);
or U10694 (N_10694,N_10076,N_9823);
nand U10695 (N_10695,N_9771,N_9863);
nor U10696 (N_10696,N_9860,N_9855);
nand U10697 (N_10697,N_10026,N_10043);
nor U10698 (N_10698,N_9988,N_9914);
nand U10699 (N_10699,N_9606,N_9741);
nor U10700 (N_10700,N_10105,N_9821);
nand U10701 (N_10701,N_9750,N_9863);
xor U10702 (N_10702,N_10064,N_9748);
and U10703 (N_10703,N_9931,N_9718);
nor U10704 (N_10704,N_10162,N_10181);
nor U10705 (N_10705,N_9613,N_9966);
and U10706 (N_10706,N_10125,N_9828);
and U10707 (N_10707,N_10140,N_9912);
nand U10708 (N_10708,N_10116,N_9649);
nand U10709 (N_10709,N_10030,N_9761);
xnor U10710 (N_10710,N_9873,N_10076);
nand U10711 (N_10711,N_9641,N_9913);
and U10712 (N_10712,N_9754,N_9988);
or U10713 (N_10713,N_9675,N_9951);
nand U10714 (N_10714,N_10099,N_10089);
or U10715 (N_10715,N_9640,N_10031);
and U10716 (N_10716,N_9957,N_10067);
and U10717 (N_10717,N_9839,N_10041);
or U10718 (N_10718,N_10069,N_9832);
nor U10719 (N_10719,N_10040,N_9675);
nor U10720 (N_10720,N_9909,N_10189);
nor U10721 (N_10721,N_9910,N_10111);
or U10722 (N_10722,N_9695,N_10164);
and U10723 (N_10723,N_9917,N_10123);
nor U10724 (N_10724,N_9848,N_10038);
and U10725 (N_10725,N_9912,N_9792);
or U10726 (N_10726,N_9798,N_9833);
and U10727 (N_10727,N_9782,N_9820);
or U10728 (N_10728,N_10185,N_9643);
nor U10729 (N_10729,N_9734,N_10107);
nor U10730 (N_10730,N_9915,N_10134);
and U10731 (N_10731,N_9772,N_9922);
nor U10732 (N_10732,N_9659,N_9901);
nand U10733 (N_10733,N_10162,N_9981);
nor U10734 (N_10734,N_9853,N_9831);
or U10735 (N_10735,N_10054,N_9600);
nor U10736 (N_10736,N_9936,N_9665);
or U10737 (N_10737,N_10043,N_9681);
nor U10738 (N_10738,N_9740,N_9959);
and U10739 (N_10739,N_9777,N_9833);
nand U10740 (N_10740,N_9631,N_9714);
nand U10741 (N_10741,N_10035,N_9949);
and U10742 (N_10742,N_9960,N_9920);
or U10743 (N_10743,N_9891,N_9847);
and U10744 (N_10744,N_9661,N_9958);
or U10745 (N_10745,N_9834,N_9746);
nand U10746 (N_10746,N_9864,N_9848);
and U10747 (N_10747,N_9748,N_9678);
nor U10748 (N_10748,N_10066,N_10045);
or U10749 (N_10749,N_10155,N_9634);
nand U10750 (N_10750,N_10176,N_9707);
and U10751 (N_10751,N_10137,N_9786);
xnor U10752 (N_10752,N_10171,N_9765);
or U10753 (N_10753,N_9819,N_9860);
or U10754 (N_10754,N_9900,N_10136);
and U10755 (N_10755,N_9785,N_10048);
nand U10756 (N_10756,N_9949,N_10044);
nor U10757 (N_10757,N_9972,N_9660);
or U10758 (N_10758,N_10181,N_9672);
nand U10759 (N_10759,N_9802,N_10152);
nand U10760 (N_10760,N_9959,N_9956);
and U10761 (N_10761,N_10188,N_9742);
nor U10762 (N_10762,N_9928,N_9867);
nor U10763 (N_10763,N_9878,N_10115);
nand U10764 (N_10764,N_10195,N_9968);
nor U10765 (N_10765,N_9794,N_9811);
nand U10766 (N_10766,N_9837,N_9768);
or U10767 (N_10767,N_9902,N_9801);
nand U10768 (N_10768,N_10026,N_9627);
nor U10769 (N_10769,N_10088,N_9602);
nor U10770 (N_10770,N_9824,N_9844);
and U10771 (N_10771,N_9649,N_9609);
nor U10772 (N_10772,N_9738,N_9975);
nor U10773 (N_10773,N_10175,N_9881);
nand U10774 (N_10774,N_9911,N_9694);
nand U10775 (N_10775,N_9857,N_9993);
nand U10776 (N_10776,N_9816,N_10199);
or U10777 (N_10777,N_9661,N_10194);
nand U10778 (N_10778,N_9804,N_9625);
or U10779 (N_10779,N_9787,N_9932);
nor U10780 (N_10780,N_10147,N_9714);
nand U10781 (N_10781,N_10002,N_9643);
nand U10782 (N_10782,N_10149,N_10040);
and U10783 (N_10783,N_9671,N_9741);
and U10784 (N_10784,N_9949,N_9995);
nor U10785 (N_10785,N_10002,N_9759);
and U10786 (N_10786,N_9937,N_9722);
nor U10787 (N_10787,N_9632,N_9673);
and U10788 (N_10788,N_9635,N_9904);
nor U10789 (N_10789,N_10162,N_10013);
and U10790 (N_10790,N_10008,N_10106);
or U10791 (N_10791,N_9779,N_9734);
xnor U10792 (N_10792,N_9754,N_9871);
or U10793 (N_10793,N_10019,N_9717);
and U10794 (N_10794,N_9726,N_9639);
xnor U10795 (N_10795,N_10144,N_9950);
or U10796 (N_10796,N_9835,N_9744);
and U10797 (N_10797,N_9831,N_10062);
and U10798 (N_10798,N_10185,N_9782);
or U10799 (N_10799,N_10078,N_9698);
or U10800 (N_10800,N_10476,N_10218);
nor U10801 (N_10801,N_10511,N_10386);
nand U10802 (N_10802,N_10616,N_10687);
or U10803 (N_10803,N_10596,N_10337);
nor U10804 (N_10804,N_10368,N_10708);
and U10805 (N_10805,N_10507,N_10308);
nor U10806 (N_10806,N_10665,N_10243);
nand U10807 (N_10807,N_10460,N_10467);
nand U10808 (N_10808,N_10454,N_10603);
or U10809 (N_10809,N_10381,N_10340);
nor U10810 (N_10810,N_10545,N_10220);
nand U10811 (N_10811,N_10746,N_10719);
nand U10812 (N_10812,N_10402,N_10542);
nor U10813 (N_10813,N_10272,N_10658);
nand U10814 (N_10814,N_10258,N_10215);
nand U10815 (N_10815,N_10271,N_10724);
or U10816 (N_10816,N_10682,N_10484);
nand U10817 (N_10817,N_10748,N_10360);
nor U10818 (N_10818,N_10413,N_10366);
and U10819 (N_10819,N_10699,N_10221);
xnor U10820 (N_10820,N_10492,N_10720);
xnor U10821 (N_10821,N_10580,N_10500);
or U10822 (N_10822,N_10644,N_10672);
nand U10823 (N_10823,N_10751,N_10445);
nand U10824 (N_10824,N_10374,N_10483);
nor U10825 (N_10825,N_10513,N_10282);
nor U10826 (N_10826,N_10641,N_10474);
nor U10827 (N_10827,N_10571,N_10225);
xor U10828 (N_10828,N_10795,N_10392);
and U10829 (N_10829,N_10534,N_10287);
or U10830 (N_10830,N_10320,N_10279);
nand U10831 (N_10831,N_10640,N_10285);
or U10832 (N_10832,N_10462,N_10559);
nor U10833 (N_10833,N_10356,N_10688);
or U10834 (N_10834,N_10239,N_10276);
nand U10835 (N_10835,N_10273,N_10395);
nand U10836 (N_10836,N_10556,N_10615);
nor U10837 (N_10837,N_10459,N_10601);
or U10838 (N_10838,N_10762,N_10697);
nand U10839 (N_10839,N_10351,N_10681);
nor U10840 (N_10840,N_10431,N_10245);
or U10841 (N_10841,N_10295,N_10291);
nor U10842 (N_10842,N_10635,N_10563);
nand U10843 (N_10843,N_10633,N_10557);
or U10844 (N_10844,N_10479,N_10261);
nand U10845 (N_10845,N_10758,N_10314);
or U10846 (N_10846,N_10451,N_10400);
xor U10847 (N_10847,N_10369,N_10367);
and U10848 (N_10848,N_10560,N_10543);
nor U10849 (N_10849,N_10458,N_10211);
and U10850 (N_10850,N_10772,N_10626);
nand U10851 (N_10851,N_10683,N_10650);
or U10852 (N_10852,N_10265,N_10561);
nand U10853 (N_10853,N_10437,N_10606);
nand U10854 (N_10854,N_10444,N_10229);
nand U10855 (N_10855,N_10551,N_10673);
or U10856 (N_10856,N_10266,N_10409);
xnor U10857 (N_10857,N_10638,N_10309);
nor U10858 (N_10858,N_10284,N_10318);
nand U10859 (N_10859,N_10254,N_10564);
nand U10860 (N_10860,N_10648,N_10625);
and U10861 (N_10861,N_10410,N_10355);
or U10862 (N_10862,N_10396,N_10750);
nand U10863 (N_10863,N_10389,N_10705);
nor U10864 (N_10864,N_10345,N_10628);
or U10865 (N_10865,N_10630,N_10624);
nor U10866 (N_10866,N_10540,N_10482);
or U10867 (N_10867,N_10422,N_10424);
and U10868 (N_10868,N_10307,N_10468);
or U10869 (N_10869,N_10394,N_10686);
or U10870 (N_10870,N_10676,N_10506);
nand U10871 (N_10871,N_10782,N_10792);
nand U10872 (N_10872,N_10446,N_10608);
and U10873 (N_10873,N_10533,N_10740);
nand U10874 (N_10874,N_10497,N_10365);
nand U10875 (N_10875,N_10696,N_10607);
or U10876 (N_10876,N_10572,N_10778);
and U10877 (N_10877,N_10494,N_10766);
or U10878 (N_10878,N_10645,N_10411);
nor U10879 (N_10879,N_10700,N_10594);
and U10880 (N_10880,N_10210,N_10486);
nand U10881 (N_10881,N_10662,N_10515);
nor U10882 (N_10882,N_10588,N_10425);
and U10883 (N_10883,N_10636,N_10722);
or U10884 (N_10884,N_10439,N_10344);
or U10885 (N_10885,N_10597,N_10579);
nor U10886 (N_10886,N_10569,N_10589);
or U10887 (N_10887,N_10327,N_10298);
or U10888 (N_10888,N_10598,N_10471);
nor U10889 (N_10889,N_10539,N_10783);
or U10890 (N_10890,N_10319,N_10775);
and U10891 (N_10891,N_10725,N_10592);
and U10892 (N_10892,N_10610,N_10779);
nand U10893 (N_10893,N_10346,N_10690);
and U10894 (N_10894,N_10657,N_10448);
nand U10895 (N_10895,N_10651,N_10599);
nor U10896 (N_10896,N_10264,N_10618);
nor U10897 (N_10897,N_10335,N_10737);
and U10898 (N_10898,N_10738,N_10678);
nor U10899 (N_10899,N_10763,N_10671);
nand U10900 (N_10900,N_10288,N_10226);
nand U10901 (N_10901,N_10242,N_10401);
nor U10902 (N_10902,N_10558,N_10537);
and U10903 (N_10903,N_10404,N_10698);
nor U10904 (N_10904,N_10277,N_10747);
or U10905 (N_10905,N_10332,N_10313);
nand U10906 (N_10906,N_10510,N_10528);
and U10907 (N_10907,N_10336,N_10350);
nand U10908 (N_10908,N_10380,N_10532);
and U10909 (N_10909,N_10518,N_10214);
and U10910 (N_10910,N_10378,N_10470);
nor U10911 (N_10911,N_10509,N_10595);
and U10912 (N_10912,N_10207,N_10364);
or U10913 (N_10913,N_10328,N_10680);
or U10914 (N_10914,N_10647,N_10734);
and U10915 (N_10915,N_10246,N_10338);
or U10916 (N_10916,N_10666,N_10372);
nand U10917 (N_10917,N_10634,N_10478);
nor U10918 (N_10918,N_10674,N_10407);
nor U10919 (N_10919,N_10612,N_10727);
or U10920 (N_10920,N_10216,N_10521);
and U10921 (N_10921,N_10416,N_10485);
and U10922 (N_10922,N_10565,N_10426);
nand U10923 (N_10923,N_10622,N_10253);
or U10924 (N_10924,N_10489,N_10793);
or U10925 (N_10925,N_10735,N_10694);
or U10926 (N_10926,N_10586,N_10428);
or U10927 (N_10927,N_10627,N_10538);
nand U10928 (N_10928,N_10656,N_10268);
nor U10929 (N_10929,N_10541,N_10693);
nand U10930 (N_10930,N_10472,N_10605);
nor U10931 (N_10931,N_10398,N_10326);
or U10932 (N_10932,N_10387,N_10611);
and U10933 (N_10933,N_10247,N_10602);
nor U10934 (N_10934,N_10679,N_10434);
or U10935 (N_10935,N_10701,N_10591);
and U10936 (N_10936,N_10726,N_10299);
xor U10937 (N_10937,N_10609,N_10774);
nor U10938 (N_10938,N_10383,N_10201);
nand U10939 (N_10939,N_10742,N_10691);
and U10940 (N_10940,N_10453,N_10512);
nor U10941 (N_10941,N_10604,N_10508);
and U10942 (N_10942,N_10375,N_10784);
nand U10943 (N_10943,N_10590,N_10728);
nand U10944 (N_10944,N_10516,N_10517);
nor U10945 (N_10945,N_10732,N_10491);
and U10946 (N_10946,N_10405,N_10452);
and U10947 (N_10947,N_10575,N_10717);
nand U10948 (N_10948,N_10224,N_10659);
nand U10949 (N_10949,N_10412,N_10323);
nand U10950 (N_10950,N_10397,N_10248);
and U10951 (N_10951,N_10522,N_10423);
nor U10952 (N_10952,N_10768,N_10790);
nor U10953 (N_10953,N_10357,N_10230);
nor U10954 (N_10954,N_10756,N_10791);
nor U10955 (N_10955,N_10436,N_10244);
or U10956 (N_10956,N_10526,N_10388);
and U10957 (N_10957,N_10233,N_10736);
and U10958 (N_10958,N_10716,N_10406);
and U10959 (N_10959,N_10469,N_10234);
nand U10960 (N_10960,N_10544,N_10524);
nor U10961 (N_10961,N_10384,N_10536);
nor U10962 (N_10962,N_10495,N_10550);
or U10963 (N_10963,N_10290,N_10730);
and U10964 (N_10964,N_10504,N_10343);
nor U10965 (N_10965,N_10450,N_10235);
or U10966 (N_10966,N_10228,N_10786);
or U10967 (N_10967,N_10713,N_10749);
nor U10968 (N_10968,N_10733,N_10353);
or U10969 (N_10969,N_10664,N_10562);
nor U10970 (N_10970,N_10721,N_10442);
nor U10971 (N_10971,N_10718,N_10223);
and U10972 (N_10972,N_10408,N_10278);
and U10973 (N_10973,N_10546,N_10256);
nor U10974 (N_10974,N_10455,N_10649);
and U10975 (N_10975,N_10731,N_10752);
nor U10976 (N_10976,N_10523,N_10619);
nand U10977 (N_10977,N_10283,N_10461);
nand U10978 (N_10978,N_10535,N_10473);
nor U10979 (N_10979,N_10370,N_10643);
nand U10980 (N_10980,N_10449,N_10270);
and U10981 (N_10981,N_10709,N_10776);
and U10982 (N_10982,N_10297,N_10227);
or U10983 (N_10983,N_10613,N_10306);
xor U10984 (N_10984,N_10785,N_10501);
or U10985 (N_10985,N_10796,N_10217);
nand U10986 (N_10986,N_10654,N_10669);
or U10987 (N_10987,N_10255,N_10677);
nor U10988 (N_10988,N_10312,N_10743);
and U10989 (N_10989,N_10767,N_10761);
and U10990 (N_10990,N_10639,N_10294);
nor U10991 (N_10991,N_10584,N_10582);
nand U10992 (N_10992,N_10250,N_10794);
nand U10993 (N_10993,N_10359,N_10661);
nor U10994 (N_10994,N_10715,N_10222);
nor U10995 (N_10995,N_10757,N_10593);
nor U10996 (N_10996,N_10237,N_10310);
and U10997 (N_10997,N_10621,N_10780);
nor U10998 (N_10998,N_10303,N_10354);
nand U10999 (N_10999,N_10689,N_10321);
or U11000 (N_11000,N_10531,N_10702);
nand U11001 (N_11001,N_10548,N_10296);
and U11002 (N_11002,N_10267,N_10311);
nor U11003 (N_11003,N_10723,N_10600);
nor U11004 (N_11004,N_10712,N_10739);
nor U11005 (N_11005,N_10668,N_10798);
nand U11006 (N_11006,N_10570,N_10463);
or U11007 (N_11007,N_10660,N_10417);
or U11008 (N_11008,N_10252,N_10617);
nor U11009 (N_11009,N_10286,N_10349);
and U11010 (N_11010,N_10393,N_10549);
and U11011 (N_11011,N_10257,N_10263);
nor U11012 (N_11012,N_10753,N_10213);
nor U11013 (N_11013,N_10711,N_10322);
and U11014 (N_11014,N_10710,N_10652);
nor U11015 (N_11015,N_10585,N_10391);
nand U11016 (N_11016,N_10200,N_10525);
or U11017 (N_11017,N_10520,N_10637);
nor U11018 (N_11018,N_10204,N_10440);
and U11019 (N_11019,N_10415,N_10347);
nand U11020 (N_11020,N_10799,N_10704);
xnor U11021 (N_11021,N_10503,N_10456);
nand U11022 (N_11022,N_10573,N_10480);
or U11023 (N_11023,N_10475,N_10623);
and U11024 (N_11024,N_10249,N_10764);
nor U11025 (N_11025,N_10376,N_10773);
nand U11026 (N_11026,N_10685,N_10275);
nand U11027 (N_11027,N_10232,N_10759);
nor U11028 (N_11028,N_10577,N_10341);
nand U11029 (N_11029,N_10302,N_10646);
or U11030 (N_11030,N_10419,N_10289);
or U11031 (N_11031,N_10385,N_10281);
nand U11032 (N_11032,N_10744,N_10342);
nand U11033 (N_11033,N_10777,N_10663);
nand U11034 (N_11034,N_10769,N_10241);
nor U11035 (N_11035,N_10552,N_10377);
and U11036 (N_11036,N_10655,N_10527);
or U11037 (N_11037,N_10466,N_10505);
and U11038 (N_11038,N_10707,N_10714);
nor U11039 (N_11039,N_10420,N_10429);
and U11040 (N_11040,N_10205,N_10447);
or U11041 (N_11041,N_10797,N_10352);
nand U11042 (N_11042,N_10293,N_10692);
or U11043 (N_11043,N_10576,N_10706);
or U11044 (N_11044,N_10519,N_10464);
nor U11045 (N_11045,N_10403,N_10427);
nor U11046 (N_11046,N_10745,N_10581);
or U11047 (N_11047,N_10330,N_10379);
nor U11048 (N_11048,N_10236,N_10667);
or U11049 (N_11049,N_10240,N_10755);
or U11050 (N_11050,N_10741,N_10765);
and U11051 (N_11051,N_10788,N_10362);
nor U11052 (N_11052,N_10771,N_10206);
and U11053 (N_11053,N_10333,N_10568);
nor U11054 (N_11054,N_10684,N_10529);
nand U11055 (N_11055,N_10490,N_10457);
or U11056 (N_11056,N_10789,N_10578);
and U11057 (N_11057,N_10305,N_10530);
or U11058 (N_11058,N_10209,N_10399);
nor U11059 (N_11059,N_10695,N_10300);
nor U11060 (N_11060,N_10202,N_10670);
and U11061 (N_11061,N_10481,N_10259);
nand U11062 (N_11062,N_10583,N_10208);
xor U11063 (N_11063,N_10781,N_10260);
or U11064 (N_11064,N_10325,N_10348);
nor U11065 (N_11065,N_10334,N_10361);
nor U11066 (N_11066,N_10433,N_10498);
nand U11067 (N_11067,N_10574,N_10219);
or U11068 (N_11068,N_10631,N_10438);
or U11069 (N_11069,N_10382,N_10547);
and U11070 (N_11070,N_10787,N_10567);
xnor U11071 (N_11071,N_10304,N_10770);
and U11072 (N_11072,N_10754,N_10432);
nand U11073 (N_11073,N_10729,N_10414);
or U11074 (N_11074,N_10371,N_10632);
and U11075 (N_11075,N_10553,N_10212);
and U11076 (N_11076,N_10587,N_10443);
or U11077 (N_11077,N_10499,N_10238);
and U11078 (N_11078,N_10373,N_10315);
and U11079 (N_11079,N_10642,N_10487);
or U11080 (N_11080,N_10496,N_10502);
nand U11081 (N_11081,N_10620,N_10231);
nand U11082 (N_11082,N_10292,N_10477);
or U11083 (N_11083,N_10251,N_10358);
or U11084 (N_11084,N_10629,N_10760);
nor U11085 (N_11085,N_10435,N_10653);
xor U11086 (N_11086,N_10465,N_10316);
nand U11087 (N_11087,N_10421,N_10493);
or U11088 (N_11088,N_10566,N_10675);
nand U11089 (N_11089,N_10280,N_10514);
or U11090 (N_11090,N_10418,N_10317);
or U11091 (N_11091,N_10301,N_10488);
or U11092 (N_11092,N_10203,N_10329);
and U11093 (N_11093,N_10262,N_10269);
or U11094 (N_11094,N_10441,N_10703);
nor U11095 (N_11095,N_10339,N_10555);
nand U11096 (N_11096,N_10363,N_10324);
nand U11097 (N_11097,N_10554,N_10614);
nand U11098 (N_11098,N_10390,N_10430);
and U11099 (N_11099,N_10274,N_10331);
or U11100 (N_11100,N_10733,N_10394);
or U11101 (N_11101,N_10212,N_10559);
or U11102 (N_11102,N_10635,N_10799);
and U11103 (N_11103,N_10734,N_10589);
nand U11104 (N_11104,N_10695,N_10277);
or U11105 (N_11105,N_10319,N_10711);
nor U11106 (N_11106,N_10382,N_10286);
or U11107 (N_11107,N_10442,N_10619);
and U11108 (N_11108,N_10688,N_10374);
nand U11109 (N_11109,N_10655,N_10269);
and U11110 (N_11110,N_10474,N_10585);
and U11111 (N_11111,N_10288,N_10479);
xor U11112 (N_11112,N_10245,N_10793);
or U11113 (N_11113,N_10390,N_10407);
nand U11114 (N_11114,N_10298,N_10326);
and U11115 (N_11115,N_10514,N_10647);
nand U11116 (N_11116,N_10700,N_10521);
or U11117 (N_11117,N_10483,N_10246);
nand U11118 (N_11118,N_10227,N_10698);
nor U11119 (N_11119,N_10236,N_10471);
and U11120 (N_11120,N_10359,N_10768);
xor U11121 (N_11121,N_10734,N_10460);
and U11122 (N_11122,N_10533,N_10628);
and U11123 (N_11123,N_10412,N_10547);
nand U11124 (N_11124,N_10503,N_10218);
nor U11125 (N_11125,N_10421,N_10256);
or U11126 (N_11126,N_10541,N_10432);
nand U11127 (N_11127,N_10744,N_10556);
nand U11128 (N_11128,N_10294,N_10298);
nor U11129 (N_11129,N_10571,N_10372);
or U11130 (N_11130,N_10549,N_10749);
nor U11131 (N_11131,N_10676,N_10568);
nand U11132 (N_11132,N_10442,N_10547);
nand U11133 (N_11133,N_10658,N_10464);
and U11134 (N_11134,N_10685,N_10490);
nor U11135 (N_11135,N_10403,N_10484);
nand U11136 (N_11136,N_10358,N_10224);
nand U11137 (N_11137,N_10704,N_10371);
and U11138 (N_11138,N_10642,N_10285);
and U11139 (N_11139,N_10791,N_10603);
or U11140 (N_11140,N_10474,N_10722);
nor U11141 (N_11141,N_10543,N_10661);
and U11142 (N_11142,N_10255,N_10797);
nor U11143 (N_11143,N_10250,N_10505);
xor U11144 (N_11144,N_10272,N_10376);
or U11145 (N_11145,N_10644,N_10361);
or U11146 (N_11146,N_10590,N_10710);
nor U11147 (N_11147,N_10389,N_10396);
and U11148 (N_11148,N_10721,N_10354);
and U11149 (N_11149,N_10425,N_10797);
nand U11150 (N_11150,N_10229,N_10795);
or U11151 (N_11151,N_10286,N_10220);
and U11152 (N_11152,N_10362,N_10514);
nand U11153 (N_11153,N_10547,N_10647);
nor U11154 (N_11154,N_10592,N_10598);
xor U11155 (N_11155,N_10784,N_10264);
nor U11156 (N_11156,N_10585,N_10508);
nand U11157 (N_11157,N_10504,N_10237);
and U11158 (N_11158,N_10201,N_10596);
and U11159 (N_11159,N_10292,N_10693);
nand U11160 (N_11160,N_10336,N_10738);
nor U11161 (N_11161,N_10794,N_10358);
or U11162 (N_11162,N_10767,N_10609);
nand U11163 (N_11163,N_10303,N_10366);
or U11164 (N_11164,N_10429,N_10776);
nor U11165 (N_11165,N_10656,N_10399);
and U11166 (N_11166,N_10284,N_10613);
nor U11167 (N_11167,N_10603,N_10474);
or U11168 (N_11168,N_10582,N_10746);
nand U11169 (N_11169,N_10565,N_10746);
or U11170 (N_11170,N_10658,N_10728);
nand U11171 (N_11171,N_10354,N_10727);
xor U11172 (N_11172,N_10392,N_10334);
nor U11173 (N_11173,N_10769,N_10648);
nand U11174 (N_11174,N_10647,N_10544);
nand U11175 (N_11175,N_10296,N_10665);
or U11176 (N_11176,N_10648,N_10626);
nor U11177 (N_11177,N_10361,N_10729);
or U11178 (N_11178,N_10342,N_10427);
and U11179 (N_11179,N_10707,N_10748);
nor U11180 (N_11180,N_10707,N_10777);
nor U11181 (N_11181,N_10316,N_10602);
or U11182 (N_11182,N_10793,N_10548);
nand U11183 (N_11183,N_10458,N_10476);
and U11184 (N_11184,N_10518,N_10547);
or U11185 (N_11185,N_10276,N_10678);
or U11186 (N_11186,N_10235,N_10773);
nor U11187 (N_11187,N_10552,N_10626);
and U11188 (N_11188,N_10731,N_10701);
and U11189 (N_11189,N_10313,N_10477);
and U11190 (N_11190,N_10770,N_10327);
nand U11191 (N_11191,N_10621,N_10557);
and U11192 (N_11192,N_10471,N_10356);
or U11193 (N_11193,N_10404,N_10600);
and U11194 (N_11194,N_10695,N_10207);
nand U11195 (N_11195,N_10460,N_10644);
xnor U11196 (N_11196,N_10266,N_10262);
nor U11197 (N_11197,N_10565,N_10466);
or U11198 (N_11198,N_10332,N_10542);
nand U11199 (N_11199,N_10509,N_10599);
or U11200 (N_11200,N_10669,N_10347);
and U11201 (N_11201,N_10378,N_10474);
nor U11202 (N_11202,N_10752,N_10712);
or U11203 (N_11203,N_10369,N_10549);
and U11204 (N_11204,N_10302,N_10570);
and U11205 (N_11205,N_10219,N_10411);
nand U11206 (N_11206,N_10366,N_10255);
or U11207 (N_11207,N_10734,N_10604);
and U11208 (N_11208,N_10703,N_10300);
or U11209 (N_11209,N_10206,N_10442);
nand U11210 (N_11210,N_10254,N_10488);
nand U11211 (N_11211,N_10267,N_10484);
nand U11212 (N_11212,N_10699,N_10377);
and U11213 (N_11213,N_10372,N_10339);
or U11214 (N_11214,N_10210,N_10740);
nor U11215 (N_11215,N_10777,N_10286);
and U11216 (N_11216,N_10470,N_10696);
nor U11217 (N_11217,N_10220,N_10380);
or U11218 (N_11218,N_10419,N_10790);
and U11219 (N_11219,N_10685,N_10230);
xnor U11220 (N_11220,N_10648,N_10689);
xnor U11221 (N_11221,N_10427,N_10757);
and U11222 (N_11222,N_10227,N_10259);
nor U11223 (N_11223,N_10414,N_10633);
or U11224 (N_11224,N_10216,N_10784);
and U11225 (N_11225,N_10566,N_10266);
and U11226 (N_11226,N_10297,N_10543);
and U11227 (N_11227,N_10622,N_10589);
nand U11228 (N_11228,N_10625,N_10529);
or U11229 (N_11229,N_10326,N_10274);
nor U11230 (N_11230,N_10383,N_10487);
or U11231 (N_11231,N_10260,N_10434);
xor U11232 (N_11232,N_10506,N_10727);
nor U11233 (N_11233,N_10616,N_10317);
nor U11234 (N_11234,N_10328,N_10209);
and U11235 (N_11235,N_10652,N_10281);
nor U11236 (N_11236,N_10415,N_10281);
xnor U11237 (N_11237,N_10273,N_10525);
and U11238 (N_11238,N_10465,N_10449);
nor U11239 (N_11239,N_10429,N_10565);
nand U11240 (N_11240,N_10645,N_10703);
nor U11241 (N_11241,N_10398,N_10257);
nor U11242 (N_11242,N_10263,N_10245);
or U11243 (N_11243,N_10643,N_10369);
nor U11244 (N_11244,N_10733,N_10761);
and U11245 (N_11245,N_10606,N_10367);
and U11246 (N_11246,N_10515,N_10359);
nor U11247 (N_11247,N_10540,N_10650);
xor U11248 (N_11248,N_10446,N_10401);
nor U11249 (N_11249,N_10721,N_10524);
nor U11250 (N_11250,N_10331,N_10728);
nor U11251 (N_11251,N_10673,N_10304);
nand U11252 (N_11252,N_10592,N_10574);
xor U11253 (N_11253,N_10264,N_10649);
or U11254 (N_11254,N_10347,N_10482);
nor U11255 (N_11255,N_10639,N_10595);
and U11256 (N_11256,N_10474,N_10726);
nand U11257 (N_11257,N_10441,N_10641);
or U11258 (N_11258,N_10713,N_10785);
and U11259 (N_11259,N_10786,N_10579);
nand U11260 (N_11260,N_10451,N_10418);
or U11261 (N_11261,N_10287,N_10377);
xor U11262 (N_11262,N_10377,N_10533);
nand U11263 (N_11263,N_10368,N_10296);
or U11264 (N_11264,N_10784,N_10568);
or U11265 (N_11265,N_10589,N_10400);
nand U11266 (N_11266,N_10355,N_10613);
or U11267 (N_11267,N_10380,N_10293);
nor U11268 (N_11268,N_10699,N_10355);
and U11269 (N_11269,N_10467,N_10419);
or U11270 (N_11270,N_10300,N_10432);
nand U11271 (N_11271,N_10225,N_10723);
nand U11272 (N_11272,N_10509,N_10206);
or U11273 (N_11273,N_10334,N_10790);
or U11274 (N_11274,N_10713,N_10361);
and U11275 (N_11275,N_10254,N_10377);
nand U11276 (N_11276,N_10286,N_10576);
nand U11277 (N_11277,N_10642,N_10486);
nand U11278 (N_11278,N_10209,N_10690);
and U11279 (N_11279,N_10778,N_10347);
nand U11280 (N_11280,N_10727,N_10204);
nor U11281 (N_11281,N_10261,N_10544);
or U11282 (N_11282,N_10438,N_10567);
nor U11283 (N_11283,N_10514,N_10614);
nor U11284 (N_11284,N_10639,N_10603);
and U11285 (N_11285,N_10411,N_10598);
or U11286 (N_11286,N_10228,N_10429);
and U11287 (N_11287,N_10758,N_10777);
nand U11288 (N_11288,N_10590,N_10297);
and U11289 (N_11289,N_10797,N_10788);
nand U11290 (N_11290,N_10679,N_10581);
or U11291 (N_11291,N_10792,N_10595);
nand U11292 (N_11292,N_10370,N_10542);
and U11293 (N_11293,N_10479,N_10406);
or U11294 (N_11294,N_10754,N_10524);
nand U11295 (N_11295,N_10227,N_10707);
nor U11296 (N_11296,N_10237,N_10724);
or U11297 (N_11297,N_10796,N_10256);
or U11298 (N_11298,N_10429,N_10559);
nor U11299 (N_11299,N_10665,N_10249);
nor U11300 (N_11300,N_10205,N_10237);
or U11301 (N_11301,N_10276,N_10581);
and U11302 (N_11302,N_10658,N_10295);
or U11303 (N_11303,N_10216,N_10556);
nor U11304 (N_11304,N_10797,N_10315);
and U11305 (N_11305,N_10415,N_10241);
or U11306 (N_11306,N_10473,N_10784);
nor U11307 (N_11307,N_10238,N_10789);
and U11308 (N_11308,N_10401,N_10350);
or U11309 (N_11309,N_10275,N_10756);
or U11310 (N_11310,N_10357,N_10695);
or U11311 (N_11311,N_10335,N_10254);
nor U11312 (N_11312,N_10732,N_10225);
and U11313 (N_11313,N_10275,N_10693);
nor U11314 (N_11314,N_10261,N_10702);
or U11315 (N_11315,N_10577,N_10644);
and U11316 (N_11316,N_10446,N_10257);
and U11317 (N_11317,N_10517,N_10419);
nor U11318 (N_11318,N_10758,N_10714);
or U11319 (N_11319,N_10289,N_10602);
nor U11320 (N_11320,N_10211,N_10303);
nor U11321 (N_11321,N_10630,N_10393);
and U11322 (N_11322,N_10274,N_10350);
nor U11323 (N_11323,N_10496,N_10552);
and U11324 (N_11324,N_10430,N_10492);
nor U11325 (N_11325,N_10506,N_10710);
and U11326 (N_11326,N_10599,N_10433);
or U11327 (N_11327,N_10606,N_10741);
or U11328 (N_11328,N_10748,N_10733);
nand U11329 (N_11329,N_10505,N_10237);
and U11330 (N_11330,N_10289,N_10339);
nor U11331 (N_11331,N_10744,N_10369);
or U11332 (N_11332,N_10386,N_10294);
and U11333 (N_11333,N_10731,N_10541);
nand U11334 (N_11334,N_10728,N_10274);
nand U11335 (N_11335,N_10442,N_10623);
nor U11336 (N_11336,N_10658,N_10480);
or U11337 (N_11337,N_10725,N_10243);
nand U11338 (N_11338,N_10483,N_10285);
nor U11339 (N_11339,N_10737,N_10602);
nand U11340 (N_11340,N_10409,N_10439);
and U11341 (N_11341,N_10579,N_10413);
nor U11342 (N_11342,N_10479,N_10334);
nor U11343 (N_11343,N_10623,N_10765);
or U11344 (N_11344,N_10490,N_10201);
nand U11345 (N_11345,N_10403,N_10276);
and U11346 (N_11346,N_10215,N_10360);
nand U11347 (N_11347,N_10757,N_10774);
and U11348 (N_11348,N_10342,N_10370);
or U11349 (N_11349,N_10340,N_10509);
and U11350 (N_11350,N_10741,N_10551);
nor U11351 (N_11351,N_10525,N_10403);
nor U11352 (N_11352,N_10568,N_10219);
nand U11353 (N_11353,N_10295,N_10215);
nand U11354 (N_11354,N_10433,N_10549);
nor U11355 (N_11355,N_10490,N_10439);
or U11356 (N_11356,N_10206,N_10352);
xor U11357 (N_11357,N_10739,N_10537);
and U11358 (N_11358,N_10272,N_10221);
and U11359 (N_11359,N_10344,N_10641);
or U11360 (N_11360,N_10244,N_10218);
and U11361 (N_11361,N_10379,N_10548);
and U11362 (N_11362,N_10366,N_10322);
and U11363 (N_11363,N_10624,N_10797);
nor U11364 (N_11364,N_10701,N_10655);
and U11365 (N_11365,N_10700,N_10321);
nor U11366 (N_11366,N_10397,N_10359);
nand U11367 (N_11367,N_10262,N_10470);
nor U11368 (N_11368,N_10508,N_10490);
or U11369 (N_11369,N_10200,N_10746);
nor U11370 (N_11370,N_10543,N_10730);
or U11371 (N_11371,N_10253,N_10230);
nand U11372 (N_11372,N_10278,N_10282);
nand U11373 (N_11373,N_10362,N_10738);
nand U11374 (N_11374,N_10722,N_10356);
nand U11375 (N_11375,N_10292,N_10236);
nor U11376 (N_11376,N_10260,N_10530);
and U11377 (N_11377,N_10427,N_10482);
or U11378 (N_11378,N_10456,N_10669);
and U11379 (N_11379,N_10298,N_10286);
xor U11380 (N_11380,N_10367,N_10252);
xnor U11381 (N_11381,N_10632,N_10437);
nand U11382 (N_11382,N_10715,N_10276);
and U11383 (N_11383,N_10403,N_10796);
nand U11384 (N_11384,N_10464,N_10278);
and U11385 (N_11385,N_10362,N_10525);
nor U11386 (N_11386,N_10724,N_10571);
nor U11387 (N_11387,N_10202,N_10724);
or U11388 (N_11388,N_10537,N_10775);
and U11389 (N_11389,N_10615,N_10561);
and U11390 (N_11390,N_10309,N_10252);
and U11391 (N_11391,N_10542,N_10484);
nand U11392 (N_11392,N_10305,N_10593);
xor U11393 (N_11393,N_10753,N_10396);
and U11394 (N_11394,N_10298,N_10770);
or U11395 (N_11395,N_10217,N_10752);
nor U11396 (N_11396,N_10323,N_10558);
or U11397 (N_11397,N_10545,N_10706);
nand U11398 (N_11398,N_10629,N_10361);
and U11399 (N_11399,N_10364,N_10710);
and U11400 (N_11400,N_11354,N_10833);
and U11401 (N_11401,N_11245,N_11134);
nand U11402 (N_11402,N_11202,N_10829);
nand U11403 (N_11403,N_10894,N_10975);
or U11404 (N_11404,N_11284,N_10839);
nand U11405 (N_11405,N_11240,N_11103);
nor U11406 (N_11406,N_10990,N_11126);
nand U11407 (N_11407,N_10875,N_11144);
and U11408 (N_11408,N_11345,N_11229);
and U11409 (N_11409,N_10972,N_11180);
nor U11410 (N_11410,N_10982,N_11380);
xnor U11411 (N_11411,N_10929,N_10911);
and U11412 (N_11412,N_10905,N_11005);
nand U11413 (N_11413,N_11095,N_11153);
or U11414 (N_11414,N_10866,N_11259);
or U11415 (N_11415,N_10967,N_11042);
or U11416 (N_11416,N_11270,N_10968);
xor U11417 (N_11417,N_10938,N_11088);
nand U11418 (N_11418,N_11030,N_10945);
and U11419 (N_11419,N_10874,N_10822);
nor U11420 (N_11420,N_11300,N_10999);
nand U11421 (N_11421,N_11043,N_11185);
or U11422 (N_11422,N_11223,N_10898);
nor U11423 (N_11423,N_11399,N_10966);
nor U11424 (N_11424,N_11241,N_11159);
nor U11425 (N_11425,N_11031,N_10997);
and U11426 (N_11426,N_10949,N_10925);
nor U11427 (N_11427,N_10873,N_10980);
nand U11428 (N_11428,N_11371,N_11288);
and U11429 (N_11429,N_11023,N_11108);
nand U11430 (N_11430,N_11091,N_11228);
and U11431 (N_11431,N_10983,N_11182);
and U11432 (N_11432,N_11295,N_11324);
nor U11433 (N_11433,N_11029,N_10915);
or U11434 (N_11434,N_11203,N_11028);
or U11435 (N_11435,N_11049,N_11332);
or U11436 (N_11436,N_10892,N_10852);
nor U11437 (N_11437,N_11056,N_10821);
and U11438 (N_11438,N_10813,N_11236);
or U11439 (N_11439,N_11131,N_11150);
nand U11440 (N_11440,N_10961,N_10823);
nand U11441 (N_11441,N_10812,N_11363);
nor U11442 (N_11442,N_11343,N_11075);
or U11443 (N_11443,N_11276,N_11096);
nor U11444 (N_11444,N_10817,N_10974);
nand U11445 (N_11445,N_11356,N_10831);
nor U11446 (N_11446,N_10806,N_11162);
and U11447 (N_11447,N_11334,N_11122);
and U11448 (N_11448,N_11289,N_11148);
nand U11449 (N_11449,N_11283,N_10828);
or U11450 (N_11450,N_11348,N_11322);
or U11451 (N_11451,N_11204,N_11372);
and U11452 (N_11452,N_11243,N_11205);
and U11453 (N_11453,N_10919,N_10973);
nor U11454 (N_11454,N_10801,N_11156);
and U11455 (N_11455,N_10927,N_11124);
or U11456 (N_11456,N_10991,N_11287);
and U11457 (N_11457,N_11141,N_11151);
and U11458 (N_11458,N_11004,N_10969);
nor U11459 (N_11459,N_11021,N_11214);
or U11460 (N_11460,N_10985,N_11158);
nand U11461 (N_11461,N_10855,N_11076);
nand U11462 (N_11462,N_11398,N_11253);
nand U11463 (N_11463,N_11367,N_11377);
and U11464 (N_11464,N_11269,N_11045);
and U11465 (N_11465,N_11020,N_11169);
and U11466 (N_11466,N_11211,N_11093);
nor U11467 (N_11467,N_11335,N_11083);
nand U11468 (N_11468,N_10917,N_10808);
nor U11469 (N_11469,N_11032,N_11138);
nand U11470 (N_11470,N_10820,N_10950);
xor U11471 (N_11471,N_10844,N_11188);
nand U11472 (N_11472,N_11050,N_11320);
nand U11473 (N_11473,N_11170,N_11206);
and U11474 (N_11474,N_11209,N_11198);
or U11475 (N_11475,N_10928,N_11107);
and U11476 (N_11476,N_10888,N_11225);
or U11477 (N_11477,N_11316,N_11341);
nand U11478 (N_11478,N_11186,N_11000);
nor U11479 (N_11479,N_11364,N_11114);
nand U11480 (N_11480,N_11081,N_11177);
nor U11481 (N_11481,N_10960,N_11145);
nand U11482 (N_11482,N_11067,N_10872);
nand U11483 (N_11483,N_11393,N_10804);
and U11484 (N_11484,N_11244,N_10887);
nand U11485 (N_11485,N_11314,N_11392);
and U11486 (N_11486,N_11331,N_11387);
or U11487 (N_11487,N_11167,N_11007);
or U11488 (N_11488,N_11113,N_11351);
nor U11489 (N_11489,N_11140,N_10996);
or U11490 (N_11490,N_11116,N_11220);
nand U11491 (N_11491,N_11040,N_10937);
nand U11492 (N_11492,N_10900,N_10935);
nand U11493 (N_11493,N_11217,N_11163);
or U11494 (N_11494,N_10908,N_10859);
nand U11495 (N_11495,N_11369,N_11313);
or U11496 (N_11496,N_10881,N_11135);
nor U11497 (N_11497,N_11157,N_11099);
nand U11498 (N_11498,N_10933,N_11390);
nor U11499 (N_11499,N_10847,N_11038);
nand U11500 (N_11500,N_11060,N_10877);
and U11501 (N_11501,N_10932,N_11058);
nand U11502 (N_11502,N_10802,N_11246);
nor U11503 (N_11503,N_10891,N_11179);
nand U11504 (N_11504,N_10998,N_11395);
nand U11505 (N_11505,N_11053,N_10864);
nand U11506 (N_11506,N_11342,N_11044);
or U11507 (N_11507,N_11216,N_10834);
or U11508 (N_11508,N_10811,N_11027);
nor U11509 (N_11509,N_10986,N_11193);
or U11510 (N_11510,N_11172,N_11082);
or U11511 (N_11511,N_11263,N_10816);
and U11512 (N_11512,N_11018,N_11368);
and U11513 (N_11513,N_10842,N_10846);
nand U11514 (N_11514,N_11176,N_10850);
nor U11515 (N_11515,N_10912,N_11366);
nand U11516 (N_11516,N_11391,N_10907);
nor U11517 (N_11517,N_10944,N_11078);
nand U11518 (N_11518,N_11226,N_11340);
nor U11519 (N_11519,N_11274,N_11128);
and U11520 (N_11520,N_11199,N_10899);
nor U11521 (N_11521,N_11352,N_11155);
or U11522 (N_11522,N_11278,N_11092);
and U11523 (N_11523,N_10869,N_11090);
nor U11524 (N_11524,N_10976,N_11349);
nor U11525 (N_11525,N_11271,N_11101);
nor U11526 (N_11526,N_11006,N_11074);
nor U11527 (N_11527,N_11080,N_11257);
nor U11528 (N_11528,N_10931,N_11299);
and U11529 (N_11529,N_11189,N_10941);
nor U11530 (N_11530,N_11059,N_11164);
and U11531 (N_11531,N_11196,N_11282);
nor U11532 (N_11532,N_10978,N_10838);
nor U11533 (N_11533,N_11111,N_11133);
nand U11534 (N_11534,N_11321,N_10836);
nand U11535 (N_11535,N_11258,N_11033);
nor U11536 (N_11536,N_11230,N_11051);
or U11537 (N_11537,N_10994,N_10964);
and U11538 (N_11538,N_11037,N_11394);
nand U11539 (N_11539,N_11277,N_11089);
or U11540 (N_11540,N_10923,N_11290);
nand U11541 (N_11541,N_11120,N_11197);
nand U11542 (N_11542,N_11190,N_11001);
nand U11543 (N_11543,N_11238,N_10971);
nor U11544 (N_11544,N_11171,N_11070);
and U11545 (N_11545,N_11362,N_11308);
and U11546 (N_11546,N_10979,N_10862);
and U11547 (N_11547,N_11275,N_11222);
or U11548 (N_11548,N_11085,N_11146);
nor U11549 (N_11549,N_11184,N_11213);
or U11550 (N_11550,N_11112,N_11130);
nor U11551 (N_11551,N_10880,N_10840);
nand U11552 (N_11552,N_11389,N_10921);
nor U11553 (N_11553,N_11381,N_11118);
and U11554 (N_11554,N_10948,N_11194);
nor U11555 (N_11555,N_11237,N_11383);
xor U11556 (N_11556,N_10884,N_10930);
nor U11557 (N_11557,N_11315,N_11046);
or U11558 (N_11558,N_10824,N_10963);
and U11559 (N_11559,N_10860,N_11055);
nor U11560 (N_11560,N_11212,N_10814);
or U11561 (N_11561,N_11154,N_11323);
nand U11562 (N_11562,N_11142,N_11117);
nand U11563 (N_11563,N_11181,N_10910);
xnor U11564 (N_11564,N_11248,N_11012);
and U11565 (N_11565,N_10882,N_11079);
nor U11566 (N_11566,N_10987,N_10807);
or U11567 (N_11567,N_10835,N_11261);
and U11568 (N_11568,N_11165,N_10954);
or U11569 (N_11569,N_11219,N_10863);
or U11570 (N_11570,N_10870,N_11234);
or U11571 (N_11571,N_10819,N_11125);
nor U11572 (N_11572,N_11298,N_10904);
or U11573 (N_11573,N_11357,N_10832);
or U11574 (N_11574,N_11011,N_10946);
or U11575 (N_11575,N_11337,N_11339);
and U11576 (N_11576,N_11132,N_10988);
nand U11577 (N_11577,N_11336,N_11260);
and U11578 (N_11578,N_11087,N_11265);
nand U11579 (N_11579,N_11396,N_11303);
and U11580 (N_11580,N_10893,N_11115);
nand U11581 (N_11581,N_11218,N_11014);
nor U11582 (N_11582,N_10913,N_11242);
nand U11583 (N_11583,N_11178,N_11015);
nand U11584 (N_11584,N_11311,N_10815);
and U11585 (N_11585,N_11294,N_10858);
or U11586 (N_11586,N_11328,N_11346);
nor U11587 (N_11587,N_11267,N_10841);
and U11588 (N_11588,N_11231,N_11256);
nor U11589 (N_11589,N_11071,N_11305);
nand U11590 (N_11590,N_10879,N_11086);
nor U11591 (N_11591,N_11227,N_10897);
nand U11592 (N_11592,N_11192,N_11036);
nand U11593 (N_11593,N_10843,N_11350);
and U11594 (N_11594,N_11378,N_11106);
nor U11595 (N_11595,N_10918,N_11183);
or U11596 (N_11596,N_11065,N_11054);
nand U11597 (N_11597,N_11013,N_11268);
xnor U11598 (N_11598,N_11123,N_11008);
nor U11599 (N_11599,N_10818,N_10854);
nor U11600 (N_11600,N_11002,N_11062);
or U11601 (N_11601,N_11039,N_11297);
and U11602 (N_11602,N_10995,N_11069);
nand U11603 (N_11603,N_11143,N_10886);
or U11604 (N_11604,N_10993,N_11152);
nor U11605 (N_11605,N_10920,N_11077);
or U11606 (N_11606,N_11104,N_11309);
xor U11607 (N_11607,N_10902,N_11384);
or U11608 (N_11608,N_10827,N_11251);
xnor U11609 (N_11609,N_10957,N_11136);
and U11610 (N_11610,N_11224,N_11310);
nor U11611 (N_11611,N_10953,N_11022);
nand U11612 (N_11612,N_11373,N_10914);
and U11613 (N_11613,N_11047,N_11382);
and U11614 (N_11614,N_11376,N_11191);
nand U11615 (N_11615,N_11221,N_11375);
or U11616 (N_11616,N_11010,N_11250);
nand U11617 (N_11617,N_11306,N_11360);
nand U11618 (N_11618,N_11266,N_10895);
and U11619 (N_11619,N_10903,N_11379);
or U11620 (N_11620,N_11129,N_11317);
nor U11621 (N_11621,N_11397,N_11304);
and U11622 (N_11622,N_11064,N_11312);
nand U11623 (N_11623,N_10965,N_11239);
nor U11624 (N_11624,N_11235,N_11307);
or U11625 (N_11625,N_11100,N_10889);
nor U11626 (N_11626,N_10956,N_11329);
and U11627 (N_11627,N_10826,N_11232);
and U11628 (N_11628,N_10992,N_11016);
or U11629 (N_11629,N_10837,N_11024);
nor U11630 (N_11630,N_11147,N_11249);
nor U11631 (N_11631,N_11127,N_11355);
nor U11632 (N_11632,N_11279,N_11291);
xnor U11633 (N_11633,N_11388,N_11121);
and U11634 (N_11634,N_11026,N_10853);
and U11635 (N_11635,N_11052,N_10943);
and U11636 (N_11636,N_10952,N_11370);
nand U11637 (N_11637,N_11347,N_11201);
and U11638 (N_11638,N_10940,N_11161);
and U11639 (N_11639,N_10800,N_11338);
or U11640 (N_11640,N_11264,N_11286);
and U11641 (N_11641,N_11326,N_10958);
nand U11642 (N_11642,N_11385,N_11207);
nor U11643 (N_11643,N_10924,N_11149);
nand U11644 (N_11644,N_11292,N_10939);
and U11645 (N_11645,N_11333,N_11374);
nor U11646 (N_11646,N_11017,N_11068);
and U11647 (N_11647,N_11272,N_11365);
nor U11648 (N_11648,N_11262,N_11208);
and U11649 (N_11649,N_11063,N_11254);
nand U11650 (N_11650,N_10984,N_10885);
nor U11651 (N_11651,N_10810,N_10845);
or U11652 (N_11652,N_11233,N_11358);
or U11653 (N_11653,N_11296,N_11102);
nand U11654 (N_11654,N_11035,N_10868);
nand U11655 (N_11655,N_10890,N_11034);
nand U11656 (N_11656,N_10867,N_10951);
nand U11657 (N_11657,N_11025,N_11325);
nand U11658 (N_11658,N_11084,N_11187);
or U11659 (N_11659,N_11273,N_11252);
or U11660 (N_11660,N_11057,N_10803);
nand U11661 (N_11661,N_11160,N_10906);
nand U11662 (N_11662,N_11166,N_11066);
nor U11663 (N_11663,N_11330,N_11098);
xnor U11664 (N_11664,N_11174,N_11318);
nor U11665 (N_11665,N_11139,N_11173);
nor U11666 (N_11666,N_10977,N_11200);
and U11667 (N_11667,N_11301,N_11302);
or U11668 (N_11668,N_10849,N_10878);
and U11669 (N_11669,N_11061,N_10865);
and U11670 (N_11670,N_10959,N_10962);
nand U11671 (N_11671,N_10947,N_11019);
nand U11672 (N_11672,N_11009,N_11210);
nor U11673 (N_11673,N_10989,N_10876);
or U11674 (N_11674,N_10916,N_11359);
nand U11675 (N_11675,N_11048,N_10830);
nor U11676 (N_11676,N_11119,N_10805);
nand U11677 (N_11677,N_10909,N_10934);
and U11678 (N_11678,N_11072,N_11280);
nand U11679 (N_11679,N_10981,N_11285);
or U11680 (N_11680,N_10861,N_11247);
or U11681 (N_11681,N_11094,N_11255);
and U11682 (N_11682,N_11105,N_10848);
and U11683 (N_11683,N_10896,N_11195);
and U11684 (N_11684,N_10857,N_10926);
nand U11685 (N_11685,N_11293,N_11168);
or U11686 (N_11686,N_11319,N_11361);
and U11687 (N_11687,N_11109,N_11175);
nor U11688 (N_11688,N_11215,N_11041);
nor U11689 (N_11689,N_11327,N_11344);
or U11690 (N_11690,N_11110,N_11137);
or U11691 (N_11691,N_11386,N_11073);
nor U11692 (N_11692,N_11353,N_10936);
nand U11693 (N_11693,N_10851,N_11281);
nand U11694 (N_11694,N_10922,N_10901);
and U11695 (N_11695,N_10809,N_10955);
nor U11696 (N_11696,N_10871,N_10883);
or U11697 (N_11697,N_10942,N_11097);
or U11698 (N_11698,N_10825,N_10970);
nor U11699 (N_11699,N_10856,N_11003);
nor U11700 (N_11700,N_10920,N_11046);
nor U11701 (N_11701,N_11169,N_10944);
nand U11702 (N_11702,N_10848,N_11049);
nand U11703 (N_11703,N_11069,N_10856);
and U11704 (N_11704,N_10942,N_10913);
or U11705 (N_11705,N_10942,N_11001);
or U11706 (N_11706,N_11054,N_11205);
or U11707 (N_11707,N_11129,N_10844);
and U11708 (N_11708,N_11081,N_11247);
nand U11709 (N_11709,N_10889,N_11011);
nand U11710 (N_11710,N_10881,N_11001);
nand U11711 (N_11711,N_11303,N_11114);
and U11712 (N_11712,N_11290,N_11161);
xnor U11713 (N_11713,N_11277,N_11138);
or U11714 (N_11714,N_11357,N_11356);
nor U11715 (N_11715,N_11283,N_11271);
nor U11716 (N_11716,N_11029,N_10980);
and U11717 (N_11717,N_11226,N_11310);
or U11718 (N_11718,N_10882,N_11245);
or U11719 (N_11719,N_10983,N_11277);
and U11720 (N_11720,N_10932,N_10806);
nor U11721 (N_11721,N_11318,N_10928);
nand U11722 (N_11722,N_11080,N_11370);
or U11723 (N_11723,N_11240,N_11167);
or U11724 (N_11724,N_11035,N_11278);
and U11725 (N_11725,N_11109,N_10825);
nor U11726 (N_11726,N_10962,N_11222);
and U11727 (N_11727,N_11119,N_11239);
or U11728 (N_11728,N_10945,N_10970);
nor U11729 (N_11729,N_10810,N_11361);
or U11730 (N_11730,N_11358,N_11066);
nor U11731 (N_11731,N_10995,N_11080);
and U11732 (N_11732,N_11245,N_10876);
or U11733 (N_11733,N_10830,N_11079);
xor U11734 (N_11734,N_11160,N_10908);
nand U11735 (N_11735,N_11251,N_11037);
nand U11736 (N_11736,N_11258,N_11206);
or U11737 (N_11737,N_10887,N_11189);
nand U11738 (N_11738,N_10930,N_10963);
or U11739 (N_11739,N_11109,N_10918);
or U11740 (N_11740,N_11393,N_11092);
or U11741 (N_11741,N_10930,N_11179);
or U11742 (N_11742,N_10827,N_10822);
nand U11743 (N_11743,N_10859,N_11056);
nor U11744 (N_11744,N_10813,N_11136);
nand U11745 (N_11745,N_11387,N_11210);
and U11746 (N_11746,N_10813,N_11199);
nand U11747 (N_11747,N_11172,N_11235);
or U11748 (N_11748,N_11002,N_10896);
and U11749 (N_11749,N_11300,N_11029);
and U11750 (N_11750,N_10923,N_10970);
nor U11751 (N_11751,N_11031,N_10882);
nor U11752 (N_11752,N_10860,N_11215);
or U11753 (N_11753,N_10898,N_11225);
nor U11754 (N_11754,N_11174,N_10899);
or U11755 (N_11755,N_11090,N_11276);
and U11756 (N_11756,N_11232,N_11181);
or U11757 (N_11757,N_11000,N_11146);
nor U11758 (N_11758,N_11393,N_10971);
nand U11759 (N_11759,N_11049,N_10876);
and U11760 (N_11760,N_10953,N_10930);
or U11761 (N_11761,N_11053,N_10897);
nor U11762 (N_11762,N_11211,N_10970);
nand U11763 (N_11763,N_11313,N_11219);
and U11764 (N_11764,N_10870,N_11392);
and U11765 (N_11765,N_11359,N_10831);
and U11766 (N_11766,N_11311,N_10871);
and U11767 (N_11767,N_10950,N_11199);
nand U11768 (N_11768,N_11161,N_11251);
nor U11769 (N_11769,N_11267,N_11297);
and U11770 (N_11770,N_11108,N_11067);
and U11771 (N_11771,N_11033,N_11330);
nand U11772 (N_11772,N_11211,N_11090);
or U11773 (N_11773,N_11013,N_10963);
nand U11774 (N_11774,N_11093,N_11087);
nor U11775 (N_11775,N_11169,N_11192);
and U11776 (N_11776,N_11159,N_11380);
xor U11777 (N_11777,N_11125,N_10904);
or U11778 (N_11778,N_10800,N_11336);
and U11779 (N_11779,N_11270,N_11008);
nor U11780 (N_11780,N_10886,N_10883);
or U11781 (N_11781,N_10994,N_11100);
nand U11782 (N_11782,N_10873,N_11288);
nand U11783 (N_11783,N_11031,N_10800);
nand U11784 (N_11784,N_10977,N_11299);
nor U11785 (N_11785,N_11327,N_10902);
nand U11786 (N_11786,N_11112,N_11350);
and U11787 (N_11787,N_10948,N_10962);
xnor U11788 (N_11788,N_11307,N_11372);
nand U11789 (N_11789,N_11128,N_11110);
or U11790 (N_11790,N_11228,N_10908);
nor U11791 (N_11791,N_11337,N_10907);
and U11792 (N_11792,N_10809,N_10823);
nor U11793 (N_11793,N_11147,N_11290);
nor U11794 (N_11794,N_10959,N_10872);
and U11795 (N_11795,N_11088,N_11270);
and U11796 (N_11796,N_11178,N_10961);
or U11797 (N_11797,N_11075,N_11326);
nor U11798 (N_11798,N_11097,N_10977);
nor U11799 (N_11799,N_10907,N_11195);
nand U11800 (N_11800,N_10983,N_10945);
and U11801 (N_11801,N_10959,N_10995);
and U11802 (N_11802,N_11309,N_11138);
nand U11803 (N_11803,N_11355,N_11384);
nor U11804 (N_11804,N_10848,N_11215);
nand U11805 (N_11805,N_10807,N_11043);
or U11806 (N_11806,N_10851,N_11341);
nor U11807 (N_11807,N_11016,N_11334);
nor U11808 (N_11808,N_11011,N_11057);
nor U11809 (N_11809,N_11103,N_10834);
or U11810 (N_11810,N_10825,N_11275);
or U11811 (N_11811,N_11353,N_11278);
nand U11812 (N_11812,N_11305,N_11327);
or U11813 (N_11813,N_11375,N_11363);
or U11814 (N_11814,N_11121,N_11348);
and U11815 (N_11815,N_11375,N_10989);
nand U11816 (N_11816,N_11019,N_11399);
and U11817 (N_11817,N_10910,N_11232);
nand U11818 (N_11818,N_11139,N_11347);
or U11819 (N_11819,N_10928,N_11222);
nor U11820 (N_11820,N_11092,N_11385);
nand U11821 (N_11821,N_11109,N_10800);
or U11822 (N_11822,N_11094,N_11231);
or U11823 (N_11823,N_11327,N_11134);
nand U11824 (N_11824,N_11200,N_11168);
nand U11825 (N_11825,N_10932,N_11245);
or U11826 (N_11826,N_10903,N_11309);
nor U11827 (N_11827,N_11102,N_11286);
nand U11828 (N_11828,N_10954,N_10994);
or U11829 (N_11829,N_11318,N_10814);
or U11830 (N_11830,N_11193,N_11016);
nand U11831 (N_11831,N_11189,N_10885);
nor U11832 (N_11832,N_10918,N_11010);
nor U11833 (N_11833,N_11087,N_10857);
or U11834 (N_11834,N_11064,N_10991);
nand U11835 (N_11835,N_11382,N_11370);
or U11836 (N_11836,N_11251,N_10995);
and U11837 (N_11837,N_11334,N_11266);
or U11838 (N_11838,N_10804,N_11293);
nand U11839 (N_11839,N_11093,N_10889);
or U11840 (N_11840,N_10991,N_10882);
or U11841 (N_11841,N_11031,N_11048);
and U11842 (N_11842,N_11156,N_11311);
nor U11843 (N_11843,N_11349,N_10892);
and U11844 (N_11844,N_11257,N_10976);
or U11845 (N_11845,N_10992,N_11384);
nand U11846 (N_11846,N_11305,N_11185);
nand U11847 (N_11847,N_11205,N_11064);
nor U11848 (N_11848,N_11293,N_11004);
nand U11849 (N_11849,N_11067,N_11276);
and U11850 (N_11850,N_11326,N_11307);
nor U11851 (N_11851,N_11147,N_10815);
nand U11852 (N_11852,N_10883,N_11035);
nand U11853 (N_11853,N_11151,N_10881);
nor U11854 (N_11854,N_10845,N_10851);
nor U11855 (N_11855,N_11059,N_11173);
or U11856 (N_11856,N_11040,N_11269);
or U11857 (N_11857,N_10839,N_11142);
or U11858 (N_11858,N_10895,N_11359);
nor U11859 (N_11859,N_11386,N_11044);
nand U11860 (N_11860,N_11195,N_11209);
or U11861 (N_11861,N_10983,N_10866);
nor U11862 (N_11862,N_10903,N_10843);
or U11863 (N_11863,N_11007,N_11199);
nor U11864 (N_11864,N_10850,N_10925);
nor U11865 (N_11865,N_10919,N_11200);
nand U11866 (N_11866,N_11238,N_11246);
or U11867 (N_11867,N_11080,N_11107);
nor U11868 (N_11868,N_11249,N_11306);
xnor U11869 (N_11869,N_11000,N_11123);
or U11870 (N_11870,N_11025,N_11083);
nand U11871 (N_11871,N_10975,N_10871);
and U11872 (N_11872,N_11025,N_11288);
and U11873 (N_11873,N_11338,N_11203);
nand U11874 (N_11874,N_11256,N_11283);
and U11875 (N_11875,N_10899,N_10905);
xnor U11876 (N_11876,N_10812,N_10824);
nand U11877 (N_11877,N_10849,N_11310);
or U11878 (N_11878,N_10948,N_11379);
or U11879 (N_11879,N_11259,N_11268);
and U11880 (N_11880,N_11089,N_11024);
nor U11881 (N_11881,N_10852,N_10972);
nand U11882 (N_11882,N_11152,N_11083);
nand U11883 (N_11883,N_10975,N_11309);
or U11884 (N_11884,N_11178,N_10983);
nor U11885 (N_11885,N_11280,N_11244);
nand U11886 (N_11886,N_10909,N_11333);
nor U11887 (N_11887,N_11093,N_10915);
or U11888 (N_11888,N_11156,N_11222);
nor U11889 (N_11889,N_10963,N_11313);
and U11890 (N_11890,N_11211,N_10942);
or U11891 (N_11891,N_11066,N_10881);
nand U11892 (N_11892,N_11161,N_11362);
or U11893 (N_11893,N_10838,N_10875);
and U11894 (N_11894,N_11160,N_10946);
and U11895 (N_11895,N_11083,N_11027);
nor U11896 (N_11896,N_11283,N_10922);
nor U11897 (N_11897,N_11061,N_11287);
nand U11898 (N_11898,N_11177,N_11313);
nand U11899 (N_11899,N_11204,N_11211);
nand U11900 (N_11900,N_11385,N_11018);
or U11901 (N_11901,N_11205,N_11072);
nand U11902 (N_11902,N_11047,N_11363);
nand U11903 (N_11903,N_11291,N_10802);
or U11904 (N_11904,N_10896,N_11207);
nand U11905 (N_11905,N_11105,N_10981);
nor U11906 (N_11906,N_10811,N_11072);
or U11907 (N_11907,N_11108,N_11232);
or U11908 (N_11908,N_11194,N_11214);
nor U11909 (N_11909,N_11118,N_11349);
or U11910 (N_11910,N_10810,N_11056);
and U11911 (N_11911,N_11149,N_10809);
nand U11912 (N_11912,N_11262,N_11124);
and U11913 (N_11913,N_11098,N_11138);
and U11914 (N_11914,N_11168,N_11127);
nor U11915 (N_11915,N_10881,N_11041);
and U11916 (N_11916,N_11085,N_10896);
and U11917 (N_11917,N_11076,N_10867);
and U11918 (N_11918,N_11279,N_11333);
nand U11919 (N_11919,N_10969,N_11068);
nand U11920 (N_11920,N_11184,N_11069);
nand U11921 (N_11921,N_11329,N_11260);
nand U11922 (N_11922,N_11079,N_11224);
nor U11923 (N_11923,N_11090,N_11267);
and U11924 (N_11924,N_11080,N_11071);
nor U11925 (N_11925,N_11035,N_11374);
nand U11926 (N_11926,N_10912,N_11232);
and U11927 (N_11927,N_11275,N_11153);
xor U11928 (N_11928,N_11279,N_11351);
and U11929 (N_11929,N_11230,N_10871);
or U11930 (N_11930,N_11050,N_11067);
or U11931 (N_11931,N_11232,N_11004);
and U11932 (N_11932,N_11193,N_11105);
or U11933 (N_11933,N_10905,N_11227);
xor U11934 (N_11934,N_10847,N_11327);
and U11935 (N_11935,N_11152,N_11208);
nor U11936 (N_11936,N_11107,N_11291);
nand U11937 (N_11937,N_11245,N_11018);
and U11938 (N_11938,N_11209,N_11246);
nor U11939 (N_11939,N_11095,N_11261);
nand U11940 (N_11940,N_11383,N_11352);
and U11941 (N_11941,N_10882,N_10958);
and U11942 (N_11942,N_10847,N_11131);
or U11943 (N_11943,N_11323,N_10942);
or U11944 (N_11944,N_10921,N_11048);
and U11945 (N_11945,N_10915,N_11306);
nand U11946 (N_11946,N_10862,N_11057);
nand U11947 (N_11947,N_11173,N_11044);
or U11948 (N_11948,N_11040,N_10851);
nand U11949 (N_11949,N_11114,N_10859);
nor U11950 (N_11950,N_10827,N_11359);
and U11951 (N_11951,N_10876,N_11039);
or U11952 (N_11952,N_11180,N_11070);
and U11953 (N_11953,N_11175,N_11013);
nand U11954 (N_11954,N_11233,N_11195);
nand U11955 (N_11955,N_11079,N_11066);
nand U11956 (N_11956,N_10988,N_11033);
and U11957 (N_11957,N_10977,N_10899);
nand U11958 (N_11958,N_11043,N_10885);
nand U11959 (N_11959,N_10879,N_11113);
nor U11960 (N_11960,N_11217,N_11078);
nand U11961 (N_11961,N_10873,N_11286);
nor U11962 (N_11962,N_11389,N_11336);
or U11963 (N_11963,N_11302,N_11299);
nand U11964 (N_11964,N_10902,N_10898);
and U11965 (N_11965,N_11061,N_10859);
or U11966 (N_11966,N_10802,N_11112);
or U11967 (N_11967,N_11034,N_11030);
and U11968 (N_11968,N_11175,N_11191);
or U11969 (N_11969,N_11108,N_10812);
nand U11970 (N_11970,N_11278,N_10837);
nand U11971 (N_11971,N_11241,N_11175);
nor U11972 (N_11972,N_11214,N_10900);
nor U11973 (N_11973,N_11076,N_11032);
nor U11974 (N_11974,N_11277,N_11135);
or U11975 (N_11975,N_10822,N_10808);
and U11976 (N_11976,N_10895,N_10919);
nand U11977 (N_11977,N_11270,N_11065);
nand U11978 (N_11978,N_11366,N_11365);
and U11979 (N_11979,N_11092,N_10986);
nand U11980 (N_11980,N_11384,N_11160);
nor U11981 (N_11981,N_11300,N_11069);
nand U11982 (N_11982,N_10962,N_10921);
nand U11983 (N_11983,N_11122,N_11063);
nor U11984 (N_11984,N_11319,N_10968);
nand U11985 (N_11985,N_11127,N_11113);
nor U11986 (N_11986,N_11051,N_10802);
nand U11987 (N_11987,N_10979,N_10877);
or U11988 (N_11988,N_10967,N_11170);
and U11989 (N_11989,N_11216,N_11240);
nand U11990 (N_11990,N_10984,N_11261);
and U11991 (N_11991,N_11023,N_11147);
or U11992 (N_11992,N_11186,N_11142);
or U11993 (N_11993,N_11252,N_10804);
or U11994 (N_11994,N_11175,N_10893);
nor U11995 (N_11995,N_11134,N_11042);
nand U11996 (N_11996,N_10813,N_11300);
or U11997 (N_11997,N_11092,N_11274);
nand U11998 (N_11998,N_11220,N_11280);
nand U11999 (N_11999,N_11217,N_11239);
nand U12000 (N_12000,N_11693,N_11652);
nor U12001 (N_12001,N_11773,N_11938);
nor U12002 (N_12002,N_11939,N_11797);
or U12003 (N_12003,N_11466,N_11803);
or U12004 (N_12004,N_11782,N_11855);
nand U12005 (N_12005,N_11557,N_11837);
nand U12006 (N_12006,N_11528,N_11794);
nor U12007 (N_12007,N_11669,N_11996);
nor U12008 (N_12008,N_11726,N_11920);
and U12009 (N_12009,N_11582,N_11640);
nor U12010 (N_12010,N_11744,N_11595);
and U12011 (N_12011,N_11403,N_11816);
nand U12012 (N_12012,N_11968,N_11845);
or U12013 (N_12013,N_11587,N_11596);
or U12014 (N_12014,N_11863,N_11432);
or U12015 (N_12015,N_11824,N_11676);
or U12016 (N_12016,N_11627,N_11666);
or U12017 (N_12017,N_11555,N_11830);
nor U12018 (N_12018,N_11672,N_11536);
and U12019 (N_12019,N_11565,N_11729);
and U12020 (N_12020,N_11420,N_11589);
and U12021 (N_12021,N_11493,N_11683);
nand U12022 (N_12022,N_11992,N_11561);
or U12023 (N_12023,N_11725,N_11911);
and U12024 (N_12024,N_11895,N_11500);
and U12025 (N_12025,N_11868,N_11784);
nor U12026 (N_12026,N_11808,N_11719);
or U12027 (N_12027,N_11846,N_11906);
and U12028 (N_12028,N_11749,N_11978);
or U12029 (N_12029,N_11825,N_11440);
or U12030 (N_12030,N_11711,N_11524);
nor U12031 (N_12031,N_11549,N_11513);
nand U12032 (N_12032,N_11748,N_11608);
and U12033 (N_12033,N_11701,N_11983);
and U12034 (N_12034,N_11780,N_11621);
nand U12035 (N_12035,N_11870,N_11722);
nor U12036 (N_12036,N_11497,N_11927);
nand U12037 (N_12037,N_11747,N_11932);
nand U12038 (N_12038,N_11743,N_11738);
nor U12039 (N_12039,N_11987,N_11761);
and U12040 (N_12040,N_11955,N_11572);
nand U12041 (N_12041,N_11428,N_11817);
nand U12042 (N_12042,N_11584,N_11698);
or U12043 (N_12043,N_11586,N_11919);
xor U12044 (N_12044,N_11455,N_11880);
or U12045 (N_12045,N_11883,N_11527);
and U12046 (N_12046,N_11574,N_11752);
nand U12047 (N_12047,N_11450,N_11998);
nor U12048 (N_12048,N_11723,N_11401);
nor U12049 (N_12049,N_11971,N_11551);
nand U12050 (N_12050,N_11771,N_11805);
nor U12051 (N_12051,N_11954,N_11459);
or U12052 (N_12052,N_11486,N_11688);
nor U12053 (N_12053,N_11661,N_11585);
xor U12054 (N_12054,N_11478,N_11458);
nor U12055 (N_12055,N_11984,N_11694);
and U12056 (N_12056,N_11490,N_11446);
nand U12057 (N_12057,N_11857,N_11681);
nand U12058 (N_12058,N_11542,N_11731);
or U12059 (N_12059,N_11734,N_11468);
nor U12060 (N_12060,N_11790,N_11579);
nand U12061 (N_12061,N_11961,N_11634);
nand U12062 (N_12062,N_11566,N_11519);
or U12063 (N_12063,N_11957,N_11687);
or U12064 (N_12064,N_11847,N_11736);
nand U12065 (N_12065,N_11943,N_11710);
nand U12066 (N_12066,N_11813,N_11503);
or U12067 (N_12067,N_11827,N_11496);
and U12068 (N_12068,N_11581,N_11509);
or U12069 (N_12069,N_11624,N_11473);
or U12070 (N_12070,N_11691,N_11707);
nor U12071 (N_12071,N_11484,N_11408);
xnor U12072 (N_12072,N_11946,N_11663);
or U12073 (N_12073,N_11461,N_11924);
or U12074 (N_12074,N_11603,N_11658);
or U12075 (N_12075,N_11424,N_11620);
nand U12076 (N_12076,N_11778,N_11914);
nor U12077 (N_12077,N_11618,N_11454);
xnor U12078 (N_12078,N_11575,N_11556);
and U12079 (N_12079,N_11717,N_11953);
and U12080 (N_12080,N_11779,N_11897);
and U12081 (N_12081,N_11560,N_11550);
xnor U12082 (N_12082,N_11737,N_11965);
nor U12083 (N_12083,N_11642,N_11653);
nor U12084 (N_12084,N_11951,N_11617);
and U12085 (N_12085,N_11430,N_11947);
and U12086 (N_12086,N_11421,N_11840);
nand U12087 (N_12087,N_11801,N_11606);
nor U12088 (N_12088,N_11604,N_11980);
nand U12089 (N_12089,N_11567,N_11525);
nand U12090 (N_12090,N_11460,N_11786);
and U12091 (N_12091,N_11487,N_11656);
or U12092 (N_12092,N_11732,N_11552);
nor U12093 (N_12093,N_11593,N_11592);
or U12094 (N_12094,N_11721,N_11940);
nand U12095 (N_12095,N_11760,N_11605);
nand U12096 (N_12096,N_11730,N_11886);
and U12097 (N_12097,N_11613,N_11819);
nand U12098 (N_12098,N_11495,N_11591);
or U12099 (N_12099,N_11999,N_11990);
or U12100 (N_12100,N_11501,N_11470);
or U12101 (N_12101,N_11506,N_11479);
and U12102 (N_12102,N_11809,N_11449);
nor U12103 (N_12103,N_11685,N_11912);
nand U12104 (N_12104,N_11896,N_11400);
nor U12105 (N_12105,N_11843,N_11643);
nand U12106 (N_12106,N_11772,N_11792);
xor U12107 (N_12107,N_11447,N_11714);
and U12108 (N_12108,N_11891,N_11783);
and U12109 (N_12109,N_11977,N_11664);
and U12110 (N_12110,N_11851,N_11807);
or U12111 (N_12111,N_11435,N_11644);
or U12112 (N_12112,N_11662,N_11504);
nand U12113 (N_12113,N_11646,N_11443);
or U12114 (N_12114,N_11937,N_11964);
nor U12115 (N_12115,N_11692,N_11485);
nand U12116 (N_12116,N_11654,N_11795);
nand U12117 (N_12117,N_11768,N_11770);
nand U12118 (N_12118,N_11690,N_11625);
or U12119 (N_12119,N_11793,N_11464);
or U12120 (N_12120,N_11724,N_11594);
and U12121 (N_12121,N_11423,N_11728);
nand U12122 (N_12122,N_11888,N_11706);
xnor U12123 (N_12123,N_11571,N_11425);
and U12124 (N_12124,N_11414,N_11601);
and U12125 (N_12125,N_11563,N_11881);
and U12126 (N_12126,N_11925,N_11441);
nand U12127 (N_12127,N_11649,N_11507);
xnor U12128 (N_12128,N_11900,N_11814);
or U12129 (N_12129,N_11452,N_11609);
and U12130 (N_12130,N_11806,N_11885);
nor U12131 (N_12131,N_11568,N_11573);
nor U12132 (N_12132,N_11483,N_11869);
nor U12133 (N_12133,N_11993,N_11530);
and U12134 (N_12134,N_11890,N_11988);
nand U12135 (N_12135,N_11766,N_11742);
and U12136 (N_12136,N_11774,N_11765);
nor U12137 (N_12137,N_11826,N_11769);
nand U12138 (N_12138,N_11926,N_11510);
or U12139 (N_12139,N_11610,N_11789);
nor U12140 (N_12140,N_11482,N_11451);
and U12141 (N_12141,N_11626,N_11907);
and U12142 (N_12142,N_11462,N_11402);
or U12143 (N_12143,N_11558,N_11602);
or U12144 (N_12144,N_11523,N_11995);
or U12145 (N_12145,N_11439,N_11829);
and U12146 (N_12146,N_11657,N_11989);
nor U12147 (N_12147,N_11514,N_11823);
or U12148 (N_12148,N_11491,N_11410);
nor U12149 (N_12149,N_11429,N_11545);
nor U12150 (N_12150,N_11546,N_11614);
or U12151 (N_12151,N_11815,N_11970);
or U12152 (N_12152,N_11583,N_11835);
nor U12153 (N_12153,N_11850,N_11628);
nor U12154 (N_12154,N_11569,N_11442);
nor U12155 (N_12155,N_11413,N_11739);
or U12156 (N_12156,N_11667,N_11876);
or U12157 (N_12157,N_11671,N_11629);
or U12158 (N_12158,N_11437,N_11521);
or U12159 (N_12159,N_11818,N_11810);
or U12160 (N_12160,N_11856,N_11598);
and U12161 (N_12161,N_11419,N_11522);
or U12162 (N_12162,N_11705,N_11944);
nor U12163 (N_12163,N_11875,N_11704);
xnor U12164 (N_12164,N_11526,N_11878);
nand U12165 (N_12165,N_11758,N_11637);
nand U12166 (N_12166,N_11918,N_11882);
and U12167 (N_12167,N_11933,N_11456);
and U12168 (N_12168,N_11763,N_11909);
or U12169 (N_12169,N_11849,N_11991);
or U12170 (N_12170,N_11848,N_11787);
nand U12171 (N_12171,N_11679,N_11969);
or U12172 (N_12172,N_11820,N_11502);
or U12173 (N_12173,N_11928,N_11630);
xor U12174 (N_12174,N_11684,N_11675);
nor U12175 (N_12175,N_11406,N_11518);
nor U12176 (N_12176,N_11699,N_11828);
nand U12177 (N_12177,N_11917,N_11975);
and U12178 (N_12178,N_11547,N_11804);
nand U12179 (N_12179,N_11543,N_11821);
nand U12180 (N_12180,N_11570,N_11979);
or U12181 (N_12181,N_11788,N_11910);
or U12182 (N_12182,N_11615,N_11822);
nor U12183 (N_12183,N_11686,N_11751);
or U12184 (N_12184,N_11986,N_11877);
or U12185 (N_12185,N_11967,N_11445);
or U12186 (N_12186,N_11715,N_11494);
or U12187 (N_12187,N_11444,N_11641);
nand U12188 (N_12188,N_11905,N_11873);
nand U12189 (N_12189,N_11492,N_11645);
nor U12190 (N_12190,N_11713,N_11405);
or U12191 (N_12191,N_11916,N_11678);
and U12192 (N_12192,N_11866,N_11677);
nand U12193 (N_12193,N_11887,N_11942);
nand U12194 (N_12194,N_11682,N_11665);
or U12195 (N_12195,N_11475,N_11799);
nand U12196 (N_12196,N_11517,N_11532);
nand U12197 (N_12197,N_11703,N_11931);
nor U12198 (N_12198,N_11436,N_11913);
and U12199 (N_12199,N_11673,N_11791);
nor U12200 (N_12200,N_11963,N_11562);
nor U12201 (N_12201,N_11884,N_11901);
or U12202 (N_12202,N_11915,N_11894);
nand U12203 (N_12203,N_11499,N_11936);
nor U12204 (N_12204,N_11531,N_11670);
nor U12205 (N_12205,N_11867,N_11520);
nand U12206 (N_12206,N_11861,N_11839);
nand U12207 (N_12207,N_11639,N_11930);
nand U12208 (N_12208,N_11636,N_11638);
or U12209 (N_12209,N_11535,N_11776);
and U12210 (N_12210,N_11465,N_11655);
nand U12211 (N_12211,N_11841,N_11689);
nor U12212 (N_12212,N_11767,N_11854);
or U12213 (N_12213,N_11529,N_11541);
nor U12214 (N_12214,N_11929,N_11700);
or U12215 (N_12215,N_11785,N_11702);
and U12216 (N_12216,N_11576,N_11812);
nand U12217 (N_12217,N_11860,N_11746);
and U12218 (N_12218,N_11834,N_11696);
nor U12219 (N_12219,N_11733,N_11457);
nor U12220 (N_12220,N_11588,N_11600);
nand U12221 (N_12221,N_11564,N_11754);
or U12222 (N_12222,N_11775,N_11431);
nor U12223 (N_12223,N_11833,N_11720);
nand U12224 (N_12224,N_11852,N_11966);
nand U12225 (N_12225,N_11434,N_11505);
or U12226 (N_12226,N_11416,N_11802);
nand U12227 (N_12227,N_11427,N_11537);
and U12228 (N_12228,N_11959,N_11836);
nand U12229 (N_12229,N_11798,N_11515);
nand U12230 (N_12230,N_11659,N_11553);
or U12231 (N_12231,N_11544,N_11548);
and U12232 (N_12232,N_11859,N_11472);
nor U12233 (N_12233,N_11612,N_11512);
and U12234 (N_12234,N_11976,N_11635);
or U12235 (N_12235,N_11477,N_11889);
nor U12236 (N_12236,N_11874,N_11745);
nor U12237 (N_12237,N_11781,N_11853);
nor U12238 (N_12238,N_11862,N_11762);
nor U12239 (N_12239,N_11879,N_11467);
nor U12240 (N_12240,N_11476,N_11488);
or U12241 (N_12241,N_11973,N_11871);
nand U12242 (N_12242,N_11577,N_11463);
and U12243 (N_12243,N_11534,N_11741);
nand U12244 (N_12244,N_11540,N_11622);
or U12245 (N_12245,N_11756,N_11831);
nor U12246 (N_12246,N_11453,N_11578);
or U12247 (N_12247,N_11415,N_11921);
nand U12248 (N_12248,N_11718,N_11632);
and U12249 (N_12249,N_11412,N_11948);
nand U12250 (N_12250,N_11433,N_11872);
and U12251 (N_12251,N_11796,N_11607);
nor U12252 (N_12252,N_11864,N_11508);
and U12253 (N_12253,N_11404,N_11935);
nand U12254 (N_12254,N_11709,N_11716);
or U12255 (N_12255,N_11899,N_11838);
and U12256 (N_12256,N_11811,N_11750);
nand U12257 (N_12257,N_11660,N_11865);
and U12258 (N_12258,N_11904,N_11777);
and U12259 (N_12259,N_11407,N_11941);
nand U12260 (N_12260,N_11481,N_11902);
and U12261 (N_12261,N_11599,N_11903);
and U12262 (N_12262,N_11832,N_11893);
or U12263 (N_12263,N_11934,N_11708);
nand U12264 (N_12264,N_11764,N_11960);
and U12265 (N_12265,N_11974,N_11997);
nor U12266 (N_12266,N_11538,N_11511);
nand U12267 (N_12267,N_11554,N_11908);
nor U12268 (N_12268,N_11712,N_11958);
nor U12269 (N_12269,N_11674,N_11489);
nand U12270 (N_12270,N_11922,N_11498);
or U12271 (N_12271,N_11409,N_11757);
and U12272 (N_12272,N_11580,N_11753);
nor U12273 (N_12273,N_11981,N_11471);
or U12274 (N_12274,N_11945,N_11755);
nand U12275 (N_12275,N_11623,N_11619);
nand U12276 (N_12276,N_11898,N_11631);
nand U12277 (N_12277,N_11735,N_11956);
nor U12278 (N_12278,N_11411,N_11844);
or U12279 (N_12279,N_11533,N_11469);
nor U12280 (N_12280,N_11448,N_11994);
xor U12281 (N_12281,N_11616,N_11480);
and U12282 (N_12282,N_11727,N_11516);
nor U12283 (N_12283,N_11842,N_11438);
nand U12284 (N_12284,N_11647,N_11611);
nand U12285 (N_12285,N_11759,N_11648);
or U12286 (N_12286,N_11982,N_11892);
or U12287 (N_12287,N_11590,N_11559);
or U12288 (N_12288,N_11651,N_11418);
nor U12289 (N_12289,N_11950,N_11952);
nand U12290 (N_12290,N_11923,N_11800);
nor U12291 (N_12291,N_11474,N_11417);
or U12292 (N_12292,N_11740,N_11650);
nand U12293 (N_12293,N_11949,N_11633);
nand U12294 (N_12294,N_11972,N_11695);
nand U12295 (N_12295,N_11426,N_11539);
xnor U12296 (N_12296,N_11680,N_11962);
or U12297 (N_12297,N_11668,N_11697);
or U12298 (N_12298,N_11985,N_11858);
nor U12299 (N_12299,N_11422,N_11597);
or U12300 (N_12300,N_11413,N_11419);
nand U12301 (N_12301,N_11751,N_11776);
nor U12302 (N_12302,N_11946,N_11858);
nor U12303 (N_12303,N_11817,N_11447);
or U12304 (N_12304,N_11419,N_11430);
nand U12305 (N_12305,N_11868,N_11871);
and U12306 (N_12306,N_11447,N_11636);
or U12307 (N_12307,N_11462,N_11447);
nor U12308 (N_12308,N_11620,N_11897);
nand U12309 (N_12309,N_11633,N_11599);
nand U12310 (N_12310,N_11803,N_11425);
nor U12311 (N_12311,N_11799,N_11716);
and U12312 (N_12312,N_11890,N_11565);
nand U12313 (N_12313,N_11432,N_11513);
or U12314 (N_12314,N_11505,N_11433);
nand U12315 (N_12315,N_11760,N_11928);
nand U12316 (N_12316,N_11987,N_11961);
nor U12317 (N_12317,N_11558,N_11922);
nand U12318 (N_12318,N_11587,N_11564);
and U12319 (N_12319,N_11683,N_11571);
nand U12320 (N_12320,N_11566,N_11464);
or U12321 (N_12321,N_11480,N_11624);
and U12322 (N_12322,N_11567,N_11897);
or U12323 (N_12323,N_11687,N_11493);
nor U12324 (N_12324,N_11998,N_11872);
nor U12325 (N_12325,N_11442,N_11950);
nand U12326 (N_12326,N_11598,N_11513);
or U12327 (N_12327,N_11464,N_11857);
or U12328 (N_12328,N_11928,N_11607);
nand U12329 (N_12329,N_11598,N_11504);
and U12330 (N_12330,N_11724,N_11949);
and U12331 (N_12331,N_11559,N_11555);
xnor U12332 (N_12332,N_11750,N_11911);
or U12333 (N_12333,N_11874,N_11703);
or U12334 (N_12334,N_11401,N_11834);
or U12335 (N_12335,N_11601,N_11906);
nor U12336 (N_12336,N_11642,N_11881);
nor U12337 (N_12337,N_11600,N_11408);
or U12338 (N_12338,N_11872,N_11755);
nor U12339 (N_12339,N_11746,N_11994);
and U12340 (N_12340,N_11653,N_11447);
nor U12341 (N_12341,N_11734,N_11467);
or U12342 (N_12342,N_11592,N_11837);
nor U12343 (N_12343,N_11540,N_11437);
nor U12344 (N_12344,N_11518,N_11632);
nor U12345 (N_12345,N_11598,N_11677);
nand U12346 (N_12346,N_11650,N_11612);
nand U12347 (N_12347,N_11892,N_11710);
or U12348 (N_12348,N_11766,N_11805);
and U12349 (N_12349,N_11434,N_11946);
and U12350 (N_12350,N_11638,N_11542);
nor U12351 (N_12351,N_11562,N_11926);
nor U12352 (N_12352,N_11723,N_11850);
nor U12353 (N_12353,N_11905,N_11696);
xor U12354 (N_12354,N_11685,N_11640);
nor U12355 (N_12355,N_11458,N_11485);
nand U12356 (N_12356,N_11806,N_11949);
and U12357 (N_12357,N_11655,N_11450);
or U12358 (N_12358,N_11735,N_11703);
and U12359 (N_12359,N_11589,N_11972);
nand U12360 (N_12360,N_11950,N_11768);
nand U12361 (N_12361,N_11938,N_11901);
or U12362 (N_12362,N_11700,N_11975);
or U12363 (N_12363,N_11584,N_11784);
nor U12364 (N_12364,N_11631,N_11583);
nor U12365 (N_12365,N_11854,N_11906);
or U12366 (N_12366,N_11613,N_11986);
nor U12367 (N_12367,N_11649,N_11683);
or U12368 (N_12368,N_11427,N_11790);
and U12369 (N_12369,N_11462,N_11675);
nand U12370 (N_12370,N_11875,N_11699);
nand U12371 (N_12371,N_11854,N_11632);
nand U12372 (N_12372,N_11458,N_11799);
and U12373 (N_12373,N_11646,N_11537);
or U12374 (N_12374,N_11883,N_11627);
nor U12375 (N_12375,N_11670,N_11781);
nor U12376 (N_12376,N_11439,N_11699);
or U12377 (N_12377,N_11902,N_11664);
xnor U12378 (N_12378,N_11704,N_11565);
or U12379 (N_12379,N_11990,N_11961);
or U12380 (N_12380,N_11793,N_11758);
or U12381 (N_12381,N_11625,N_11473);
nand U12382 (N_12382,N_11856,N_11517);
or U12383 (N_12383,N_11888,N_11733);
xor U12384 (N_12384,N_11760,N_11611);
nor U12385 (N_12385,N_11754,N_11678);
nor U12386 (N_12386,N_11999,N_11460);
nand U12387 (N_12387,N_11944,N_11684);
and U12388 (N_12388,N_11777,N_11738);
nor U12389 (N_12389,N_11910,N_11913);
and U12390 (N_12390,N_11457,N_11816);
or U12391 (N_12391,N_11499,N_11845);
nand U12392 (N_12392,N_11849,N_11672);
or U12393 (N_12393,N_11818,N_11632);
and U12394 (N_12394,N_11527,N_11564);
xnor U12395 (N_12395,N_11890,N_11521);
nor U12396 (N_12396,N_11530,N_11453);
nor U12397 (N_12397,N_11420,N_11692);
nor U12398 (N_12398,N_11500,N_11543);
nor U12399 (N_12399,N_11952,N_11742);
or U12400 (N_12400,N_11675,N_11933);
and U12401 (N_12401,N_11894,N_11804);
and U12402 (N_12402,N_11619,N_11950);
or U12403 (N_12403,N_11436,N_11506);
and U12404 (N_12404,N_11953,N_11601);
and U12405 (N_12405,N_11469,N_11877);
and U12406 (N_12406,N_11943,N_11971);
and U12407 (N_12407,N_11681,N_11719);
nand U12408 (N_12408,N_11620,N_11837);
nand U12409 (N_12409,N_11690,N_11888);
or U12410 (N_12410,N_11922,N_11989);
nor U12411 (N_12411,N_11877,N_11968);
nor U12412 (N_12412,N_11692,N_11448);
or U12413 (N_12413,N_11988,N_11955);
xnor U12414 (N_12414,N_11415,N_11882);
xor U12415 (N_12415,N_11527,N_11472);
and U12416 (N_12416,N_11811,N_11932);
nor U12417 (N_12417,N_11679,N_11734);
and U12418 (N_12418,N_11813,N_11475);
and U12419 (N_12419,N_11433,N_11468);
nand U12420 (N_12420,N_11672,N_11422);
or U12421 (N_12421,N_11815,N_11543);
nor U12422 (N_12422,N_11627,N_11546);
nor U12423 (N_12423,N_11576,N_11704);
or U12424 (N_12424,N_11559,N_11864);
or U12425 (N_12425,N_11618,N_11791);
nor U12426 (N_12426,N_11566,N_11604);
or U12427 (N_12427,N_11738,N_11599);
nand U12428 (N_12428,N_11439,N_11785);
or U12429 (N_12429,N_11696,N_11917);
or U12430 (N_12430,N_11712,N_11692);
or U12431 (N_12431,N_11873,N_11490);
nor U12432 (N_12432,N_11725,N_11917);
or U12433 (N_12433,N_11552,N_11733);
or U12434 (N_12434,N_11967,N_11936);
and U12435 (N_12435,N_11513,N_11689);
and U12436 (N_12436,N_11851,N_11760);
nand U12437 (N_12437,N_11971,N_11662);
nor U12438 (N_12438,N_11421,N_11998);
or U12439 (N_12439,N_11828,N_11486);
nor U12440 (N_12440,N_11586,N_11727);
or U12441 (N_12441,N_11875,N_11450);
and U12442 (N_12442,N_11698,N_11434);
nand U12443 (N_12443,N_11545,N_11666);
and U12444 (N_12444,N_11938,N_11657);
nand U12445 (N_12445,N_11938,N_11888);
or U12446 (N_12446,N_11655,N_11912);
or U12447 (N_12447,N_11536,N_11933);
nor U12448 (N_12448,N_11546,N_11400);
nand U12449 (N_12449,N_11799,N_11586);
and U12450 (N_12450,N_11814,N_11545);
or U12451 (N_12451,N_11837,N_11608);
nor U12452 (N_12452,N_11434,N_11723);
or U12453 (N_12453,N_11424,N_11567);
and U12454 (N_12454,N_11891,N_11753);
or U12455 (N_12455,N_11800,N_11628);
nand U12456 (N_12456,N_11832,N_11527);
or U12457 (N_12457,N_11540,N_11831);
nor U12458 (N_12458,N_11528,N_11825);
or U12459 (N_12459,N_11663,N_11801);
and U12460 (N_12460,N_11743,N_11908);
nand U12461 (N_12461,N_11404,N_11955);
and U12462 (N_12462,N_11886,N_11757);
and U12463 (N_12463,N_11899,N_11598);
nor U12464 (N_12464,N_11593,N_11755);
or U12465 (N_12465,N_11818,N_11854);
nand U12466 (N_12466,N_11952,N_11408);
nor U12467 (N_12467,N_11940,N_11634);
nand U12468 (N_12468,N_11485,N_11767);
nor U12469 (N_12469,N_11715,N_11849);
nand U12470 (N_12470,N_11427,N_11556);
nor U12471 (N_12471,N_11796,N_11981);
nand U12472 (N_12472,N_11992,N_11875);
or U12473 (N_12473,N_11933,N_11736);
nand U12474 (N_12474,N_11845,N_11439);
and U12475 (N_12475,N_11539,N_11418);
nor U12476 (N_12476,N_11947,N_11905);
or U12477 (N_12477,N_11662,N_11541);
and U12478 (N_12478,N_11616,N_11809);
and U12479 (N_12479,N_11918,N_11964);
and U12480 (N_12480,N_11896,N_11749);
nor U12481 (N_12481,N_11566,N_11456);
nor U12482 (N_12482,N_11844,N_11858);
and U12483 (N_12483,N_11882,N_11402);
nor U12484 (N_12484,N_11794,N_11753);
xor U12485 (N_12485,N_11977,N_11593);
nand U12486 (N_12486,N_11446,N_11827);
nand U12487 (N_12487,N_11758,N_11674);
nand U12488 (N_12488,N_11425,N_11482);
or U12489 (N_12489,N_11872,N_11888);
nand U12490 (N_12490,N_11819,N_11713);
or U12491 (N_12491,N_11451,N_11573);
nor U12492 (N_12492,N_11783,N_11713);
and U12493 (N_12493,N_11668,N_11536);
nor U12494 (N_12494,N_11830,N_11547);
and U12495 (N_12495,N_11659,N_11570);
or U12496 (N_12496,N_11432,N_11947);
or U12497 (N_12497,N_11894,N_11401);
and U12498 (N_12498,N_11560,N_11844);
nand U12499 (N_12499,N_11606,N_11736);
or U12500 (N_12500,N_11885,N_11844);
nor U12501 (N_12501,N_11599,N_11777);
or U12502 (N_12502,N_11942,N_11423);
and U12503 (N_12503,N_11761,N_11696);
nand U12504 (N_12504,N_11629,N_11445);
nor U12505 (N_12505,N_11902,N_11428);
or U12506 (N_12506,N_11899,N_11609);
nand U12507 (N_12507,N_11746,N_11498);
nand U12508 (N_12508,N_11521,N_11493);
or U12509 (N_12509,N_11981,N_11866);
nor U12510 (N_12510,N_11917,N_11791);
nor U12511 (N_12511,N_11746,N_11902);
nand U12512 (N_12512,N_11919,N_11732);
and U12513 (N_12513,N_11991,N_11939);
nor U12514 (N_12514,N_11666,N_11980);
and U12515 (N_12515,N_11907,N_11850);
nor U12516 (N_12516,N_11552,N_11781);
or U12517 (N_12517,N_11490,N_11959);
nand U12518 (N_12518,N_11816,N_11664);
or U12519 (N_12519,N_11640,N_11644);
nand U12520 (N_12520,N_11977,N_11492);
and U12521 (N_12521,N_11532,N_11692);
nor U12522 (N_12522,N_11601,N_11574);
nor U12523 (N_12523,N_11825,N_11515);
or U12524 (N_12524,N_11635,N_11408);
nor U12525 (N_12525,N_11904,N_11467);
nor U12526 (N_12526,N_11563,N_11941);
nor U12527 (N_12527,N_11744,N_11601);
nand U12528 (N_12528,N_11513,N_11872);
nand U12529 (N_12529,N_11405,N_11791);
nor U12530 (N_12530,N_11717,N_11744);
nor U12531 (N_12531,N_11546,N_11577);
or U12532 (N_12532,N_11491,N_11889);
and U12533 (N_12533,N_11402,N_11655);
and U12534 (N_12534,N_11933,N_11823);
and U12535 (N_12535,N_11511,N_11962);
nor U12536 (N_12536,N_11854,N_11808);
and U12537 (N_12537,N_11986,N_11483);
or U12538 (N_12538,N_11712,N_11452);
and U12539 (N_12539,N_11664,N_11712);
or U12540 (N_12540,N_11702,N_11673);
nand U12541 (N_12541,N_11732,N_11729);
nand U12542 (N_12542,N_11988,N_11606);
and U12543 (N_12543,N_11795,N_11415);
and U12544 (N_12544,N_11534,N_11676);
nor U12545 (N_12545,N_11857,N_11610);
nand U12546 (N_12546,N_11997,N_11714);
and U12547 (N_12547,N_11715,N_11521);
nor U12548 (N_12548,N_11559,N_11787);
and U12549 (N_12549,N_11750,N_11485);
and U12550 (N_12550,N_11520,N_11971);
nor U12551 (N_12551,N_11988,N_11474);
or U12552 (N_12552,N_11567,N_11486);
and U12553 (N_12553,N_11871,N_11782);
nand U12554 (N_12554,N_11790,N_11949);
or U12555 (N_12555,N_11809,N_11618);
nand U12556 (N_12556,N_11469,N_11785);
nand U12557 (N_12557,N_11919,N_11528);
and U12558 (N_12558,N_11683,N_11709);
nand U12559 (N_12559,N_11960,N_11800);
nor U12560 (N_12560,N_11934,N_11646);
nand U12561 (N_12561,N_11477,N_11688);
and U12562 (N_12562,N_11527,N_11869);
nand U12563 (N_12563,N_11828,N_11559);
xor U12564 (N_12564,N_11832,N_11938);
nand U12565 (N_12565,N_11691,N_11446);
and U12566 (N_12566,N_11400,N_11634);
and U12567 (N_12567,N_11918,N_11746);
and U12568 (N_12568,N_11896,N_11601);
and U12569 (N_12569,N_11884,N_11447);
nor U12570 (N_12570,N_11891,N_11403);
and U12571 (N_12571,N_11700,N_11999);
and U12572 (N_12572,N_11571,N_11947);
nand U12573 (N_12573,N_11890,N_11444);
and U12574 (N_12574,N_11931,N_11452);
nand U12575 (N_12575,N_11583,N_11855);
xor U12576 (N_12576,N_11869,N_11992);
and U12577 (N_12577,N_11849,N_11576);
and U12578 (N_12578,N_11419,N_11697);
or U12579 (N_12579,N_11558,N_11449);
or U12580 (N_12580,N_11999,N_11964);
or U12581 (N_12581,N_11499,N_11542);
or U12582 (N_12582,N_11987,N_11638);
nor U12583 (N_12583,N_11872,N_11962);
nor U12584 (N_12584,N_11745,N_11402);
and U12585 (N_12585,N_11697,N_11488);
or U12586 (N_12586,N_11638,N_11735);
nand U12587 (N_12587,N_11762,N_11511);
nor U12588 (N_12588,N_11814,N_11993);
nand U12589 (N_12589,N_11595,N_11811);
nand U12590 (N_12590,N_11879,N_11619);
nand U12591 (N_12591,N_11664,N_11656);
and U12592 (N_12592,N_11458,N_11990);
nand U12593 (N_12593,N_11619,N_11911);
or U12594 (N_12594,N_11589,N_11876);
nand U12595 (N_12595,N_11542,N_11548);
or U12596 (N_12596,N_11437,N_11493);
nand U12597 (N_12597,N_11687,N_11461);
nand U12598 (N_12598,N_11569,N_11810);
nor U12599 (N_12599,N_11896,N_11564);
nand U12600 (N_12600,N_12510,N_12148);
or U12601 (N_12601,N_12251,N_12222);
and U12602 (N_12602,N_12257,N_12368);
and U12603 (N_12603,N_12339,N_12562);
and U12604 (N_12604,N_12460,N_12202);
nor U12605 (N_12605,N_12144,N_12367);
nor U12606 (N_12606,N_12082,N_12231);
or U12607 (N_12607,N_12513,N_12407);
nand U12608 (N_12608,N_12312,N_12211);
nor U12609 (N_12609,N_12084,N_12459);
or U12610 (N_12610,N_12261,N_12524);
nor U12611 (N_12611,N_12110,N_12100);
nor U12612 (N_12612,N_12147,N_12160);
or U12613 (N_12613,N_12479,N_12493);
nor U12614 (N_12614,N_12187,N_12370);
nor U12615 (N_12615,N_12078,N_12131);
nand U12616 (N_12616,N_12363,N_12327);
nand U12617 (N_12617,N_12039,N_12053);
nor U12618 (N_12618,N_12549,N_12530);
nor U12619 (N_12619,N_12470,N_12298);
or U12620 (N_12620,N_12263,N_12528);
nor U12621 (N_12621,N_12595,N_12518);
xnor U12622 (N_12622,N_12324,N_12168);
or U12623 (N_12623,N_12041,N_12464);
or U12624 (N_12624,N_12394,N_12296);
and U12625 (N_12625,N_12121,N_12300);
nand U12626 (N_12626,N_12031,N_12564);
and U12627 (N_12627,N_12097,N_12319);
or U12628 (N_12628,N_12467,N_12068);
and U12629 (N_12629,N_12204,N_12125);
and U12630 (N_12630,N_12259,N_12405);
nand U12631 (N_12631,N_12194,N_12551);
nor U12632 (N_12632,N_12005,N_12027);
nor U12633 (N_12633,N_12042,N_12426);
or U12634 (N_12634,N_12448,N_12278);
or U12635 (N_12635,N_12580,N_12219);
or U12636 (N_12636,N_12072,N_12353);
and U12637 (N_12637,N_12279,N_12250);
nor U12638 (N_12638,N_12019,N_12299);
xnor U12639 (N_12639,N_12489,N_12152);
or U12640 (N_12640,N_12526,N_12445);
nor U12641 (N_12641,N_12566,N_12588);
nand U12642 (N_12642,N_12054,N_12589);
nor U12643 (N_12643,N_12456,N_12217);
and U12644 (N_12644,N_12401,N_12535);
or U12645 (N_12645,N_12547,N_12276);
xnor U12646 (N_12646,N_12396,N_12398);
nand U12647 (N_12647,N_12375,N_12506);
or U12648 (N_12648,N_12335,N_12040);
and U12649 (N_12649,N_12377,N_12007);
or U12650 (N_12650,N_12229,N_12343);
nor U12651 (N_12651,N_12453,N_12381);
and U12652 (N_12652,N_12388,N_12461);
and U12653 (N_12653,N_12362,N_12124);
or U12654 (N_12654,N_12395,N_12013);
or U12655 (N_12655,N_12273,N_12378);
or U12656 (N_12656,N_12102,N_12272);
or U12657 (N_12657,N_12289,N_12006);
and U12658 (N_12658,N_12174,N_12206);
or U12659 (N_12659,N_12157,N_12421);
and U12660 (N_12660,N_12063,N_12200);
and U12661 (N_12661,N_12010,N_12462);
nand U12662 (N_12662,N_12351,N_12075);
nor U12663 (N_12663,N_12226,N_12244);
or U12664 (N_12664,N_12403,N_12391);
and U12665 (N_12665,N_12062,N_12357);
or U12666 (N_12666,N_12466,N_12109);
or U12667 (N_12667,N_12049,N_12000);
or U12668 (N_12668,N_12571,N_12503);
and U12669 (N_12669,N_12590,N_12587);
or U12670 (N_12670,N_12491,N_12267);
nor U12671 (N_12671,N_12163,N_12034);
and U12672 (N_12672,N_12140,N_12112);
and U12673 (N_12673,N_12020,N_12582);
and U12674 (N_12674,N_12585,N_12220);
nand U12675 (N_12675,N_12099,N_12282);
or U12676 (N_12676,N_12520,N_12365);
and U12677 (N_12677,N_12500,N_12234);
nor U12678 (N_12678,N_12314,N_12225);
nor U12679 (N_12679,N_12207,N_12149);
and U12680 (N_12680,N_12419,N_12090);
nor U12681 (N_12681,N_12344,N_12292);
and U12682 (N_12682,N_12281,N_12138);
nor U12683 (N_12683,N_12498,N_12565);
nor U12684 (N_12684,N_12169,N_12508);
xor U12685 (N_12685,N_12228,N_12095);
nor U12686 (N_12686,N_12457,N_12155);
and U12687 (N_12687,N_12232,N_12141);
or U12688 (N_12688,N_12023,N_12531);
nand U12689 (N_12689,N_12570,N_12258);
and U12690 (N_12690,N_12191,N_12360);
or U12691 (N_12691,N_12444,N_12047);
and U12692 (N_12692,N_12304,N_12196);
nand U12693 (N_12693,N_12540,N_12178);
nand U12694 (N_12694,N_12323,N_12165);
or U12695 (N_12695,N_12415,N_12235);
nor U12696 (N_12696,N_12208,N_12372);
nor U12697 (N_12697,N_12071,N_12076);
or U12698 (N_12698,N_12497,N_12573);
or U12699 (N_12699,N_12424,N_12598);
nor U12700 (N_12700,N_12086,N_12043);
nand U12701 (N_12701,N_12478,N_12432);
nor U12702 (N_12702,N_12104,N_12030);
or U12703 (N_12703,N_12472,N_12067);
nor U12704 (N_12704,N_12545,N_12354);
nor U12705 (N_12705,N_12009,N_12516);
and U12706 (N_12706,N_12065,N_12369);
nor U12707 (N_12707,N_12105,N_12091);
nor U12708 (N_12708,N_12488,N_12197);
xor U12709 (N_12709,N_12532,N_12429);
or U12710 (N_12710,N_12523,N_12213);
or U12711 (N_12711,N_12242,N_12449);
or U12712 (N_12712,N_12212,N_12115);
or U12713 (N_12713,N_12318,N_12249);
nor U12714 (N_12714,N_12546,N_12463);
and U12715 (N_12715,N_12195,N_12575);
or U12716 (N_12716,N_12237,N_12413);
or U12717 (N_12717,N_12128,N_12172);
and U12718 (N_12718,N_12061,N_12480);
nor U12719 (N_12719,N_12294,N_12297);
nor U12720 (N_12720,N_12270,N_12440);
nand U12721 (N_12721,N_12153,N_12451);
and U12722 (N_12722,N_12166,N_12181);
nand U12723 (N_12723,N_12179,N_12502);
and U12724 (N_12724,N_12268,N_12120);
nor U12725 (N_12725,N_12476,N_12118);
nor U12726 (N_12726,N_12356,N_12254);
and U12727 (N_12727,N_12406,N_12494);
nand U12728 (N_12728,N_12058,N_12156);
or U12729 (N_12729,N_12239,N_12435);
or U12730 (N_12730,N_12064,N_12586);
nor U12731 (N_12731,N_12055,N_12527);
or U12732 (N_12732,N_12085,N_12584);
and U12733 (N_12733,N_12485,N_12262);
nand U12734 (N_12734,N_12114,N_12486);
nand U12735 (N_12735,N_12490,N_12216);
nor U12736 (N_12736,N_12233,N_12142);
or U12737 (N_12737,N_12317,N_12230);
or U12738 (N_12738,N_12224,N_12384);
nor U12739 (N_12739,N_12350,N_12143);
nor U12740 (N_12740,N_12046,N_12409);
or U12741 (N_12741,N_12550,N_12596);
or U12742 (N_12742,N_12519,N_12471);
nor U12743 (N_12743,N_12180,N_12495);
or U12744 (N_12744,N_12175,N_12420);
or U12745 (N_12745,N_12475,N_12011);
nor U12746 (N_12746,N_12022,N_12411);
and U12747 (N_12747,N_12277,N_12008);
nand U12748 (N_12748,N_12484,N_12126);
nor U12749 (N_12749,N_12438,N_12223);
or U12750 (N_12750,N_12482,N_12477);
nor U12751 (N_12751,N_12132,N_12539);
nand U12752 (N_12752,N_12248,N_12521);
and U12753 (N_12753,N_12400,N_12364);
nand U12754 (N_12754,N_12271,N_12321);
nand U12755 (N_12755,N_12433,N_12492);
or U12756 (N_12756,N_12410,N_12417);
nand U12757 (N_12757,N_12517,N_12560);
nor U12758 (N_12758,N_12119,N_12569);
nor U12759 (N_12759,N_12285,N_12541);
xor U12760 (N_12760,N_12103,N_12483);
nor U12761 (N_12761,N_12499,N_12003);
nor U12762 (N_12762,N_12515,N_12416);
and U12763 (N_12763,N_12045,N_12305);
or U12764 (N_12764,N_12328,N_12552);
nor U12765 (N_12765,N_12504,N_12574);
or U12766 (N_12766,N_12096,N_12139);
and U12767 (N_12767,N_12496,N_12245);
and U12768 (N_12768,N_12301,N_12361);
or U12769 (N_12769,N_12252,N_12056);
xnor U12770 (N_12770,N_12346,N_12016);
and U12771 (N_12771,N_12184,N_12542);
nor U12772 (N_12772,N_12189,N_12487);
nand U12773 (N_12773,N_12255,N_12193);
xor U12774 (N_12774,N_12349,N_12468);
and U12775 (N_12775,N_12389,N_12447);
nand U12776 (N_12776,N_12218,N_12455);
nand U12777 (N_12777,N_12287,N_12033);
and U12778 (N_12778,N_12347,N_12465);
nor U12779 (N_12779,N_12501,N_12146);
and U12780 (N_12780,N_12340,N_12326);
nor U12781 (N_12781,N_12348,N_12026);
and U12782 (N_12782,N_12537,N_12111);
and U12783 (N_12783,N_12553,N_12345);
xor U12784 (N_12784,N_12094,N_12288);
and U12785 (N_12785,N_12423,N_12028);
and U12786 (N_12786,N_12341,N_12366);
and U12787 (N_12787,N_12306,N_12544);
and U12788 (N_12788,N_12543,N_12408);
nor U12789 (N_12789,N_12001,N_12437);
and U12790 (N_12790,N_12522,N_12116);
or U12791 (N_12791,N_12302,N_12002);
nor U12792 (N_12792,N_12159,N_12536);
nand U12793 (N_12793,N_12201,N_12597);
or U12794 (N_12794,N_12374,N_12469);
or U12795 (N_12795,N_12529,N_12568);
nand U12796 (N_12796,N_12358,N_12599);
and U12797 (N_12797,N_12352,N_12037);
nand U12798 (N_12798,N_12422,N_12088);
nand U12799 (N_12799,N_12093,N_12557);
nand U12800 (N_12800,N_12576,N_12556);
nand U12801 (N_12801,N_12113,N_12592);
nor U12802 (N_12802,N_12291,N_12074);
nor U12803 (N_12803,N_12048,N_12260);
and U12804 (N_12804,N_12025,N_12591);
and U12805 (N_12805,N_12514,N_12015);
and U12806 (N_12806,N_12402,N_12129);
nor U12807 (N_12807,N_12450,N_12134);
or U12808 (N_12808,N_12117,N_12164);
or U12809 (N_12809,N_12436,N_12563);
and U12810 (N_12810,N_12371,N_12538);
and U12811 (N_12811,N_12376,N_12342);
nand U12812 (N_12812,N_12081,N_12265);
and U12813 (N_12813,N_12167,N_12004);
or U12814 (N_12814,N_12581,N_12188);
nor U12815 (N_12815,N_12320,N_12205);
and U12816 (N_12816,N_12241,N_12238);
nor U12817 (N_12817,N_12387,N_12051);
nor U12818 (N_12818,N_12247,N_12428);
and U12819 (N_12819,N_12017,N_12069);
or U12820 (N_12820,N_12154,N_12380);
nor U12821 (N_12821,N_12209,N_12145);
or U12822 (N_12822,N_12583,N_12578);
and U12823 (N_12823,N_12024,N_12038);
nand U12824 (N_12824,N_12577,N_12192);
or U12825 (N_12825,N_12280,N_12087);
nand U12826 (N_12826,N_12331,N_12161);
and U12827 (N_12827,N_12430,N_12322);
nand U12828 (N_12828,N_12452,N_12315);
or U12829 (N_12829,N_12337,N_12227);
or U12830 (N_12830,N_12533,N_12303);
or U12831 (N_12831,N_12379,N_12177);
nor U12832 (N_12832,N_12186,N_12057);
nor U12833 (N_12833,N_12431,N_12052);
nor U12834 (N_12834,N_12183,N_12284);
xor U12835 (N_12835,N_12332,N_12080);
nor U12836 (N_12836,N_12283,N_12418);
and U12837 (N_12837,N_12275,N_12221);
nor U12838 (N_12838,N_12509,N_12135);
nand U12839 (N_12839,N_12481,N_12399);
nor U12840 (N_12840,N_12199,N_12106);
nand U12841 (N_12841,N_12256,N_12264);
nor U12842 (N_12842,N_12338,N_12579);
and U12843 (N_12843,N_12133,N_12123);
nor U12844 (N_12844,N_12505,N_12397);
nand U12845 (N_12845,N_12425,N_12246);
or U12846 (N_12846,N_12434,N_12309);
and U12847 (N_12847,N_12070,N_12032);
nand U12848 (N_12848,N_12359,N_12383);
nand U12849 (N_12849,N_12441,N_12029);
or U12850 (N_12850,N_12559,N_12414);
and U12851 (N_12851,N_12214,N_12373);
and U12852 (N_12852,N_12266,N_12083);
or U12853 (N_12853,N_12127,N_12190);
nor U12854 (N_12854,N_12329,N_12511);
or U12855 (N_12855,N_12130,N_12253);
nand U12856 (N_12856,N_12310,N_12018);
nand U12857 (N_12857,N_12150,N_12036);
or U12858 (N_12858,N_12439,N_12473);
or U12859 (N_12859,N_12060,N_12393);
and U12860 (N_12860,N_12059,N_12385);
and U12861 (N_12861,N_12215,N_12210);
and U12862 (N_12862,N_12313,N_12330);
and U12863 (N_12863,N_12333,N_12092);
nor U12864 (N_12864,N_12446,N_12098);
nand U12865 (N_12865,N_12151,N_12021);
nand U12866 (N_12866,N_12355,N_12185);
nand U12867 (N_12867,N_12286,N_12173);
or U12868 (N_12868,N_12198,N_12101);
nor U12869 (N_12869,N_12392,N_12240);
nor U12870 (N_12870,N_12176,N_12073);
or U12871 (N_12871,N_12334,N_12454);
nor U12872 (N_12872,N_12170,N_12336);
nand U12873 (N_12873,N_12325,N_12274);
or U12874 (N_12874,N_12404,N_12554);
nor U12875 (N_12875,N_12269,N_12203);
or U12876 (N_12876,N_12594,N_12572);
or U12877 (N_12877,N_12442,N_12311);
or U12878 (N_12878,N_12443,N_12382);
or U12879 (N_12879,N_12534,N_12014);
or U12880 (N_12880,N_12079,N_12171);
or U12881 (N_12881,N_12308,N_12050);
nor U12882 (N_12882,N_12561,N_12108);
nand U12883 (N_12883,N_12548,N_12593);
or U12884 (N_12884,N_12137,N_12066);
nor U12885 (N_12885,N_12044,N_12507);
or U12886 (N_12886,N_12412,N_12295);
and U12887 (N_12887,N_12035,N_12512);
nand U12888 (N_12888,N_12136,N_12307);
xor U12889 (N_12889,N_12089,N_12427);
xnor U12890 (N_12890,N_12122,N_12236);
xnor U12891 (N_12891,N_12525,N_12290);
and U12892 (N_12892,N_12107,N_12555);
or U12893 (N_12893,N_12386,N_12390);
and U12894 (N_12894,N_12474,N_12243);
nor U12895 (N_12895,N_12012,N_12558);
nand U12896 (N_12896,N_12158,N_12458);
or U12897 (N_12897,N_12567,N_12182);
xor U12898 (N_12898,N_12162,N_12077);
nor U12899 (N_12899,N_12316,N_12293);
or U12900 (N_12900,N_12542,N_12488);
xnor U12901 (N_12901,N_12572,N_12173);
nand U12902 (N_12902,N_12171,N_12230);
and U12903 (N_12903,N_12490,N_12588);
nand U12904 (N_12904,N_12008,N_12078);
and U12905 (N_12905,N_12083,N_12084);
nor U12906 (N_12906,N_12303,N_12420);
and U12907 (N_12907,N_12215,N_12453);
nor U12908 (N_12908,N_12127,N_12035);
nor U12909 (N_12909,N_12008,N_12268);
or U12910 (N_12910,N_12148,N_12413);
and U12911 (N_12911,N_12196,N_12122);
nor U12912 (N_12912,N_12523,N_12024);
or U12913 (N_12913,N_12153,N_12497);
nand U12914 (N_12914,N_12370,N_12167);
nand U12915 (N_12915,N_12596,N_12256);
nor U12916 (N_12916,N_12388,N_12217);
nand U12917 (N_12917,N_12243,N_12595);
nand U12918 (N_12918,N_12511,N_12062);
and U12919 (N_12919,N_12236,N_12120);
and U12920 (N_12920,N_12525,N_12232);
nand U12921 (N_12921,N_12216,N_12120);
nor U12922 (N_12922,N_12363,N_12284);
and U12923 (N_12923,N_12195,N_12112);
nand U12924 (N_12924,N_12413,N_12467);
and U12925 (N_12925,N_12294,N_12524);
and U12926 (N_12926,N_12229,N_12383);
xnor U12927 (N_12927,N_12515,N_12246);
nand U12928 (N_12928,N_12303,N_12253);
and U12929 (N_12929,N_12334,N_12426);
and U12930 (N_12930,N_12327,N_12529);
nand U12931 (N_12931,N_12524,N_12391);
and U12932 (N_12932,N_12236,N_12280);
and U12933 (N_12933,N_12178,N_12357);
xor U12934 (N_12934,N_12430,N_12502);
or U12935 (N_12935,N_12189,N_12356);
nand U12936 (N_12936,N_12506,N_12276);
or U12937 (N_12937,N_12558,N_12014);
nor U12938 (N_12938,N_12052,N_12189);
nor U12939 (N_12939,N_12103,N_12545);
nand U12940 (N_12940,N_12185,N_12505);
nor U12941 (N_12941,N_12283,N_12256);
nand U12942 (N_12942,N_12380,N_12296);
nor U12943 (N_12943,N_12403,N_12125);
nand U12944 (N_12944,N_12551,N_12128);
nor U12945 (N_12945,N_12178,N_12114);
nand U12946 (N_12946,N_12157,N_12599);
or U12947 (N_12947,N_12265,N_12210);
nor U12948 (N_12948,N_12590,N_12538);
xor U12949 (N_12949,N_12133,N_12599);
nor U12950 (N_12950,N_12214,N_12260);
nand U12951 (N_12951,N_12188,N_12289);
nor U12952 (N_12952,N_12283,N_12231);
nand U12953 (N_12953,N_12476,N_12430);
or U12954 (N_12954,N_12080,N_12382);
nor U12955 (N_12955,N_12521,N_12212);
nand U12956 (N_12956,N_12378,N_12270);
nand U12957 (N_12957,N_12068,N_12411);
xnor U12958 (N_12958,N_12415,N_12006);
nor U12959 (N_12959,N_12085,N_12137);
nor U12960 (N_12960,N_12234,N_12300);
nor U12961 (N_12961,N_12456,N_12503);
and U12962 (N_12962,N_12114,N_12155);
nor U12963 (N_12963,N_12199,N_12557);
xor U12964 (N_12964,N_12526,N_12357);
nand U12965 (N_12965,N_12233,N_12543);
or U12966 (N_12966,N_12001,N_12036);
nor U12967 (N_12967,N_12241,N_12542);
nor U12968 (N_12968,N_12194,N_12366);
and U12969 (N_12969,N_12047,N_12217);
and U12970 (N_12970,N_12046,N_12365);
nor U12971 (N_12971,N_12079,N_12414);
and U12972 (N_12972,N_12196,N_12299);
and U12973 (N_12973,N_12121,N_12187);
nor U12974 (N_12974,N_12254,N_12573);
nand U12975 (N_12975,N_12535,N_12378);
nand U12976 (N_12976,N_12225,N_12191);
and U12977 (N_12977,N_12487,N_12366);
or U12978 (N_12978,N_12564,N_12202);
nand U12979 (N_12979,N_12480,N_12594);
and U12980 (N_12980,N_12068,N_12537);
or U12981 (N_12981,N_12429,N_12386);
or U12982 (N_12982,N_12514,N_12302);
nor U12983 (N_12983,N_12133,N_12158);
and U12984 (N_12984,N_12354,N_12443);
nor U12985 (N_12985,N_12318,N_12562);
and U12986 (N_12986,N_12034,N_12539);
or U12987 (N_12987,N_12542,N_12231);
nor U12988 (N_12988,N_12440,N_12124);
nand U12989 (N_12989,N_12259,N_12297);
nor U12990 (N_12990,N_12204,N_12587);
or U12991 (N_12991,N_12413,N_12254);
nand U12992 (N_12992,N_12048,N_12474);
nand U12993 (N_12993,N_12150,N_12160);
or U12994 (N_12994,N_12284,N_12409);
xor U12995 (N_12995,N_12343,N_12288);
and U12996 (N_12996,N_12128,N_12505);
and U12997 (N_12997,N_12469,N_12398);
and U12998 (N_12998,N_12144,N_12028);
nor U12999 (N_12999,N_12347,N_12413);
or U13000 (N_13000,N_12437,N_12591);
nor U13001 (N_13001,N_12246,N_12014);
and U13002 (N_13002,N_12141,N_12169);
or U13003 (N_13003,N_12069,N_12578);
or U13004 (N_13004,N_12596,N_12311);
or U13005 (N_13005,N_12599,N_12004);
and U13006 (N_13006,N_12186,N_12411);
nand U13007 (N_13007,N_12098,N_12485);
nor U13008 (N_13008,N_12105,N_12078);
nand U13009 (N_13009,N_12055,N_12215);
nor U13010 (N_13010,N_12292,N_12163);
nor U13011 (N_13011,N_12570,N_12493);
nor U13012 (N_13012,N_12113,N_12089);
or U13013 (N_13013,N_12395,N_12187);
nand U13014 (N_13014,N_12379,N_12345);
nor U13015 (N_13015,N_12585,N_12077);
or U13016 (N_13016,N_12010,N_12245);
nand U13017 (N_13017,N_12101,N_12230);
and U13018 (N_13018,N_12479,N_12521);
nand U13019 (N_13019,N_12182,N_12443);
or U13020 (N_13020,N_12073,N_12386);
and U13021 (N_13021,N_12153,N_12307);
nor U13022 (N_13022,N_12002,N_12297);
and U13023 (N_13023,N_12212,N_12451);
or U13024 (N_13024,N_12135,N_12442);
nand U13025 (N_13025,N_12167,N_12500);
or U13026 (N_13026,N_12108,N_12456);
nor U13027 (N_13027,N_12507,N_12126);
nand U13028 (N_13028,N_12290,N_12198);
or U13029 (N_13029,N_12537,N_12289);
nor U13030 (N_13030,N_12042,N_12027);
and U13031 (N_13031,N_12236,N_12115);
or U13032 (N_13032,N_12405,N_12531);
and U13033 (N_13033,N_12179,N_12481);
and U13034 (N_13034,N_12395,N_12558);
or U13035 (N_13035,N_12131,N_12304);
xor U13036 (N_13036,N_12245,N_12286);
or U13037 (N_13037,N_12511,N_12239);
or U13038 (N_13038,N_12560,N_12580);
nand U13039 (N_13039,N_12565,N_12091);
or U13040 (N_13040,N_12489,N_12075);
or U13041 (N_13041,N_12296,N_12053);
nor U13042 (N_13042,N_12101,N_12470);
nor U13043 (N_13043,N_12129,N_12364);
nor U13044 (N_13044,N_12588,N_12054);
or U13045 (N_13045,N_12555,N_12007);
nor U13046 (N_13046,N_12251,N_12394);
and U13047 (N_13047,N_12014,N_12474);
or U13048 (N_13048,N_12241,N_12219);
or U13049 (N_13049,N_12554,N_12424);
nor U13050 (N_13050,N_12263,N_12558);
nor U13051 (N_13051,N_12202,N_12507);
nand U13052 (N_13052,N_12067,N_12413);
or U13053 (N_13053,N_12526,N_12459);
or U13054 (N_13054,N_12378,N_12175);
nand U13055 (N_13055,N_12379,N_12499);
and U13056 (N_13056,N_12057,N_12016);
nand U13057 (N_13057,N_12505,N_12018);
and U13058 (N_13058,N_12372,N_12214);
or U13059 (N_13059,N_12175,N_12388);
and U13060 (N_13060,N_12331,N_12259);
or U13061 (N_13061,N_12563,N_12463);
or U13062 (N_13062,N_12159,N_12093);
and U13063 (N_13063,N_12214,N_12049);
or U13064 (N_13064,N_12136,N_12435);
nor U13065 (N_13065,N_12135,N_12431);
nor U13066 (N_13066,N_12200,N_12333);
or U13067 (N_13067,N_12439,N_12425);
or U13068 (N_13068,N_12327,N_12045);
nor U13069 (N_13069,N_12244,N_12083);
or U13070 (N_13070,N_12339,N_12559);
or U13071 (N_13071,N_12171,N_12347);
or U13072 (N_13072,N_12136,N_12161);
nor U13073 (N_13073,N_12178,N_12014);
and U13074 (N_13074,N_12303,N_12296);
or U13075 (N_13075,N_12565,N_12536);
nor U13076 (N_13076,N_12217,N_12300);
and U13077 (N_13077,N_12267,N_12053);
nand U13078 (N_13078,N_12219,N_12108);
or U13079 (N_13079,N_12175,N_12529);
nand U13080 (N_13080,N_12553,N_12141);
or U13081 (N_13081,N_12538,N_12030);
and U13082 (N_13082,N_12564,N_12177);
nor U13083 (N_13083,N_12505,N_12319);
or U13084 (N_13084,N_12331,N_12083);
nor U13085 (N_13085,N_12248,N_12451);
or U13086 (N_13086,N_12090,N_12099);
and U13087 (N_13087,N_12469,N_12121);
nand U13088 (N_13088,N_12460,N_12524);
and U13089 (N_13089,N_12070,N_12290);
nor U13090 (N_13090,N_12356,N_12543);
or U13091 (N_13091,N_12577,N_12144);
nor U13092 (N_13092,N_12475,N_12533);
and U13093 (N_13093,N_12077,N_12446);
nor U13094 (N_13094,N_12247,N_12507);
and U13095 (N_13095,N_12173,N_12568);
or U13096 (N_13096,N_12455,N_12277);
nor U13097 (N_13097,N_12155,N_12531);
nand U13098 (N_13098,N_12080,N_12419);
nand U13099 (N_13099,N_12483,N_12547);
and U13100 (N_13100,N_12021,N_12249);
or U13101 (N_13101,N_12544,N_12426);
or U13102 (N_13102,N_12044,N_12225);
nand U13103 (N_13103,N_12020,N_12167);
nor U13104 (N_13104,N_12030,N_12402);
nor U13105 (N_13105,N_12030,N_12233);
nor U13106 (N_13106,N_12156,N_12227);
or U13107 (N_13107,N_12496,N_12019);
nand U13108 (N_13108,N_12181,N_12466);
nand U13109 (N_13109,N_12509,N_12544);
or U13110 (N_13110,N_12125,N_12158);
nor U13111 (N_13111,N_12126,N_12449);
nand U13112 (N_13112,N_12493,N_12555);
nor U13113 (N_13113,N_12324,N_12074);
or U13114 (N_13114,N_12142,N_12228);
or U13115 (N_13115,N_12502,N_12223);
or U13116 (N_13116,N_12404,N_12443);
nor U13117 (N_13117,N_12174,N_12586);
or U13118 (N_13118,N_12493,N_12159);
nand U13119 (N_13119,N_12250,N_12199);
and U13120 (N_13120,N_12432,N_12399);
and U13121 (N_13121,N_12417,N_12484);
or U13122 (N_13122,N_12467,N_12054);
and U13123 (N_13123,N_12358,N_12284);
nand U13124 (N_13124,N_12245,N_12506);
nand U13125 (N_13125,N_12439,N_12125);
and U13126 (N_13126,N_12126,N_12249);
and U13127 (N_13127,N_12518,N_12428);
or U13128 (N_13128,N_12317,N_12172);
nor U13129 (N_13129,N_12104,N_12135);
nand U13130 (N_13130,N_12318,N_12458);
nor U13131 (N_13131,N_12069,N_12422);
nand U13132 (N_13132,N_12272,N_12359);
and U13133 (N_13133,N_12091,N_12577);
nand U13134 (N_13134,N_12198,N_12138);
or U13135 (N_13135,N_12273,N_12592);
and U13136 (N_13136,N_12081,N_12125);
and U13137 (N_13137,N_12377,N_12067);
nand U13138 (N_13138,N_12216,N_12579);
nand U13139 (N_13139,N_12034,N_12196);
or U13140 (N_13140,N_12447,N_12255);
or U13141 (N_13141,N_12421,N_12080);
and U13142 (N_13142,N_12400,N_12461);
or U13143 (N_13143,N_12126,N_12166);
or U13144 (N_13144,N_12478,N_12281);
nand U13145 (N_13145,N_12276,N_12126);
nand U13146 (N_13146,N_12304,N_12054);
nand U13147 (N_13147,N_12267,N_12363);
nor U13148 (N_13148,N_12440,N_12009);
nor U13149 (N_13149,N_12526,N_12015);
and U13150 (N_13150,N_12034,N_12094);
nor U13151 (N_13151,N_12576,N_12524);
or U13152 (N_13152,N_12282,N_12464);
or U13153 (N_13153,N_12496,N_12294);
nor U13154 (N_13154,N_12196,N_12256);
nand U13155 (N_13155,N_12259,N_12531);
nand U13156 (N_13156,N_12517,N_12218);
nor U13157 (N_13157,N_12029,N_12457);
nand U13158 (N_13158,N_12438,N_12205);
and U13159 (N_13159,N_12334,N_12586);
xor U13160 (N_13160,N_12209,N_12520);
or U13161 (N_13161,N_12264,N_12207);
or U13162 (N_13162,N_12061,N_12354);
nand U13163 (N_13163,N_12543,N_12542);
nand U13164 (N_13164,N_12544,N_12226);
xor U13165 (N_13165,N_12246,N_12417);
nor U13166 (N_13166,N_12596,N_12355);
or U13167 (N_13167,N_12018,N_12191);
nand U13168 (N_13168,N_12276,N_12267);
or U13169 (N_13169,N_12141,N_12183);
or U13170 (N_13170,N_12213,N_12417);
xor U13171 (N_13171,N_12029,N_12380);
or U13172 (N_13172,N_12138,N_12064);
or U13173 (N_13173,N_12348,N_12258);
nor U13174 (N_13174,N_12324,N_12188);
or U13175 (N_13175,N_12497,N_12108);
and U13176 (N_13176,N_12281,N_12155);
nor U13177 (N_13177,N_12569,N_12400);
nor U13178 (N_13178,N_12197,N_12466);
and U13179 (N_13179,N_12052,N_12051);
or U13180 (N_13180,N_12185,N_12217);
nor U13181 (N_13181,N_12470,N_12369);
xnor U13182 (N_13182,N_12227,N_12165);
and U13183 (N_13183,N_12511,N_12460);
nand U13184 (N_13184,N_12336,N_12412);
nand U13185 (N_13185,N_12420,N_12145);
nand U13186 (N_13186,N_12086,N_12015);
nand U13187 (N_13187,N_12407,N_12366);
nand U13188 (N_13188,N_12257,N_12180);
and U13189 (N_13189,N_12244,N_12424);
nor U13190 (N_13190,N_12128,N_12106);
nand U13191 (N_13191,N_12019,N_12150);
nor U13192 (N_13192,N_12478,N_12072);
or U13193 (N_13193,N_12158,N_12297);
nor U13194 (N_13194,N_12027,N_12429);
nand U13195 (N_13195,N_12184,N_12566);
or U13196 (N_13196,N_12022,N_12528);
nand U13197 (N_13197,N_12321,N_12090);
and U13198 (N_13198,N_12456,N_12508);
or U13199 (N_13199,N_12016,N_12460);
nand U13200 (N_13200,N_12996,N_13139);
and U13201 (N_13201,N_12867,N_13029);
nand U13202 (N_13202,N_13134,N_12997);
and U13203 (N_13203,N_12721,N_12913);
or U13204 (N_13204,N_12677,N_12839);
and U13205 (N_13205,N_12736,N_13001);
or U13206 (N_13206,N_13176,N_12968);
nor U13207 (N_13207,N_12609,N_13118);
nand U13208 (N_13208,N_12704,N_13083);
nand U13209 (N_13209,N_12714,N_13132);
nand U13210 (N_13210,N_13079,N_13062);
or U13211 (N_13211,N_12754,N_12779);
nand U13212 (N_13212,N_12826,N_12735);
nor U13213 (N_13213,N_12883,N_13126);
and U13214 (N_13214,N_12957,N_13099);
and U13215 (N_13215,N_12795,N_13145);
nor U13216 (N_13216,N_12875,N_13193);
nand U13217 (N_13217,N_13188,N_13190);
nor U13218 (N_13218,N_12855,N_12756);
nand U13219 (N_13219,N_12682,N_12724);
or U13220 (N_13220,N_13178,N_12964);
or U13221 (N_13221,N_12917,N_12882);
and U13222 (N_13222,N_12653,N_12678);
nand U13223 (N_13223,N_12841,N_12743);
or U13224 (N_13224,N_12765,N_13045);
and U13225 (N_13225,N_13010,N_13124);
or U13226 (N_13226,N_12711,N_12665);
nor U13227 (N_13227,N_12651,N_12930);
nand U13228 (N_13228,N_12628,N_12999);
and U13229 (N_13229,N_13056,N_13112);
nand U13230 (N_13230,N_12733,N_13011);
or U13231 (N_13231,N_13129,N_12695);
nand U13232 (N_13232,N_12837,N_12858);
or U13233 (N_13233,N_13180,N_13050);
nor U13234 (N_13234,N_13031,N_13000);
or U13235 (N_13235,N_12831,N_13059);
xnor U13236 (N_13236,N_12949,N_12904);
or U13237 (N_13237,N_13194,N_13092);
and U13238 (N_13238,N_12786,N_12862);
and U13239 (N_13239,N_13035,N_13192);
or U13240 (N_13240,N_13021,N_13068);
and U13241 (N_13241,N_13130,N_13199);
or U13242 (N_13242,N_13156,N_13012);
nor U13243 (N_13243,N_12873,N_13164);
or U13244 (N_13244,N_12702,N_12832);
xnor U13245 (N_13245,N_12891,N_13127);
nor U13246 (N_13246,N_12921,N_12749);
nand U13247 (N_13247,N_12829,N_13122);
nor U13248 (N_13248,N_13002,N_12920);
or U13249 (N_13249,N_12800,N_13087);
and U13250 (N_13250,N_12849,N_12960);
xor U13251 (N_13251,N_12819,N_13168);
and U13252 (N_13252,N_13096,N_12720);
nor U13253 (N_13253,N_13057,N_13090);
or U13254 (N_13254,N_12990,N_13166);
or U13255 (N_13255,N_13151,N_13114);
nor U13256 (N_13256,N_12636,N_13007);
nand U13257 (N_13257,N_12851,N_12911);
nand U13258 (N_13258,N_13133,N_12899);
nor U13259 (N_13259,N_12692,N_12923);
nor U13260 (N_13260,N_12966,N_12722);
and U13261 (N_13261,N_13154,N_12901);
nand U13262 (N_13262,N_12944,N_12965);
or U13263 (N_13263,N_12885,N_12633);
nor U13264 (N_13264,N_12974,N_12778);
or U13265 (N_13265,N_12980,N_13028);
or U13266 (N_13266,N_12767,N_13069);
and U13267 (N_13267,N_12621,N_12947);
nand U13268 (N_13268,N_12739,N_12657);
or U13269 (N_13269,N_12670,N_13044);
xnor U13270 (N_13270,N_13063,N_12798);
and U13271 (N_13271,N_12614,N_13033);
nand U13272 (N_13272,N_13171,N_12672);
and U13273 (N_13273,N_12925,N_12744);
and U13274 (N_13274,N_12706,N_13058);
nor U13275 (N_13275,N_12856,N_12707);
nor U13276 (N_13276,N_13146,N_12846);
or U13277 (N_13277,N_12802,N_12690);
or U13278 (N_13278,N_13017,N_13136);
nand U13279 (N_13279,N_12908,N_12649);
or U13280 (N_13280,N_12812,N_12822);
nand U13281 (N_13281,N_12834,N_13172);
and U13282 (N_13282,N_12955,N_12658);
nor U13283 (N_13283,N_12729,N_12763);
or U13284 (N_13284,N_12630,N_12638);
nor U13285 (N_13285,N_12945,N_12626);
nor U13286 (N_13286,N_12660,N_12809);
nor U13287 (N_13287,N_13117,N_12619);
nor U13288 (N_13288,N_12853,N_12751);
nand U13289 (N_13289,N_12631,N_13177);
or U13290 (N_13290,N_12728,N_12994);
nand U13291 (N_13291,N_12680,N_13187);
or U13292 (N_13292,N_13159,N_12813);
or U13293 (N_13293,N_12953,N_13179);
or U13294 (N_13294,N_13170,N_13003);
and U13295 (N_13295,N_12664,N_13073);
xnor U13296 (N_13296,N_12725,N_12848);
or U13297 (N_13297,N_12652,N_13064);
nor U13298 (N_13298,N_12869,N_12732);
nor U13299 (N_13299,N_13191,N_12622);
nor U13300 (N_13300,N_12662,N_12854);
nand U13301 (N_13301,N_12956,N_12629);
and U13302 (N_13302,N_13152,N_13088);
nor U13303 (N_13303,N_12892,N_12773);
and U13304 (N_13304,N_12713,N_13004);
nand U13305 (N_13305,N_13006,N_13026);
xnor U13306 (N_13306,N_12742,N_12723);
nor U13307 (N_13307,N_13037,N_12691);
nand U13308 (N_13308,N_12700,N_12808);
xor U13309 (N_13309,N_12864,N_12650);
nand U13310 (N_13310,N_12865,N_12632);
nor U13311 (N_13311,N_12878,N_12993);
or U13312 (N_13312,N_12698,N_12654);
nand U13313 (N_13313,N_12717,N_13076);
nor U13314 (N_13314,N_12909,N_12746);
and U13315 (N_13315,N_13169,N_13052);
nand U13316 (N_13316,N_13105,N_12696);
and U13317 (N_13317,N_12967,N_13153);
nor U13318 (N_13318,N_12676,N_13110);
and U13319 (N_13319,N_13030,N_13144);
nor U13320 (N_13320,N_12675,N_12606);
nand U13321 (N_13321,N_13077,N_12718);
or U13322 (N_13322,N_12868,N_12794);
or U13323 (N_13323,N_13121,N_13027);
or U13324 (N_13324,N_12973,N_12852);
nor U13325 (N_13325,N_12770,N_12982);
or U13326 (N_13326,N_12975,N_13198);
nor U13327 (N_13327,N_12612,N_12948);
and U13328 (N_13328,N_12979,N_13125);
or U13329 (N_13329,N_13113,N_12991);
nor U13330 (N_13330,N_13183,N_12915);
nor U13331 (N_13331,N_12668,N_13115);
or U13332 (N_13332,N_12874,N_12978);
nand U13333 (N_13333,N_12792,N_12821);
and U13334 (N_13334,N_13085,N_12893);
or U13335 (N_13335,N_12719,N_13135);
nand U13336 (N_13336,N_13023,N_12656);
or U13337 (N_13337,N_12823,N_12842);
nor U13338 (N_13338,N_12916,N_12799);
nand U13339 (N_13339,N_12835,N_12818);
nand U13340 (N_13340,N_13071,N_12634);
and U13341 (N_13341,N_13070,N_12946);
or U13342 (N_13342,N_12937,N_12914);
nand U13343 (N_13343,N_12666,N_12881);
and U13344 (N_13344,N_12860,N_12667);
nand U13345 (N_13345,N_13078,N_12608);
nor U13346 (N_13346,N_13014,N_13024);
or U13347 (N_13347,N_13015,N_12663);
and U13348 (N_13348,N_12686,N_12764);
nand U13349 (N_13349,N_13082,N_12811);
nor U13350 (N_13350,N_13100,N_13197);
and U13351 (N_13351,N_13039,N_12694);
nand U13352 (N_13352,N_13175,N_12603);
nor U13353 (N_13353,N_12640,N_12963);
nor U13354 (N_13354,N_12731,N_12709);
nand U13355 (N_13355,N_13111,N_12827);
nand U13356 (N_13356,N_12726,N_12984);
nor U13357 (N_13357,N_12986,N_12772);
xor U13358 (N_13358,N_13061,N_12992);
nor U13359 (N_13359,N_12624,N_12645);
or U13360 (N_13360,N_13161,N_13138);
or U13361 (N_13361,N_12872,N_12816);
and U13362 (N_13362,N_12679,N_12616);
nand U13363 (N_13363,N_12783,N_13089);
nand U13364 (N_13364,N_12897,N_12604);
and U13365 (N_13365,N_12693,N_13141);
and U13366 (N_13366,N_12820,N_13009);
and U13367 (N_13367,N_13109,N_12791);
or U13368 (N_13368,N_12617,N_13137);
or U13369 (N_13369,N_12906,N_12647);
or U13370 (N_13370,N_12871,N_13038);
nand U13371 (N_13371,N_12922,N_13140);
or U13372 (N_13372,N_13086,N_13098);
nand U13373 (N_13373,N_12951,N_12902);
nor U13374 (N_13374,N_13107,N_13067);
xnor U13375 (N_13375,N_13036,N_12927);
nand U13376 (N_13376,N_12699,N_12924);
nand U13377 (N_13377,N_12903,N_12785);
nand U13378 (N_13378,N_12788,N_13055);
or U13379 (N_13379,N_13163,N_13160);
nor U13380 (N_13380,N_12635,N_12907);
nor U13381 (N_13381,N_13155,N_13147);
and U13382 (N_13382,N_12689,N_12790);
nor U13383 (N_13383,N_13041,N_13157);
nor U13384 (N_13384,N_12807,N_13025);
nor U13385 (N_13385,N_12988,N_13074);
and U13386 (N_13386,N_13196,N_12870);
nor U13387 (N_13387,N_12970,N_13149);
and U13388 (N_13388,N_12697,N_12659);
nand U13389 (N_13389,N_12936,N_12737);
or U13390 (N_13390,N_12952,N_12701);
nand U13391 (N_13391,N_13123,N_12727);
or U13392 (N_13392,N_13120,N_12833);
and U13393 (N_13393,N_12752,N_13150);
and U13394 (N_13394,N_12781,N_13143);
nor U13395 (N_13395,N_12895,N_13013);
nor U13396 (N_13396,N_12712,N_12888);
and U13397 (N_13397,N_13018,N_13048);
nand U13398 (N_13398,N_12750,N_12912);
nor U13399 (N_13399,N_12615,N_12815);
nand U13400 (N_13400,N_12942,N_12933);
nand U13401 (N_13401,N_13060,N_12646);
or U13402 (N_13402,N_12977,N_12806);
and U13403 (N_13403,N_13148,N_12859);
nor U13404 (N_13404,N_13075,N_12740);
nand U13405 (N_13405,N_12681,N_12757);
nor U13406 (N_13406,N_12863,N_12618);
nor U13407 (N_13407,N_13020,N_12669);
or U13408 (N_13408,N_12890,N_13049);
nor U13409 (N_13409,N_13174,N_12610);
or U13410 (N_13410,N_12685,N_12989);
and U13411 (N_13411,N_12661,N_12880);
nand U13412 (N_13412,N_12810,N_12828);
nor U13413 (N_13413,N_12745,N_12793);
and U13414 (N_13414,N_12887,N_12777);
and U13415 (N_13415,N_12708,N_12918);
and U13416 (N_13416,N_12998,N_12961);
nand U13417 (N_13417,N_12959,N_12969);
and U13418 (N_13418,N_12929,N_13065);
or U13419 (N_13419,N_12730,N_12847);
nand U13420 (N_13420,N_12748,N_13116);
and U13421 (N_13421,N_13158,N_12814);
or U13422 (N_13422,N_13189,N_12771);
or U13423 (N_13423,N_12639,N_13032);
or U13424 (N_13424,N_12776,N_12759);
and U13425 (N_13425,N_13042,N_12983);
nor U13426 (N_13426,N_13022,N_12910);
or U13427 (N_13427,N_12716,N_12843);
or U13428 (N_13428,N_12671,N_12840);
nor U13429 (N_13429,N_12919,N_12766);
and U13430 (N_13430,N_12705,N_12905);
nand U13431 (N_13431,N_12782,N_12688);
nor U13432 (N_13432,N_12643,N_12644);
nor U13433 (N_13433,N_12876,N_13103);
and U13434 (N_13434,N_12932,N_12796);
nand U13435 (N_13435,N_13094,N_12939);
or U13436 (N_13436,N_13054,N_12894);
nor U13437 (N_13437,N_13016,N_13091);
xnor U13438 (N_13438,N_13008,N_12747);
and U13439 (N_13439,N_12801,N_12935);
nor U13440 (N_13440,N_13072,N_12673);
nor U13441 (N_13441,N_12940,N_12769);
nor U13442 (N_13442,N_12981,N_12602);
or U13443 (N_13443,N_12805,N_13173);
and U13444 (N_13444,N_12753,N_13181);
or U13445 (N_13445,N_12607,N_12755);
nor U13446 (N_13446,N_12987,N_12687);
and U13447 (N_13447,N_12803,N_12710);
or U13448 (N_13448,N_12641,N_12784);
or U13449 (N_13449,N_12683,N_12972);
nor U13450 (N_13450,N_13104,N_13162);
and U13451 (N_13451,N_12738,N_12601);
and U13452 (N_13452,N_13081,N_13142);
nor U13453 (N_13453,N_13051,N_12938);
and U13454 (N_13454,N_12958,N_12886);
nand U13455 (N_13455,N_12941,N_12758);
nor U13456 (N_13456,N_13097,N_12625);
xor U13457 (N_13457,N_12866,N_12787);
nor U13458 (N_13458,N_12824,N_12762);
or U13459 (N_13459,N_13066,N_12962);
or U13460 (N_13460,N_12844,N_12703);
nor U13461 (N_13461,N_13182,N_12825);
and U13462 (N_13462,N_13184,N_12934);
nor U13463 (N_13463,N_12775,N_13165);
nand U13464 (N_13464,N_12954,N_12741);
nor U13465 (N_13465,N_13053,N_13043);
nor U13466 (N_13466,N_12613,N_12928);
nand U13467 (N_13467,N_12734,N_12611);
nor U13468 (N_13468,N_12877,N_12768);
nand U13469 (N_13469,N_13101,N_12623);
nor U13470 (N_13470,N_12637,N_12889);
nor U13471 (N_13471,N_13108,N_12884);
xnor U13472 (N_13472,N_12830,N_12896);
and U13473 (N_13473,N_13131,N_12780);
or U13474 (N_13474,N_13102,N_12898);
and U13475 (N_13475,N_13128,N_13186);
nor U13476 (N_13476,N_12620,N_12861);
xor U13477 (N_13477,N_12850,N_13119);
nor U13478 (N_13478,N_13167,N_13005);
or U13479 (N_13479,N_12838,N_12857);
nor U13480 (N_13480,N_13093,N_12605);
nand U13481 (N_13481,N_12715,N_12797);
and U13482 (N_13482,N_12600,N_12789);
nand U13483 (N_13483,N_12976,N_12648);
or U13484 (N_13484,N_13034,N_12804);
and U13485 (N_13485,N_13046,N_12985);
or U13486 (N_13486,N_12684,N_13040);
nor U13487 (N_13487,N_12943,N_12674);
and U13488 (N_13488,N_13047,N_12950);
nor U13489 (N_13489,N_12642,N_12879);
or U13490 (N_13490,N_12627,N_13106);
or U13491 (N_13491,N_13080,N_12931);
nor U13492 (N_13492,N_12971,N_12760);
nand U13493 (N_13493,N_12926,N_13095);
and U13494 (N_13494,N_13195,N_12774);
or U13495 (N_13495,N_12761,N_13084);
or U13496 (N_13496,N_12817,N_13019);
nor U13497 (N_13497,N_12900,N_13185);
nand U13498 (N_13498,N_12995,N_12655);
nand U13499 (N_13499,N_12836,N_12845);
or U13500 (N_13500,N_12762,N_12955);
or U13501 (N_13501,N_12626,N_12882);
nor U13502 (N_13502,N_13051,N_12939);
nand U13503 (N_13503,N_12654,N_12755);
nor U13504 (N_13504,N_13102,N_13013);
or U13505 (N_13505,N_12855,N_13045);
nand U13506 (N_13506,N_13139,N_12613);
or U13507 (N_13507,N_12919,N_12715);
or U13508 (N_13508,N_12710,N_12891);
nand U13509 (N_13509,N_13155,N_12998);
nand U13510 (N_13510,N_12958,N_12681);
and U13511 (N_13511,N_12690,N_12951);
and U13512 (N_13512,N_12670,N_12956);
and U13513 (N_13513,N_12946,N_13103);
nor U13514 (N_13514,N_12916,N_12977);
or U13515 (N_13515,N_12713,N_13014);
or U13516 (N_13516,N_12638,N_13162);
or U13517 (N_13517,N_12609,N_12981);
or U13518 (N_13518,N_12614,N_12718);
nor U13519 (N_13519,N_12717,N_13135);
and U13520 (N_13520,N_12655,N_12801);
nor U13521 (N_13521,N_13023,N_12686);
or U13522 (N_13522,N_12750,N_13048);
and U13523 (N_13523,N_12893,N_12767);
or U13524 (N_13524,N_13128,N_13190);
or U13525 (N_13525,N_12877,N_13096);
xor U13526 (N_13526,N_12780,N_13176);
and U13527 (N_13527,N_13076,N_12826);
and U13528 (N_13528,N_12669,N_12827);
nor U13529 (N_13529,N_13043,N_13154);
nand U13530 (N_13530,N_12895,N_12630);
or U13531 (N_13531,N_12677,N_12712);
nor U13532 (N_13532,N_13057,N_12683);
or U13533 (N_13533,N_12838,N_12734);
nor U13534 (N_13534,N_12820,N_12905);
or U13535 (N_13535,N_13047,N_12988);
nand U13536 (N_13536,N_12652,N_13091);
and U13537 (N_13537,N_12817,N_13104);
and U13538 (N_13538,N_12650,N_12617);
nand U13539 (N_13539,N_12691,N_12882);
and U13540 (N_13540,N_12885,N_13007);
nor U13541 (N_13541,N_12771,N_12726);
nand U13542 (N_13542,N_12677,N_12899);
or U13543 (N_13543,N_12785,N_12768);
or U13544 (N_13544,N_12937,N_12918);
nand U13545 (N_13545,N_12886,N_13157);
nor U13546 (N_13546,N_13034,N_13010);
or U13547 (N_13547,N_12924,N_12830);
and U13548 (N_13548,N_12765,N_12655);
or U13549 (N_13549,N_12728,N_12646);
nor U13550 (N_13550,N_12988,N_13096);
xor U13551 (N_13551,N_13067,N_13096);
or U13552 (N_13552,N_12932,N_12665);
and U13553 (N_13553,N_12921,N_13128);
or U13554 (N_13554,N_12693,N_13095);
nor U13555 (N_13555,N_13088,N_12928);
xnor U13556 (N_13556,N_12866,N_12691);
nand U13557 (N_13557,N_13195,N_12675);
or U13558 (N_13558,N_13155,N_12831);
nor U13559 (N_13559,N_12742,N_13117);
or U13560 (N_13560,N_12726,N_12911);
or U13561 (N_13561,N_12789,N_12605);
or U13562 (N_13562,N_13182,N_12915);
and U13563 (N_13563,N_13099,N_12659);
nand U13564 (N_13564,N_12831,N_12955);
nand U13565 (N_13565,N_12682,N_13036);
nand U13566 (N_13566,N_12821,N_12822);
and U13567 (N_13567,N_12761,N_13108);
and U13568 (N_13568,N_13073,N_13119);
or U13569 (N_13569,N_12633,N_12848);
and U13570 (N_13570,N_12943,N_12878);
nor U13571 (N_13571,N_12769,N_12904);
nor U13572 (N_13572,N_13132,N_12777);
nor U13573 (N_13573,N_12781,N_13000);
or U13574 (N_13574,N_12632,N_13144);
nand U13575 (N_13575,N_12629,N_12977);
nor U13576 (N_13576,N_12699,N_12883);
and U13577 (N_13577,N_12692,N_13156);
nand U13578 (N_13578,N_12906,N_12811);
and U13579 (N_13579,N_13183,N_12814);
or U13580 (N_13580,N_12727,N_13186);
or U13581 (N_13581,N_12692,N_12717);
nor U13582 (N_13582,N_12905,N_12811);
and U13583 (N_13583,N_12893,N_13069);
nor U13584 (N_13584,N_12611,N_12607);
nor U13585 (N_13585,N_13134,N_12823);
or U13586 (N_13586,N_12757,N_13160);
xor U13587 (N_13587,N_12848,N_12884);
or U13588 (N_13588,N_13034,N_13046);
and U13589 (N_13589,N_12960,N_13154);
nor U13590 (N_13590,N_12902,N_12883);
xor U13591 (N_13591,N_13021,N_12708);
nand U13592 (N_13592,N_12751,N_12811);
nand U13593 (N_13593,N_13011,N_12616);
nor U13594 (N_13594,N_12835,N_13196);
nor U13595 (N_13595,N_13089,N_13057);
or U13596 (N_13596,N_12688,N_12989);
nand U13597 (N_13597,N_12680,N_13016);
and U13598 (N_13598,N_13180,N_12789);
nand U13599 (N_13599,N_12956,N_12971);
or U13600 (N_13600,N_13108,N_12737);
nand U13601 (N_13601,N_13039,N_12763);
and U13602 (N_13602,N_12635,N_12605);
nand U13603 (N_13603,N_12887,N_12812);
and U13604 (N_13604,N_12678,N_12715);
and U13605 (N_13605,N_12631,N_13164);
and U13606 (N_13606,N_13032,N_12740);
nand U13607 (N_13607,N_12926,N_13067);
xnor U13608 (N_13608,N_12769,N_12944);
nand U13609 (N_13609,N_12794,N_13117);
nand U13610 (N_13610,N_13067,N_12765);
nor U13611 (N_13611,N_13016,N_12880);
nand U13612 (N_13612,N_12619,N_13141);
nor U13613 (N_13613,N_12938,N_12612);
nand U13614 (N_13614,N_12788,N_12713);
nor U13615 (N_13615,N_13027,N_12706);
and U13616 (N_13616,N_12820,N_13119);
nor U13617 (N_13617,N_12628,N_12768);
nand U13618 (N_13618,N_12875,N_12971);
nor U13619 (N_13619,N_13193,N_13110);
nor U13620 (N_13620,N_13130,N_12649);
nand U13621 (N_13621,N_13184,N_13029);
nor U13622 (N_13622,N_12964,N_12617);
or U13623 (N_13623,N_13014,N_12780);
nand U13624 (N_13624,N_12819,N_13173);
nand U13625 (N_13625,N_12786,N_12710);
nand U13626 (N_13626,N_13043,N_12613);
and U13627 (N_13627,N_12635,N_13120);
or U13628 (N_13628,N_12684,N_12836);
and U13629 (N_13629,N_12696,N_12713);
and U13630 (N_13630,N_12743,N_13167);
or U13631 (N_13631,N_12914,N_13150);
and U13632 (N_13632,N_12872,N_12807);
or U13633 (N_13633,N_12681,N_12977);
nor U13634 (N_13634,N_12995,N_13050);
nor U13635 (N_13635,N_12687,N_12902);
nor U13636 (N_13636,N_12967,N_13076);
and U13637 (N_13637,N_12705,N_12866);
nand U13638 (N_13638,N_13146,N_12884);
nor U13639 (N_13639,N_12913,N_12613);
nor U13640 (N_13640,N_12696,N_12886);
and U13641 (N_13641,N_12862,N_13142);
nand U13642 (N_13642,N_12835,N_12868);
or U13643 (N_13643,N_12958,N_12649);
nor U13644 (N_13644,N_12804,N_12996);
and U13645 (N_13645,N_12600,N_12856);
and U13646 (N_13646,N_12765,N_12701);
and U13647 (N_13647,N_13060,N_12864);
nand U13648 (N_13648,N_13025,N_13139);
and U13649 (N_13649,N_13073,N_12738);
or U13650 (N_13650,N_12777,N_13063);
nand U13651 (N_13651,N_12970,N_13019);
nor U13652 (N_13652,N_12984,N_12686);
and U13653 (N_13653,N_12731,N_12739);
and U13654 (N_13654,N_12966,N_13154);
and U13655 (N_13655,N_13160,N_12884);
nand U13656 (N_13656,N_13075,N_12621);
nand U13657 (N_13657,N_13015,N_13117);
nor U13658 (N_13658,N_12625,N_13066);
xnor U13659 (N_13659,N_12963,N_13196);
or U13660 (N_13660,N_12940,N_12719);
nor U13661 (N_13661,N_12618,N_12675);
nand U13662 (N_13662,N_12820,N_12695);
or U13663 (N_13663,N_12882,N_12665);
nand U13664 (N_13664,N_12975,N_12645);
and U13665 (N_13665,N_12883,N_12610);
or U13666 (N_13666,N_12699,N_12651);
and U13667 (N_13667,N_12651,N_12998);
nand U13668 (N_13668,N_13093,N_12746);
nand U13669 (N_13669,N_12746,N_12804);
and U13670 (N_13670,N_12808,N_13057);
nor U13671 (N_13671,N_13089,N_12923);
or U13672 (N_13672,N_13063,N_12682);
xnor U13673 (N_13673,N_13006,N_12791);
nand U13674 (N_13674,N_13180,N_12618);
nor U13675 (N_13675,N_13089,N_12983);
or U13676 (N_13676,N_13010,N_12993);
and U13677 (N_13677,N_12770,N_12847);
or U13678 (N_13678,N_12914,N_12641);
or U13679 (N_13679,N_12926,N_12977);
nand U13680 (N_13680,N_12737,N_12848);
and U13681 (N_13681,N_12732,N_12953);
nand U13682 (N_13682,N_12977,N_13095);
or U13683 (N_13683,N_12735,N_12702);
and U13684 (N_13684,N_12686,N_12805);
and U13685 (N_13685,N_12664,N_12760);
nor U13686 (N_13686,N_12749,N_13092);
or U13687 (N_13687,N_12640,N_12992);
or U13688 (N_13688,N_12704,N_12797);
and U13689 (N_13689,N_12781,N_13079);
or U13690 (N_13690,N_12861,N_12983);
nor U13691 (N_13691,N_12761,N_12716);
and U13692 (N_13692,N_12861,N_12993);
and U13693 (N_13693,N_12720,N_12905);
xor U13694 (N_13694,N_12677,N_12646);
or U13695 (N_13695,N_12889,N_12964);
nand U13696 (N_13696,N_12841,N_12989);
and U13697 (N_13697,N_12670,N_12632);
nor U13698 (N_13698,N_13089,N_12623);
nand U13699 (N_13699,N_13003,N_12954);
nor U13700 (N_13700,N_13069,N_12647);
and U13701 (N_13701,N_13110,N_12617);
nand U13702 (N_13702,N_12736,N_13053);
and U13703 (N_13703,N_13196,N_12704);
and U13704 (N_13704,N_13159,N_12781);
or U13705 (N_13705,N_13082,N_13097);
or U13706 (N_13706,N_12966,N_12737);
and U13707 (N_13707,N_13081,N_13066);
or U13708 (N_13708,N_12899,N_12889);
nand U13709 (N_13709,N_12834,N_12886);
and U13710 (N_13710,N_13151,N_13099);
nand U13711 (N_13711,N_13015,N_12661);
or U13712 (N_13712,N_12678,N_12884);
xor U13713 (N_13713,N_12698,N_13050);
nand U13714 (N_13714,N_12778,N_13042);
and U13715 (N_13715,N_13075,N_12883);
nand U13716 (N_13716,N_12699,N_13141);
nand U13717 (N_13717,N_13193,N_12958);
nand U13718 (N_13718,N_13119,N_12789);
and U13719 (N_13719,N_12786,N_12760);
nor U13720 (N_13720,N_13107,N_13073);
or U13721 (N_13721,N_12633,N_12773);
nand U13722 (N_13722,N_12963,N_12684);
nor U13723 (N_13723,N_13028,N_13093);
and U13724 (N_13724,N_12631,N_12892);
or U13725 (N_13725,N_12636,N_12712);
nand U13726 (N_13726,N_13114,N_12856);
or U13727 (N_13727,N_12924,N_12883);
or U13728 (N_13728,N_12969,N_13040);
or U13729 (N_13729,N_12833,N_13090);
xnor U13730 (N_13730,N_12719,N_12875);
nor U13731 (N_13731,N_12870,N_12609);
or U13732 (N_13732,N_13172,N_12674);
or U13733 (N_13733,N_12755,N_12733);
and U13734 (N_13734,N_12632,N_13199);
nor U13735 (N_13735,N_13083,N_13122);
or U13736 (N_13736,N_12984,N_12676);
nand U13737 (N_13737,N_12817,N_12741);
and U13738 (N_13738,N_12887,N_12732);
and U13739 (N_13739,N_12776,N_13145);
or U13740 (N_13740,N_12821,N_12811);
nor U13741 (N_13741,N_12812,N_12734);
nor U13742 (N_13742,N_13009,N_12726);
or U13743 (N_13743,N_12660,N_12894);
nand U13744 (N_13744,N_13048,N_12743);
and U13745 (N_13745,N_13044,N_12726);
nand U13746 (N_13746,N_12619,N_13073);
and U13747 (N_13747,N_12806,N_12852);
or U13748 (N_13748,N_12801,N_12719);
and U13749 (N_13749,N_12947,N_13136);
nor U13750 (N_13750,N_13016,N_12828);
nand U13751 (N_13751,N_13111,N_12865);
and U13752 (N_13752,N_12876,N_12716);
nand U13753 (N_13753,N_12825,N_13038);
or U13754 (N_13754,N_13080,N_12841);
nand U13755 (N_13755,N_12759,N_12740);
nand U13756 (N_13756,N_13190,N_12651);
nor U13757 (N_13757,N_12682,N_12643);
or U13758 (N_13758,N_13031,N_12602);
nor U13759 (N_13759,N_12780,N_12674);
or U13760 (N_13760,N_13042,N_13098);
nand U13761 (N_13761,N_13009,N_12692);
nand U13762 (N_13762,N_12630,N_12672);
nand U13763 (N_13763,N_13018,N_12740);
nand U13764 (N_13764,N_12611,N_13129);
nand U13765 (N_13765,N_13115,N_13036);
nand U13766 (N_13766,N_12967,N_13005);
nand U13767 (N_13767,N_13166,N_12838);
nand U13768 (N_13768,N_13134,N_12846);
and U13769 (N_13769,N_13021,N_12778);
nand U13770 (N_13770,N_12627,N_13082);
nor U13771 (N_13771,N_12687,N_12766);
or U13772 (N_13772,N_12611,N_13111);
nand U13773 (N_13773,N_13025,N_12849);
nor U13774 (N_13774,N_12968,N_13080);
and U13775 (N_13775,N_12742,N_12924);
nor U13776 (N_13776,N_12831,N_12652);
and U13777 (N_13777,N_12814,N_12676);
and U13778 (N_13778,N_12849,N_12710);
nand U13779 (N_13779,N_12604,N_12717);
nand U13780 (N_13780,N_12765,N_12801);
or U13781 (N_13781,N_12677,N_12728);
or U13782 (N_13782,N_12920,N_12744);
or U13783 (N_13783,N_13172,N_12875);
nand U13784 (N_13784,N_12822,N_13081);
nand U13785 (N_13785,N_12714,N_12600);
or U13786 (N_13786,N_12788,N_13059);
nand U13787 (N_13787,N_12784,N_12920);
nand U13788 (N_13788,N_12848,N_13156);
nand U13789 (N_13789,N_12648,N_13144);
and U13790 (N_13790,N_12724,N_12617);
and U13791 (N_13791,N_12937,N_13074);
and U13792 (N_13792,N_13017,N_12889);
nand U13793 (N_13793,N_12621,N_12862);
and U13794 (N_13794,N_12860,N_12709);
or U13795 (N_13795,N_12663,N_12992);
nor U13796 (N_13796,N_12735,N_12834);
xor U13797 (N_13797,N_13118,N_12759);
nor U13798 (N_13798,N_13117,N_13196);
or U13799 (N_13799,N_12917,N_13041);
nand U13800 (N_13800,N_13617,N_13375);
or U13801 (N_13801,N_13433,N_13605);
nand U13802 (N_13802,N_13358,N_13292);
or U13803 (N_13803,N_13792,N_13265);
nand U13804 (N_13804,N_13590,N_13296);
nand U13805 (N_13805,N_13780,N_13319);
nand U13806 (N_13806,N_13514,N_13232);
nor U13807 (N_13807,N_13418,N_13364);
nor U13808 (N_13808,N_13528,N_13220);
and U13809 (N_13809,N_13578,N_13636);
and U13810 (N_13810,N_13260,N_13356);
or U13811 (N_13811,N_13659,N_13299);
and U13812 (N_13812,N_13350,N_13304);
nor U13813 (N_13813,N_13287,N_13487);
nor U13814 (N_13814,N_13774,N_13349);
or U13815 (N_13815,N_13286,N_13308);
nor U13816 (N_13816,N_13750,N_13703);
and U13817 (N_13817,N_13718,N_13523);
and U13818 (N_13818,N_13236,N_13243);
or U13819 (N_13819,N_13479,N_13744);
nor U13820 (N_13820,N_13687,N_13682);
xnor U13821 (N_13821,N_13639,N_13776);
nor U13822 (N_13822,N_13627,N_13383);
nand U13823 (N_13823,N_13655,N_13615);
nand U13824 (N_13824,N_13362,N_13507);
nor U13825 (N_13825,N_13440,N_13318);
nor U13826 (N_13826,N_13297,N_13225);
and U13827 (N_13827,N_13711,N_13737);
or U13828 (N_13828,N_13587,N_13591);
nor U13829 (N_13829,N_13261,N_13445);
nor U13830 (N_13830,N_13281,N_13421);
xor U13831 (N_13831,N_13395,N_13416);
nor U13832 (N_13832,N_13326,N_13565);
nand U13833 (N_13833,N_13501,N_13549);
or U13834 (N_13834,N_13380,N_13669);
nor U13835 (N_13835,N_13798,N_13443);
nand U13836 (N_13836,N_13724,N_13613);
or U13837 (N_13837,N_13557,N_13508);
nand U13838 (N_13838,N_13213,N_13715);
or U13839 (N_13839,N_13392,N_13765);
nand U13840 (N_13840,N_13469,N_13431);
nor U13841 (N_13841,N_13527,N_13746);
nor U13842 (N_13842,N_13394,N_13520);
nor U13843 (N_13843,N_13531,N_13550);
nor U13844 (N_13844,N_13716,N_13676);
nand U13845 (N_13845,N_13321,N_13403);
and U13846 (N_13846,N_13582,N_13420);
nor U13847 (N_13847,N_13742,N_13256);
and U13848 (N_13848,N_13496,N_13770);
and U13849 (N_13849,N_13200,N_13551);
nand U13850 (N_13850,N_13450,N_13233);
nand U13851 (N_13851,N_13301,N_13782);
or U13852 (N_13852,N_13570,N_13690);
xor U13853 (N_13853,N_13778,N_13572);
and U13854 (N_13854,N_13675,N_13543);
nor U13855 (N_13855,N_13309,N_13263);
or U13856 (N_13856,N_13542,N_13365);
nand U13857 (N_13857,N_13670,N_13234);
nor U13858 (N_13858,N_13732,N_13315);
nand U13859 (N_13859,N_13586,N_13568);
and U13860 (N_13860,N_13325,N_13579);
nand U13861 (N_13861,N_13666,N_13235);
and U13862 (N_13862,N_13632,N_13757);
nand U13863 (N_13863,N_13665,N_13417);
nor U13864 (N_13864,N_13427,N_13722);
nor U13865 (N_13865,N_13538,N_13288);
or U13866 (N_13866,N_13547,N_13646);
or U13867 (N_13867,N_13644,N_13686);
nand U13868 (N_13868,N_13228,N_13303);
nand U13869 (N_13869,N_13794,N_13634);
and U13870 (N_13870,N_13731,N_13552);
nor U13871 (N_13871,N_13624,N_13787);
or U13872 (N_13872,N_13674,N_13477);
nor U13873 (N_13873,N_13426,N_13516);
nor U13874 (N_13874,N_13635,N_13734);
and U13875 (N_13875,N_13316,N_13663);
and U13876 (N_13876,N_13555,N_13580);
or U13877 (N_13877,N_13495,N_13460);
and U13878 (N_13878,N_13244,N_13438);
or U13879 (N_13879,N_13505,N_13444);
or U13880 (N_13880,N_13667,N_13337);
or U13881 (N_13881,N_13467,N_13313);
nand U13882 (N_13882,N_13201,N_13209);
nand U13883 (N_13883,N_13473,N_13569);
or U13884 (N_13884,N_13249,N_13652);
nor U13885 (N_13885,N_13370,N_13564);
or U13886 (N_13886,N_13504,N_13502);
nand U13887 (N_13887,N_13619,N_13402);
nand U13888 (N_13888,N_13493,N_13576);
and U13889 (N_13889,N_13498,N_13475);
nor U13890 (N_13890,N_13781,N_13728);
nor U13891 (N_13891,N_13412,N_13736);
nand U13892 (N_13892,N_13259,N_13419);
and U13893 (N_13893,N_13341,N_13541);
and U13894 (N_13894,N_13471,N_13526);
or U13895 (N_13895,N_13215,N_13255);
nand U13896 (N_13896,N_13406,N_13714);
and U13897 (N_13897,N_13689,N_13784);
nand U13898 (N_13898,N_13449,N_13306);
nand U13899 (N_13899,N_13628,N_13293);
nor U13900 (N_13900,N_13747,N_13295);
and U13901 (N_13901,N_13310,N_13739);
nand U13902 (N_13902,N_13767,N_13465);
nand U13903 (N_13903,N_13462,N_13434);
nor U13904 (N_13904,N_13422,N_13575);
nor U13905 (N_13905,N_13257,N_13393);
nand U13906 (N_13906,N_13603,N_13229);
and U13907 (N_13907,N_13764,N_13616);
and U13908 (N_13908,N_13577,N_13359);
or U13909 (N_13909,N_13691,N_13441);
and U13910 (N_13910,N_13353,N_13436);
and U13911 (N_13911,N_13335,N_13611);
nand U13912 (N_13912,N_13322,N_13548);
nor U13913 (N_13913,N_13683,N_13214);
nand U13914 (N_13914,N_13583,N_13481);
or U13915 (N_13915,N_13702,N_13269);
or U13916 (N_13916,N_13745,N_13783);
and U13917 (N_13917,N_13428,N_13361);
and U13918 (N_13918,N_13251,N_13276);
nand U13919 (N_13919,N_13668,N_13741);
and U13920 (N_13920,N_13388,N_13283);
nand U13921 (N_13921,N_13696,N_13290);
or U13922 (N_13922,N_13328,N_13386);
and U13923 (N_13923,N_13323,N_13753);
nand U13924 (N_13924,N_13594,N_13777);
or U13925 (N_13925,N_13489,N_13492);
or U13926 (N_13926,N_13414,N_13553);
or U13927 (N_13927,N_13329,N_13484);
and U13928 (N_13928,N_13539,N_13795);
nor U13929 (N_13929,N_13461,N_13435);
nor U13930 (N_13930,N_13270,N_13275);
and U13931 (N_13931,N_13756,N_13793);
and U13932 (N_13932,N_13685,N_13372);
nor U13933 (N_13933,N_13697,N_13749);
nand U13934 (N_13934,N_13314,N_13253);
nor U13935 (N_13935,N_13342,N_13252);
xnor U13936 (N_13936,N_13763,N_13203);
nor U13937 (N_13937,N_13529,N_13410);
or U13938 (N_13938,N_13456,N_13404);
nand U13939 (N_13939,N_13357,N_13369);
or U13940 (N_13940,N_13254,N_13720);
nand U13941 (N_13941,N_13710,N_13660);
or U13942 (N_13942,N_13478,N_13595);
nor U13943 (N_13943,N_13592,N_13684);
or U13944 (N_13944,N_13791,N_13240);
or U13945 (N_13945,N_13327,N_13339);
and U13946 (N_13946,N_13540,N_13497);
or U13947 (N_13947,N_13797,N_13648);
and U13948 (N_13948,N_13250,N_13554);
nand U13949 (N_13949,N_13559,N_13399);
and U13950 (N_13950,N_13298,N_13588);
and U13951 (N_13951,N_13614,N_13246);
and U13952 (N_13952,N_13637,N_13500);
nor U13953 (N_13953,N_13355,N_13786);
and U13954 (N_13954,N_13439,N_13681);
and U13955 (N_13955,N_13464,N_13740);
and U13956 (N_13956,N_13212,N_13647);
nor U13957 (N_13957,N_13704,N_13352);
nand U13958 (N_13958,N_13799,N_13300);
or U13959 (N_13959,N_13340,N_13302);
or U13960 (N_13960,N_13307,N_13790);
xor U13961 (N_13961,N_13241,N_13272);
nor U13962 (N_13962,N_13672,N_13522);
or U13963 (N_13963,N_13772,N_13626);
and U13964 (N_13964,N_13454,N_13205);
nor U13965 (N_13965,N_13796,N_13332);
nor U13966 (N_13966,N_13503,N_13680);
nor U13967 (N_13967,N_13248,N_13584);
xnor U13968 (N_13968,N_13788,N_13204);
or U13969 (N_13969,N_13743,N_13247);
and U13970 (N_13970,N_13769,N_13597);
and U13971 (N_13971,N_13346,N_13515);
or U13972 (N_13972,N_13486,N_13472);
or U13973 (N_13973,N_13566,N_13625);
xor U13974 (N_13974,N_13752,N_13596);
or U13975 (N_13975,N_13537,N_13709);
nor U13976 (N_13976,N_13719,N_13407);
nor U13977 (N_13977,N_13231,N_13482);
nor U13978 (N_13978,N_13649,N_13536);
and U13979 (N_13979,N_13699,N_13760);
or U13980 (N_13980,N_13398,N_13600);
and U13981 (N_13981,N_13618,N_13400);
nor U13982 (N_13982,N_13599,N_13331);
and U13983 (N_13983,N_13723,N_13284);
nand U13984 (N_13984,N_13330,N_13448);
nand U13985 (N_13985,N_13560,N_13242);
and U13986 (N_13986,N_13677,N_13612);
nand U13987 (N_13987,N_13609,N_13266);
or U13988 (N_13988,N_13606,N_13671);
or U13989 (N_13989,N_13621,N_13376);
nand U13990 (N_13990,N_13513,N_13218);
nand U13991 (N_13991,N_13695,N_13657);
nand U13992 (N_13992,N_13707,N_13558);
or U13993 (N_13993,N_13607,N_13294);
or U13994 (N_13994,N_13661,N_13608);
or U13995 (N_13995,N_13447,N_13348);
nor U13996 (N_13996,N_13262,N_13650);
nor U13997 (N_13997,N_13499,N_13207);
nand U13998 (N_13998,N_13645,N_13762);
or U13999 (N_13999,N_13678,N_13629);
nand U14000 (N_14000,N_13239,N_13338);
xnor U14001 (N_14001,N_13396,N_13759);
nand U14002 (N_14002,N_13567,N_13480);
nand U14003 (N_14003,N_13692,N_13382);
nor U14004 (N_14004,N_13509,N_13725);
or U14005 (N_14005,N_13424,N_13491);
nor U14006 (N_14006,N_13630,N_13506);
nand U14007 (N_14007,N_13532,N_13277);
nor U14008 (N_14008,N_13423,N_13571);
and U14009 (N_14009,N_13415,N_13391);
or U14010 (N_14010,N_13589,N_13466);
nor U14011 (N_14011,N_13768,N_13379);
or U14012 (N_14012,N_13384,N_13654);
nor U14013 (N_14013,N_13733,N_13278);
nor U14014 (N_14014,N_13701,N_13221);
and U14015 (N_14015,N_13333,N_13457);
and U14016 (N_14016,N_13688,N_13345);
and U14017 (N_14017,N_13409,N_13754);
or U14018 (N_14018,N_13267,N_13425);
and U14019 (N_14019,N_13642,N_13381);
nand U14020 (N_14020,N_13279,N_13641);
nor U14021 (N_14021,N_13653,N_13713);
or U14022 (N_14022,N_13429,N_13411);
nor U14023 (N_14023,N_13217,N_13490);
or U14024 (N_14024,N_13602,N_13771);
and U14025 (N_14025,N_13620,N_13282);
nor U14026 (N_14026,N_13700,N_13534);
and U14027 (N_14027,N_13755,N_13775);
nor U14028 (N_14028,N_13694,N_13389);
and U14029 (N_14029,N_13698,N_13758);
nor U14030 (N_14030,N_13658,N_13773);
nand U14031 (N_14031,N_13216,N_13211);
or U14032 (N_14032,N_13387,N_13459);
nand U14033 (N_14033,N_13623,N_13374);
and U14034 (N_14034,N_13633,N_13738);
xor U14035 (N_14035,N_13408,N_13285);
nor U14036 (N_14036,N_13727,N_13610);
nand U14037 (N_14037,N_13785,N_13779);
or U14038 (N_14038,N_13224,N_13271);
or U14039 (N_14039,N_13320,N_13483);
and U14040 (N_14040,N_13521,N_13470);
or U14041 (N_14041,N_13226,N_13643);
nand U14042 (N_14042,N_13761,N_13468);
nor U14043 (N_14043,N_13730,N_13206);
and U14044 (N_14044,N_13343,N_13601);
nand U14045 (N_14045,N_13789,N_13706);
or U14046 (N_14046,N_13367,N_13517);
and U14047 (N_14047,N_13237,N_13693);
or U14048 (N_14048,N_13662,N_13377);
nor U14049 (N_14049,N_13351,N_13494);
and U14050 (N_14050,N_13258,N_13453);
xor U14051 (N_14051,N_13360,N_13530);
or U14052 (N_14052,N_13413,N_13485);
and U14053 (N_14053,N_13452,N_13230);
nor U14054 (N_14054,N_13268,N_13312);
nor U14055 (N_14055,N_13368,N_13474);
and U14056 (N_14056,N_13510,N_13446);
nand U14057 (N_14057,N_13581,N_13317);
or U14058 (N_14058,N_13430,N_13533);
nor U14059 (N_14059,N_13476,N_13324);
and U14060 (N_14060,N_13712,N_13638);
and U14061 (N_14061,N_13721,N_13545);
nor U14062 (N_14062,N_13640,N_13664);
or U14063 (N_14063,N_13405,N_13598);
or U14064 (N_14064,N_13524,N_13651);
nand U14065 (N_14065,N_13378,N_13766);
nand U14066 (N_14066,N_13202,N_13673);
or U14067 (N_14067,N_13544,N_13535);
nor U14068 (N_14068,N_13280,N_13726);
nor U14069 (N_14069,N_13305,N_13735);
nor U14070 (N_14070,N_13748,N_13622);
and U14071 (N_14071,N_13390,N_13344);
nand U14072 (N_14072,N_13366,N_13291);
and U14073 (N_14073,N_13401,N_13512);
nor U14074 (N_14074,N_13631,N_13373);
nor U14075 (N_14075,N_13238,N_13311);
nor U14076 (N_14076,N_13593,N_13455);
nor U14077 (N_14077,N_13463,N_13264);
or U14078 (N_14078,N_13708,N_13371);
nor U14079 (N_14079,N_13511,N_13518);
nand U14080 (N_14080,N_13556,N_13432);
nand U14081 (N_14081,N_13385,N_13222);
and U14082 (N_14082,N_13397,N_13574);
and U14083 (N_14083,N_13519,N_13458);
and U14084 (N_14084,N_13563,N_13437);
and U14085 (N_14085,N_13223,N_13227);
or U14086 (N_14086,N_13573,N_13525);
nor U14087 (N_14087,N_13336,N_13219);
nand U14088 (N_14088,N_13585,N_13546);
nor U14089 (N_14089,N_13717,N_13656);
nand U14090 (N_14090,N_13751,N_13488);
nor U14091 (N_14091,N_13363,N_13347);
and U14092 (N_14092,N_13210,N_13354);
nor U14093 (N_14093,N_13334,N_13274);
and U14094 (N_14094,N_13451,N_13679);
or U14095 (N_14095,N_13729,N_13208);
nor U14096 (N_14096,N_13442,N_13245);
and U14097 (N_14097,N_13273,N_13289);
nand U14098 (N_14098,N_13604,N_13561);
or U14099 (N_14099,N_13705,N_13562);
nor U14100 (N_14100,N_13712,N_13688);
nor U14101 (N_14101,N_13666,N_13466);
and U14102 (N_14102,N_13309,N_13602);
nor U14103 (N_14103,N_13400,N_13238);
nand U14104 (N_14104,N_13263,N_13207);
nand U14105 (N_14105,N_13397,N_13265);
nor U14106 (N_14106,N_13518,N_13369);
nand U14107 (N_14107,N_13463,N_13403);
nor U14108 (N_14108,N_13321,N_13654);
nor U14109 (N_14109,N_13792,N_13412);
nand U14110 (N_14110,N_13544,N_13423);
and U14111 (N_14111,N_13313,N_13348);
nand U14112 (N_14112,N_13629,N_13436);
nor U14113 (N_14113,N_13693,N_13269);
and U14114 (N_14114,N_13442,N_13345);
or U14115 (N_14115,N_13350,N_13520);
nand U14116 (N_14116,N_13283,N_13641);
or U14117 (N_14117,N_13756,N_13500);
nor U14118 (N_14118,N_13244,N_13459);
and U14119 (N_14119,N_13212,N_13566);
nor U14120 (N_14120,N_13474,N_13288);
nand U14121 (N_14121,N_13498,N_13779);
nor U14122 (N_14122,N_13742,N_13522);
nor U14123 (N_14123,N_13609,N_13344);
and U14124 (N_14124,N_13308,N_13395);
nand U14125 (N_14125,N_13683,N_13578);
or U14126 (N_14126,N_13726,N_13470);
xnor U14127 (N_14127,N_13754,N_13633);
or U14128 (N_14128,N_13394,N_13628);
or U14129 (N_14129,N_13522,N_13675);
and U14130 (N_14130,N_13546,N_13772);
or U14131 (N_14131,N_13776,N_13233);
xor U14132 (N_14132,N_13629,N_13588);
and U14133 (N_14133,N_13366,N_13558);
nand U14134 (N_14134,N_13411,N_13273);
nand U14135 (N_14135,N_13510,N_13758);
nand U14136 (N_14136,N_13323,N_13525);
or U14137 (N_14137,N_13231,N_13704);
or U14138 (N_14138,N_13356,N_13330);
and U14139 (N_14139,N_13671,N_13431);
nand U14140 (N_14140,N_13784,N_13458);
or U14141 (N_14141,N_13688,N_13298);
and U14142 (N_14142,N_13248,N_13609);
and U14143 (N_14143,N_13435,N_13667);
nand U14144 (N_14144,N_13232,N_13395);
nand U14145 (N_14145,N_13721,N_13367);
nor U14146 (N_14146,N_13443,N_13505);
or U14147 (N_14147,N_13645,N_13502);
nor U14148 (N_14148,N_13595,N_13352);
or U14149 (N_14149,N_13709,N_13601);
nor U14150 (N_14150,N_13457,N_13362);
and U14151 (N_14151,N_13246,N_13676);
nor U14152 (N_14152,N_13523,N_13510);
and U14153 (N_14153,N_13398,N_13444);
and U14154 (N_14154,N_13270,N_13608);
and U14155 (N_14155,N_13774,N_13438);
nor U14156 (N_14156,N_13742,N_13322);
and U14157 (N_14157,N_13591,N_13293);
or U14158 (N_14158,N_13516,N_13333);
or U14159 (N_14159,N_13751,N_13613);
nand U14160 (N_14160,N_13345,N_13716);
or U14161 (N_14161,N_13701,N_13318);
nor U14162 (N_14162,N_13701,N_13749);
nand U14163 (N_14163,N_13791,N_13392);
and U14164 (N_14164,N_13270,N_13469);
nand U14165 (N_14165,N_13421,N_13777);
nand U14166 (N_14166,N_13476,N_13628);
nand U14167 (N_14167,N_13352,N_13706);
nor U14168 (N_14168,N_13512,N_13293);
nand U14169 (N_14169,N_13659,N_13751);
nand U14170 (N_14170,N_13354,N_13564);
xnor U14171 (N_14171,N_13493,N_13395);
nor U14172 (N_14172,N_13261,N_13544);
nand U14173 (N_14173,N_13574,N_13559);
and U14174 (N_14174,N_13434,N_13448);
nand U14175 (N_14175,N_13410,N_13697);
or U14176 (N_14176,N_13681,N_13545);
nand U14177 (N_14177,N_13481,N_13759);
or U14178 (N_14178,N_13752,N_13706);
and U14179 (N_14179,N_13632,N_13489);
nor U14180 (N_14180,N_13299,N_13212);
and U14181 (N_14181,N_13474,N_13627);
or U14182 (N_14182,N_13589,N_13554);
nor U14183 (N_14183,N_13480,N_13592);
or U14184 (N_14184,N_13779,N_13747);
or U14185 (N_14185,N_13339,N_13711);
nor U14186 (N_14186,N_13774,N_13295);
or U14187 (N_14187,N_13213,N_13302);
nand U14188 (N_14188,N_13694,N_13471);
nand U14189 (N_14189,N_13329,N_13247);
or U14190 (N_14190,N_13329,N_13440);
nand U14191 (N_14191,N_13461,N_13689);
nor U14192 (N_14192,N_13794,N_13554);
nor U14193 (N_14193,N_13338,N_13636);
nand U14194 (N_14194,N_13424,N_13279);
xor U14195 (N_14195,N_13409,N_13782);
nor U14196 (N_14196,N_13371,N_13637);
xor U14197 (N_14197,N_13485,N_13491);
nor U14198 (N_14198,N_13281,N_13729);
or U14199 (N_14199,N_13608,N_13645);
and U14200 (N_14200,N_13712,N_13622);
nand U14201 (N_14201,N_13222,N_13711);
and U14202 (N_14202,N_13527,N_13426);
or U14203 (N_14203,N_13709,N_13606);
or U14204 (N_14204,N_13555,N_13422);
nor U14205 (N_14205,N_13780,N_13222);
or U14206 (N_14206,N_13449,N_13443);
and U14207 (N_14207,N_13751,N_13276);
and U14208 (N_14208,N_13485,N_13322);
or U14209 (N_14209,N_13590,N_13233);
or U14210 (N_14210,N_13711,N_13271);
nand U14211 (N_14211,N_13685,N_13464);
nor U14212 (N_14212,N_13466,N_13552);
and U14213 (N_14213,N_13459,N_13499);
and U14214 (N_14214,N_13638,N_13413);
or U14215 (N_14215,N_13294,N_13639);
and U14216 (N_14216,N_13258,N_13203);
nand U14217 (N_14217,N_13437,N_13643);
and U14218 (N_14218,N_13329,N_13286);
or U14219 (N_14219,N_13733,N_13581);
nand U14220 (N_14220,N_13448,N_13258);
and U14221 (N_14221,N_13694,N_13209);
nor U14222 (N_14222,N_13244,N_13355);
or U14223 (N_14223,N_13419,N_13785);
or U14224 (N_14224,N_13617,N_13725);
nand U14225 (N_14225,N_13793,N_13629);
and U14226 (N_14226,N_13787,N_13312);
and U14227 (N_14227,N_13283,N_13475);
and U14228 (N_14228,N_13654,N_13503);
and U14229 (N_14229,N_13786,N_13290);
nor U14230 (N_14230,N_13517,N_13552);
and U14231 (N_14231,N_13497,N_13262);
nand U14232 (N_14232,N_13558,N_13278);
and U14233 (N_14233,N_13531,N_13650);
nor U14234 (N_14234,N_13292,N_13734);
nand U14235 (N_14235,N_13546,N_13318);
and U14236 (N_14236,N_13228,N_13339);
nand U14237 (N_14237,N_13569,N_13210);
and U14238 (N_14238,N_13583,N_13732);
nor U14239 (N_14239,N_13328,N_13654);
and U14240 (N_14240,N_13476,N_13378);
or U14241 (N_14241,N_13268,N_13261);
nor U14242 (N_14242,N_13489,N_13271);
or U14243 (N_14243,N_13698,N_13331);
or U14244 (N_14244,N_13631,N_13259);
and U14245 (N_14245,N_13264,N_13399);
or U14246 (N_14246,N_13473,N_13556);
nand U14247 (N_14247,N_13729,N_13206);
and U14248 (N_14248,N_13595,N_13327);
and U14249 (N_14249,N_13423,N_13649);
and U14250 (N_14250,N_13315,N_13492);
and U14251 (N_14251,N_13233,N_13661);
nor U14252 (N_14252,N_13723,N_13763);
nand U14253 (N_14253,N_13232,N_13262);
nand U14254 (N_14254,N_13218,N_13746);
nand U14255 (N_14255,N_13597,N_13687);
and U14256 (N_14256,N_13619,N_13468);
and U14257 (N_14257,N_13375,N_13764);
and U14258 (N_14258,N_13409,N_13639);
and U14259 (N_14259,N_13375,N_13663);
nor U14260 (N_14260,N_13736,N_13477);
xnor U14261 (N_14261,N_13250,N_13643);
or U14262 (N_14262,N_13380,N_13304);
and U14263 (N_14263,N_13237,N_13389);
xnor U14264 (N_14264,N_13500,N_13338);
and U14265 (N_14265,N_13551,N_13556);
nand U14266 (N_14266,N_13284,N_13302);
nor U14267 (N_14267,N_13669,N_13282);
nand U14268 (N_14268,N_13651,N_13415);
or U14269 (N_14269,N_13640,N_13250);
nor U14270 (N_14270,N_13548,N_13483);
or U14271 (N_14271,N_13643,N_13319);
and U14272 (N_14272,N_13679,N_13405);
and U14273 (N_14273,N_13526,N_13538);
and U14274 (N_14274,N_13505,N_13775);
nand U14275 (N_14275,N_13448,N_13624);
nor U14276 (N_14276,N_13767,N_13277);
xor U14277 (N_14277,N_13788,N_13430);
and U14278 (N_14278,N_13591,N_13780);
nor U14279 (N_14279,N_13505,N_13496);
nor U14280 (N_14280,N_13608,N_13244);
or U14281 (N_14281,N_13208,N_13397);
nor U14282 (N_14282,N_13275,N_13312);
nor U14283 (N_14283,N_13734,N_13377);
nand U14284 (N_14284,N_13393,N_13755);
or U14285 (N_14285,N_13218,N_13566);
or U14286 (N_14286,N_13565,N_13620);
xnor U14287 (N_14287,N_13720,N_13545);
and U14288 (N_14288,N_13565,N_13364);
nand U14289 (N_14289,N_13332,N_13236);
nand U14290 (N_14290,N_13665,N_13387);
nand U14291 (N_14291,N_13429,N_13508);
and U14292 (N_14292,N_13718,N_13211);
nand U14293 (N_14293,N_13253,N_13693);
or U14294 (N_14294,N_13388,N_13721);
nand U14295 (N_14295,N_13693,N_13601);
or U14296 (N_14296,N_13700,N_13525);
nor U14297 (N_14297,N_13545,N_13252);
and U14298 (N_14298,N_13574,N_13381);
nor U14299 (N_14299,N_13611,N_13479);
nand U14300 (N_14300,N_13750,N_13359);
or U14301 (N_14301,N_13570,N_13776);
nand U14302 (N_14302,N_13226,N_13652);
nand U14303 (N_14303,N_13382,N_13555);
nor U14304 (N_14304,N_13470,N_13669);
and U14305 (N_14305,N_13552,N_13433);
and U14306 (N_14306,N_13608,N_13289);
and U14307 (N_14307,N_13427,N_13586);
nor U14308 (N_14308,N_13678,N_13641);
nor U14309 (N_14309,N_13518,N_13424);
nor U14310 (N_14310,N_13521,N_13529);
or U14311 (N_14311,N_13369,N_13720);
nor U14312 (N_14312,N_13648,N_13221);
nand U14313 (N_14313,N_13588,N_13766);
and U14314 (N_14314,N_13746,N_13613);
or U14315 (N_14315,N_13302,N_13682);
nand U14316 (N_14316,N_13563,N_13220);
nand U14317 (N_14317,N_13473,N_13524);
or U14318 (N_14318,N_13664,N_13319);
or U14319 (N_14319,N_13655,N_13671);
or U14320 (N_14320,N_13400,N_13437);
and U14321 (N_14321,N_13477,N_13263);
nand U14322 (N_14322,N_13591,N_13789);
nor U14323 (N_14323,N_13598,N_13294);
nor U14324 (N_14324,N_13778,N_13725);
nand U14325 (N_14325,N_13509,N_13768);
and U14326 (N_14326,N_13743,N_13389);
or U14327 (N_14327,N_13563,N_13423);
nor U14328 (N_14328,N_13688,N_13758);
nor U14329 (N_14329,N_13738,N_13609);
nand U14330 (N_14330,N_13799,N_13460);
or U14331 (N_14331,N_13683,N_13661);
nor U14332 (N_14332,N_13640,N_13415);
nor U14333 (N_14333,N_13301,N_13688);
nor U14334 (N_14334,N_13313,N_13540);
or U14335 (N_14335,N_13468,N_13719);
nand U14336 (N_14336,N_13537,N_13504);
nor U14337 (N_14337,N_13358,N_13356);
nor U14338 (N_14338,N_13755,N_13398);
or U14339 (N_14339,N_13561,N_13437);
or U14340 (N_14340,N_13603,N_13793);
or U14341 (N_14341,N_13211,N_13624);
nand U14342 (N_14342,N_13336,N_13211);
or U14343 (N_14343,N_13360,N_13434);
and U14344 (N_14344,N_13201,N_13706);
xnor U14345 (N_14345,N_13445,N_13615);
or U14346 (N_14346,N_13756,N_13798);
or U14347 (N_14347,N_13494,N_13226);
and U14348 (N_14348,N_13703,N_13337);
nand U14349 (N_14349,N_13526,N_13600);
nand U14350 (N_14350,N_13305,N_13464);
and U14351 (N_14351,N_13489,N_13490);
or U14352 (N_14352,N_13706,N_13307);
nand U14353 (N_14353,N_13488,N_13323);
nand U14354 (N_14354,N_13323,N_13583);
or U14355 (N_14355,N_13379,N_13344);
nor U14356 (N_14356,N_13635,N_13344);
and U14357 (N_14357,N_13382,N_13224);
or U14358 (N_14358,N_13393,N_13267);
and U14359 (N_14359,N_13262,N_13713);
nor U14360 (N_14360,N_13291,N_13566);
and U14361 (N_14361,N_13396,N_13412);
nand U14362 (N_14362,N_13480,N_13683);
nand U14363 (N_14363,N_13300,N_13266);
and U14364 (N_14364,N_13705,N_13753);
xor U14365 (N_14365,N_13558,N_13789);
nand U14366 (N_14366,N_13356,N_13208);
or U14367 (N_14367,N_13494,N_13304);
or U14368 (N_14368,N_13628,N_13581);
or U14369 (N_14369,N_13372,N_13388);
or U14370 (N_14370,N_13603,N_13726);
and U14371 (N_14371,N_13639,N_13299);
or U14372 (N_14372,N_13755,N_13780);
or U14373 (N_14373,N_13497,N_13794);
or U14374 (N_14374,N_13785,N_13315);
nand U14375 (N_14375,N_13587,N_13597);
and U14376 (N_14376,N_13631,N_13395);
and U14377 (N_14377,N_13753,N_13219);
nor U14378 (N_14378,N_13557,N_13552);
and U14379 (N_14379,N_13554,N_13679);
and U14380 (N_14380,N_13767,N_13709);
and U14381 (N_14381,N_13532,N_13580);
or U14382 (N_14382,N_13532,N_13544);
or U14383 (N_14383,N_13628,N_13700);
nand U14384 (N_14384,N_13775,N_13285);
nand U14385 (N_14385,N_13621,N_13304);
nand U14386 (N_14386,N_13342,N_13242);
nor U14387 (N_14387,N_13723,N_13342);
and U14388 (N_14388,N_13299,N_13308);
nor U14389 (N_14389,N_13583,N_13492);
and U14390 (N_14390,N_13746,N_13637);
or U14391 (N_14391,N_13726,N_13707);
or U14392 (N_14392,N_13328,N_13245);
nand U14393 (N_14393,N_13684,N_13245);
and U14394 (N_14394,N_13713,N_13201);
or U14395 (N_14395,N_13629,N_13774);
nor U14396 (N_14396,N_13590,N_13500);
nor U14397 (N_14397,N_13324,N_13625);
nor U14398 (N_14398,N_13360,N_13512);
or U14399 (N_14399,N_13631,N_13323);
nand U14400 (N_14400,N_14259,N_14302);
or U14401 (N_14401,N_14159,N_13965);
nand U14402 (N_14402,N_14037,N_14080);
nor U14403 (N_14403,N_13942,N_14209);
and U14404 (N_14404,N_14333,N_14366);
nor U14405 (N_14405,N_13984,N_13996);
or U14406 (N_14406,N_14177,N_13820);
and U14407 (N_14407,N_14065,N_14072);
and U14408 (N_14408,N_14237,N_14018);
xor U14409 (N_14409,N_14172,N_13828);
or U14410 (N_14410,N_14033,N_14120);
or U14411 (N_14411,N_14055,N_14389);
or U14412 (N_14412,N_14359,N_14283);
and U14413 (N_14413,N_14145,N_14232);
or U14414 (N_14414,N_14305,N_14211);
nor U14415 (N_14415,N_14287,N_13811);
nand U14416 (N_14416,N_14139,N_14016);
and U14417 (N_14417,N_13903,N_14027);
nor U14418 (N_14418,N_13954,N_14187);
or U14419 (N_14419,N_14311,N_14089);
nand U14420 (N_14420,N_14167,N_14102);
nor U14421 (N_14421,N_14024,N_14032);
nor U14422 (N_14422,N_14298,N_13936);
nand U14423 (N_14423,N_14056,N_13815);
nor U14424 (N_14424,N_13976,N_14173);
or U14425 (N_14425,N_13899,N_14214);
and U14426 (N_14426,N_14003,N_14260);
and U14427 (N_14427,N_14193,N_14281);
nor U14428 (N_14428,N_14247,N_13836);
and U14429 (N_14429,N_14251,N_13999);
or U14430 (N_14430,N_14157,N_14184);
and U14431 (N_14431,N_14023,N_14227);
nor U14432 (N_14432,N_14367,N_14108);
or U14433 (N_14433,N_14257,N_14236);
or U14434 (N_14434,N_14069,N_14061);
or U14435 (N_14435,N_14011,N_14097);
nor U14436 (N_14436,N_14132,N_14352);
nor U14437 (N_14437,N_14385,N_14291);
or U14438 (N_14438,N_14078,N_14031);
or U14439 (N_14439,N_14250,N_14158);
or U14440 (N_14440,N_14319,N_13978);
nand U14441 (N_14441,N_14354,N_14077);
and U14442 (N_14442,N_14253,N_13961);
or U14443 (N_14443,N_14240,N_14142);
or U14444 (N_14444,N_14269,N_14345);
or U14445 (N_14445,N_14264,N_14249);
and U14446 (N_14446,N_14096,N_14046);
nor U14447 (N_14447,N_14383,N_13947);
and U14448 (N_14448,N_13931,N_13887);
nor U14449 (N_14449,N_14397,N_13925);
nand U14450 (N_14450,N_14064,N_13983);
or U14451 (N_14451,N_13987,N_14121);
nor U14452 (N_14452,N_14161,N_14165);
and U14453 (N_14453,N_14369,N_14112);
or U14454 (N_14454,N_13813,N_14106);
nor U14455 (N_14455,N_14190,N_13902);
and U14456 (N_14456,N_13824,N_13840);
nor U14457 (N_14457,N_13918,N_14054);
or U14458 (N_14458,N_14030,N_13881);
nand U14459 (N_14459,N_14109,N_13846);
or U14460 (N_14460,N_14143,N_14356);
nor U14461 (N_14461,N_13974,N_14379);
nor U14462 (N_14462,N_14344,N_14169);
nor U14463 (N_14463,N_13821,N_14199);
nand U14464 (N_14464,N_14289,N_14196);
nand U14465 (N_14465,N_13885,N_13952);
nor U14466 (N_14466,N_13938,N_14194);
nand U14467 (N_14467,N_14085,N_14215);
nand U14468 (N_14468,N_14323,N_14270);
or U14469 (N_14469,N_13837,N_13805);
and U14470 (N_14470,N_14244,N_14342);
nand U14471 (N_14471,N_14198,N_14039);
or U14472 (N_14472,N_14206,N_14268);
nand U14473 (N_14473,N_14006,N_14233);
or U14474 (N_14474,N_13893,N_13891);
nor U14475 (N_14475,N_14241,N_14375);
nand U14476 (N_14476,N_13964,N_13913);
nand U14477 (N_14477,N_14224,N_14315);
nand U14478 (N_14478,N_14144,N_13814);
nand U14479 (N_14479,N_14163,N_14294);
nor U14480 (N_14480,N_14252,N_14380);
and U14481 (N_14481,N_13872,N_13868);
or U14482 (N_14482,N_13997,N_14047);
nand U14483 (N_14483,N_14357,N_14266);
xnor U14484 (N_14484,N_13839,N_14365);
nor U14485 (N_14485,N_13924,N_14392);
and U14486 (N_14486,N_14149,N_14125);
nor U14487 (N_14487,N_13803,N_14063);
nand U14488 (N_14488,N_14374,N_14160);
nor U14489 (N_14489,N_14044,N_13843);
or U14490 (N_14490,N_13800,N_13930);
nand U14491 (N_14491,N_14141,N_13934);
and U14492 (N_14492,N_14221,N_14022);
or U14493 (N_14493,N_14098,N_13898);
nor U14494 (N_14494,N_14310,N_14295);
and U14495 (N_14495,N_14175,N_14092);
nor U14496 (N_14496,N_14238,N_14256);
or U14497 (N_14497,N_14088,N_14373);
or U14498 (N_14498,N_14148,N_13829);
and U14499 (N_14499,N_14179,N_13856);
nor U14500 (N_14500,N_14384,N_13919);
and U14501 (N_14501,N_13994,N_13900);
and U14502 (N_14502,N_14317,N_13946);
or U14503 (N_14503,N_14395,N_13897);
nand U14504 (N_14504,N_14231,N_14245);
nand U14505 (N_14505,N_14126,N_14279);
nor U14506 (N_14506,N_13816,N_14396);
and U14507 (N_14507,N_13857,N_13859);
nand U14508 (N_14508,N_13962,N_14363);
and U14509 (N_14509,N_14318,N_14189);
or U14510 (N_14510,N_14082,N_13890);
and U14511 (N_14511,N_13990,N_13949);
nand U14512 (N_14512,N_13831,N_14192);
nor U14513 (N_14513,N_13826,N_13921);
nand U14514 (N_14514,N_13993,N_14049);
nor U14515 (N_14515,N_14201,N_14288);
nand U14516 (N_14516,N_14176,N_13810);
nand U14517 (N_14517,N_14019,N_14242);
nor U14518 (N_14518,N_14079,N_13982);
nor U14519 (N_14519,N_14327,N_14262);
and U14520 (N_14520,N_14335,N_14329);
nor U14521 (N_14521,N_13928,N_13876);
and U14522 (N_14522,N_14219,N_14336);
nand U14523 (N_14523,N_14355,N_14217);
nand U14524 (N_14524,N_13827,N_13933);
and U14525 (N_14525,N_13822,N_14312);
nand U14526 (N_14526,N_14068,N_14014);
or U14527 (N_14527,N_14113,N_14324);
and U14528 (N_14528,N_14071,N_14301);
nor U14529 (N_14529,N_13972,N_14292);
nor U14530 (N_14530,N_14028,N_14343);
nor U14531 (N_14531,N_14183,N_13943);
nor U14532 (N_14532,N_14050,N_14337);
or U14533 (N_14533,N_13851,N_14076);
or U14534 (N_14534,N_14115,N_14204);
xnor U14535 (N_14535,N_13960,N_14225);
or U14536 (N_14536,N_13869,N_14099);
nor U14537 (N_14537,N_14186,N_14391);
nor U14538 (N_14538,N_14012,N_13927);
and U14539 (N_14539,N_13825,N_14104);
nand U14540 (N_14540,N_14146,N_13904);
or U14541 (N_14541,N_14358,N_14191);
and U14542 (N_14542,N_14107,N_13920);
nor U14543 (N_14543,N_14307,N_14368);
and U14544 (N_14544,N_13873,N_14001);
and U14545 (N_14545,N_13807,N_13981);
nor U14546 (N_14546,N_14029,N_13830);
nand U14547 (N_14547,N_14210,N_14116);
or U14548 (N_14548,N_13998,N_14205);
nor U14549 (N_14549,N_13923,N_13854);
nand U14550 (N_14550,N_13939,N_14220);
nor U14551 (N_14551,N_13917,N_14338);
and U14552 (N_14552,N_13958,N_14004);
or U14553 (N_14553,N_14300,N_13833);
or U14554 (N_14554,N_13888,N_13915);
nor U14555 (N_14555,N_14273,N_14168);
nor U14556 (N_14556,N_13907,N_14276);
nor U14557 (N_14557,N_14372,N_14185);
nand U14558 (N_14558,N_13845,N_13989);
nor U14559 (N_14559,N_14258,N_14015);
or U14560 (N_14560,N_14347,N_14330);
nand U14561 (N_14561,N_14025,N_13971);
nor U14562 (N_14562,N_14008,N_14341);
and U14563 (N_14563,N_13986,N_13944);
or U14564 (N_14564,N_14156,N_14362);
nor U14565 (N_14565,N_14293,N_14129);
nand U14566 (N_14566,N_14314,N_14361);
or U14567 (N_14567,N_14017,N_14285);
nor U14568 (N_14568,N_14026,N_14133);
nand U14569 (N_14569,N_14306,N_14328);
or U14570 (N_14570,N_13973,N_13916);
nor U14571 (N_14571,N_14043,N_14095);
nand U14572 (N_14572,N_14230,N_13975);
nor U14573 (N_14573,N_14000,N_13855);
nand U14574 (N_14574,N_14267,N_14325);
or U14575 (N_14575,N_14042,N_14218);
or U14576 (N_14576,N_13980,N_13844);
nor U14577 (N_14577,N_13867,N_13860);
or U14578 (N_14578,N_14331,N_13848);
and U14579 (N_14579,N_13883,N_14213);
nand U14580 (N_14580,N_14282,N_14274);
nand U14581 (N_14581,N_14111,N_14370);
and U14582 (N_14582,N_13849,N_14087);
or U14583 (N_14583,N_13992,N_14309);
nand U14584 (N_14584,N_13922,N_13968);
nor U14585 (N_14585,N_13834,N_14075);
or U14586 (N_14586,N_14313,N_13852);
nor U14587 (N_14587,N_13911,N_14128);
and U14588 (N_14588,N_13870,N_13967);
or U14589 (N_14589,N_14284,N_13926);
or U14590 (N_14590,N_14135,N_13901);
and U14591 (N_14591,N_14265,N_13841);
nand U14592 (N_14592,N_13863,N_13945);
or U14593 (N_14593,N_14094,N_14182);
or U14594 (N_14594,N_14181,N_13853);
nor U14595 (N_14595,N_14122,N_14140);
or U14596 (N_14596,N_14091,N_14348);
or U14597 (N_14597,N_13877,N_14195);
and U14598 (N_14598,N_14239,N_14084);
nand U14599 (N_14599,N_14388,N_13858);
and U14600 (N_14600,N_14137,N_13953);
nor U14601 (N_14601,N_14235,N_13985);
nor U14602 (N_14602,N_14154,N_14067);
and U14603 (N_14603,N_13995,N_14171);
or U14604 (N_14604,N_14150,N_13879);
nor U14605 (N_14605,N_14390,N_14286);
nor U14606 (N_14606,N_13874,N_14166);
and U14607 (N_14607,N_14304,N_14349);
or U14608 (N_14608,N_14117,N_13909);
and U14609 (N_14609,N_14321,N_13929);
or U14610 (N_14610,N_13801,N_14200);
and U14611 (N_14611,N_13865,N_13894);
or U14612 (N_14612,N_14299,N_13875);
and U14613 (N_14613,N_14114,N_14280);
nand U14614 (N_14614,N_13948,N_14290);
and U14615 (N_14615,N_13864,N_14353);
nor U14616 (N_14616,N_14188,N_14332);
or U14617 (N_14617,N_14234,N_14035);
or U14618 (N_14618,N_14151,N_14038);
and U14619 (N_14619,N_14013,N_14060);
or U14620 (N_14620,N_14197,N_14398);
and U14621 (N_14621,N_13850,N_14351);
nand U14622 (N_14622,N_14222,N_14131);
and U14623 (N_14623,N_13808,N_14387);
or U14624 (N_14624,N_13861,N_14105);
or U14625 (N_14625,N_14316,N_13959);
nor U14626 (N_14626,N_14058,N_13832);
nor U14627 (N_14627,N_14254,N_14386);
nor U14628 (N_14628,N_13963,N_14320);
and U14629 (N_14629,N_14303,N_13842);
or U14630 (N_14630,N_14066,N_13804);
nor U14631 (N_14631,N_14136,N_13940);
nor U14632 (N_14632,N_14382,N_14360);
nor U14633 (N_14633,N_13979,N_14339);
and U14634 (N_14634,N_14377,N_14263);
or U14635 (N_14635,N_13880,N_14378);
or U14636 (N_14636,N_14346,N_13809);
nand U14637 (N_14637,N_14053,N_14101);
nand U14638 (N_14638,N_14223,N_14248);
and U14639 (N_14639,N_14174,N_13819);
and U14640 (N_14640,N_14119,N_14261);
nand U14641 (N_14641,N_13866,N_13812);
or U14642 (N_14642,N_13882,N_14010);
or U14643 (N_14643,N_14052,N_13802);
and U14644 (N_14644,N_14045,N_14005);
and U14645 (N_14645,N_14041,N_13878);
nor U14646 (N_14646,N_14226,N_14229);
nor U14647 (N_14647,N_14255,N_14170);
nor U14648 (N_14648,N_14147,N_14110);
nor U14649 (N_14649,N_14399,N_14326);
xor U14650 (N_14650,N_14164,N_14103);
nand U14651 (N_14651,N_13817,N_14070);
nor U14652 (N_14652,N_14272,N_14334);
nand U14653 (N_14653,N_13908,N_14216);
or U14654 (N_14654,N_14124,N_14162);
nor U14655 (N_14655,N_13884,N_14034);
or U14656 (N_14656,N_13951,N_14340);
nor U14657 (N_14657,N_13892,N_14073);
or U14658 (N_14658,N_14093,N_14394);
and U14659 (N_14659,N_13835,N_13906);
or U14660 (N_14660,N_13905,N_13823);
nor U14661 (N_14661,N_13991,N_14203);
nand U14662 (N_14662,N_13896,N_14036);
nor U14663 (N_14663,N_14090,N_14376);
nor U14664 (N_14664,N_13950,N_14083);
or U14665 (N_14665,N_13886,N_13932);
or U14666 (N_14666,N_14155,N_13969);
and U14667 (N_14667,N_14296,N_14062);
and U14668 (N_14668,N_14350,N_14020);
nand U14669 (N_14669,N_13955,N_14202);
xnor U14670 (N_14670,N_14178,N_14100);
nor U14671 (N_14671,N_14051,N_14371);
xnor U14672 (N_14672,N_13956,N_14009);
nor U14673 (N_14673,N_14130,N_14081);
nor U14674 (N_14674,N_14278,N_14322);
nor U14675 (N_14675,N_13806,N_13818);
or U14676 (N_14676,N_14040,N_14007);
nor U14677 (N_14677,N_14275,N_13871);
nand U14678 (N_14678,N_14074,N_14381);
or U14679 (N_14679,N_14243,N_13889);
nor U14680 (N_14680,N_13935,N_14048);
and U14681 (N_14681,N_14057,N_14308);
nand U14682 (N_14682,N_13977,N_14152);
or U14683 (N_14683,N_14277,N_14246);
nand U14684 (N_14684,N_13914,N_14212);
nand U14685 (N_14685,N_14207,N_14393);
and U14686 (N_14686,N_13847,N_14364);
or U14687 (N_14687,N_14127,N_14118);
or U14688 (N_14688,N_14134,N_13988);
and U14689 (N_14689,N_13838,N_14021);
nand U14690 (N_14690,N_14271,N_13941);
nand U14691 (N_14691,N_14228,N_14297);
and U14692 (N_14692,N_13966,N_13912);
nand U14693 (N_14693,N_13970,N_13895);
or U14694 (N_14694,N_13862,N_14086);
and U14695 (N_14695,N_14138,N_13957);
and U14696 (N_14696,N_13910,N_14180);
nor U14697 (N_14697,N_14123,N_14153);
or U14698 (N_14698,N_14002,N_13937);
nor U14699 (N_14699,N_14059,N_14208);
and U14700 (N_14700,N_14334,N_14015);
or U14701 (N_14701,N_14116,N_14203);
or U14702 (N_14702,N_14234,N_13900);
nand U14703 (N_14703,N_14184,N_14219);
nor U14704 (N_14704,N_13883,N_13895);
or U14705 (N_14705,N_14388,N_13995);
and U14706 (N_14706,N_13994,N_13852);
and U14707 (N_14707,N_14343,N_13928);
xor U14708 (N_14708,N_14027,N_13993);
and U14709 (N_14709,N_14160,N_14065);
or U14710 (N_14710,N_14252,N_14369);
or U14711 (N_14711,N_14157,N_14191);
nor U14712 (N_14712,N_13962,N_13968);
nand U14713 (N_14713,N_14343,N_14085);
and U14714 (N_14714,N_14396,N_14193);
nor U14715 (N_14715,N_14289,N_14087);
nor U14716 (N_14716,N_14049,N_13827);
nor U14717 (N_14717,N_14096,N_14298);
nor U14718 (N_14718,N_14248,N_13979);
xor U14719 (N_14719,N_14145,N_14325);
nor U14720 (N_14720,N_14366,N_13997);
or U14721 (N_14721,N_14276,N_13964);
xnor U14722 (N_14722,N_14139,N_13912);
and U14723 (N_14723,N_13841,N_14294);
nand U14724 (N_14724,N_13978,N_14272);
or U14725 (N_14725,N_14203,N_14234);
or U14726 (N_14726,N_14074,N_14019);
nor U14727 (N_14727,N_14168,N_13910);
and U14728 (N_14728,N_13858,N_14247);
nand U14729 (N_14729,N_14351,N_13887);
and U14730 (N_14730,N_13845,N_13849);
and U14731 (N_14731,N_14205,N_13968);
nand U14732 (N_14732,N_14278,N_14221);
xor U14733 (N_14733,N_14301,N_14092);
nor U14734 (N_14734,N_14274,N_13901);
or U14735 (N_14735,N_14396,N_14352);
xnor U14736 (N_14736,N_14247,N_14235);
nand U14737 (N_14737,N_14075,N_14036);
or U14738 (N_14738,N_14176,N_14294);
and U14739 (N_14739,N_14003,N_14349);
xor U14740 (N_14740,N_14306,N_13876);
nor U14741 (N_14741,N_13861,N_13822);
and U14742 (N_14742,N_14325,N_14067);
xnor U14743 (N_14743,N_14152,N_13869);
or U14744 (N_14744,N_13993,N_14335);
and U14745 (N_14745,N_14129,N_14387);
or U14746 (N_14746,N_13912,N_14101);
nand U14747 (N_14747,N_14041,N_14123);
nand U14748 (N_14748,N_14095,N_14363);
nor U14749 (N_14749,N_14303,N_14160);
and U14750 (N_14750,N_13967,N_13905);
and U14751 (N_14751,N_14284,N_13889);
nor U14752 (N_14752,N_14210,N_13951);
nand U14753 (N_14753,N_14236,N_13904);
nand U14754 (N_14754,N_14189,N_13883);
and U14755 (N_14755,N_14297,N_14337);
nand U14756 (N_14756,N_14198,N_13890);
nand U14757 (N_14757,N_14352,N_14113);
nand U14758 (N_14758,N_14273,N_14098);
nand U14759 (N_14759,N_14227,N_14313);
or U14760 (N_14760,N_13876,N_13830);
or U14761 (N_14761,N_14214,N_13990);
xnor U14762 (N_14762,N_14042,N_13824);
nor U14763 (N_14763,N_14387,N_13893);
and U14764 (N_14764,N_14027,N_14236);
and U14765 (N_14765,N_13903,N_14022);
nor U14766 (N_14766,N_13807,N_14095);
nor U14767 (N_14767,N_14181,N_14137);
nand U14768 (N_14768,N_14115,N_14077);
nor U14769 (N_14769,N_14391,N_14049);
or U14770 (N_14770,N_14054,N_14217);
and U14771 (N_14771,N_14329,N_13974);
or U14772 (N_14772,N_14038,N_13897);
and U14773 (N_14773,N_13896,N_14098);
or U14774 (N_14774,N_14267,N_14168);
nand U14775 (N_14775,N_14121,N_14099);
nor U14776 (N_14776,N_13816,N_14256);
or U14777 (N_14777,N_14186,N_13869);
nand U14778 (N_14778,N_14132,N_14300);
nor U14779 (N_14779,N_13970,N_14003);
nor U14780 (N_14780,N_14152,N_14287);
nor U14781 (N_14781,N_14101,N_14315);
nand U14782 (N_14782,N_13948,N_13933);
or U14783 (N_14783,N_14323,N_13884);
nand U14784 (N_14784,N_13977,N_14348);
nor U14785 (N_14785,N_14194,N_14112);
nor U14786 (N_14786,N_14236,N_14084);
nand U14787 (N_14787,N_14270,N_14340);
nand U14788 (N_14788,N_13966,N_14216);
and U14789 (N_14789,N_14130,N_14258);
nand U14790 (N_14790,N_14315,N_13934);
nand U14791 (N_14791,N_13895,N_14064);
and U14792 (N_14792,N_14087,N_14338);
xnor U14793 (N_14793,N_13819,N_14249);
nand U14794 (N_14794,N_14192,N_14352);
or U14795 (N_14795,N_14369,N_13901);
nand U14796 (N_14796,N_14042,N_14135);
and U14797 (N_14797,N_14261,N_13949);
and U14798 (N_14798,N_13853,N_14162);
or U14799 (N_14799,N_14208,N_14175);
or U14800 (N_14800,N_14253,N_14162);
nor U14801 (N_14801,N_14330,N_14105);
nand U14802 (N_14802,N_14393,N_13896);
or U14803 (N_14803,N_13877,N_13855);
nor U14804 (N_14804,N_13997,N_13822);
and U14805 (N_14805,N_14092,N_13906);
and U14806 (N_14806,N_14153,N_14392);
and U14807 (N_14807,N_14020,N_14320);
and U14808 (N_14808,N_14331,N_14012);
and U14809 (N_14809,N_14182,N_13820);
nand U14810 (N_14810,N_14354,N_14271);
and U14811 (N_14811,N_14170,N_13840);
and U14812 (N_14812,N_14026,N_14337);
nor U14813 (N_14813,N_14153,N_14255);
and U14814 (N_14814,N_14039,N_13823);
and U14815 (N_14815,N_14214,N_14324);
or U14816 (N_14816,N_14366,N_14344);
and U14817 (N_14817,N_14391,N_14362);
and U14818 (N_14818,N_13883,N_14129);
nand U14819 (N_14819,N_14270,N_13901);
and U14820 (N_14820,N_13855,N_13817);
or U14821 (N_14821,N_13867,N_13823);
and U14822 (N_14822,N_14258,N_13853);
or U14823 (N_14823,N_13975,N_14353);
nor U14824 (N_14824,N_14102,N_14097);
and U14825 (N_14825,N_13937,N_14337);
and U14826 (N_14826,N_14185,N_13846);
nand U14827 (N_14827,N_14096,N_14132);
and U14828 (N_14828,N_14213,N_13950);
nand U14829 (N_14829,N_13963,N_14091);
nand U14830 (N_14830,N_13918,N_13883);
or U14831 (N_14831,N_14384,N_13897);
nand U14832 (N_14832,N_13976,N_14028);
or U14833 (N_14833,N_14014,N_13814);
nand U14834 (N_14834,N_13821,N_13990);
and U14835 (N_14835,N_13991,N_14081);
and U14836 (N_14836,N_14293,N_14237);
nor U14837 (N_14837,N_14370,N_14042);
and U14838 (N_14838,N_14232,N_13887);
and U14839 (N_14839,N_14342,N_14279);
or U14840 (N_14840,N_13911,N_13915);
nand U14841 (N_14841,N_14288,N_14240);
nand U14842 (N_14842,N_14339,N_14001);
nand U14843 (N_14843,N_13812,N_14150);
nor U14844 (N_14844,N_13915,N_13883);
nor U14845 (N_14845,N_13933,N_14260);
and U14846 (N_14846,N_13947,N_13877);
and U14847 (N_14847,N_14357,N_14349);
nor U14848 (N_14848,N_13832,N_14061);
nor U14849 (N_14849,N_14110,N_13824);
nand U14850 (N_14850,N_14179,N_14055);
nor U14851 (N_14851,N_14121,N_13902);
nand U14852 (N_14852,N_14173,N_13917);
and U14853 (N_14853,N_14214,N_13978);
nand U14854 (N_14854,N_13940,N_13918);
nand U14855 (N_14855,N_13922,N_14099);
nor U14856 (N_14856,N_13857,N_13864);
or U14857 (N_14857,N_14011,N_13840);
nor U14858 (N_14858,N_14122,N_14039);
or U14859 (N_14859,N_14188,N_14305);
nor U14860 (N_14860,N_14111,N_14039);
or U14861 (N_14861,N_13953,N_14146);
nand U14862 (N_14862,N_13880,N_14225);
or U14863 (N_14863,N_13916,N_14096);
and U14864 (N_14864,N_14247,N_14060);
and U14865 (N_14865,N_14248,N_13949);
and U14866 (N_14866,N_13923,N_14019);
nor U14867 (N_14867,N_14396,N_13856);
or U14868 (N_14868,N_14214,N_14046);
nand U14869 (N_14869,N_14299,N_14088);
nor U14870 (N_14870,N_13963,N_14162);
nand U14871 (N_14871,N_14182,N_14301);
nor U14872 (N_14872,N_14312,N_14278);
and U14873 (N_14873,N_14016,N_13851);
and U14874 (N_14874,N_13852,N_14348);
nor U14875 (N_14875,N_13804,N_13901);
and U14876 (N_14876,N_14185,N_14289);
or U14877 (N_14877,N_13937,N_13852);
nand U14878 (N_14878,N_14173,N_14310);
nand U14879 (N_14879,N_14065,N_13918);
and U14880 (N_14880,N_14200,N_13923);
xor U14881 (N_14881,N_13968,N_14108);
and U14882 (N_14882,N_14308,N_14023);
nand U14883 (N_14883,N_14187,N_13873);
or U14884 (N_14884,N_13979,N_14018);
nand U14885 (N_14885,N_14201,N_14325);
and U14886 (N_14886,N_14071,N_14340);
and U14887 (N_14887,N_14210,N_13831);
nor U14888 (N_14888,N_14139,N_13876);
or U14889 (N_14889,N_14224,N_13922);
and U14890 (N_14890,N_13853,N_14334);
nand U14891 (N_14891,N_13979,N_14399);
nor U14892 (N_14892,N_14340,N_14272);
and U14893 (N_14893,N_13981,N_14082);
or U14894 (N_14894,N_14060,N_14053);
nor U14895 (N_14895,N_13854,N_13834);
or U14896 (N_14896,N_13889,N_14030);
and U14897 (N_14897,N_14163,N_14280);
nor U14898 (N_14898,N_14372,N_14017);
or U14899 (N_14899,N_14084,N_14076);
and U14900 (N_14900,N_13983,N_14192);
nand U14901 (N_14901,N_14001,N_14347);
nor U14902 (N_14902,N_14045,N_13881);
nand U14903 (N_14903,N_14271,N_14172);
or U14904 (N_14904,N_13993,N_14129);
and U14905 (N_14905,N_14259,N_14020);
nand U14906 (N_14906,N_14205,N_14051);
or U14907 (N_14907,N_14327,N_13978);
nand U14908 (N_14908,N_14205,N_14109);
or U14909 (N_14909,N_13978,N_14235);
and U14910 (N_14910,N_13815,N_14273);
or U14911 (N_14911,N_14146,N_14051);
nor U14912 (N_14912,N_13902,N_14253);
nor U14913 (N_14913,N_14078,N_13808);
and U14914 (N_14914,N_14302,N_13869);
nor U14915 (N_14915,N_14366,N_14353);
and U14916 (N_14916,N_14249,N_14230);
nor U14917 (N_14917,N_14031,N_13851);
nand U14918 (N_14918,N_14160,N_14109);
and U14919 (N_14919,N_14211,N_14003);
or U14920 (N_14920,N_14298,N_13940);
and U14921 (N_14921,N_14210,N_13935);
nor U14922 (N_14922,N_14047,N_14220);
nor U14923 (N_14923,N_14055,N_14106);
or U14924 (N_14924,N_13893,N_13892);
and U14925 (N_14925,N_13960,N_14137);
nor U14926 (N_14926,N_13928,N_14075);
or U14927 (N_14927,N_14071,N_13844);
nand U14928 (N_14928,N_14106,N_13917);
or U14929 (N_14929,N_14070,N_13835);
or U14930 (N_14930,N_13895,N_14395);
or U14931 (N_14931,N_14394,N_14043);
nor U14932 (N_14932,N_14148,N_14278);
or U14933 (N_14933,N_13907,N_14302);
and U14934 (N_14934,N_13941,N_14137);
and U14935 (N_14935,N_14176,N_14355);
nand U14936 (N_14936,N_14387,N_13821);
nand U14937 (N_14937,N_13825,N_14273);
or U14938 (N_14938,N_14063,N_14154);
nand U14939 (N_14939,N_13950,N_13807);
and U14940 (N_14940,N_14094,N_13919);
nand U14941 (N_14941,N_14039,N_14245);
and U14942 (N_14942,N_14392,N_13863);
nor U14943 (N_14943,N_14188,N_13998);
nor U14944 (N_14944,N_14161,N_14290);
and U14945 (N_14945,N_13949,N_14021);
and U14946 (N_14946,N_14345,N_14244);
nor U14947 (N_14947,N_14178,N_14101);
and U14948 (N_14948,N_14050,N_14332);
and U14949 (N_14949,N_14111,N_13808);
nand U14950 (N_14950,N_13852,N_13897);
nor U14951 (N_14951,N_13909,N_14348);
nor U14952 (N_14952,N_14154,N_14198);
nand U14953 (N_14953,N_13930,N_14366);
and U14954 (N_14954,N_13870,N_13960);
and U14955 (N_14955,N_13851,N_14371);
nand U14956 (N_14956,N_14129,N_13973);
nor U14957 (N_14957,N_14046,N_13805);
nand U14958 (N_14958,N_14103,N_14305);
nor U14959 (N_14959,N_13867,N_14174);
nor U14960 (N_14960,N_13969,N_14183);
xnor U14961 (N_14961,N_13966,N_14284);
and U14962 (N_14962,N_13954,N_14087);
nor U14963 (N_14963,N_14144,N_14262);
nor U14964 (N_14964,N_14373,N_14295);
nand U14965 (N_14965,N_14000,N_14066);
and U14966 (N_14966,N_13902,N_13958);
and U14967 (N_14967,N_13923,N_13821);
nand U14968 (N_14968,N_14176,N_13891);
xnor U14969 (N_14969,N_13803,N_14311);
nand U14970 (N_14970,N_14098,N_14077);
nand U14971 (N_14971,N_14126,N_13992);
or U14972 (N_14972,N_14352,N_14152);
or U14973 (N_14973,N_14199,N_14296);
or U14974 (N_14974,N_14284,N_13891);
nor U14975 (N_14975,N_14113,N_14368);
nand U14976 (N_14976,N_14240,N_14118);
or U14977 (N_14977,N_14393,N_14268);
or U14978 (N_14978,N_14009,N_14158);
and U14979 (N_14979,N_14322,N_14182);
or U14980 (N_14980,N_14262,N_13966);
nand U14981 (N_14981,N_13942,N_14350);
or U14982 (N_14982,N_13817,N_14379);
and U14983 (N_14983,N_14026,N_13820);
and U14984 (N_14984,N_14260,N_13975);
nand U14985 (N_14985,N_14060,N_13818);
or U14986 (N_14986,N_13811,N_14353);
and U14987 (N_14987,N_13872,N_13835);
or U14988 (N_14988,N_13879,N_13871);
and U14989 (N_14989,N_13995,N_14014);
nand U14990 (N_14990,N_14092,N_14091);
or U14991 (N_14991,N_13961,N_14279);
nand U14992 (N_14992,N_14372,N_14337);
nand U14993 (N_14993,N_14112,N_14215);
or U14994 (N_14994,N_14303,N_14033);
nand U14995 (N_14995,N_14249,N_13817);
and U14996 (N_14996,N_14122,N_13949);
nor U14997 (N_14997,N_13992,N_14169);
nand U14998 (N_14998,N_14077,N_14277);
or U14999 (N_14999,N_14238,N_14035);
and U15000 (N_15000,N_14737,N_14410);
and U15001 (N_15001,N_14450,N_14746);
or U15002 (N_15002,N_14752,N_14472);
or U15003 (N_15003,N_14872,N_14400);
and U15004 (N_15004,N_14840,N_14757);
nor U15005 (N_15005,N_14877,N_14862);
and U15006 (N_15006,N_14914,N_14692);
nor U15007 (N_15007,N_14618,N_14792);
nor U15008 (N_15008,N_14694,N_14874);
nand U15009 (N_15009,N_14656,N_14449);
or U15010 (N_15010,N_14731,N_14582);
nand U15011 (N_15011,N_14493,N_14622);
nor U15012 (N_15012,N_14721,N_14961);
nand U15013 (N_15013,N_14853,N_14465);
nor U15014 (N_15014,N_14575,N_14913);
and U15015 (N_15015,N_14445,N_14697);
and U15016 (N_15016,N_14654,N_14875);
or U15017 (N_15017,N_14548,N_14490);
and U15018 (N_15018,N_14911,N_14606);
nor U15019 (N_15019,N_14866,N_14933);
nor U15020 (N_15020,N_14550,N_14458);
or U15021 (N_15021,N_14940,N_14412);
or U15022 (N_15022,N_14748,N_14659);
nand U15023 (N_15023,N_14819,N_14507);
nor U15024 (N_15024,N_14971,N_14716);
or U15025 (N_15025,N_14763,N_14451);
or U15026 (N_15026,N_14597,N_14546);
and U15027 (N_15027,N_14639,N_14588);
and U15028 (N_15028,N_14753,N_14585);
nand U15029 (N_15029,N_14952,N_14577);
nor U15030 (N_15030,N_14584,N_14718);
or U15031 (N_15031,N_14554,N_14568);
nor U15032 (N_15032,N_14719,N_14836);
and U15033 (N_15033,N_14565,N_14802);
nand U15034 (N_15034,N_14631,N_14453);
or U15035 (N_15035,N_14759,N_14591);
nand U15036 (N_15036,N_14513,N_14993);
nor U15037 (N_15037,N_14804,N_14648);
or U15038 (N_15038,N_14436,N_14809);
nor U15039 (N_15039,N_14534,N_14803);
or U15040 (N_15040,N_14770,N_14953);
and U15041 (N_15041,N_14972,N_14402);
nor U15042 (N_15042,N_14881,N_14724);
or U15043 (N_15043,N_14523,N_14482);
or U15044 (N_15044,N_14477,N_14787);
and U15045 (N_15045,N_14766,N_14690);
or U15046 (N_15046,N_14587,N_14830);
or U15047 (N_15047,N_14901,N_14406);
and U15048 (N_15048,N_14794,N_14838);
nor U15049 (N_15049,N_14567,N_14852);
and U15050 (N_15050,N_14888,N_14774);
nand U15051 (N_15051,N_14646,N_14668);
nor U15052 (N_15052,N_14825,N_14667);
and U15053 (N_15053,N_14779,N_14791);
nor U15054 (N_15054,N_14435,N_14761);
nand U15055 (N_15055,N_14665,N_14943);
xnor U15056 (N_15056,N_14706,N_14636);
or U15057 (N_15057,N_14906,N_14886);
and U15058 (N_15058,N_14421,N_14921);
and U15059 (N_15059,N_14885,N_14745);
nor U15060 (N_15060,N_14832,N_14891);
nand U15061 (N_15061,N_14569,N_14851);
and U15062 (N_15062,N_14843,N_14768);
or U15063 (N_15063,N_14492,N_14564);
and U15064 (N_15064,N_14725,N_14617);
and U15065 (N_15065,N_14863,N_14699);
nor U15066 (N_15066,N_14858,N_14531);
and U15067 (N_15067,N_14896,N_14789);
nor U15068 (N_15068,N_14844,N_14994);
or U15069 (N_15069,N_14711,N_14658);
or U15070 (N_15070,N_14855,N_14430);
or U15071 (N_15071,N_14603,N_14570);
and U15072 (N_15072,N_14540,N_14965);
nor U15073 (N_15073,N_14799,N_14643);
or U15074 (N_15074,N_14894,N_14583);
or U15075 (N_15075,N_14882,N_14714);
nor U15076 (N_15076,N_14439,N_14762);
xnor U15077 (N_15077,N_14992,N_14645);
and U15078 (N_15078,N_14483,N_14728);
nand U15079 (N_15079,N_14635,N_14563);
nor U15080 (N_15080,N_14782,N_14826);
nor U15081 (N_15081,N_14424,N_14558);
and U15082 (N_15082,N_14519,N_14625);
and U15083 (N_15083,N_14726,N_14754);
or U15084 (N_15084,N_14898,N_14544);
nor U15085 (N_15085,N_14817,N_14590);
or U15086 (N_15086,N_14937,N_14468);
or U15087 (N_15087,N_14765,N_14604);
or U15088 (N_15088,N_14974,N_14626);
or U15089 (N_15089,N_14509,N_14890);
and U15090 (N_15090,N_14664,N_14771);
nand U15091 (N_15091,N_14671,N_14413);
nand U15092 (N_15092,N_14627,N_14904);
or U15093 (N_15093,N_14884,N_14437);
nor U15094 (N_15094,N_14600,N_14557);
nand U15095 (N_15095,N_14497,N_14772);
nand U15096 (N_15096,N_14644,N_14938);
nor U15097 (N_15097,N_14611,N_14735);
nand U15098 (N_15098,N_14729,N_14685);
and U15099 (N_15099,N_14788,N_14983);
nand U15100 (N_15100,N_14653,N_14623);
and U15101 (N_15101,N_14580,N_14592);
nand U15102 (N_15102,N_14823,N_14871);
or U15103 (N_15103,N_14680,N_14813);
nand U15104 (N_15104,N_14669,N_14542);
nand U15105 (N_15105,N_14463,N_14876);
or U15106 (N_15106,N_14910,N_14526);
xnor U15107 (N_15107,N_14741,N_14756);
nor U15108 (N_15108,N_14598,N_14968);
or U15109 (N_15109,N_14525,N_14883);
nor U15110 (N_15110,N_14522,N_14801);
nor U15111 (N_15111,N_14417,N_14909);
nand U15112 (N_15112,N_14740,N_14814);
nand U15113 (N_15113,N_14977,N_14764);
or U15114 (N_15114,N_14723,N_14491);
nor U15115 (N_15115,N_14957,N_14734);
and U15116 (N_15116,N_14432,N_14790);
and U15117 (N_15117,N_14695,N_14988);
nand U15118 (N_15118,N_14552,N_14868);
nor U15119 (N_15119,N_14709,N_14828);
and U15120 (N_15120,N_14556,N_14796);
and U15121 (N_15121,N_14747,N_14429);
and U15122 (N_15122,N_14727,N_14925);
or U15123 (N_15123,N_14446,N_14677);
and U15124 (N_15124,N_14707,N_14902);
nand U15125 (N_15125,N_14459,N_14989);
nor U15126 (N_15126,N_14879,N_14551);
nor U15127 (N_15127,N_14918,N_14601);
nand U15128 (N_15128,N_14481,N_14433);
nor U15129 (N_15129,N_14613,N_14831);
and U15130 (N_15130,N_14688,N_14423);
nand U15131 (N_15131,N_14608,N_14889);
or U15132 (N_15132,N_14924,N_14524);
or U15133 (N_15133,N_14466,N_14899);
nand U15134 (N_15134,N_14793,N_14660);
nand U15135 (N_15135,N_14955,N_14521);
or U15136 (N_15136,N_14930,N_14810);
nand U15137 (N_15137,N_14683,N_14928);
or U15138 (N_15138,N_14454,N_14506);
or U15139 (N_15139,N_14640,N_14543);
nand U15140 (N_15140,N_14441,N_14777);
nor U15141 (N_15141,N_14573,N_14900);
nand U15142 (N_15142,N_14649,N_14457);
nor U15143 (N_15143,N_14686,N_14508);
nand U15144 (N_15144,N_14405,N_14530);
or U15145 (N_15145,N_14775,N_14945);
nand U15146 (N_15146,N_14923,N_14673);
or U15147 (N_15147,N_14738,N_14538);
and U15148 (N_15148,N_14448,N_14712);
or U15149 (N_15149,N_14970,N_14839);
and U15150 (N_15150,N_14474,N_14783);
nor U15151 (N_15151,N_14517,N_14431);
or U15152 (N_15152,N_14541,N_14687);
nor U15153 (N_15153,N_14999,N_14998);
and U15154 (N_15154,N_14566,N_14818);
and U15155 (N_15155,N_14964,N_14837);
and U15156 (N_15156,N_14946,N_14520);
nor U15157 (N_15157,N_14705,N_14717);
nor U15158 (N_15158,N_14722,N_14462);
nand U15159 (N_15159,N_14750,N_14786);
nor U15160 (N_15160,N_14773,N_14966);
and U15161 (N_15161,N_14976,N_14661);
nand U15162 (N_15162,N_14401,N_14652);
nor U15163 (N_15163,N_14931,N_14848);
or U15164 (N_15164,N_14984,N_14869);
nand U15165 (N_15165,N_14942,N_14720);
nor U15166 (N_15166,N_14847,N_14471);
and U15167 (N_15167,N_14878,N_14950);
nor U15168 (N_15168,N_14973,N_14807);
and U15169 (N_15169,N_14963,N_14939);
nor U15170 (N_15170,N_14473,N_14895);
nand U15171 (N_15171,N_14978,N_14675);
nand U15172 (N_15172,N_14919,N_14547);
or U15173 (N_15173,N_14982,N_14981);
or U15174 (N_15174,N_14561,N_14452);
nand U15175 (N_15175,N_14461,N_14678);
or U15176 (N_15176,N_14571,N_14553);
nor U15177 (N_15177,N_14438,N_14751);
and U15178 (N_15178,N_14713,N_14480);
nor U15179 (N_15179,N_14867,N_14487);
nand U15180 (N_15180,N_14785,N_14489);
nor U15181 (N_15181,N_14760,N_14778);
or U15182 (N_15182,N_14532,N_14641);
nand U15183 (N_15183,N_14932,N_14529);
and U15184 (N_15184,N_14927,N_14574);
xor U15185 (N_15185,N_14478,N_14859);
nand U15186 (N_15186,N_14861,N_14975);
nor U15187 (N_15187,N_14510,N_14505);
or U15188 (N_15188,N_14479,N_14776);
nor U15189 (N_15189,N_14516,N_14536);
or U15190 (N_15190,N_14502,N_14800);
nand U15191 (N_15191,N_14986,N_14833);
nor U15192 (N_15192,N_14907,N_14846);
or U15193 (N_15193,N_14467,N_14655);
nor U15194 (N_15194,N_14504,N_14624);
nand U15195 (N_15195,N_14460,N_14829);
and U15196 (N_15196,N_14958,N_14620);
or U15197 (N_15197,N_14593,N_14893);
and U15198 (N_15198,N_14944,N_14684);
nand U15199 (N_15199,N_14954,N_14609);
or U15200 (N_15200,N_14812,N_14610);
and U15201 (N_15201,N_14411,N_14769);
and U15202 (N_15202,N_14865,N_14811);
or U15203 (N_15203,N_14404,N_14647);
nor U15204 (N_15204,N_14651,N_14630);
nand U15205 (N_15205,N_14420,N_14442);
and U15206 (N_15206,N_14632,N_14702);
or U15207 (N_15207,N_14425,N_14710);
nor U15208 (N_15208,N_14579,N_14860);
or U15209 (N_15209,N_14498,N_14864);
or U15210 (N_15210,N_14595,N_14511);
and U15211 (N_15211,N_14758,N_14755);
nor U15212 (N_15212,N_14730,N_14698);
and U15213 (N_15213,N_14960,N_14485);
nor U15214 (N_15214,N_14681,N_14503);
xnor U15215 (N_15215,N_14670,N_14555);
nor U15216 (N_15216,N_14934,N_14701);
and U15217 (N_15217,N_14842,N_14619);
nand U15218 (N_15218,N_14912,N_14434);
nor U15219 (N_15219,N_14821,N_14739);
xnor U15220 (N_15220,N_14951,N_14815);
and U15221 (N_15221,N_14822,N_14841);
and U15222 (N_15222,N_14935,N_14880);
and U15223 (N_15223,N_14419,N_14850);
or U15224 (N_15224,N_14736,N_14559);
xnor U15225 (N_15225,N_14537,N_14615);
and U15226 (N_15226,N_14500,N_14476);
nand U15227 (N_15227,N_14805,N_14936);
or U15228 (N_15228,N_14605,N_14674);
and U15229 (N_15229,N_14696,N_14518);
nand U15230 (N_15230,N_14856,N_14447);
and U15231 (N_15231,N_14545,N_14501);
nand U15232 (N_15232,N_14979,N_14469);
or U15233 (N_15233,N_14576,N_14409);
and U15234 (N_15234,N_14629,N_14455);
and U15235 (N_15235,N_14854,N_14486);
and U15236 (N_15236,N_14422,N_14456);
nor U15237 (N_15237,N_14996,N_14515);
and U15238 (N_15238,N_14512,N_14638);
nand U15239 (N_15239,N_14589,N_14637);
nand U15240 (N_15240,N_14427,N_14594);
nand U15241 (N_15241,N_14549,N_14835);
nand U15242 (N_15242,N_14693,N_14672);
or U15243 (N_15243,N_14887,N_14873);
and U15244 (N_15244,N_14586,N_14897);
or U15245 (N_15245,N_14744,N_14599);
and U15246 (N_15246,N_14663,N_14484);
nor U15247 (N_15247,N_14602,N_14784);
and U15248 (N_15248,N_14691,N_14806);
nor U15249 (N_15249,N_14642,N_14428);
nor U15250 (N_15250,N_14689,N_14915);
nor U15251 (N_15251,N_14824,N_14715);
and U15252 (N_15252,N_14908,N_14780);
nand U15253 (N_15253,N_14849,N_14742);
nand U15254 (N_15254,N_14949,N_14816);
nand U15255 (N_15255,N_14464,N_14581);
nor U15256 (N_15256,N_14708,N_14616);
and U15257 (N_15257,N_14967,N_14941);
nor U15258 (N_15258,N_14560,N_14948);
and U15259 (N_15259,N_14857,N_14767);
and U15260 (N_15260,N_14990,N_14403);
nand U15261 (N_15261,N_14920,N_14749);
nand U15262 (N_15262,N_14415,N_14916);
and U15263 (N_15263,N_14682,N_14845);
or U15264 (N_15264,N_14798,N_14987);
nand U15265 (N_15265,N_14470,N_14892);
nand U15266 (N_15266,N_14488,N_14612);
nand U15267 (N_15267,N_14418,N_14596);
or U15268 (N_15268,N_14650,N_14494);
or U15269 (N_15269,N_14607,N_14827);
xnor U15270 (N_15270,N_14743,N_14917);
nand U15271 (N_15271,N_14980,N_14533);
or U15272 (N_15272,N_14408,N_14499);
or U15273 (N_15273,N_14676,N_14926);
nor U15274 (N_15274,N_14732,N_14407);
and U15275 (N_15275,N_14704,N_14527);
or U15276 (N_15276,N_14795,N_14562);
nor U15277 (N_15277,N_14416,N_14634);
nor U15278 (N_15278,N_14820,N_14947);
or U15279 (N_15279,N_14679,N_14614);
or U15280 (N_15280,N_14905,N_14444);
and U15281 (N_15281,N_14572,N_14539);
nor U15282 (N_15282,N_14808,N_14703);
and U15283 (N_15283,N_14903,N_14991);
or U15284 (N_15284,N_14956,N_14959);
nor U15285 (N_15285,N_14578,N_14514);
nor U15286 (N_15286,N_14985,N_14700);
nor U15287 (N_15287,N_14662,N_14628);
nor U15288 (N_15288,N_14995,N_14922);
nand U15289 (N_15289,N_14969,N_14997);
or U15290 (N_15290,N_14929,N_14496);
or U15291 (N_15291,N_14440,N_14621);
nor U15292 (N_15292,N_14475,N_14426);
and U15293 (N_15293,N_14443,N_14528);
or U15294 (N_15294,N_14495,N_14535);
nor U15295 (N_15295,N_14870,N_14834);
and U15296 (N_15296,N_14414,N_14962);
and U15297 (N_15297,N_14797,N_14781);
and U15298 (N_15298,N_14666,N_14657);
nor U15299 (N_15299,N_14633,N_14733);
nand U15300 (N_15300,N_14785,N_14788);
or U15301 (N_15301,N_14926,N_14409);
and U15302 (N_15302,N_14696,N_14712);
nand U15303 (N_15303,N_14960,N_14610);
nor U15304 (N_15304,N_14604,N_14416);
nor U15305 (N_15305,N_14421,N_14730);
and U15306 (N_15306,N_14658,N_14956);
nor U15307 (N_15307,N_14914,N_14729);
nand U15308 (N_15308,N_14778,N_14794);
and U15309 (N_15309,N_14466,N_14943);
and U15310 (N_15310,N_14952,N_14685);
nand U15311 (N_15311,N_14446,N_14459);
nand U15312 (N_15312,N_14589,N_14832);
nand U15313 (N_15313,N_14904,N_14711);
nand U15314 (N_15314,N_14944,N_14809);
nor U15315 (N_15315,N_14736,N_14615);
nor U15316 (N_15316,N_14837,N_14528);
and U15317 (N_15317,N_14554,N_14644);
and U15318 (N_15318,N_14638,N_14457);
and U15319 (N_15319,N_14901,N_14782);
or U15320 (N_15320,N_14772,N_14749);
and U15321 (N_15321,N_14553,N_14868);
and U15322 (N_15322,N_14555,N_14499);
and U15323 (N_15323,N_14877,N_14509);
nand U15324 (N_15324,N_14901,N_14445);
nand U15325 (N_15325,N_14401,N_14703);
nor U15326 (N_15326,N_14753,N_14544);
nand U15327 (N_15327,N_14862,N_14727);
nor U15328 (N_15328,N_14498,N_14963);
and U15329 (N_15329,N_14869,N_14996);
and U15330 (N_15330,N_14413,N_14546);
nand U15331 (N_15331,N_14457,N_14781);
nand U15332 (N_15332,N_14816,N_14941);
nor U15333 (N_15333,N_14924,N_14977);
nand U15334 (N_15334,N_14515,N_14750);
or U15335 (N_15335,N_14912,N_14932);
or U15336 (N_15336,N_14910,N_14632);
nor U15337 (N_15337,N_14697,N_14783);
and U15338 (N_15338,N_14799,N_14936);
nor U15339 (N_15339,N_14950,N_14723);
nor U15340 (N_15340,N_14536,N_14808);
and U15341 (N_15341,N_14455,N_14413);
and U15342 (N_15342,N_14980,N_14589);
xnor U15343 (N_15343,N_14986,N_14849);
nor U15344 (N_15344,N_14734,N_14451);
and U15345 (N_15345,N_14710,N_14889);
nor U15346 (N_15346,N_14676,N_14478);
nand U15347 (N_15347,N_14470,N_14871);
nor U15348 (N_15348,N_14440,N_14686);
nand U15349 (N_15349,N_14798,N_14874);
or U15350 (N_15350,N_14740,N_14719);
or U15351 (N_15351,N_14709,N_14449);
and U15352 (N_15352,N_14712,N_14827);
nand U15353 (N_15353,N_14804,N_14570);
and U15354 (N_15354,N_14442,N_14872);
nand U15355 (N_15355,N_14577,N_14924);
nor U15356 (N_15356,N_14891,N_14834);
nand U15357 (N_15357,N_14780,N_14810);
and U15358 (N_15358,N_14485,N_14820);
and U15359 (N_15359,N_14974,N_14722);
and U15360 (N_15360,N_14509,N_14842);
or U15361 (N_15361,N_14455,N_14784);
and U15362 (N_15362,N_14477,N_14517);
and U15363 (N_15363,N_14648,N_14915);
and U15364 (N_15364,N_14683,N_14572);
xnor U15365 (N_15365,N_14952,N_14509);
or U15366 (N_15366,N_14485,N_14471);
nor U15367 (N_15367,N_14666,N_14670);
or U15368 (N_15368,N_14581,N_14625);
or U15369 (N_15369,N_14962,N_14807);
nor U15370 (N_15370,N_14696,N_14795);
nor U15371 (N_15371,N_14563,N_14433);
nand U15372 (N_15372,N_14622,N_14987);
nor U15373 (N_15373,N_14670,N_14776);
and U15374 (N_15374,N_14993,N_14999);
or U15375 (N_15375,N_14428,N_14572);
nand U15376 (N_15376,N_14933,N_14782);
and U15377 (N_15377,N_14518,N_14967);
nor U15378 (N_15378,N_14963,N_14793);
or U15379 (N_15379,N_14486,N_14877);
or U15380 (N_15380,N_14897,N_14813);
nand U15381 (N_15381,N_14507,N_14603);
xor U15382 (N_15382,N_14881,N_14654);
nand U15383 (N_15383,N_14888,N_14511);
or U15384 (N_15384,N_14826,N_14940);
xnor U15385 (N_15385,N_14770,N_14927);
nor U15386 (N_15386,N_14555,N_14874);
nor U15387 (N_15387,N_14414,N_14521);
nand U15388 (N_15388,N_14964,N_14657);
nor U15389 (N_15389,N_14651,N_14513);
or U15390 (N_15390,N_14540,N_14603);
and U15391 (N_15391,N_14402,N_14406);
and U15392 (N_15392,N_14804,N_14501);
nand U15393 (N_15393,N_14725,N_14428);
nand U15394 (N_15394,N_14688,N_14526);
or U15395 (N_15395,N_14790,N_14993);
xnor U15396 (N_15396,N_14644,N_14989);
and U15397 (N_15397,N_14470,N_14653);
nand U15398 (N_15398,N_14951,N_14408);
and U15399 (N_15399,N_14606,N_14705);
or U15400 (N_15400,N_14881,N_14681);
nand U15401 (N_15401,N_14483,N_14844);
nand U15402 (N_15402,N_14875,N_14643);
xor U15403 (N_15403,N_14419,N_14910);
or U15404 (N_15404,N_14826,N_14653);
and U15405 (N_15405,N_14501,N_14754);
nand U15406 (N_15406,N_14621,N_14618);
nor U15407 (N_15407,N_14685,N_14842);
and U15408 (N_15408,N_14501,N_14543);
nand U15409 (N_15409,N_14472,N_14883);
nor U15410 (N_15410,N_14566,N_14497);
nor U15411 (N_15411,N_14465,N_14448);
or U15412 (N_15412,N_14827,N_14421);
nor U15413 (N_15413,N_14508,N_14955);
nor U15414 (N_15414,N_14657,N_14840);
nand U15415 (N_15415,N_14601,N_14676);
or U15416 (N_15416,N_14717,N_14435);
xnor U15417 (N_15417,N_14513,N_14822);
nor U15418 (N_15418,N_14595,N_14663);
and U15419 (N_15419,N_14919,N_14587);
and U15420 (N_15420,N_14784,N_14521);
nor U15421 (N_15421,N_14569,N_14626);
nand U15422 (N_15422,N_14669,N_14889);
or U15423 (N_15423,N_14425,N_14727);
or U15424 (N_15424,N_14595,N_14584);
nor U15425 (N_15425,N_14547,N_14715);
and U15426 (N_15426,N_14555,N_14572);
or U15427 (N_15427,N_14521,N_14665);
or U15428 (N_15428,N_14692,N_14591);
and U15429 (N_15429,N_14849,N_14672);
nand U15430 (N_15430,N_14663,N_14413);
or U15431 (N_15431,N_14839,N_14683);
nor U15432 (N_15432,N_14910,N_14952);
or U15433 (N_15433,N_14899,N_14578);
or U15434 (N_15434,N_14805,N_14498);
and U15435 (N_15435,N_14822,N_14861);
nor U15436 (N_15436,N_14988,N_14667);
or U15437 (N_15437,N_14871,N_14627);
and U15438 (N_15438,N_14492,N_14770);
and U15439 (N_15439,N_14480,N_14543);
nand U15440 (N_15440,N_14676,N_14858);
or U15441 (N_15441,N_14700,N_14913);
nor U15442 (N_15442,N_14401,N_14552);
xnor U15443 (N_15443,N_14422,N_14408);
or U15444 (N_15444,N_14963,N_14450);
nor U15445 (N_15445,N_14470,N_14679);
and U15446 (N_15446,N_14522,N_14844);
nand U15447 (N_15447,N_14444,N_14870);
nand U15448 (N_15448,N_14856,N_14759);
nand U15449 (N_15449,N_14912,N_14923);
nor U15450 (N_15450,N_14556,N_14449);
and U15451 (N_15451,N_14681,N_14994);
nand U15452 (N_15452,N_14656,N_14834);
and U15453 (N_15453,N_14703,N_14507);
nand U15454 (N_15454,N_14484,N_14733);
nor U15455 (N_15455,N_14506,N_14882);
nor U15456 (N_15456,N_14838,N_14520);
and U15457 (N_15457,N_14411,N_14816);
nor U15458 (N_15458,N_14432,N_14494);
or U15459 (N_15459,N_14432,N_14970);
nand U15460 (N_15460,N_14857,N_14542);
or U15461 (N_15461,N_14450,N_14900);
nor U15462 (N_15462,N_14640,N_14837);
nand U15463 (N_15463,N_14925,N_14956);
nand U15464 (N_15464,N_14692,N_14701);
and U15465 (N_15465,N_14957,N_14431);
or U15466 (N_15466,N_14468,N_14491);
nand U15467 (N_15467,N_14772,N_14884);
and U15468 (N_15468,N_14455,N_14484);
nor U15469 (N_15469,N_14609,N_14798);
nand U15470 (N_15470,N_14898,N_14749);
or U15471 (N_15471,N_14764,N_14721);
or U15472 (N_15472,N_14707,N_14857);
nand U15473 (N_15473,N_14822,N_14498);
or U15474 (N_15474,N_14583,N_14401);
nor U15475 (N_15475,N_14511,N_14587);
nand U15476 (N_15476,N_14538,N_14434);
and U15477 (N_15477,N_14965,N_14951);
nor U15478 (N_15478,N_14581,N_14920);
or U15479 (N_15479,N_14468,N_14666);
or U15480 (N_15480,N_14714,N_14523);
nor U15481 (N_15481,N_14630,N_14635);
nand U15482 (N_15482,N_14917,N_14836);
nand U15483 (N_15483,N_14958,N_14516);
nor U15484 (N_15484,N_14781,N_14508);
nand U15485 (N_15485,N_14700,N_14446);
nand U15486 (N_15486,N_14713,N_14414);
nor U15487 (N_15487,N_14867,N_14948);
nand U15488 (N_15488,N_14518,N_14535);
nor U15489 (N_15489,N_14606,N_14837);
nor U15490 (N_15490,N_14689,N_14776);
or U15491 (N_15491,N_14928,N_14571);
nor U15492 (N_15492,N_14790,N_14851);
nand U15493 (N_15493,N_14640,N_14484);
and U15494 (N_15494,N_14834,N_14437);
nor U15495 (N_15495,N_14567,N_14804);
or U15496 (N_15496,N_14908,N_14485);
or U15497 (N_15497,N_14458,N_14991);
or U15498 (N_15498,N_14906,N_14913);
and U15499 (N_15499,N_14636,N_14683);
nand U15500 (N_15500,N_14736,N_14683);
nand U15501 (N_15501,N_14811,N_14514);
or U15502 (N_15502,N_14607,N_14927);
xor U15503 (N_15503,N_14533,N_14994);
and U15504 (N_15504,N_14569,N_14951);
and U15505 (N_15505,N_14465,N_14862);
xnor U15506 (N_15506,N_14873,N_14580);
and U15507 (N_15507,N_14810,N_14914);
nand U15508 (N_15508,N_14979,N_14571);
nand U15509 (N_15509,N_14695,N_14457);
or U15510 (N_15510,N_14460,N_14920);
nand U15511 (N_15511,N_14877,N_14656);
and U15512 (N_15512,N_14936,N_14678);
nor U15513 (N_15513,N_14894,N_14812);
nand U15514 (N_15514,N_14749,N_14850);
nor U15515 (N_15515,N_14676,N_14877);
nand U15516 (N_15516,N_14602,N_14786);
and U15517 (N_15517,N_14986,N_14424);
nand U15518 (N_15518,N_14688,N_14406);
and U15519 (N_15519,N_14591,N_14778);
or U15520 (N_15520,N_14532,N_14777);
or U15521 (N_15521,N_14545,N_14958);
nand U15522 (N_15522,N_14426,N_14468);
or U15523 (N_15523,N_14852,N_14887);
or U15524 (N_15524,N_14587,N_14590);
and U15525 (N_15525,N_14913,N_14963);
nor U15526 (N_15526,N_14847,N_14834);
nand U15527 (N_15527,N_14556,N_14954);
nor U15528 (N_15528,N_14974,N_14661);
and U15529 (N_15529,N_14678,N_14400);
and U15530 (N_15530,N_14593,N_14869);
nand U15531 (N_15531,N_14642,N_14410);
nand U15532 (N_15532,N_14493,N_14688);
or U15533 (N_15533,N_14756,N_14755);
nor U15534 (N_15534,N_14500,N_14420);
and U15535 (N_15535,N_14496,N_14738);
or U15536 (N_15536,N_14828,N_14795);
nor U15537 (N_15537,N_14906,N_14640);
and U15538 (N_15538,N_14434,N_14956);
nor U15539 (N_15539,N_14737,N_14870);
nand U15540 (N_15540,N_14726,N_14583);
and U15541 (N_15541,N_14656,N_14434);
nand U15542 (N_15542,N_14644,N_14833);
and U15543 (N_15543,N_14826,N_14978);
or U15544 (N_15544,N_14946,N_14781);
and U15545 (N_15545,N_14466,N_14502);
nor U15546 (N_15546,N_14441,N_14842);
or U15547 (N_15547,N_14444,N_14681);
nor U15548 (N_15548,N_14671,N_14412);
nand U15549 (N_15549,N_14615,N_14651);
nor U15550 (N_15550,N_14508,N_14433);
nand U15551 (N_15551,N_14528,N_14913);
nand U15552 (N_15552,N_14873,N_14518);
or U15553 (N_15553,N_14767,N_14973);
nand U15554 (N_15554,N_14789,N_14782);
and U15555 (N_15555,N_14711,N_14769);
nand U15556 (N_15556,N_14771,N_14963);
and U15557 (N_15557,N_14440,N_14980);
or U15558 (N_15558,N_14576,N_14635);
nand U15559 (N_15559,N_14623,N_14678);
nand U15560 (N_15560,N_14440,N_14635);
nor U15561 (N_15561,N_14706,N_14502);
or U15562 (N_15562,N_14463,N_14880);
nor U15563 (N_15563,N_14565,N_14666);
or U15564 (N_15564,N_14624,N_14899);
or U15565 (N_15565,N_14592,N_14504);
and U15566 (N_15566,N_14532,N_14657);
nor U15567 (N_15567,N_14501,N_14480);
nor U15568 (N_15568,N_14477,N_14947);
nor U15569 (N_15569,N_14778,N_14639);
nand U15570 (N_15570,N_14613,N_14515);
or U15571 (N_15571,N_14593,N_14923);
xnor U15572 (N_15572,N_14899,N_14421);
and U15573 (N_15573,N_14925,N_14637);
and U15574 (N_15574,N_14878,N_14539);
and U15575 (N_15575,N_14668,N_14935);
nand U15576 (N_15576,N_14927,N_14413);
and U15577 (N_15577,N_14913,N_14785);
or U15578 (N_15578,N_14611,N_14764);
or U15579 (N_15579,N_14775,N_14434);
nand U15580 (N_15580,N_14557,N_14773);
nor U15581 (N_15581,N_14460,N_14789);
or U15582 (N_15582,N_14514,N_14936);
or U15583 (N_15583,N_14611,N_14664);
or U15584 (N_15584,N_14404,N_14898);
nand U15585 (N_15585,N_14924,N_14926);
nor U15586 (N_15586,N_14494,N_14957);
or U15587 (N_15587,N_14546,N_14973);
and U15588 (N_15588,N_14999,N_14758);
nand U15589 (N_15589,N_14824,N_14573);
and U15590 (N_15590,N_14582,N_14930);
nand U15591 (N_15591,N_14715,N_14738);
or U15592 (N_15592,N_14816,N_14885);
nand U15593 (N_15593,N_14494,N_14841);
or U15594 (N_15594,N_14653,N_14996);
nand U15595 (N_15595,N_14437,N_14603);
nor U15596 (N_15596,N_14737,N_14861);
or U15597 (N_15597,N_14976,N_14400);
nand U15598 (N_15598,N_14709,N_14782);
nand U15599 (N_15599,N_14712,N_14490);
and U15600 (N_15600,N_15244,N_15451);
or U15601 (N_15601,N_15230,N_15257);
nor U15602 (N_15602,N_15071,N_15590);
nor U15603 (N_15603,N_15054,N_15465);
nor U15604 (N_15604,N_15048,N_15216);
and U15605 (N_15605,N_15219,N_15192);
or U15606 (N_15606,N_15481,N_15079);
nand U15607 (N_15607,N_15583,N_15405);
xor U15608 (N_15608,N_15328,N_15169);
or U15609 (N_15609,N_15092,N_15524);
nor U15610 (N_15610,N_15565,N_15027);
or U15611 (N_15611,N_15443,N_15452);
nor U15612 (N_15612,N_15040,N_15287);
and U15613 (N_15613,N_15401,N_15100);
nand U15614 (N_15614,N_15359,N_15528);
and U15615 (N_15615,N_15435,N_15099);
or U15616 (N_15616,N_15517,N_15539);
nor U15617 (N_15617,N_15274,N_15156);
and U15618 (N_15618,N_15260,N_15205);
or U15619 (N_15619,N_15547,N_15407);
and U15620 (N_15620,N_15128,N_15397);
and U15621 (N_15621,N_15327,N_15095);
or U15622 (N_15622,N_15352,N_15000);
nand U15623 (N_15623,N_15320,N_15179);
and U15624 (N_15624,N_15564,N_15024);
nand U15625 (N_15625,N_15368,N_15271);
nor U15626 (N_15626,N_15259,N_15508);
or U15627 (N_15627,N_15002,N_15090);
nand U15628 (N_15628,N_15548,N_15431);
nand U15629 (N_15629,N_15258,N_15017);
or U15630 (N_15630,N_15356,N_15218);
or U15631 (N_15631,N_15323,N_15595);
nand U15632 (N_15632,N_15113,N_15588);
nand U15633 (N_15633,N_15266,N_15275);
or U15634 (N_15634,N_15006,N_15228);
nor U15635 (N_15635,N_15083,N_15396);
nor U15636 (N_15636,N_15341,N_15459);
or U15637 (N_15637,N_15206,N_15007);
nand U15638 (N_15638,N_15303,N_15560);
and U15639 (N_15639,N_15240,N_15331);
nand U15640 (N_15640,N_15150,N_15133);
and U15641 (N_15641,N_15387,N_15585);
or U15642 (N_15642,N_15297,N_15020);
nor U15643 (N_15643,N_15505,N_15313);
nor U15644 (N_15644,N_15005,N_15335);
nor U15645 (N_15645,N_15582,N_15183);
nand U15646 (N_15646,N_15542,N_15164);
and U15647 (N_15647,N_15449,N_15509);
nor U15648 (N_15648,N_15042,N_15393);
nand U15649 (N_15649,N_15533,N_15536);
nand U15650 (N_15650,N_15062,N_15468);
and U15651 (N_15651,N_15483,N_15569);
and U15652 (N_15652,N_15032,N_15383);
nand U15653 (N_15653,N_15281,N_15476);
and U15654 (N_15654,N_15082,N_15510);
nand U15655 (N_15655,N_15428,N_15105);
nor U15656 (N_15656,N_15047,N_15364);
or U15657 (N_15657,N_15031,N_15186);
nand U15658 (N_15658,N_15446,N_15529);
or U15659 (N_15659,N_15370,N_15298);
nand U15660 (N_15660,N_15424,N_15068);
nand U15661 (N_15661,N_15417,N_15550);
nor U15662 (N_15662,N_15035,N_15125);
or U15663 (N_15663,N_15361,N_15430);
and U15664 (N_15664,N_15110,N_15175);
xnor U15665 (N_15665,N_15333,N_15367);
and U15666 (N_15666,N_15294,N_15208);
nand U15667 (N_15667,N_15112,N_15315);
and U15668 (N_15668,N_15347,N_15339);
or U15669 (N_15669,N_15130,N_15447);
nand U15670 (N_15670,N_15530,N_15104);
and U15671 (N_15671,N_15085,N_15592);
nor U15672 (N_15672,N_15060,N_15144);
nor U15673 (N_15673,N_15302,N_15344);
nand U15674 (N_15674,N_15563,N_15498);
nor U15675 (N_15675,N_15028,N_15190);
or U15676 (N_15676,N_15391,N_15295);
nor U15677 (N_15677,N_15038,N_15423);
or U15678 (N_15678,N_15107,N_15593);
or U15679 (N_15679,N_15490,N_15010);
or U15680 (N_15680,N_15078,N_15037);
and U15681 (N_15681,N_15293,N_15012);
and U15682 (N_15682,N_15545,N_15157);
or U15683 (N_15683,N_15167,N_15403);
or U15684 (N_15684,N_15185,N_15375);
and U15685 (N_15685,N_15504,N_15402);
nand U15686 (N_15686,N_15210,N_15337);
and U15687 (N_15687,N_15362,N_15189);
and U15688 (N_15688,N_15366,N_15102);
or U15689 (N_15689,N_15022,N_15577);
nand U15690 (N_15690,N_15457,N_15586);
or U15691 (N_15691,N_15077,N_15571);
and U15692 (N_15692,N_15096,N_15482);
or U15693 (N_15693,N_15534,N_15348);
and U15694 (N_15694,N_15045,N_15154);
nor U15695 (N_15695,N_15118,N_15248);
xor U15696 (N_15696,N_15225,N_15426);
and U15697 (N_15697,N_15301,N_15217);
and U15698 (N_15698,N_15199,N_15381);
nand U15699 (N_15699,N_15233,N_15029);
or U15700 (N_15700,N_15404,N_15312);
nand U15701 (N_15701,N_15440,N_15261);
nor U15702 (N_15702,N_15345,N_15254);
or U15703 (N_15703,N_15554,N_15001);
and U15704 (N_15704,N_15235,N_15292);
or U15705 (N_15705,N_15306,N_15086);
nor U15706 (N_15706,N_15149,N_15455);
nor U15707 (N_15707,N_15013,N_15142);
and U15708 (N_15708,N_15052,N_15456);
or U15709 (N_15709,N_15329,N_15231);
nand U15710 (N_15710,N_15507,N_15474);
nor U15711 (N_15711,N_15273,N_15503);
nor U15712 (N_15712,N_15145,N_15497);
and U15713 (N_15713,N_15172,N_15053);
and U15714 (N_15714,N_15553,N_15194);
and U15715 (N_15715,N_15514,N_15538);
nand U15716 (N_15716,N_15296,N_15245);
nor U15717 (N_15717,N_15413,N_15420);
nor U15718 (N_15718,N_15502,N_15477);
and U15719 (N_15719,N_15117,N_15270);
nor U15720 (N_15720,N_15523,N_15392);
and U15721 (N_15721,N_15147,N_15226);
or U15722 (N_15722,N_15436,N_15023);
and U15723 (N_15723,N_15203,N_15171);
nand U15724 (N_15724,N_15044,N_15198);
or U15725 (N_15725,N_15450,N_15251);
nand U15726 (N_15726,N_15232,N_15444);
or U15727 (N_15727,N_15527,N_15304);
or U15728 (N_15728,N_15276,N_15019);
and U15729 (N_15729,N_15499,N_15568);
nand U15730 (N_15730,N_15526,N_15419);
nor U15731 (N_15731,N_15464,N_15166);
or U15732 (N_15732,N_15097,N_15200);
and U15733 (N_15733,N_15575,N_15491);
nand U15734 (N_15734,N_15136,N_15058);
nor U15735 (N_15735,N_15003,N_15411);
nor U15736 (N_15736,N_15134,N_15546);
or U15737 (N_15737,N_15265,N_15390);
nor U15738 (N_15738,N_15253,N_15242);
nor U15739 (N_15739,N_15434,N_15406);
xnor U15740 (N_15740,N_15472,N_15422);
nor U15741 (N_15741,N_15063,N_15429);
nand U15742 (N_15742,N_15358,N_15181);
or U15743 (N_15743,N_15234,N_15321);
or U15744 (N_15744,N_15469,N_15425);
nand U15745 (N_15745,N_15478,N_15594);
or U15746 (N_15746,N_15014,N_15256);
nor U15747 (N_15747,N_15552,N_15069);
and U15748 (N_15748,N_15215,N_15353);
or U15749 (N_15749,N_15123,N_15089);
nor U15750 (N_15750,N_15140,N_15525);
nor U15751 (N_15751,N_15573,N_15070);
and U15752 (N_15752,N_15109,N_15088);
or U15753 (N_15753,N_15416,N_15541);
nor U15754 (N_15754,N_15414,N_15162);
and U15755 (N_15755,N_15350,N_15284);
nand U15756 (N_15756,N_15369,N_15039);
nand U15757 (N_15757,N_15138,N_15555);
or U15758 (N_15758,N_15151,N_15501);
and U15759 (N_15759,N_15388,N_15243);
or U15760 (N_15760,N_15379,N_15229);
and U15761 (N_15761,N_15036,N_15222);
and U15762 (N_15762,N_15394,N_15008);
and U15763 (N_15763,N_15378,N_15280);
and U15764 (N_15764,N_15374,N_15050);
nor U15765 (N_15765,N_15597,N_15250);
or U15766 (N_15766,N_15584,N_15355);
nor U15767 (N_15767,N_15141,N_15579);
or U15768 (N_15768,N_15561,N_15343);
nand U15769 (N_15769,N_15471,N_15241);
or U15770 (N_15770,N_15439,N_15021);
and U15771 (N_15771,N_15400,N_15371);
nand U15772 (N_15772,N_15496,N_15268);
xor U15773 (N_15773,N_15290,N_15463);
nand U15774 (N_15774,N_15227,N_15389);
nor U15775 (N_15775,N_15380,N_15349);
nand U15776 (N_15776,N_15066,N_15191);
and U15777 (N_15777,N_15460,N_15453);
nand U15778 (N_15778,N_15532,N_15055);
nand U15779 (N_15779,N_15318,N_15148);
nor U15780 (N_15780,N_15516,N_15272);
and U15781 (N_15781,N_15016,N_15466);
and U15782 (N_15782,N_15330,N_15484);
nand U15783 (N_15783,N_15412,N_15515);
and U15784 (N_15784,N_15076,N_15269);
nor U15785 (N_15785,N_15421,N_15121);
and U15786 (N_15786,N_15566,N_15540);
or U15787 (N_15787,N_15357,N_15521);
nand U15788 (N_15788,N_15018,N_15286);
or U15789 (N_15789,N_15173,N_15415);
nor U15790 (N_15790,N_15363,N_15493);
nand U15791 (N_15791,N_15311,N_15500);
or U15792 (N_15792,N_15061,N_15152);
and U15793 (N_15793,N_15091,N_15159);
nand U15794 (N_15794,N_15116,N_15596);
nand U15795 (N_15795,N_15084,N_15108);
and U15796 (N_15796,N_15188,N_15127);
nor U15797 (N_15797,N_15432,N_15479);
nand U15798 (N_15798,N_15213,N_15139);
nand U15799 (N_15799,N_15262,N_15283);
xnor U15800 (N_15800,N_15319,N_15506);
or U15801 (N_15801,N_15065,N_15174);
nand U15802 (N_15802,N_15454,N_15067);
nand U15803 (N_15803,N_15193,N_15072);
and U15804 (N_15804,N_15543,N_15161);
xor U15805 (N_15805,N_15520,N_15236);
and U15806 (N_15806,N_15305,N_15030);
or U15807 (N_15807,N_15373,N_15209);
or U15808 (N_15808,N_15160,N_15587);
and U15809 (N_15809,N_15338,N_15537);
nor U15810 (N_15810,N_15122,N_15187);
and U15811 (N_15811,N_15438,N_15458);
nor U15812 (N_15812,N_15080,N_15201);
nand U15813 (N_15813,N_15342,N_15212);
nand U15814 (N_15814,N_15289,N_15559);
or U15815 (N_15815,N_15049,N_15336);
nor U15816 (N_15816,N_15599,N_15309);
nand U15817 (N_15817,N_15247,N_15015);
or U15818 (N_15818,N_15448,N_15011);
and U15819 (N_15819,N_15511,N_15211);
and U15820 (N_15820,N_15299,N_15494);
and U15821 (N_15821,N_15376,N_15427);
or U15822 (N_15822,N_15317,N_15103);
nor U15823 (N_15823,N_15581,N_15155);
and U15824 (N_15824,N_15470,N_15278);
and U15825 (N_15825,N_15180,N_15495);
and U15826 (N_15826,N_15467,N_15195);
nor U15827 (N_15827,N_15398,N_15382);
nor U15828 (N_15828,N_15132,N_15489);
and U15829 (N_15829,N_15170,N_15143);
nor U15830 (N_15830,N_15246,N_15480);
nand U15831 (N_15831,N_15551,N_15360);
or U15832 (N_15832,N_15239,N_15372);
nand U15833 (N_15833,N_15549,N_15314);
or U15834 (N_15834,N_15519,N_15263);
nand U15835 (N_15835,N_15129,N_15324);
nand U15836 (N_15836,N_15325,N_15051);
or U15837 (N_15837,N_15056,N_15334);
or U15838 (N_15838,N_15114,N_15267);
xnor U15839 (N_15839,N_15081,N_15558);
nand U15840 (N_15840,N_15340,N_15316);
and U15841 (N_15841,N_15163,N_15461);
and U15842 (N_15842,N_15310,N_15308);
or U15843 (N_15843,N_15101,N_15043);
nand U15844 (N_15844,N_15445,N_15223);
nand U15845 (N_15845,N_15395,N_15153);
nor U15846 (N_15846,N_15473,N_15146);
nor U15847 (N_15847,N_15197,N_15282);
nand U15848 (N_15848,N_15238,N_15557);
nor U15849 (N_15849,N_15074,N_15093);
nand U15850 (N_15850,N_15572,N_15377);
nor U15851 (N_15851,N_15576,N_15598);
nand U15852 (N_15852,N_15437,N_15409);
nor U15853 (N_15853,N_15111,N_15513);
and U15854 (N_15854,N_15556,N_15106);
nand U15855 (N_15855,N_15224,N_15580);
and U15856 (N_15856,N_15041,N_15589);
or U15857 (N_15857,N_15574,N_15119);
or U15858 (N_15858,N_15518,N_15178);
nor U15859 (N_15859,N_15120,N_15567);
or U15860 (N_15860,N_15064,N_15326);
and U15861 (N_15861,N_15291,N_15264);
or U15862 (N_15862,N_15182,N_15237);
or U15863 (N_15863,N_15535,N_15591);
or U15864 (N_15864,N_15399,N_15196);
nand U15865 (N_15865,N_15220,N_15418);
and U15866 (N_15866,N_15386,N_15512);
and U15867 (N_15867,N_15137,N_15073);
or U15868 (N_15868,N_15255,N_15578);
nand U15869 (N_15869,N_15351,N_15184);
nor U15870 (N_15870,N_15462,N_15279);
nand U15871 (N_15871,N_15562,N_15485);
nand U15872 (N_15872,N_15094,N_15026);
and U15873 (N_15873,N_15300,N_15075);
or U15874 (N_15874,N_15115,N_15441);
and U15875 (N_15875,N_15098,N_15408);
or U15876 (N_15876,N_15214,N_15277);
nor U15877 (N_15877,N_15135,N_15009);
xnor U15878 (N_15878,N_15033,N_15488);
or U15879 (N_15879,N_15177,N_15131);
and U15880 (N_15880,N_15087,N_15046);
nor U15881 (N_15881,N_15354,N_15176);
or U15882 (N_15882,N_15034,N_15249);
or U15883 (N_15883,N_15531,N_15486);
or U15884 (N_15884,N_15365,N_15433);
and U15885 (N_15885,N_15285,N_15025);
xnor U15886 (N_15886,N_15322,N_15252);
nand U15887 (N_15887,N_15126,N_15207);
nor U15888 (N_15888,N_15384,N_15570);
and U15889 (N_15889,N_15492,N_15544);
or U15890 (N_15890,N_15165,N_15158);
xor U15891 (N_15891,N_15124,N_15059);
nor U15892 (N_15892,N_15221,N_15332);
nor U15893 (N_15893,N_15307,N_15057);
and U15894 (N_15894,N_15522,N_15202);
nor U15895 (N_15895,N_15346,N_15204);
or U15896 (N_15896,N_15487,N_15410);
nand U15897 (N_15897,N_15385,N_15004);
or U15898 (N_15898,N_15475,N_15442);
and U15899 (N_15899,N_15288,N_15168);
nand U15900 (N_15900,N_15119,N_15161);
xor U15901 (N_15901,N_15368,N_15409);
and U15902 (N_15902,N_15195,N_15455);
or U15903 (N_15903,N_15268,N_15293);
nor U15904 (N_15904,N_15596,N_15233);
nand U15905 (N_15905,N_15496,N_15061);
nor U15906 (N_15906,N_15272,N_15393);
and U15907 (N_15907,N_15094,N_15557);
and U15908 (N_15908,N_15569,N_15053);
and U15909 (N_15909,N_15300,N_15331);
xor U15910 (N_15910,N_15556,N_15184);
or U15911 (N_15911,N_15442,N_15150);
and U15912 (N_15912,N_15238,N_15559);
nand U15913 (N_15913,N_15243,N_15329);
nand U15914 (N_15914,N_15012,N_15250);
and U15915 (N_15915,N_15299,N_15360);
and U15916 (N_15916,N_15391,N_15099);
nand U15917 (N_15917,N_15362,N_15404);
nor U15918 (N_15918,N_15583,N_15058);
or U15919 (N_15919,N_15067,N_15495);
or U15920 (N_15920,N_15333,N_15301);
or U15921 (N_15921,N_15554,N_15357);
nand U15922 (N_15922,N_15396,N_15398);
and U15923 (N_15923,N_15233,N_15089);
and U15924 (N_15924,N_15052,N_15491);
nand U15925 (N_15925,N_15257,N_15038);
nand U15926 (N_15926,N_15190,N_15554);
or U15927 (N_15927,N_15406,N_15225);
or U15928 (N_15928,N_15154,N_15340);
or U15929 (N_15929,N_15119,N_15342);
nor U15930 (N_15930,N_15385,N_15010);
and U15931 (N_15931,N_15134,N_15282);
and U15932 (N_15932,N_15317,N_15014);
or U15933 (N_15933,N_15519,N_15325);
nor U15934 (N_15934,N_15505,N_15447);
nor U15935 (N_15935,N_15378,N_15105);
nor U15936 (N_15936,N_15585,N_15444);
and U15937 (N_15937,N_15518,N_15052);
or U15938 (N_15938,N_15055,N_15416);
and U15939 (N_15939,N_15470,N_15413);
or U15940 (N_15940,N_15194,N_15572);
or U15941 (N_15941,N_15066,N_15394);
and U15942 (N_15942,N_15057,N_15067);
and U15943 (N_15943,N_15528,N_15458);
nor U15944 (N_15944,N_15079,N_15061);
xnor U15945 (N_15945,N_15045,N_15464);
xnor U15946 (N_15946,N_15122,N_15035);
nand U15947 (N_15947,N_15356,N_15135);
or U15948 (N_15948,N_15263,N_15191);
nand U15949 (N_15949,N_15271,N_15511);
or U15950 (N_15950,N_15209,N_15187);
or U15951 (N_15951,N_15582,N_15563);
nor U15952 (N_15952,N_15300,N_15089);
or U15953 (N_15953,N_15198,N_15318);
nand U15954 (N_15954,N_15338,N_15410);
or U15955 (N_15955,N_15530,N_15541);
nand U15956 (N_15956,N_15314,N_15566);
xor U15957 (N_15957,N_15513,N_15039);
nor U15958 (N_15958,N_15144,N_15203);
nand U15959 (N_15959,N_15214,N_15365);
nand U15960 (N_15960,N_15227,N_15406);
nand U15961 (N_15961,N_15092,N_15543);
or U15962 (N_15962,N_15370,N_15553);
nand U15963 (N_15963,N_15554,N_15303);
nand U15964 (N_15964,N_15284,N_15580);
nor U15965 (N_15965,N_15077,N_15446);
and U15966 (N_15966,N_15265,N_15113);
nor U15967 (N_15967,N_15031,N_15371);
nor U15968 (N_15968,N_15217,N_15424);
or U15969 (N_15969,N_15098,N_15344);
nor U15970 (N_15970,N_15437,N_15347);
or U15971 (N_15971,N_15066,N_15048);
or U15972 (N_15972,N_15115,N_15496);
or U15973 (N_15973,N_15204,N_15284);
and U15974 (N_15974,N_15095,N_15483);
or U15975 (N_15975,N_15356,N_15148);
nand U15976 (N_15976,N_15498,N_15119);
or U15977 (N_15977,N_15098,N_15224);
and U15978 (N_15978,N_15133,N_15529);
nor U15979 (N_15979,N_15426,N_15535);
and U15980 (N_15980,N_15089,N_15401);
nor U15981 (N_15981,N_15474,N_15288);
or U15982 (N_15982,N_15555,N_15000);
and U15983 (N_15983,N_15516,N_15447);
or U15984 (N_15984,N_15252,N_15557);
nor U15985 (N_15985,N_15011,N_15322);
nand U15986 (N_15986,N_15292,N_15586);
or U15987 (N_15987,N_15459,N_15188);
and U15988 (N_15988,N_15258,N_15405);
nand U15989 (N_15989,N_15546,N_15394);
nand U15990 (N_15990,N_15352,N_15073);
nand U15991 (N_15991,N_15169,N_15324);
and U15992 (N_15992,N_15362,N_15471);
nor U15993 (N_15993,N_15213,N_15083);
or U15994 (N_15994,N_15392,N_15076);
nor U15995 (N_15995,N_15197,N_15180);
nand U15996 (N_15996,N_15544,N_15593);
or U15997 (N_15997,N_15587,N_15084);
and U15998 (N_15998,N_15228,N_15089);
or U15999 (N_15999,N_15337,N_15235);
xor U16000 (N_16000,N_15087,N_15240);
nand U16001 (N_16001,N_15311,N_15455);
nor U16002 (N_16002,N_15005,N_15452);
nor U16003 (N_16003,N_15228,N_15533);
nand U16004 (N_16004,N_15387,N_15549);
and U16005 (N_16005,N_15291,N_15589);
and U16006 (N_16006,N_15013,N_15413);
nor U16007 (N_16007,N_15438,N_15334);
and U16008 (N_16008,N_15268,N_15528);
nand U16009 (N_16009,N_15366,N_15144);
or U16010 (N_16010,N_15500,N_15297);
nand U16011 (N_16011,N_15248,N_15535);
xor U16012 (N_16012,N_15495,N_15248);
nor U16013 (N_16013,N_15213,N_15432);
or U16014 (N_16014,N_15295,N_15227);
nor U16015 (N_16015,N_15091,N_15082);
xnor U16016 (N_16016,N_15113,N_15208);
nor U16017 (N_16017,N_15411,N_15422);
nor U16018 (N_16018,N_15296,N_15380);
or U16019 (N_16019,N_15231,N_15057);
and U16020 (N_16020,N_15582,N_15232);
and U16021 (N_16021,N_15222,N_15115);
nor U16022 (N_16022,N_15151,N_15131);
or U16023 (N_16023,N_15186,N_15178);
or U16024 (N_16024,N_15552,N_15176);
xnor U16025 (N_16025,N_15384,N_15184);
and U16026 (N_16026,N_15339,N_15302);
nor U16027 (N_16027,N_15561,N_15260);
nand U16028 (N_16028,N_15358,N_15110);
and U16029 (N_16029,N_15321,N_15168);
nor U16030 (N_16030,N_15309,N_15067);
nand U16031 (N_16031,N_15575,N_15431);
nand U16032 (N_16032,N_15208,N_15157);
nand U16033 (N_16033,N_15043,N_15075);
nand U16034 (N_16034,N_15278,N_15453);
nor U16035 (N_16035,N_15145,N_15385);
or U16036 (N_16036,N_15336,N_15005);
nand U16037 (N_16037,N_15403,N_15544);
nand U16038 (N_16038,N_15214,N_15088);
and U16039 (N_16039,N_15107,N_15337);
nand U16040 (N_16040,N_15485,N_15247);
and U16041 (N_16041,N_15075,N_15051);
xnor U16042 (N_16042,N_15217,N_15533);
nor U16043 (N_16043,N_15180,N_15396);
and U16044 (N_16044,N_15472,N_15375);
and U16045 (N_16045,N_15532,N_15189);
nand U16046 (N_16046,N_15359,N_15403);
and U16047 (N_16047,N_15118,N_15117);
or U16048 (N_16048,N_15138,N_15310);
or U16049 (N_16049,N_15296,N_15597);
or U16050 (N_16050,N_15512,N_15195);
and U16051 (N_16051,N_15161,N_15513);
and U16052 (N_16052,N_15548,N_15405);
nand U16053 (N_16053,N_15016,N_15213);
or U16054 (N_16054,N_15538,N_15061);
nor U16055 (N_16055,N_15572,N_15519);
nor U16056 (N_16056,N_15287,N_15014);
nor U16057 (N_16057,N_15210,N_15563);
and U16058 (N_16058,N_15536,N_15428);
xnor U16059 (N_16059,N_15013,N_15426);
and U16060 (N_16060,N_15245,N_15461);
or U16061 (N_16061,N_15507,N_15050);
nor U16062 (N_16062,N_15048,N_15457);
or U16063 (N_16063,N_15518,N_15187);
or U16064 (N_16064,N_15484,N_15585);
or U16065 (N_16065,N_15587,N_15564);
nand U16066 (N_16066,N_15443,N_15548);
and U16067 (N_16067,N_15367,N_15324);
nand U16068 (N_16068,N_15469,N_15556);
or U16069 (N_16069,N_15459,N_15026);
nand U16070 (N_16070,N_15326,N_15194);
and U16071 (N_16071,N_15458,N_15126);
xor U16072 (N_16072,N_15592,N_15052);
nand U16073 (N_16073,N_15214,N_15183);
nand U16074 (N_16074,N_15264,N_15224);
xor U16075 (N_16075,N_15019,N_15082);
and U16076 (N_16076,N_15164,N_15529);
and U16077 (N_16077,N_15278,N_15538);
or U16078 (N_16078,N_15021,N_15029);
nand U16079 (N_16079,N_15119,N_15409);
and U16080 (N_16080,N_15499,N_15306);
nor U16081 (N_16081,N_15161,N_15090);
nand U16082 (N_16082,N_15452,N_15052);
nor U16083 (N_16083,N_15136,N_15402);
or U16084 (N_16084,N_15336,N_15213);
nand U16085 (N_16085,N_15300,N_15456);
and U16086 (N_16086,N_15308,N_15170);
nand U16087 (N_16087,N_15593,N_15015);
nand U16088 (N_16088,N_15320,N_15496);
nor U16089 (N_16089,N_15308,N_15262);
and U16090 (N_16090,N_15332,N_15181);
or U16091 (N_16091,N_15210,N_15495);
and U16092 (N_16092,N_15344,N_15485);
nand U16093 (N_16093,N_15286,N_15546);
nand U16094 (N_16094,N_15297,N_15042);
nand U16095 (N_16095,N_15383,N_15592);
and U16096 (N_16096,N_15327,N_15379);
or U16097 (N_16097,N_15224,N_15299);
or U16098 (N_16098,N_15586,N_15102);
and U16099 (N_16099,N_15264,N_15510);
or U16100 (N_16100,N_15289,N_15506);
nor U16101 (N_16101,N_15283,N_15386);
or U16102 (N_16102,N_15194,N_15396);
nand U16103 (N_16103,N_15489,N_15560);
or U16104 (N_16104,N_15324,N_15200);
nand U16105 (N_16105,N_15359,N_15363);
or U16106 (N_16106,N_15312,N_15210);
nor U16107 (N_16107,N_15374,N_15575);
nand U16108 (N_16108,N_15267,N_15323);
nor U16109 (N_16109,N_15245,N_15043);
or U16110 (N_16110,N_15413,N_15519);
and U16111 (N_16111,N_15576,N_15476);
nor U16112 (N_16112,N_15083,N_15391);
nand U16113 (N_16113,N_15557,N_15051);
nor U16114 (N_16114,N_15480,N_15391);
and U16115 (N_16115,N_15255,N_15202);
or U16116 (N_16116,N_15534,N_15030);
nor U16117 (N_16117,N_15332,N_15444);
nand U16118 (N_16118,N_15560,N_15507);
and U16119 (N_16119,N_15402,N_15568);
nor U16120 (N_16120,N_15459,N_15062);
or U16121 (N_16121,N_15383,N_15379);
nor U16122 (N_16122,N_15198,N_15239);
nor U16123 (N_16123,N_15084,N_15595);
nor U16124 (N_16124,N_15437,N_15581);
nand U16125 (N_16125,N_15205,N_15279);
or U16126 (N_16126,N_15306,N_15529);
or U16127 (N_16127,N_15032,N_15466);
or U16128 (N_16128,N_15090,N_15130);
and U16129 (N_16129,N_15225,N_15107);
nor U16130 (N_16130,N_15010,N_15005);
nor U16131 (N_16131,N_15247,N_15348);
nand U16132 (N_16132,N_15298,N_15484);
nand U16133 (N_16133,N_15415,N_15265);
nor U16134 (N_16134,N_15015,N_15378);
and U16135 (N_16135,N_15410,N_15555);
nor U16136 (N_16136,N_15052,N_15401);
or U16137 (N_16137,N_15373,N_15291);
or U16138 (N_16138,N_15288,N_15109);
xnor U16139 (N_16139,N_15461,N_15585);
nand U16140 (N_16140,N_15573,N_15441);
nand U16141 (N_16141,N_15570,N_15514);
and U16142 (N_16142,N_15203,N_15108);
and U16143 (N_16143,N_15414,N_15222);
nor U16144 (N_16144,N_15447,N_15030);
or U16145 (N_16145,N_15529,N_15182);
and U16146 (N_16146,N_15179,N_15475);
nor U16147 (N_16147,N_15062,N_15038);
or U16148 (N_16148,N_15433,N_15161);
nand U16149 (N_16149,N_15003,N_15122);
nand U16150 (N_16150,N_15394,N_15069);
or U16151 (N_16151,N_15148,N_15500);
nand U16152 (N_16152,N_15449,N_15285);
or U16153 (N_16153,N_15539,N_15516);
nor U16154 (N_16154,N_15380,N_15282);
nor U16155 (N_16155,N_15157,N_15356);
and U16156 (N_16156,N_15284,N_15330);
or U16157 (N_16157,N_15527,N_15378);
and U16158 (N_16158,N_15355,N_15435);
nand U16159 (N_16159,N_15224,N_15121);
nand U16160 (N_16160,N_15596,N_15297);
or U16161 (N_16161,N_15101,N_15091);
nand U16162 (N_16162,N_15388,N_15341);
xnor U16163 (N_16163,N_15018,N_15120);
nor U16164 (N_16164,N_15388,N_15205);
and U16165 (N_16165,N_15342,N_15122);
or U16166 (N_16166,N_15513,N_15557);
and U16167 (N_16167,N_15214,N_15341);
and U16168 (N_16168,N_15181,N_15132);
nor U16169 (N_16169,N_15575,N_15331);
or U16170 (N_16170,N_15591,N_15569);
nand U16171 (N_16171,N_15360,N_15273);
or U16172 (N_16172,N_15269,N_15380);
nand U16173 (N_16173,N_15325,N_15363);
and U16174 (N_16174,N_15153,N_15308);
nor U16175 (N_16175,N_15202,N_15185);
and U16176 (N_16176,N_15157,N_15411);
and U16177 (N_16177,N_15234,N_15419);
nor U16178 (N_16178,N_15204,N_15199);
or U16179 (N_16179,N_15377,N_15319);
nor U16180 (N_16180,N_15358,N_15543);
and U16181 (N_16181,N_15508,N_15277);
and U16182 (N_16182,N_15163,N_15188);
and U16183 (N_16183,N_15221,N_15018);
or U16184 (N_16184,N_15505,N_15390);
and U16185 (N_16185,N_15598,N_15197);
and U16186 (N_16186,N_15030,N_15041);
nand U16187 (N_16187,N_15092,N_15319);
nand U16188 (N_16188,N_15502,N_15081);
nor U16189 (N_16189,N_15015,N_15089);
nand U16190 (N_16190,N_15453,N_15493);
nor U16191 (N_16191,N_15579,N_15222);
nand U16192 (N_16192,N_15579,N_15278);
and U16193 (N_16193,N_15357,N_15506);
or U16194 (N_16194,N_15587,N_15559);
nand U16195 (N_16195,N_15333,N_15097);
and U16196 (N_16196,N_15130,N_15519);
nor U16197 (N_16197,N_15078,N_15569);
or U16198 (N_16198,N_15490,N_15045);
nand U16199 (N_16199,N_15051,N_15284);
or U16200 (N_16200,N_15972,N_16116);
or U16201 (N_16201,N_15632,N_15794);
and U16202 (N_16202,N_16191,N_15959);
nor U16203 (N_16203,N_16176,N_15873);
nor U16204 (N_16204,N_16074,N_15858);
nand U16205 (N_16205,N_15692,N_15609);
or U16206 (N_16206,N_16146,N_15960);
and U16207 (N_16207,N_15804,N_16034);
and U16208 (N_16208,N_15778,N_15900);
and U16209 (N_16209,N_15660,N_15760);
nor U16210 (N_16210,N_16183,N_15709);
or U16211 (N_16211,N_15623,N_15779);
and U16212 (N_16212,N_15711,N_15832);
xor U16213 (N_16213,N_15841,N_15734);
nand U16214 (N_16214,N_15975,N_15830);
nor U16215 (N_16215,N_16150,N_15670);
or U16216 (N_16216,N_15761,N_16157);
or U16217 (N_16217,N_15718,N_16114);
xor U16218 (N_16218,N_15849,N_15968);
and U16219 (N_16219,N_15710,N_15661);
nor U16220 (N_16220,N_16024,N_16035);
nor U16221 (N_16221,N_15921,N_15973);
nand U16222 (N_16222,N_16152,N_15684);
xor U16223 (N_16223,N_15913,N_16133);
or U16224 (N_16224,N_16067,N_16138);
or U16225 (N_16225,N_15757,N_15895);
nor U16226 (N_16226,N_16042,N_15792);
nand U16227 (N_16227,N_15813,N_15705);
or U16228 (N_16228,N_16055,N_15756);
nor U16229 (N_16229,N_15643,N_15624);
nand U16230 (N_16230,N_15826,N_16109);
nor U16231 (N_16231,N_15985,N_15912);
nand U16232 (N_16232,N_15769,N_15821);
nand U16233 (N_16233,N_15868,N_15680);
nor U16234 (N_16234,N_16120,N_15677);
or U16235 (N_16235,N_15945,N_15658);
nor U16236 (N_16236,N_15874,N_15907);
and U16237 (N_16237,N_15864,N_15822);
nor U16238 (N_16238,N_15948,N_15893);
or U16239 (N_16239,N_15630,N_15631);
xnor U16240 (N_16240,N_15862,N_15754);
nand U16241 (N_16241,N_16130,N_15818);
and U16242 (N_16242,N_15729,N_15820);
and U16243 (N_16243,N_15927,N_16196);
nand U16244 (N_16244,N_15694,N_15886);
or U16245 (N_16245,N_16148,N_15923);
and U16246 (N_16246,N_15990,N_15614);
nor U16247 (N_16247,N_15675,N_15721);
nor U16248 (N_16248,N_16032,N_16087);
nand U16249 (N_16249,N_16073,N_15938);
and U16250 (N_16250,N_15950,N_15621);
or U16251 (N_16251,N_16081,N_15723);
or U16252 (N_16252,N_15622,N_15884);
nor U16253 (N_16253,N_16180,N_15798);
or U16254 (N_16254,N_15674,N_15665);
nor U16255 (N_16255,N_15742,N_16164);
nand U16256 (N_16256,N_16190,N_15967);
nand U16257 (N_16257,N_15753,N_15640);
or U16258 (N_16258,N_15915,N_15982);
xor U16259 (N_16259,N_15612,N_15641);
and U16260 (N_16260,N_15663,N_16136);
or U16261 (N_16261,N_16007,N_15625);
and U16262 (N_16262,N_15827,N_16145);
or U16263 (N_16263,N_15936,N_16003);
and U16264 (N_16264,N_15897,N_15745);
and U16265 (N_16265,N_15800,N_15655);
nor U16266 (N_16266,N_15943,N_15823);
nand U16267 (N_16267,N_16175,N_15838);
nor U16268 (N_16268,N_16083,N_15853);
nand U16269 (N_16269,N_15777,N_16017);
nor U16270 (N_16270,N_15994,N_16044);
or U16271 (N_16271,N_16009,N_16107);
nor U16272 (N_16272,N_16173,N_16004);
and U16273 (N_16273,N_15740,N_15810);
and U16274 (N_16274,N_15683,N_15766);
and U16275 (N_16275,N_15628,N_15870);
nor U16276 (N_16276,N_15918,N_16147);
and U16277 (N_16277,N_15946,N_15771);
and U16278 (N_16278,N_15876,N_15808);
or U16279 (N_16279,N_16002,N_15966);
or U16280 (N_16280,N_16198,N_15891);
nor U16281 (N_16281,N_15840,N_16079);
and U16282 (N_16282,N_15726,N_15678);
and U16283 (N_16283,N_16025,N_15706);
or U16284 (N_16284,N_15958,N_16066);
and U16285 (N_16285,N_15957,N_16001);
or U16286 (N_16286,N_15928,N_15676);
and U16287 (N_16287,N_15793,N_16050);
nand U16288 (N_16288,N_15981,N_15656);
and U16289 (N_16289,N_16135,N_16140);
and U16290 (N_16290,N_15965,N_15940);
and U16291 (N_16291,N_16162,N_16106);
nand U16292 (N_16292,N_15882,N_16108);
or U16293 (N_16293,N_16195,N_15889);
xnor U16294 (N_16294,N_16181,N_15824);
or U16295 (N_16295,N_15629,N_15865);
nand U16296 (N_16296,N_16013,N_15932);
and U16297 (N_16297,N_15815,N_15664);
or U16298 (N_16298,N_15668,N_15775);
or U16299 (N_16299,N_15998,N_15930);
or U16300 (N_16300,N_16018,N_16099);
nor U16301 (N_16301,N_15790,N_15807);
and U16302 (N_16302,N_15704,N_16089);
or U16303 (N_16303,N_16048,N_16052);
or U16304 (N_16304,N_16072,N_15963);
or U16305 (N_16305,N_15883,N_15620);
or U16306 (N_16306,N_15781,N_16093);
nand U16307 (N_16307,N_15787,N_15910);
and U16308 (N_16308,N_15925,N_16049);
or U16309 (N_16309,N_16155,N_15847);
or U16310 (N_16310,N_16185,N_15758);
or U16311 (N_16311,N_15601,N_15690);
nand U16312 (N_16312,N_15802,N_15716);
nor U16313 (N_16313,N_15949,N_15871);
nor U16314 (N_16314,N_16121,N_15866);
and U16315 (N_16315,N_15613,N_15842);
and U16316 (N_16316,N_16122,N_16092);
nor U16317 (N_16317,N_15837,N_15686);
or U16318 (N_16318,N_15894,N_15746);
nor U16319 (N_16319,N_15652,N_15816);
nand U16320 (N_16320,N_15699,N_15717);
and U16321 (N_16321,N_15616,N_16038);
or U16322 (N_16322,N_15682,N_15770);
or U16323 (N_16323,N_16062,N_15696);
and U16324 (N_16324,N_16171,N_15911);
nor U16325 (N_16325,N_15722,N_16075);
and U16326 (N_16326,N_15695,N_15714);
nand U16327 (N_16327,N_15843,N_15752);
nand U16328 (N_16328,N_15848,N_15860);
or U16329 (N_16329,N_15984,N_15644);
or U16330 (N_16330,N_16033,N_15920);
nor U16331 (N_16331,N_15996,N_16086);
or U16332 (N_16332,N_16056,N_16161);
nand U16333 (N_16333,N_15801,N_15617);
nand U16334 (N_16334,N_15869,N_15892);
or U16335 (N_16335,N_15627,N_15735);
nor U16336 (N_16336,N_15607,N_15785);
nand U16337 (N_16337,N_15797,N_15743);
and U16338 (N_16338,N_16134,N_15780);
or U16339 (N_16339,N_15750,N_15922);
nor U16340 (N_16340,N_15877,N_16153);
nand U16341 (N_16341,N_15600,N_15834);
nand U16342 (N_16342,N_15728,N_16082);
or U16343 (N_16343,N_16127,N_16174);
nand U16344 (N_16344,N_15651,N_16059);
and U16345 (N_16345,N_16168,N_16102);
nand U16346 (N_16346,N_16101,N_15755);
nor U16347 (N_16347,N_15817,N_15909);
nor U16348 (N_16348,N_15654,N_15917);
nor U16349 (N_16349,N_16045,N_15899);
or U16350 (N_16350,N_16139,N_15805);
xnor U16351 (N_16351,N_15914,N_16169);
nor U16352 (N_16352,N_15713,N_16036);
nand U16353 (N_16353,N_15993,N_15989);
nand U16354 (N_16354,N_15691,N_15855);
nand U16355 (N_16355,N_15979,N_16047);
or U16356 (N_16356,N_15875,N_16193);
nor U16357 (N_16357,N_15795,N_15980);
or U16358 (N_16358,N_16151,N_16143);
xnor U16359 (N_16359,N_15926,N_15857);
and U16360 (N_16360,N_16124,N_16071);
and U16361 (N_16361,N_16077,N_15896);
nor U16362 (N_16362,N_15744,N_16021);
and U16363 (N_16363,N_16125,N_15712);
and U16364 (N_16364,N_16137,N_15947);
nor U16365 (N_16365,N_15955,N_16149);
and U16366 (N_16366,N_15806,N_15637);
nand U16367 (N_16367,N_16158,N_16119);
nand U16368 (N_16368,N_15854,N_15971);
and U16369 (N_16369,N_15783,N_15944);
nand U16370 (N_16370,N_16126,N_15698);
nor U16371 (N_16371,N_16080,N_15764);
or U16372 (N_16372,N_15905,N_15606);
or U16373 (N_16373,N_15693,N_15741);
and U16374 (N_16374,N_15952,N_15636);
and U16375 (N_16375,N_15653,N_15747);
and U16376 (N_16376,N_16179,N_16061);
or U16377 (N_16377,N_15732,N_15825);
and U16378 (N_16378,N_16057,N_16113);
nor U16379 (N_16379,N_15737,N_16065);
and U16380 (N_16380,N_15836,N_15799);
or U16381 (N_16381,N_15605,N_16117);
or U16382 (N_16382,N_15811,N_15681);
nor U16383 (N_16383,N_15672,N_15618);
nand U16384 (N_16384,N_16040,N_15774);
and U16385 (N_16385,N_15685,N_15916);
nand U16386 (N_16386,N_16156,N_16132);
nor U16387 (N_16387,N_16129,N_16010);
or U16388 (N_16388,N_16097,N_15978);
nor U16389 (N_16389,N_16166,N_16199);
nand U16390 (N_16390,N_16111,N_15669);
xor U16391 (N_16391,N_15772,N_16165);
nor U16392 (N_16392,N_15953,N_15679);
and U16393 (N_16393,N_15991,N_15724);
nand U16394 (N_16394,N_15715,N_15733);
or U16395 (N_16395,N_15969,N_15786);
nand U16396 (N_16396,N_16115,N_15645);
or U16397 (N_16397,N_15974,N_16068);
nor U16398 (N_16398,N_15935,N_16159);
and U16399 (N_16399,N_15687,N_16046);
nor U16400 (N_16400,N_16178,N_16016);
nand U16401 (N_16401,N_16053,N_16184);
nand U16402 (N_16402,N_15642,N_15610);
nor U16403 (N_16403,N_15852,N_15867);
nand U16404 (N_16404,N_15977,N_16085);
and U16405 (N_16405,N_16141,N_15878);
xor U16406 (N_16406,N_16000,N_16118);
nor U16407 (N_16407,N_15796,N_16028);
nand U16408 (N_16408,N_16142,N_15880);
nor U16409 (N_16409,N_15850,N_15689);
nor U16410 (N_16410,N_15863,N_16029);
nand U16411 (N_16411,N_15934,N_16076);
nand U16412 (N_16412,N_15619,N_16112);
nand U16413 (N_16413,N_16104,N_16197);
or U16414 (N_16414,N_16063,N_16012);
nand U16415 (N_16415,N_16058,N_16069);
nor U16416 (N_16416,N_15648,N_16022);
and U16417 (N_16417,N_16094,N_15872);
nand U16418 (N_16418,N_15831,N_15666);
nand U16419 (N_16419,N_15859,N_16041);
and U16420 (N_16420,N_16051,N_15997);
or U16421 (N_16421,N_15688,N_15673);
xnor U16422 (N_16422,N_15608,N_15906);
nor U16423 (N_16423,N_15707,N_15861);
and U16424 (N_16424,N_15649,N_16160);
or U16425 (N_16425,N_15839,N_15789);
nor U16426 (N_16426,N_15701,N_16070);
nor U16427 (N_16427,N_15931,N_16019);
nand U16428 (N_16428,N_15703,N_15962);
or U16429 (N_16429,N_15773,N_16163);
and U16430 (N_16430,N_15879,N_16154);
nand U16431 (N_16431,N_15941,N_15851);
and U16432 (N_16432,N_15784,N_16031);
and U16433 (N_16433,N_16030,N_15828);
nor U16434 (N_16434,N_15763,N_15759);
nand U16435 (N_16435,N_16186,N_16144);
xor U16436 (N_16436,N_16014,N_15720);
xor U16437 (N_16437,N_15833,N_16039);
nand U16438 (N_16438,N_15908,N_15727);
nor U16439 (N_16439,N_16090,N_15667);
and U16440 (N_16440,N_15888,N_15782);
nor U16441 (N_16441,N_15626,N_15788);
xnor U16442 (N_16442,N_15904,N_15748);
and U16443 (N_16443,N_15671,N_15898);
or U16444 (N_16444,N_16037,N_16105);
nand U16445 (N_16445,N_15819,N_15970);
and U16446 (N_16446,N_15803,N_16027);
xnor U16447 (N_16447,N_15767,N_15604);
nor U16448 (N_16448,N_15700,N_15738);
nand U16449 (N_16449,N_15885,N_15995);
nand U16450 (N_16450,N_15736,N_16172);
nor U16451 (N_16451,N_15647,N_15812);
nand U16452 (N_16452,N_15987,N_16103);
or U16453 (N_16453,N_15992,N_16194);
xor U16454 (N_16454,N_16098,N_15697);
or U16455 (N_16455,N_15919,N_16177);
or U16456 (N_16456,N_16011,N_16167);
nand U16457 (N_16457,N_15983,N_15603);
nand U16458 (N_16458,N_15829,N_15961);
nor U16459 (N_16459,N_16128,N_15988);
or U16460 (N_16460,N_16084,N_15951);
nand U16461 (N_16461,N_15942,N_16015);
nor U16462 (N_16462,N_15662,N_15731);
and U16463 (N_16463,N_15762,N_16110);
nor U16464 (N_16464,N_15791,N_16131);
or U16465 (N_16465,N_16170,N_15844);
nor U16466 (N_16466,N_15768,N_15902);
or U16467 (N_16467,N_16123,N_15924);
or U16468 (N_16468,N_16188,N_15730);
or U16469 (N_16469,N_15887,N_16006);
or U16470 (N_16470,N_16023,N_15954);
and U16471 (N_16471,N_15776,N_15708);
nor U16472 (N_16472,N_15856,N_15634);
or U16473 (N_16473,N_15956,N_16043);
nor U16474 (N_16474,N_16054,N_15638);
or U16475 (N_16475,N_15702,N_15881);
nand U16476 (N_16476,N_15976,N_16100);
nand U16477 (N_16477,N_15964,N_16005);
nand U16478 (N_16478,N_16020,N_15615);
or U16479 (N_16479,N_15890,N_15639);
nand U16480 (N_16480,N_16088,N_16064);
nor U16481 (N_16481,N_16060,N_15814);
or U16482 (N_16482,N_15602,N_15635);
and U16483 (N_16483,N_15719,N_15835);
nand U16484 (N_16484,N_15986,N_15999);
nand U16485 (N_16485,N_16187,N_15903);
and U16486 (N_16486,N_16182,N_15739);
or U16487 (N_16487,N_16096,N_15929);
nor U16488 (N_16488,N_15901,N_15749);
xnor U16489 (N_16489,N_16008,N_16091);
and U16490 (N_16490,N_15939,N_15933);
and U16491 (N_16491,N_15765,N_16078);
or U16492 (N_16492,N_15845,N_15650);
and U16493 (N_16493,N_16026,N_15611);
or U16494 (N_16494,N_16189,N_15659);
or U16495 (N_16495,N_16095,N_15937);
and U16496 (N_16496,N_15809,N_16192);
nor U16497 (N_16497,N_15751,N_15646);
and U16498 (N_16498,N_15657,N_15633);
or U16499 (N_16499,N_15725,N_15846);
xnor U16500 (N_16500,N_16022,N_16010);
or U16501 (N_16501,N_15635,N_15782);
nor U16502 (N_16502,N_15835,N_15634);
nor U16503 (N_16503,N_15651,N_16113);
or U16504 (N_16504,N_16044,N_15997);
nor U16505 (N_16505,N_15703,N_15743);
nand U16506 (N_16506,N_15871,N_15666);
nor U16507 (N_16507,N_15908,N_15995);
nand U16508 (N_16508,N_15695,N_15975);
nor U16509 (N_16509,N_15781,N_15783);
or U16510 (N_16510,N_15859,N_15806);
and U16511 (N_16511,N_15981,N_15643);
and U16512 (N_16512,N_15860,N_15856);
or U16513 (N_16513,N_15887,N_15982);
or U16514 (N_16514,N_16113,N_15670);
nand U16515 (N_16515,N_16072,N_15995);
nor U16516 (N_16516,N_16030,N_15968);
or U16517 (N_16517,N_16051,N_15636);
and U16518 (N_16518,N_15922,N_15686);
nand U16519 (N_16519,N_15737,N_16169);
and U16520 (N_16520,N_15646,N_15722);
xor U16521 (N_16521,N_16036,N_15880);
nand U16522 (N_16522,N_15977,N_15837);
nor U16523 (N_16523,N_15653,N_15941);
and U16524 (N_16524,N_16097,N_15839);
and U16525 (N_16525,N_15965,N_16017);
and U16526 (N_16526,N_15930,N_15908);
nand U16527 (N_16527,N_16070,N_15629);
xor U16528 (N_16528,N_16167,N_15834);
and U16529 (N_16529,N_15815,N_16163);
or U16530 (N_16530,N_15836,N_15627);
nor U16531 (N_16531,N_16195,N_16061);
nor U16532 (N_16532,N_15912,N_16169);
nand U16533 (N_16533,N_15807,N_15680);
or U16534 (N_16534,N_15705,N_16040);
nor U16535 (N_16535,N_15937,N_15700);
or U16536 (N_16536,N_16018,N_15648);
or U16537 (N_16537,N_15973,N_15602);
nand U16538 (N_16538,N_15603,N_15738);
nor U16539 (N_16539,N_16117,N_15920);
nand U16540 (N_16540,N_16175,N_15714);
and U16541 (N_16541,N_15642,N_16183);
and U16542 (N_16542,N_16086,N_15701);
and U16543 (N_16543,N_15938,N_15616);
nand U16544 (N_16544,N_15761,N_15866);
or U16545 (N_16545,N_15697,N_16057);
and U16546 (N_16546,N_15974,N_16076);
nor U16547 (N_16547,N_15934,N_16127);
and U16548 (N_16548,N_16088,N_16021);
or U16549 (N_16549,N_16024,N_15943);
and U16550 (N_16550,N_16197,N_16014);
nor U16551 (N_16551,N_15607,N_16141);
nand U16552 (N_16552,N_16177,N_15880);
or U16553 (N_16553,N_16088,N_15767);
and U16554 (N_16554,N_15631,N_16012);
or U16555 (N_16555,N_15751,N_15813);
and U16556 (N_16556,N_15846,N_16027);
or U16557 (N_16557,N_16145,N_16078);
and U16558 (N_16558,N_15888,N_15672);
nor U16559 (N_16559,N_16117,N_15900);
or U16560 (N_16560,N_15837,N_16043);
xor U16561 (N_16561,N_15679,N_16056);
nand U16562 (N_16562,N_16121,N_16140);
nand U16563 (N_16563,N_15672,N_15682);
nand U16564 (N_16564,N_15715,N_16062);
xnor U16565 (N_16565,N_15940,N_15979);
or U16566 (N_16566,N_15611,N_16145);
nand U16567 (N_16567,N_16061,N_15676);
nor U16568 (N_16568,N_15803,N_16148);
nor U16569 (N_16569,N_16017,N_15851);
nor U16570 (N_16570,N_16058,N_15790);
nor U16571 (N_16571,N_16187,N_15669);
nand U16572 (N_16572,N_16047,N_16168);
xnor U16573 (N_16573,N_15794,N_16160);
nand U16574 (N_16574,N_15825,N_15954);
or U16575 (N_16575,N_15775,N_15687);
or U16576 (N_16576,N_16044,N_15947);
nand U16577 (N_16577,N_15858,N_16109);
nand U16578 (N_16578,N_15918,N_15892);
and U16579 (N_16579,N_16034,N_15637);
and U16580 (N_16580,N_15737,N_15659);
or U16581 (N_16581,N_16109,N_16186);
nor U16582 (N_16582,N_15936,N_16081);
or U16583 (N_16583,N_16174,N_15983);
or U16584 (N_16584,N_16041,N_15999);
or U16585 (N_16585,N_15947,N_16123);
and U16586 (N_16586,N_15899,N_16193);
or U16587 (N_16587,N_15922,N_15961);
nand U16588 (N_16588,N_15748,N_16011);
xor U16589 (N_16589,N_15750,N_15977);
nor U16590 (N_16590,N_16059,N_15908);
and U16591 (N_16591,N_15984,N_16122);
nand U16592 (N_16592,N_16048,N_15877);
and U16593 (N_16593,N_15988,N_15847);
and U16594 (N_16594,N_16002,N_16056);
nand U16595 (N_16595,N_15722,N_16108);
nor U16596 (N_16596,N_15715,N_15976);
and U16597 (N_16597,N_15707,N_15737);
nor U16598 (N_16598,N_15932,N_15662);
or U16599 (N_16599,N_15863,N_16184);
nand U16600 (N_16600,N_16130,N_15733);
and U16601 (N_16601,N_15881,N_16028);
and U16602 (N_16602,N_15622,N_16106);
and U16603 (N_16603,N_15690,N_15859);
and U16604 (N_16604,N_16000,N_15834);
and U16605 (N_16605,N_15903,N_15696);
nand U16606 (N_16606,N_15890,N_16045);
and U16607 (N_16607,N_16037,N_16148);
nand U16608 (N_16608,N_15914,N_15801);
nor U16609 (N_16609,N_16129,N_16153);
nand U16610 (N_16610,N_15993,N_15617);
and U16611 (N_16611,N_16082,N_15760);
and U16612 (N_16612,N_15754,N_15982);
and U16613 (N_16613,N_15768,N_15860);
and U16614 (N_16614,N_16189,N_15893);
nand U16615 (N_16615,N_15781,N_15795);
or U16616 (N_16616,N_15954,N_15901);
nor U16617 (N_16617,N_16010,N_15762);
and U16618 (N_16618,N_15856,N_15627);
or U16619 (N_16619,N_16028,N_16092);
nor U16620 (N_16620,N_16056,N_15944);
nor U16621 (N_16621,N_16097,N_15670);
nand U16622 (N_16622,N_15985,N_16168);
nand U16623 (N_16623,N_15951,N_15751);
and U16624 (N_16624,N_16051,N_15780);
and U16625 (N_16625,N_15756,N_15913);
nor U16626 (N_16626,N_15870,N_15637);
nand U16627 (N_16627,N_16059,N_15793);
nand U16628 (N_16628,N_16179,N_15608);
nor U16629 (N_16629,N_15898,N_16126);
or U16630 (N_16630,N_15821,N_15684);
nor U16631 (N_16631,N_15943,N_15920);
nand U16632 (N_16632,N_16049,N_15952);
nand U16633 (N_16633,N_16006,N_16014);
nand U16634 (N_16634,N_15956,N_15664);
nor U16635 (N_16635,N_15849,N_15872);
xnor U16636 (N_16636,N_16122,N_15990);
nand U16637 (N_16637,N_15682,N_16035);
and U16638 (N_16638,N_16106,N_16115);
or U16639 (N_16639,N_16133,N_16053);
nand U16640 (N_16640,N_15728,N_16187);
or U16641 (N_16641,N_16192,N_15934);
and U16642 (N_16642,N_16016,N_16132);
and U16643 (N_16643,N_16111,N_16064);
xor U16644 (N_16644,N_15933,N_15676);
nand U16645 (N_16645,N_15860,N_16131);
nor U16646 (N_16646,N_15832,N_15654);
nand U16647 (N_16647,N_16016,N_16082);
or U16648 (N_16648,N_15705,N_15642);
nor U16649 (N_16649,N_15632,N_15636);
nand U16650 (N_16650,N_15734,N_15654);
or U16651 (N_16651,N_15983,N_16144);
nor U16652 (N_16652,N_16109,N_16184);
nand U16653 (N_16653,N_15909,N_16181);
nand U16654 (N_16654,N_15986,N_15736);
or U16655 (N_16655,N_16076,N_15758);
nor U16656 (N_16656,N_15940,N_15763);
nor U16657 (N_16657,N_16119,N_16094);
nor U16658 (N_16658,N_15866,N_15783);
nor U16659 (N_16659,N_16152,N_15760);
or U16660 (N_16660,N_15947,N_16129);
or U16661 (N_16661,N_15649,N_15994);
or U16662 (N_16662,N_15655,N_15806);
xor U16663 (N_16663,N_15672,N_15991);
nor U16664 (N_16664,N_15662,N_15669);
or U16665 (N_16665,N_16181,N_15734);
nand U16666 (N_16666,N_16006,N_15766);
nor U16667 (N_16667,N_15758,N_15912);
or U16668 (N_16668,N_15814,N_15616);
nand U16669 (N_16669,N_15614,N_15804);
and U16670 (N_16670,N_15650,N_15950);
nand U16671 (N_16671,N_15961,N_15819);
nor U16672 (N_16672,N_16113,N_15942);
nand U16673 (N_16673,N_15820,N_15924);
and U16674 (N_16674,N_15985,N_16048);
nand U16675 (N_16675,N_15676,N_15791);
nand U16676 (N_16676,N_16094,N_15857);
and U16677 (N_16677,N_15602,N_15657);
and U16678 (N_16678,N_15675,N_15743);
nor U16679 (N_16679,N_15934,N_15750);
and U16680 (N_16680,N_15613,N_15664);
or U16681 (N_16681,N_15804,N_16104);
nand U16682 (N_16682,N_15940,N_15617);
or U16683 (N_16683,N_15949,N_15831);
nor U16684 (N_16684,N_16125,N_16128);
or U16685 (N_16685,N_15631,N_15950);
xnor U16686 (N_16686,N_15762,N_16157);
or U16687 (N_16687,N_15818,N_16004);
nand U16688 (N_16688,N_15955,N_16196);
or U16689 (N_16689,N_16128,N_15850);
nor U16690 (N_16690,N_15678,N_16160);
nand U16691 (N_16691,N_15905,N_16143);
nor U16692 (N_16692,N_15831,N_16147);
or U16693 (N_16693,N_15888,N_16164);
xnor U16694 (N_16694,N_16198,N_15940);
or U16695 (N_16695,N_15909,N_16106);
or U16696 (N_16696,N_16118,N_16179);
nand U16697 (N_16697,N_16057,N_16176);
nand U16698 (N_16698,N_15610,N_15764);
nand U16699 (N_16699,N_15652,N_15762);
and U16700 (N_16700,N_15834,N_15897);
nor U16701 (N_16701,N_16180,N_15772);
xnor U16702 (N_16702,N_16100,N_16125);
nor U16703 (N_16703,N_16075,N_16134);
or U16704 (N_16704,N_15787,N_16061);
or U16705 (N_16705,N_16075,N_15667);
xnor U16706 (N_16706,N_16175,N_16008);
nor U16707 (N_16707,N_15750,N_15762);
or U16708 (N_16708,N_16120,N_16080);
nand U16709 (N_16709,N_15804,N_15760);
and U16710 (N_16710,N_15697,N_15931);
nor U16711 (N_16711,N_15609,N_16135);
or U16712 (N_16712,N_15735,N_15932);
or U16713 (N_16713,N_16020,N_15863);
and U16714 (N_16714,N_15618,N_15888);
and U16715 (N_16715,N_15662,N_16188);
nand U16716 (N_16716,N_15892,N_15645);
and U16717 (N_16717,N_16083,N_15626);
nor U16718 (N_16718,N_15691,N_15804);
nor U16719 (N_16719,N_15875,N_16174);
nand U16720 (N_16720,N_15851,N_15919);
nor U16721 (N_16721,N_15617,N_15734);
and U16722 (N_16722,N_15644,N_15834);
and U16723 (N_16723,N_16188,N_15873);
and U16724 (N_16724,N_16036,N_15850);
and U16725 (N_16725,N_15876,N_15854);
or U16726 (N_16726,N_15700,N_15930);
and U16727 (N_16727,N_16051,N_15600);
nor U16728 (N_16728,N_15951,N_15830);
and U16729 (N_16729,N_15802,N_15692);
xor U16730 (N_16730,N_16054,N_16074);
and U16731 (N_16731,N_16192,N_15735);
or U16732 (N_16732,N_15989,N_15839);
and U16733 (N_16733,N_15987,N_15716);
nor U16734 (N_16734,N_15839,N_16044);
nor U16735 (N_16735,N_15670,N_16007);
or U16736 (N_16736,N_15675,N_15853);
nand U16737 (N_16737,N_15799,N_15940);
xnor U16738 (N_16738,N_15902,N_15731);
or U16739 (N_16739,N_16085,N_15791);
nor U16740 (N_16740,N_15792,N_16116);
nor U16741 (N_16741,N_15941,N_16000);
nand U16742 (N_16742,N_15662,N_16149);
nor U16743 (N_16743,N_15878,N_15648);
nor U16744 (N_16744,N_15613,N_16115);
nand U16745 (N_16745,N_15835,N_15776);
xor U16746 (N_16746,N_15920,N_15834);
or U16747 (N_16747,N_15975,N_16197);
or U16748 (N_16748,N_15924,N_15819);
and U16749 (N_16749,N_15904,N_16038);
nand U16750 (N_16750,N_15602,N_15901);
or U16751 (N_16751,N_15970,N_15855);
nor U16752 (N_16752,N_16192,N_16181);
and U16753 (N_16753,N_16144,N_15648);
and U16754 (N_16754,N_15617,N_15914);
nor U16755 (N_16755,N_16010,N_15882);
or U16756 (N_16756,N_15845,N_16182);
nand U16757 (N_16757,N_15798,N_15724);
nor U16758 (N_16758,N_16008,N_15710);
and U16759 (N_16759,N_15965,N_15614);
and U16760 (N_16760,N_16157,N_15895);
nand U16761 (N_16761,N_15943,N_15877);
and U16762 (N_16762,N_16000,N_16004);
or U16763 (N_16763,N_16032,N_15695);
nand U16764 (N_16764,N_15756,N_15801);
and U16765 (N_16765,N_15676,N_16045);
nand U16766 (N_16766,N_16007,N_15737);
nand U16767 (N_16767,N_16145,N_15747);
nor U16768 (N_16768,N_15871,N_15733);
nor U16769 (N_16769,N_15878,N_16107);
nor U16770 (N_16770,N_15624,N_16197);
and U16771 (N_16771,N_15814,N_16013);
nor U16772 (N_16772,N_15779,N_15958);
xor U16773 (N_16773,N_15782,N_16185);
and U16774 (N_16774,N_15623,N_15797);
nand U16775 (N_16775,N_15981,N_15925);
and U16776 (N_16776,N_16140,N_15775);
and U16777 (N_16777,N_15604,N_15648);
nand U16778 (N_16778,N_15965,N_16168);
and U16779 (N_16779,N_15730,N_15707);
or U16780 (N_16780,N_15614,N_15708);
or U16781 (N_16781,N_15833,N_15700);
or U16782 (N_16782,N_15970,N_15991);
or U16783 (N_16783,N_16161,N_16014);
nor U16784 (N_16784,N_15731,N_16157);
nand U16785 (N_16785,N_16158,N_15848);
or U16786 (N_16786,N_15756,N_15733);
or U16787 (N_16787,N_16175,N_15642);
nand U16788 (N_16788,N_15844,N_15774);
or U16789 (N_16789,N_15791,N_15815);
nand U16790 (N_16790,N_15958,N_15839);
or U16791 (N_16791,N_16132,N_15825);
and U16792 (N_16792,N_16075,N_15957);
nor U16793 (N_16793,N_16096,N_15845);
and U16794 (N_16794,N_15605,N_15984);
and U16795 (N_16795,N_15653,N_15796);
and U16796 (N_16796,N_15932,N_15613);
or U16797 (N_16797,N_15881,N_16161);
and U16798 (N_16798,N_15881,N_15992);
nor U16799 (N_16799,N_15729,N_16035);
nand U16800 (N_16800,N_16676,N_16463);
and U16801 (N_16801,N_16765,N_16318);
or U16802 (N_16802,N_16624,N_16430);
nor U16803 (N_16803,N_16670,N_16791);
nand U16804 (N_16804,N_16393,N_16326);
or U16805 (N_16805,N_16209,N_16606);
nand U16806 (N_16806,N_16271,N_16353);
or U16807 (N_16807,N_16493,N_16457);
and U16808 (N_16808,N_16614,N_16354);
and U16809 (N_16809,N_16520,N_16277);
nand U16810 (N_16810,N_16434,N_16369);
nand U16811 (N_16811,N_16554,N_16748);
or U16812 (N_16812,N_16729,N_16545);
and U16813 (N_16813,N_16320,N_16695);
nor U16814 (N_16814,N_16527,N_16404);
nand U16815 (N_16815,N_16462,N_16469);
nand U16816 (N_16816,N_16645,N_16665);
or U16817 (N_16817,N_16454,N_16505);
nand U16818 (N_16818,N_16339,N_16573);
nand U16819 (N_16819,N_16452,N_16661);
or U16820 (N_16820,N_16641,N_16411);
or U16821 (N_16821,N_16262,N_16567);
nor U16822 (N_16822,N_16747,N_16337);
or U16823 (N_16823,N_16403,N_16479);
or U16824 (N_16824,N_16544,N_16599);
nor U16825 (N_16825,N_16701,N_16364);
and U16826 (N_16826,N_16443,N_16475);
or U16827 (N_16827,N_16540,N_16564);
and U16828 (N_16828,N_16603,N_16276);
nor U16829 (N_16829,N_16588,N_16553);
and U16830 (N_16830,N_16572,N_16459);
and U16831 (N_16831,N_16223,N_16472);
and U16832 (N_16832,N_16466,N_16626);
nor U16833 (N_16833,N_16376,N_16696);
and U16834 (N_16834,N_16694,N_16655);
nor U16835 (N_16835,N_16391,N_16287);
or U16836 (N_16836,N_16292,N_16372);
or U16837 (N_16837,N_16733,N_16557);
and U16838 (N_16838,N_16448,N_16321);
nand U16839 (N_16839,N_16640,N_16525);
nand U16840 (N_16840,N_16647,N_16332);
and U16841 (N_16841,N_16504,N_16771);
nor U16842 (N_16842,N_16598,N_16489);
or U16843 (N_16843,N_16619,N_16220);
or U16844 (N_16844,N_16308,N_16461);
nor U16845 (N_16845,N_16618,N_16421);
nor U16846 (N_16846,N_16286,N_16345);
or U16847 (N_16847,N_16232,N_16713);
nor U16848 (N_16848,N_16428,N_16724);
and U16849 (N_16849,N_16392,N_16431);
nand U16850 (N_16850,N_16578,N_16638);
nand U16851 (N_16851,N_16280,N_16485);
or U16852 (N_16852,N_16705,N_16565);
nand U16853 (N_16853,N_16203,N_16437);
nand U16854 (N_16854,N_16648,N_16674);
nor U16855 (N_16855,N_16248,N_16615);
xnor U16856 (N_16856,N_16290,N_16478);
nor U16857 (N_16857,N_16390,N_16241);
xor U16858 (N_16858,N_16324,N_16570);
or U16859 (N_16859,N_16215,N_16343);
and U16860 (N_16860,N_16759,N_16338);
or U16861 (N_16861,N_16418,N_16651);
nand U16862 (N_16862,N_16245,N_16779);
nand U16863 (N_16863,N_16726,N_16703);
or U16864 (N_16864,N_16356,N_16377);
xor U16865 (N_16865,N_16427,N_16507);
nand U16866 (N_16866,N_16758,N_16467);
and U16867 (N_16867,N_16219,N_16658);
nor U16868 (N_16868,N_16274,N_16438);
nand U16869 (N_16869,N_16789,N_16228);
and U16870 (N_16870,N_16208,N_16742);
nand U16871 (N_16871,N_16798,N_16582);
nand U16872 (N_16872,N_16494,N_16576);
nor U16873 (N_16873,N_16351,N_16200);
and U16874 (N_16874,N_16601,N_16600);
nand U16875 (N_16875,N_16387,N_16773);
and U16876 (N_16876,N_16777,N_16562);
and U16877 (N_16877,N_16768,N_16442);
or U16878 (N_16878,N_16796,N_16301);
nor U16879 (N_16879,N_16649,N_16378);
or U16880 (N_16880,N_16566,N_16218);
or U16881 (N_16881,N_16639,N_16523);
or U16882 (N_16882,N_16365,N_16293);
nand U16883 (N_16883,N_16445,N_16756);
nand U16884 (N_16884,N_16451,N_16312);
and U16885 (N_16885,N_16456,N_16363);
or U16886 (N_16886,N_16741,N_16333);
or U16887 (N_16887,N_16263,N_16737);
nor U16888 (N_16888,N_16305,N_16740);
and U16889 (N_16889,N_16613,N_16233);
nor U16890 (N_16890,N_16374,N_16336);
and U16891 (N_16891,N_16715,N_16652);
nor U16892 (N_16892,N_16323,N_16636);
or U16893 (N_16893,N_16357,N_16691);
nand U16894 (N_16894,N_16447,N_16348);
xnor U16895 (N_16895,N_16420,N_16731);
nand U16896 (N_16896,N_16524,N_16628);
nor U16897 (N_16897,N_16531,N_16528);
and U16898 (N_16898,N_16304,N_16563);
nand U16899 (N_16899,N_16385,N_16782);
nand U16900 (N_16900,N_16744,N_16711);
or U16901 (N_16901,N_16642,N_16739);
or U16902 (N_16902,N_16587,N_16379);
nand U16903 (N_16903,N_16416,N_16723);
nor U16904 (N_16904,N_16269,N_16755);
or U16905 (N_16905,N_16264,N_16571);
or U16906 (N_16906,N_16380,N_16552);
or U16907 (N_16907,N_16498,N_16368);
or U16908 (N_16908,N_16240,N_16714);
nor U16909 (N_16909,N_16707,N_16201);
nand U16910 (N_16910,N_16797,N_16311);
nand U16911 (N_16911,N_16397,N_16327);
nor U16912 (N_16912,N_16586,N_16684);
nor U16913 (N_16913,N_16346,N_16322);
and U16914 (N_16914,N_16629,N_16254);
or U16915 (N_16915,N_16202,N_16754);
nand U16916 (N_16916,N_16272,N_16699);
nand U16917 (N_16917,N_16222,N_16560);
xnor U16918 (N_16918,N_16298,N_16558);
and U16919 (N_16919,N_16488,N_16687);
nor U16920 (N_16920,N_16750,N_16384);
nand U16921 (N_16921,N_16307,N_16501);
and U16922 (N_16922,N_16410,N_16712);
nand U16923 (N_16923,N_16730,N_16362);
nor U16924 (N_16924,N_16704,N_16500);
or U16925 (N_16925,N_16518,N_16511);
and U16926 (N_16926,N_16584,N_16611);
nand U16927 (N_16927,N_16671,N_16444);
nor U16928 (N_16928,N_16602,N_16604);
nand U16929 (N_16929,N_16289,N_16697);
nor U16930 (N_16930,N_16270,N_16361);
nand U16931 (N_16931,N_16236,N_16516);
and U16932 (N_16932,N_16266,N_16722);
nor U16933 (N_16933,N_16784,N_16743);
nor U16934 (N_16934,N_16482,N_16440);
or U16935 (N_16935,N_16646,N_16621);
and U16936 (N_16936,N_16344,N_16710);
nor U16937 (N_16937,N_16660,N_16519);
or U16938 (N_16938,N_16590,N_16745);
or U16939 (N_16939,N_16788,N_16347);
nand U16940 (N_16940,N_16595,N_16609);
or U16941 (N_16941,N_16279,N_16213);
and U16942 (N_16942,N_16718,N_16546);
and U16943 (N_16943,N_16429,N_16751);
nor U16944 (N_16944,N_16306,N_16281);
xnor U16945 (N_16945,N_16341,N_16550);
or U16946 (N_16946,N_16794,N_16529);
or U16947 (N_16947,N_16559,N_16650);
or U16948 (N_16948,N_16439,N_16698);
nor U16949 (N_16949,N_16772,N_16253);
nor U16950 (N_16950,N_16468,N_16762);
nand U16951 (N_16951,N_16453,N_16503);
or U16952 (N_16952,N_16473,N_16366);
nand U16953 (N_16953,N_16792,N_16217);
or U16954 (N_16954,N_16388,N_16549);
nand U16955 (N_16955,N_16734,N_16334);
nand U16956 (N_16956,N_16373,N_16725);
nor U16957 (N_16957,N_16409,N_16594);
nand U16958 (N_16958,N_16294,N_16367);
and U16959 (N_16959,N_16465,N_16335);
nand U16960 (N_16960,N_16486,N_16631);
nand U16961 (N_16961,N_16719,N_16510);
nor U16962 (N_16962,N_16763,N_16764);
nor U16963 (N_16963,N_16425,N_16408);
or U16964 (N_16964,N_16314,N_16688);
nor U16965 (N_16965,N_16477,N_16288);
nor U16966 (N_16966,N_16548,N_16370);
or U16967 (N_16967,N_16689,N_16535);
and U16968 (N_16968,N_16593,N_16786);
nand U16969 (N_16969,N_16291,N_16799);
and U16970 (N_16970,N_16358,N_16679);
or U16971 (N_16971,N_16303,N_16580);
nor U16972 (N_16972,N_16605,N_16533);
and U16973 (N_16973,N_16246,N_16746);
nor U16974 (N_16974,N_16250,N_16783);
or U16975 (N_16975,N_16455,N_16449);
or U16976 (N_16976,N_16412,N_16513);
or U16977 (N_16977,N_16583,N_16749);
or U16978 (N_16978,N_16686,N_16426);
nor U16979 (N_16979,N_16706,N_16702);
nand U16980 (N_16980,N_16591,N_16608);
or U16981 (N_16981,N_16417,N_16677);
nand U16982 (N_16982,N_16774,N_16669);
nand U16983 (N_16983,N_16781,N_16509);
or U16984 (N_16984,N_16278,N_16212);
xor U16985 (N_16985,N_16753,N_16683);
and U16986 (N_16986,N_16654,N_16766);
and U16987 (N_16987,N_16476,N_16775);
nand U16988 (N_16988,N_16526,N_16574);
or U16989 (N_16989,N_16487,N_16414);
and U16990 (N_16990,N_16752,N_16508);
or U16991 (N_16991,N_16389,N_16675);
or U16992 (N_16992,N_16625,N_16300);
nor U16993 (N_16993,N_16506,N_16319);
or U16994 (N_16994,N_16672,N_16204);
or U16995 (N_16995,N_16585,N_16235);
and U16996 (N_16996,N_16350,N_16207);
or U16997 (N_16997,N_16709,N_16268);
and U16998 (N_16998,N_16716,N_16433);
nand U16999 (N_16999,N_16653,N_16496);
and U17000 (N_17000,N_16568,N_16721);
nand U17001 (N_17001,N_16757,N_16259);
nand U17002 (N_17002,N_16371,N_16537);
and U17003 (N_17003,N_16577,N_16302);
nor U17004 (N_17004,N_16732,N_16261);
and U17005 (N_17005,N_16678,N_16239);
and U17006 (N_17006,N_16682,N_16728);
and U17007 (N_17007,N_16407,N_16446);
nand U17008 (N_17008,N_16483,N_16258);
nor U17009 (N_17009,N_16230,N_16395);
nor U17010 (N_17010,N_16243,N_16521);
nand U17011 (N_17011,N_16539,N_16785);
nor U17012 (N_17012,N_16382,N_16330);
nor U17013 (N_17013,N_16205,N_16252);
nand U17014 (N_17014,N_16795,N_16666);
nand U17015 (N_17015,N_16267,N_16355);
nand U17016 (N_17016,N_16659,N_16257);
nand U17017 (N_17017,N_16470,N_16579);
nand U17018 (N_17018,N_16441,N_16490);
and U17019 (N_17019,N_16386,N_16597);
or U17020 (N_17020,N_16592,N_16667);
nand U17021 (N_17021,N_16299,N_16681);
nor U17022 (N_17022,N_16673,N_16657);
nand U17023 (N_17023,N_16422,N_16708);
or U17024 (N_17024,N_16260,N_16249);
nand U17025 (N_17025,N_16575,N_16360);
and U17026 (N_17026,N_16242,N_16406);
nor U17027 (N_17027,N_16297,N_16396);
nand U17028 (N_17028,N_16402,N_16325);
nand U17029 (N_17029,N_16538,N_16315);
or U17030 (N_17030,N_16225,N_16282);
nor U17031 (N_17031,N_16760,N_16787);
and U17032 (N_17032,N_16329,N_16480);
or U17033 (N_17033,N_16484,N_16761);
nand U17034 (N_17034,N_16664,N_16491);
and U17035 (N_17035,N_16663,N_16342);
and U17036 (N_17036,N_16778,N_16214);
nand U17037 (N_17037,N_16690,N_16275);
and U17038 (N_17038,N_16569,N_16229);
nand U17039 (N_17039,N_16512,N_16502);
and U17040 (N_17040,N_16394,N_16635);
nor U17041 (N_17041,N_16283,N_16770);
and U17042 (N_17042,N_16295,N_16693);
and U17043 (N_17043,N_16405,N_16541);
and U17044 (N_17044,N_16244,N_16432);
nand U17045 (N_17045,N_16623,N_16692);
or U17046 (N_17046,N_16617,N_16555);
nor U17047 (N_17047,N_16551,N_16514);
nand U17048 (N_17048,N_16612,N_16727);
nor U17049 (N_17049,N_16596,N_16359);
nor U17050 (N_17050,N_16206,N_16450);
or U17051 (N_17051,N_16227,N_16530);
or U17052 (N_17052,N_16460,N_16399);
or U17053 (N_17053,N_16481,N_16738);
nor U17054 (N_17054,N_16221,N_16309);
or U17055 (N_17055,N_16637,N_16400);
and U17056 (N_17056,N_16284,N_16375);
or U17057 (N_17057,N_16622,N_16216);
xor U17058 (N_17058,N_16536,N_16471);
and U17059 (N_17059,N_16720,N_16401);
or U17060 (N_17060,N_16328,N_16662);
nor U17061 (N_17061,N_16668,N_16340);
and U17062 (N_17062,N_16735,N_16464);
or U17063 (N_17063,N_16607,N_16310);
and U17064 (N_17064,N_16780,N_16620);
or U17065 (N_17065,N_16685,N_16643);
or U17066 (N_17066,N_16769,N_16633);
and U17067 (N_17067,N_16352,N_16331);
and U17068 (N_17068,N_16316,N_16383);
and U17069 (N_17069,N_16237,N_16542);
or U17070 (N_17070,N_16522,N_16210);
and U17071 (N_17071,N_16255,N_16265);
nand U17072 (N_17072,N_16644,N_16543);
nor U17073 (N_17073,N_16313,N_16436);
nor U17074 (N_17074,N_16517,N_16767);
and U17075 (N_17075,N_16790,N_16458);
and U17076 (N_17076,N_16634,N_16231);
and U17077 (N_17077,N_16656,N_16616);
or U17078 (N_17078,N_16700,N_16413);
and U17079 (N_17079,N_16561,N_16680);
and U17080 (N_17080,N_16581,N_16497);
and U17081 (N_17081,N_16349,N_16556);
nor U17082 (N_17082,N_16630,N_16515);
nand U17083 (N_17083,N_16398,N_16296);
nand U17084 (N_17084,N_16589,N_16423);
or U17085 (N_17085,N_16211,N_16736);
and U17086 (N_17086,N_16499,N_16793);
nand U17087 (N_17087,N_16224,N_16547);
or U17088 (N_17088,N_16273,N_16317);
nand U17089 (N_17089,N_16532,N_16474);
and U17090 (N_17090,N_16424,N_16534);
nor U17091 (N_17091,N_16226,N_16419);
nor U17092 (N_17092,N_16251,N_16627);
nand U17093 (N_17093,N_16632,N_16610);
or U17094 (N_17094,N_16495,N_16776);
nor U17095 (N_17095,N_16717,N_16381);
and U17096 (N_17096,N_16247,N_16256);
or U17097 (N_17097,N_16234,N_16492);
or U17098 (N_17098,N_16435,N_16415);
and U17099 (N_17099,N_16285,N_16238);
and U17100 (N_17100,N_16746,N_16799);
or U17101 (N_17101,N_16607,N_16337);
and U17102 (N_17102,N_16798,N_16224);
nor U17103 (N_17103,N_16381,N_16770);
or U17104 (N_17104,N_16595,N_16785);
nand U17105 (N_17105,N_16438,N_16721);
and U17106 (N_17106,N_16260,N_16697);
and U17107 (N_17107,N_16369,N_16511);
and U17108 (N_17108,N_16587,N_16284);
nand U17109 (N_17109,N_16759,N_16522);
nand U17110 (N_17110,N_16342,N_16577);
or U17111 (N_17111,N_16369,N_16762);
nor U17112 (N_17112,N_16224,N_16729);
nor U17113 (N_17113,N_16560,N_16451);
and U17114 (N_17114,N_16266,N_16629);
and U17115 (N_17115,N_16778,N_16223);
or U17116 (N_17116,N_16349,N_16289);
nor U17117 (N_17117,N_16376,N_16560);
nor U17118 (N_17118,N_16640,N_16470);
nor U17119 (N_17119,N_16254,N_16247);
or U17120 (N_17120,N_16608,N_16427);
or U17121 (N_17121,N_16516,N_16257);
and U17122 (N_17122,N_16638,N_16672);
nor U17123 (N_17123,N_16227,N_16598);
or U17124 (N_17124,N_16648,N_16447);
and U17125 (N_17125,N_16521,N_16688);
and U17126 (N_17126,N_16259,N_16392);
or U17127 (N_17127,N_16548,N_16216);
nor U17128 (N_17128,N_16608,N_16606);
nand U17129 (N_17129,N_16787,N_16601);
or U17130 (N_17130,N_16726,N_16210);
or U17131 (N_17131,N_16403,N_16778);
nand U17132 (N_17132,N_16462,N_16261);
nor U17133 (N_17133,N_16412,N_16543);
or U17134 (N_17134,N_16468,N_16428);
or U17135 (N_17135,N_16550,N_16661);
or U17136 (N_17136,N_16691,N_16260);
and U17137 (N_17137,N_16396,N_16370);
nor U17138 (N_17138,N_16636,N_16781);
nor U17139 (N_17139,N_16730,N_16363);
and U17140 (N_17140,N_16733,N_16252);
nor U17141 (N_17141,N_16393,N_16380);
and U17142 (N_17142,N_16300,N_16659);
nor U17143 (N_17143,N_16302,N_16460);
xnor U17144 (N_17144,N_16698,N_16555);
or U17145 (N_17145,N_16643,N_16651);
and U17146 (N_17146,N_16325,N_16412);
or U17147 (N_17147,N_16602,N_16505);
xor U17148 (N_17148,N_16488,N_16422);
nor U17149 (N_17149,N_16258,N_16712);
nor U17150 (N_17150,N_16211,N_16582);
nand U17151 (N_17151,N_16638,N_16720);
or U17152 (N_17152,N_16785,N_16668);
nor U17153 (N_17153,N_16582,N_16479);
and U17154 (N_17154,N_16493,N_16365);
nand U17155 (N_17155,N_16254,N_16232);
nor U17156 (N_17156,N_16387,N_16416);
xor U17157 (N_17157,N_16509,N_16376);
nand U17158 (N_17158,N_16411,N_16757);
nand U17159 (N_17159,N_16614,N_16521);
or U17160 (N_17160,N_16609,N_16246);
nand U17161 (N_17161,N_16246,N_16350);
nor U17162 (N_17162,N_16604,N_16234);
nand U17163 (N_17163,N_16208,N_16664);
nand U17164 (N_17164,N_16400,N_16279);
nor U17165 (N_17165,N_16629,N_16510);
nand U17166 (N_17166,N_16565,N_16762);
and U17167 (N_17167,N_16449,N_16390);
and U17168 (N_17168,N_16551,N_16521);
and U17169 (N_17169,N_16676,N_16464);
nand U17170 (N_17170,N_16752,N_16463);
nand U17171 (N_17171,N_16433,N_16540);
nand U17172 (N_17172,N_16710,N_16282);
or U17173 (N_17173,N_16279,N_16538);
and U17174 (N_17174,N_16525,N_16347);
nand U17175 (N_17175,N_16312,N_16564);
and U17176 (N_17176,N_16320,N_16273);
and U17177 (N_17177,N_16488,N_16683);
or U17178 (N_17178,N_16616,N_16378);
nor U17179 (N_17179,N_16634,N_16348);
or U17180 (N_17180,N_16600,N_16473);
nand U17181 (N_17181,N_16231,N_16414);
and U17182 (N_17182,N_16347,N_16697);
and U17183 (N_17183,N_16226,N_16672);
nand U17184 (N_17184,N_16596,N_16717);
nor U17185 (N_17185,N_16567,N_16524);
nor U17186 (N_17186,N_16552,N_16259);
or U17187 (N_17187,N_16593,N_16462);
or U17188 (N_17188,N_16351,N_16508);
or U17189 (N_17189,N_16722,N_16774);
and U17190 (N_17190,N_16530,N_16535);
and U17191 (N_17191,N_16473,N_16736);
nor U17192 (N_17192,N_16658,N_16336);
nand U17193 (N_17193,N_16545,N_16632);
and U17194 (N_17194,N_16333,N_16575);
and U17195 (N_17195,N_16704,N_16329);
or U17196 (N_17196,N_16540,N_16792);
nand U17197 (N_17197,N_16292,N_16278);
or U17198 (N_17198,N_16774,N_16393);
or U17199 (N_17199,N_16586,N_16278);
or U17200 (N_17200,N_16543,N_16634);
nand U17201 (N_17201,N_16328,N_16422);
or U17202 (N_17202,N_16798,N_16511);
nand U17203 (N_17203,N_16718,N_16626);
or U17204 (N_17204,N_16708,N_16207);
and U17205 (N_17205,N_16533,N_16489);
nor U17206 (N_17206,N_16397,N_16480);
and U17207 (N_17207,N_16338,N_16445);
nor U17208 (N_17208,N_16670,N_16615);
nor U17209 (N_17209,N_16773,N_16675);
nor U17210 (N_17210,N_16224,N_16653);
xor U17211 (N_17211,N_16765,N_16705);
nand U17212 (N_17212,N_16308,N_16770);
nand U17213 (N_17213,N_16692,N_16619);
nand U17214 (N_17214,N_16703,N_16292);
nor U17215 (N_17215,N_16709,N_16394);
nand U17216 (N_17216,N_16728,N_16310);
nand U17217 (N_17217,N_16217,N_16691);
or U17218 (N_17218,N_16517,N_16751);
nor U17219 (N_17219,N_16397,N_16646);
and U17220 (N_17220,N_16649,N_16673);
and U17221 (N_17221,N_16216,N_16634);
nor U17222 (N_17222,N_16271,N_16658);
nand U17223 (N_17223,N_16496,N_16229);
nor U17224 (N_17224,N_16745,N_16506);
and U17225 (N_17225,N_16634,N_16292);
and U17226 (N_17226,N_16770,N_16787);
or U17227 (N_17227,N_16407,N_16747);
nand U17228 (N_17228,N_16392,N_16508);
or U17229 (N_17229,N_16311,N_16663);
or U17230 (N_17230,N_16526,N_16661);
nor U17231 (N_17231,N_16553,N_16694);
xor U17232 (N_17232,N_16651,N_16645);
or U17233 (N_17233,N_16616,N_16344);
nand U17234 (N_17234,N_16790,N_16643);
xor U17235 (N_17235,N_16226,N_16327);
nand U17236 (N_17236,N_16624,N_16476);
nand U17237 (N_17237,N_16773,N_16578);
nor U17238 (N_17238,N_16240,N_16609);
nand U17239 (N_17239,N_16343,N_16686);
and U17240 (N_17240,N_16478,N_16411);
or U17241 (N_17241,N_16601,N_16262);
or U17242 (N_17242,N_16669,N_16466);
and U17243 (N_17243,N_16587,N_16644);
nor U17244 (N_17244,N_16651,N_16510);
nand U17245 (N_17245,N_16615,N_16707);
and U17246 (N_17246,N_16229,N_16761);
and U17247 (N_17247,N_16551,N_16312);
and U17248 (N_17248,N_16664,N_16337);
and U17249 (N_17249,N_16345,N_16664);
nand U17250 (N_17250,N_16579,N_16522);
nor U17251 (N_17251,N_16380,N_16250);
nor U17252 (N_17252,N_16747,N_16262);
nand U17253 (N_17253,N_16667,N_16717);
nor U17254 (N_17254,N_16670,N_16408);
and U17255 (N_17255,N_16792,N_16349);
nor U17256 (N_17256,N_16536,N_16438);
nand U17257 (N_17257,N_16635,N_16245);
nand U17258 (N_17258,N_16572,N_16763);
or U17259 (N_17259,N_16378,N_16215);
or U17260 (N_17260,N_16479,N_16707);
or U17261 (N_17261,N_16475,N_16650);
or U17262 (N_17262,N_16293,N_16329);
nor U17263 (N_17263,N_16340,N_16510);
or U17264 (N_17264,N_16317,N_16380);
and U17265 (N_17265,N_16689,N_16678);
and U17266 (N_17266,N_16334,N_16748);
xor U17267 (N_17267,N_16403,N_16747);
nand U17268 (N_17268,N_16545,N_16533);
nor U17269 (N_17269,N_16418,N_16417);
and U17270 (N_17270,N_16347,N_16640);
and U17271 (N_17271,N_16666,N_16270);
and U17272 (N_17272,N_16365,N_16353);
or U17273 (N_17273,N_16700,N_16666);
nand U17274 (N_17274,N_16475,N_16689);
and U17275 (N_17275,N_16496,N_16288);
and U17276 (N_17276,N_16276,N_16444);
or U17277 (N_17277,N_16442,N_16327);
or U17278 (N_17278,N_16554,N_16340);
nor U17279 (N_17279,N_16405,N_16754);
or U17280 (N_17280,N_16276,N_16711);
nor U17281 (N_17281,N_16586,N_16620);
nand U17282 (N_17282,N_16234,N_16655);
or U17283 (N_17283,N_16695,N_16372);
or U17284 (N_17284,N_16533,N_16477);
and U17285 (N_17285,N_16463,N_16391);
or U17286 (N_17286,N_16334,N_16428);
nor U17287 (N_17287,N_16768,N_16202);
nor U17288 (N_17288,N_16646,N_16317);
or U17289 (N_17289,N_16440,N_16539);
nor U17290 (N_17290,N_16237,N_16309);
and U17291 (N_17291,N_16557,N_16716);
nand U17292 (N_17292,N_16772,N_16636);
and U17293 (N_17293,N_16355,N_16558);
nand U17294 (N_17294,N_16379,N_16499);
or U17295 (N_17295,N_16795,N_16358);
or U17296 (N_17296,N_16593,N_16585);
nand U17297 (N_17297,N_16253,N_16282);
and U17298 (N_17298,N_16274,N_16295);
or U17299 (N_17299,N_16783,N_16655);
or U17300 (N_17300,N_16699,N_16560);
xor U17301 (N_17301,N_16253,N_16494);
nor U17302 (N_17302,N_16588,N_16792);
and U17303 (N_17303,N_16542,N_16413);
nor U17304 (N_17304,N_16546,N_16450);
nand U17305 (N_17305,N_16300,N_16787);
or U17306 (N_17306,N_16697,N_16759);
nor U17307 (N_17307,N_16689,N_16400);
nand U17308 (N_17308,N_16692,N_16700);
nand U17309 (N_17309,N_16424,N_16391);
nand U17310 (N_17310,N_16425,N_16781);
nand U17311 (N_17311,N_16390,N_16443);
or U17312 (N_17312,N_16661,N_16786);
nand U17313 (N_17313,N_16414,N_16476);
nor U17314 (N_17314,N_16362,N_16637);
and U17315 (N_17315,N_16284,N_16603);
nand U17316 (N_17316,N_16426,N_16619);
and U17317 (N_17317,N_16683,N_16370);
xnor U17318 (N_17318,N_16672,N_16239);
and U17319 (N_17319,N_16798,N_16592);
and U17320 (N_17320,N_16666,N_16442);
nand U17321 (N_17321,N_16564,N_16243);
xor U17322 (N_17322,N_16579,N_16334);
nand U17323 (N_17323,N_16224,N_16540);
nand U17324 (N_17324,N_16719,N_16451);
nand U17325 (N_17325,N_16417,N_16743);
or U17326 (N_17326,N_16345,N_16598);
nand U17327 (N_17327,N_16298,N_16582);
and U17328 (N_17328,N_16259,N_16456);
and U17329 (N_17329,N_16648,N_16343);
nor U17330 (N_17330,N_16396,N_16708);
nor U17331 (N_17331,N_16529,N_16375);
and U17332 (N_17332,N_16596,N_16518);
and U17333 (N_17333,N_16772,N_16324);
nand U17334 (N_17334,N_16780,N_16698);
nor U17335 (N_17335,N_16415,N_16635);
nor U17336 (N_17336,N_16330,N_16443);
nor U17337 (N_17337,N_16728,N_16441);
and U17338 (N_17338,N_16220,N_16457);
or U17339 (N_17339,N_16596,N_16239);
nand U17340 (N_17340,N_16712,N_16284);
nand U17341 (N_17341,N_16223,N_16400);
and U17342 (N_17342,N_16627,N_16404);
and U17343 (N_17343,N_16471,N_16299);
nor U17344 (N_17344,N_16218,N_16262);
nand U17345 (N_17345,N_16319,N_16203);
or U17346 (N_17346,N_16699,N_16717);
and U17347 (N_17347,N_16587,N_16447);
and U17348 (N_17348,N_16581,N_16654);
and U17349 (N_17349,N_16282,N_16236);
nor U17350 (N_17350,N_16797,N_16422);
nor U17351 (N_17351,N_16643,N_16494);
nor U17352 (N_17352,N_16639,N_16552);
nor U17353 (N_17353,N_16346,N_16267);
nor U17354 (N_17354,N_16497,N_16287);
nor U17355 (N_17355,N_16513,N_16470);
and U17356 (N_17356,N_16227,N_16659);
nor U17357 (N_17357,N_16239,N_16392);
or U17358 (N_17358,N_16587,N_16233);
or U17359 (N_17359,N_16307,N_16282);
nor U17360 (N_17360,N_16286,N_16799);
nand U17361 (N_17361,N_16526,N_16488);
nand U17362 (N_17362,N_16756,N_16423);
or U17363 (N_17363,N_16552,N_16515);
and U17364 (N_17364,N_16646,N_16380);
or U17365 (N_17365,N_16671,N_16697);
and U17366 (N_17366,N_16769,N_16462);
and U17367 (N_17367,N_16555,N_16209);
and U17368 (N_17368,N_16666,N_16282);
xnor U17369 (N_17369,N_16534,N_16660);
nor U17370 (N_17370,N_16545,N_16380);
xor U17371 (N_17371,N_16303,N_16310);
nand U17372 (N_17372,N_16365,N_16210);
nor U17373 (N_17373,N_16233,N_16740);
nor U17374 (N_17374,N_16667,N_16599);
nor U17375 (N_17375,N_16691,N_16218);
nand U17376 (N_17376,N_16751,N_16730);
or U17377 (N_17377,N_16403,N_16473);
or U17378 (N_17378,N_16601,N_16472);
nor U17379 (N_17379,N_16390,N_16661);
nor U17380 (N_17380,N_16231,N_16442);
nor U17381 (N_17381,N_16380,N_16686);
and U17382 (N_17382,N_16289,N_16798);
and U17383 (N_17383,N_16359,N_16379);
and U17384 (N_17384,N_16580,N_16793);
nor U17385 (N_17385,N_16217,N_16467);
and U17386 (N_17386,N_16615,N_16797);
nor U17387 (N_17387,N_16615,N_16591);
or U17388 (N_17388,N_16772,N_16226);
nand U17389 (N_17389,N_16501,N_16383);
and U17390 (N_17390,N_16563,N_16533);
nand U17391 (N_17391,N_16340,N_16669);
nor U17392 (N_17392,N_16759,N_16680);
nand U17393 (N_17393,N_16366,N_16456);
or U17394 (N_17394,N_16783,N_16240);
nand U17395 (N_17395,N_16376,N_16768);
and U17396 (N_17396,N_16701,N_16689);
and U17397 (N_17397,N_16743,N_16602);
and U17398 (N_17398,N_16663,N_16599);
xnor U17399 (N_17399,N_16741,N_16677);
or U17400 (N_17400,N_17007,N_17261);
nor U17401 (N_17401,N_16813,N_17016);
and U17402 (N_17402,N_17234,N_16971);
or U17403 (N_17403,N_17282,N_17116);
nor U17404 (N_17404,N_17009,N_17134);
and U17405 (N_17405,N_17080,N_17389);
and U17406 (N_17406,N_17123,N_17191);
or U17407 (N_17407,N_17301,N_17033);
or U17408 (N_17408,N_17373,N_16820);
nand U17409 (N_17409,N_17317,N_17110);
and U17410 (N_17410,N_17018,N_17113);
xnor U17411 (N_17411,N_16948,N_16902);
nor U17412 (N_17412,N_16803,N_17197);
and U17413 (N_17413,N_17241,N_17184);
or U17414 (N_17414,N_17387,N_17199);
and U17415 (N_17415,N_16827,N_17326);
nand U17416 (N_17416,N_16977,N_16976);
and U17417 (N_17417,N_17127,N_17036);
or U17418 (N_17418,N_16967,N_16841);
nor U17419 (N_17419,N_17354,N_17152);
nand U17420 (N_17420,N_17194,N_16887);
nor U17421 (N_17421,N_16915,N_17390);
nand U17422 (N_17422,N_17190,N_17265);
nand U17423 (N_17423,N_17329,N_17256);
nand U17424 (N_17424,N_17132,N_16914);
nor U17425 (N_17425,N_16812,N_16920);
xnor U17426 (N_17426,N_17070,N_16945);
and U17427 (N_17427,N_17114,N_16873);
and U17428 (N_17428,N_17362,N_16933);
or U17429 (N_17429,N_17300,N_17200);
and U17430 (N_17430,N_17124,N_17195);
or U17431 (N_17431,N_16882,N_17082);
nand U17432 (N_17432,N_16996,N_17005);
and U17433 (N_17433,N_17306,N_16900);
nand U17434 (N_17434,N_16935,N_17312);
nor U17435 (N_17435,N_16867,N_17364);
nor U17436 (N_17436,N_17164,N_17183);
and U17437 (N_17437,N_16930,N_16944);
nand U17438 (N_17438,N_17398,N_16905);
xnor U17439 (N_17439,N_17353,N_17271);
nor U17440 (N_17440,N_17231,N_17020);
nor U17441 (N_17441,N_17382,N_17165);
nor U17442 (N_17442,N_16968,N_17103);
nand U17443 (N_17443,N_17055,N_17204);
nand U17444 (N_17444,N_17022,N_17245);
nor U17445 (N_17445,N_16839,N_16868);
nor U17446 (N_17446,N_17085,N_17064);
or U17447 (N_17447,N_17289,N_17276);
nor U17448 (N_17448,N_17159,N_17130);
or U17449 (N_17449,N_16872,N_17324);
nor U17450 (N_17450,N_16907,N_17146);
nand U17451 (N_17451,N_16881,N_16942);
nand U17452 (N_17452,N_16884,N_16831);
nand U17453 (N_17453,N_16940,N_16895);
or U17454 (N_17454,N_17333,N_16891);
xnor U17455 (N_17455,N_17001,N_17313);
nor U17456 (N_17456,N_17102,N_17286);
or U17457 (N_17457,N_17263,N_17338);
and U17458 (N_17458,N_17360,N_17314);
or U17459 (N_17459,N_17088,N_17223);
or U17460 (N_17460,N_17295,N_16848);
nor U17461 (N_17461,N_17210,N_16864);
and U17462 (N_17462,N_17397,N_17267);
and U17463 (N_17463,N_16987,N_17305);
and U17464 (N_17464,N_17322,N_17321);
nand U17465 (N_17465,N_17225,N_16998);
nand U17466 (N_17466,N_17355,N_17066);
or U17467 (N_17467,N_16931,N_16857);
and U17468 (N_17468,N_17140,N_16874);
nor U17469 (N_17469,N_17294,N_16952);
or U17470 (N_17470,N_16893,N_16877);
nor U17471 (N_17471,N_17008,N_17045);
nor U17472 (N_17472,N_16880,N_17094);
and U17473 (N_17473,N_17264,N_17298);
or U17474 (N_17474,N_17266,N_17292);
and U17475 (N_17475,N_16982,N_17077);
xnor U17476 (N_17476,N_16981,N_17028);
and U17477 (N_17477,N_17236,N_17391);
and U17478 (N_17478,N_17073,N_16834);
nand U17479 (N_17479,N_17023,N_17303);
and U17480 (N_17480,N_17219,N_16972);
nand U17481 (N_17481,N_17117,N_17216);
and U17482 (N_17482,N_17034,N_16963);
or U17483 (N_17483,N_17238,N_17273);
nor U17484 (N_17484,N_17148,N_16852);
or U17485 (N_17485,N_17378,N_16853);
or U17486 (N_17486,N_16821,N_17220);
nand U17487 (N_17487,N_17176,N_17125);
nand U17488 (N_17488,N_16883,N_17232);
and U17489 (N_17489,N_16934,N_16833);
nand U17490 (N_17490,N_16815,N_17221);
nor U17491 (N_17491,N_17186,N_17101);
nor U17492 (N_17492,N_17142,N_16991);
nand U17493 (N_17493,N_17188,N_16879);
and U17494 (N_17494,N_16814,N_17166);
and U17495 (N_17495,N_17192,N_17086);
nor U17496 (N_17496,N_17330,N_16961);
or U17497 (N_17497,N_16937,N_17297);
nor U17498 (N_17498,N_17270,N_17071);
nand U17499 (N_17499,N_17193,N_16953);
nand U17500 (N_17500,N_17366,N_17227);
nor U17501 (N_17501,N_17187,N_16949);
and U17502 (N_17502,N_17021,N_17318);
or U17503 (N_17503,N_17097,N_17006);
or U17504 (N_17504,N_16936,N_16871);
or U17505 (N_17505,N_17067,N_17161);
or U17506 (N_17506,N_17174,N_17032);
or U17507 (N_17507,N_17052,N_17272);
nand U17508 (N_17508,N_17115,N_17035);
nor U17509 (N_17509,N_17120,N_16854);
nor U17510 (N_17510,N_17049,N_17202);
nand U17511 (N_17511,N_16983,N_16990);
or U17512 (N_17512,N_17156,N_16927);
nand U17513 (N_17513,N_16875,N_17323);
nand U17514 (N_17514,N_17057,N_17230);
or U17515 (N_17515,N_17310,N_16951);
and U17516 (N_17516,N_16906,N_17167);
nand U17517 (N_17517,N_17104,N_17178);
nor U17518 (N_17518,N_16818,N_16886);
and U17519 (N_17519,N_17243,N_17240);
or U17520 (N_17520,N_17143,N_16837);
and U17521 (N_17521,N_17044,N_17218);
nor U17522 (N_17522,N_17000,N_17208);
nor U17523 (N_17523,N_17121,N_17371);
nor U17524 (N_17524,N_16889,N_16970);
nor U17525 (N_17525,N_17315,N_17361);
nand U17526 (N_17526,N_16885,N_17065);
or U17527 (N_17527,N_17072,N_17068);
nor U17528 (N_17528,N_16957,N_16817);
and U17529 (N_17529,N_17268,N_17010);
or U17530 (N_17530,N_17380,N_16851);
nand U17531 (N_17531,N_17244,N_17285);
and U17532 (N_17532,N_17061,N_17201);
nor U17533 (N_17533,N_16959,N_16850);
nor U17534 (N_17534,N_17356,N_17106);
nand U17535 (N_17535,N_16908,N_17341);
nand U17536 (N_17536,N_17248,N_17189);
and U17537 (N_17537,N_16954,N_16964);
and U17538 (N_17538,N_16994,N_17128);
and U17539 (N_17539,N_16912,N_17100);
and U17540 (N_17540,N_16985,N_16805);
nor U17541 (N_17541,N_16956,N_17395);
or U17542 (N_17542,N_17346,N_17098);
nor U17543 (N_17543,N_16979,N_17388);
nand U17544 (N_17544,N_17396,N_17274);
and U17545 (N_17545,N_17251,N_16925);
or U17546 (N_17546,N_17351,N_16913);
or U17547 (N_17547,N_17136,N_17048);
nand U17548 (N_17548,N_17368,N_17031);
nand U17549 (N_17549,N_16911,N_17149);
and U17550 (N_17550,N_17304,N_17290);
and U17551 (N_17551,N_17027,N_16896);
nor U17552 (N_17552,N_17058,N_17054);
nand U17553 (N_17553,N_17175,N_16829);
nand U17554 (N_17554,N_17062,N_17163);
nand U17555 (N_17555,N_17332,N_16816);
and U17556 (N_17556,N_17316,N_16997);
nor U17557 (N_17557,N_16941,N_17129);
xor U17558 (N_17558,N_16819,N_17091);
nor U17559 (N_17559,N_16921,N_17169);
or U17560 (N_17560,N_17119,N_17255);
or U17561 (N_17561,N_16986,N_17039);
and U17562 (N_17562,N_17030,N_17377);
and U17563 (N_17563,N_17059,N_17096);
nand U17564 (N_17564,N_16843,N_17348);
nand U17565 (N_17565,N_17047,N_17237);
or U17566 (N_17566,N_17019,N_16988);
nand U17567 (N_17567,N_17041,N_17042);
nor U17568 (N_17568,N_16950,N_16844);
or U17569 (N_17569,N_17038,N_17384);
nor U17570 (N_17570,N_17253,N_16811);
nor U17571 (N_17571,N_17092,N_17074);
or U17572 (N_17572,N_17081,N_16962);
or U17573 (N_17573,N_17226,N_17307);
nand U17574 (N_17574,N_17337,N_17242);
or U17575 (N_17575,N_17087,N_17011);
or U17576 (N_17576,N_17385,N_17112);
or U17577 (N_17577,N_16822,N_17399);
or U17578 (N_17578,N_17206,N_17108);
nor U17579 (N_17579,N_17235,N_16869);
or U17580 (N_17580,N_17173,N_16806);
and U17581 (N_17581,N_17162,N_17372);
or U17582 (N_17582,N_17060,N_17376);
and U17583 (N_17583,N_16870,N_17247);
and U17584 (N_17584,N_16958,N_17144);
nor U17585 (N_17585,N_16928,N_17158);
nor U17586 (N_17586,N_17325,N_16845);
nor U17587 (N_17587,N_17004,N_17171);
and U17588 (N_17588,N_17350,N_16892);
nand U17589 (N_17589,N_17214,N_16865);
or U17590 (N_17590,N_16926,N_17258);
and U17591 (N_17591,N_17283,N_16924);
or U17592 (N_17592,N_16894,N_17090);
nand U17593 (N_17593,N_16918,N_17254);
and U17594 (N_17594,N_16955,N_17099);
or U17595 (N_17595,N_17138,N_17288);
nor U17596 (N_17596,N_17180,N_17111);
or U17597 (N_17597,N_17250,N_17217);
or U17598 (N_17598,N_17257,N_17275);
or U17599 (N_17599,N_16922,N_17252);
nor U17600 (N_17600,N_17299,N_17046);
nor U17601 (N_17601,N_17196,N_17154);
xnor U17602 (N_17602,N_16866,N_16842);
nand U17603 (N_17603,N_16861,N_17336);
xor U17604 (N_17604,N_17155,N_17246);
or U17605 (N_17605,N_17012,N_17093);
and U17606 (N_17606,N_16923,N_16975);
nand U17607 (N_17607,N_16899,N_17365);
nand U17608 (N_17608,N_17037,N_16992);
nor U17609 (N_17609,N_17229,N_17278);
nand U17610 (N_17610,N_16840,N_17050);
nand U17611 (N_17611,N_17133,N_16823);
or U17612 (N_17612,N_17259,N_17358);
or U17613 (N_17613,N_17014,N_17141);
nor U17614 (N_17614,N_16999,N_16858);
nand U17615 (N_17615,N_16824,N_17053);
and U17616 (N_17616,N_17109,N_16863);
or U17617 (N_17617,N_17172,N_16939);
and U17618 (N_17618,N_17291,N_17284);
nand U17619 (N_17619,N_17122,N_17340);
xnor U17620 (N_17620,N_17383,N_16862);
or U17621 (N_17621,N_17040,N_17359);
nor U17622 (N_17622,N_17177,N_16943);
and U17623 (N_17623,N_16909,N_17370);
and U17624 (N_17624,N_17139,N_17345);
nor U17625 (N_17625,N_17179,N_16810);
and U17626 (N_17626,N_17320,N_16993);
or U17627 (N_17627,N_16878,N_17280);
and U17628 (N_17628,N_16938,N_17212);
or U17629 (N_17629,N_17157,N_17228);
or U17630 (N_17630,N_16974,N_17207);
and U17631 (N_17631,N_16859,N_17084);
nand U17632 (N_17632,N_17002,N_17392);
nor U17633 (N_17633,N_17293,N_17344);
or U17634 (N_17634,N_16847,N_17369);
or U17635 (N_17635,N_17013,N_17198);
and U17636 (N_17636,N_17357,N_17381);
nand U17637 (N_17637,N_17269,N_17349);
and U17638 (N_17638,N_17363,N_16855);
nor U17639 (N_17639,N_17095,N_17302);
or U17640 (N_17640,N_17056,N_16830);
or U17641 (N_17641,N_16808,N_17296);
or U17642 (N_17642,N_17083,N_17379);
or U17643 (N_17643,N_16916,N_17352);
nor U17644 (N_17644,N_17025,N_17393);
nor U17645 (N_17645,N_16973,N_17024);
nand U17646 (N_17646,N_17215,N_16860);
or U17647 (N_17647,N_17137,N_16838);
nor U17648 (N_17648,N_17029,N_17311);
nand U17649 (N_17649,N_17262,N_16804);
and U17650 (N_17650,N_16980,N_16978);
nand U17651 (N_17651,N_17287,N_17233);
nor U17652 (N_17652,N_17339,N_16809);
nand U17653 (N_17653,N_17147,N_16929);
or U17654 (N_17654,N_16828,N_17182);
or U17655 (N_17655,N_16965,N_16888);
nand U17656 (N_17656,N_16826,N_17145);
nor U17657 (N_17657,N_17211,N_16910);
nor U17658 (N_17658,N_17319,N_16825);
or U17659 (N_17659,N_16835,N_17015);
and U17660 (N_17660,N_17170,N_17394);
or U17661 (N_17661,N_16917,N_16849);
nand U17662 (N_17662,N_17069,N_16932);
and U17663 (N_17663,N_17277,N_17181);
and U17664 (N_17664,N_17209,N_16904);
or U17665 (N_17665,N_17089,N_17135);
nand U17666 (N_17666,N_16995,N_17153);
nand U17667 (N_17667,N_17075,N_17281);
nor U17668 (N_17668,N_17308,N_17222);
nand U17669 (N_17669,N_16903,N_17118);
nand U17670 (N_17670,N_17386,N_17079);
nand U17671 (N_17671,N_17078,N_17105);
nand U17672 (N_17672,N_17213,N_17239);
and U17673 (N_17673,N_17327,N_17375);
nor U17674 (N_17674,N_17205,N_17343);
nor U17675 (N_17675,N_17347,N_16897);
or U17676 (N_17676,N_16969,N_17335);
nor U17677 (N_17677,N_16901,N_17051);
and U17678 (N_17678,N_17131,N_17043);
xnor U17679 (N_17679,N_16890,N_17328);
nor U17680 (N_17680,N_17342,N_16946);
nand U17681 (N_17681,N_16898,N_16984);
and U17682 (N_17682,N_17367,N_16800);
nor U17683 (N_17683,N_17374,N_16960);
nand U17684 (N_17684,N_16989,N_16832);
nor U17685 (N_17685,N_17063,N_17160);
or U17686 (N_17686,N_17076,N_17126);
or U17687 (N_17687,N_16801,N_16836);
nor U17688 (N_17688,N_16856,N_17249);
and U17689 (N_17689,N_16802,N_17168);
and U17690 (N_17690,N_17150,N_17331);
and U17691 (N_17691,N_17224,N_17003);
nor U17692 (N_17692,N_17017,N_17203);
nor U17693 (N_17693,N_17107,N_16947);
and U17694 (N_17694,N_17260,N_16966);
or U17695 (N_17695,N_16846,N_17334);
nor U17696 (N_17696,N_16919,N_17185);
nor U17697 (N_17697,N_17151,N_16807);
and U17698 (N_17698,N_17279,N_16876);
or U17699 (N_17699,N_17026,N_17309);
nor U17700 (N_17700,N_17037,N_17110);
nor U17701 (N_17701,N_17214,N_16880);
or U17702 (N_17702,N_17017,N_16954);
nand U17703 (N_17703,N_17225,N_17323);
nor U17704 (N_17704,N_17313,N_16902);
or U17705 (N_17705,N_17131,N_16920);
nor U17706 (N_17706,N_17116,N_17223);
or U17707 (N_17707,N_17009,N_16884);
or U17708 (N_17708,N_17232,N_16936);
nand U17709 (N_17709,N_17074,N_17126);
nand U17710 (N_17710,N_16920,N_17372);
nor U17711 (N_17711,N_16956,N_17116);
or U17712 (N_17712,N_17345,N_17093);
and U17713 (N_17713,N_17003,N_17238);
nand U17714 (N_17714,N_17067,N_17227);
xor U17715 (N_17715,N_17219,N_17205);
nand U17716 (N_17716,N_17158,N_16800);
nand U17717 (N_17717,N_17199,N_17244);
and U17718 (N_17718,N_16826,N_17291);
nor U17719 (N_17719,N_16956,N_17266);
or U17720 (N_17720,N_17312,N_17121);
nor U17721 (N_17721,N_17320,N_16859);
and U17722 (N_17722,N_17311,N_17288);
and U17723 (N_17723,N_17043,N_16921);
nor U17724 (N_17724,N_17368,N_16863);
nand U17725 (N_17725,N_17089,N_17186);
xor U17726 (N_17726,N_16844,N_17361);
nor U17727 (N_17727,N_17376,N_17220);
nor U17728 (N_17728,N_17007,N_17340);
or U17729 (N_17729,N_17123,N_17347);
xnor U17730 (N_17730,N_16916,N_17209);
or U17731 (N_17731,N_16941,N_16892);
and U17732 (N_17732,N_17149,N_17051);
xor U17733 (N_17733,N_17205,N_17223);
or U17734 (N_17734,N_16963,N_17332);
and U17735 (N_17735,N_17084,N_16992);
or U17736 (N_17736,N_17178,N_17079);
nor U17737 (N_17737,N_17341,N_17302);
nor U17738 (N_17738,N_17340,N_17394);
or U17739 (N_17739,N_16924,N_16810);
or U17740 (N_17740,N_17157,N_16866);
or U17741 (N_17741,N_17359,N_17348);
nor U17742 (N_17742,N_17157,N_16884);
or U17743 (N_17743,N_17091,N_17185);
nor U17744 (N_17744,N_17268,N_17138);
and U17745 (N_17745,N_17094,N_16891);
or U17746 (N_17746,N_17285,N_16869);
nand U17747 (N_17747,N_16920,N_17094);
or U17748 (N_17748,N_16851,N_17175);
nor U17749 (N_17749,N_17157,N_16937);
nand U17750 (N_17750,N_17295,N_17166);
nand U17751 (N_17751,N_16886,N_16873);
nand U17752 (N_17752,N_16948,N_17163);
nand U17753 (N_17753,N_17008,N_16936);
nor U17754 (N_17754,N_16832,N_16879);
or U17755 (N_17755,N_17172,N_17383);
or U17756 (N_17756,N_16918,N_16884);
nor U17757 (N_17757,N_17381,N_17189);
or U17758 (N_17758,N_17200,N_16942);
nand U17759 (N_17759,N_17348,N_17047);
nor U17760 (N_17760,N_17250,N_17125);
nand U17761 (N_17761,N_16853,N_17186);
nand U17762 (N_17762,N_17068,N_17158);
and U17763 (N_17763,N_17209,N_17145);
or U17764 (N_17764,N_16962,N_17226);
nand U17765 (N_17765,N_16936,N_17202);
and U17766 (N_17766,N_16841,N_17047);
nor U17767 (N_17767,N_17165,N_16823);
nor U17768 (N_17768,N_17091,N_16909);
nor U17769 (N_17769,N_16964,N_16988);
or U17770 (N_17770,N_17086,N_17060);
or U17771 (N_17771,N_17035,N_17311);
and U17772 (N_17772,N_17136,N_17119);
or U17773 (N_17773,N_17081,N_17114);
or U17774 (N_17774,N_17076,N_17002);
nand U17775 (N_17775,N_17254,N_17036);
nand U17776 (N_17776,N_17384,N_17330);
or U17777 (N_17777,N_16944,N_17373);
and U17778 (N_17778,N_16802,N_17281);
or U17779 (N_17779,N_17146,N_17022);
and U17780 (N_17780,N_17127,N_17013);
xor U17781 (N_17781,N_17276,N_17333);
or U17782 (N_17782,N_17347,N_16899);
or U17783 (N_17783,N_17195,N_17276);
and U17784 (N_17784,N_17366,N_17201);
and U17785 (N_17785,N_16915,N_16885);
or U17786 (N_17786,N_17302,N_17327);
and U17787 (N_17787,N_17040,N_17282);
nand U17788 (N_17788,N_16989,N_17056);
and U17789 (N_17789,N_16977,N_16986);
nor U17790 (N_17790,N_17001,N_17212);
nand U17791 (N_17791,N_17337,N_17041);
nand U17792 (N_17792,N_16832,N_16994);
nor U17793 (N_17793,N_17290,N_17248);
nor U17794 (N_17794,N_17170,N_17100);
nand U17795 (N_17795,N_17099,N_16894);
nor U17796 (N_17796,N_17061,N_16856);
or U17797 (N_17797,N_17161,N_17379);
or U17798 (N_17798,N_16937,N_16846);
and U17799 (N_17799,N_16985,N_17388);
nor U17800 (N_17800,N_16886,N_17296);
nor U17801 (N_17801,N_17189,N_17026);
or U17802 (N_17802,N_17205,N_17118);
and U17803 (N_17803,N_17298,N_17358);
xnor U17804 (N_17804,N_17249,N_17198);
and U17805 (N_17805,N_17179,N_17116);
nor U17806 (N_17806,N_17072,N_17391);
and U17807 (N_17807,N_16834,N_17239);
nand U17808 (N_17808,N_17061,N_16994);
nor U17809 (N_17809,N_16840,N_17221);
nand U17810 (N_17810,N_16876,N_17120);
nand U17811 (N_17811,N_17056,N_17235);
or U17812 (N_17812,N_16868,N_16887);
and U17813 (N_17813,N_17025,N_16835);
and U17814 (N_17814,N_16959,N_17298);
nor U17815 (N_17815,N_17005,N_17328);
and U17816 (N_17816,N_17284,N_17316);
nor U17817 (N_17817,N_17256,N_17146);
nor U17818 (N_17818,N_17358,N_17021);
nor U17819 (N_17819,N_17074,N_17163);
and U17820 (N_17820,N_16809,N_16823);
or U17821 (N_17821,N_16852,N_16819);
xor U17822 (N_17822,N_16966,N_17187);
nor U17823 (N_17823,N_16890,N_17376);
or U17824 (N_17824,N_17373,N_16911);
nand U17825 (N_17825,N_17038,N_17211);
and U17826 (N_17826,N_17187,N_17193);
and U17827 (N_17827,N_17350,N_16813);
nor U17828 (N_17828,N_17084,N_17139);
and U17829 (N_17829,N_17055,N_17112);
nor U17830 (N_17830,N_16904,N_17093);
nor U17831 (N_17831,N_17047,N_16813);
nand U17832 (N_17832,N_17056,N_17348);
or U17833 (N_17833,N_17232,N_17162);
nor U17834 (N_17834,N_17370,N_16926);
xnor U17835 (N_17835,N_17260,N_17195);
xnor U17836 (N_17836,N_16949,N_17365);
nand U17837 (N_17837,N_17381,N_17187);
nor U17838 (N_17838,N_16804,N_17366);
nor U17839 (N_17839,N_17214,N_16964);
and U17840 (N_17840,N_17084,N_16893);
or U17841 (N_17841,N_17357,N_16987);
nor U17842 (N_17842,N_17322,N_16994);
or U17843 (N_17843,N_17059,N_16881);
nor U17844 (N_17844,N_17390,N_16888);
nor U17845 (N_17845,N_16846,N_16845);
nand U17846 (N_17846,N_17384,N_17197);
xnor U17847 (N_17847,N_16937,N_17373);
nor U17848 (N_17848,N_17238,N_17375);
nor U17849 (N_17849,N_17114,N_16890);
nand U17850 (N_17850,N_16868,N_17110);
nand U17851 (N_17851,N_16980,N_17209);
nor U17852 (N_17852,N_16943,N_17003);
or U17853 (N_17853,N_17087,N_17244);
and U17854 (N_17854,N_16833,N_16841);
xnor U17855 (N_17855,N_17248,N_17391);
or U17856 (N_17856,N_17127,N_17145);
nand U17857 (N_17857,N_16880,N_17187);
nor U17858 (N_17858,N_16892,N_17166);
nor U17859 (N_17859,N_16888,N_17382);
nor U17860 (N_17860,N_17180,N_17155);
nand U17861 (N_17861,N_17369,N_17179);
or U17862 (N_17862,N_17036,N_17020);
and U17863 (N_17863,N_17366,N_16848);
nand U17864 (N_17864,N_16889,N_17214);
nand U17865 (N_17865,N_16883,N_16930);
and U17866 (N_17866,N_17285,N_17166);
or U17867 (N_17867,N_16957,N_16992);
nand U17868 (N_17868,N_16962,N_17236);
and U17869 (N_17869,N_17015,N_17397);
or U17870 (N_17870,N_17136,N_17375);
nand U17871 (N_17871,N_17125,N_17259);
nor U17872 (N_17872,N_16895,N_17223);
nor U17873 (N_17873,N_16964,N_17076);
or U17874 (N_17874,N_17393,N_17254);
nand U17875 (N_17875,N_17014,N_16809);
nor U17876 (N_17876,N_16927,N_16965);
nor U17877 (N_17877,N_17015,N_17010);
and U17878 (N_17878,N_16819,N_16848);
and U17879 (N_17879,N_17399,N_17310);
nand U17880 (N_17880,N_17113,N_17254);
nand U17881 (N_17881,N_17035,N_17085);
nor U17882 (N_17882,N_16998,N_17360);
nor U17883 (N_17883,N_17053,N_16979);
nor U17884 (N_17884,N_16845,N_17346);
or U17885 (N_17885,N_17347,N_17186);
nand U17886 (N_17886,N_16882,N_16887);
nand U17887 (N_17887,N_16872,N_16892);
and U17888 (N_17888,N_17056,N_17076);
nand U17889 (N_17889,N_16840,N_16874);
and U17890 (N_17890,N_17137,N_17023);
nor U17891 (N_17891,N_16934,N_17237);
and U17892 (N_17892,N_16909,N_17313);
nor U17893 (N_17893,N_17147,N_17235);
nand U17894 (N_17894,N_17095,N_17290);
or U17895 (N_17895,N_17248,N_17124);
or U17896 (N_17896,N_16871,N_17063);
and U17897 (N_17897,N_17135,N_16854);
or U17898 (N_17898,N_17090,N_17084);
and U17899 (N_17899,N_16823,N_17259);
or U17900 (N_17900,N_17333,N_17054);
xor U17901 (N_17901,N_16903,N_16874);
nand U17902 (N_17902,N_16901,N_17165);
xor U17903 (N_17903,N_16999,N_16887);
nand U17904 (N_17904,N_16991,N_16889);
nand U17905 (N_17905,N_17307,N_17064);
nand U17906 (N_17906,N_17070,N_17030);
nor U17907 (N_17907,N_17103,N_17338);
or U17908 (N_17908,N_17038,N_17176);
and U17909 (N_17909,N_16894,N_16842);
or U17910 (N_17910,N_16990,N_17078);
xnor U17911 (N_17911,N_17020,N_16891);
or U17912 (N_17912,N_17040,N_16856);
nand U17913 (N_17913,N_16868,N_16863);
nor U17914 (N_17914,N_16980,N_17365);
nor U17915 (N_17915,N_17014,N_17111);
nor U17916 (N_17916,N_17033,N_16899);
nand U17917 (N_17917,N_17182,N_16959);
and U17918 (N_17918,N_17174,N_16916);
nand U17919 (N_17919,N_16801,N_17396);
nand U17920 (N_17920,N_16887,N_17006);
or U17921 (N_17921,N_17208,N_17388);
or U17922 (N_17922,N_16931,N_16980);
and U17923 (N_17923,N_16996,N_17379);
nor U17924 (N_17924,N_17058,N_16881);
and U17925 (N_17925,N_17214,N_17013);
and U17926 (N_17926,N_17153,N_17015);
and U17927 (N_17927,N_16869,N_17155);
nor U17928 (N_17928,N_17130,N_17049);
or U17929 (N_17929,N_16899,N_17231);
nor U17930 (N_17930,N_17282,N_17225);
nor U17931 (N_17931,N_17170,N_17330);
or U17932 (N_17932,N_17313,N_16841);
nor U17933 (N_17933,N_17201,N_17047);
or U17934 (N_17934,N_17345,N_16981);
or U17935 (N_17935,N_16998,N_16973);
nand U17936 (N_17936,N_17057,N_16845);
or U17937 (N_17937,N_17278,N_17031);
nand U17938 (N_17938,N_17216,N_17074);
nor U17939 (N_17939,N_17355,N_17104);
nor U17940 (N_17940,N_17275,N_16989);
nor U17941 (N_17941,N_16881,N_17044);
nand U17942 (N_17942,N_16954,N_16872);
and U17943 (N_17943,N_17207,N_17158);
or U17944 (N_17944,N_17281,N_16889);
nand U17945 (N_17945,N_16914,N_17051);
nand U17946 (N_17946,N_17246,N_17017);
or U17947 (N_17947,N_17244,N_16848);
or U17948 (N_17948,N_17306,N_17026);
and U17949 (N_17949,N_17095,N_17296);
or U17950 (N_17950,N_17178,N_16824);
nor U17951 (N_17951,N_17242,N_16892);
nand U17952 (N_17952,N_16821,N_17106);
nor U17953 (N_17953,N_16917,N_17199);
nand U17954 (N_17954,N_17277,N_17001);
nor U17955 (N_17955,N_17062,N_16876);
and U17956 (N_17956,N_16864,N_16918);
nand U17957 (N_17957,N_17277,N_16906);
nor U17958 (N_17958,N_17302,N_17224);
nor U17959 (N_17959,N_16848,N_17248);
or U17960 (N_17960,N_16911,N_16878);
nor U17961 (N_17961,N_17140,N_17312);
xor U17962 (N_17962,N_17100,N_17232);
nand U17963 (N_17963,N_17045,N_17373);
nor U17964 (N_17964,N_17252,N_17103);
and U17965 (N_17965,N_17288,N_16895);
and U17966 (N_17966,N_17047,N_16876);
or U17967 (N_17967,N_17130,N_17092);
or U17968 (N_17968,N_17248,N_17395);
nor U17969 (N_17969,N_17098,N_17320);
xor U17970 (N_17970,N_16938,N_17150);
nor U17971 (N_17971,N_17074,N_17113);
xnor U17972 (N_17972,N_17029,N_17272);
and U17973 (N_17973,N_17134,N_17341);
nor U17974 (N_17974,N_17313,N_17134);
nor U17975 (N_17975,N_17023,N_16984);
nand U17976 (N_17976,N_16885,N_17173);
nand U17977 (N_17977,N_17072,N_16896);
or U17978 (N_17978,N_17201,N_17093);
nor U17979 (N_17979,N_17099,N_17397);
and U17980 (N_17980,N_17018,N_17281);
nand U17981 (N_17981,N_17303,N_16922);
and U17982 (N_17982,N_17311,N_17204);
or U17983 (N_17983,N_17131,N_16864);
nand U17984 (N_17984,N_17300,N_16984);
nor U17985 (N_17985,N_17038,N_17154);
or U17986 (N_17986,N_17251,N_16929);
nor U17987 (N_17987,N_16984,N_16928);
nand U17988 (N_17988,N_17318,N_17019);
nor U17989 (N_17989,N_16927,N_17031);
or U17990 (N_17990,N_17374,N_17338);
and U17991 (N_17991,N_17103,N_16856);
and U17992 (N_17992,N_17197,N_17375);
or U17993 (N_17993,N_17302,N_17311);
and U17994 (N_17994,N_17297,N_16837);
or U17995 (N_17995,N_17020,N_16832);
nand U17996 (N_17996,N_16878,N_17049);
nand U17997 (N_17997,N_16872,N_16923);
nand U17998 (N_17998,N_17149,N_17343);
nor U17999 (N_17999,N_16985,N_16974);
or U18000 (N_18000,N_17854,N_17827);
nand U18001 (N_18001,N_17817,N_17555);
or U18002 (N_18002,N_17882,N_17762);
and U18003 (N_18003,N_17510,N_17716);
nor U18004 (N_18004,N_17464,N_17443);
nor U18005 (N_18005,N_17576,N_17933);
or U18006 (N_18006,N_17564,N_17631);
nor U18007 (N_18007,N_17805,N_17522);
or U18008 (N_18008,N_17757,N_17847);
and U18009 (N_18009,N_17936,N_17872);
and U18010 (N_18010,N_17893,N_17704);
or U18011 (N_18011,N_17569,N_17519);
or U18012 (N_18012,N_17639,N_17620);
or U18013 (N_18013,N_17518,N_17635);
and U18014 (N_18014,N_17850,N_17766);
nor U18015 (N_18015,N_17923,N_17410);
or U18016 (N_18016,N_17862,N_17965);
or U18017 (N_18017,N_17498,N_17483);
nand U18018 (N_18018,N_17504,N_17680);
nor U18019 (N_18019,N_17954,N_17619);
and U18020 (N_18020,N_17688,N_17864);
nor U18021 (N_18021,N_17903,N_17673);
or U18022 (N_18022,N_17646,N_17616);
and U18023 (N_18023,N_17986,N_17694);
or U18024 (N_18024,N_17445,N_17552);
nand U18025 (N_18025,N_17718,N_17804);
nor U18026 (N_18026,N_17562,N_17963);
or U18027 (N_18027,N_17982,N_17431);
and U18028 (N_18028,N_17558,N_17831);
or U18029 (N_18029,N_17597,N_17481);
nand U18030 (N_18030,N_17434,N_17934);
and U18031 (N_18031,N_17846,N_17784);
nor U18032 (N_18032,N_17949,N_17835);
and U18033 (N_18033,N_17623,N_17977);
or U18034 (N_18034,N_17890,N_17681);
nand U18035 (N_18035,N_17806,N_17426);
nor U18036 (N_18036,N_17580,N_17606);
and U18037 (N_18037,N_17826,N_17417);
and U18038 (N_18038,N_17726,N_17617);
or U18039 (N_18039,N_17554,N_17799);
or U18040 (N_18040,N_17689,N_17414);
nand U18041 (N_18041,N_17700,N_17750);
nand U18042 (N_18042,N_17975,N_17989);
and U18043 (N_18043,N_17733,N_17676);
xor U18044 (N_18044,N_17520,N_17674);
or U18045 (N_18045,N_17690,N_17729);
and U18046 (N_18046,N_17730,N_17735);
or U18047 (N_18047,N_17720,N_17664);
or U18048 (N_18048,N_17636,N_17840);
or U18049 (N_18049,N_17715,N_17752);
nor U18050 (N_18050,N_17601,N_17480);
or U18051 (N_18051,N_17560,N_17915);
nand U18052 (N_18052,N_17845,N_17849);
nand U18053 (N_18053,N_17906,N_17657);
nand U18054 (N_18054,N_17599,N_17789);
nor U18055 (N_18055,N_17472,N_17615);
nand U18056 (N_18056,N_17914,N_17887);
nor U18057 (N_18057,N_17839,N_17880);
nor U18058 (N_18058,N_17910,N_17433);
nor U18059 (N_18059,N_17878,N_17452);
and U18060 (N_18060,N_17979,N_17763);
or U18061 (N_18061,N_17419,N_17496);
nand U18062 (N_18062,N_17721,N_17425);
nor U18063 (N_18063,N_17473,N_17595);
nor U18064 (N_18064,N_17465,N_17753);
and U18065 (N_18065,N_17941,N_17810);
and U18066 (N_18066,N_17413,N_17886);
nor U18067 (N_18067,N_17405,N_17874);
or U18068 (N_18068,N_17660,N_17503);
nor U18069 (N_18069,N_17786,N_17513);
nand U18070 (N_18070,N_17628,N_17900);
and U18071 (N_18071,N_17950,N_17953);
or U18072 (N_18072,N_17633,N_17454);
nor U18073 (N_18073,N_17883,N_17524);
and U18074 (N_18074,N_17561,N_17427);
and U18075 (N_18075,N_17695,N_17816);
nor U18076 (N_18076,N_17798,N_17820);
or U18077 (N_18077,N_17958,N_17921);
xor U18078 (N_18078,N_17647,N_17858);
or U18079 (N_18079,N_17962,N_17719);
nand U18080 (N_18080,N_17844,N_17671);
and U18081 (N_18081,N_17570,N_17612);
and U18082 (N_18082,N_17998,N_17706);
nand U18083 (N_18083,N_17439,N_17546);
and U18084 (N_18084,N_17904,N_17774);
nand U18085 (N_18085,N_17404,N_17794);
or U18086 (N_18086,N_17604,N_17709);
nor U18087 (N_18087,N_17743,N_17731);
or U18088 (N_18088,N_17575,N_17655);
nor U18089 (N_18089,N_17551,N_17931);
nand U18090 (N_18090,N_17705,N_17521);
and U18091 (N_18091,N_17768,N_17912);
or U18092 (N_18092,N_17767,N_17744);
and U18093 (N_18093,N_17765,N_17782);
and U18094 (N_18094,N_17453,N_17486);
nand U18095 (N_18095,N_17583,N_17833);
nor U18096 (N_18096,N_17420,N_17780);
nor U18097 (N_18097,N_17402,N_17468);
and U18098 (N_18098,N_17867,N_17838);
nor U18099 (N_18099,N_17710,N_17937);
and U18100 (N_18100,N_17544,N_17972);
or U18101 (N_18101,N_17778,N_17692);
or U18102 (N_18102,N_17699,N_17578);
and U18103 (N_18103,N_17907,N_17935);
and U18104 (N_18104,N_17819,N_17701);
nand U18105 (N_18105,N_17632,N_17802);
nand U18106 (N_18106,N_17484,N_17531);
nor U18107 (N_18107,N_17600,N_17999);
and U18108 (N_18108,N_17523,N_17591);
or U18109 (N_18109,N_17856,N_17916);
nand U18110 (N_18110,N_17788,N_17447);
nand U18111 (N_18111,N_17538,N_17500);
and U18112 (N_18112,N_17714,N_17793);
or U18113 (N_18113,N_17543,N_17581);
and U18114 (N_18114,N_17622,N_17913);
or U18115 (N_18115,N_17529,N_17897);
nor U18116 (N_18116,N_17942,N_17997);
nand U18117 (N_18117,N_17456,N_17458);
and U18118 (N_18118,N_17667,N_17888);
nand U18119 (N_18119,N_17516,N_17596);
and U18120 (N_18120,N_17951,N_17961);
nand U18121 (N_18121,N_17938,N_17821);
nand U18122 (N_18122,N_17514,N_17926);
or U18123 (N_18123,N_17625,N_17918);
nor U18124 (N_18124,N_17848,N_17577);
xor U18125 (N_18125,N_17853,N_17917);
or U18126 (N_18126,N_17421,N_17542);
or U18127 (N_18127,N_17870,N_17640);
nor U18128 (N_18128,N_17801,N_17852);
nor U18129 (N_18129,N_17851,N_17995);
nand U18130 (N_18130,N_17505,N_17672);
nand U18131 (N_18131,N_17517,N_17829);
and U18132 (N_18132,N_17613,N_17602);
nand U18133 (N_18133,N_17808,N_17892);
nor U18134 (N_18134,N_17584,N_17637);
nor U18135 (N_18135,N_17841,N_17857);
or U18136 (N_18136,N_17448,N_17630);
or U18137 (N_18137,N_17968,N_17740);
or U18138 (N_18138,N_17828,N_17470);
and U18139 (N_18139,N_17509,N_17830);
nand U18140 (N_18140,N_17945,N_17708);
nand U18141 (N_18141,N_17755,N_17476);
nand U18142 (N_18142,N_17573,N_17587);
and U18143 (N_18143,N_17738,N_17537);
nand U18144 (N_18144,N_17873,N_17653);
nor U18145 (N_18145,N_17444,N_17588);
and U18146 (N_18146,N_17506,N_17812);
or U18147 (N_18147,N_17651,N_17732);
nor U18148 (N_18148,N_17556,N_17693);
nand U18149 (N_18149,N_17928,N_17787);
nand U18150 (N_18150,N_17605,N_17607);
and U18151 (N_18151,N_17990,N_17462);
and U18152 (N_18152,N_17559,N_17776);
nor U18153 (N_18153,N_17495,N_17956);
or U18154 (N_18154,N_17791,N_17512);
nand U18155 (N_18155,N_17884,N_17834);
xor U18156 (N_18156,N_17469,N_17525);
or U18157 (N_18157,N_17869,N_17980);
xnor U18158 (N_18158,N_17401,N_17547);
and U18159 (N_18159,N_17482,N_17624);
or U18160 (N_18160,N_17978,N_17803);
or U18161 (N_18161,N_17837,N_17698);
and U18162 (N_18162,N_17984,N_17885);
and U18163 (N_18163,N_17568,N_17492);
nor U18164 (N_18164,N_17611,N_17594);
and U18165 (N_18165,N_17534,N_17407);
nor U18166 (N_18166,N_17415,N_17683);
nor U18167 (N_18167,N_17641,N_17758);
nand U18168 (N_18168,N_17796,N_17756);
nand U18169 (N_18169,N_17955,N_17603);
and U18170 (N_18170,N_17761,N_17855);
or U18171 (N_18171,N_17939,N_17675);
nor U18172 (N_18172,N_17638,N_17440);
nor U18173 (N_18173,N_17571,N_17739);
and U18174 (N_18174,N_17457,N_17707);
or U18175 (N_18175,N_17927,N_17842);
nor U18176 (N_18176,N_17993,N_17662);
or U18177 (N_18177,N_17973,N_17467);
or U18178 (N_18178,N_17889,N_17745);
and U18179 (N_18179,N_17811,N_17661);
and U18180 (N_18180,N_17749,N_17746);
or U18181 (N_18181,N_17553,N_17988);
nor U18182 (N_18182,N_17932,N_17679);
xor U18183 (N_18183,N_17654,N_17530);
and U18184 (N_18184,N_17741,N_17742);
and U18185 (N_18185,N_17723,N_17435);
and U18186 (N_18186,N_17860,N_17686);
and U18187 (N_18187,N_17795,N_17574);
or U18188 (N_18188,N_17712,N_17943);
nand U18189 (N_18189,N_17894,N_17441);
and U18190 (N_18190,N_17899,N_17919);
or U18191 (N_18191,N_17754,N_17960);
nor U18192 (N_18192,N_17987,N_17772);
nand U18193 (N_18193,N_17650,N_17843);
or U18194 (N_18194,N_17976,N_17540);
nand U18195 (N_18195,N_17461,N_17877);
or U18196 (N_18196,N_17901,N_17929);
xnor U18197 (N_18197,N_17409,N_17466);
or U18198 (N_18198,N_17471,N_17866);
nand U18199 (N_18199,N_17515,N_17450);
nor U18200 (N_18200,N_17511,N_17737);
nand U18201 (N_18201,N_17947,N_17930);
nor U18202 (N_18202,N_17609,N_17593);
xnor U18203 (N_18203,N_17626,N_17643);
or U18204 (N_18204,N_17598,N_17487);
nor U18205 (N_18205,N_17891,N_17996);
nor U18206 (N_18206,N_17896,N_17687);
nor U18207 (N_18207,N_17861,N_17663);
nor U18208 (N_18208,N_17474,N_17533);
nor U18209 (N_18209,N_17983,N_17711);
or U18210 (N_18210,N_17898,N_17644);
and U18211 (N_18211,N_17779,N_17528);
nand U18212 (N_18212,N_17957,N_17446);
or U18213 (N_18213,N_17436,N_17814);
or U18214 (N_18214,N_17771,N_17432);
or U18215 (N_18215,N_17684,N_17502);
nand U18216 (N_18216,N_17437,N_17621);
and U18217 (N_18217,N_17769,N_17557);
nand U18218 (N_18218,N_17460,N_17909);
nor U18219 (N_18219,N_17497,N_17734);
nor U18220 (N_18220,N_17614,N_17634);
nor U18221 (N_18221,N_17964,N_17567);
nand U18222 (N_18222,N_17871,N_17902);
or U18223 (N_18223,N_17728,N_17759);
nor U18224 (N_18224,N_17985,N_17566);
nand U18225 (N_18225,N_17809,N_17682);
or U18226 (N_18226,N_17781,N_17920);
nor U18227 (N_18227,N_17549,N_17944);
and U18228 (N_18228,N_17823,N_17775);
and U18229 (N_18229,N_17717,N_17665);
nand U18230 (N_18230,N_17959,N_17565);
and U18231 (N_18231,N_17760,N_17792);
nand U18232 (N_18232,N_17590,N_17535);
nand U18233 (N_18233,N_17971,N_17800);
or U18234 (N_18234,N_17668,N_17627);
xnor U18235 (N_18235,N_17491,N_17526);
or U18236 (N_18236,N_17952,N_17488);
nand U18237 (N_18237,N_17429,N_17659);
nor U18238 (N_18238,N_17875,N_17748);
nand U18239 (N_18239,N_17449,N_17418);
nor U18240 (N_18240,N_17783,N_17969);
nand U18241 (N_18241,N_17966,N_17656);
or U18242 (N_18242,N_17702,N_17642);
nand U18243 (N_18243,N_17863,N_17697);
and U18244 (N_18244,N_17489,N_17548);
and U18245 (N_18245,N_17770,N_17691);
and U18246 (N_18246,N_17992,N_17807);
nor U18247 (N_18247,N_17677,N_17494);
or U18248 (N_18248,N_17493,N_17545);
nor U18249 (N_18249,N_17678,N_17824);
or U18250 (N_18250,N_17940,N_17868);
or U18251 (N_18251,N_17648,N_17724);
or U18252 (N_18252,N_17881,N_17400);
or U18253 (N_18253,N_17991,N_17406);
or U18254 (N_18254,N_17785,N_17879);
and U18255 (N_18255,N_17508,N_17696);
or U18256 (N_18256,N_17713,N_17685);
and U18257 (N_18257,N_17618,N_17475);
or U18258 (N_18258,N_17725,N_17666);
and U18259 (N_18259,N_17922,N_17925);
nand U18260 (N_18260,N_17527,N_17859);
and U18261 (N_18261,N_17790,N_17490);
or U18262 (N_18262,N_17946,N_17585);
and U18263 (N_18263,N_17722,N_17563);
and U18264 (N_18264,N_17411,N_17451);
nor U18265 (N_18265,N_17536,N_17815);
or U18266 (N_18266,N_17478,N_17797);
nand U18267 (N_18267,N_17610,N_17550);
nand U18268 (N_18268,N_17412,N_17736);
nor U18269 (N_18269,N_17658,N_17582);
xor U18270 (N_18270,N_17455,N_17994);
nand U18271 (N_18271,N_17645,N_17438);
nor U18272 (N_18272,N_17572,N_17485);
nor U18273 (N_18273,N_17608,N_17477);
nand U18274 (N_18274,N_17422,N_17579);
and U18275 (N_18275,N_17905,N_17813);
nand U18276 (N_18276,N_17592,N_17541);
or U18277 (N_18277,N_17430,N_17408);
nor U18278 (N_18278,N_17764,N_17442);
nand U18279 (N_18279,N_17825,N_17747);
nor U18280 (N_18280,N_17818,N_17539);
nor U18281 (N_18281,N_17501,N_17970);
or U18282 (N_18282,N_17924,N_17586);
nor U18283 (N_18283,N_17865,N_17832);
nor U18284 (N_18284,N_17499,N_17703);
or U18285 (N_18285,N_17967,N_17911);
and U18286 (N_18286,N_17652,N_17777);
or U18287 (N_18287,N_17751,N_17416);
nand U18288 (N_18288,N_17428,N_17876);
nor U18289 (N_18289,N_17424,N_17507);
nor U18290 (N_18290,N_17629,N_17403);
nand U18291 (N_18291,N_17773,N_17948);
or U18292 (N_18292,N_17727,N_17532);
and U18293 (N_18293,N_17974,N_17836);
and U18294 (N_18294,N_17423,N_17981);
xor U18295 (N_18295,N_17459,N_17463);
and U18296 (N_18296,N_17479,N_17822);
nor U18297 (N_18297,N_17895,N_17670);
nor U18298 (N_18298,N_17908,N_17589);
or U18299 (N_18299,N_17669,N_17649);
or U18300 (N_18300,N_17494,N_17724);
or U18301 (N_18301,N_17772,N_17515);
nor U18302 (N_18302,N_17868,N_17986);
and U18303 (N_18303,N_17962,N_17646);
nand U18304 (N_18304,N_17646,N_17813);
nor U18305 (N_18305,N_17915,N_17755);
or U18306 (N_18306,N_17552,N_17527);
nor U18307 (N_18307,N_17535,N_17851);
or U18308 (N_18308,N_17685,N_17615);
nor U18309 (N_18309,N_17559,N_17916);
or U18310 (N_18310,N_17516,N_17986);
nand U18311 (N_18311,N_17885,N_17441);
nand U18312 (N_18312,N_17925,N_17438);
nor U18313 (N_18313,N_17835,N_17549);
and U18314 (N_18314,N_17661,N_17796);
nor U18315 (N_18315,N_17509,N_17809);
or U18316 (N_18316,N_17843,N_17498);
nand U18317 (N_18317,N_17974,N_17941);
or U18318 (N_18318,N_17608,N_17633);
xor U18319 (N_18319,N_17588,N_17849);
nor U18320 (N_18320,N_17712,N_17562);
nand U18321 (N_18321,N_17645,N_17671);
nor U18322 (N_18322,N_17808,N_17611);
nand U18323 (N_18323,N_17608,N_17406);
and U18324 (N_18324,N_17697,N_17955);
and U18325 (N_18325,N_17971,N_17583);
and U18326 (N_18326,N_17759,N_17705);
and U18327 (N_18327,N_17952,N_17550);
and U18328 (N_18328,N_17589,N_17523);
nor U18329 (N_18329,N_17466,N_17902);
and U18330 (N_18330,N_17769,N_17961);
or U18331 (N_18331,N_17743,N_17733);
nand U18332 (N_18332,N_17681,N_17706);
or U18333 (N_18333,N_17539,N_17792);
or U18334 (N_18334,N_17811,N_17791);
and U18335 (N_18335,N_17872,N_17454);
nor U18336 (N_18336,N_17759,N_17723);
and U18337 (N_18337,N_17729,N_17989);
nor U18338 (N_18338,N_17487,N_17677);
nor U18339 (N_18339,N_17626,N_17546);
nor U18340 (N_18340,N_17589,N_17834);
and U18341 (N_18341,N_17666,N_17750);
nor U18342 (N_18342,N_17467,N_17524);
nand U18343 (N_18343,N_17532,N_17747);
nor U18344 (N_18344,N_17553,N_17505);
nand U18345 (N_18345,N_17995,N_17472);
nor U18346 (N_18346,N_17725,N_17664);
nor U18347 (N_18347,N_17509,N_17541);
and U18348 (N_18348,N_17463,N_17643);
and U18349 (N_18349,N_17590,N_17938);
nor U18350 (N_18350,N_17692,N_17938);
xor U18351 (N_18351,N_17659,N_17675);
or U18352 (N_18352,N_17492,N_17473);
nand U18353 (N_18353,N_17748,N_17918);
and U18354 (N_18354,N_17741,N_17944);
nor U18355 (N_18355,N_17770,N_17680);
nand U18356 (N_18356,N_17749,N_17617);
or U18357 (N_18357,N_17519,N_17779);
and U18358 (N_18358,N_17451,N_17497);
and U18359 (N_18359,N_17606,N_17827);
or U18360 (N_18360,N_17542,N_17600);
nor U18361 (N_18361,N_17850,N_17999);
or U18362 (N_18362,N_17770,N_17571);
and U18363 (N_18363,N_17816,N_17800);
or U18364 (N_18364,N_17801,N_17437);
or U18365 (N_18365,N_17434,N_17871);
or U18366 (N_18366,N_17445,N_17871);
nand U18367 (N_18367,N_17649,N_17926);
nor U18368 (N_18368,N_17730,N_17782);
and U18369 (N_18369,N_17424,N_17449);
or U18370 (N_18370,N_17956,N_17467);
nor U18371 (N_18371,N_17551,N_17847);
or U18372 (N_18372,N_17766,N_17839);
nand U18373 (N_18373,N_17773,N_17593);
and U18374 (N_18374,N_17681,N_17914);
nand U18375 (N_18375,N_17826,N_17567);
and U18376 (N_18376,N_17440,N_17411);
nand U18377 (N_18377,N_17982,N_17656);
and U18378 (N_18378,N_17946,N_17552);
or U18379 (N_18379,N_17613,N_17833);
or U18380 (N_18380,N_17577,N_17828);
nor U18381 (N_18381,N_17675,N_17624);
and U18382 (N_18382,N_17518,N_17705);
nand U18383 (N_18383,N_17608,N_17987);
nand U18384 (N_18384,N_17871,N_17413);
or U18385 (N_18385,N_17827,N_17665);
or U18386 (N_18386,N_17836,N_17522);
nor U18387 (N_18387,N_17444,N_17416);
nand U18388 (N_18388,N_17423,N_17792);
and U18389 (N_18389,N_17465,N_17760);
nor U18390 (N_18390,N_17464,N_17782);
or U18391 (N_18391,N_17933,N_17863);
nor U18392 (N_18392,N_17662,N_17623);
and U18393 (N_18393,N_17730,N_17513);
nor U18394 (N_18394,N_17897,N_17848);
and U18395 (N_18395,N_17751,N_17418);
nor U18396 (N_18396,N_17675,N_17471);
nand U18397 (N_18397,N_17644,N_17848);
and U18398 (N_18398,N_17526,N_17884);
nor U18399 (N_18399,N_17828,N_17474);
nor U18400 (N_18400,N_17775,N_17452);
nor U18401 (N_18401,N_17942,N_17474);
nand U18402 (N_18402,N_17988,N_17722);
nor U18403 (N_18403,N_17486,N_17483);
nand U18404 (N_18404,N_17929,N_17939);
nand U18405 (N_18405,N_17900,N_17922);
and U18406 (N_18406,N_17661,N_17847);
and U18407 (N_18407,N_17964,N_17773);
nand U18408 (N_18408,N_17606,N_17795);
nor U18409 (N_18409,N_17688,N_17423);
and U18410 (N_18410,N_17933,N_17902);
nand U18411 (N_18411,N_17657,N_17537);
or U18412 (N_18412,N_17959,N_17902);
nand U18413 (N_18413,N_17918,N_17628);
nand U18414 (N_18414,N_17825,N_17938);
nor U18415 (N_18415,N_17968,N_17433);
nor U18416 (N_18416,N_17448,N_17540);
and U18417 (N_18417,N_17522,N_17949);
and U18418 (N_18418,N_17831,N_17727);
or U18419 (N_18419,N_17750,N_17680);
nor U18420 (N_18420,N_17517,N_17999);
and U18421 (N_18421,N_17757,N_17932);
nand U18422 (N_18422,N_17680,N_17854);
and U18423 (N_18423,N_17534,N_17701);
xnor U18424 (N_18424,N_17419,N_17756);
nand U18425 (N_18425,N_17778,N_17511);
nand U18426 (N_18426,N_17748,N_17715);
or U18427 (N_18427,N_17510,N_17843);
nand U18428 (N_18428,N_17417,N_17433);
and U18429 (N_18429,N_17788,N_17980);
or U18430 (N_18430,N_17460,N_17988);
nand U18431 (N_18431,N_17661,N_17894);
or U18432 (N_18432,N_17706,N_17518);
nand U18433 (N_18433,N_17709,N_17814);
nor U18434 (N_18434,N_17456,N_17637);
and U18435 (N_18435,N_17475,N_17446);
nor U18436 (N_18436,N_17911,N_17820);
or U18437 (N_18437,N_17673,N_17545);
and U18438 (N_18438,N_17679,N_17836);
or U18439 (N_18439,N_17487,N_17602);
and U18440 (N_18440,N_17652,N_17439);
or U18441 (N_18441,N_17494,N_17625);
or U18442 (N_18442,N_17660,N_17546);
or U18443 (N_18443,N_17716,N_17658);
nand U18444 (N_18444,N_17823,N_17828);
and U18445 (N_18445,N_17630,N_17944);
or U18446 (N_18446,N_17755,N_17953);
or U18447 (N_18447,N_17926,N_17977);
nand U18448 (N_18448,N_17428,N_17674);
and U18449 (N_18449,N_17521,N_17779);
or U18450 (N_18450,N_17870,N_17423);
nand U18451 (N_18451,N_17482,N_17865);
or U18452 (N_18452,N_17411,N_17696);
nand U18453 (N_18453,N_17870,N_17818);
nand U18454 (N_18454,N_17812,N_17453);
or U18455 (N_18455,N_17894,N_17592);
or U18456 (N_18456,N_17857,N_17836);
xnor U18457 (N_18457,N_17945,N_17859);
or U18458 (N_18458,N_17813,N_17751);
nand U18459 (N_18459,N_17427,N_17870);
or U18460 (N_18460,N_17657,N_17409);
or U18461 (N_18461,N_17847,N_17841);
nor U18462 (N_18462,N_17704,N_17905);
nor U18463 (N_18463,N_17816,N_17947);
nor U18464 (N_18464,N_17430,N_17822);
nand U18465 (N_18465,N_17757,N_17902);
nand U18466 (N_18466,N_17627,N_17865);
nor U18467 (N_18467,N_17961,N_17866);
and U18468 (N_18468,N_17702,N_17739);
nand U18469 (N_18469,N_17597,N_17839);
or U18470 (N_18470,N_17917,N_17799);
and U18471 (N_18471,N_17715,N_17929);
nand U18472 (N_18472,N_17698,N_17959);
and U18473 (N_18473,N_17878,N_17837);
nand U18474 (N_18474,N_17978,N_17758);
nand U18475 (N_18475,N_17642,N_17911);
nand U18476 (N_18476,N_17430,N_17653);
or U18477 (N_18477,N_17900,N_17929);
or U18478 (N_18478,N_17736,N_17841);
nor U18479 (N_18479,N_17981,N_17984);
nand U18480 (N_18480,N_17461,N_17428);
nor U18481 (N_18481,N_17466,N_17590);
and U18482 (N_18482,N_17652,N_17419);
or U18483 (N_18483,N_17606,N_17475);
nand U18484 (N_18484,N_17964,N_17837);
or U18485 (N_18485,N_17512,N_17475);
nor U18486 (N_18486,N_17852,N_17716);
and U18487 (N_18487,N_17635,N_17709);
nor U18488 (N_18488,N_17489,N_17871);
nand U18489 (N_18489,N_17739,N_17855);
nand U18490 (N_18490,N_17937,N_17818);
nand U18491 (N_18491,N_17410,N_17476);
nor U18492 (N_18492,N_17462,N_17404);
nand U18493 (N_18493,N_17863,N_17526);
nand U18494 (N_18494,N_17442,N_17992);
and U18495 (N_18495,N_17525,N_17831);
nor U18496 (N_18496,N_17836,N_17624);
nor U18497 (N_18497,N_17789,N_17847);
nor U18498 (N_18498,N_17764,N_17467);
xor U18499 (N_18499,N_17649,N_17482);
and U18500 (N_18500,N_17753,N_17735);
and U18501 (N_18501,N_17552,N_17501);
and U18502 (N_18502,N_17654,N_17432);
nand U18503 (N_18503,N_17482,N_17607);
nand U18504 (N_18504,N_17827,N_17466);
and U18505 (N_18505,N_17691,N_17478);
nand U18506 (N_18506,N_17914,N_17595);
nand U18507 (N_18507,N_17639,N_17786);
nand U18508 (N_18508,N_17821,N_17450);
or U18509 (N_18509,N_17645,N_17792);
nand U18510 (N_18510,N_17741,N_17942);
nor U18511 (N_18511,N_17812,N_17701);
nand U18512 (N_18512,N_17965,N_17781);
or U18513 (N_18513,N_17408,N_17491);
nand U18514 (N_18514,N_17783,N_17743);
and U18515 (N_18515,N_17688,N_17889);
xor U18516 (N_18516,N_17880,N_17679);
xnor U18517 (N_18517,N_17740,N_17646);
or U18518 (N_18518,N_17893,N_17840);
and U18519 (N_18519,N_17516,N_17770);
xnor U18520 (N_18520,N_17956,N_17917);
nand U18521 (N_18521,N_17950,N_17712);
nand U18522 (N_18522,N_17724,N_17942);
and U18523 (N_18523,N_17865,N_17420);
and U18524 (N_18524,N_17434,N_17786);
nor U18525 (N_18525,N_17994,N_17464);
nand U18526 (N_18526,N_17509,N_17446);
and U18527 (N_18527,N_17957,N_17948);
or U18528 (N_18528,N_17407,N_17849);
or U18529 (N_18529,N_17795,N_17588);
nor U18530 (N_18530,N_17847,N_17927);
nand U18531 (N_18531,N_17864,N_17880);
and U18532 (N_18532,N_17782,N_17511);
nor U18533 (N_18533,N_17966,N_17427);
or U18534 (N_18534,N_17731,N_17809);
nand U18535 (N_18535,N_17650,N_17603);
or U18536 (N_18536,N_17981,N_17923);
nand U18537 (N_18537,N_17580,N_17715);
nand U18538 (N_18538,N_17925,N_17460);
nand U18539 (N_18539,N_17881,N_17787);
nand U18540 (N_18540,N_17797,N_17918);
and U18541 (N_18541,N_17764,N_17718);
nor U18542 (N_18542,N_17717,N_17588);
or U18543 (N_18543,N_17913,N_17737);
nand U18544 (N_18544,N_17805,N_17686);
and U18545 (N_18545,N_17432,N_17668);
nor U18546 (N_18546,N_17644,N_17821);
and U18547 (N_18547,N_17856,N_17770);
nor U18548 (N_18548,N_17752,N_17415);
xnor U18549 (N_18549,N_17605,N_17944);
nor U18550 (N_18550,N_17465,N_17562);
or U18551 (N_18551,N_17604,N_17743);
or U18552 (N_18552,N_17661,N_17669);
or U18553 (N_18553,N_17806,N_17764);
nor U18554 (N_18554,N_17895,N_17553);
nand U18555 (N_18555,N_17770,N_17498);
and U18556 (N_18556,N_17565,N_17527);
xor U18557 (N_18557,N_17938,N_17699);
nand U18558 (N_18558,N_17999,N_17488);
nand U18559 (N_18559,N_17527,N_17628);
and U18560 (N_18560,N_17765,N_17790);
nand U18561 (N_18561,N_17864,N_17640);
nand U18562 (N_18562,N_17812,N_17804);
or U18563 (N_18563,N_17428,N_17784);
nand U18564 (N_18564,N_17642,N_17850);
nand U18565 (N_18565,N_17513,N_17647);
and U18566 (N_18566,N_17400,N_17439);
nand U18567 (N_18567,N_17461,N_17674);
nand U18568 (N_18568,N_17654,N_17428);
nand U18569 (N_18569,N_17457,N_17975);
nor U18570 (N_18570,N_17705,N_17534);
and U18571 (N_18571,N_17731,N_17759);
and U18572 (N_18572,N_17789,N_17930);
and U18573 (N_18573,N_17619,N_17537);
xor U18574 (N_18574,N_17646,N_17636);
xor U18575 (N_18575,N_17614,N_17476);
nor U18576 (N_18576,N_17919,N_17968);
nor U18577 (N_18577,N_17749,N_17776);
nand U18578 (N_18578,N_17445,N_17918);
and U18579 (N_18579,N_17451,N_17766);
nand U18580 (N_18580,N_17708,N_17465);
nand U18581 (N_18581,N_17878,N_17470);
nand U18582 (N_18582,N_17999,N_17562);
or U18583 (N_18583,N_17918,N_17447);
nand U18584 (N_18584,N_17989,N_17590);
xor U18585 (N_18585,N_17942,N_17653);
nand U18586 (N_18586,N_17891,N_17528);
or U18587 (N_18587,N_17887,N_17918);
nand U18588 (N_18588,N_17491,N_17745);
and U18589 (N_18589,N_17832,N_17645);
or U18590 (N_18590,N_17747,N_17935);
nand U18591 (N_18591,N_17709,N_17639);
and U18592 (N_18592,N_17645,N_17817);
or U18593 (N_18593,N_17871,N_17961);
and U18594 (N_18594,N_17707,N_17836);
nand U18595 (N_18595,N_17749,N_17847);
nand U18596 (N_18596,N_17907,N_17547);
and U18597 (N_18597,N_17999,N_17691);
or U18598 (N_18598,N_17616,N_17833);
nor U18599 (N_18599,N_17662,N_17951);
nand U18600 (N_18600,N_18487,N_18215);
or U18601 (N_18601,N_18159,N_18370);
nand U18602 (N_18602,N_18194,N_18076);
and U18603 (N_18603,N_18123,N_18516);
or U18604 (N_18604,N_18517,N_18584);
and U18605 (N_18605,N_18548,N_18237);
nand U18606 (N_18606,N_18325,N_18431);
or U18607 (N_18607,N_18497,N_18475);
or U18608 (N_18608,N_18334,N_18445);
or U18609 (N_18609,N_18054,N_18234);
and U18610 (N_18610,N_18522,N_18449);
nor U18611 (N_18611,N_18221,N_18037);
nor U18612 (N_18612,N_18326,N_18205);
and U18613 (N_18613,N_18314,N_18147);
nand U18614 (N_18614,N_18319,N_18353);
or U18615 (N_18615,N_18161,N_18316);
nor U18616 (N_18616,N_18012,N_18141);
nor U18617 (N_18617,N_18398,N_18381);
and U18618 (N_18618,N_18294,N_18178);
nand U18619 (N_18619,N_18007,N_18503);
and U18620 (N_18620,N_18592,N_18324);
xor U18621 (N_18621,N_18167,N_18179);
or U18622 (N_18622,N_18013,N_18391);
or U18623 (N_18623,N_18373,N_18127);
nor U18624 (N_18624,N_18439,N_18595);
or U18625 (N_18625,N_18590,N_18002);
and U18626 (N_18626,N_18022,N_18130);
nand U18627 (N_18627,N_18155,N_18392);
and U18628 (N_18628,N_18483,N_18533);
nor U18629 (N_18629,N_18502,N_18303);
or U18630 (N_18630,N_18200,N_18249);
nor U18631 (N_18631,N_18597,N_18171);
nand U18632 (N_18632,N_18331,N_18121);
and U18633 (N_18633,N_18586,N_18486);
and U18634 (N_18634,N_18419,N_18132);
or U18635 (N_18635,N_18423,N_18558);
nand U18636 (N_18636,N_18114,N_18403);
and U18637 (N_18637,N_18466,N_18096);
or U18638 (N_18638,N_18542,N_18067);
nor U18639 (N_18639,N_18387,N_18573);
nor U18640 (N_18640,N_18153,N_18519);
nand U18641 (N_18641,N_18404,N_18014);
nand U18642 (N_18642,N_18284,N_18248);
or U18643 (N_18643,N_18520,N_18115);
and U18644 (N_18644,N_18189,N_18490);
nand U18645 (N_18645,N_18023,N_18426);
or U18646 (N_18646,N_18265,N_18357);
and U18647 (N_18647,N_18446,N_18031);
or U18648 (N_18648,N_18344,N_18036);
or U18649 (N_18649,N_18062,N_18436);
or U18650 (N_18650,N_18264,N_18024);
nand U18651 (N_18651,N_18228,N_18238);
xnor U18652 (N_18652,N_18382,N_18322);
nor U18653 (N_18653,N_18343,N_18187);
nand U18654 (N_18654,N_18409,N_18274);
nand U18655 (N_18655,N_18420,N_18296);
and U18656 (N_18656,N_18244,N_18534);
and U18657 (N_18657,N_18152,N_18511);
nand U18658 (N_18658,N_18256,N_18089);
nor U18659 (N_18659,N_18253,N_18546);
nand U18660 (N_18660,N_18126,N_18488);
or U18661 (N_18661,N_18226,N_18307);
nor U18662 (N_18662,N_18437,N_18364);
nand U18663 (N_18663,N_18148,N_18113);
or U18664 (N_18664,N_18273,N_18090);
nor U18665 (N_18665,N_18050,N_18207);
and U18666 (N_18666,N_18251,N_18321);
nand U18667 (N_18667,N_18538,N_18415);
or U18668 (N_18668,N_18111,N_18416);
or U18669 (N_18669,N_18323,N_18480);
nor U18670 (N_18670,N_18544,N_18169);
or U18671 (N_18671,N_18367,N_18242);
nor U18672 (N_18672,N_18125,N_18029);
nand U18673 (N_18673,N_18046,N_18588);
nand U18674 (N_18674,N_18421,N_18471);
or U18675 (N_18675,N_18317,N_18020);
nand U18676 (N_18676,N_18192,N_18501);
or U18677 (N_18677,N_18241,N_18377);
nand U18678 (N_18678,N_18025,N_18260);
nor U18679 (N_18679,N_18414,N_18330);
nor U18680 (N_18680,N_18550,N_18509);
and U18681 (N_18681,N_18453,N_18202);
and U18682 (N_18682,N_18191,N_18557);
or U18683 (N_18683,N_18079,N_18175);
nand U18684 (N_18684,N_18341,N_18227);
nand U18685 (N_18685,N_18578,N_18120);
or U18686 (N_18686,N_18271,N_18482);
nand U18687 (N_18687,N_18231,N_18400);
xor U18688 (N_18688,N_18019,N_18374);
and U18689 (N_18689,N_18072,N_18492);
nand U18690 (N_18690,N_18252,N_18094);
nor U18691 (N_18691,N_18363,N_18554);
nand U18692 (N_18692,N_18468,N_18240);
or U18693 (N_18693,N_18073,N_18560);
nand U18694 (N_18694,N_18499,N_18267);
or U18695 (N_18695,N_18407,N_18218);
and U18696 (N_18696,N_18591,N_18572);
nand U18697 (N_18697,N_18006,N_18394);
or U18698 (N_18698,N_18185,N_18411);
nand U18699 (N_18699,N_18477,N_18320);
or U18700 (N_18700,N_18077,N_18430);
nand U18701 (N_18701,N_18478,N_18461);
nor U18702 (N_18702,N_18318,N_18124);
nand U18703 (N_18703,N_18368,N_18385);
nand U18704 (N_18704,N_18513,N_18579);
and U18705 (N_18705,N_18122,N_18063);
nand U18706 (N_18706,N_18236,N_18432);
nand U18707 (N_18707,N_18038,N_18360);
and U18708 (N_18708,N_18220,N_18366);
or U18709 (N_18709,N_18386,N_18058);
nor U18710 (N_18710,N_18258,N_18304);
nand U18711 (N_18711,N_18261,N_18042);
or U18712 (N_18712,N_18116,N_18406);
nor U18713 (N_18713,N_18379,N_18075);
nand U18714 (N_18714,N_18301,N_18535);
nand U18715 (N_18715,N_18547,N_18243);
or U18716 (N_18716,N_18064,N_18142);
and U18717 (N_18717,N_18388,N_18532);
nand U18718 (N_18718,N_18108,N_18540);
nand U18719 (N_18719,N_18145,N_18092);
nor U18720 (N_18720,N_18206,N_18541);
nor U18721 (N_18721,N_18225,N_18199);
and U18722 (N_18722,N_18340,N_18208);
nand U18723 (N_18723,N_18348,N_18515);
nor U18724 (N_18724,N_18310,N_18279);
nand U18725 (N_18725,N_18582,N_18137);
nand U18726 (N_18726,N_18055,N_18507);
and U18727 (N_18727,N_18418,N_18447);
or U18728 (N_18728,N_18168,N_18444);
or U18729 (N_18729,N_18508,N_18051);
and U18730 (N_18730,N_18091,N_18107);
nand U18731 (N_18731,N_18160,N_18245);
nor U18732 (N_18732,N_18278,N_18459);
and U18733 (N_18733,N_18395,N_18569);
xnor U18734 (N_18734,N_18052,N_18441);
and U18735 (N_18735,N_18448,N_18427);
and U18736 (N_18736,N_18552,N_18559);
and U18737 (N_18737,N_18181,N_18371);
nor U18738 (N_18738,N_18105,N_18018);
or U18739 (N_18739,N_18287,N_18170);
and U18740 (N_18740,N_18543,N_18496);
or U18741 (N_18741,N_18053,N_18070);
xnor U18742 (N_18742,N_18306,N_18095);
nand U18743 (N_18743,N_18425,N_18040);
and U18744 (N_18744,N_18383,N_18537);
nor U18745 (N_18745,N_18526,N_18250);
or U18746 (N_18746,N_18442,N_18378);
nor U18747 (N_18747,N_18246,N_18026);
or U18748 (N_18748,N_18282,N_18044);
and U18749 (N_18749,N_18080,N_18346);
nand U18750 (N_18750,N_18131,N_18570);
or U18751 (N_18751,N_18109,N_18596);
or U18752 (N_18752,N_18585,N_18097);
and U18753 (N_18753,N_18083,N_18259);
nor U18754 (N_18754,N_18283,N_18299);
or U18755 (N_18755,N_18372,N_18438);
nor U18756 (N_18756,N_18295,N_18566);
nor U18757 (N_18757,N_18350,N_18078);
and U18758 (N_18758,N_18197,N_18232);
nand U18759 (N_18759,N_18165,N_18593);
nand U18760 (N_18760,N_18001,N_18521);
and U18761 (N_18761,N_18104,N_18587);
nor U18762 (N_18762,N_18233,N_18146);
or U18763 (N_18763,N_18361,N_18337);
nor U18764 (N_18764,N_18086,N_18292);
nand U18765 (N_18765,N_18247,N_18057);
or U18766 (N_18766,N_18598,N_18305);
nand U18767 (N_18767,N_18158,N_18276);
or U18768 (N_18768,N_18405,N_18136);
nand U18769 (N_18769,N_18429,N_18450);
or U18770 (N_18770,N_18525,N_18069);
or U18771 (N_18771,N_18129,N_18150);
nand U18772 (N_18772,N_18216,N_18098);
nor U18773 (N_18773,N_18166,N_18177);
nor U18774 (N_18774,N_18047,N_18465);
or U18775 (N_18775,N_18163,N_18365);
nor U18776 (N_18776,N_18359,N_18494);
or U18777 (N_18777,N_18568,N_18571);
nor U18778 (N_18778,N_18529,N_18339);
and U18779 (N_18779,N_18134,N_18384);
and U18780 (N_18780,N_18354,N_18204);
nand U18781 (N_18781,N_18143,N_18190);
nand U18782 (N_18782,N_18201,N_18369);
or U18783 (N_18783,N_18003,N_18255);
nor U18784 (N_18784,N_18176,N_18342);
nand U18785 (N_18785,N_18224,N_18327);
nor U18786 (N_18786,N_18032,N_18068);
nand U18787 (N_18787,N_18281,N_18180);
nand U18788 (N_18788,N_18017,N_18056);
and U18789 (N_18789,N_18476,N_18061);
nor U18790 (N_18790,N_18308,N_18085);
xnor U18791 (N_18791,N_18352,N_18048);
nand U18792 (N_18792,N_18112,N_18151);
and U18793 (N_18793,N_18523,N_18100);
or U18794 (N_18794,N_18375,N_18581);
or U18795 (N_18795,N_18117,N_18213);
and U18796 (N_18796,N_18157,N_18034);
or U18797 (N_18797,N_18211,N_18082);
xor U18798 (N_18798,N_18272,N_18060);
nor U18799 (N_18799,N_18333,N_18280);
nand U18800 (N_18800,N_18580,N_18474);
or U18801 (N_18801,N_18088,N_18144);
or U18802 (N_18802,N_18410,N_18235);
or U18803 (N_18803,N_18209,N_18135);
nor U18804 (N_18804,N_18495,N_18196);
nor U18805 (N_18805,N_18536,N_18210);
or U18806 (N_18806,N_18000,N_18093);
nand U18807 (N_18807,N_18473,N_18099);
or U18808 (N_18808,N_18349,N_18084);
nor U18809 (N_18809,N_18285,N_18428);
nand U18810 (N_18810,N_18277,N_18239);
xnor U18811 (N_18811,N_18556,N_18356);
or U18812 (N_18812,N_18298,N_18589);
and U18813 (N_18813,N_18291,N_18101);
nand U18814 (N_18814,N_18103,N_18469);
xor U18815 (N_18815,N_18574,N_18005);
and U18816 (N_18816,N_18183,N_18376);
or U18817 (N_18817,N_18312,N_18186);
and U18818 (N_18818,N_18565,N_18045);
nor U18819 (N_18819,N_18545,N_18182);
nand U18820 (N_18820,N_18351,N_18119);
and U18821 (N_18821,N_18254,N_18464);
nor U18822 (N_18822,N_18010,N_18214);
nor U18823 (N_18823,N_18358,N_18309);
or U18824 (N_18824,N_18266,N_18493);
or U18825 (N_18825,N_18128,N_18451);
and U18826 (N_18826,N_18066,N_18422);
nand U18827 (N_18827,N_18412,N_18164);
or U18828 (N_18828,N_18454,N_18424);
nor U18829 (N_18829,N_18230,N_18049);
or U18830 (N_18830,N_18399,N_18564);
nand U18831 (N_18831,N_18184,N_18195);
and U18832 (N_18832,N_18397,N_18462);
nor U18833 (N_18833,N_18173,N_18472);
or U18834 (N_18834,N_18527,N_18401);
and U18835 (N_18835,N_18539,N_18059);
nor U18836 (N_18836,N_18288,N_18463);
nor U18837 (N_18837,N_18222,N_18498);
nand U18838 (N_18838,N_18074,N_18408);
and U18839 (N_18839,N_18268,N_18455);
or U18840 (N_18840,N_18355,N_18203);
nor U18841 (N_18841,N_18149,N_18393);
nor U18842 (N_18842,N_18081,N_18110);
nor U18843 (N_18843,N_18484,N_18016);
nor U18844 (N_18844,N_18599,N_18440);
and U18845 (N_18845,N_18457,N_18506);
nor U18846 (N_18846,N_18332,N_18275);
nor U18847 (N_18847,N_18362,N_18435);
xnor U18848 (N_18848,N_18188,N_18315);
and U18849 (N_18849,N_18479,N_18156);
nor U18850 (N_18850,N_18027,N_18297);
or U18851 (N_18851,N_18500,N_18302);
or U18852 (N_18852,N_18300,N_18417);
nand U18853 (N_18853,N_18561,N_18229);
and U18854 (N_18854,N_18467,N_18594);
and U18855 (N_18855,N_18345,N_18021);
or U18856 (N_18856,N_18139,N_18504);
nand U18857 (N_18857,N_18217,N_18133);
or U18858 (N_18858,N_18293,N_18286);
nand U18859 (N_18859,N_18434,N_18174);
nor U18860 (N_18860,N_18263,N_18270);
and U18861 (N_18861,N_18172,N_18512);
nand U18862 (N_18862,N_18389,N_18329);
nor U18863 (N_18863,N_18396,N_18162);
nand U18864 (N_18864,N_18562,N_18481);
and U18865 (N_18865,N_18269,N_18118);
nor U18866 (N_18866,N_18380,N_18262);
and U18867 (N_18867,N_18518,N_18553);
nor U18868 (N_18868,N_18413,N_18030);
xor U18869 (N_18869,N_18402,N_18071);
or U18870 (N_18870,N_18335,N_18290);
nand U18871 (N_18871,N_18041,N_18140);
and U18872 (N_18872,N_18530,N_18456);
nor U18873 (N_18873,N_18313,N_18138);
and U18874 (N_18874,N_18154,N_18555);
nand U18875 (N_18875,N_18433,N_18039);
nor U18876 (N_18876,N_18328,N_18524);
nor U18877 (N_18877,N_18011,N_18458);
nor U18878 (N_18878,N_18087,N_18193);
xor U18879 (N_18879,N_18452,N_18491);
nand U18880 (N_18880,N_18485,N_18549);
or U18881 (N_18881,N_18575,N_18223);
nand U18882 (N_18882,N_18576,N_18460);
nand U18883 (N_18883,N_18583,N_18028);
and U18884 (N_18884,N_18008,N_18514);
and U18885 (N_18885,N_18338,N_18489);
nand U18886 (N_18886,N_18443,N_18567);
nand U18887 (N_18887,N_18004,N_18065);
and U18888 (N_18888,N_18336,N_18505);
or U18889 (N_18889,N_18219,N_18531);
nor U18890 (N_18890,N_18289,N_18510);
and U18891 (N_18891,N_18106,N_18043);
nor U18892 (N_18892,N_18033,N_18347);
nor U18893 (N_18893,N_18563,N_18390);
and U18894 (N_18894,N_18311,N_18015);
or U18895 (N_18895,N_18577,N_18551);
nor U18896 (N_18896,N_18212,N_18198);
or U18897 (N_18897,N_18009,N_18035);
or U18898 (N_18898,N_18257,N_18528);
and U18899 (N_18899,N_18470,N_18102);
nand U18900 (N_18900,N_18165,N_18067);
and U18901 (N_18901,N_18259,N_18207);
nor U18902 (N_18902,N_18170,N_18258);
nor U18903 (N_18903,N_18483,N_18556);
nor U18904 (N_18904,N_18358,N_18433);
or U18905 (N_18905,N_18483,N_18221);
or U18906 (N_18906,N_18494,N_18219);
nor U18907 (N_18907,N_18300,N_18333);
or U18908 (N_18908,N_18083,N_18078);
nor U18909 (N_18909,N_18022,N_18008);
nand U18910 (N_18910,N_18115,N_18021);
nand U18911 (N_18911,N_18370,N_18136);
nor U18912 (N_18912,N_18386,N_18086);
or U18913 (N_18913,N_18262,N_18357);
nor U18914 (N_18914,N_18312,N_18090);
and U18915 (N_18915,N_18332,N_18203);
and U18916 (N_18916,N_18548,N_18560);
and U18917 (N_18917,N_18428,N_18336);
nor U18918 (N_18918,N_18303,N_18211);
nand U18919 (N_18919,N_18522,N_18277);
and U18920 (N_18920,N_18218,N_18168);
and U18921 (N_18921,N_18485,N_18116);
nand U18922 (N_18922,N_18465,N_18449);
nor U18923 (N_18923,N_18485,N_18274);
nand U18924 (N_18924,N_18042,N_18555);
nor U18925 (N_18925,N_18565,N_18108);
xnor U18926 (N_18926,N_18577,N_18455);
nand U18927 (N_18927,N_18035,N_18098);
and U18928 (N_18928,N_18104,N_18008);
or U18929 (N_18929,N_18496,N_18426);
or U18930 (N_18930,N_18142,N_18400);
nand U18931 (N_18931,N_18219,N_18544);
nand U18932 (N_18932,N_18203,N_18177);
or U18933 (N_18933,N_18284,N_18012);
or U18934 (N_18934,N_18081,N_18233);
and U18935 (N_18935,N_18419,N_18371);
nand U18936 (N_18936,N_18008,N_18279);
nor U18937 (N_18937,N_18351,N_18504);
nor U18938 (N_18938,N_18500,N_18436);
nor U18939 (N_18939,N_18510,N_18472);
nand U18940 (N_18940,N_18547,N_18392);
nand U18941 (N_18941,N_18318,N_18553);
nand U18942 (N_18942,N_18197,N_18312);
or U18943 (N_18943,N_18216,N_18596);
and U18944 (N_18944,N_18170,N_18044);
nor U18945 (N_18945,N_18097,N_18061);
nand U18946 (N_18946,N_18545,N_18363);
or U18947 (N_18947,N_18555,N_18279);
and U18948 (N_18948,N_18548,N_18148);
nor U18949 (N_18949,N_18265,N_18189);
nand U18950 (N_18950,N_18012,N_18072);
and U18951 (N_18951,N_18347,N_18332);
nor U18952 (N_18952,N_18492,N_18143);
xnor U18953 (N_18953,N_18269,N_18166);
and U18954 (N_18954,N_18369,N_18055);
nor U18955 (N_18955,N_18224,N_18589);
or U18956 (N_18956,N_18538,N_18308);
and U18957 (N_18957,N_18424,N_18548);
or U18958 (N_18958,N_18038,N_18090);
nor U18959 (N_18959,N_18007,N_18183);
and U18960 (N_18960,N_18354,N_18576);
nand U18961 (N_18961,N_18201,N_18342);
and U18962 (N_18962,N_18321,N_18183);
and U18963 (N_18963,N_18371,N_18473);
nand U18964 (N_18964,N_18476,N_18404);
and U18965 (N_18965,N_18251,N_18160);
nand U18966 (N_18966,N_18415,N_18571);
nor U18967 (N_18967,N_18519,N_18108);
or U18968 (N_18968,N_18548,N_18326);
and U18969 (N_18969,N_18351,N_18202);
nand U18970 (N_18970,N_18020,N_18098);
nand U18971 (N_18971,N_18139,N_18091);
nor U18972 (N_18972,N_18160,N_18588);
nor U18973 (N_18973,N_18033,N_18103);
and U18974 (N_18974,N_18300,N_18337);
and U18975 (N_18975,N_18498,N_18455);
and U18976 (N_18976,N_18088,N_18038);
or U18977 (N_18977,N_18577,N_18576);
or U18978 (N_18978,N_18416,N_18351);
and U18979 (N_18979,N_18267,N_18132);
nor U18980 (N_18980,N_18236,N_18026);
and U18981 (N_18981,N_18118,N_18240);
nor U18982 (N_18982,N_18127,N_18300);
and U18983 (N_18983,N_18342,N_18395);
and U18984 (N_18984,N_18159,N_18386);
nor U18985 (N_18985,N_18089,N_18552);
or U18986 (N_18986,N_18189,N_18227);
nand U18987 (N_18987,N_18450,N_18101);
and U18988 (N_18988,N_18330,N_18343);
and U18989 (N_18989,N_18303,N_18534);
and U18990 (N_18990,N_18046,N_18525);
nor U18991 (N_18991,N_18149,N_18398);
xor U18992 (N_18992,N_18356,N_18491);
and U18993 (N_18993,N_18151,N_18208);
and U18994 (N_18994,N_18574,N_18347);
nor U18995 (N_18995,N_18456,N_18192);
nand U18996 (N_18996,N_18334,N_18349);
nand U18997 (N_18997,N_18135,N_18581);
xor U18998 (N_18998,N_18409,N_18500);
or U18999 (N_18999,N_18454,N_18595);
xor U19000 (N_19000,N_18359,N_18074);
nor U19001 (N_19001,N_18548,N_18356);
nand U19002 (N_19002,N_18429,N_18425);
or U19003 (N_19003,N_18080,N_18599);
and U19004 (N_19004,N_18122,N_18464);
or U19005 (N_19005,N_18408,N_18244);
or U19006 (N_19006,N_18029,N_18582);
nand U19007 (N_19007,N_18308,N_18171);
xnor U19008 (N_19008,N_18248,N_18224);
nand U19009 (N_19009,N_18457,N_18256);
or U19010 (N_19010,N_18513,N_18590);
nand U19011 (N_19011,N_18199,N_18045);
and U19012 (N_19012,N_18225,N_18118);
and U19013 (N_19013,N_18206,N_18268);
and U19014 (N_19014,N_18170,N_18322);
or U19015 (N_19015,N_18477,N_18373);
nand U19016 (N_19016,N_18517,N_18102);
nand U19017 (N_19017,N_18343,N_18361);
and U19018 (N_19018,N_18512,N_18450);
nor U19019 (N_19019,N_18523,N_18073);
and U19020 (N_19020,N_18564,N_18143);
and U19021 (N_19021,N_18030,N_18259);
and U19022 (N_19022,N_18403,N_18045);
or U19023 (N_19023,N_18118,N_18157);
or U19024 (N_19024,N_18365,N_18221);
nand U19025 (N_19025,N_18360,N_18255);
or U19026 (N_19026,N_18048,N_18040);
or U19027 (N_19027,N_18459,N_18000);
and U19028 (N_19028,N_18125,N_18445);
or U19029 (N_19029,N_18409,N_18503);
or U19030 (N_19030,N_18096,N_18509);
nand U19031 (N_19031,N_18475,N_18383);
nand U19032 (N_19032,N_18562,N_18207);
or U19033 (N_19033,N_18552,N_18450);
or U19034 (N_19034,N_18279,N_18465);
nor U19035 (N_19035,N_18218,N_18332);
or U19036 (N_19036,N_18371,N_18138);
and U19037 (N_19037,N_18489,N_18425);
or U19038 (N_19038,N_18542,N_18281);
nand U19039 (N_19039,N_18106,N_18529);
or U19040 (N_19040,N_18426,N_18593);
nor U19041 (N_19041,N_18489,N_18530);
and U19042 (N_19042,N_18395,N_18176);
and U19043 (N_19043,N_18288,N_18338);
nor U19044 (N_19044,N_18513,N_18536);
nand U19045 (N_19045,N_18210,N_18318);
nor U19046 (N_19046,N_18435,N_18442);
nor U19047 (N_19047,N_18585,N_18530);
nor U19048 (N_19048,N_18126,N_18038);
nand U19049 (N_19049,N_18321,N_18463);
nor U19050 (N_19050,N_18278,N_18241);
or U19051 (N_19051,N_18116,N_18214);
nand U19052 (N_19052,N_18495,N_18480);
or U19053 (N_19053,N_18447,N_18202);
nor U19054 (N_19054,N_18132,N_18342);
nor U19055 (N_19055,N_18487,N_18243);
and U19056 (N_19056,N_18086,N_18077);
or U19057 (N_19057,N_18512,N_18170);
and U19058 (N_19058,N_18383,N_18384);
and U19059 (N_19059,N_18117,N_18457);
and U19060 (N_19060,N_18217,N_18584);
and U19061 (N_19061,N_18239,N_18406);
nor U19062 (N_19062,N_18234,N_18561);
and U19063 (N_19063,N_18507,N_18333);
or U19064 (N_19064,N_18004,N_18326);
and U19065 (N_19065,N_18431,N_18299);
and U19066 (N_19066,N_18517,N_18556);
and U19067 (N_19067,N_18001,N_18353);
nor U19068 (N_19068,N_18494,N_18403);
nand U19069 (N_19069,N_18022,N_18364);
and U19070 (N_19070,N_18069,N_18255);
nand U19071 (N_19071,N_18429,N_18390);
or U19072 (N_19072,N_18149,N_18569);
or U19073 (N_19073,N_18470,N_18345);
and U19074 (N_19074,N_18143,N_18151);
xnor U19075 (N_19075,N_18044,N_18598);
and U19076 (N_19076,N_18089,N_18257);
or U19077 (N_19077,N_18311,N_18319);
xnor U19078 (N_19078,N_18539,N_18071);
xnor U19079 (N_19079,N_18494,N_18228);
nor U19080 (N_19080,N_18301,N_18201);
and U19081 (N_19081,N_18588,N_18253);
and U19082 (N_19082,N_18198,N_18495);
and U19083 (N_19083,N_18124,N_18257);
nor U19084 (N_19084,N_18524,N_18372);
and U19085 (N_19085,N_18578,N_18421);
nor U19086 (N_19086,N_18454,N_18234);
nand U19087 (N_19087,N_18106,N_18523);
nor U19088 (N_19088,N_18228,N_18290);
nand U19089 (N_19089,N_18415,N_18201);
nand U19090 (N_19090,N_18285,N_18045);
or U19091 (N_19091,N_18130,N_18270);
nand U19092 (N_19092,N_18388,N_18306);
nor U19093 (N_19093,N_18578,N_18230);
nand U19094 (N_19094,N_18395,N_18467);
or U19095 (N_19095,N_18172,N_18124);
nor U19096 (N_19096,N_18458,N_18002);
or U19097 (N_19097,N_18108,N_18452);
nand U19098 (N_19098,N_18214,N_18033);
nor U19099 (N_19099,N_18117,N_18235);
or U19100 (N_19100,N_18016,N_18403);
and U19101 (N_19101,N_18024,N_18327);
and U19102 (N_19102,N_18286,N_18198);
nand U19103 (N_19103,N_18555,N_18032);
or U19104 (N_19104,N_18573,N_18393);
or U19105 (N_19105,N_18520,N_18289);
nor U19106 (N_19106,N_18189,N_18371);
xnor U19107 (N_19107,N_18117,N_18376);
and U19108 (N_19108,N_18070,N_18123);
and U19109 (N_19109,N_18158,N_18031);
nand U19110 (N_19110,N_18265,N_18100);
nor U19111 (N_19111,N_18529,N_18207);
or U19112 (N_19112,N_18149,N_18375);
nand U19113 (N_19113,N_18331,N_18117);
xor U19114 (N_19114,N_18260,N_18332);
xor U19115 (N_19115,N_18496,N_18243);
or U19116 (N_19116,N_18043,N_18283);
and U19117 (N_19117,N_18249,N_18127);
nor U19118 (N_19118,N_18029,N_18555);
and U19119 (N_19119,N_18441,N_18369);
nand U19120 (N_19120,N_18308,N_18290);
xnor U19121 (N_19121,N_18103,N_18097);
or U19122 (N_19122,N_18040,N_18442);
or U19123 (N_19123,N_18205,N_18223);
nand U19124 (N_19124,N_18256,N_18370);
xor U19125 (N_19125,N_18188,N_18340);
nand U19126 (N_19126,N_18342,N_18044);
nor U19127 (N_19127,N_18033,N_18583);
and U19128 (N_19128,N_18423,N_18404);
and U19129 (N_19129,N_18279,N_18296);
nor U19130 (N_19130,N_18517,N_18423);
and U19131 (N_19131,N_18576,N_18597);
nand U19132 (N_19132,N_18049,N_18569);
nand U19133 (N_19133,N_18594,N_18464);
or U19134 (N_19134,N_18050,N_18196);
or U19135 (N_19135,N_18453,N_18138);
and U19136 (N_19136,N_18534,N_18542);
or U19137 (N_19137,N_18372,N_18319);
nor U19138 (N_19138,N_18187,N_18277);
nor U19139 (N_19139,N_18007,N_18040);
nor U19140 (N_19140,N_18369,N_18402);
or U19141 (N_19141,N_18124,N_18018);
or U19142 (N_19142,N_18445,N_18072);
nand U19143 (N_19143,N_18137,N_18139);
and U19144 (N_19144,N_18598,N_18273);
nor U19145 (N_19145,N_18034,N_18335);
and U19146 (N_19146,N_18449,N_18153);
and U19147 (N_19147,N_18307,N_18529);
nor U19148 (N_19148,N_18304,N_18203);
nor U19149 (N_19149,N_18019,N_18354);
nand U19150 (N_19150,N_18263,N_18006);
nand U19151 (N_19151,N_18057,N_18404);
nor U19152 (N_19152,N_18456,N_18136);
nor U19153 (N_19153,N_18175,N_18003);
nor U19154 (N_19154,N_18247,N_18471);
nor U19155 (N_19155,N_18157,N_18025);
or U19156 (N_19156,N_18296,N_18348);
nand U19157 (N_19157,N_18202,N_18194);
nand U19158 (N_19158,N_18157,N_18012);
nor U19159 (N_19159,N_18286,N_18347);
nor U19160 (N_19160,N_18158,N_18242);
and U19161 (N_19161,N_18075,N_18450);
or U19162 (N_19162,N_18373,N_18081);
nand U19163 (N_19163,N_18042,N_18004);
nand U19164 (N_19164,N_18465,N_18297);
nand U19165 (N_19165,N_18475,N_18247);
and U19166 (N_19166,N_18403,N_18451);
and U19167 (N_19167,N_18324,N_18314);
and U19168 (N_19168,N_18006,N_18448);
nor U19169 (N_19169,N_18186,N_18025);
or U19170 (N_19170,N_18361,N_18415);
nor U19171 (N_19171,N_18270,N_18474);
nand U19172 (N_19172,N_18498,N_18194);
or U19173 (N_19173,N_18255,N_18477);
nor U19174 (N_19174,N_18146,N_18252);
nand U19175 (N_19175,N_18176,N_18013);
xor U19176 (N_19176,N_18115,N_18043);
nand U19177 (N_19177,N_18154,N_18208);
nor U19178 (N_19178,N_18186,N_18145);
nand U19179 (N_19179,N_18246,N_18132);
and U19180 (N_19180,N_18209,N_18575);
or U19181 (N_19181,N_18019,N_18538);
and U19182 (N_19182,N_18462,N_18596);
and U19183 (N_19183,N_18330,N_18357);
nor U19184 (N_19184,N_18119,N_18198);
nand U19185 (N_19185,N_18418,N_18124);
or U19186 (N_19186,N_18478,N_18557);
nand U19187 (N_19187,N_18444,N_18079);
or U19188 (N_19188,N_18455,N_18211);
nor U19189 (N_19189,N_18041,N_18438);
nand U19190 (N_19190,N_18011,N_18002);
nor U19191 (N_19191,N_18023,N_18111);
and U19192 (N_19192,N_18327,N_18296);
or U19193 (N_19193,N_18242,N_18101);
or U19194 (N_19194,N_18049,N_18163);
or U19195 (N_19195,N_18041,N_18340);
or U19196 (N_19196,N_18385,N_18272);
nand U19197 (N_19197,N_18275,N_18315);
and U19198 (N_19198,N_18011,N_18581);
or U19199 (N_19199,N_18101,N_18054);
or U19200 (N_19200,N_18750,N_19005);
and U19201 (N_19201,N_18606,N_19142);
and U19202 (N_19202,N_19059,N_18670);
nand U19203 (N_19203,N_18863,N_19130);
xnor U19204 (N_19204,N_18788,N_18809);
and U19205 (N_19205,N_19182,N_18915);
nor U19206 (N_19206,N_18773,N_19069);
or U19207 (N_19207,N_18767,N_18785);
nor U19208 (N_19208,N_18725,N_18802);
and U19209 (N_19209,N_18826,N_18717);
nand U19210 (N_19210,N_19195,N_18793);
nand U19211 (N_19211,N_18679,N_18964);
or U19212 (N_19212,N_18739,N_18937);
xor U19213 (N_19213,N_18860,N_18790);
nand U19214 (N_19214,N_18660,N_18945);
or U19215 (N_19215,N_19099,N_18897);
nand U19216 (N_19216,N_18821,N_18962);
and U19217 (N_19217,N_18768,N_19157);
nand U19218 (N_19218,N_18819,N_18783);
nor U19219 (N_19219,N_19028,N_18676);
nand U19220 (N_19220,N_18707,N_18686);
xor U19221 (N_19221,N_18630,N_18856);
and U19222 (N_19222,N_18623,N_18695);
nand U19223 (N_19223,N_19150,N_18702);
or U19224 (N_19224,N_18633,N_18723);
and U19225 (N_19225,N_19160,N_18611);
nor U19226 (N_19226,N_18830,N_18703);
nor U19227 (N_19227,N_19025,N_18841);
and U19228 (N_19228,N_18997,N_19014);
and U19229 (N_19229,N_18942,N_19100);
and U19230 (N_19230,N_18610,N_18643);
and U19231 (N_19231,N_18982,N_19117);
and U19232 (N_19232,N_18846,N_18842);
nand U19233 (N_19233,N_19077,N_19189);
nand U19234 (N_19234,N_18824,N_18727);
or U19235 (N_19235,N_19043,N_18835);
nor U19236 (N_19236,N_18825,N_18941);
nor U19237 (N_19237,N_18672,N_18999);
xnor U19238 (N_19238,N_19023,N_18921);
or U19239 (N_19239,N_19064,N_18906);
or U19240 (N_19240,N_19048,N_18722);
and U19241 (N_19241,N_18740,N_19062);
and U19242 (N_19242,N_18614,N_19173);
nand U19243 (N_19243,N_18666,N_18652);
or U19244 (N_19244,N_18622,N_18936);
or U19245 (N_19245,N_18859,N_19111);
nor U19246 (N_19246,N_18928,N_18758);
nor U19247 (N_19247,N_19139,N_18864);
xor U19248 (N_19248,N_19041,N_18948);
nor U19249 (N_19249,N_18680,N_18957);
nor U19250 (N_19250,N_19122,N_18700);
nand U19251 (N_19251,N_18851,N_19147);
nand U19252 (N_19252,N_19013,N_18720);
and U19253 (N_19253,N_18884,N_19026);
nand U19254 (N_19254,N_19197,N_18625);
and U19255 (N_19255,N_18708,N_18668);
nor U19256 (N_19256,N_19083,N_18934);
xor U19257 (N_19257,N_18832,N_18711);
and U19258 (N_19258,N_18735,N_18744);
nand U19259 (N_19259,N_18965,N_18747);
nor U19260 (N_19260,N_19003,N_18973);
xor U19261 (N_19261,N_18857,N_19018);
nor U19262 (N_19262,N_19184,N_18728);
xnor U19263 (N_19263,N_18861,N_19183);
or U19264 (N_19264,N_19072,N_18632);
and U19265 (N_19265,N_18766,N_18724);
and U19266 (N_19266,N_19135,N_18638);
nor U19267 (N_19267,N_18902,N_18690);
or U19268 (N_19268,N_18924,N_18910);
or U19269 (N_19269,N_18960,N_19022);
nor U19270 (N_19270,N_18791,N_18913);
nor U19271 (N_19271,N_18692,N_18947);
nand U19272 (N_19272,N_18834,N_19075);
nand U19273 (N_19273,N_19019,N_18829);
or U19274 (N_19274,N_18677,N_18998);
and U19275 (N_19275,N_19109,N_18799);
nor U19276 (N_19276,N_18904,N_19012);
and U19277 (N_19277,N_18624,N_18868);
nor U19278 (N_19278,N_18866,N_19121);
nand U19279 (N_19279,N_18991,N_19124);
nor U19280 (N_19280,N_19031,N_18877);
nand U19281 (N_19281,N_18887,N_19112);
or U19282 (N_19282,N_19131,N_18975);
and U19283 (N_19283,N_19180,N_19106);
nor U19284 (N_19284,N_18737,N_19058);
and U19285 (N_19285,N_18992,N_19052);
and U19286 (N_19286,N_19015,N_19107);
nand U19287 (N_19287,N_19093,N_18981);
or U19288 (N_19288,N_18961,N_18933);
nor U19289 (N_19289,N_18971,N_19155);
or U19290 (N_19290,N_18639,N_18903);
nor U19291 (N_19291,N_18979,N_18986);
or U19292 (N_19292,N_18800,N_19020);
or U19293 (N_19293,N_19082,N_18770);
and U19294 (N_19294,N_19181,N_18881);
nor U19295 (N_19295,N_18794,N_18605);
nand U19296 (N_19296,N_18726,N_18721);
or U19297 (N_19297,N_18811,N_18876);
or U19298 (N_19298,N_19110,N_19108);
and U19299 (N_19299,N_18718,N_18810);
or U19300 (N_19300,N_19127,N_18813);
and U19301 (N_19301,N_18629,N_19071);
or U19302 (N_19302,N_19070,N_18644);
and U19303 (N_19303,N_19199,N_18763);
nor U19304 (N_19304,N_18663,N_19174);
nor U19305 (N_19305,N_18781,N_19076);
or U19306 (N_19306,N_19042,N_18940);
nand U19307 (N_19307,N_18706,N_18609);
nand U19308 (N_19308,N_18943,N_18651);
nand U19309 (N_19309,N_19159,N_18696);
or U19310 (N_19310,N_19004,N_19163);
nor U19311 (N_19311,N_18715,N_18642);
nand U19312 (N_19312,N_18917,N_18949);
and U19313 (N_19313,N_18798,N_18888);
and U19314 (N_19314,N_19033,N_18966);
and U19315 (N_19315,N_18759,N_18855);
and U19316 (N_19316,N_18963,N_18691);
and U19317 (N_19317,N_18925,N_19161);
or U19318 (N_19318,N_19191,N_18955);
or U19319 (N_19319,N_18661,N_18968);
nor U19320 (N_19320,N_18844,N_18875);
and U19321 (N_19321,N_18608,N_19177);
or U19322 (N_19322,N_18815,N_18688);
or U19323 (N_19323,N_18729,N_18653);
and U19324 (N_19324,N_18836,N_19144);
and U19325 (N_19325,N_19103,N_19166);
nand U19326 (N_19326,N_18780,N_18673);
nand U19327 (N_19327,N_18607,N_19011);
nor U19328 (N_19328,N_18847,N_18929);
and U19329 (N_19329,N_18618,N_18699);
or U19330 (N_19330,N_19178,N_19035);
nand U19331 (N_19331,N_18710,N_19185);
nor U19332 (N_19332,N_18905,N_19101);
nand U19333 (N_19333,N_18993,N_19030);
and U19334 (N_19334,N_18985,N_19009);
nor U19335 (N_19335,N_19097,N_18647);
nand U19336 (N_19336,N_18930,N_18900);
and U19337 (N_19337,N_18901,N_18619);
or U19338 (N_19338,N_18689,N_18657);
nand U19339 (N_19339,N_19128,N_18762);
nand U19340 (N_19340,N_18967,N_19036);
or U19341 (N_19341,N_18775,N_18867);
or U19342 (N_19342,N_18890,N_19024);
or U19343 (N_19343,N_18914,N_18693);
xor U19344 (N_19344,N_18922,N_18746);
nand U19345 (N_19345,N_19198,N_19039);
and U19346 (N_19346,N_18848,N_19171);
or U19347 (N_19347,N_18797,N_19186);
nor U19348 (N_19348,N_19046,N_18764);
nand U19349 (N_19349,N_19040,N_18704);
nand U19350 (N_19350,N_18786,N_19187);
nor U19351 (N_19351,N_19125,N_19190);
and U19352 (N_19352,N_18731,N_18935);
and U19353 (N_19353,N_18681,N_18812);
and U19354 (N_19354,N_18637,N_18898);
nor U19355 (N_19355,N_18946,N_18849);
or U19356 (N_19356,N_19055,N_19001);
nand U19357 (N_19357,N_18635,N_19080);
nand U19358 (N_19358,N_18926,N_18616);
nor U19359 (N_19359,N_18658,N_18678);
or U19360 (N_19360,N_18953,N_18796);
and U19361 (N_19361,N_18789,N_19169);
or U19362 (N_19362,N_18988,N_19068);
or U19363 (N_19363,N_18909,N_19132);
nand U19364 (N_19364,N_18659,N_18822);
nor U19365 (N_19365,N_18719,N_18617);
nand U19366 (N_19366,N_18886,N_18969);
and U19367 (N_19367,N_19067,N_18743);
nor U19368 (N_19368,N_19074,N_19118);
nor U19369 (N_19369,N_18774,N_18989);
and U19370 (N_19370,N_18634,N_18801);
xnor U19371 (N_19371,N_18772,N_19152);
xor U19372 (N_19372,N_18769,N_18870);
or U19373 (N_19373,N_18927,N_18983);
nand U19374 (N_19374,N_19049,N_18956);
or U19375 (N_19375,N_19193,N_18894);
or U19376 (N_19376,N_18628,N_18853);
or U19377 (N_19377,N_18734,N_19089);
and U19378 (N_19378,N_19092,N_18756);
or U19379 (N_19379,N_19148,N_18779);
nor U19380 (N_19380,N_19063,N_18880);
and U19381 (N_19381,N_18959,N_18865);
nor U19382 (N_19382,N_18854,N_18858);
nor U19383 (N_19383,N_19179,N_18776);
or U19384 (N_19384,N_19141,N_18923);
or U19385 (N_19385,N_18664,N_18741);
xnor U19386 (N_19386,N_18603,N_18732);
or U19387 (N_19387,N_18883,N_18978);
and U19388 (N_19388,N_19167,N_19104);
or U19389 (N_19389,N_18970,N_19170);
and U19390 (N_19390,N_18850,N_18814);
and U19391 (N_19391,N_18852,N_18675);
or U19392 (N_19392,N_18807,N_18804);
nand U19393 (N_19393,N_18827,N_19151);
nand U19394 (N_19394,N_19090,N_19138);
nor U19395 (N_19395,N_19114,N_19056);
and U19396 (N_19396,N_18733,N_18650);
and U19397 (N_19397,N_19010,N_19140);
nor U19398 (N_19398,N_18602,N_18871);
nor U19399 (N_19399,N_19000,N_18604);
and U19400 (N_19400,N_18908,N_18885);
nor U19401 (N_19401,N_18899,N_19137);
nor U19402 (N_19402,N_18754,N_18896);
and U19403 (N_19403,N_19057,N_19168);
nand U19404 (N_19404,N_18760,N_18795);
nand U19405 (N_19405,N_18820,N_18918);
nand U19406 (N_19406,N_18631,N_19154);
and U19407 (N_19407,N_18771,N_18777);
nor U19408 (N_19408,N_18778,N_19119);
nand U19409 (N_19409,N_18787,N_19094);
nor U19410 (N_19410,N_18843,N_19156);
or U19411 (N_19411,N_19066,N_18984);
nor U19412 (N_19412,N_18891,N_18752);
nor U19413 (N_19413,N_18757,N_18736);
nand U19414 (N_19414,N_18919,N_18669);
or U19415 (N_19415,N_18615,N_19084);
or U19416 (N_19416,N_19172,N_18730);
or U19417 (N_19417,N_18792,N_18697);
and U19418 (N_19418,N_18805,N_19027);
and U19419 (N_19419,N_19129,N_18685);
or U19420 (N_19420,N_19164,N_18972);
and U19421 (N_19421,N_19032,N_19113);
nor U19422 (N_19422,N_19085,N_18837);
and U19423 (N_19423,N_18698,N_19123);
and U19424 (N_19424,N_18874,N_19016);
or U19425 (N_19425,N_18684,N_18716);
and U19426 (N_19426,N_18782,N_18765);
and U19427 (N_19427,N_18873,N_18816);
nor U19428 (N_19428,N_19060,N_18862);
nor U19429 (N_19429,N_18705,N_19102);
or U19430 (N_19430,N_18709,N_18738);
or U19431 (N_19431,N_18892,N_19034);
nor U19432 (N_19432,N_18636,N_18995);
nand U19433 (N_19433,N_19091,N_19134);
nand U19434 (N_19434,N_18831,N_18713);
nand U19435 (N_19435,N_18980,N_19162);
and U19436 (N_19436,N_18671,N_19002);
nand U19437 (N_19437,N_18655,N_18755);
or U19438 (N_19438,N_19088,N_19196);
or U19439 (N_19439,N_18938,N_19146);
xnor U19440 (N_19440,N_18687,N_19038);
nor U19441 (N_19441,N_19158,N_19008);
nand U19442 (N_19442,N_18745,N_18620);
nand U19443 (N_19443,N_18818,N_18654);
nor U19444 (N_19444,N_19115,N_18916);
nand U19445 (N_19445,N_18976,N_19029);
nand U19446 (N_19446,N_18751,N_19050);
and U19447 (N_19447,N_19047,N_19053);
nand U19448 (N_19448,N_18665,N_18612);
nor U19449 (N_19449,N_18889,N_18806);
or U19450 (N_19450,N_19061,N_18621);
and U19451 (N_19451,N_19116,N_18833);
nand U19452 (N_19452,N_19194,N_19081);
or U19453 (N_19453,N_18641,N_18748);
xnor U19454 (N_19454,N_18958,N_18682);
or U19455 (N_19455,N_18656,N_18912);
and U19456 (N_19456,N_18879,N_18817);
or U19457 (N_19457,N_19078,N_19096);
nand U19458 (N_19458,N_19044,N_18667);
or U19459 (N_19459,N_18828,N_18872);
or U19460 (N_19460,N_18683,N_18648);
nand U19461 (N_19461,N_19136,N_18839);
or U19462 (N_19462,N_18753,N_18840);
nor U19463 (N_19463,N_18895,N_18990);
nand U19464 (N_19464,N_19149,N_18761);
nor U19465 (N_19465,N_18893,N_18977);
and U19466 (N_19466,N_19086,N_18950);
xor U19467 (N_19467,N_19051,N_18712);
xnor U19468 (N_19468,N_18601,N_18626);
nor U19469 (N_19469,N_18600,N_18838);
or U19470 (N_19470,N_18996,N_19054);
nor U19471 (N_19471,N_19120,N_18987);
nand U19472 (N_19472,N_18974,N_18674);
xor U19473 (N_19473,N_19126,N_19188);
or U19474 (N_19474,N_18878,N_19079);
or U19475 (N_19475,N_18939,N_19045);
or U19476 (N_19476,N_19175,N_19007);
or U19477 (N_19477,N_18944,N_18742);
or U19478 (N_19478,N_19073,N_19087);
nand U19479 (N_19479,N_19095,N_19098);
or U19480 (N_19480,N_18640,N_19021);
and U19481 (N_19481,N_18627,N_18808);
nor U19482 (N_19482,N_19192,N_18869);
nand U19483 (N_19483,N_19017,N_18954);
and U19484 (N_19484,N_19105,N_19006);
nand U19485 (N_19485,N_18662,N_18920);
nor U19486 (N_19486,N_18845,N_18613);
nand U19487 (N_19487,N_19153,N_19037);
nand U19488 (N_19488,N_18749,N_18932);
nand U19489 (N_19489,N_19143,N_18694);
nor U19490 (N_19490,N_18714,N_18649);
and U19491 (N_19491,N_18951,N_18931);
nor U19492 (N_19492,N_18994,N_19176);
nand U19493 (N_19493,N_18803,N_18907);
or U19494 (N_19494,N_18645,N_18952);
or U19495 (N_19495,N_18784,N_18701);
and U19496 (N_19496,N_18911,N_19065);
nor U19497 (N_19497,N_18823,N_18646);
or U19498 (N_19498,N_19165,N_19145);
nor U19499 (N_19499,N_18882,N_19133);
and U19500 (N_19500,N_18957,N_18956);
or U19501 (N_19501,N_18628,N_18992);
or U19502 (N_19502,N_19044,N_18883);
and U19503 (N_19503,N_18919,N_18832);
and U19504 (N_19504,N_18829,N_18705);
xor U19505 (N_19505,N_19026,N_18805);
nand U19506 (N_19506,N_19032,N_19040);
nand U19507 (N_19507,N_18862,N_18719);
or U19508 (N_19508,N_18687,N_18672);
xor U19509 (N_19509,N_19166,N_18717);
or U19510 (N_19510,N_18931,N_18809);
or U19511 (N_19511,N_18672,N_18735);
or U19512 (N_19512,N_19095,N_18634);
nor U19513 (N_19513,N_18817,N_18699);
and U19514 (N_19514,N_19032,N_18758);
and U19515 (N_19515,N_18975,N_19153);
nor U19516 (N_19516,N_19031,N_18643);
nor U19517 (N_19517,N_18751,N_18828);
nand U19518 (N_19518,N_18620,N_18858);
or U19519 (N_19519,N_18707,N_19143);
nor U19520 (N_19520,N_18656,N_18966);
nor U19521 (N_19521,N_19070,N_18823);
or U19522 (N_19522,N_18655,N_18979);
and U19523 (N_19523,N_18855,N_18813);
nand U19524 (N_19524,N_18839,N_19064);
or U19525 (N_19525,N_18879,N_19037);
nor U19526 (N_19526,N_18771,N_18822);
nor U19527 (N_19527,N_19061,N_19068);
nor U19528 (N_19528,N_19170,N_18941);
and U19529 (N_19529,N_19187,N_18693);
nor U19530 (N_19530,N_18987,N_18798);
nor U19531 (N_19531,N_19009,N_18998);
nor U19532 (N_19532,N_19176,N_19120);
or U19533 (N_19533,N_18751,N_18718);
or U19534 (N_19534,N_18795,N_19146);
or U19535 (N_19535,N_19039,N_18730);
nor U19536 (N_19536,N_18784,N_18957);
nand U19537 (N_19537,N_18915,N_19020);
or U19538 (N_19538,N_19008,N_18826);
and U19539 (N_19539,N_18663,N_19019);
nor U19540 (N_19540,N_18937,N_18968);
or U19541 (N_19541,N_18759,N_19163);
nor U19542 (N_19542,N_18917,N_18971);
nand U19543 (N_19543,N_18697,N_19068);
nor U19544 (N_19544,N_18871,N_19031);
nor U19545 (N_19545,N_18742,N_18615);
nor U19546 (N_19546,N_19056,N_19185);
or U19547 (N_19547,N_19109,N_19024);
or U19548 (N_19548,N_19171,N_18908);
nor U19549 (N_19549,N_19125,N_18708);
nand U19550 (N_19550,N_18839,N_18882);
nand U19551 (N_19551,N_19130,N_19016);
and U19552 (N_19552,N_18686,N_19086);
or U19553 (N_19553,N_18876,N_18602);
nor U19554 (N_19554,N_18989,N_19009);
and U19555 (N_19555,N_18739,N_18820);
and U19556 (N_19556,N_18964,N_18896);
or U19557 (N_19557,N_18626,N_19184);
nor U19558 (N_19558,N_18830,N_19170);
and U19559 (N_19559,N_18610,N_18684);
and U19560 (N_19560,N_18965,N_18670);
and U19561 (N_19561,N_19014,N_19075);
or U19562 (N_19562,N_18905,N_18683);
and U19563 (N_19563,N_19059,N_18907);
or U19564 (N_19564,N_19062,N_18654);
and U19565 (N_19565,N_18873,N_18658);
nor U19566 (N_19566,N_18878,N_19014);
and U19567 (N_19567,N_18739,N_19065);
or U19568 (N_19568,N_18756,N_18686);
and U19569 (N_19569,N_18781,N_18769);
or U19570 (N_19570,N_19180,N_18932);
or U19571 (N_19571,N_18889,N_19102);
nand U19572 (N_19572,N_19199,N_18621);
nand U19573 (N_19573,N_18889,N_18701);
nand U19574 (N_19574,N_18658,N_18902);
nor U19575 (N_19575,N_19091,N_18709);
nor U19576 (N_19576,N_19132,N_18915);
nand U19577 (N_19577,N_19069,N_19117);
nand U19578 (N_19578,N_18906,N_19083);
nand U19579 (N_19579,N_19004,N_18699);
nand U19580 (N_19580,N_19191,N_18766);
nand U19581 (N_19581,N_18769,N_19090);
or U19582 (N_19582,N_19099,N_19039);
and U19583 (N_19583,N_19151,N_18783);
or U19584 (N_19584,N_18707,N_19128);
or U19585 (N_19585,N_18660,N_18607);
nand U19586 (N_19586,N_18647,N_19105);
or U19587 (N_19587,N_18895,N_18733);
nor U19588 (N_19588,N_18647,N_18970);
nand U19589 (N_19589,N_19114,N_19168);
nor U19590 (N_19590,N_18760,N_18891);
nor U19591 (N_19591,N_19032,N_19021);
and U19592 (N_19592,N_18856,N_18703);
and U19593 (N_19593,N_19019,N_18816);
and U19594 (N_19594,N_18932,N_18936);
or U19595 (N_19595,N_18856,N_19018);
nand U19596 (N_19596,N_19060,N_18611);
nor U19597 (N_19597,N_18996,N_18839);
and U19598 (N_19598,N_18621,N_18970);
and U19599 (N_19599,N_18976,N_19077);
and U19600 (N_19600,N_19056,N_18722);
or U19601 (N_19601,N_19028,N_18938);
or U19602 (N_19602,N_18654,N_18864);
nand U19603 (N_19603,N_19014,N_19143);
nand U19604 (N_19604,N_19149,N_19055);
and U19605 (N_19605,N_19170,N_19190);
or U19606 (N_19606,N_19065,N_18609);
nand U19607 (N_19607,N_19053,N_19114);
nor U19608 (N_19608,N_18688,N_18808);
nand U19609 (N_19609,N_19111,N_19046);
nand U19610 (N_19610,N_18805,N_19179);
nand U19611 (N_19611,N_19124,N_18917);
or U19612 (N_19612,N_18845,N_18827);
nand U19613 (N_19613,N_19079,N_19012);
or U19614 (N_19614,N_19106,N_18646);
and U19615 (N_19615,N_19043,N_18877);
nor U19616 (N_19616,N_18602,N_19109);
nor U19617 (N_19617,N_18712,N_18897);
or U19618 (N_19618,N_18618,N_18934);
nor U19619 (N_19619,N_19121,N_18813);
nand U19620 (N_19620,N_18810,N_19100);
and U19621 (N_19621,N_18968,N_18913);
or U19622 (N_19622,N_18831,N_18907);
nand U19623 (N_19623,N_19095,N_18720);
nor U19624 (N_19624,N_18930,N_18721);
and U19625 (N_19625,N_18697,N_18721);
nand U19626 (N_19626,N_19174,N_19008);
or U19627 (N_19627,N_18837,N_18736);
or U19628 (N_19628,N_19008,N_18831);
and U19629 (N_19629,N_18997,N_18907);
xor U19630 (N_19630,N_18742,N_18733);
nor U19631 (N_19631,N_18640,N_18626);
and U19632 (N_19632,N_19139,N_18619);
xnor U19633 (N_19633,N_18905,N_18978);
nor U19634 (N_19634,N_18622,N_19089);
nor U19635 (N_19635,N_19082,N_18928);
xor U19636 (N_19636,N_18950,N_18845);
and U19637 (N_19637,N_19036,N_18844);
nor U19638 (N_19638,N_18905,N_18723);
and U19639 (N_19639,N_18789,N_18949);
or U19640 (N_19640,N_19093,N_19124);
or U19641 (N_19641,N_18662,N_18901);
and U19642 (N_19642,N_18785,N_18708);
and U19643 (N_19643,N_19074,N_18632);
or U19644 (N_19644,N_18876,N_18858);
nand U19645 (N_19645,N_19087,N_18672);
or U19646 (N_19646,N_19001,N_19132);
or U19647 (N_19647,N_19112,N_18963);
or U19648 (N_19648,N_18618,N_18979);
nand U19649 (N_19649,N_19092,N_19123);
nor U19650 (N_19650,N_19113,N_18893);
nand U19651 (N_19651,N_18943,N_19112);
or U19652 (N_19652,N_19013,N_19003);
and U19653 (N_19653,N_18627,N_18892);
nand U19654 (N_19654,N_18756,N_18653);
and U19655 (N_19655,N_19070,N_19104);
or U19656 (N_19656,N_18900,N_18757);
and U19657 (N_19657,N_18833,N_18788);
and U19658 (N_19658,N_18792,N_18839);
and U19659 (N_19659,N_19081,N_18787);
nor U19660 (N_19660,N_18795,N_18746);
and U19661 (N_19661,N_18614,N_18995);
or U19662 (N_19662,N_18993,N_19151);
nor U19663 (N_19663,N_18822,N_19097);
nand U19664 (N_19664,N_18817,N_18940);
nor U19665 (N_19665,N_18870,N_18970);
nor U19666 (N_19666,N_18858,N_18628);
and U19667 (N_19667,N_19017,N_18722);
nor U19668 (N_19668,N_19006,N_19080);
nor U19669 (N_19669,N_18882,N_19053);
or U19670 (N_19670,N_18678,N_18865);
nor U19671 (N_19671,N_18734,N_19168);
and U19672 (N_19672,N_19105,N_18622);
or U19673 (N_19673,N_18883,N_18952);
or U19674 (N_19674,N_18680,N_19071);
and U19675 (N_19675,N_18761,N_18949);
and U19676 (N_19676,N_18976,N_19119);
and U19677 (N_19677,N_18646,N_19075);
or U19678 (N_19678,N_18761,N_18810);
nand U19679 (N_19679,N_18682,N_19008);
and U19680 (N_19680,N_18881,N_18632);
or U19681 (N_19681,N_18853,N_18766);
or U19682 (N_19682,N_18811,N_18654);
or U19683 (N_19683,N_18678,N_19124);
nand U19684 (N_19684,N_18886,N_18613);
and U19685 (N_19685,N_18677,N_19041);
or U19686 (N_19686,N_19014,N_18903);
xnor U19687 (N_19687,N_18909,N_18643);
or U19688 (N_19688,N_19196,N_18919);
nand U19689 (N_19689,N_18826,N_18839);
or U19690 (N_19690,N_18986,N_18858);
nand U19691 (N_19691,N_19004,N_18934);
nand U19692 (N_19692,N_19109,N_18984);
or U19693 (N_19693,N_19180,N_18686);
or U19694 (N_19694,N_18774,N_19095);
or U19695 (N_19695,N_18695,N_18839);
or U19696 (N_19696,N_18670,N_19069);
or U19697 (N_19697,N_18726,N_18643);
nand U19698 (N_19698,N_19047,N_18767);
nor U19699 (N_19699,N_18651,N_19055);
nor U19700 (N_19700,N_18793,N_18914);
or U19701 (N_19701,N_18887,N_19091);
nand U19702 (N_19702,N_18851,N_18944);
and U19703 (N_19703,N_18609,N_18926);
xnor U19704 (N_19704,N_19128,N_19179);
nor U19705 (N_19705,N_18775,N_19177);
and U19706 (N_19706,N_19144,N_18994);
nor U19707 (N_19707,N_19071,N_18677);
nor U19708 (N_19708,N_19119,N_18720);
or U19709 (N_19709,N_18702,N_18733);
nor U19710 (N_19710,N_19063,N_18799);
nand U19711 (N_19711,N_19000,N_18929);
and U19712 (N_19712,N_18985,N_18695);
nand U19713 (N_19713,N_19131,N_19199);
nor U19714 (N_19714,N_18924,N_18858);
and U19715 (N_19715,N_18651,N_18807);
or U19716 (N_19716,N_18771,N_18617);
or U19717 (N_19717,N_18686,N_19054);
and U19718 (N_19718,N_18687,N_18936);
nand U19719 (N_19719,N_19090,N_18823);
or U19720 (N_19720,N_18991,N_18814);
or U19721 (N_19721,N_19072,N_19106);
nor U19722 (N_19722,N_18948,N_18807);
nor U19723 (N_19723,N_18607,N_18847);
nand U19724 (N_19724,N_18881,N_18640);
and U19725 (N_19725,N_18960,N_19167);
nor U19726 (N_19726,N_18666,N_19124);
nand U19727 (N_19727,N_18887,N_18904);
and U19728 (N_19728,N_18877,N_19144);
or U19729 (N_19729,N_18967,N_18847);
and U19730 (N_19730,N_18830,N_18810);
nor U19731 (N_19731,N_18849,N_18768);
nor U19732 (N_19732,N_18616,N_18867);
nand U19733 (N_19733,N_18977,N_18887);
nand U19734 (N_19734,N_19138,N_19084);
and U19735 (N_19735,N_19109,N_19087);
and U19736 (N_19736,N_19031,N_19174);
and U19737 (N_19737,N_19169,N_18843);
nand U19738 (N_19738,N_19010,N_18894);
or U19739 (N_19739,N_19195,N_18867);
or U19740 (N_19740,N_19050,N_19143);
nand U19741 (N_19741,N_19090,N_19182);
and U19742 (N_19742,N_18645,N_18759);
and U19743 (N_19743,N_18702,N_19080);
nor U19744 (N_19744,N_19048,N_19065);
and U19745 (N_19745,N_18619,N_18807);
nand U19746 (N_19746,N_18987,N_18976);
or U19747 (N_19747,N_19189,N_18890);
nor U19748 (N_19748,N_19185,N_19158);
nor U19749 (N_19749,N_19047,N_18758);
nand U19750 (N_19750,N_19199,N_19115);
nand U19751 (N_19751,N_19186,N_19155);
or U19752 (N_19752,N_18952,N_18691);
or U19753 (N_19753,N_19095,N_19086);
or U19754 (N_19754,N_18646,N_18609);
nand U19755 (N_19755,N_18888,N_18872);
and U19756 (N_19756,N_18759,N_19126);
nand U19757 (N_19757,N_18949,N_18757);
and U19758 (N_19758,N_18738,N_18708);
and U19759 (N_19759,N_18606,N_18730);
or U19760 (N_19760,N_18654,N_18646);
nor U19761 (N_19761,N_18922,N_18652);
nand U19762 (N_19762,N_19058,N_19128);
nand U19763 (N_19763,N_18911,N_19197);
xnor U19764 (N_19764,N_19086,N_18645);
or U19765 (N_19765,N_18908,N_18626);
and U19766 (N_19766,N_18865,N_18669);
nand U19767 (N_19767,N_19097,N_18844);
nand U19768 (N_19768,N_18838,N_19183);
nand U19769 (N_19769,N_19029,N_18682);
xnor U19770 (N_19770,N_18783,N_18813);
nor U19771 (N_19771,N_19024,N_18695);
nand U19772 (N_19772,N_18720,N_18620);
nand U19773 (N_19773,N_18660,N_19022);
or U19774 (N_19774,N_19109,N_18787);
and U19775 (N_19775,N_19155,N_18910);
nand U19776 (N_19776,N_18828,N_18684);
or U19777 (N_19777,N_18682,N_18925);
or U19778 (N_19778,N_19138,N_18841);
nor U19779 (N_19779,N_18728,N_19164);
xnor U19780 (N_19780,N_18791,N_19040);
xor U19781 (N_19781,N_18940,N_18791);
and U19782 (N_19782,N_18611,N_19142);
nand U19783 (N_19783,N_18983,N_18891);
nand U19784 (N_19784,N_18841,N_18996);
nand U19785 (N_19785,N_18704,N_18830);
nor U19786 (N_19786,N_19124,N_18749);
nor U19787 (N_19787,N_18853,N_18911);
and U19788 (N_19788,N_19035,N_18692);
xor U19789 (N_19789,N_18776,N_18864);
and U19790 (N_19790,N_19076,N_18822);
and U19791 (N_19791,N_19192,N_19066);
and U19792 (N_19792,N_19096,N_18600);
nand U19793 (N_19793,N_18731,N_18846);
and U19794 (N_19794,N_19156,N_18811);
xor U19795 (N_19795,N_19000,N_19098);
or U19796 (N_19796,N_19088,N_19146);
nor U19797 (N_19797,N_18881,N_18899);
or U19798 (N_19798,N_18889,N_18916);
nand U19799 (N_19799,N_18785,N_18756);
and U19800 (N_19800,N_19289,N_19722);
nor U19801 (N_19801,N_19261,N_19573);
nand U19802 (N_19802,N_19756,N_19449);
and U19803 (N_19803,N_19501,N_19411);
and U19804 (N_19804,N_19584,N_19668);
nand U19805 (N_19805,N_19201,N_19500);
nand U19806 (N_19806,N_19364,N_19224);
and U19807 (N_19807,N_19544,N_19207);
nor U19808 (N_19808,N_19484,N_19563);
and U19809 (N_19809,N_19533,N_19318);
or U19810 (N_19810,N_19695,N_19431);
xnor U19811 (N_19811,N_19259,N_19476);
and U19812 (N_19812,N_19412,N_19527);
nand U19813 (N_19813,N_19684,N_19331);
xnor U19814 (N_19814,N_19534,N_19227);
nand U19815 (N_19815,N_19418,N_19294);
nor U19816 (N_19816,N_19304,N_19220);
and U19817 (N_19817,N_19792,N_19234);
nor U19818 (N_19818,N_19767,N_19350);
and U19819 (N_19819,N_19583,N_19319);
nand U19820 (N_19820,N_19376,N_19219);
nand U19821 (N_19821,N_19675,N_19473);
nand U19822 (N_19822,N_19607,N_19326);
and U19823 (N_19823,N_19754,N_19265);
and U19824 (N_19824,N_19337,N_19508);
nand U19825 (N_19825,N_19783,N_19249);
or U19826 (N_19826,N_19665,N_19549);
and U19827 (N_19827,N_19378,N_19755);
or U19828 (N_19828,N_19644,N_19585);
nand U19829 (N_19829,N_19316,N_19540);
nand U19830 (N_19830,N_19594,N_19794);
or U19831 (N_19831,N_19639,N_19360);
or U19832 (N_19832,N_19687,N_19642);
nor U19833 (N_19833,N_19263,N_19238);
nand U19834 (N_19834,N_19321,N_19662);
and U19835 (N_19835,N_19497,N_19398);
nor U19836 (N_19836,N_19513,N_19221);
or U19837 (N_19837,N_19509,N_19303);
xnor U19838 (N_19838,N_19773,N_19752);
nand U19839 (N_19839,N_19424,N_19499);
or U19840 (N_19840,N_19517,N_19613);
and U19841 (N_19841,N_19658,N_19299);
nand U19842 (N_19842,N_19264,N_19298);
or U19843 (N_19843,N_19590,N_19787);
and U19844 (N_19844,N_19737,N_19377);
nor U19845 (N_19845,N_19515,N_19223);
nor U19846 (N_19846,N_19570,N_19554);
nor U19847 (N_19847,N_19553,N_19243);
and U19848 (N_19848,N_19325,N_19560);
nor U19849 (N_19849,N_19339,N_19771);
or U19850 (N_19850,N_19362,N_19680);
nand U19851 (N_19851,N_19649,N_19693);
nand U19852 (N_19852,N_19237,N_19539);
nor U19853 (N_19853,N_19248,N_19366);
and U19854 (N_19854,N_19620,N_19548);
or U19855 (N_19855,N_19525,N_19724);
nor U19856 (N_19856,N_19797,N_19694);
xor U19857 (N_19857,N_19487,N_19222);
and U19858 (N_19858,N_19233,N_19429);
nand U19859 (N_19859,N_19335,N_19381);
or U19860 (N_19860,N_19716,N_19660);
and U19861 (N_19861,N_19516,N_19683);
and U19862 (N_19862,N_19511,N_19438);
and U19863 (N_19863,N_19469,N_19205);
nand U19864 (N_19864,N_19543,N_19251);
nor U19865 (N_19865,N_19556,N_19498);
nor U19866 (N_19866,N_19715,N_19640);
or U19867 (N_19867,N_19312,N_19464);
nand U19868 (N_19868,N_19349,N_19460);
nand U19869 (N_19869,N_19228,N_19440);
and U19870 (N_19870,N_19267,N_19605);
or U19871 (N_19871,N_19442,N_19632);
nand U19872 (N_19872,N_19647,N_19652);
nand U19873 (N_19873,N_19707,N_19531);
and U19874 (N_19874,N_19271,N_19296);
or U19875 (N_19875,N_19396,N_19608);
or U19876 (N_19876,N_19455,N_19575);
nor U19877 (N_19877,N_19677,N_19285);
nand U19878 (N_19878,N_19609,N_19699);
nand U19879 (N_19879,N_19612,N_19358);
xor U19880 (N_19880,N_19468,N_19778);
nor U19881 (N_19881,N_19764,N_19242);
and U19882 (N_19882,N_19505,N_19306);
and U19883 (N_19883,N_19439,N_19519);
and U19884 (N_19884,N_19718,N_19555);
nor U19885 (N_19885,N_19232,N_19399);
and U19886 (N_19886,N_19686,N_19307);
xor U19887 (N_19887,N_19580,N_19616);
and U19888 (N_19888,N_19689,N_19314);
nor U19889 (N_19889,N_19777,N_19581);
nand U19890 (N_19890,N_19546,N_19388);
or U19891 (N_19891,N_19256,N_19655);
xor U19892 (N_19892,N_19338,N_19493);
nor U19893 (N_19893,N_19372,N_19557);
nor U19894 (N_19894,N_19212,N_19365);
nor U19895 (N_19895,N_19610,N_19636);
nor U19896 (N_19896,N_19714,N_19203);
nor U19897 (N_19897,N_19214,N_19788);
or U19898 (N_19898,N_19759,N_19322);
nand U19899 (N_19899,N_19281,N_19384);
or U19900 (N_19900,N_19369,N_19762);
nand U19901 (N_19901,N_19280,N_19309);
and U19902 (N_19902,N_19209,N_19416);
nand U19903 (N_19903,N_19713,N_19290);
nor U19904 (N_19904,N_19295,N_19648);
nor U19905 (N_19905,N_19269,N_19542);
or U19906 (N_19906,N_19451,N_19629);
or U19907 (N_19907,N_19611,N_19391);
nor U19908 (N_19908,N_19731,N_19749);
or U19909 (N_19909,N_19472,N_19262);
or U19910 (N_19910,N_19617,N_19300);
and U19911 (N_19911,N_19336,N_19245);
nand U19912 (N_19912,N_19567,N_19743);
nand U19913 (N_19913,N_19547,N_19490);
nor U19914 (N_19914,N_19667,N_19415);
nand U19915 (N_19915,N_19389,N_19456);
and U19916 (N_19916,N_19623,N_19387);
or U19917 (N_19917,N_19385,N_19635);
or U19918 (N_19918,N_19491,N_19332);
and U19919 (N_19919,N_19448,N_19382);
and U19920 (N_19920,N_19286,N_19650);
nand U19921 (N_19921,N_19458,N_19638);
and U19922 (N_19922,N_19481,N_19796);
or U19923 (N_19923,N_19340,N_19457);
nor U19924 (N_19924,N_19272,N_19466);
and U19925 (N_19925,N_19241,N_19780);
nor U19926 (N_19926,N_19690,N_19681);
and U19927 (N_19927,N_19673,N_19239);
and U19928 (N_19928,N_19253,N_19346);
nor U19929 (N_19929,N_19218,N_19293);
nor U19930 (N_19930,N_19748,N_19732);
or U19931 (N_19931,N_19663,N_19661);
nor U19932 (N_19932,N_19216,N_19370);
or U19933 (N_19933,N_19202,N_19363);
or U19934 (N_19934,N_19521,N_19786);
nand U19935 (N_19935,N_19447,N_19402);
nor U19936 (N_19936,N_19266,N_19761);
and U19937 (N_19937,N_19664,N_19735);
or U19938 (N_19938,N_19592,N_19624);
nor U19939 (N_19939,N_19344,N_19204);
nor U19940 (N_19940,N_19669,N_19551);
nand U19941 (N_19941,N_19628,N_19368);
nor U19942 (N_19942,N_19710,N_19333);
and U19943 (N_19943,N_19784,N_19518);
nand U19944 (N_19944,N_19357,N_19618);
nor U19945 (N_19945,N_19751,N_19329);
or U19946 (N_19946,N_19702,N_19302);
or U19947 (N_19947,N_19225,N_19785);
nand U19948 (N_19948,N_19565,N_19659);
or U19949 (N_19949,N_19602,N_19646);
and U19950 (N_19950,N_19297,N_19507);
and U19951 (N_19951,N_19591,N_19676);
nor U19952 (N_19952,N_19414,N_19211);
and U19953 (N_19953,N_19409,N_19478);
and U19954 (N_19954,N_19729,N_19723);
nor U19955 (N_19955,N_19558,N_19528);
nor U19956 (N_19956,N_19781,N_19705);
nor U19957 (N_19957,N_19657,N_19696);
and U19958 (N_19958,N_19494,N_19282);
and U19959 (N_19959,N_19571,N_19395);
or U19960 (N_19960,N_19206,N_19593);
nor U19961 (N_19961,N_19257,N_19356);
or U19962 (N_19962,N_19443,N_19471);
and U19963 (N_19963,N_19461,N_19479);
or U19964 (N_19964,N_19404,N_19597);
nor U19965 (N_19965,N_19670,N_19229);
or U19966 (N_19966,N_19305,N_19782);
and U19967 (N_19967,N_19361,N_19480);
or U19968 (N_19968,N_19450,N_19217);
or U19969 (N_19969,N_19578,N_19279);
nor U19970 (N_19970,N_19627,N_19445);
or U19971 (N_19971,N_19273,N_19758);
nor U19972 (N_19972,N_19483,N_19727);
xnor U19973 (N_19973,N_19600,N_19656);
nand U19974 (N_19974,N_19400,N_19526);
or U19975 (N_19975,N_19524,N_19621);
or U19976 (N_19976,N_19236,N_19572);
nand U19977 (N_19977,N_19379,N_19576);
or U19978 (N_19978,N_19579,N_19599);
or U19979 (N_19979,N_19341,N_19353);
nor U19980 (N_19980,N_19765,N_19700);
nor U19981 (N_19981,N_19252,N_19308);
and U19982 (N_19982,N_19348,N_19691);
and U19983 (N_19983,N_19441,N_19453);
and U19984 (N_19984,N_19733,N_19422);
and U19985 (N_19985,N_19313,N_19405);
nor U19986 (N_19986,N_19492,N_19408);
nand U19987 (N_19987,N_19512,N_19383);
and U19988 (N_19988,N_19529,N_19601);
nor U19989 (N_19989,N_19488,N_19742);
or U19990 (N_19990,N_19744,N_19446);
xnor U19991 (N_19991,N_19327,N_19347);
or U19992 (N_19992,N_19489,N_19246);
nand U19993 (N_19993,N_19775,N_19247);
xor U19994 (N_19994,N_19776,N_19631);
and U19995 (N_19995,N_19688,N_19351);
and U19996 (N_19996,N_19393,N_19432);
nand U19997 (N_19997,N_19495,N_19770);
nand U19998 (N_19998,N_19698,N_19403);
or U19999 (N_19999,N_19274,N_19626);
or U20000 (N_20000,N_19793,N_19437);
and U20001 (N_20001,N_19725,N_19779);
nor U20002 (N_20002,N_19359,N_19730);
nand U20003 (N_20003,N_19287,N_19763);
nand U20004 (N_20004,N_19425,N_19428);
or U20005 (N_20005,N_19200,N_19426);
or U20006 (N_20006,N_19514,N_19284);
and U20007 (N_20007,N_19772,N_19709);
and U20008 (N_20008,N_19355,N_19401);
nor U20009 (N_20009,N_19739,N_19231);
nor U20010 (N_20010,N_19774,N_19712);
or U20011 (N_20011,N_19587,N_19750);
or U20012 (N_20012,N_19255,N_19208);
nand U20013 (N_20013,N_19697,N_19604);
and U20014 (N_20014,N_19380,N_19790);
or U20015 (N_20015,N_19603,N_19561);
and U20016 (N_20016,N_19760,N_19423);
and U20017 (N_20017,N_19462,N_19334);
nor U20018 (N_20018,N_19522,N_19477);
and U20019 (N_20019,N_19520,N_19719);
nand U20020 (N_20020,N_19747,N_19538);
nand U20021 (N_20021,N_19268,N_19354);
and U20022 (N_20022,N_19666,N_19769);
or U20023 (N_20023,N_19430,N_19250);
nand U20024 (N_20024,N_19679,N_19586);
nand U20025 (N_20025,N_19503,N_19275);
and U20026 (N_20026,N_19226,N_19535);
or U20027 (N_20027,N_19277,N_19345);
and U20028 (N_20028,N_19736,N_19745);
nand U20029 (N_20029,N_19530,N_19685);
or U20030 (N_20030,N_19215,N_19435);
xor U20031 (N_20031,N_19766,N_19682);
and U20032 (N_20032,N_19276,N_19343);
nor U20033 (N_20033,N_19552,N_19454);
nand U20034 (N_20034,N_19213,N_19496);
nor U20035 (N_20035,N_19537,N_19562);
nor U20036 (N_20036,N_19598,N_19651);
xor U20037 (N_20037,N_19566,N_19753);
or U20038 (N_20038,N_19734,N_19260);
nor U20039 (N_20039,N_19394,N_19371);
nor U20040 (N_20040,N_19452,N_19474);
and U20041 (N_20041,N_19559,N_19320);
xnor U20042 (N_20042,N_19577,N_19475);
nand U20043 (N_20043,N_19704,N_19324);
nand U20044 (N_20044,N_19485,N_19392);
nand U20045 (N_20045,N_19757,N_19619);
and U20046 (N_20046,N_19502,N_19596);
nand U20047 (N_20047,N_19614,N_19568);
and U20048 (N_20048,N_19671,N_19653);
and U20049 (N_20049,N_19315,N_19692);
nand U20050 (N_20050,N_19564,N_19390);
and U20051 (N_20051,N_19291,N_19436);
nand U20052 (N_20052,N_19654,N_19630);
nor U20053 (N_20053,N_19482,N_19615);
nor U20054 (N_20054,N_19406,N_19791);
nor U20055 (N_20055,N_19463,N_19574);
nor U20056 (N_20056,N_19589,N_19467);
nor U20057 (N_20057,N_19768,N_19470);
or U20058 (N_20058,N_19292,N_19410);
and U20059 (N_20059,N_19740,N_19421);
nand U20060 (N_20060,N_19545,N_19323);
nand U20061 (N_20061,N_19798,N_19633);
or U20062 (N_20062,N_19459,N_19637);
or U20063 (N_20063,N_19342,N_19352);
nand U20064 (N_20064,N_19721,N_19717);
nor U20065 (N_20065,N_19510,N_19795);
nor U20066 (N_20066,N_19532,N_19678);
xnor U20067 (N_20067,N_19301,N_19328);
xor U20068 (N_20068,N_19258,N_19708);
nand U20069 (N_20069,N_19595,N_19444);
or U20070 (N_20070,N_19645,N_19210);
nor U20071 (N_20071,N_19278,N_19375);
or U20072 (N_20072,N_19311,N_19703);
and U20073 (N_20073,N_19569,N_19407);
nor U20074 (N_20074,N_19420,N_19799);
or U20075 (N_20075,N_19728,N_19506);
nor U20076 (N_20076,N_19606,N_19504);
or U20077 (N_20077,N_19720,N_19701);
and U20078 (N_20078,N_19367,N_19434);
and U20079 (N_20079,N_19741,N_19550);
and U20080 (N_20080,N_19625,N_19672);
nor U20081 (N_20081,N_19746,N_19283);
nor U20082 (N_20082,N_19588,N_19386);
or U20083 (N_20083,N_19541,N_19373);
nand U20084 (N_20084,N_19465,N_19536);
nor U20085 (N_20085,N_19330,N_19738);
and U20086 (N_20086,N_19417,N_19789);
or U20087 (N_20087,N_19419,N_19235);
nor U20088 (N_20088,N_19270,N_19706);
and U20089 (N_20089,N_19726,N_19240);
nand U20090 (N_20090,N_19433,N_19643);
nor U20091 (N_20091,N_19310,N_19230);
nor U20092 (N_20092,N_19486,N_19413);
or U20093 (N_20093,N_19674,N_19374);
xnor U20094 (N_20094,N_19397,N_19427);
and U20095 (N_20095,N_19244,N_19254);
or U20096 (N_20096,N_19634,N_19641);
nand U20097 (N_20097,N_19622,N_19582);
nor U20098 (N_20098,N_19288,N_19317);
and U20099 (N_20099,N_19711,N_19523);
nor U20100 (N_20100,N_19753,N_19793);
or U20101 (N_20101,N_19759,N_19251);
nand U20102 (N_20102,N_19790,N_19797);
and U20103 (N_20103,N_19320,N_19460);
and U20104 (N_20104,N_19589,N_19388);
or U20105 (N_20105,N_19310,N_19643);
and U20106 (N_20106,N_19221,N_19252);
and U20107 (N_20107,N_19696,N_19308);
nand U20108 (N_20108,N_19590,N_19705);
nor U20109 (N_20109,N_19407,N_19431);
and U20110 (N_20110,N_19591,N_19525);
nand U20111 (N_20111,N_19231,N_19766);
nand U20112 (N_20112,N_19732,N_19792);
nor U20113 (N_20113,N_19242,N_19308);
nand U20114 (N_20114,N_19419,N_19238);
nand U20115 (N_20115,N_19281,N_19799);
or U20116 (N_20116,N_19659,N_19717);
or U20117 (N_20117,N_19287,N_19564);
nand U20118 (N_20118,N_19769,N_19396);
and U20119 (N_20119,N_19299,N_19368);
and U20120 (N_20120,N_19737,N_19795);
nand U20121 (N_20121,N_19489,N_19650);
nor U20122 (N_20122,N_19635,N_19561);
nor U20123 (N_20123,N_19269,N_19672);
or U20124 (N_20124,N_19762,N_19436);
or U20125 (N_20125,N_19688,N_19726);
nand U20126 (N_20126,N_19513,N_19790);
and U20127 (N_20127,N_19217,N_19761);
nand U20128 (N_20128,N_19516,N_19233);
nand U20129 (N_20129,N_19422,N_19703);
and U20130 (N_20130,N_19693,N_19541);
and U20131 (N_20131,N_19215,N_19332);
and U20132 (N_20132,N_19747,N_19607);
nor U20133 (N_20133,N_19390,N_19299);
nand U20134 (N_20134,N_19551,N_19781);
or U20135 (N_20135,N_19241,N_19706);
or U20136 (N_20136,N_19373,N_19215);
nand U20137 (N_20137,N_19575,N_19646);
nand U20138 (N_20138,N_19258,N_19616);
xor U20139 (N_20139,N_19537,N_19782);
nand U20140 (N_20140,N_19347,N_19787);
nor U20141 (N_20141,N_19459,N_19475);
nand U20142 (N_20142,N_19258,N_19341);
nor U20143 (N_20143,N_19449,N_19696);
or U20144 (N_20144,N_19247,N_19332);
nand U20145 (N_20145,N_19311,N_19649);
nor U20146 (N_20146,N_19302,N_19781);
or U20147 (N_20147,N_19481,N_19731);
xnor U20148 (N_20148,N_19538,N_19594);
and U20149 (N_20149,N_19335,N_19334);
and U20150 (N_20150,N_19417,N_19257);
nand U20151 (N_20151,N_19498,N_19433);
and U20152 (N_20152,N_19284,N_19260);
nor U20153 (N_20153,N_19727,N_19796);
nor U20154 (N_20154,N_19670,N_19693);
nor U20155 (N_20155,N_19622,N_19785);
nor U20156 (N_20156,N_19492,N_19235);
nor U20157 (N_20157,N_19388,N_19590);
or U20158 (N_20158,N_19659,N_19722);
and U20159 (N_20159,N_19301,N_19377);
or U20160 (N_20160,N_19774,N_19289);
nor U20161 (N_20161,N_19565,N_19790);
and U20162 (N_20162,N_19770,N_19327);
nand U20163 (N_20163,N_19718,N_19358);
nor U20164 (N_20164,N_19546,N_19452);
and U20165 (N_20165,N_19495,N_19287);
or U20166 (N_20166,N_19309,N_19453);
nor U20167 (N_20167,N_19667,N_19663);
nand U20168 (N_20168,N_19489,N_19775);
nor U20169 (N_20169,N_19478,N_19481);
nand U20170 (N_20170,N_19262,N_19640);
or U20171 (N_20171,N_19213,N_19702);
and U20172 (N_20172,N_19341,N_19656);
and U20173 (N_20173,N_19528,N_19389);
nand U20174 (N_20174,N_19233,N_19261);
and U20175 (N_20175,N_19368,N_19708);
and U20176 (N_20176,N_19555,N_19594);
nor U20177 (N_20177,N_19429,N_19711);
or U20178 (N_20178,N_19396,N_19420);
nand U20179 (N_20179,N_19343,N_19790);
and U20180 (N_20180,N_19377,N_19696);
nand U20181 (N_20181,N_19366,N_19735);
nor U20182 (N_20182,N_19462,N_19386);
nor U20183 (N_20183,N_19400,N_19674);
nand U20184 (N_20184,N_19291,N_19239);
and U20185 (N_20185,N_19599,N_19687);
or U20186 (N_20186,N_19581,N_19744);
nand U20187 (N_20187,N_19207,N_19782);
and U20188 (N_20188,N_19315,N_19237);
or U20189 (N_20189,N_19699,N_19552);
nor U20190 (N_20190,N_19568,N_19248);
nand U20191 (N_20191,N_19714,N_19459);
or U20192 (N_20192,N_19508,N_19583);
or U20193 (N_20193,N_19245,N_19265);
nand U20194 (N_20194,N_19656,N_19751);
nand U20195 (N_20195,N_19316,N_19455);
and U20196 (N_20196,N_19623,N_19505);
nand U20197 (N_20197,N_19413,N_19366);
nand U20198 (N_20198,N_19258,N_19491);
nor U20199 (N_20199,N_19734,N_19490);
and U20200 (N_20200,N_19331,N_19757);
and U20201 (N_20201,N_19532,N_19609);
nand U20202 (N_20202,N_19602,N_19695);
or U20203 (N_20203,N_19758,N_19589);
nor U20204 (N_20204,N_19436,N_19543);
nor U20205 (N_20205,N_19202,N_19542);
xnor U20206 (N_20206,N_19740,N_19792);
and U20207 (N_20207,N_19579,N_19431);
nand U20208 (N_20208,N_19694,N_19698);
nand U20209 (N_20209,N_19229,N_19458);
or U20210 (N_20210,N_19521,N_19558);
nand U20211 (N_20211,N_19789,N_19792);
nand U20212 (N_20212,N_19325,N_19353);
nand U20213 (N_20213,N_19425,N_19696);
nor U20214 (N_20214,N_19219,N_19361);
nand U20215 (N_20215,N_19511,N_19213);
and U20216 (N_20216,N_19358,N_19759);
nand U20217 (N_20217,N_19552,N_19651);
nand U20218 (N_20218,N_19760,N_19770);
nor U20219 (N_20219,N_19595,N_19278);
or U20220 (N_20220,N_19728,N_19503);
nand U20221 (N_20221,N_19485,N_19734);
and U20222 (N_20222,N_19734,N_19423);
nand U20223 (N_20223,N_19224,N_19718);
or U20224 (N_20224,N_19441,N_19770);
nor U20225 (N_20225,N_19270,N_19794);
or U20226 (N_20226,N_19441,N_19274);
and U20227 (N_20227,N_19500,N_19415);
nand U20228 (N_20228,N_19363,N_19411);
nor U20229 (N_20229,N_19240,N_19217);
and U20230 (N_20230,N_19447,N_19438);
and U20231 (N_20231,N_19709,N_19368);
or U20232 (N_20232,N_19438,N_19339);
or U20233 (N_20233,N_19291,N_19797);
nor U20234 (N_20234,N_19754,N_19779);
and U20235 (N_20235,N_19656,N_19400);
and U20236 (N_20236,N_19697,N_19636);
xnor U20237 (N_20237,N_19356,N_19618);
or U20238 (N_20238,N_19566,N_19543);
nand U20239 (N_20239,N_19707,N_19527);
nand U20240 (N_20240,N_19502,N_19613);
nor U20241 (N_20241,N_19232,N_19410);
nor U20242 (N_20242,N_19201,N_19277);
nand U20243 (N_20243,N_19245,N_19325);
or U20244 (N_20244,N_19721,N_19305);
or U20245 (N_20245,N_19222,N_19713);
nand U20246 (N_20246,N_19634,N_19458);
and U20247 (N_20247,N_19491,N_19688);
nor U20248 (N_20248,N_19504,N_19316);
and U20249 (N_20249,N_19420,N_19492);
or U20250 (N_20250,N_19252,N_19430);
nand U20251 (N_20251,N_19420,N_19576);
nor U20252 (N_20252,N_19475,N_19219);
nor U20253 (N_20253,N_19450,N_19643);
and U20254 (N_20254,N_19275,N_19361);
and U20255 (N_20255,N_19557,N_19698);
nor U20256 (N_20256,N_19507,N_19263);
or U20257 (N_20257,N_19552,N_19368);
nand U20258 (N_20258,N_19574,N_19337);
or U20259 (N_20259,N_19702,N_19709);
or U20260 (N_20260,N_19717,N_19626);
nor U20261 (N_20261,N_19324,N_19264);
nor U20262 (N_20262,N_19520,N_19359);
and U20263 (N_20263,N_19529,N_19537);
and U20264 (N_20264,N_19677,N_19387);
nor U20265 (N_20265,N_19716,N_19511);
or U20266 (N_20266,N_19688,N_19720);
or U20267 (N_20267,N_19682,N_19611);
and U20268 (N_20268,N_19283,N_19286);
xor U20269 (N_20269,N_19730,N_19380);
nor U20270 (N_20270,N_19449,N_19440);
or U20271 (N_20271,N_19476,N_19222);
or U20272 (N_20272,N_19325,N_19209);
xor U20273 (N_20273,N_19756,N_19299);
nor U20274 (N_20274,N_19314,N_19257);
or U20275 (N_20275,N_19562,N_19393);
and U20276 (N_20276,N_19324,N_19399);
or U20277 (N_20277,N_19339,N_19454);
xor U20278 (N_20278,N_19740,N_19571);
nor U20279 (N_20279,N_19640,N_19327);
nor U20280 (N_20280,N_19493,N_19460);
and U20281 (N_20281,N_19729,N_19397);
or U20282 (N_20282,N_19736,N_19645);
nand U20283 (N_20283,N_19286,N_19210);
or U20284 (N_20284,N_19745,N_19289);
or U20285 (N_20285,N_19729,N_19403);
nor U20286 (N_20286,N_19342,N_19750);
or U20287 (N_20287,N_19356,N_19752);
nor U20288 (N_20288,N_19637,N_19300);
nand U20289 (N_20289,N_19552,N_19281);
nand U20290 (N_20290,N_19793,N_19496);
nor U20291 (N_20291,N_19514,N_19666);
nand U20292 (N_20292,N_19235,N_19521);
nor U20293 (N_20293,N_19348,N_19283);
nand U20294 (N_20294,N_19697,N_19724);
nand U20295 (N_20295,N_19361,N_19335);
xnor U20296 (N_20296,N_19490,N_19514);
or U20297 (N_20297,N_19411,N_19289);
nor U20298 (N_20298,N_19498,N_19524);
nor U20299 (N_20299,N_19577,N_19290);
or U20300 (N_20300,N_19745,N_19485);
or U20301 (N_20301,N_19542,N_19798);
or U20302 (N_20302,N_19442,N_19265);
and U20303 (N_20303,N_19665,N_19419);
nor U20304 (N_20304,N_19766,N_19600);
nor U20305 (N_20305,N_19375,N_19337);
nand U20306 (N_20306,N_19490,N_19652);
or U20307 (N_20307,N_19596,N_19250);
or U20308 (N_20308,N_19679,N_19730);
nand U20309 (N_20309,N_19584,N_19295);
nand U20310 (N_20310,N_19293,N_19397);
or U20311 (N_20311,N_19370,N_19411);
nor U20312 (N_20312,N_19641,N_19687);
and U20313 (N_20313,N_19239,N_19476);
nand U20314 (N_20314,N_19257,N_19659);
or U20315 (N_20315,N_19587,N_19545);
nor U20316 (N_20316,N_19228,N_19702);
or U20317 (N_20317,N_19224,N_19499);
xor U20318 (N_20318,N_19250,N_19499);
nor U20319 (N_20319,N_19207,N_19629);
nor U20320 (N_20320,N_19670,N_19796);
or U20321 (N_20321,N_19581,N_19272);
nand U20322 (N_20322,N_19578,N_19431);
nand U20323 (N_20323,N_19641,N_19386);
or U20324 (N_20324,N_19308,N_19214);
and U20325 (N_20325,N_19798,N_19525);
xnor U20326 (N_20326,N_19763,N_19390);
or U20327 (N_20327,N_19277,N_19466);
nand U20328 (N_20328,N_19547,N_19635);
or U20329 (N_20329,N_19544,N_19295);
nor U20330 (N_20330,N_19229,N_19570);
nor U20331 (N_20331,N_19207,N_19420);
and U20332 (N_20332,N_19717,N_19379);
nand U20333 (N_20333,N_19372,N_19615);
nand U20334 (N_20334,N_19519,N_19751);
nand U20335 (N_20335,N_19456,N_19423);
or U20336 (N_20336,N_19624,N_19370);
and U20337 (N_20337,N_19226,N_19249);
nor U20338 (N_20338,N_19608,N_19212);
nor U20339 (N_20339,N_19757,N_19412);
xnor U20340 (N_20340,N_19369,N_19302);
and U20341 (N_20341,N_19501,N_19482);
and U20342 (N_20342,N_19515,N_19378);
nand U20343 (N_20343,N_19322,N_19642);
nand U20344 (N_20344,N_19556,N_19224);
nand U20345 (N_20345,N_19574,N_19243);
or U20346 (N_20346,N_19768,N_19792);
or U20347 (N_20347,N_19583,N_19385);
and U20348 (N_20348,N_19436,N_19690);
and U20349 (N_20349,N_19722,N_19526);
nor U20350 (N_20350,N_19592,N_19600);
or U20351 (N_20351,N_19305,N_19338);
and U20352 (N_20352,N_19225,N_19610);
or U20353 (N_20353,N_19787,N_19657);
and U20354 (N_20354,N_19501,N_19713);
nor U20355 (N_20355,N_19260,N_19584);
and U20356 (N_20356,N_19564,N_19342);
or U20357 (N_20357,N_19497,N_19255);
or U20358 (N_20358,N_19210,N_19250);
and U20359 (N_20359,N_19502,N_19343);
nor U20360 (N_20360,N_19213,N_19322);
and U20361 (N_20361,N_19331,N_19701);
nand U20362 (N_20362,N_19447,N_19317);
xnor U20363 (N_20363,N_19672,N_19603);
and U20364 (N_20364,N_19417,N_19697);
or U20365 (N_20365,N_19367,N_19458);
nand U20366 (N_20366,N_19293,N_19717);
nand U20367 (N_20367,N_19624,N_19734);
and U20368 (N_20368,N_19634,N_19526);
or U20369 (N_20369,N_19658,N_19561);
or U20370 (N_20370,N_19581,N_19684);
nand U20371 (N_20371,N_19308,N_19744);
or U20372 (N_20372,N_19376,N_19636);
and U20373 (N_20373,N_19429,N_19473);
and U20374 (N_20374,N_19223,N_19268);
and U20375 (N_20375,N_19230,N_19634);
or U20376 (N_20376,N_19420,N_19529);
nand U20377 (N_20377,N_19581,N_19488);
or U20378 (N_20378,N_19718,N_19277);
nor U20379 (N_20379,N_19417,N_19566);
nor U20380 (N_20380,N_19516,N_19586);
nand U20381 (N_20381,N_19375,N_19419);
and U20382 (N_20382,N_19694,N_19370);
and U20383 (N_20383,N_19318,N_19556);
nor U20384 (N_20384,N_19635,N_19632);
or U20385 (N_20385,N_19698,N_19289);
or U20386 (N_20386,N_19327,N_19400);
and U20387 (N_20387,N_19303,N_19622);
nand U20388 (N_20388,N_19475,N_19277);
nor U20389 (N_20389,N_19503,N_19650);
or U20390 (N_20390,N_19739,N_19506);
nor U20391 (N_20391,N_19468,N_19620);
or U20392 (N_20392,N_19362,N_19498);
or U20393 (N_20393,N_19723,N_19559);
nor U20394 (N_20394,N_19223,N_19546);
or U20395 (N_20395,N_19746,N_19528);
nor U20396 (N_20396,N_19270,N_19729);
nor U20397 (N_20397,N_19458,N_19218);
nand U20398 (N_20398,N_19345,N_19638);
nor U20399 (N_20399,N_19397,N_19407);
nand U20400 (N_20400,N_19851,N_20340);
nand U20401 (N_20401,N_20316,N_20235);
nor U20402 (N_20402,N_20039,N_20212);
xnor U20403 (N_20403,N_20311,N_19945);
nor U20404 (N_20404,N_19988,N_20180);
nor U20405 (N_20405,N_19983,N_20252);
or U20406 (N_20406,N_20390,N_20102);
and U20407 (N_20407,N_20004,N_20392);
nand U20408 (N_20408,N_20128,N_20114);
or U20409 (N_20409,N_20055,N_20136);
nand U20410 (N_20410,N_20115,N_20154);
nand U20411 (N_20411,N_19866,N_20083);
and U20412 (N_20412,N_20260,N_20216);
nor U20413 (N_20413,N_20150,N_20188);
nand U20414 (N_20414,N_20146,N_19944);
nor U20415 (N_20415,N_19981,N_19970);
nand U20416 (N_20416,N_19976,N_20249);
nor U20417 (N_20417,N_19919,N_19957);
and U20418 (N_20418,N_19831,N_19872);
nand U20419 (N_20419,N_20112,N_20286);
nand U20420 (N_20420,N_20242,N_20138);
nand U20421 (N_20421,N_20284,N_19877);
nand U20422 (N_20422,N_19911,N_20091);
and U20423 (N_20423,N_20008,N_19826);
xnor U20424 (N_20424,N_19842,N_20043);
and U20425 (N_20425,N_20054,N_20086);
and U20426 (N_20426,N_19952,N_20258);
and U20427 (N_20427,N_20240,N_20289);
nand U20428 (N_20428,N_20191,N_19884);
nand U20429 (N_20429,N_20326,N_20171);
or U20430 (N_20430,N_20342,N_19832);
nand U20431 (N_20431,N_20245,N_20141);
or U20432 (N_20432,N_20085,N_19838);
nand U20433 (N_20433,N_20337,N_20384);
or U20434 (N_20434,N_20122,N_19951);
nor U20435 (N_20435,N_20359,N_19978);
nand U20436 (N_20436,N_20155,N_20302);
nor U20437 (N_20437,N_20101,N_20177);
nand U20438 (N_20438,N_20264,N_20388);
or U20439 (N_20439,N_20028,N_20121);
nand U20440 (N_20440,N_20126,N_19928);
nand U20441 (N_20441,N_20183,N_20058);
nand U20442 (N_20442,N_20360,N_20296);
or U20443 (N_20443,N_20084,N_20009);
or U20444 (N_20444,N_20005,N_20147);
nand U20445 (N_20445,N_20132,N_20109);
and U20446 (N_20446,N_19990,N_19930);
and U20447 (N_20447,N_20068,N_19926);
nor U20448 (N_20448,N_20149,N_20229);
nor U20449 (N_20449,N_20287,N_20019);
nand U20450 (N_20450,N_20387,N_20305);
nor U20451 (N_20451,N_20098,N_19847);
nor U20452 (N_20452,N_20354,N_20320);
nand U20453 (N_20453,N_20381,N_19873);
nor U20454 (N_20454,N_19963,N_20351);
nor U20455 (N_20455,N_19856,N_20133);
and U20456 (N_20456,N_20394,N_20124);
and U20457 (N_20457,N_20293,N_20162);
or U20458 (N_20458,N_20110,N_19876);
nor U20459 (N_20459,N_20194,N_20012);
and U20460 (N_20460,N_20193,N_20233);
or U20461 (N_20461,N_20324,N_20017);
nand U20462 (N_20462,N_20376,N_20172);
or U20463 (N_20463,N_20176,N_20108);
or U20464 (N_20464,N_20160,N_20315);
nand U20465 (N_20465,N_20181,N_20358);
nor U20466 (N_20466,N_20209,N_20199);
nor U20467 (N_20467,N_20041,N_20158);
nand U20468 (N_20468,N_19937,N_20203);
or U20469 (N_20469,N_19849,N_19871);
and U20470 (N_20470,N_20190,N_19992);
or U20471 (N_20471,N_20288,N_20369);
or U20472 (N_20472,N_20088,N_20100);
nor U20473 (N_20473,N_20333,N_20001);
or U20474 (N_20474,N_20299,N_20330);
nand U20475 (N_20475,N_20053,N_20192);
and U20476 (N_20476,N_20165,N_20319);
nand U20477 (N_20477,N_19829,N_20372);
and U20478 (N_20478,N_20161,N_20064);
and U20479 (N_20479,N_19996,N_19896);
nor U20480 (N_20480,N_20187,N_20391);
nand U20481 (N_20481,N_20185,N_20285);
nor U20482 (N_20482,N_19878,N_20234);
and U20483 (N_20483,N_19865,N_20297);
or U20484 (N_20484,N_20259,N_19935);
nand U20485 (N_20485,N_20395,N_20000);
and U20486 (N_20486,N_20228,N_19912);
nand U20487 (N_20487,N_19997,N_20021);
and U20488 (N_20488,N_20230,N_19823);
nor U20489 (N_20489,N_20134,N_20250);
or U20490 (N_20490,N_19800,N_19903);
nor U20491 (N_20491,N_19835,N_19984);
nor U20492 (N_20492,N_20167,N_20006);
nor U20493 (N_20493,N_19875,N_19994);
or U20494 (N_20494,N_20170,N_20220);
or U20495 (N_20495,N_19922,N_20398);
nor U20496 (N_20496,N_19867,N_20221);
or U20497 (N_20497,N_20257,N_20156);
nor U20498 (N_20498,N_19844,N_20075);
nor U20499 (N_20499,N_19809,N_20377);
and U20500 (N_20500,N_20061,N_19942);
nor U20501 (N_20501,N_20151,N_19815);
or U20502 (N_20502,N_20385,N_20350);
and U20503 (N_20503,N_19850,N_20349);
nand U20504 (N_20504,N_20238,N_20353);
or U20505 (N_20505,N_19939,N_20262);
or U20506 (N_20506,N_19870,N_20366);
or U20507 (N_20507,N_20003,N_19953);
xor U20508 (N_20508,N_20168,N_20018);
nor U20509 (N_20509,N_19991,N_20037);
nand U20510 (N_20510,N_19910,N_20062);
nor U20511 (N_20511,N_20087,N_20274);
or U20512 (N_20512,N_19892,N_19959);
nor U20513 (N_20513,N_20261,N_20033);
and U20514 (N_20514,N_20304,N_20137);
and U20515 (N_20515,N_20208,N_19813);
nor U20516 (N_20516,N_19916,N_20131);
nand U20517 (N_20517,N_20202,N_20135);
xnor U20518 (N_20518,N_19880,N_20211);
nand U20519 (N_20519,N_19936,N_20065);
nor U20520 (N_20520,N_20280,N_20010);
nor U20521 (N_20521,N_20306,N_20219);
and U20522 (N_20522,N_20218,N_20362);
nand U20523 (N_20523,N_20111,N_20081);
xnor U20524 (N_20524,N_20036,N_20357);
or U20525 (N_20525,N_20107,N_19989);
nand U20526 (N_20526,N_20241,N_20105);
nand U20527 (N_20527,N_20094,N_19914);
nor U20528 (N_20528,N_20397,N_19900);
nand U20529 (N_20529,N_20117,N_20380);
or U20530 (N_20530,N_20182,N_19854);
or U20531 (N_20531,N_19925,N_20368);
nand U20532 (N_20532,N_19886,N_19968);
or U20533 (N_20533,N_20074,N_20092);
and U20534 (N_20534,N_19923,N_20367);
or U20535 (N_20535,N_20282,N_19974);
nor U20536 (N_20536,N_20383,N_20214);
xnor U20537 (N_20537,N_19965,N_20347);
or U20538 (N_20538,N_20356,N_20157);
nor U20539 (N_20539,N_19819,N_20374);
nand U20540 (N_20540,N_19915,N_20196);
nor U20541 (N_20541,N_19830,N_20370);
or U20542 (N_20542,N_20227,N_20035);
nand U20543 (N_20543,N_20312,N_20130);
nand U20544 (N_20544,N_20278,N_20236);
or U20545 (N_20545,N_19921,N_20224);
nand U20546 (N_20546,N_20267,N_19917);
and U20547 (N_20547,N_20051,N_19918);
nor U20548 (N_20548,N_20014,N_19999);
and U20549 (N_20549,N_20078,N_20071);
nand U20550 (N_20550,N_20332,N_19883);
and U20551 (N_20551,N_19868,N_20022);
or U20552 (N_20552,N_20263,N_20123);
or U20553 (N_20553,N_19879,N_20118);
or U20554 (N_20554,N_20063,N_19899);
nand U20555 (N_20555,N_20011,N_19967);
nor U20556 (N_20556,N_20113,N_19855);
nor U20557 (N_20557,N_20279,N_19979);
or U20558 (N_20558,N_20034,N_20029);
nor U20559 (N_20559,N_19853,N_20069);
nor U20560 (N_20560,N_20056,N_20294);
and U20561 (N_20561,N_19816,N_20104);
nand U20562 (N_20562,N_19904,N_20273);
or U20563 (N_20563,N_20116,N_20222);
nand U20564 (N_20564,N_19874,N_20059);
xnor U20565 (N_20565,N_20256,N_20057);
nand U20566 (N_20566,N_19966,N_20244);
nor U20567 (N_20567,N_19846,N_19821);
or U20568 (N_20568,N_19948,N_19827);
and U20569 (N_20569,N_19982,N_20335);
and U20570 (N_20570,N_19843,N_20313);
nand U20571 (N_20571,N_19859,N_20097);
and U20572 (N_20572,N_19962,N_20140);
or U20573 (N_20573,N_20148,N_20246);
or U20574 (N_20574,N_20310,N_20298);
nand U20575 (N_20575,N_20292,N_20247);
or U20576 (N_20576,N_20103,N_20072);
nand U20577 (N_20577,N_20243,N_19972);
and U20578 (N_20578,N_20321,N_20205);
and U20579 (N_20579,N_20231,N_19803);
and U20580 (N_20580,N_19805,N_19811);
nor U20581 (N_20581,N_20291,N_20106);
and U20582 (N_20582,N_20201,N_20031);
nor U20583 (N_20583,N_20082,N_20237);
nand U20584 (N_20584,N_20076,N_19901);
nand U20585 (N_20585,N_19993,N_20204);
nor U20586 (N_20586,N_20364,N_20327);
xnor U20587 (N_20587,N_20142,N_19940);
nand U20588 (N_20588,N_20144,N_20189);
nand U20589 (N_20589,N_19888,N_20253);
nand U20590 (N_20590,N_20079,N_20026);
nor U20591 (N_20591,N_20308,N_20166);
or U20592 (N_20592,N_20046,N_20174);
and U20593 (N_20593,N_19906,N_20015);
nand U20594 (N_20594,N_20346,N_19958);
nand U20595 (N_20595,N_20127,N_19905);
nor U20596 (N_20596,N_20382,N_20255);
nand U20597 (N_20597,N_20341,N_19863);
and U20598 (N_20598,N_19858,N_20195);
nor U20599 (N_20599,N_19947,N_20027);
or U20600 (N_20600,N_20373,N_20032);
or U20601 (N_20601,N_19824,N_19987);
or U20602 (N_20602,N_20329,N_19834);
and U20603 (N_20603,N_20119,N_20339);
and U20604 (N_20604,N_19845,N_20270);
and U20605 (N_20605,N_20251,N_19810);
nand U20606 (N_20606,N_20050,N_20265);
nand U20607 (N_20607,N_20307,N_19857);
or U20608 (N_20608,N_20225,N_20328);
xor U20609 (N_20609,N_20396,N_19961);
or U20610 (N_20610,N_20399,N_19828);
or U20611 (N_20611,N_20200,N_19969);
nand U20612 (N_20612,N_20023,N_19802);
nor U20613 (N_20613,N_19927,N_20314);
and U20614 (N_20614,N_19932,N_20040);
nand U20615 (N_20615,N_20207,N_20334);
or U20616 (N_20616,N_19822,N_20232);
nand U20617 (N_20617,N_19924,N_20363);
nor U20618 (N_20618,N_20038,N_20020);
nand U20619 (N_20619,N_20143,N_20052);
or U20620 (N_20620,N_20338,N_20090);
or U20621 (N_20621,N_19909,N_20013);
nand U20622 (N_20622,N_20344,N_19889);
nor U20623 (N_20623,N_20348,N_20355);
nand U20624 (N_20624,N_20044,N_20365);
or U20625 (N_20625,N_19956,N_20066);
and U20626 (N_20626,N_19975,N_20047);
and U20627 (N_20627,N_19833,N_20371);
nand U20628 (N_20628,N_20268,N_19887);
and U20629 (N_20629,N_20145,N_19931);
nor U20630 (N_20630,N_19929,N_19864);
nor U20631 (N_20631,N_19971,N_20169);
and U20632 (N_20632,N_20336,N_20317);
nor U20633 (N_20633,N_20318,N_20378);
nand U20634 (N_20634,N_20322,N_19861);
nand U20635 (N_20635,N_20159,N_20325);
nand U20636 (N_20636,N_20352,N_19941);
and U20637 (N_20637,N_19949,N_20178);
or U20638 (N_20638,N_20060,N_20269);
nor U20639 (N_20639,N_20173,N_20226);
and U20640 (N_20640,N_19806,N_19933);
or U20641 (N_20641,N_20120,N_19980);
or U20642 (N_20642,N_19946,N_20096);
or U20643 (N_20643,N_19938,N_20125);
nor U20644 (N_20644,N_20080,N_20266);
nand U20645 (N_20645,N_20300,N_19986);
and U20646 (N_20646,N_19894,N_20077);
nand U20647 (N_20647,N_19985,N_20217);
or U20648 (N_20648,N_19804,N_20016);
nor U20649 (N_20649,N_20301,N_20045);
or U20650 (N_20650,N_20272,N_19841);
and U20651 (N_20651,N_20070,N_19869);
or U20652 (N_20652,N_19907,N_20276);
and U20653 (N_20653,N_19817,N_20048);
nand U20654 (N_20654,N_20331,N_20223);
nor U20655 (N_20655,N_19890,N_19995);
and U20656 (N_20656,N_19848,N_20303);
or U20657 (N_20657,N_20271,N_20095);
and U20658 (N_20658,N_19862,N_20186);
nor U20659 (N_20659,N_19950,N_19885);
or U20660 (N_20660,N_20206,N_19998);
nor U20661 (N_20661,N_20309,N_20093);
and U20662 (N_20662,N_20213,N_20375);
or U20663 (N_20663,N_19825,N_20361);
or U20664 (N_20664,N_20393,N_19908);
nor U20665 (N_20665,N_19882,N_20002);
nand U20666 (N_20666,N_20290,N_20067);
or U20667 (N_20667,N_20215,N_19902);
and U20668 (N_20668,N_19860,N_19840);
nor U20669 (N_20669,N_20283,N_20281);
nor U20670 (N_20670,N_20389,N_20210);
nand U20671 (N_20671,N_19897,N_20254);
nand U20672 (N_20672,N_20024,N_19954);
nand U20673 (N_20673,N_20379,N_20198);
nor U20674 (N_20674,N_20153,N_19898);
and U20675 (N_20675,N_20179,N_20343);
or U20676 (N_20676,N_19812,N_19955);
and U20677 (N_20677,N_20345,N_19891);
and U20678 (N_20678,N_19814,N_19820);
nand U20679 (N_20679,N_19837,N_19895);
xor U20680 (N_20680,N_19852,N_20295);
nor U20681 (N_20681,N_20089,N_19807);
and U20682 (N_20682,N_20073,N_20277);
nor U20683 (N_20683,N_20099,N_19920);
or U20684 (N_20684,N_20139,N_20152);
and U20685 (N_20685,N_20197,N_20248);
nor U20686 (N_20686,N_20042,N_20386);
or U20687 (N_20687,N_19977,N_20275);
nor U20688 (N_20688,N_19801,N_20030);
and U20689 (N_20689,N_19893,N_19818);
nor U20690 (N_20690,N_20129,N_19960);
and U20691 (N_20691,N_19973,N_19839);
or U20692 (N_20692,N_20007,N_20164);
or U20693 (N_20693,N_20239,N_19934);
and U20694 (N_20694,N_20184,N_20323);
or U20695 (N_20695,N_20049,N_19836);
and U20696 (N_20696,N_20163,N_19964);
or U20697 (N_20697,N_19881,N_19943);
xor U20698 (N_20698,N_19808,N_20025);
nand U20699 (N_20699,N_19913,N_20175);
and U20700 (N_20700,N_20289,N_20223);
nor U20701 (N_20701,N_20229,N_19862);
nor U20702 (N_20702,N_20284,N_20235);
or U20703 (N_20703,N_20165,N_19964);
or U20704 (N_20704,N_20110,N_19979);
nand U20705 (N_20705,N_20374,N_20083);
and U20706 (N_20706,N_20360,N_20244);
nand U20707 (N_20707,N_19843,N_20314);
nor U20708 (N_20708,N_20234,N_20233);
nor U20709 (N_20709,N_20347,N_20132);
and U20710 (N_20710,N_19959,N_20385);
nand U20711 (N_20711,N_19925,N_20099);
nor U20712 (N_20712,N_20356,N_20153);
nand U20713 (N_20713,N_19949,N_20296);
or U20714 (N_20714,N_20202,N_19964);
or U20715 (N_20715,N_19832,N_19974);
nor U20716 (N_20716,N_20353,N_20069);
nor U20717 (N_20717,N_20163,N_19915);
or U20718 (N_20718,N_19977,N_20144);
nand U20719 (N_20719,N_19814,N_20245);
and U20720 (N_20720,N_20009,N_19993);
or U20721 (N_20721,N_20120,N_20153);
nor U20722 (N_20722,N_19956,N_20089);
nor U20723 (N_20723,N_20050,N_20228);
nor U20724 (N_20724,N_20087,N_19982);
xnor U20725 (N_20725,N_19833,N_20392);
or U20726 (N_20726,N_20210,N_20002);
nor U20727 (N_20727,N_20146,N_20134);
nand U20728 (N_20728,N_19981,N_20229);
nand U20729 (N_20729,N_20270,N_20317);
and U20730 (N_20730,N_19890,N_20093);
nor U20731 (N_20731,N_19860,N_19985);
nand U20732 (N_20732,N_20281,N_20236);
nand U20733 (N_20733,N_20146,N_20373);
and U20734 (N_20734,N_20347,N_20362);
nor U20735 (N_20735,N_19834,N_20040);
or U20736 (N_20736,N_20297,N_20264);
or U20737 (N_20737,N_20303,N_19864);
nor U20738 (N_20738,N_19902,N_20348);
nand U20739 (N_20739,N_20029,N_20026);
xor U20740 (N_20740,N_19835,N_20240);
and U20741 (N_20741,N_19906,N_19804);
nor U20742 (N_20742,N_19865,N_20307);
and U20743 (N_20743,N_20061,N_20320);
and U20744 (N_20744,N_20275,N_19963);
nor U20745 (N_20745,N_19937,N_19867);
nand U20746 (N_20746,N_20020,N_20362);
and U20747 (N_20747,N_20335,N_19937);
or U20748 (N_20748,N_20164,N_20112);
or U20749 (N_20749,N_19900,N_20246);
or U20750 (N_20750,N_20361,N_20159);
and U20751 (N_20751,N_20306,N_19901);
xor U20752 (N_20752,N_20159,N_20145);
and U20753 (N_20753,N_20260,N_20385);
or U20754 (N_20754,N_20177,N_19800);
and U20755 (N_20755,N_20391,N_20361);
xnor U20756 (N_20756,N_20322,N_20200);
nor U20757 (N_20757,N_19838,N_20129);
nand U20758 (N_20758,N_20051,N_20274);
nor U20759 (N_20759,N_19915,N_20191);
or U20760 (N_20760,N_20171,N_20329);
or U20761 (N_20761,N_20337,N_19826);
nand U20762 (N_20762,N_20343,N_20255);
and U20763 (N_20763,N_19917,N_20184);
nor U20764 (N_20764,N_19982,N_20097);
nor U20765 (N_20765,N_19947,N_19844);
and U20766 (N_20766,N_19883,N_20320);
or U20767 (N_20767,N_19847,N_20390);
or U20768 (N_20768,N_20147,N_20326);
nand U20769 (N_20769,N_20253,N_20269);
nor U20770 (N_20770,N_20395,N_19929);
or U20771 (N_20771,N_19952,N_20029);
nand U20772 (N_20772,N_20204,N_20212);
and U20773 (N_20773,N_19930,N_19928);
or U20774 (N_20774,N_20023,N_19833);
xnor U20775 (N_20775,N_19801,N_20370);
nand U20776 (N_20776,N_20253,N_19965);
or U20777 (N_20777,N_20177,N_20107);
nor U20778 (N_20778,N_20372,N_19865);
and U20779 (N_20779,N_20386,N_20312);
nor U20780 (N_20780,N_20238,N_20389);
nor U20781 (N_20781,N_20227,N_19969);
and U20782 (N_20782,N_20061,N_19984);
nand U20783 (N_20783,N_20099,N_20142);
or U20784 (N_20784,N_20214,N_20056);
and U20785 (N_20785,N_20252,N_19854);
nor U20786 (N_20786,N_19861,N_20022);
nor U20787 (N_20787,N_20177,N_19811);
nor U20788 (N_20788,N_19939,N_19981);
nor U20789 (N_20789,N_19947,N_20023);
and U20790 (N_20790,N_20250,N_20032);
and U20791 (N_20791,N_20043,N_20391);
nor U20792 (N_20792,N_20383,N_19877);
xnor U20793 (N_20793,N_20203,N_20257);
nand U20794 (N_20794,N_20020,N_20223);
nor U20795 (N_20795,N_20036,N_20102);
or U20796 (N_20796,N_20382,N_20257);
nand U20797 (N_20797,N_19874,N_19918);
nor U20798 (N_20798,N_20200,N_20239);
or U20799 (N_20799,N_19892,N_20093);
or U20800 (N_20800,N_20001,N_20390);
nor U20801 (N_20801,N_19831,N_20384);
or U20802 (N_20802,N_20349,N_20246);
nand U20803 (N_20803,N_20328,N_19896);
and U20804 (N_20804,N_20392,N_19809);
or U20805 (N_20805,N_20003,N_20212);
or U20806 (N_20806,N_20048,N_20180);
nor U20807 (N_20807,N_20026,N_20008);
or U20808 (N_20808,N_20026,N_19927);
and U20809 (N_20809,N_20256,N_20044);
nand U20810 (N_20810,N_20350,N_20397);
xnor U20811 (N_20811,N_20386,N_20086);
nor U20812 (N_20812,N_20052,N_20342);
or U20813 (N_20813,N_20220,N_20012);
xor U20814 (N_20814,N_19904,N_19942);
or U20815 (N_20815,N_19966,N_19824);
nor U20816 (N_20816,N_19981,N_20051);
and U20817 (N_20817,N_20179,N_20030);
and U20818 (N_20818,N_19929,N_19836);
and U20819 (N_20819,N_20098,N_20182);
or U20820 (N_20820,N_20175,N_19861);
or U20821 (N_20821,N_19825,N_19923);
nor U20822 (N_20822,N_19829,N_19851);
nor U20823 (N_20823,N_20202,N_20390);
and U20824 (N_20824,N_20005,N_20026);
nor U20825 (N_20825,N_20027,N_20266);
or U20826 (N_20826,N_19897,N_19975);
or U20827 (N_20827,N_20244,N_20296);
and U20828 (N_20828,N_19933,N_20034);
nor U20829 (N_20829,N_19883,N_20267);
nand U20830 (N_20830,N_20253,N_19912);
or U20831 (N_20831,N_20261,N_19914);
nand U20832 (N_20832,N_20342,N_20359);
and U20833 (N_20833,N_20011,N_19880);
and U20834 (N_20834,N_20369,N_19992);
nor U20835 (N_20835,N_20009,N_20265);
and U20836 (N_20836,N_20279,N_20168);
and U20837 (N_20837,N_20152,N_20241);
or U20838 (N_20838,N_19856,N_19951);
and U20839 (N_20839,N_20287,N_20310);
and U20840 (N_20840,N_19844,N_19925);
nand U20841 (N_20841,N_20065,N_19968);
or U20842 (N_20842,N_20351,N_20123);
nand U20843 (N_20843,N_20214,N_20191);
or U20844 (N_20844,N_19936,N_20086);
xor U20845 (N_20845,N_20292,N_20234);
nand U20846 (N_20846,N_20060,N_20010);
nor U20847 (N_20847,N_20329,N_19907);
and U20848 (N_20848,N_20122,N_20294);
nor U20849 (N_20849,N_19899,N_20141);
or U20850 (N_20850,N_20270,N_19881);
and U20851 (N_20851,N_20019,N_19993);
and U20852 (N_20852,N_19843,N_19996);
and U20853 (N_20853,N_20078,N_20188);
and U20854 (N_20854,N_20260,N_20075);
or U20855 (N_20855,N_20002,N_20308);
or U20856 (N_20856,N_20192,N_20113);
nand U20857 (N_20857,N_20347,N_20131);
nor U20858 (N_20858,N_20397,N_19909);
nand U20859 (N_20859,N_20022,N_20186);
and U20860 (N_20860,N_20309,N_19802);
nand U20861 (N_20861,N_20070,N_20290);
nand U20862 (N_20862,N_20091,N_20007);
or U20863 (N_20863,N_20062,N_19867);
xor U20864 (N_20864,N_20265,N_20066);
nand U20865 (N_20865,N_19939,N_20029);
nor U20866 (N_20866,N_19986,N_20036);
nor U20867 (N_20867,N_19929,N_20025);
nor U20868 (N_20868,N_20270,N_19870);
or U20869 (N_20869,N_20166,N_20358);
or U20870 (N_20870,N_19838,N_19973);
and U20871 (N_20871,N_20237,N_19811);
nor U20872 (N_20872,N_19951,N_20368);
nand U20873 (N_20873,N_19920,N_19857);
nand U20874 (N_20874,N_20218,N_19936);
nand U20875 (N_20875,N_20280,N_20270);
nand U20876 (N_20876,N_20279,N_20380);
or U20877 (N_20877,N_20065,N_20168);
xnor U20878 (N_20878,N_20395,N_20381);
or U20879 (N_20879,N_20110,N_20317);
nor U20880 (N_20880,N_20149,N_20313);
nor U20881 (N_20881,N_20208,N_19901);
nand U20882 (N_20882,N_20152,N_20394);
nor U20883 (N_20883,N_20261,N_19910);
and U20884 (N_20884,N_20245,N_20007);
nor U20885 (N_20885,N_19928,N_20183);
nor U20886 (N_20886,N_19815,N_20039);
nand U20887 (N_20887,N_20029,N_20346);
and U20888 (N_20888,N_20397,N_20133);
nor U20889 (N_20889,N_20239,N_19866);
or U20890 (N_20890,N_19856,N_20105);
and U20891 (N_20891,N_19881,N_20359);
or U20892 (N_20892,N_20040,N_20192);
and U20893 (N_20893,N_20072,N_20170);
nor U20894 (N_20894,N_19894,N_19803);
or U20895 (N_20895,N_20038,N_19889);
nor U20896 (N_20896,N_20324,N_20038);
nor U20897 (N_20897,N_20114,N_20115);
or U20898 (N_20898,N_20031,N_20296);
or U20899 (N_20899,N_19993,N_20161);
nor U20900 (N_20900,N_20075,N_20253);
nor U20901 (N_20901,N_19920,N_20299);
and U20902 (N_20902,N_20286,N_19836);
nand U20903 (N_20903,N_20061,N_19970);
or U20904 (N_20904,N_20168,N_20029);
nand U20905 (N_20905,N_20074,N_19926);
nand U20906 (N_20906,N_20375,N_20341);
nor U20907 (N_20907,N_20204,N_19967);
or U20908 (N_20908,N_19835,N_20309);
and U20909 (N_20909,N_20223,N_19943);
or U20910 (N_20910,N_20325,N_19982);
nand U20911 (N_20911,N_20311,N_20049);
xor U20912 (N_20912,N_20247,N_19815);
nor U20913 (N_20913,N_19960,N_19978);
or U20914 (N_20914,N_19839,N_20025);
and U20915 (N_20915,N_19841,N_20312);
and U20916 (N_20916,N_20198,N_20047);
nand U20917 (N_20917,N_20234,N_19858);
nand U20918 (N_20918,N_20259,N_19952);
or U20919 (N_20919,N_20054,N_19997);
and U20920 (N_20920,N_20003,N_19999);
or U20921 (N_20921,N_20366,N_20358);
and U20922 (N_20922,N_20305,N_20141);
nand U20923 (N_20923,N_20317,N_20015);
nor U20924 (N_20924,N_20032,N_19949);
nand U20925 (N_20925,N_20180,N_20039);
and U20926 (N_20926,N_19875,N_20317);
nand U20927 (N_20927,N_20203,N_20264);
and U20928 (N_20928,N_20330,N_19982);
or U20929 (N_20929,N_20077,N_20303);
and U20930 (N_20930,N_20131,N_20085);
nor U20931 (N_20931,N_20175,N_20213);
nor U20932 (N_20932,N_19941,N_20256);
and U20933 (N_20933,N_20055,N_20127);
nand U20934 (N_20934,N_20163,N_20296);
and U20935 (N_20935,N_20285,N_20326);
or U20936 (N_20936,N_20145,N_20024);
nor U20937 (N_20937,N_20323,N_20018);
nor U20938 (N_20938,N_20193,N_20002);
and U20939 (N_20939,N_20298,N_20047);
nand U20940 (N_20940,N_19848,N_19822);
nand U20941 (N_20941,N_20241,N_20090);
or U20942 (N_20942,N_20047,N_20385);
and U20943 (N_20943,N_20133,N_20100);
nand U20944 (N_20944,N_20263,N_20116);
nand U20945 (N_20945,N_20322,N_19833);
and U20946 (N_20946,N_19947,N_20346);
nor U20947 (N_20947,N_19800,N_20193);
nand U20948 (N_20948,N_20132,N_20020);
and U20949 (N_20949,N_19845,N_20096);
and U20950 (N_20950,N_20137,N_20154);
nor U20951 (N_20951,N_20358,N_20020);
or U20952 (N_20952,N_19981,N_20097);
or U20953 (N_20953,N_20054,N_20394);
and U20954 (N_20954,N_19954,N_19873);
xnor U20955 (N_20955,N_19863,N_19942);
nand U20956 (N_20956,N_20084,N_20289);
nand U20957 (N_20957,N_20013,N_19994);
or U20958 (N_20958,N_19805,N_20004);
nor U20959 (N_20959,N_19830,N_19916);
or U20960 (N_20960,N_19958,N_20302);
and U20961 (N_20961,N_20182,N_20230);
nand U20962 (N_20962,N_19816,N_20387);
nand U20963 (N_20963,N_20259,N_20201);
xor U20964 (N_20964,N_19978,N_20043);
or U20965 (N_20965,N_19925,N_20325);
xor U20966 (N_20966,N_20241,N_19984);
and U20967 (N_20967,N_20194,N_20197);
nand U20968 (N_20968,N_20333,N_19820);
nand U20969 (N_20969,N_20342,N_20170);
nor U20970 (N_20970,N_20159,N_20375);
xor U20971 (N_20971,N_20056,N_20312);
and U20972 (N_20972,N_19873,N_20043);
and U20973 (N_20973,N_20309,N_19812);
nor U20974 (N_20974,N_20134,N_20013);
nand U20975 (N_20975,N_20166,N_20345);
and U20976 (N_20976,N_19839,N_19880);
and U20977 (N_20977,N_20178,N_20080);
nor U20978 (N_20978,N_19997,N_20010);
and U20979 (N_20979,N_20191,N_20371);
nand U20980 (N_20980,N_20361,N_20310);
or U20981 (N_20981,N_19950,N_19843);
xnor U20982 (N_20982,N_20235,N_20292);
nand U20983 (N_20983,N_19917,N_19843);
nor U20984 (N_20984,N_19995,N_20301);
nand U20985 (N_20985,N_19941,N_20349);
and U20986 (N_20986,N_20378,N_20035);
nand U20987 (N_20987,N_20183,N_20237);
nor U20988 (N_20988,N_20195,N_20394);
or U20989 (N_20989,N_19909,N_20212);
and U20990 (N_20990,N_20001,N_20245);
nand U20991 (N_20991,N_19959,N_20307);
nor U20992 (N_20992,N_20374,N_20330);
and U20993 (N_20993,N_19936,N_19920);
and U20994 (N_20994,N_19865,N_20344);
and U20995 (N_20995,N_20247,N_20356);
or U20996 (N_20996,N_20224,N_19858);
nand U20997 (N_20997,N_19914,N_19984);
or U20998 (N_20998,N_20168,N_19890);
or U20999 (N_20999,N_20116,N_20220);
nor U21000 (N_21000,N_20788,N_20467);
nor U21001 (N_21001,N_20742,N_20975);
nand U21002 (N_21002,N_20821,N_20765);
nand U21003 (N_21003,N_20564,N_20546);
nand U21004 (N_21004,N_20567,N_20422);
nand U21005 (N_21005,N_20496,N_20851);
nor U21006 (N_21006,N_20426,N_20405);
or U21007 (N_21007,N_20433,N_20540);
nand U21008 (N_21008,N_20593,N_20949);
or U21009 (N_21009,N_20648,N_20704);
nand U21010 (N_21010,N_20900,N_20558);
nor U21011 (N_21011,N_20459,N_20718);
and U21012 (N_21012,N_20635,N_20573);
or U21013 (N_21013,N_20694,N_20752);
nand U21014 (N_21014,N_20962,N_20557);
and U21015 (N_21015,N_20741,N_20491);
nand U21016 (N_21016,N_20645,N_20676);
and U21017 (N_21017,N_20611,N_20672);
nand U21018 (N_21018,N_20650,N_20753);
nand U21019 (N_21019,N_20657,N_20413);
or U21020 (N_21020,N_20563,N_20612);
nand U21021 (N_21021,N_20745,N_20907);
and U21022 (N_21022,N_20685,N_20568);
or U21023 (N_21023,N_20526,N_20522);
nor U21024 (N_21024,N_20455,N_20503);
nor U21025 (N_21025,N_20549,N_20743);
and U21026 (N_21026,N_20910,N_20968);
nand U21027 (N_21027,N_20516,N_20936);
or U21028 (N_21028,N_20410,N_20776);
and U21029 (N_21029,N_20875,N_20780);
and U21030 (N_21030,N_20616,N_20458);
and U21031 (N_21031,N_20690,N_20716);
nand U21032 (N_21032,N_20669,N_20946);
nor U21033 (N_21033,N_20698,N_20956);
and U21034 (N_21034,N_20644,N_20565);
or U21035 (N_21035,N_20935,N_20556);
or U21036 (N_21036,N_20592,N_20789);
nor U21037 (N_21037,N_20888,N_20518);
and U21038 (N_21038,N_20701,N_20705);
or U21039 (N_21039,N_20823,N_20554);
nand U21040 (N_21040,N_20819,N_20841);
nor U21041 (N_21041,N_20508,N_20476);
nor U21042 (N_21042,N_20871,N_20889);
nor U21043 (N_21043,N_20808,N_20586);
nor U21044 (N_21044,N_20629,N_20997);
and U21045 (N_21045,N_20805,N_20509);
nor U21046 (N_21046,N_20533,N_20983);
nand U21047 (N_21047,N_20506,N_20853);
nand U21048 (N_21048,N_20735,N_20639);
or U21049 (N_21049,N_20661,N_20763);
or U21050 (N_21050,N_20646,N_20441);
nor U21051 (N_21051,N_20621,N_20991);
xor U21052 (N_21052,N_20712,N_20996);
or U21053 (N_21053,N_20677,N_20489);
or U21054 (N_21054,N_20981,N_20670);
and U21055 (N_21055,N_20472,N_20658);
and U21056 (N_21056,N_20688,N_20449);
or U21057 (N_21057,N_20604,N_20757);
or U21058 (N_21058,N_20845,N_20969);
nor U21059 (N_21059,N_20746,N_20933);
or U21060 (N_21060,N_20487,N_20810);
nor U21061 (N_21061,N_20543,N_20477);
nand U21062 (N_21062,N_20750,N_20766);
or U21063 (N_21063,N_20758,N_20723);
xnor U21064 (N_21064,N_20727,N_20703);
or U21065 (N_21065,N_20793,N_20938);
or U21066 (N_21066,N_20964,N_20919);
xor U21067 (N_21067,N_20647,N_20811);
and U21068 (N_21068,N_20702,N_20451);
nor U21069 (N_21069,N_20905,N_20479);
nor U21070 (N_21070,N_20782,N_20597);
nor U21071 (N_21071,N_20667,N_20637);
or U21072 (N_21072,N_20510,N_20497);
and U21073 (N_21073,N_20867,N_20733);
and U21074 (N_21074,N_20896,N_20816);
or U21075 (N_21075,N_20992,N_20717);
nor U21076 (N_21076,N_20908,N_20885);
or U21077 (N_21077,N_20863,N_20493);
nand U21078 (N_21078,N_20801,N_20940);
or U21079 (N_21079,N_20684,N_20613);
nand U21080 (N_21080,N_20598,N_20777);
nand U21081 (N_21081,N_20686,N_20760);
and U21082 (N_21082,N_20924,N_20640);
and U21083 (N_21083,N_20427,N_20544);
nor U21084 (N_21084,N_20957,N_20580);
nand U21085 (N_21085,N_20502,N_20790);
nor U21086 (N_21086,N_20420,N_20706);
and U21087 (N_21087,N_20562,N_20797);
or U21088 (N_21088,N_20898,N_20680);
or U21089 (N_21089,N_20719,N_20673);
and U21090 (N_21090,N_20715,N_20649);
nor U21091 (N_21091,N_20878,N_20591);
nor U21092 (N_21092,N_20762,N_20600);
nand U21093 (N_21093,N_20903,N_20973);
or U21094 (N_21094,N_20605,N_20772);
nor U21095 (N_21095,N_20986,N_20585);
nor U21096 (N_21096,N_20577,N_20876);
or U21097 (N_21097,N_20833,N_20462);
or U21098 (N_21098,N_20836,N_20634);
or U21099 (N_21099,N_20707,N_20499);
nor U21100 (N_21100,N_20445,N_20967);
and U21101 (N_21101,N_20897,N_20872);
or U21102 (N_21102,N_20482,N_20978);
or U21103 (N_21103,N_20904,N_20525);
nand U21104 (N_21104,N_20572,N_20447);
and U21105 (N_21105,N_20662,N_20627);
nand U21106 (N_21106,N_20912,N_20636);
nor U21107 (N_21107,N_20504,N_20665);
nor U21108 (N_21108,N_20517,N_20831);
nor U21109 (N_21109,N_20976,N_20998);
and U21110 (N_21110,N_20434,N_20490);
nand U21111 (N_21111,N_20569,N_20519);
nand U21112 (N_21112,N_20521,N_20892);
and U21113 (N_21113,N_20838,N_20535);
nor U21114 (N_21114,N_20412,N_20681);
nand U21115 (N_21115,N_20817,N_20806);
nand U21116 (N_21116,N_20581,N_20773);
nor U21117 (N_21117,N_20980,N_20601);
nand U21118 (N_21118,N_20860,N_20800);
and U21119 (N_21119,N_20820,N_20920);
nand U21120 (N_21120,N_20843,N_20638);
or U21121 (N_21121,N_20982,N_20902);
xnor U21122 (N_21122,N_20664,N_20498);
nand U21123 (N_21123,N_20945,N_20767);
and U21124 (N_21124,N_20632,N_20439);
or U21125 (N_21125,N_20858,N_20622);
and U21126 (N_21126,N_20930,N_20401);
nand U21127 (N_21127,N_20740,N_20937);
or U21128 (N_21128,N_20744,N_20560);
xnor U21129 (N_21129,N_20881,N_20755);
and U21130 (N_21130,N_20775,N_20618);
nand U21131 (N_21131,N_20958,N_20660);
nor U21132 (N_21132,N_20927,N_20768);
nand U21133 (N_21133,N_20520,N_20666);
or U21134 (N_21134,N_20542,N_20751);
or U21135 (N_21135,N_20578,N_20699);
and U21136 (N_21136,N_20454,N_20834);
or U21137 (N_21137,N_20671,N_20737);
or U21138 (N_21138,N_20523,N_20785);
and U21139 (N_21139,N_20990,N_20424);
or U21140 (N_21140,N_20423,N_20994);
nand U21141 (N_21141,N_20692,N_20880);
nor U21142 (N_21142,N_20859,N_20915);
or U21143 (N_21143,N_20495,N_20473);
nand U21144 (N_21144,N_20720,N_20886);
nand U21145 (N_21145,N_20583,N_20448);
nor U21146 (N_21146,N_20799,N_20874);
nand U21147 (N_21147,N_20861,N_20494);
and U21148 (N_21148,N_20415,N_20784);
nand U21149 (N_21149,N_20961,N_20923);
and U21150 (N_21150,N_20713,N_20615);
or U21151 (N_21151,N_20804,N_20955);
nand U21152 (N_21152,N_20865,N_20548);
or U21153 (N_21153,N_20468,N_20759);
and U21154 (N_21154,N_20619,N_20417);
and U21155 (N_21155,N_20406,N_20608);
or U21156 (N_21156,N_20419,N_20749);
or U21157 (N_21157,N_20952,N_20827);
nand U21158 (N_21158,N_20626,N_20942);
nor U21159 (N_21159,N_20870,N_20890);
and U21160 (N_21160,N_20623,N_20478);
nor U21161 (N_21161,N_20628,N_20895);
or U21162 (N_21162,N_20527,N_20553);
or U21163 (N_21163,N_20989,N_20999);
nor U21164 (N_21164,N_20972,N_20798);
nand U21165 (N_21165,N_20446,N_20995);
nor U21166 (N_21166,N_20916,N_20435);
nand U21167 (N_21167,N_20862,N_20971);
and U21168 (N_21168,N_20954,N_20655);
nand U21169 (N_21169,N_20943,N_20425);
and U21170 (N_21170,N_20959,N_20812);
nand U21171 (N_21171,N_20529,N_20839);
xnor U21172 (N_21172,N_20595,N_20921);
xor U21173 (N_21173,N_20442,N_20829);
nor U21174 (N_21174,N_20480,N_20802);
nand U21175 (N_21175,N_20721,N_20579);
or U21176 (N_21176,N_20869,N_20436);
or U21177 (N_21177,N_20857,N_20584);
nor U21178 (N_21178,N_20963,N_20469);
nand U21179 (N_21179,N_20761,N_20939);
and U21180 (N_21180,N_20754,N_20475);
and U21181 (N_21181,N_20794,N_20428);
and U21182 (N_21182,N_20842,N_20643);
and U21183 (N_21183,N_20471,N_20465);
and U21184 (N_21184,N_20709,N_20879);
or U21185 (N_21185,N_20787,N_20414);
nor U21186 (N_21186,N_20620,N_20710);
and U21187 (N_21187,N_20732,N_20864);
or U21188 (N_21188,N_20965,N_20679);
or U21189 (N_21189,N_20404,N_20588);
nor U21190 (N_21190,N_20764,N_20736);
nand U21191 (N_21191,N_20697,N_20726);
nand U21192 (N_21192,N_20941,N_20734);
nor U21193 (N_21193,N_20505,N_20779);
nor U21194 (N_21194,N_20695,N_20411);
or U21195 (N_21195,N_20729,N_20571);
nand U21196 (N_21196,N_20599,N_20714);
nor U21197 (N_21197,N_20944,N_20663);
nor U21198 (N_21198,N_20534,N_20429);
nand U21199 (N_21199,N_20609,N_20481);
nand U21200 (N_21200,N_20748,N_20848);
and U21201 (N_21201,N_20687,N_20607);
or U21202 (N_21202,N_20537,N_20711);
nand U21203 (N_21203,N_20625,N_20561);
and U21204 (N_21204,N_20887,N_20911);
or U21205 (N_21205,N_20402,N_20722);
nor U21206 (N_21206,N_20840,N_20913);
nor U21207 (N_21207,N_20450,N_20691);
nor U21208 (N_21208,N_20539,N_20877);
nor U21209 (N_21209,N_20738,N_20431);
and U21210 (N_21210,N_20574,N_20500);
nand U21211 (N_21211,N_20416,N_20929);
or U21212 (N_21212,N_20984,N_20654);
or U21213 (N_21213,N_20977,N_20769);
or U21214 (N_21214,N_20594,N_20814);
nor U21215 (N_21215,N_20513,N_20507);
or U21216 (N_21216,N_20683,N_20825);
nor U21217 (N_21217,N_20771,N_20678);
or U21218 (N_21218,N_20795,N_20970);
and U21219 (N_21219,N_20610,N_20855);
and U21220 (N_21220,N_20545,N_20486);
or U21221 (N_21221,N_20532,N_20856);
nor U21222 (N_21222,N_20979,N_20642);
and U21223 (N_21223,N_20882,N_20925);
and U21224 (N_21224,N_20514,N_20570);
and U21225 (N_21225,N_20409,N_20974);
and U21226 (N_21226,N_20809,N_20541);
or U21227 (N_21227,N_20854,N_20488);
and U21228 (N_21228,N_20786,N_20651);
nor U21229 (N_21229,N_20689,N_20866);
or U21230 (N_21230,N_20538,N_20728);
and U21231 (N_21231,N_20682,N_20624);
nand U21232 (N_21232,N_20602,N_20407);
nand U21233 (N_21233,N_20403,N_20774);
or U21234 (N_21234,N_20452,N_20551);
nor U21235 (N_21235,N_20948,N_20928);
nor U21236 (N_21236,N_20512,N_20559);
nor U21237 (N_21237,N_20483,N_20575);
nor U21238 (N_21238,N_20674,N_20492);
nand U21239 (N_21239,N_20950,N_20832);
or U21240 (N_21240,N_20835,N_20536);
nor U21241 (N_21241,N_20756,N_20576);
nor U21242 (N_21242,N_20453,N_20530);
or U21243 (N_21243,N_20531,N_20653);
nor U21244 (N_21244,N_20730,N_20437);
nor U21245 (N_21245,N_20951,N_20985);
or U21246 (N_21246,N_20641,N_20466);
nand U21247 (N_21247,N_20914,N_20603);
nor U21248 (N_21248,N_20899,N_20747);
xnor U21249 (N_21249,N_20550,N_20891);
nor U21250 (N_21250,N_20731,N_20792);
and U21251 (N_21251,N_20852,N_20953);
nor U21252 (N_21252,N_20484,N_20659);
and U21253 (N_21253,N_20630,N_20515);
nor U21254 (N_21254,N_20818,N_20547);
or U21255 (N_21255,N_20693,N_20614);
and U21256 (N_21256,N_20807,N_20652);
or U21257 (N_21257,N_20464,N_20988);
xor U21258 (N_21258,N_20457,N_20668);
or U21259 (N_21259,N_20850,N_20778);
or U21260 (N_21260,N_20873,N_20883);
and U21261 (N_21261,N_20906,N_20631);
or U21262 (N_21262,N_20987,N_20418);
or U21263 (N_21263,N_20617,N_20931);
or U21264 (N_21264,N_20926,N_20606);
and U21265 (N_21265,N_20894,N_20633);
and U21266 (N_21266,N_20922,N_20770);
and U21267 (N_21267,N_20934,N_20511);
or U21268 (N_21268,N_20893,N_20708);
nand U21269 (N_21269,N_20917,N_20847);
nand U21270 (N_21270,N_20796,N_20824);
nor U21271 (N_21271,N_20444,N_20739);
nand U21272 (N_21272,N_20474,N_20837);
and U21273 (N_21273,N_20868,N_20781);
nor U21274 (N_21274,N_20918,N_20443);
and U21275 (N_21275,N_20590,N_20725);
or U21276 (N_21276,N_20438,N_20552);
or U21277 (N_21277,N_20589,N_20849);
or U21278 (N_21278,N_20815,N_20696);
nor U21279 (N_21279,N_20791,N_20966);
nor U21280 (N_21280,N_20528,N_20932);
and U21281 (N_21281,N_20408,N_20901);
or U21282 (N_21282,N_20461,N_20587);
xnor U21283 (N_21283,N_20460,N_20566);
nor U21284 (N_21284,N_20700,N_20485);
and U21285 (N_21285,N_20555,N_20844);
or U21286 (N_21286,N_20675,N_20993);
nor U21287 (N_21287,N_20947,N_20724);
nor U21288 (N_21288,N_20456,N_20432);
nand U21289 (N_21289,N_20846,N_20421);
xor U21290 (N_21290,N_20400,N_20830);
xnor U21291 (N_21291,N_20960,N_20440);
nand U21292 (N_21292,N_20596,N_20430);
nand U21293 (N_21293,N_20822,N_20463);
nand U21294 (N_21294,N_20470,N_20884);
nand U21295 (N_21295,N_20828,N_20909);
nor U21296 (N_21296,N_20813,N_20803);
nand U21297 (N_21297,N_20582,N_20656);
or U21298 (N_21298,N_20524,N_20501);
and U21299 (N_21299,N_20826,N_20783);
or U21300 (N_21300,N_20630,N_20559);
nand U21301 (N_21301,N_20920,N_20609);
nor U21302 (N_21302,N_20698,N_20614);
nand U21303 (N_21303,N_20553,N_20675);
and U21304 (N_21304,N_20831,N_20694);
nand U21305 (N_21305,N_20666,N_20441);
nor U21306 (N_21306,N_20439,N_20440);
or U21307 (N_21307,N_20453,N_20808);
or U21308 (N_21308,N_20904,N_20411);
and U21309 (N_21309,N_20460,N_20839);
nand U21310 (N_21310,N_20669,N_20912);
xnor U21311 (N_21311,N_20471,N_20692);
nor U21312 (N_21312,N_20775,N_20443);
and U21313 (N_21313,N_20750,N_20893);
and U21314 (N_21314,N_20554,N_20970);
and U21315 (N_21315,N_20801,N_20486);
xor U21316 (N_21316,N_20457,N_20416);
nor U21317 (N_21317,N_20625,N_20671);
nand U21318 (N_21318,N_20622,N_20612);
or U21319 (N_21319,N_20977,N_20788);
nand U21320 (N_21320,N_20979,N_20515);
or U21321 (N_21321,N_20531,N_20419);
nor U21322 (N_21322,N_20580,N_20801);
nor U21323 (N_21323,N_20872,N_20634);
or U21324 (N_21324,N_20971,N_20514);
and U21325 (N_21325,N_20521,N_20538);
nand U21326 (N_21326,N_20600,N_20470);
and U21327 (N_21327,N_20444,N_20894);
nor U21328 (N_21328,N_20486,N_20757);
or U21329 (N_21329,N_20780,N_20882);
nor U21330 (N_21330,N_20909,N_20576);
nor U21331 (N_21331,N_20865,N_20889);
and U21332 (N_21332,N_20921,N_20500);
nor U21333 (N_21333,N_20990,N_20471);
nor U21334 (N_21334,N_20976,N_20994);
and U21335 (N_21335,N_20893,N_20748);
or U21336 (N_21336,N_20731,N_20852);
nand U21337 (N_21337,N_20518,N_20751);
nor U21338 (N_21338,N_20902,N_20553);
and U21339 (N_21339,N_20824,N_20645);
and U21340 (N_21340,N_20510,N_20804);
nor U21341 (N_21341,N_20913,N_20625);
xor U21342 (N_21342,N_20877,N_20518);
or U21343 (N_21343,N_20630,N_20555);
and U21344 (N_21344,N_20945,N_20632);
or U21345 (N_21345,N_20917,N_20674);
and U21346 (N_21346,N_20903,N_20632);
and U21347 (N_21347,N_20797,N_20891);
and U21348 (N_21348,N_20911,N_20460);
xnor U21349 (N_21349,N_20925,N_20878);
and U21350 (N_21350,N_20570,N_20540);
or U21351 (N_21351,N_20797,N_20896);
or U21352 (N_21352,N_20828,N_20957);
and U21353 (N_21353,N_20907,N_20582);
or U21354 (N_21354,N_20744,N_20666);
nor U21355 (N_21355,N_20618,N_20504);
and U21356 (N_21356,N_20910,N_20672);
and U21357 (N_21357,N_20686,N_20784);
or U21358 (N_21358,N_20490,N_20675);
nor U21359 (N_21359,N_20818,N_20763);
and U21360 (N_21360,N_20608,N_20898);
nor U21361 (N_21361,N_20720,N_20461);
nor U21362 (N_21362,N_20923,N_20840);
or U21363 (N_21363,N_20647,N_20899);
nand U21364 (N_21364,N_20433,N_20454);
or U21365 (N_21365,N_20611,N_20858);
nor U21366 (N_21366,N_20911,N_20953);
nand U21367 (N_21367,N_20725,N_20929);
nand U21368 (N_21368,N_20473,N_20979);
and U21369 (N_21369,N_20458,N_20878);
nand U21370 (N_21370,N_20955,N_20607);
and U21371 (N_21371,N_20964,N_20848);
and U21372 (N_21372,N_20615,N_20816);
and U21373 (N_21373,N_20655,N_20647);
nand U21374 (N_21374,N_20684,N_20495);
or U21375 (N_21375,N_20870,N_20881);
or U21376 (N_21376,N_20816,N_20611);
nand U21377 (N_21377,N_20852,N_20565);
nor U21378 (N_21378,N_20707,N_20954);
nand U21379 (N_21379,N_20682,N_20928);
nand U21380 (N_21380,N_20645,N_20467);
or U21381 (N_21381,N_20422,N_20784);
nand U21382 (N_21382,N_20629,N_20682);
nor U21383 (N_21383,N_20759,N_20646);
nand U21384 (N_21384,N_20521,N_20996);
nand U21385 (N_21385,N_20963,N_20562);
nor U21386 (N_21386,N_20929,N_20620);
nor U21387 (N_21387,N_20489,N_20436);
nand U21388 (N_21388,N_20943,N_20607);
or U21389 (N_21389,N_20762,N_20752);
or U21390 (N_21390,N_20444,N_20994);
nand U21391 (N_21391,N_20535,N_20936);
nand U21392 (N_21392,N_20520,N_20578);
nand U21393 (N_21393,N_20959,N_20750);
and U21394 (N_21394,N_20791,N_20856);
or U21395 (N_21395,N_20507,N_20993);
nand U21396 (N_21396,N_20442,N_20710);
and U21397 (N_21397,N_20659,N_20628);
and U21398 (N_21398,N_20451,N_20813);
or U21399 (N_21399,N_20639,N_20885);
nand U21400 (N_21400,N_20853,N_20602);
nor U21401 (N_21401,N_20439,N_20615);
nor U21402 (N_21402,N_20807,N_20693);
and U21403 (N_21403,N_20699,N_20508);
xor U21404 (N_21404,N_20932,N_20612);
and U21405 (N_21405,N_20498,N_20522);
nor U21406 (N_21406,N_20753,N_20498);
nor U21407 (N_21407,N_20675,N_20486);
xor U21408 (N_21408,N_20602,N_20638);
nand U21409 (N_21409,N_20868,N_20761);
and U21410 (N_21410,N_20608,N_20750);
nor U21411 (N_21411,N_20830,N_20555);
or U21412 (N_21412,N_20467,N_20631);
or U21413 (N_21413,N_20974,N_20780);
nand U21414 (N_21414,N_20883,N_20512);
and U21415 (N_21415,N_20520,N_20734);
or U21416 (N_21416,N_20563,N_20429);
or U21417 (N_21417,N_20993,N_20645);
nand U21418 (N_21418,N_20707,N_20946);
nand U21419 (N_21419,N_20494,N_20751);
and U21420 (N_21420,N_20474,N_20911);
or U21421 (N_21421,N_20545,N_20889);
nor U21422 (N_21422,N_20495,N_20790);
nor U21423 (N_21423,N_20450,N_20628);
and U21424 (N_21424,N_20775,N_20855);
nor U21425 (N_21425,N_20624,N_20869);
and U21426 (N_21426,N_20926,N_20887);
or U21427 (N_21427,N_20904,N_20809);
nand U21428 (N_21428,N_20673,N_20406);
or U21429 (N_21429,N_20845,N_20775);
or U21430 (N_21430,N_20802,N_20883);
nand U21431 (N_21431,N_20493,N_20864);
nand U21432 (N_21432,N_20886,N_20860);
nand U21433 (N_21433,N_20909,N_20888);
or U21434 (N_21434,N_20951,N_20452);
and U21435 (N_21435,N_20752,N_20742);
nand U21436 (N_21436,N_20657,N_20485);
and U21437 (N_21437,N_20699,N_20524);
and U21438 (N_21438,N_20552,N_20886);
nor U21439 (N_21439,N_20505,N_20752);
nand U21440 (N_21440,N_20913,N_20830);
and U21441 (N_21441,N_20675,N_20878);
and U21442 (N_21442,N_20925,N_20843);
nand U21443 (N_21443,N_20475,N_20430);
nor U21444 (N_21444,N_20666,N_20435);
nand U21445 (N_21445,N_20504,N_20472);
and U21446 (N_21446,N_20778,N_20411);
and U21447 (N_21447,N_20647,N_20671);
or U21448 (N_21448,N_20938,N_20956);
and U21449 (N_21449,N_20411,N_20797);
or U21450 (N_21450,N_20797,N_20771);
nand U21451 (N_21451,N_20419,N_20409);
nand U21452 (N_21452,N_20930,N_20945);
or U21453 (N_21453,N_20754,N_20474);
and U21454 (N_21454,N_20599,N_20550);
nor U21455 (N_21455,N_20401,N_20438);
and U21456 (N_21456,N_20738,N_20710);
nand U21457 (N_21457,N_20725,N_20424);
and U21458 (N_21458,N_20495,N_20789);
nand U21459 (N_21459,N_20416,N_20893);
nor U21460 (N_21460,N_20953,N_20896);
and U21461 (N_21461,N_20601,N_20447);
or U21462 (N_21462,N_20928,N_20548);
and U21463 (N_21463,N_20921,N_20758);
and U21464 (N_21464,N_20556,N_20927);
nor U21465 (N_21465,N_20627,N_20832);
nand U21466 (N_21466,N_20657,N_20990);
nand U21467 (N_21467,N_20670,N_20936);
nand U21468 (N_21468,N_20952,N_20440);
nand U21469 (N_21469,N_20516,N_20932);
and U21470 (N_21470,N_20961,N_20445);
nand U21471 (N_21471,N_20466,N_20646);
or U21472 (N_21472,N_20648,N_20439);
or U21473 (N_21473,N_20401,N_20601);
and U21474 (N_21474,N_20887,N_20661);
or U21475 (N_21475,N_20751,N_20823);
nor U21476 (N_21476,N_20850,N_20631);
and U21477 (N_21477,N_20818,N_20441);
nor U21478 (N_21478,N_20608,N_20763);
nand U21479 (N_21479,N_20460,N_20407);
nand U21480 (N_21480,N_20527,N_20476);
nor U21481 (N_21481,N_20487,N_20982);
and U21482 (N_21482,N_20906,N_20553);
nand U21483 (N_21483,N_20579,N_20964);
nor U21484 (N_21484,N_20910,N_20464);
xnor U21485 (N_21485,N_20894,N_20675);
and U21486 (N_21486,N_20972,N_20855);
or U21487 (N_21487,N_20496,N_20959);
nor U21488 (N_21488,N_20616,N_20674);
or U21489 (N_21489,N_20470,N_20415);
nor U21490 (N_21490,N_20663,N_20657);
or U21491 (N_21491,N_20518,N_20684);
nor U21492 (N_21492,N_20829,N_20612);
nand U21493 (N_21493,N_20400,N_20516);
or U21494 (N_21494,N_20489,N_20708);
and U21495 (N_21495,N_20766,N_20546);
and U21496 (N_21496,N_20687,N_20760);
and U21497 (N_21497,N_20836,N_20873);
and U21498 (N_21498,N_20562,N_20594);
and U21499 (N_21499,N_20601,N_20969);
nand U21500 (N_21500,N_20422,N_20507);
xor U21501 (N_21501,N_20768,N_20612);
nor U21502 (N_21502,N_20937,N_20405);
nand U21503 (N_21503,N_20916,N_20795);
nand U21504 (N_21504,N_20466,N_20983);
nand U21505 (N_21505,N_20708,N_20776);
and U21506 (N_21506,N_20599,N_20517);
nor U21507 (N_21507,N_20808,N_20757);
nor U21508 (N_21508,N_20689,N_20451);
nand U21509 (N_21509,N_20602,N_20657);
nand U21510 (N_21510,N_20924,N_20776);
nand U21511 (N_21511,N_20763,N_20901);
and U21512 (N_21512,N_20588,N_20983);
nand U21513 (N_21513,N_20519,N_20857);
or U21514 (N_21514,N_20448,N_20682);
and U21515 (N_21515,N_20566,N_20846);
nor U21516 (N_21516,N_20751,N_20798);
nor U21517 (N_21517,N_20912,N_20533);
nor U21518 (N_21518,N_20846,N_20854);
or U21519 (N_21519,N_20612,N_20865);
xor U21520 (N_21520,N_20403,N_20467);
nor U21521 (N_21521,N_20702,N_20540);
nor U21522 (N_21522,N_20656,N_20980);
or U21523 (N_21523,N_20868,N_20875);
or U21524 (N_21524,N_20837,N_20572);
and U21525 (N_21525,N_20790,N_20428);
nor U21526 (N_21526,N_20697,N_20653);
or U21527 (N_21527,N_20601,N_20571);
xor U21528 (N_21528,N_20683,N_20662);
and U21529 (N_21529,N_20734,N_20564);
or U21530 (N_21530,N_20477,N_20875);
nand U21531 (N_21531,N_20665,N_20501);
and U21532 (N_21532,N_20997,N_20967);
nand U21533 (N_21533,N_20623,N_20405);
nand U21534 (N_21534,N_20655,N_20981);
nor U21535 (N_21535,N_20931,N_20614);
nand U21536 (N_21536,N_20565,N_20993);
nand U21537 (N_21537,N_20634,N_20510);
nand U21538 (N_21538,N_20753,N_20969);
or U21539 (N_21539,N_20648,N_20444);
nor U21540 (N_21540,N_20669,N_20942);
and U21541 (N_21541,N_20822,N_20612);
or U21542 (N_21542,N_20681,N_20481);
nor U21543 (N_21543,N_20721,N_20736);
or U21544 (N_21544,N_20479,N_20440);
or U21545 (N_21545,N_20608,N_20593);
or U21546 (N_21546,N_20630,N_20807);
nor U21547 (N_21547,N_20906,N_20984);
xnor U21548 (N_21548,N_20402,N_20858);
nor U21549 (N_21549,N_20451,N_20542);
nor U21550 (N_21550,N_20930,N_20859);
and U21551 (N_21551,N_20721,N_20824);
nor U21552 (N_21552,N_20837,N_20834);
nand U21553 (N_21553,N_20558,N_20433);
or U21554 (N_21554,N_20612,N_20648);
and U21555 (N_21555,N_20412,N_20798);
nand U21556 (N_21556,N_20975,N_20666);
xnor U21557 (N_21557,N_20552,N_20596);
nand U21558 (N_21558,N_20888,N_20603);
nand U21559 (N_21559,N_20788,N_20749);
nor U21560 (N_21560,N_20889,N_20635);
nor U21561 (N_21561,N_20563,N_20646);
or U21562 (N_21562,N_20463,N_20736);
or U21563 (N_21563,N_20885,N_20477);
and U21564 (N_21564,N_20744,N_20861);
nand U21565 (N_21565,N_20966,N_20970);
and U21566 (N_21566,N_20943,N_20511);
nand U21567 (N_21567,N_20827,N_20937);
nand U21568 (N_21568,N_20943,N_20416);
xnor U21569 (N_21569,N_20989,N_20925);
and U21570 (N_21570,N_20682,N_20413);
nor U21571 (N_21571,N_20843,N_20471);
or U21572 (N_21572,N_20604,N_20639);
and U21573 (N_21573,N_20678,N_20458);
or U21574 (N_21574,N_20471,N_20481);
nor U21575 (N_21575,N_20882,N_20550);
or U21576 (N_21576,N_20939,N_20869);
nor U21577 (N_21577,N_20907,N_20733);
or U21578 (N_21578,N_20416,N_20608);
nand U21579 (N_21579,N_20903,N_20782);
and U21580 (N_21580,N_20686,N_20879);
or U21581 (N_21581,N_20624,N_20489);
nand U21582 (N_21582,N_20850,N_20567);
nor U21583 (N_21583,N_20973,N_20727);
xor U21584 (N_21584,N_20620,N_20488);
and U21585 (N_21585,N_20958,N_20763);
or U21586 (N_21586,N_20860,N_20453);
and U21587 (N_21587,N_20811,N_20723);
nor U21588 (N_21588,N_20444,N_20792);
or U21589 (N_21589,N_20695,N_20832);
or U21590 (N_21590,N_20658,N_20564);
and U21591 (N_21591,N_20600,N_20759);
and U21592 (N_21592,N_20491,N_20863);
nand U21593 (N_21593,N_20959,N_20589);
or U21594 (N_21594,N_20466,N_20495);
and U21595 (N_21595,N_20510,N_20480);
and U21596 (N_21596,N_20599,N_20540);
or U21597 (N_21597,N_20776,N_20878);
nand U21598 (N_21598,N_20922,N_20893);
nor U21599 (N_21599,N_20938,N_20922);
nor U21600 (N_21600,N_21244,N_21175);
or U21601 (N_21601,N_21193,N_21549);
and U21602 (N_21602,N_21509,N_21168);
or U21603 (N_21603,N_21017,N_21043);
and U21604 (N_21604,N_21054,N_21026);
nor U21605 (N_21605,N_21520,N_21273);
nor U21606 (N_21606,N_21476,N_21535);
and U21607 (N_21607,N_21416,N_21167);
nand U21608 (N_21608,N_21100,N_21363);
nand U21609 (N_21609,N_21231,N_21032);
and U21610 (N_21610,N_21492,N_21178);
and U21611 (N_21611,N_21420,N_21539);
or U21612 (N_21612,N_21162,N_21091);
and U21613 (N_21613,N_21240,N_21551);
and U21614 (N_21614,N_21394,N_21134);
nand U21615 (N_21615,N_21560,N_21269);
nor U21616 (N_21616,N_21357,N_21454);
and U21617 (N_21617,N_21112,N_21409);
and U21618 (N_21618,N_21428,N_21086);
and U21619 (N_21619,N_21139,N_21505);
xor U21620 (N_21620,N_21197,N_21374);
xnor U21621 (N_21621,N_21141,N_21270);
or U21622 (N_21622,N_21070,N_21384);
nor U21623 (N_21623,N_21326,N_21439);
nand U21624 (N_21624,N_21554,N_21500);
nor U21625 (N_21625,N_21351,N_21506);
nor U21626 (N_21626,N_21576,N_21315);
and U21627 (N_21627,N_21460,N_21275);
xnor U21628 (N_21628,N_21307,N_21120);
or U21629 (N_21629,N_21172,N_21272);
nor U21630 (N_21630,N_21446,N_21156);
xnor U21631 (N_21631,N_21138,N_21569);
nor U21632 (N_21632,N_21195,N_21425);
nor U21633 (N_21633,N_21128,N_21053);
nand U21634 (N_21634,N_21084,N_21410);
and U21635 (N_21635,N_21513,N_21572);
nand U21636 (N_21636,N_21190,N_21408);
nand U21637 (N_21637,N_21573,N_21238);
nand U21638 (N_21638,N_21228,N_21164);
or U21639 (N_21639,N_21342,N_21267);
nor U21640 (N_21640,N_21057,N_21562);
and U21641 (N_21641,N_21237,N_21246);
nor U21642 (N_21642,N_21419,N_21458);
nor U21643 (N_21643,N_21119,N_21504);
nand U21644 (N_21644,N_21249,N_21241);
or U21645 (N_21645,N_21113,N_21177);
nor U21646 (N_21646,N_21438,N_21290);
nand U21647 (N_21647,N_21591,N_21180);
nand U21648 (N_21648,N_21466,N_21088);
or U21649 (N_21649,N_21482,N_21372);
and U21650 (N_21650,N_21470,N_21581);
nand U21651 (N_21651,N_21340,N_21108);
or U21652 (N_21652,N_21004,N_21255);
and U21653 (N_21653,N_21503,N_21391);
nor U21654 (N_21654,N_21523,N_21035);
and U21655 (N_21655,N_21336,N_21015);
nor U21656 (N_21656,N_21265,N_21214);
and U21657 (N_21657,N_21296,N_21349);
and U21658 (N_21658,N_21499,N_21327);
or U21659 (N_21659,N_21400,N_21486);
nor U21660 (N_21660,N_21395,N_21516);
xnor U21661 (N_21661,N_21302,N_21297);
and U21662 (N_21662,N_21510,N_21188);
nor U21663 (N_21663,N_21056,N_21397);
and U21664 (N_21664,N_21335,N_21060);
nor U21665 (N_21665,N_21239,N_21300);
and U21666 (N_21666,N_21203,N_21483);
and U21667 (N_21667,N_21117,N_21089);
nor U21668 (N_21668,N_21079,N_21271);
or U21669 (N_21669,N_21251,N_21532);
and U21670 (N_21670,N_21110,N_21046);
xor U21671 (N_21671,N_21555,N_21437);
nand U21672 (N_21672,N_21588,N_21536);
or U21673 (N_21673,N_21316,N_21266);
nor U21674 (N_21674,N_21192,N_21430);
nand U21675 (N_21675,N_21145,N_21033);
and U21676 (N_21676,N_21081,N_21051);
and U21677 (N_21677,N_21559,N_21348);
or U21678 (N_21678,N_21097,N_21455);
nand U21679 (N_21679,N_21518,N_21501);
or U21680 (N_21680,N_21194,N_21163);
nor U21681 (N_21681,N_21008,N_21161);
nand U21682 (N_21682,N_21260,N_21373);
nor U21683 (N_21683,N_21223,N_21078);
nor U21684 (N_21684,N_21441,N_21107);
nand U21685 (N_21685,N_21157,N_21567);
nand U21686 (N_21686,N_21146,N_21544);
nor U21687 (N_21687,N_21289,N_21069);
nor U21688 (N_21688,N_21375,N_21392);
nor U21689 (N_21689,N_21538,N_21218);
and U21690 (N_21690,N_21072,N_21371);
nor U21691 (N_21691,N_21450,N_21390);
nor U21692 (N_21692,N_21250,N_21147);
and U21693 (N_21693,N_21012,N_21528);
and U21694 (N_21694,N_21073,N_21417);
and U21695 (N_21695,N_21023,N_21028);
or U21696 (N_21696,N_21599,N_21596);
and U21697 (N_21697,N_21489,N_21341);
and U21698 (N_21698,N_21323,N_21337);
nand U21699 (N_21699,N_21338,N_21074);
or U21700 (N_21700,N_21469,N_21024);
and U21701 (N_21701,N_21031,N_21103);
nand U21702 (N_21702,N_21062,N_21405);
nor U21703 (N_21703,N_21354,N_21122);
nor U21704 (N_21704,N_21463,N_21537);
nor U21705 (N_21705,N_21459,N_21189);
nor U21706 (N_21706,N_21521,N_21461);
or U21707 (N_21707,N_21176,N_21093);
nand U21708 (N_21708,N_21383,N_21075);
nand U21709 (N_21709,N_21123,N_21243);
nor U21710 (N_21710,N_21570,N_21380);
or U21711 (N_21711,N_21472,N_21369);
nor U21712 (N_21712,N_21515,N_21467);
and U21713 (N_21713,N_21159,N_21215);
or U21714 (N_21714,N_21477,N_21353);
nand U21715 (N_21715,N_21452,N_21333);
nor U21716 (N_21716,N_21552,N_21487);
xor U21717 (N_21717,N_21519,N_21421);
nand U21718 (N_21718,N_21011,N_21099);
nor U21719 (N_21719,N_21213,N_21038);
nor U21720 (N_21720,N_21232,N_21433);
and U21721 (N_21721,N_21451,N_21435);
nor U21722 (N_21722,N_21236,N_21235);
xnor U21723 (N_21723,N_21334,N_21484);
nand U21724 (N_21724,N_21402,N_21136);
or U21725 (N_21725,N_21245,N_21283);
nand U21726 (N_21726,N_21474,N_21185);
nand U21727 (N_21727,N_21140,N_21366);
nor U21728 (N_21728,N_21219,N_21564);
nor U21729 (N_21729,N_21036,N_21007);
nand U21730 (N_21730,N_21277,N_21558);
nand U21731 (N_21731,N_21264,N_21048);
or U21732 (N_21732,N_21382,N_21115);
or U21733 (N_21733,N_21594,N_21456);
or U21734 (N_21734,N_21016,N_21527);
or U21735 (N_21735,N_21018,N_21149);
nor U21736 (N_21736,N_21102,N_21131);
nand U21737 (N_21737,N_21111,N_21066);
or U21738 (N_21738,N_21044,N_21095);
xnor U21739 (N_21739,N_21059,N_21339);
nand U21740 (N_21740,N_21013,N_21222);
nor U21741 (N_21741,N_21049,N_21396);
nor U21742 (N_21742,N_21352,N_21155);
nor U21743 (N_21743,N_21135,N_21288);
nor U21744 (N_21744,N_21406,N_21005);
nor U21745 (N_21745,N_21468,N_21313);
and U21746 (N_21746,N_21432,N_21385);
nand U21747 (N_21747,N_21173,N_21531);
nand U21748 (N_21748,N_21186,N_21129);
nand U21749 (N_21749,N_21256,N_21566);
nand U21750 (N_21750,N_21478,N_21465);
or U21751 (N_21751,N_21006,N_21442);
or U21752 (N_21752,N_21169,N_21423);
nor U21753 (N_21753,N_21584,N_21052);
and U21754 (N_21754,N_21359,N_21233);
and U21755 (N_21755,N_21087,N_21497);
and U21756 (N_21756,N_21152,N_21144);
and U21757 (N_21757,N_21041,N_21199);
nor U21758 (N_21758,N_21029,N_21274);
and U21759 (N_21759,N_21565,N_21325);
nand U21760 (N_21760,N_21511,N_21597);
or U21761 (N_21761,N_21258,N_21303);
and U21762 (N_21762,N_21047,N_21291);
and U21763 (N_21763,N_21488,N_21183);
nand U21764 (N_21764,N_21512,N_21116);
nand U21765 (N_21765,N_21356,N_21347);
nor U21766 (N_21766,N_21401,N_21317);
nand U21767 (N_21767,N_21328,N_21431);
nand U21768 (N_21768,N_21127,N_21225);
xor U21769 (N_21769,N_21201,N_21496);
and U21770 (N_21770,N_21436,N_21118);
or U21771 (N_21771,N_21321,N_21252);
or U21772 (N_21772,N_21298,N_21226);
or U21773 (N_21773,N_21083,N_21211);
and U21774 (N_21774,N_21076,N_21418);
or U21775 (N_21775,N_21548,N_21268);
or U21776 (N_21776,N_21310,N_21479);
nor U21777 (N_21777,N_21216,N_21114);
or U21778 (N_21778,N_21568,N_21301);
nand U21779 (N_21779,N_21593,N_21386);
nand U21780 (N_21780,N_21376,N_21200);
or U21781 (N_21781,N_21541,N_21229);
or U21782 (N_21782,N_21257,N_21247);
or U21783 (N_21783,N_21098,N_21507);
nand U21784 (N_21784,N_21227,N_21556);
nand U21785 (N_21785,N_21282,N_21133);
or U21786 (N_21786,N_21319,N_21485);
and U21787 (N_21787,N_21377,N_21404);
and U21788 (N_21788,N_21312,N_21368);
nor U21789 (N_21789,N_21475,N_21457);
or U21790 (N_21790,N_21039,N_21550);
and U21791 (N_21791,N_21045,N_21585);
or U21792 (N_21792,N_21151,N_21050);
nand U21793 (N_21793,N_21294,N_21305);
nor U21794 (N_21794,N_21579,N_21153);
and U21795 (N_21795,N_21025,N_21329);
and U21796 (N_21796,N_21055,N_21170);
and U21797 (N_21797,N_21571,N_21158);
nor U21798 (N_21798,N_21480,N_21582);
and U21799 (N_21799,N_21595,N_21242);
and U21800 (N_21800,N_21105,N_21292);
xnor U21801 (N_21801,N_21525,N_21148);
and U21802 (N_21802,N_21022,N_21137);
xnor U21803 (N_21803,N_21132,N_21592);
xor U21804 (N_21804,N_21577,N_21355);
and U21805 (N_21805,N_21540,N_21104);
nand U21806 (N_21806,N_21322,N_21003);
nor U21807 (N_21807,N_21142,N_21449);
or U21808 (N_21808,N_21443,N_21171);
or U21809 (N_21809,N_21524,N_21030);
nor U21810 (N_21810,N_21473,N_21403);
or U21811 (N_21811,N_21364,N_21434);
nand U21812 (N_21812,N_21285,N_21165);
nand U21813 (N_21813,N_21224,N_21278);
or U21814 (N_21814,N_21557,N_21179);
nor U21815 (N_21815,N_21002,N_21209);
and U21816 (N_21816,N_21064,N_21414);
nor U21817 (N_21817,N_21365,N_21314);
nand U21818 (N_21818,N_21346,N_21308);
or U21819 (N_21819,N_21514,N_21220);
nand U21820 (N_21820,N_21561,N_21361);
nand U21821 (N_21821,N_21208,N_21206);
nand U21822 (N_21822,N_21553,N_21331);
nand U21823 (N_21823,N_21526,N_21563);
nand U21824 (N_21824,N_21306,N_21412);
and U21825 (N_21825,N_21261,N_21543);
or U21826 (N_21826,N_21362,N_21077);
and U21827 (N_21827,N_21350,N_21534);
nor U21828 (N_21828,N_21590,N_21181);
nor U21829 (N_21829,N_21445,N_21299);
nand U21830 (N_21830,N_21085,N_21109);
nand U21831 (N_21831,N_21575,N_21174);
nand U21832 (N_21832,N_21040,N_21295);
nor U21833 (N_21833,N_21533,N_21106);
nor U21834 (N_21834,N_21330,N_21580);
nand U21835 (N_21835,N_21094,N_21517);
and U21836 (N_21836,N_21286,N_21530);
nor U21837 (N_21837,N_21453,N_21014);
nand U21838 (N_21838,N_21370,N_21000);
and U21839 (N_21839,N_21358,N_21399);
nand U21840 (N_21840,N_21279,N_21124);
nor U21841 (N_21841,N_21184,N_21393);
or U21842 (N_21842,N_21490,N_21378);
and U21843 (N_21843,N_21276,N_21034);
or U21844 (N_21844,N_21589,N_21198);
nand U21845 (N_21845,N_21191,N_21262);
and U21846 (N_21846,N_21293,N_21481);
or U21847 (N_21847,N_21101,N_21381);
nand U21848 (N_21848,N_21387,N_21360);
and U21849 (N_21849,N_21429,N_21529);
xor U21850 (N_21850,N_21212,N_21210);
or U21851 (N_21851,N_21065,N_21154);
nor U21852 (N_21852,N_21494,N_21063);
and U21853 (N_21853,N_21121,N_21281);
and U21854 (N_21854,N_21096,N_21587);
nand U21855 (N_21855,N_21187,N_21042);
nand U21856 (N_21856,N_21309,N_21440);
and U21857 (N_21857,N_21068,N_21166);
and U21858 (N_21858,N_21343,N_21304);
or U21859 (N_21859,N_21259,N_21160);
nor U21860 (N_21860,N_21027,N_21471);
or U21861 (N_21861,N_21508,N_21082);
nand U21862 (N_21862,N_21125,N_21495);
or U21863 (N_21863,N_21324,N_21345);
nor U21864 (N_21864,N_21126,N_21221);
and U21865 (N_21865,N_21407,N_21411);
or U21866 (N_21866,N_21422,N_21586);
nand U21867 (N_21867,N_21502,N_21067);
nand U21868 (N_21868,N_21462,N_21379);
or U21869 (N_21869,N_21598,N_21444);
or U21870 (N_21870,N_21021,N_21574);
nand U21871 (N_21871,N_21010,N_21020);
or U21872 (N_21872,N_21253,N_21071);
and U21873 (N_21873,N_21204,N_21143);
nor U21874 (N_21874,N_21332,N_21398);
or U21875 (N_21875,N_21284,N_21583);
nor U21876 (N_21876,N_21424,N_21546);
xnor U21877 (N_21877,N_21522,N_21447);
or U21878 (N_21878,N_21130,N_21311);
and U21879 (N_21879,N_21254,N_21320);
or U21880 (N_21880,N_21196,N_21318);
nor U21881 (N_21881,N_21263,N_21578);
or U21882 (N_21882,N_21230,N_21090);
or U21883 (N_21883,N_21448,N_21037);
or U21884 (N_21884,N_21217,N_21427);
nand U21885 (N_21885,N_21545,N_21344);
or U21886 (N_21886,N_21202,N_21415);
nor U21887 (N_21887,N_21493,N_21498);
and U21888 (N_21888,N_21001,N_21058);
nand U21889 (N_21889,N_21019,N_21092);
nand U21890 (N_21890,N_21426,N_21280);
or U21891 (N_21891,N_21464,N_21080);
and U21892 (N_21892,N_21061,N_21389);
or U21893 (N_21893,N_21367,N_21491);
and U21894 (N_21894,N_21388,N_21207);
and U21895 (N_21895,N_21234,N_21150);
nand U21896 (N_21896,N_21248,N_21287);
or U21897 (N_21897,N_21547,N_21542);
or U21898 (N_21898,N_21205,N_21009);
or U21899 (N_21899,N_21413,N_21182);
or U21900 (N_21900,N_21597,N_21285);
nand U21901 (N_21901,N_21406,N_21540);
and U21902 (N_21902,N_21583,N_21372);
and U21903 (N_21903,N_21029,N_21239);
or U21904 (N_21904,N_21462,N_21132);
and U21905 (N_21905,N_21239,N_21383);
nor U21906 (N_21906,N_21455,N_21152);
nor U21907 (N_21907,N_21459,N_21524);
xor U21908 (N_21908,N_21030,N_21010);
or U21909 (N_21909,N_21549,N_21512);
and U21910 (N_21910,N_21142,N_21545);
or U21911 (N_21911,N_21330,N_21419);
or U21912 (N_21912,N_21444,N_21334);
and U21913 (N_21913,N_21319,N_21373);
or U21914 (N_21914,N_21328,N_21300);
and U21915 (N_21915,N_21574,N_21482);
or U21916 (N_21916,N_21435,N_21340);
and U21917 (N_21917,N_21236,N_21033);
and U21918 (N_21918,N_21003,N_21500);
or U21919 (N_21919,N_21218,N_21007);
and U21920 (N_21920,N_21305,N_21487);
nor U21921 (N_21921,N_21067,N_21252);
nand U21922 (N_21922,N_21263,N_21235);
nor U21923 (N_21923,N_21410,N_21209);
nor U21924 (N_21924,N_21546,N_21289);
nand U21925 (N_21925,N_21092,N_21188);
or U21926 (N_21926,N_21529,N_21005);
and U21927 (N_21927,N_21429,N_21359);
nor U21928 (N_21928,N_21363,N_21028);
nor U21929 (N_21929,N_21545,N_21051);
nand U21930 (N_21930,N_21498,N_21031);
nand U21931 (N_21931,N_21598,N_21184);
or U21932 (N_21932,N_21435,N_21421);
or U21933 (N_21933,N_21413,N_21119);
nor U21934 (N_21934,N_21113,N_21296);
or U21935 (N_21935,N_21249,N_21523);
and U21936 (N_21936,N_21312,N_21156);
and U21937 (N_21937,N_21050,N_21384);
nor U21938 (N_21938,N_21318,N_21467);
nor U21939 (N_21939,N_21106,N_21215);
nand U21940 (N_21940,N_21564,N_21469);
nor U21941 (N_21941,N_21529,N_21287);
and U21942 (N_21942,N_21485,N_21445);
or U21943 (N_21943,N_21525,N_21147);
and U21944 (N_21944,N_21580,N_21219);
nor U21945 (N_21945,N_21127,N_21440);
nand U21946 (N_21946,N_21195,N_21230);
and U21947 (N_21947,N_21424,N_21112);
and U21948 (N_21948,N_21405,N_21235);
or U21949 (N_21949,N_21088,N_21440);
nand U21950 (N_21950,N_21034,N_21260);
nor U21951 (N_21951,N_21443,N_21565);
and U21952 (N_21952,N_21563,N_21207);
nor U21953 (N_21953,N_21265,N_21309);
nor U21954 (N_21954,N_21468,N_21170);
nor U21955 (N_21955,N_21073,N_21598);
nand U21956 (N_21956,N_21552,N_21075);
or U21957 (N_21957,N_21237,N_21215);
xor U21958 (N_21958,N_21340,N_21406);
or U21959 (N_21959,N_21123,N_21474);
and U21960 (N_21960,N_21313,N_21124);
and U21961 (N_21961,N_21104,N_21208);
nor U21962 (N_21962,N_21598,N_21337);
nand U21963 (N_21963,N_21044,N_21119);
nand U21964 (N_21964,N_21170,N_21009);
nand U21965 (N_21965,N_21180,N_21406);
nor U21966 (N_21966,N_21392,N_21338);
or U21967 (N_21967,N_21097,N_21365);
nor U21968 (N_21968,N_21021,N_21334);
nand U21969 (N_21969,N_21375,N_21036);
or U21970 (N_21970,N_21198,N_21278);
xnor U21971 (N_21971,N_21159,N_21150);
or U21972 (N_21972,N_21147,N_21411);
nor U21973 (N_21973,N_21315,N_21050);
nand U21974 (N_21974,N_21194,N_21406);
or U21975 (N_21975,N_21176,N_21453);
or U21976 (N_21976,N_21048,N_21009);
and U21977 (N_21977,N_21485,N_21171);
and U21978 (N_21978,N_21300,N_21445);
nor U21979 (N_21979,N_21250,N_21141);
and U21980 (N_21980,N_21096,N_21365);
xor U21981 (N_21981,N_21561,N_21051);
and U21982 (N_21982,N_21012,N_21535);
nand U21983 (N_21983,N_21027,N_21510);
nor U21984 (N_21984,N_21121,N_21474);
or U21985 (N_21985,N_21421,N_21002);
and U21986 (N_21986,N_21267,N_21485);
or U21987 (N_21987,N_21288,N_21019);
nor U21988 (N_21988,N_21233,N_21006);
and U21989 (N_21989,N_21077,N_21402);
and U21990 (N_21990,N_21114,N_21101);
and U21991 (N_21991,N_21355,N_21069);
or U21992 (N_21992,N_21465,N_21338);
nand U21993 (N_21993,N_21386,N_21186);
nor U21994 (N_21994,N_21422,N_21123);
or U21995 (N_21995,N_21264,N_21533);
nor U21996 (N_21996,N_21476,N_21064);
and U21997 (N_21997,N_21427,N_21070);
nor U21998 (N_21998,N_21332,N_21267);
or U21999 (N_21999,N_21135,N_21491);
nand U22000 (N_22000,N_21571,N_21070);
xnor U22001 (N_22001,N_21512,N_21548);
nor U22002 (N_22002,N_21394,N_21013);
nand U22003 (N_22003,N_21189,N_21303);
nor U22004 (N_22004,N_21462,N_21529);
or U22005 (N_22005,N_21159,N_21372);
and U22006 (N_22006,N_21150,N_21187);
nand U22007 (N_22007,N_21036,N_21024);
nor U22008 (N_22008,N_21434,N_21554);
and U22009 (N_22009,N_21147,N_21474);
nor U22010 (N_22010,N_21204,N_21314);
nor U22011 (N_22011,N_21363,N_21343);
nor U22012 (N_22012,N_21176,N_21327);
nor U22013 (N_22013,N_21257,N_21098);
nand U22014 (N_22014,N_21165,N_21221);
or U22015 (N_22015,N_21142,N_21362);
or U22016 (N_22016,N_21161,N_21470);
nor U22017 (N_22017,N_21559,N_21070);
or U22018 (N_22018,N_21484,N_21209);
nand U22019 (N_22019,N_21594,N_21428);
and U22020 (N_22020,N_21024,N_21430);
nand U22021 (N_22021,N_21233,N_21535);
nor U22022 (N_22022,N_21526,N_21193);
or U22023 (N_22023,N_21564,N_21152);
nand U22024 (N_22024,N_21472,N_21408);
xnor U22025 (N_22025,N_21182,N_21586);
nor U22026 (N_22026,N_21292,N_21252);
nor U22027 (N_22027,N_21083,N_21226);
nand U22028 (N_22028,N_21478,N_21401);
nor U22029 (N_22029,N_21381,N_21020);
nand U22030 (N_22030,N_21137,N_21553);
and U22031 (N_22031,N_21103,N_21410);
nor U22032 (N_22032,N_21449,N_21072);
and U22033 (N_22033,N_21265,N_21371);
or U22034 (N_22034,N_21191,N_21159);
nand U22035 (N_22035,N_21247,N_21127);
nand U22036 (N_22036,N_21246,N_21507);
and U22037 (N_22037,N_21336,N_21134);
nand U22038 (N_22038,N_21559,N_21358);
nor U22039 (N_22039,N_21165,N_21235);
or U22040 (N_22040,N_21039,N_21584);
nand U22041 (N_22041,N_21114,N_21248);
nand U22042 (N_22042,N_21103,N_21098);
nor U22043 (N_22043,N_21271,N_21120);
and U22044 (N_22044,N_21372,N_21080);
and U22045 (N_22045,N_21221,N_21498);
or U22046 (N_22046,N_21367,N_21590);
or U22047 (N_22047,N_21142,N_21133);
or U22048 (N_22048,N_21452,N_21154);
or U22049 (N_22049,N_21146,N_21356);
and U22050 (N_22050,N_21342,N_21573);
nand U22051 (N_22051,N_21511,N_21521);
nor U22052 (N_22052,N_21220,N_21579);
nand U22053 (N_22053,N_21538,N_21539);
xor U22054 (N_22054,N_21207,N_21014);
nand U22055 (N_22055,N_21404,N_21462);
and U22056 (N_22056,N_21452,N_21430);
or U22057 (N_22057,N_21288,N_21533);
or U22058 (N_22058,N_21420,N_21598);
nor U22059 (N_22059,N_21083,N_21023);
and U22060 (N_22060,N_21161,N_21395);
nand U22061 (N_22061,N_21135,N_21363);
nand U22062 (N_22062,N_21070,N_21304);
nor U22063 (N_22063,N_21211,N_21220);
nor U22064 (N_22064,N_21383,N_21398);
nor U22065 (N_22065,N_21574,N_21596);
or U22066 (N_22066,N_21207,N_21127);
or U22067 (N_22067,N_21215,N_21208);
or U22068 (N_22068,N_21068,N_21410);
or U22069 (N_22069,N_21508,N_21164);
and U22070 (N_22070,N_21140,N_21510);
or U22071 (N_22071,N_21518,N_21018);
nor U22072 (N_22072,N_21403,N_21379);
nand U22073 (N_22073,N_21453,N_21443);
and U22074 (N_22074,N_21226,N_21383);
nor U22075 (N_22075,N_21040,N_21555);
and U22076 (N_22076,N_21142,N_21127);
nor U22077 (N_22077,N_21110,N_21286);
and U22078 (N_22078,N_21410,N_21378);
nand U22079 (N_22079,N_21490,N_21273);
nor U22080 (N_22080,N_21036,N_21560);
and U22081 (N_22081,N_21413,N_21106);
and U22082 (N_22082,N_21389,N_21451);
nand U22083 (N_22083,N_21016,N_21229);
or U22084 (N_22084,N_21377,N_21596);
and U22085 (N_22085,N_21123,N_21410);
and U22086 (N_22086,N_21495,N_21238);
nand U22087 (N_22087,N_21400,N_21291);
or U22088 (N_22088,N_21342,N_21218);
or U22089 (N_22089,N_21397,N_21129);
nor U22090 (N_22090,N_21076,N_21423);
or U22091 (N_22091,N_21164,N_21426);
or U22092 (N_22092,N_21497,N_21509);
or U22093 (N_22093,N_21486,N_21260);
nor U22094 (N_22094,N_21367,N_21513);
nand U22095 (N_22095,N_21163,N_21528);
or U22096 (N_22096,N_21067,N_21018);
nor U22097 (N_22097,N_21459,N_21413);
and U22098 (N_22098,N_21358,N_21528);
nor U22099 (N_22099,N_21588,N_21424);
or U22100 (N_22100,N_21421,N_21502);
nor U22101 (N_22101,N_21556,N_21195);
nand U22102 (N_22102,N_21383,N_21421);
and U22103 (N_22103,N_21569,N_21392);
nor U22104 (N_22104,N_21597,N_21072);
or U22105 (N_22105,N_21267,N_21442);
and U22106 (N_22106,N_21072,N_21328);
nand U22107 (N_22107,N_21459,N_21209);
nor U22108 (N_22108,N_21427,N_21315);
nor U22109 (N_22109,N_21509,N_21017);
xor U22110 (N_22110,N_21435,N_21459);
and U22111 (N_22111,N_21387,N_21096);
nor U22112 (N_22112,N_21387,N_21468);
nand U22113 (N_22113,N_21285,N_21425);
nand U22114 (N_22114,N_21248,N_21459);
nor U22115 (N_22115,N_21578,N_21274);
or U22116 (N_22116,N_21112,N_21193);
xor U22117 (N_22117,N_21468,N_21543);
xnor U22118 (N_22118,N_21326,N_21370);
nor U22119 (N_22119,N_21023,N_21411);
or U22120 (N_22120,N_21012,N_21372);
and U22121 (N_22121,N_21476,N_21247);
or U22122 (N_22122,N_21121,N_21091);
or U22123 (N_22123,N_21565,N_21596);
nand U22124 (N_22124,N_21300,N_21122);
and U22125 (N_22125,N_21550,N_21460);
nand U22126 (N_22126,N_21005,N_21197);
or U22127 (N_22127,N_21209,N_21211);
nor U22128 (N_22128,N_21319,N_21571);
or U22129 (N_22129,N_21586,N_21028);
nor U22130 (N_22130,N_21228,N_21427);
xor U22131 (N_22131,N_21354,N_21043);
or U22132 (N_22132,N_21561,N_21181);
nand U22133 (N_22133,N_21100,N_21233);
nand U22134 (N_22134,N_21426,N_21578);
and U22135 (N_22135,N_21477,N_21487);
and U22136 (N_22136,N_21084,N_21043);
nor U22137 (N_22137,N_21331,N_21419);
or U22138 (N_22138,N_21460,N_21137);
and U22139 (N_22139,N_21228,N_21288);
or U22140 (N_22140,N_21299,N_21206);
or U22141 (N_22141,N_21543,N_21008);
nand U22142 (N_22142,N_21411,N_21566);
and U22143 (N_22143,N_21043,N_21115);
or U22144 (N_22144,N_21108,N_21271);
and U22145 (N_22145,N_21545,N_21290);
and U22146 (N_22146,N_21373,N_21115);
nand U22147 (N_22147,N_21006,N_21556);
nand U22148 (N_22148,N_21379,N_21546);
or U22149 (N_22149,N_21035,N_21345);
and U22150 (N_22150,N_21087,N_21090);
nor U22151 (N_22151,N_21373,N_21503);
nand U22152 (N_22152,N_21448,N_21230);
nand U22153 (N_22153,N_21326,N_21084);
or U22154 (N_22154,N_21531,N_21285);
and U22155 (N_22155,N_21005,N_21582);
nand U22156 (N_22156,N_21438,N_21217);
and U22157 (N_22157,N_21474,N_21373);
and U22158 (N_22158,N_21405,N_21598);
nor U22159 (N_22159,N_21386,N_21445);
or U22160 (N_22160,N_21139,N_21190);
and U22161 (N_22161,N_21360,N_21317);
nor U22162 (N_22162,N_21231,N_21202);
and U22163 (N_22163,N_21441,N_21286);
nor U22164 (N_22164,N_21291,N_21490);
nor U22165 (N_22165,N_21535,N_21459);
or U22166 (N_22166,N_21290,N_21116);
or U22167 (N_22167,N_21491,N_21036);
nand U22168 (N_22168,N_21482,N_21408);
nand U22169 (N_22169,N_21525,N_21113);
nor U22170 (N_22170,N_21373,N_21104);
or U22171 (N_22171,N_21259,N_21360);
nor U22172 (N_22172,N_21314,N_21429);
nand U22173 (N_22173,N_21120,N_21194);
nor U22174 (N_22174,N_21135,N_21591);
nor U22175 (N_22175,N_21465,N_21591);
nand U22176 (N_22176,N_21384,N_21267);
and U22177 (N_22177,N_21343,N_21027);
or U22178 (N_22178,N_21365,N_21019);
or U22179 (N_22179,N_21391,N_21082);
nand U22180 (N_22180,N_21409,N_21045);
and U22181 (N_22181,N_21123,N_21395);
nor U22182 (N_22182,N_21274,N_21060);
and U22183 (N_22183,N_21141,N_21138);
and U22184 (N_22184,N_21201,N_21442);
nor U22185 (N_22185,N_21526,N_21410);
and U22186 (N_22186,N_21299,N_21534);
nand U22187 (N_22187,N_21574,N_21591);
and U22188 (N_22188,N_21215,N_21473);
nand U22189 (N_22189,N_21143,N_21173);
and U22190 (N_22190,N_21004,N_21095);
and U22191 (N_22191,N_21495,N_21360);
nand U22192 (N_22192,N_21558,N_21354);
or U22193 (N_22193,N_21514,N_21487);
or U22194 (N_22194,N_21289,N_21093);
nor U22195 (N_22195,N_21353,N_21062);
and U22196 (N_22196,N_21092,N_21121);
and U22197 (N_22197,N_21495,N_21166);
nor U22198 (N_22198,N_21041,N_21224);
or U22199 (N_22199,N_21061,N_21352);
nor U22200 (N_22200,N_22145,N_21838);
or U22201 (N_22201,N_21878,N_21609);
or U22202 (N_22202,N_22113,N_22169);
nand U22203 (N_22203,N_21905,N_21887);
and U22204 (N_22204,N_22108,N_22072);
and U22205 (N_22205,N_21890,N_22018);
nor U22206 (N_22206,N_22112,N_21603);
nor U22207 (N_22207,N_21825,N_22063);
or U22208 (N_22208,N_22051,N_21813);
nand U22209 (N_22209,N_22037,N_22118);
or U22210 (N_22210,N_21649,N_22167);
nand U22211 (N_22211,N_21952,N_21855);
or U22212 (N_22212,N_21894,N_21729);
and U22213 (N_22213,N_21832,N_21882);
or U22214 (N_22214,N_21973,N_21995);
or U22215 (N_22215,N_21921,N_21714);
nand U22216 (N_22216,N_21904,N_22001);
or U22217 (N_22217,N_21960,N_21760);
nand U22218 (N_22218,N_21869,N_21680);
nor U22219 (N_22219,N_22164,N_21764);
nand U22220 (N_22220,N_21705,N_21853);
and U22221 (N_22221,N_21840,N_22013);
xnor U22222 (N_22222,N_22146,N_21994);
nand U22223 (N_22223,N_21901,N_21648);
nor U22224 (N_22224,N_21713,N_21930);
or U22225 (N_22225,N_22186,N_21981);
nand U22226 (N_22226,N_21681,N_21924);
nor U22227 (N_22227,N_21629,N_21826);
nand U22228 (N_22228,N_21834,N_21993);
and U22229 (N_22229,N_22198,N_21966);
and U22230 (N_22230,N_22153,N_22010);
nor U22231 (N_22231,N_22110,N_21687);
nand U22232 (N_22232,N_21667,N_22193);
or U22233 (N_22233,N_21642,N_22129);
or U22234 (N_22234,N_21803,N_21636);
or U22235 (N_22235,N_22194,N_21935);
nor U22236 (N_22236,N_21639,N_21748);
nor U22237 (N_22237,N_21936,N_21659);
or U22238 (N_22238,N_22172,N_22178);
or U22239 (N_22239,N_21661,N_21922);
nor U22240 (N_22240,N_21925,N_21688);
xor U22241 (N_22241,N_22124,N_22041);
nor U22242 (N_22242,N_21669,N_21800);
nor U22243 (N_22243,N_22133,N_21982);
xor U22244 (N_22244,N_21738,N_22103);
nor U22245 (N_22245,N_21690,N_22168);
and U22246 (N_22246,N_21926,N_21651);
or U22247 (N_22247,N_21739,N_22002);
nor U22248 (N_22248,N_22105,N_21616);
nand U22249 (N_22249,N_21785,N_22029);
or U22250 (N_22250,N_21723,N_22137);
nor U22251 (N_22251,N_21843,N_21810);
or U22252 (N_22252,N_21902,N_21865);
nor U22253 (N_22253,N_22014,N_21691);
nor U22254 (N_22254,N_22050,N_22141);
nor U22255 (N_22255,N_22114,N_21766);
nand U22256 (N_22256,N_21816,N_21671);
nor U22257 (N_22257,N_22087,N_22082);
nand U22258 (N_22258,N_21913,N_21716);
nand U22259 (N_22259,N_21818,N_21980);
and U22260 (N_22260,N_22158,N_22045);
and U22261 (N_22261,N_22068,N_21678);
nor U22262 (N_22262,N_21910,N_22101);
nor U22263 (N_22263,N_21896,N_21961);
nand U22264 (N_22264,N_21806,N_21941);
or U22265 (N_22265,N_21954,N_21815);
nor U22266 (N_22266,N_21842,N_22192);
or U22267 (N_22267,N_21916,N_21797);
nor U22268 (N_22268,N_21807,N_21751);
nand U22269 (N_22269,N_22174,N_21617);
or U22270 (N_22270,N_22119,N_21854);
nand U22271 (N_22271,N_21889,N_22017);
nor U22272 (N_22272,N_22085,N_21725);
xor U22273 (N_22273,N_21728,N_21884);
nand U22274 (N_22274,N_21976,N_21962);
and U22275 (N_22275,N_21695,N_21817);
or U22276 (N_22276,N_21822,N_21864);
nor U22277 (N_22277,N_21903,N_21731);
and U22278 (N_22278,N_21875,N_22044);
nor U22279 (N_22279,N_21770,N_22161);
nand U22280 (N_22280,N_21602,N_22032);
and U22281 (N_22281,N_22100,N_21844);
nand U22282 (N_22282,N_22154,N_21915);
or U22283 (N_22283,N_21786,N_21963);
nor U22284 (N_22284,N_22189,N_21634);
or U22285 (N_22285,N_21654,N_22058);
or U22286 (N_22286,N_21622,N_22175);
nor U22287 (N_22287,N_21612,N_22173);
xnor U22288 (N_22288,N_21771,N_21735);
and U22289 (N_22289,N_21969,N_21992);
xnor U22290 (N_22290,N_21758,N_21920);
nand U22291 (N_22291,N_22182,N_21666);
or U22292 (N_22292,N_22000,N_21988);
nand U22293 (N_22293,N_22030,N_21808);
nor U22294 (N_22294,N_21945,N_21638);
nor U22295 (N_22295,N_21633,N_22084);
nor U22296 (N_22296,N_22109,N_21620);
nor U22297 (N_22297,N_21676,N_21944);
or U22298 (N_22298,N_21823,N_22092);
or U22299 (N_22299,N_21759,N_22107);
or U22300 (N_22300,N_21950,N_22160);
nand U22301 (N_22301,N_21958,N_21977);
nor U22302 (N_22302,N_21707,N_21917);
nand U22303 (N_22303,N_22055,N_21900);
nand U22304 (N_22304,N_21720,N_22008);
nand U22305 (N_22305,N_21856,N_21778);
or U22306 (N_22306,N_22156,N_21641);
or U22307 (N_22307,N_21814,N_21604);
or U22308 (N_22308,N_21971,N_22023);
or U22309 (N_22309,N_21697,N_21608);
nand U22310 (N_22310,N_21722,N_21835);
or U22311 (N_22311,N_21883,N_21805);
nor U22312 (N_22312,N_21677,N_22006);
or U22313 (N_22313,N_21983,N_21628);
and U22314 (N_22314,N_21940,N_22170);
and U22315 (N_22315,N_21712,N_21951);
and U22316 (N_22316,N_21696,N_21744);
or U22317 (N_22317,N_21837,N_22197);
or U22318 (N_22318,N_21607,N_21821);
nand U22319 (N_22319,N_21702,N_22056);
or U22320 (N_22320,N_22039,N_22117);
nor U22321 (N_22321,N_22021,N_21750);
nor U22322 (N_22322,N_22040,N_21999);
nand U22323 (N_22323,N_21779,N_21600);
nor U22324 (N_22324,N_21955,N_22116);
or U22325 (N_22325,N_21730,N_22093);
nor U22326 (N_22326,N_22122,N_21879);
nor U22327 (N_22327,N_21857,N_22185);
nor U22328 (N_22328,N_21601,N_22150);
and U22329 (N_22329,N_21749,N_21726);
nand U22330 (N_22330,N_21895,N_22005);
and U22331 (N_22331,N_21717,N_21610);
and U22332 (N_22332,N_22131,N_21605);
nand U22333 (N_22333,N_22078,N_21784);
nor U22334 (N_22334,N_21799,N_21798);
and U22335 (N_22335,N_22049,N_21847);
nand U22336 (N_22336,N_21942,N_22195);
or U22337 (N_22337,N_22076,N_21701);
and U22338 (N_22338,N_21790,N_21984);
xnor U22339 (N_22339,N_21754,N_22035);
nand U22340 (N_22340,N_21795,N_22097);
nor U22341 (N_22341,N_22069,N_21820);
nor U22342 (N_22342,N_21987,N_21665);
nand U22343 (N_22343,N_22057,N_21861);
nand U22344 (N_22344,N_22152,N_22019);
and U22345 (N_22345,N_22099,N_22083);
and U22346 (N_22346,N_22139,N_21774);
nand U22347 (N_22347,N_21783,N_21689);
and U22348 (N_22348,N_21970,N_21899);
or U22349 (N_22349,N_21753,N_21793);
or U22350 (N_22350,N_21929,N_21870);
or U22351 (N_22351,N_22136,N_22180);
nor U22352 (N_22352,N_21827,N_21640);
nor U22353 (N_22353,N_21836,N_21703);
nor U22354 (N_22354,N_21830,N_21625);
nor U22355 (N_22355,N_21668,N_21775);
nand U22356 (N_22356,N_21781,N_22098);
nand U22357 (N_22357,N_21989,N_21611);
nand U22358 (N_22358,N_21692,N_21646);
xnor U22359 (N_22359,N_21907,N_21788);
nor U22360 (N_22360,N_22071,N_21831);
nand U22361 (N_22361,N_22015,N_22187);
nand U22362 (N_22362,N_21968,N_21979);
nand U22363 (N_22363,N_22090,N_21630);
nand U22364 (N_22364,N_22003,N_21967);
nand U22365 (N_22365,N_22179,N_22148);
nor U22366 (N_22366,N_22053,N_22196);
or U22367 (N_22367,N_21755,N_22096);
nand U22368 (N_22368,N_21886,N_22134);
or U22369 (N_22369,N_21972,N_21909);
or U22370 (N_22370,N_21621,N_21647);
or U22371 (N_22371,N_21746,N_21672);
or U22372 (N_22372,N_21943,N_21663);
and U22373 (N_22373,N_21732,N_21736);
or U22374 (N_22374,N_21923,N_21897);
or U22375 (N_22375,N_21711,N_21845);
xor U22376 (N_22376,N_21655,N_22086);
or U22377 (N_22377,N_21933,N_22126);
and U22378 (N_22378,N_21947,N_21829);
nor U22379 (N_22379,N_21719,N_21777);
nand U22380 (N_22380,N_21762,N_21990);
nand U22381 (N_22381,N_22162,N_22125);
or U22382 (N_22382,N_22091,N_21776);
nor U22383 (N_22383,N_22159,N_21998);
or U22384 (N_22384,N_22038,N_21975);
nor U22385 (N_22385,N_21794,N_21811);
nand U22386 (N_22386,N_21848,N_22166);
nor U22387 (N_22387,N_22052,N_21938);
or U22388 (N_22388,N_22144,N_21700);
or U22389 (N_22389,N_22027,N_21957);
nor U22390 (N_22390,N_21733,N_22054);
and U22391 (N_22391,N_21740,N_22048);
nand U22392 (N_22392,N_21839,N_22127);
nand U22393 (N_22393,N_22181,N_22011);
and U22394 (N_22394,N_22188,N_22157);
and U22395 (N_22395,N_21849,N_22075);
nor U22396 (N_22396,N_21708,N_21657);
and U22397 (N_22397,N_21615,N_22081);
nand U22398 (N_22398,N_22183,N_21862);
and U22399 (N_22399,N_21769,N_21768);
and U22400 (N_22400,N_21670,N_22177);
xor U22401 (N_22401,N_21928,N_21694);
nand U22402 (N_22402,N_21888,N_21743);
nand U22403 (N_22403,N_21693,N_21635);
nor U22404 (N_22404,N_21812,N_21792);
nor U22405 (N_22405,N_22009,N_21898);
xor U22406 (N_22406,N_21757,N_21637);
or U22407 (N_22407,N_21685,N_22088);
and U22408 (N_22408,N_21906,N_22142);
and U22409 (N_22409,N_21802,N_21965);
and U22410 (N_22410,N_21787,N_22059);
and U22411 (N_22411,N_22079,N_22120);
nor U22412 (N_22412,N_21846,N_21718);
nor U22413 (N_22413,N_22065,N_21644);
nor U22414 (N_22414,N_21664,N_21643);
nand U22415 (N_22415,N_22024,N_21946);
or U22416 (N_22416,N_21858,N_22151);
or U22417 (N_22417,N_21885,N_22012);
nor U22418 (N_22418,N_21745,N_21978);
or U22419 (N_22419,N_21618,N_21780);
nor U22420 (N_22420,N_22080,N_21804);
nor U22421 (N_22421,N_22064,N_21741);
xor U22422 (N_22422,N_22191,N_22016);
nor U22423 (N_22423,N_22140,N_22089);
nor U22424 (N_22424,N_21833,N_21852);
or U22425 (N_22425,N_22025,N_21704);
or U22426 (N_22426,N_22135,N_21653);
nand U22427 (N_22427,N_22165,N_21863);
and U22428 (N_22428,N_22073,N_21860);
nor U22429 (N_22429,N_21809,N_21721);
nor U22430 (N_22430,N_21819,N_21715);
nand U22431 (N_22431,N_21912,N_22077);
and U22432 (N_22432,N_22007,N_21660);
nor U22433 (N_22433,N_21656,N_21986);
and U22434 (N_22434,N_21828,N_21892);
nand U22435 (N_22435,N_21763,N_22066);
nand U22436 (N_22436,N_21772,N_21619);
nor U22437 (N_22437,N_22070,N_21614);
or U22438 (N_22438,N_22095,N_21918);
and U22439 (N_22439,N_21752,N_21765);
and U22440 (N_22440,N_21937,N_21891);
nand U22441 (N_22441,N_22115,N_21871);
or U22442 (N_22442,N_21662,N_21796);
or U22443 (N_22443,N_21724,N_22163);
and U22444 (N_22444,N_21841,N_21626);
or U22445 (N_22445,N_22033,N_21674);
nor U22446 (N_22446,N_21908,N_22043);
nor U22447 (N_22447,N_21881,N_21956);
nor U22448 (N_22448,N_21706,N_21756);
and U22449 (N_22449,N_21872,N_22121);
nand U22450 (N_22450,N_21868,N_22046);
xnor U22451 (N_22451,N_21613,N_22111);
or U22452 (N_22452,N_21632,N_21791);
xnor U22453 (N_22453,N_21919,N_22061);
or U22454 (N_22454,N_22042,N_22036);
nand U22455 (N_22455,N_22138,N_21876);
nand U22456 (N_22456,N_21710,N_21734);
and U22457 (N_22457,N_21737,N_21880);
nand U22458 (N_22458,N_22123,N_22104);
and U22459 (N_22459,N_21985,N_22004);
and U22460 (N_22460,N_21974,N_21699);
or U22461 (N_22461,N_22130,N_21873);
nand U22462 (N_22462,N_22176,N_22102);
and U22463 (N_22463,N_21658,N_21773);
and U22464 (N_22464,N_22149,N_21824);
or U22465 (N_22465,N_22143,N_21934);
nor U22466 (N_22466,N_21727,N_21948);
nand U22467 (N_22467,N_21709,N_21742);
nor U22468 (N_22468,N_21997,N_21682);
and U22469 (N_22469,N_21866,N_22034);
and U22470 (N_22470,N_22022,N_22132);
nand U22471 (N_22471,N_22047,N_21675);
or U22472 (N_22472,N_21927,N_22155);
nor U22473 (N_22473,N_21673,N_22128);
nand U22474 (N_22474,N_21911,N_21874);
nand U22475 (N_22475,N_21683,N_22074);
or U22476 (N_22476,N_21996,N_22184);
or U22477 (N_22477,N_21624,N_21949);
or U22478 (N_22478,N_22067,N_21686);
or U22479 (N_22479,N_21914,N_22020);
nand U22480 (N_22480,N_21939,N_21850);
nand U22481 (N_22481,N_22147,N_21991);
or U22482 (N_22482,N_22026,N_21867);
nand U22483 (N_22483,N_21684,N_21761);
nor U22484 (N_22484,N_21623,N_22106);
nand U22485 (N_22485,N_21859,N_21893);
nor U22486 (N_22486,N_21964,N_21953);
or U22487 (N_22487,N_21932,N_21801);
nor U22488 (N_22488,N_21652,N_21679);
and U22489 (N_22489,N_21606,N_21631);
or U22490 (N_22490,N_21782,N_21627);
or U22491 (N_22491,N_21789,N_21698);
and U22492 (N_22492,N_22031,N_22028);
or U22493 (N_22493,N_21877,N_22094);
or U22494 (N_22494,N_22062,N_22190);
nor U22495 (N_22495,N_22171,N_21959);
xnor U22496 (N_22496,N_22199,N_21645);
or U22497 (N_22497,N_22060,N_21851);
nor U22498 (N_22498,N_21931,N_21767);
nand U22499 (N_22499,N_21747,N_21650);
and U22500 (N_22500,N_22012,N_21982);
or U22501 (N_22501,N_21794,N_21626);
nand U22502 (N_22502,N_21773,N_21860);
nand U22503 (N_22503,N_21700,N_21876);
and U22504 (N_22504,N_21945,N_21840);
nand U22505 (N_22505,N_21843,N_22176);
or U22506 (N_22506,N_21899,N_21806);
nand U22507 (N_22507,N_22020,N_21840);
and U22508 (N_22508,N_21706,N_21788);
and U22509 (N_22509,N_21798,N_21691);
and U22510 (N_22510,N_22137,N_21765);
nor U22511 (N_22511,N_21914,N_22164);
or U22512 (N_22512,N_22098,N_22129);
or U22513 (N_22513,N_21698,N_21704);
nand U22514 (N_22514,N_22074,N_22072);
or U22515 (N_22515,N_21697,N_21829);
and U22516 (N_22516,N_21829,N_21717);
nand U22517 (N_22517,N_22054,N_21614);
nand U22518 (N_22518,N_21780,N_21792);
nand U22519 (N_22519,N_22023,N_21858);
or U22520 (N_22520,N_21818,N_21853);
and U22521 (N_22521,N_21850,N_21975);
or U22522 (N_22522,N_22004,N_21825);
nand U22523 (N_22523,N_21682,N_22198);
and U22524 (N_22524,N_21661,N_21869);
nand U22525 (N_22525,N_22178,N_21791);
or U22526 (N_22526,N_21670,N_21793);
nand U22527 (N_22527,N_22025,N_21962);
nand U22528 (N_22528,N_21611,N_22085);
nand U22529 (N_22529,N_21749,N_21969);
nor U22530 (N_22530,N_21917,N_22165);
nor U22531 (N_22531,N_21925,N_21799);
xor U22532 (N_22532,N_22108,N_22037);
nor U22533 (N_22533,N_22049,N_21815);
or U22534 (N_22534,N_21744,N_21896);
xor U22535 (N_22535,N_21950,N_22152);
or U22536 (N_22536,N_22140,N_21722);
nor U22537 (N_22537,N_21980,N_21736);
or U22538 (N_22538,N_21621,N_22074);
nor U22539 (N_22539,N_21912,N_22087);
xor U22540 (N_22540,N_22065,N_21687);
and U22541 (N_22541,N_21723,N_21809);
or U22542 (N_22542,N_22140,N_21817);
nor U22543 (N_22543,N_21830,N_22108);
or U22544 (N_22544,N_21996,N_21951);
nand U22545 (N_22545,N_21984,N_22154);
nand U22546 (N_22546,N_21980,N_22117);
nand U22547 (N_22547,N_22069,N_22102);
and U22548 (N_22548,N_21780,N_21829);
or U22549 (N_22549,N_22057,N_21973);
and U22550 (N_22550,N_21726,N_21877);
nor U22551 (N_22551,N_21643,N_21955);
nor U22552 (N_22552,N_21606,N_21904);
nor U22553 (N_22553,N_21924,N_21726);
nand U22554 (N_22554,N_21956,N_21708);
and U22555 (N_22555,N_22071,N_21755);
or U22556 (N_22556,N_22003,N_22084);
nor U22557 (N_22557,N_22094,N_21603);
and U22558 (N_22558,N_21912,N_22049);
or U22559 (N_22559,N_21796,N_21984);
or U22560 (N_22560,N_21876,N_21882);
and U22561 (N_22561,N_22086,N_22109);
or U22562 (N_22562,N_21690,N_22080);
nor U22563 (N_22563,N_22038,N_22051);
nor U22564 (N_22564,N_21746,N_21654);
and U22565 (N_22565,N_21798,N_22021);
and U22566 (N_22566,N_22001,N_21983);
and U22567 (N_22567,N_21694,N_21828);
or U22568 (N_22568,N_22169,N_21827);
nand U22569 (N_22569,N_22119,N_22149);
or U22570 (N_22570,N_21771,N_22043);
and U22571 (N_22571,N_21816,N_21892);
nand U22572 (N_22572,N_21654,N_21668);
or U22573 (N_22573,N_22030,N_21655);
nor U22574 (N_22574,N_22115,N_21962);
nand U22575 (N_22575,N_21629,N_21718);
nor U22576 (N_22576,N_21892,N_21749);
and U22577 (N_22577,N_21867,N_22169);
nor U22578 (N_22578,N_22191,N_21628);
or U22579 (N_22579,N_21655,N_21801);
nand U22580 (N_22580,N_21877,N_21601);
xor U22581 (N_22581,N_21647,N_22178);
and U22582 (N_22582,N_21610,N_21719);
nand U22583 (N_22583,N_21748,N_21656);
nor U22584 (N_22584,N_21865,N_21745);
and U22585 (N_22585,N_22013,N_21816);
xor U22586 (N_22586,N_22046,N_22076);
and U22587 (N_22587,N_21711,N_22109);
or U22588 (N_22588,N_21646,N_22027);
nor U22589 (N_22589,N_22115,N_21954);
nor U22590 (N_22590,N_22123,N_21734);
nor U22591 (N_22591,N_21932,N_21854);
nand U22592 (N_22592,N_21992,N_21918);
nor U22593 (N_22593,N_22005,N_21699);
or U22594 (N_22594,N_22108,N_21836);
nor U22595 (N_22595,N_21844,N_22003);
and U22596 (N_22596,N_21868,N_21720);
nor U22597 (N_22597,N_22008,N_21827);
nor U22598 (N_22598,N_21810,N_21884);
nor U22599 (N_22599,N_22008,N_21796);
and U22600 (N_22600,N_21896,N_21909);
or U22601 (N_22601,N_21901,N_21915);
or U22602 (N_22602,N_21835,N_21619);
nor U22603 (N_22603,N_21792,N_21864);
nand U22604 (N_22604,N_21700,N_22022);
or U22605 (N_22605,N_21917,N_21900);
nor U22606 (N_22606,N_21869,N_21677);
nand U22607 (N_22607,N_21629,N_21980);
and U22608 (N_22608,N_21675,N_22015);
nand U22609 (N_22609,N_21741,N_21930);
nor U22610 (N_22610,N_21898,N_21656);
and U22611 (N_22611,N_21868,N_22112);
and U22612 (N_22612,N_21998,N_22107);
xnor U22613 (N_22613,N_22142,N_22085);
nor U22614 (N_22614,N_21988,N_21876);
or U22615 (N_22615,N_22183,N_21897);
and U22616 (N_22616,N_21844,N_21616);
nor U22617 (N_22617,N_22042,N_21997);
nand U22618 (N_22618,N_22154,N_21636);
nand U22619 (N_22619,N_22118,N_22116);
and U22620 (N_22620,N_22079,N_21769);
and U22621 (N_22621,N_22178,N_21760);
nand U22622 (N_22622,N_21624,N_21787);
and U22623 (N_22623,N_22009,N_22086);
or U22624 (N_22624,N_21607,N_22132);
or U22625 (N_22625,N_21906,N_21983);
and U22626 (N_22626,N_22120,N_22174);
nand U22627 (N_22627,N_21658,N_21872);
or U22628 (N_22628,N_22148,N_21985);
and U22629 (N_22629,N_22194,N_22158);
or U22630 (N_22630,N_22118,N_21941);
nor U22631 (N_22631,N_21687,N_21912);
nor U22632 (N_22632,N_21954,N_21854);
nand U22633 (N_22633,N_21666,N_21834);
nand U22634 (N_22634,N_22043,N_21819);
and U22635 (N_22635,N_21663,N_21802);
or U22636 (N_22636,N_22091,N_21648);
or U22637 (N_22637,N_21774,N_22031);
xor U22638 (N_22638,N_21963,N_21741);
nand U22639 (N_22639,N_21600,N_21843);
or U22640 (N_22640,N_22182,N_21747);
and U22641 (N_22641,N_21812,N_21747);
nor U22642 (N_22642,N_21613,N_21890);
or U22643 (N_22643,N_21617,N_22054);
nor U22644 (N_22644,N_21831,N_22048);
or U22645 (N_22645,N_21973,N_22041);
nor U22646 (N_22646,N_22155,N_21706);
or U22647 (N_22647,N_21966,N_21612);
and U22648 (N_22648,N_21901,N_22013);
nand U22649 (N_22649,N_21913,N_21873);
nand U22650 (N_22650,N_22160,N_21736);
and U22651 (N_22651,N_22195,N_22101);
or U22652 (N_22652,N_21642,N_21740);
nor U22653 (N_22653,N_21978,N_22017);
nand U22654 (N_22654,N_21986,N_21893);
nor U22655 (N_22655,N_22081,N_21645);
nand U22656 (N_22656,N_21699,N_21737);
and U22657 (N_22657,N_21814,N_22190);
nor U22658 (N_22658,N_21823,N_21878);
nor U22659 (N_22659,N_22122,N_22001);
nor U22660 (N_22660,N_21695,N_21770);
and U22661 (N_22661,N_21953,N_22158);
nor U22662 (N_22662,N_22137,N_21770);
or U22663 (N_22663,N_21671,N_22070);
nor U22664 (N_22664,N_21631,N_21650);
nand U22665 (N_22665,N_21722,N_22134);
or U22666 (N_22666,N_22017,N_21904);
and U22667 (N_22667,N_22051,N_22112);
nor U22668 (N_22668,N_21717,N_22164);
and U22669 (N_22669,N_22081,N_22102);
nor U22670 (N_22670,N_21662,N_21848);
nor U22671 (N_22671,N_21872,N_21738);
xnor U22672 (N_22672,N_22097,N_22000);
nand U22673 (N_22673,N_21893,N_21926);
nand U22674 (N_22674,N_22176,N_21921);
and U22675 (N_22675,N_21823,N_21694);
nand U22676 (N_22676,N_21814,N_21897);
xnor U22677 (N_22677,N_21912,N_21788);
nor U22678 (N_22678,N_21609,N_22092);
nor U22679 (N_22679,N_21897,N_22152);
nand U22680 (N_22680,N_22093,N_21694);
or U22681 (N_22681,N_22089,N_22065);
and U22682 (N_22682,N_22045,N_21804);
nor U22683 (N_22683,N_21679,N_22161);
or U22684 (N_22684,N_21907,N_21944);
or U22685 (N_22685,N_22041,N_21999);
nand U22686 (N_22686,N_21761,N_21773);
nand U22687 (N_22687,N_21938,N_22121);
nand U22688 (N_22688,N_21679,N_22151);
nand U22689 (N_22689,N_21856,N_21730);
nor U22690 (N_22690,N_22024,N_21941);
or U22691 (N_22691,N_22052,N_22161);
or U22692 (N_22692,N_21888,N_21622);
and U22693 (N_22693,N_21928,N_21841);
and U22694 (N_22694,N_22065,N_21963);
nand U22695 (N_22695,N_21876,N_22032);
nor U22696 (N_22696,N_21637,N_21860);
nand U22697 (N_22697,N_21957,N_21940);
or U22698 (N_22698,N_22153,N_22125);
nand U22699 (N_22699,N_21834,N_21848);
or U22700 (N_22700,N_22073,N_22061);
or U22701 (N_22701,N_22034,N_21876);
nand U22702 (N_22702,N_21971,N_22001);
or U22703 (N_22703,N_21827,N_22150);
or U22704 (N_22704,N_21720,N_21997);
nand U22705 (N_22705,N_21817,N_21996);
nor U22706 (N_22706,N_21971,N_21600);
or U22707 (N_22707,N_21666,N_21810);
or U22708 (N_22708,N_22153,N_21686);
nor U22709 (N_22709,N_22113,N_21661);
nand U22710 (N_22710,N_21780,N_21748);
nor U22711 (N_22711,N_22016,N_21723);
or U22712 (N_22712,N_21879,N_21800);
and U22713 (N_22713,N_21732,N_21645);
nand U22714 (N_22714,N_22114,N_22017);
nand U22715 (N_22715,N_21712,N_22018);
nor U22716 (N_22716,N_21656,N_21800);
nand U22717 (N_22717,N_21713,N_21727);
nor U22718 (N_22718,N_22013,N_22019);
nor U22719 (N_22719,N_21821,N_21902);
nand U22720 (N_22720,N_21958,N_21851);
or U22721 (N_22721,N_22014,N_22134);
nor U22722 (N_22722,N_21998,N_22147);
nor U22723 (N_22723,N_21739,N_21978);
nor U22724 (N_22724,N_21789,N_21845);
nand U22725 (N_22725,N_22098,N_22144);
and U22726 (N_22726,N_22120,N_21847);
nor U22727 (N_22727,N_21769,N_22187);
nor U22728 (N_22728,N_21788,N_22127);
or U22729 (N_22729,N_21894,N_22089);
or U22730 (N_22730,N_21931,N_21612);
nor U22731 (N_22731,N_21900,N_22143);
and U22732 (N_22732,N_22100,N_22029);
and U22733 (N_22733,N_22037,N_21852);
or U22734 (N_22734,N_21793,N_21981);
nor U22735 (N_22735,N_21791,N_21674);
and U22736 (N_22736,N_21778,N_21984);
or U22737 (N_22737,N_21739,N_21934);
nor U22738 (N_22738,N_21618,N_21849);
nand U22739 (N_22739,N_21636,N_21931);
or U22740 (N_22740,N_21702,N_21745);
or U22741 (N_22741,N_21737,N_21611);
nor U22742 (N_22742,N_21984,N_22009);
nor U22743 (N_22743,N_22013,N_21874);
or U22744 (N_22744,N_22094,N_21907);
or U22745 (N_22745,N_22000,N_21789);
nand U22746 (N_22746,N_22104,N_21755);
or U22747 (N_22747,N_21818,N_22119);
or U22748 (N_22748,N_21803,N_21877);
and U22749 (N_22749,N_22134,N_22160);
and U22750 (N_22750,N_22014,N_21812);
nand U22751 (N_22751,N_22001,N_21651);
nor U22752 (N_22752,N_22174,N_21913);
nand U22753 (N_22753,N_22039,N_21605);
nor U22754 (N_22754,N_21943,N_21959);
nand U22755 (N_22755,N_21790,N_22159);
xnor U22756 (N_22756,N_21942,N_22069);
and U22757 (N_22757,N_21713,N_22043);
and U22758 (N_22758,N_21943,N_21973);
nor U22759 (N_22759,N_22068,N_21775);
nand U22760 (N_22760,N_21722,N_21630);
nand U22761 (N_22761,N_21835,N_21979);
and U22762 (N_22762,N_22190,N_21680);
and U22763 (N_22763,N_21894,N_22101);
and U22764 (N_22764,N_22134,N_22147);
nor U22765 (N_22765,N_21805,N_22015);
and U22766 (N_22766,N_22172,N_22064);
nand U22767 (N_22767,N_21829,N_22188);
or U22768 (N_22768,N_21837,N_21625);
or U22769 (N_22769,N_22143,N_22090);
nor U22770 (N_22770,N_21971,N_21910);
nand U22771 (N_22771,N_22090,N_21702);
nand U22772 (N_22772,N_21615,N_21964);
or U22773 (N_22773,N_22171,N_21741);
nand U22774 (N_22774,N_22062,N_21958);
nand U22775 (N_22775,N_22052,N_21668);
and U22776 (N_22776,N_21727,N_22182);
or U22777 (N_22777,N_21625,N_22092);
or U22778 (N_22778,N_21892,N_21671);
and U22779 (N_22779,N_21898,N_22146);
and U22780 (N_22780,N_21621,N_21968);
and U22781 (N_22781,N_21918,N_21621);
and U22782 (N_22782,N_21887,N_22064);
nand U22783 (N_22783,N_21706,N_21760);
nand U22784 (N_22784,N_22134,N_21795);
or U22785 (N_22785,N_21840,N_21939);
or U22786 (N_22786,N_21911,N_22015);
or U22787 (N_22787,N_21813,N_22030);
or U22788 (N_22788,N_22116,N_21957);
nand U22789 (N_22789,N_22002,N_22128);
nor U22790 (N_22790,N_22185,N_21628);
nor U22791 (N_22791,N_22025,N_21679);
and U22792 (N_22792,N_21682,N_21921);
and U22793 (N_22793,N_22092,N_21989);
nand U22794 (N_22794,N_22054,N_21811);
nand U22795 (N_22795,N_21906,N_21643);
nor U22796 (N_22796,N_21966,N_21601);
or U22797 (N_22797,N_21932,N_21878);
nor U22798 (N_22798,N_21766,N_21845);
nand U22799 (N_22799,N_22110,N_21716);
or U22800 (N_22800,N_22668,N_22418);
nand U22801 (N_22801,N_22308,N_22493);
nor U22802 (N_22802,N_22249,N_22798);
xor U22803 (N_22803,N_22456,N_22565);
nand U22804 (N_22804,N_22662,N_22378);
or U22805 (N_22805,N_22209,N_22555);
nand U22806 (N_22806,N_22789,N_22245);
nand U22807 (N_22807,N_22707,N_22517);
or U22808 (N_22808,N_22415,N_22756);
nor U22809 (N_22809,N_22568,N_22763);
nor U22810 (N_22810,N_22506,N_22320);
nor U22811 (N_22811,N_22566,N_22206);
nand U22812 (N_22812,N_22236,N_22533);
nand U22813 (N_22813,N_22760,N_22422);
nand U22814 (N_22814,N_22612,N_22451);
or U22815 (N_22815,N_22325,N_22393);
or U22816 (N_22816,N_22289,N_22223);
and U22817 (N_22817,N_22504,N_22375);
nand U22818 (N_22818,N_22297,N_22480);
nand U22819 (N_22819,N_22688,N_22498);
or U22820 (N_22820,N_22695,N_22720);
nand U22821 (N_22821,N_22277,N_22674);
and U22822 (N_22822,N_22401,N_22483);
nor U22823 (N_22823,N_22344,N_22270);
xor U22824 (N_22824,N_22491,N_22341);
or U22825 (N_22825,N_22439,N_22347);
xor U22826 (N_22826,N_22680,N_22352);
and U22827 (N_22827,N_22266,N_22602);
or U22828 (N_22828,N_22716,N_22471);
nand U22829 (N_22829,N_22294,N_22449);
nand U22830 (N_22830,N_22564,N_22637);
nor U22831 (N_22831,N_22241,N_22601);
nor U22832 (N_22832,N_22587,N_22200);
nand U22833 (N_22833,N_22394,N_22560);
or U22834 (N_22834,N_22364,N_22424);
and U22835 (N_22835,N_22461,N_22397);
nand U22836 (N_22836,N_22321,N_22793);
nand U22837 (N_22837,N_22543,N_22252);
or U22838 (N_22838,N_22784,N_22381);
xor U22839 (N_22839,N_22492,N_22304);
or U22840 (N_22840,N_22311,N_22474);
and U22841 (N_22841,N_22448,N_22272);
nand U22842 (N_22842,N_22232,N_22282);
or U22843 (N_22843,N_22728,N_22257);
nor U22844 (N_22844,N_22512,N_22616);
nand U22845 (N_22845,N_22576,N_22554);
nor U22846 (N_22846,N_22453,N_22500);
nand U22847 (N_22847,N_22284,N_22351);
nor U22848 (N_22848,N_22508,N_22408);
or U22849 (N_22849,N_22589,N_22704);
nor U22850 (N_22850,N_22534,N_22787);
and U22851 (N_22851,N_22698,N_22332);
or U22852 (N_22852,N_22753,N_22356);
or U22853 (N_22853,N_22440,N_22268);
nand U22854 (N_22854,N_22211,N_22447);
xor U22855 (N_22855,N_22590,N_22628);
nor U22856 (N_22856,N_22363,N_22340);
xnor U22857 (N_22857,N_22313,N_22201);
nand U22858 (N_22858,N_22339,N_22629);
or U22859 (N_22859,N_22573,N_22202);
nor U22860 (N_22860,N_22791,N_22694);
nand U22861 (N_22861,N_22368,N_22567);
or U22862 (N_22862,N_22464,N_22608);
nor U22863 (N_22863,N_22444,N_22317);
nor U22864 (N_22864,N_22389,N_22306);
nor U22865 (N_22865,N_22288,N_22656);
nor U22866 (N_22866,N_22583,N_22499);
nor U22867 (N_22867,N_22640,N_22652);
and U22868 (N_22868,N_22614,N_22705);
and U22869 (N_22869,N_22692,N_22213);
nand U22870 (N_22870,N_22666,N_22349);
nand U22871 (N_22871,N_22273,N_22469);
nor U22872 (N_22872,N_22665,N_22334);
nor U22873 (N_22873,N_22786,N_22595);
nor U22874 (N_22874,N_22617,N_22519);
or U22875 (N_22875,N_22767,N_22434);
or U22876 (N_22876,N_22669,N_22632);
and U22877 (N_22877,N_22501,N_22598);
nor U22878 (N_22878,N_22230,N_22515);
or U22879 (N_22879,N_22354,N_22623);
nand U22880 (N_22880,N_22660,N_22396);
nand U22881 (N_22881,N_22714,N_22719);
nand U22882 (N_22882,N_22400,N_22721);
and U22883 (N_22883,N_22635,N_22205);
and U22884 (N_22884,N_22369,N_22412);
xnor U22885 (N_22885,N_22234,N_22675);
xor U22886 (N_22886,N_22409,N_22299);
nand U22887 (N_22887,N_22641,N_22718);
nand U22888 (N_22888,N_22677,N_22757);
and U22889 (N_22889,N_22502,N_22420);
nand U22890 (N_22890,N_22649,N_22615);
and U22891 (N_22891,N_22657,N_22774);
and U22892 (N_22892,N_22391,N_22734);
nand U22893 (N_22893,N_22331,N_22222);
nand U22894 (N_22894,N_22293,N_22379);
or U22895 (N_22895,N_22562,N_22646);
nand U22896 (N_22896,N_22359,N_22276);
or U22897 (N_22897,N_22437,N_22281);
and U22898 (N_22898,N_22450,N_22445);
or U22899 (N_22899,N_22505,N_22550);
or U22900 (N_22900,N_22658,N_22460);
nor U22901 (N_22901,N_22759,N_22526);
nor U22902 (N_22902,N_22507,N_22374);
or U22903 (N_22903,N_22686,N_22676);
nand U22904 (N_22904,N_22588,N_22575);
and U22905 (N_22905,N_22766,N_22626);
or U22906 (N_22906,N_22383,N_22584);
or U22907 (N_22907,N_22485,N_22510);
nor U22908 (N_22908,N_22552,N_22639);
nand U22909 (N_22909,N_22305,N_22650);
or U22910 (N_22910,N_22659,N_22540);
nor U22911 (N_22911,N_22631,N_22476);
or U22912 (N_22912,N_22285,N_22664);
nand U22913 (N_22913,N_22337,N_22723);
and U22914 (N_22914,N_22772,N_22636);
or U22915 (N_22915,N_22261,N_22428);
nor U22916 (N_22916,N_22246,N_22452);
nor U22917 (N_22917,N_22537,N_22593);
nand U22918 (N_22918,N_22580,N_22746);
or U22919 (N_22919,N_22240,N_22689);
and U22920 (N_22920,N_22413,N_22366);
or U22921 (N_22921,N_22373,N_22532);
and U22922 (N_22922,N_22738,N_22758);
nand U22923 (N_22923,N_22619,N_22535);
nand U22924 (N_22924,N_22633,N_22696);
nand U22925 (N_22925,N_22741,N_22745);
and U22926 (N_22926,N_22538,N_22730);
nand U22927 (N_22927,N_22634,N_22678);
nor U22928 (N_22928,N_22775,N_22579);
xor U22929 (N_22929,N_22292,N_22663);
nand U22930 (N_22930,N_22737,N_22585);
or U22931 (N_22931,N_22613,N_22654);
or U22932 (N_22932,N_22229,N_22385);
xnor U22933 (N_22933,N_22431,N_22582);
and U22934 (N_22934,N_22473,N_22384);
or U22935 (N_22935,N_22353,N_22467);
or U22936 (N_22936,N_22513,N_22630);
nand U22937 (N_22937,N_22683,N_22235);
and U22938 (N_22938,N_22312,N_22548);
or U22939 (N_22939,N_22423,N_22733);
nor U22940 (N_22940,N_22788,N_22402);
or U22941 (N_22941,N_22527,N_22214);
xor U22942 (N_22942,N_22486,N_22372);
and U22943 (N_22943,N_22732,N_22706);
or U22944 (N_22944,N_22778,N_22322);
nand U22945 (N_22945,N_22242,N_22316);
or U22946 (N_22946,N_22260,N_22609);
or U22947 (N_22947,N_22735,N_22520);
and U22948 (N_22948,N_22404,N_22603);
nand U22949 (N_22949,N_22307,N_22524);
and U22950 (N_22950,N_22790,N_22362);
and U22951 (N_22951,N_22795,N_22301);
and U22952 (N_22952,N_22586,N_22648);
or U22953 (N_22953,N_22411,N_22370);
or U22954 (N_22954,N_22446,N_22463);
nand U22955 (N_22955,N_22208,N_22380);
nand U22956 (N_22956,N_22279,N_22570);
nand U22957 (N_22957,N_22751,N_22712);
nand U22958 (N_22958,N_22395,N_22781);
nor U22959 (N_22959,N_22699,N_22667);
and U22960 (N_22960,N_22244,N_22670);
xnor U22961 (N_22961,N_22462,N_22740);
or U22962 (N_22962,N_22509,N_22782);
and U22963 (N_22963,N_22624,N_22386);
nor U22964 (N_22964,N_22729,N_22326);
or U22965 (N_22965,N_22421,N_22643);
xnor U22966 (N_22966,N_22769,N_22203);
nor U22967 (N_22967,N_22419,N_22429);
nor U22968 (N_22968,N_22651,N_22255);
or U22969 (N_22969,N_22283,N_22553);
or U22970 (N_22970,N_22403,N_22779);
nand U22971 (N_22971,N_22539,N_22425);
and U22972 (N_22972,N_22607,N_22233);
xnor U22973 (N_22973,N_22216,N_22300);
nor U22974 (N_22974,N_22574,N_22708);
nand U22975 (N_22975,N_22490,N_22606);
or U22976 (N_22976,N_22350,N_22217);
nand U22977 (N_22977,N_22497,N_22594);
and U22978 (N_22978,N_22472,N_22653);
nor U22979 (N_22979,N_22773,N_22592);
nor U22980 (N_22980,N_22376,N_22258);
or U22981 (N_22981,N_22360,N_22336);
xor U22982 (N_22982,N_22342,N_22221);
nand U22983 (N_22983,N_22388,N_22750);
and U22984 (N_22984,N_22549,N_22672);
nand U22985 (N_22985,N_22345,N_22679);
and U22986 (N_22986,N_22355,N_22237);
or U22987 (N_22987,N_22530,N_22416);
and U22988 (N_22988,N_22253,N_22346);
nor U22989 (N_22989,N_22365,N_22765);
nor U22990 (N_22990,N_22335,N_22547);
or U22991 (N_22991,N_22310,N_22571);
and U22992 (N_22992,N_22536,N_22495);
nand U22993 (N_22993,N_22228,N_22367);
nand U22994 (N_22994,N_22302,N_22399);
nor U22995 (N_22995,N_22458,N_22703);
and U22996 (N_22996,N_22248,N_22600);
and U22997 (N_22997,N_22559,N_22514);
and U22998 (N_22998,N_22701,N_22693);
nor U22999 (N_22999,N_22263,N_22618);
and U23000 (N_23000,N_22792,N_22479);
or U23001 (N_23001,N_22597,N_22685);
nor U23002 (N_23002,N_22644,N_22432);
xnor U23003 (N_23003,N_22457,N_22722);
or U23004 (N_23004,N_22259,N_22328);
nand U23005 (N_23005,N_22433,N_22459);
nand U23006 (N_23006,N_22673,N_22238);
and U23007 (N_23007,N_22777,N_22487);
or U23008 (N_23008,N_22466,N_22796);
nand U23009 (N_23009,N_22414,N_22611);
and U23010 (N_23010,N_22687,N_22551);
and U23011 (N_23011,N_22219,N_22755);
nand U23012 (N_23012,N_22531,N_22770);
nand U23013 (N_23013,N_22661,N_22742);
nand U23014 (N_23014,N_22290,N_22731);
and U23015 (N_23015,N_22747,N_22357);
nand U23016 (N_23016,N_22478,N_22761);
or U23017 (N_23017,N_22682,N_22768);
nand U23018 (N_23018,N_22256,N_22470);
nor U23019 (N_23019,N_22227,N_22642);
and U23020 (N_23020,N_22250,N_22443);
nor U23021 (N_23021,N_22286,N_22488);
nand U23022 (N_23022,N_22684,N_22215);
and U23023 (N_23023,N_22455,N_22436);
and U23024 (N_23024,N_22744,N_22605);
nor U23025 (N_23025,N_22622,N_22799);
nand U23026 (N_23026,N_22655,N_22435);
and U23027 (N_23027,N_22717,N_22523);
nor U23028 (N_23028,N_22207,N_22727);
nand U23029 (N_23029,N_22610,N_22578);
or U23030 (N_23030,N_22465,N_22407);
and U23031 (N_23031,N_22780,N_22544);
or U23032 (N_23032,N_22762,N_22280);
or U23033 (N_23033,N_22724,N_22481);
nand U23034 (N_23034,N_22715,N_22556);
or U23035 (N_23035,N_22545,N_22697);
and U23036 (N_23036,N_22291,N_22262);
and U23037 (N_23037,N_22361,N_22410);
nor U23038 (N_23038,N_22713,N_22314);
nand U23039 (N_23039,N_22681,N_22371);
nand U23040 (N_23040,N_22330,N_22269);
xor U23041 (N_23041,N_22620,N_22645);
and U23042 (N_23042,N_22542,N_22702);
and U23043 (N_23043,N_22743,N_22477);
nand U23044 (N_23044,N_22343,N_22442);
and U23045 (N_23045,N_22333,N_22516);
and U23046 (N_23046,N_22406,N_22621);
or U23047 (N_23047,N_22518,N_22405);
or U23048 (N_23048,N_22794,N_22691);
nor U23049 (N_23049,N_22387,N_22764);
and U23050 (N_23050,N_22752,N_22392);
and U23051 (N_23051,N_22591,N_22329);
nand U23052 (N_23052,N_22625,N_22525);
and U23053 (N_23053,N_22569,N_22247);
and U23054 (N_23054,N_22771,N_22604);
nor U23055 (N_23055,N_22521,N_22754);
or U23056 (N_23056,N_22690,N_22204);
and U23057 (N_23057,N_22239,N_22503);
and U23058 (N_23058,N_22541,N_22348);
nand U23059 (N_23059,N_22441,N_22558);
and U23060 (N_23060,N_22468,N_22496);
nor U23061 (N_23061,N_22482,N_22581);
or U23062 (N_23062,N_22295,N_22319);
and U23063 (N_23063,N_22298,N_22427);
nand U23064 (N_23064,N_22671,N_22267);
nand U23065 (N_23065,N_22577,N_22426);
nor U23066 (N_23066,N_22475,N_22390);
or U23067 (N_23067,N_22254,N_22726);
or U23068 (N_23068,N_22783,N_22315);
and U23069 (N_23069,N_22382,N_22309);
and U23070 (N_23070,N_22274,N_22220);
and U23071 (N_23071,N_22797,N_22511);
nor U23072 (N_23072,N_22318,N_22710);
and U23073 (N_23073,N_22748,N_22264);
nand U23074 (N_23074,N_22647,N_22776);
and U23075 (N_23075,N_22251,N_22212);
nor U23076 (N_23076,N_22324,N_22736);
and U23077 (N_23077,N_22563,N_22296);
nor U23078 (N_23078,N_22599,N_22224);
and U23079 (N_23079,N_22303,N_22323);
nor U23080 (N_23080,N_22489,N_22638);
nor U23081 (N_23081,N_22278,N_22785);
nor U23082 (N_23082,N_22725,N_22243);
nor U23083 (N_23083,N_22226,N_22627);
and U23084 (N_23084,N_22231,N_22711);
and U23085 (N_23085,N_22271,N_22417);
or U23086 (N_23086,N_22700,N_22218);
nand U23087 (N_23087,N_22484,N_22275);
and U23088 (N_23088,N_22529,N_22572);
and U23089 (N_23089,N_22494,N_22338);
nor U23090 (N_23090,N_22709,N_22358);
nand U23091 (N_23091,N_22557,N_22528);
nand U23092 (N_23092,N_22225,N_22377);
nor U23093 (N_23093,N_22739,N_22398);
nor U23094 (N_23094,N_22287,N_22546);
nor U23095 (N_23095,N_22210,N_22596);
and U23096 (N_23096,N_22749,N_22265);
and U23097 (N_23097,N_22430,N_22522);
or U23098 (N_23098,N_22327,N_22561);
nand U23099 (N_23099,N_22438,N_22454);
nor U23100 (N_23100,N_22592,N_22454);
xor U23101 (N_23101,N_22603,N_22488);
nor U23102 (N_23102,N_22440,N_22342);
nor U23103 (N_23103,N_22700,N_22269);
nand U23104 (N_23104,N_22301,N_22243);
and U23105 (N_23105,N_22225,N_22558);
nor U23106 (N_23106,N_22496,N_22315);
and U23107 (N_23107,N_22460,N_22427);
nor U23108 (N_23108,N_22221,N_22768);
nor U23109 (N_23109,N_22207,N_22565);
or U23110 (N_23110,N_22576,N_22402);
nand U23111 (N_23111,N_22483,N_22661);
or U23112 (N_23112,N_22554,N_22473);
or U23113 (N_23113,N_22516,N_22484);
and U23114 (N_23114,N_22306,N_22792);
nand U23115 (N_23115,N_22282,N_22402);
and U23116 (N_23116,N_22767,N_22391);
nand U23117 (N_23117,N_22621,N_22410);
and U23118 (N_23118,N_22453,N_22615);
and U23119 (N_23119,N_22525,N_22502);
nand U23120 (N_23120,N_22605,N_22405);
nand U23121 (N_23121,N_22274,N_22737);
nor U23122 (N_23122,N_22333,N_22667);
xnor U23123 (N_23123,N_22791,N_22538);
or U23124 (N_23124,N_22455,N_22468);
nor U23125 (N_23125,N_22502,N_22528);
and U23126 (N_23126,N_22254,N_22204);
nand U23127 (N_23127,N_22267,N_22792);
or U23128 (N_23128,N_22276,N_22542);
nand U23129 (N_23129,N_22404,N_22610);
nor U23130 (N_23130,N_22453,N_22599);
and U23131 (N_23131,N_22441,N_22367);
and U23132 (N_23132,N_22765,N_22330);
or U23133 (N_23133,N_22539,N_22209);
nand U23134 (N_23134,N_22773,N_22437);
and U23135 (N_23135,N_22724,N_22728);
nor U23136 (N_23136,N_22466,N_22574);
or U23137 (N_23137,N_22418,N_22459);
or U23138 (N_23138,N_22410,N_22425);
nor U23139 (N_23139,N_22376,N_22721);
and U23140 (N_23140,N_22373,N_22513);
nor U23141 (N_23141,N_22271,N_22280);
nand U23142 (N_23142,N_22477,N_22771);
nand U23143 (N_23143,N_22523,N_22232);
or U23144 (N_23144,N_22240,N_22367);
and U23145 (N_23145,N_22230,N_22717);
and U23146 (N_23146,N_22369,N_22513);
nor U23147 (N_23147,N_22737,N_22475);
nand U23148 (N_23148,N_22580,N_22317);
nand U23149 (N_23149,N_22220,N_22676);
and U23150 (N_23150,N_22587,N_22240);
and U23151 (N_23151,N_22427,N_22753);
nand U23152 (N_23152,N_22654,N_22653);
nor U23153 (N_23153,N_22216,N_22619);
or U23154 (N_23154,N_22481,N_22402);
or U23155 (N_23155,N_22682,N_22703);
and U23156 (N_23156,N_22386,N_22728);
or U23157 (N_23157,N_22500,N_22785);
and U23158 (N_23158,N_22736,N_22607);
nand U23159 (N_23159,N_22700,N_22342);
and U23160 (N_23160,N_22264,N_22594);
or U23161 (N_23161,N_22669,N_22333);
nor U23162 (N_23162,N_22510,N_22455);
and U23163 (N_23163,N_22794,N_22333);
or U23164 (N_23164,N_22698,N_22478);
or U23165 (N_23165,N_22657,N_22419);
and U23166 (N_23166,N_22440,N_22571);
or U23167 (N_23167,N_22240,N_22481);
or U23168 (N_23168,N_22398,N_22201);
and U23169 (N_23169,N_22380,N_22550);
and U23170 (N_23170,N_22446,N_22423);
nand U23171 (N_23171,N_22795,N_22392);
and U23172 (N_23172,N_22494,N_22568);
nand U23173 (N_23173,N_22357,N_22603);
nand U23174 (N_23174,N_22259,N_22612);
nor U23175 (N_23175,N_22570,N_22691);
nand U23176 (N_23176,N_22640,N_22734);
nand U23177 (N_23177,N_22683,N_22443);
nand U23178 (N_23178,N_22735,N_22236);
nand U23179 (N_23179,N_22238,N_22293);
nand U23180 (N_23180,N_22486,N_22374);
nor U23181 (N_23181,N_22226,N_22631);
and U23182 (N_23182,N_22279,N_22497);
nand U23183 (N_23183,N_22610,N_22598);
nand U23184 (N_23184,N_22564,N_22338);
and U23185 (N_23185,N_22328,N_22221);
and U23186 (N_23186,N_22434,N_22382);
or U23187 (N_23187,N_22559,N_22268);
and U23188 (N_23188,N_22607,N_22705);
nand U23189 (N_23189,N_22516,N_22278);
nor U23190 (N_23190,N_22245,N_22746);
and U23191 (N_23191,N_22224,N_22321);
nand U23192 (N_23192,N_22719,N_22707);
nor U23193 (N_23193,N_22516,N_22613);
and U23194 (N_23194,N_22587,N_22416);
and U23195 (N_23195,N_22635,N_22788);
nor U23196 (N_23196,N_22302,N_22691);
nor U23197 (N_23197,N_22537,N_22663);
or U23198 (N_23198,N_22752,N_22726);
or U23199 (N_23199,N_22718,N_22229);
or U23200 (N_23200,N_22503,N_22221);
nand U23201 (N_23201,N_22373,N_22575);
nand U23202 (N_23202,N_22436,N_22725);
nand U23203 (N_23203,N_22454,N_22255);
or U23204 (N_23204,N_22543,N_22626);
and U23205 (N_23205,N_22488,N_22381);
or U23206 (N_23206,N_22374,N_22469);
nand U23207 (N_23207,N_22560,N_22615);
and U23208 (N_23208,N_22454,N_22771);
and U23209 (N_23209,N_22589,N_22319);
nor U23210 (N_23210,N_22235,N_22510);
nand U23211 (N_23211,N_22654,N_22498);
xor U23212 (N_23212,N_22207,N_22231);
nand U23213 (N_23213,N_22307,N_22296);
nand U23214 (N_23214,N_22558,N_22762);
nand U23215 (N_23215,N_22728,N_22340);
or U23216 (N_23216,N_22549,N_22753);
nand U23217 (N_23217,N_22430,N_22714);
nor U23218 (N_23218,N_22523,N_22253);
and U23219 (N_23219,N_22222,N_22582);
and U23220 (N_23220,N_22293,N_22739);
nand U23221 (N_23221,N_22219,N_22235);
or U23222 (N_23222,N_22511,N_22698);
and U23223 (N_23223,N_22343,N_22474);
or U23224 (N_23224,N_22449,N_22227);
nor U23225 (N_23225,N_22676,N_22420);
and U23226 (N_23226,N_22760,N_22330);
xor U23227 (N_23227,N_22462,N_22245);
xnor U23228 (N_23228,N_22424,N_22251);
nor U23229 (N_23229,N_22614,N_22497);
nor U23230 (N_23230,N_22520,N_22703);
nand U23231 (N_23231,N_22492,N_22329);
or U23232 (N_23232,N_22760,N_22706);
and U23233 (N_23233,N_22531,N_22661);
and U23234 (N_23234,N_22754,N_22328);
nor U23235 (N_23235,N_22690,N_22499);
or U23236 (N_23236,N_22214,N_22218);
and U23237 (N_23237,N_22325,N_22437);
and U23238 (N_23238,N_22222,N_22734);
or U23239 (N_23239,N_22380,N_22218);
or U23240 (N_23240,N_22769,N_22693);
xnor U23241 (N_23241,N_22553,N_22768);
and U23242 (N_23242,N_22387,N_22261);
nor U23243 (N_23243,N_22280,N_22210);
nand U23244 (N_23244,N_22201,N_22345);
nor U23245 (N_23245,N_22503,N_22711);
nand U23246 (N_23246,N_22623,N_22531);
nand U23247 (N_23247,N_22234,N_22305);
or U23248 (N_23248,N_22333,N_22250);
nand U23249 (N_23249,N_22503,N_22623);
nor U23250 (N_23250,N_22732,N_22603);
nor U23251 (N_23251,N_22688,N_22316);
nand U23252 (N_23252,N_22587,N_22405);
nor U23253 (N_23253,N_22203,N_22668);
and U23254 (N_23254,N_22716,N_22571);
nor U23255 (N_23255,N_22484,N_22607);
nor U23256 (N_23256,N_22646,N_22356);
nand U23257 (N_23257,N_22394,N_22325);
and U23258 (N_23258,N_22651,N_22358);
nor U23259 (N_23259,N_22398,N_22677);
nand U23260 (N_23260,N_22648,N_22568);
and U23261 (N_23261,N_22598,N_22590);
and U23262 (N_23262,N_22239,N_22245);
nor U23263 (N_23263,N_22320,N_22543);
nor U23264 (N_23264,N_22472,N_22453);
or U23265 (N_23265,N_22445,N_22649);
nand U23266 (N_23266,N_22667,N_22640);
nand U23267 (N_23267,N_22412,N_22458);
nand U23268 (N_23268,N_22538,N_22548);
nor U23269 (N_23269,N_22240,N_22624);
and U23270 (N_23270,N_22736,N_22394);
or U23271 (N_23271,N_22238,N_22239);
or U23272 (N_23272,N_22682,N_22573);
nor U23273 (N_23273,N_22345,N_22735);
nor U23274 (N_23274,N_22663,N_22368);
nor U23275 (N_23275,N_22489,N_22445);
and U23276 (N_23276,N_22755,N_22227);
nor U23277 (N_23277,N_22261,N_22377);
nor U23278 (N_23278,N_22797,N_22613);
and U23279 (N_23279,N_22307,N_22654);
nor U23280 (N_23280,N_22697,N_22314);
or U23281 (N_23281,N_22501,N_22633);
and U23282 (N_23282,N_22407,N_22590);
nor U23283 (N_23283,N_22774,N_22237);
and U23284 (N_23284,N_22227,N_22340);
nand U23285 (N_23285,N_22431,N_22217);
or U23286 (N_23286,N_22351,N_22402);
nor U23287 (N_23287,N_22677,N_22653);
nor U23288 (N_23288,N_22737,N_22726);
nor U23289 (N_23289,N_22482,N_22337);
or U23290 (N_23290,N_22626,N_22521);
nor U23291 (N_23291,N_22710,N_22243);
and U23292 (N_23292,N_22566,N_22410);
or U23293 (N_23293,N_22489,N_22436);
and U23294 (N_23294,N_22769,N_22620);
nor U23295 (N_23295,N_22693,N_22623);
nand U23296 (N_23296,N_22408,N_22275);
nand U23297 (N_23297,N_22226,N_22433);
nor U23298 (N_23298,N_22305,N_22280);
or U23299 (N_23299,N_22502,N_22302);
nor U23300 (N_23300,N_22206,N_22597);
or U23301 (N_23301,N_22317,N_22320);
or U23302 (N_23302,N_22686,N_22480);
and U23303 (N_23303,N_22287,N_22734);
and U23304 (N_23304,N_22651,N_22592);
or U23305 (N_23305,N_22508,N_22670);
and U23306 (N_23306,N_22488,N_22484);
or U23307 (N_23307,N_22600,N_22587);
or U23308 (N_23308,N_22582,N_22253);
or U23309 (N_23309,N_22745,N_22409);
nand U23310 (N_23310,N_22424,N_22227);
nand U23311 (N_23311,N_22421,N_22272);
and U23312 (N_23312,N_22598,N_22260);
xor U23313 (N_23313,N_22681,N_22556);
nor U23314 (N_23314,N_22280,N_22535);
or U23315 (N_23315,N_22241,N_22480);
and U23316 (N_23316,N_22677,N_22532);
or U23317 (N_23317,N_22461,N_22601);
or U23318 (N_23318,N_22360,N_22330);
nor U23319 (N_23319,N_22742,N_22574);
nor U23320 (N_23320,N_22510,N_22296);
and U23321 (N_23321,N_22524,N_22451);
and U23322 (N_23322,N_22420,N_22436);
nand U23323 (N_23323,N_22290,N_22484);
or U23324 (N_23324,N_22599,N_22272);
nand U23325 (N_23325,N_22757,N_22226);
nand U23326 (N_23326,N_22319,N_22408);
nand U23327 (N_23327,N_22450,N_22376);
and U23328 (N_23328,N_22447,N_22746);
xnor U23329 (N_23329,N_22523,N_22244);
and U23330 (N_23330,N_22635,N_22544);
nor U23331 (N_23331,N_22779,N_22783);
nor U23332 (N_23332,N_22235,N_22764);
nand U23333 (N_23333,N_22574,N_22343);
or U23334 (N_23334,N_22625,N_22512);
or U23335 (N_23335,N_22373,N_22348);
nand U23336 (N_23336,N_22301,N_22553);
and U23337 (N_23337,N_22638,N_22213);
or U23338 (N_23338,N_22475,N_22434);
nand U23339 (N_23339,N_22444,N_22451);
and U23340 (N_23340,N_22409,N_22289);
and U23341 (N_23341,N_22351,N_22503);
nor U23342 (N_23342,N_22202,N_22762);
xor U23343 (N_23343,N_22715,N_22463);
and U23344 (N_23344,N_22694,N_22262);
and U23345 (N_23345,N_22388,N_22541);
and U23346 (N_23346,N_22770,N_22728);
and U23347 (N_23347,N_22418,N_22633);
nand U23348 (N_23348,N_22799,N_22607);
nor U23349 (N_23349,N_22301,N_22575);
nor U23350 (N_23350,N_22426,N_22433);
or U23351 (N_23351,N_22311,N_22633);
and U23352 (N_23352,N_22421,N_22247);
and U23353 (N_23353,N_22400,N_22439);
nor U23354 (N_23354,N_22741,N_22598);
nand U23355 (N_23355,N_22684,N_22550);
nor U23356 (N_23356,N_22201,N_22764);
nand U23357 (N_23357,N_22446,N_22551);
and U23358 (N_23358,N_22665,N_22231);
nor U23359 (N_23359,N_22237,N_22657);
or U23360 (N_23360,N_22737,N_22356);
and U23361 (N_23361,N_22427,N_22273);
nand U23362 (N_23362,N_22598,N_22769);
nor U23363 (N_23363,N_22364,N_22239);
nand U23364 (N_23364,N_22481,N_22205);
nand U23365 (N_23365,N_22592,N_22656);
nor U23366 (N_23366,N_22416,N_22743);
nor U23367 (N_23367,N_22222,N_22463);
or U23368 (N_23368,N_22234,N_22689);
or U23369 (N_23369,N_22658,N_22424);
nand U23370 (N_23370,N_22733,N_22305);
nor U23371 (N_23371,N_22576,N_22424);
nor U23372 (N_23372,N_22590,N_22365);
nor U23373 (N_23373,N_22589,N_22632);
and U23374 (N_23374,N_22476,N_22740);
and U23375 (N_23375,N_22614,N_22691);
nor U23376 (N_23376,N_22780,N_22700);
nand U23377 (N_23377,N_22254,N_22319);
nand U23378 (N_23378,N_22361,N_22724);
or U23379 (N_23379,N_22274,N_22333);
nor U23380 (N_23380,N_22768,N_22694);
nor U23381 (N_23381,N_22763,N_22401);
or U23382 (N_23382,N_22625,N_22541);
or U23383 (N_23383,N_22632,N_22567);
nor U23384 (N_23384,N_22216,N_22640);
and U23385 (N_23385,N_22285,N_22420);
or U23386 (N_23386,N_22419,N_22437);
nor U23387 (N_23387,N_22243,N_22586);
and U23388 (N_23388,N_22771,N_22223);
or U23389 (N_23389,N_22652,N_22478);
nand U23390 (N_23390,N_22257,N_22521);
nand U23391 (N_23391,N_22500,N_22218);
nor U23392 (N_23392,N_22269,N_22746);
nor U23393 (N_23393,N_22398,N_22368);
or U23394 (N_23394,N_22599,N_22691);
nand U23395 (N_23395,N_22281,N_22629);
nand U23396 (N_23396,N_22414,N_22218);
and U23397 (N_23397,N_22506,N_22685);
and U23398 (N_23398,N_22560,N_22249);
nor U23399 (N_23399,N_22550,N_22359);
or U23400 (N_23400,N_23201,N_23324);
and U23401 (N_23401,N_22948,N_23273);
nand U23402 (N_23402,N_23236,N_22936);
nor U23403 (N_23403,N_22988,N_23178);
nor U23404 (N_23404,N_23154,N_23058);
or U23405 (N_23405,N_23361,N_22895);
nor U23406 (N_23406,N_22943,N_23169);
and U23407 (N_23407,N_22894,N_23312);
or U23408 (N_23408,N_23174,N_22966);
nor U23409 (N_23409,N_23101,N_23334);
and U23410 (N_23410,N_22876,N_22823);
nand U23411 (N_23411,N_22932,N_22928);
and U23412 (N_23412,N_22801,N_23213);
nor U23413 (N_23413,N_23184,N_22973);
and U23414 (N_23414,N_23149,N_23374);
nor U23415 (N_23415,N_22884,N_23151);
nand U23416 (N_23416,N_23067,N_23311);
or U23417 (N_23417,N_23116,N_23243);
nor U23418 (N_23418,N_23392,N_22912);
or U23419 (N_23419,N_22864,N_23259);
or U23420 (N_23420,N_23124,N_22870);
and U23421 (N_23421,N_23382,N_23349);
nor U23422 (N_23422,N_23222,N_23113);
or U23423 (N_23423,N_23145,N_22947);
and U23424 (N_23424,N_23224,N_23341);
and U23425 (N_23425,N_23132,N_23207);
and U23426 (N_23426,N_23269,N_22938);
nor U23427 (N_23427,N_23246,N_23363);
or U23428 (N_23428,N_23338,N_22962);
or U23429 (N_23429,N_22828,N_23195);
or U23430 (N_23430,N_23142,N_22993);
and U23431 (N_23431,N_22940,N_23267);
nand U23432 (N_23432,N_22907,N_23054);
xnor U23433 (N_23433,N_23331,N_23390);
nand U23434 (N_23434,N_23255,N_23032);
nor U23435 (N_23435,N_23176,N_23278);
or U23436 (N_23436,N_23394,N_23097);
or U23437 (N_23437,N_23064,N_23025);
nor U23438 (N_23438,N_23036,N_23128);
and U23439 (N_23439,N_22979,N_23021);
or U23440 (N_23440,N_23396,N_22808);
nor U23441 (N_23441,N_23035,N_23281);
nor U23442 (N_23442,N_22920,N_22904);
nand U23443 (N_23443,N_22980,N_23297);
and U23444 (N_23444,N_23196,N_23130);
or U23445 (N_23445,N_22891,N_22924);
or U23446 (N_23446,N_22939,N_23364);
and U23447 (N_23447,N_22995,N_23314);
and U23448 (N_23448,N_22969,N_22976);
and U23449 (N_23449,N_23099,N_23003);
nor U23450 (N_23450,N_23013,N_22923);
and U23451 (N_23451,N_23117,N_22992);
and U23452 (N_23452,N_23354,N_22862);
and U23453 (N_23453,N_23308,N_23004);
and U23454 (N_23454,N_23048,N_22883);
nor U23455 (N_23455,N_23275,N_23114);
and U23456 (N_23456,N_22825,N_22889);
or U23457 (N_23457,N_23010,N_22816);
and U23458 (N_23458,N_23147,N_22986);
and U23459 (N_23459,N_22925,N_23052);
or U23460 (N_23460,N_22837,N_22944);
and U23461 (N_23461,N_23371,N_23328);
nand U23462 (N_23462,N_22952,N_23194);
nand U23463 (N_23463,N_23143,N_23031);
nand U23464 (N_23464,N_22873,N_23288);
nand U23465 (N_23465,N_23106,N_23172);
nor U23466 (N_23466,N_23138,N_23105);
nand U23467 (N_23467,N_22908,N_23001);
nand U23468 (N_23468,N_22896,N_23082);
or U23469 (N_23469,N_23070,N_23129);
nand U23470 (N_23470,N_23379,N_22983);
or U23471 (N_23471,N_23245,N_23313);
or U23472 (N_23472,N_23310,N_22856);
nand U23473 (N_23473,N_22806,N_22874);
nand U23474 (N_23474,N_23388,N_23103);
nor U23475 (N_23475,N_23009,N_23357);
and U23476 (N_23476,N_23237,N_23330);
nor U23477 (N_23477,N_23265,N_23285);
and U23478 (N_23478,N_23059,N_22974);
and U23479 (N_23479,N_22892,N_22968);
nand U23480 (N_23480,N_22833,N_22842);
nor U23481 (N_23481,N_23333,N_23266);
nor U23482 (N_23482,N_23044,N_23295);
or U23483 (N_23483,N_23040,N_23309);
nand U23484 (N_23484,N_23028,N_23321);
and U23485 (N_23485,N_23034,N_23289);
nor U23486 (N_23486,N_23370,N_23080);
nand U23487 (N_23487,N_22849,N_22865);
nor U23488 (N_23488,N_22846,N_23220);
or U23489 (N_23489,N_23042,N_23022);
or U23490 (N_23490,N_23387,N_22970);
nand U23491 (N_23491,N_23024,N_23152);
or U23492 (N_23492,N_22918,N_23107);
and U23493 (N_23493,N_22893,N_23230);
and U23494 (N_23494,N_22934,N_23376);
nor U23495 (N_23495,N_23386,N_23261);
nand U23496 (N_23496,N_23346,N_22963);
nor U23497 (N_23497,N_23134,N_22814);
and U23498 (N_23498,N_23131,N_23298);
nand U23499 (N_23499,N_22991,N_23206);
or U23500 (N_23500,N_22840,N_22852);
nand U23501 (N_23501,N_23316,N_23326);
or U23502 (N_23502,N_23011,N_22949);
and U23503 (N_23503,N_23305,N_23214);
nand U23504 (N_23504,N_22809,N_23381);
and U23505 (N_23505,N_23204,N_23320);
nor U23506 (N_23506,N_22946,N_22901);
and U23507 (N_23507,N_22804,N_23368);
nor U23508 (N_23508,N_23358,N_22917);
and U23509 (N_23509,N_23175,N_23192);
nand U23510 (N_23510,N_23228,N_23292);
nand U23511 (N_23511,N_22942,N_23125);
or U23512 (N_23512,N_23060,N_22855);
nand U23513 (N_23513,N_22960,N_23203);
or U23514 (N_23514,N_23133,N_23257);
nor U23515 (N_23515,N_23232,N_23280);
nor U23516 (N_23516,N_23247,N_22848);
nor U23517 (N_23517,N_23355,N_23144);
and U23518 (N_23518,N_23264,N_23209);
or U23519 (N_23519,N_23072,N_23344);
nand U23520 (N_23520,N_23014,N_23348);
nor U23521 (N_23521,N_22909,N_23015);
nand U23522 (N_23522,N_23084,N_22810);
nand U23523 (N_23523,N_23197,N_23187);
nand U23524 (N_23524,N_23023,N_22826);
or U23525 (N_23525,N_23073,N_23063);
or U23526 (N_23526,N_23367,N_22857);
or U23527 (N_23527,N_22898,N_23115);
and U23528 (N_23528,N_23337,N_22836);
nor U23529 (N_23529,N_22956,N_22994);
nand U23530 (N_23530,N_23171,N_22835);
nor U23531 (N_23531,N_23141,N_22916);
or U23532 (N_23532,N_23353,N_22868);
nor U23533 (N_23533,N_23110,N_23085);
xor U23534 (N_23534,N_22999,N_22841);
and U23535 (N_23535,N_22875,N_22978);
or U23536 (N_23536,N_23233,N_23239);
or U23537 (N_23537,N_22933,N_22921);
nor U23538 (N_23538,N_23057,N_23329);
or U23539 (N_23539,N_22813,N_23244);
nand U23540 (N_23540,N_23210,N_23002);
nand U23541 (N_23541,N_22900,N_23083);
nor U23542 (N_23542,N_23166,N_22977);
nor U23543 (N_23543,N_23254,N_22812);
or U23544 (N_23544,N_23339,N_23350);
or U23545 (N_23545,N_22869,N_22905);
xnor U23546 (N_23546,N_23325,N_23007);
nor U23547 (N_23547,N_22850,N_22866);
nand U23548 (N_23548,N_22955,N_23343);
nor U23549 (N_23549,N_23071,N_22987);
or U23550 (N_23550,N_23157,N_23263);
nor U23551 (N_23551,N_23074,N_23167);
nand U23552 (N_23552,N_22890,N_23050);
nor U23553 (N_23553,N_23322,N_23177);
nor U23554 (N_23554,N_22819,N_23109);
nor U23555 (N_23555,N_22984,N_22871);
or U23556 (N_23556,N_23347,N_23284);
or U23557 (N_23557,N_22821,N_23090);
and U23558 (N_23558,N_22996,N_23282);
and U23559 (N_23559,N_22843,N_23356);
and U23560 (N_23560,N_23231,N_23122);
or U23561 (N_23561,N_22967,N_23291);
or U23562 (N_23562,N_23121,N_23340);
and U23563 (N_23563,N_22919,N_22975);
nor U23564 (N_23564,N_22827,N_22863);
or U23565 (N_23565,N_23006,N_23108);
and U23566 (N_23566,N_23079,N_22867);
nand U23567 (N_23567,N_23127,N_22844);
and U23568 (N_23568,N_23148,N_22926);
nor U23569 (N_23569,N_23218,N_23077);
nand U23570 (N_23570,N_22990,N_23216);
nand U23571 (N_23571,N_23181,N_23037);
nor U23572 (N_23572,N_23159,N_23153);
nor U23573 (N_23573,N_23190,N_22805);
or U23574 (N_23574,N_23179,N_22950);
and U23575 (N_23575,N_23193,N_23053);
nor U23576 (N_23576,N_23241,N_23251);
xor U23577 (N_23577,N_22811,N_22817);
xor U23578 (N_23578,N_23199,N_22982);
and U23579 (N_23579,N_23307,N_23317);
and U23580 (N_23580,N_22954,N_23296);
and U23581 (N_23581,N_23091,N_22965);
nand U23582 (N_23582,N_23018,N_23252);
or U23583 (N_23583,N_22861,N_22911);
or U23584 (N_23584,N_23345,N_22830);
nor U23585 (N_23585,N_23397,N_23158);
and U23586 (N_23586,N_23260,N_22929);
and U23587 (N_23587,N_23399,N_23253);
or U23588 (N_23588,N_23198,N_23319);
and U23589 (N_23589,N_23258,N_22910);
xor U23590 (N_23590,N_23069,N_23182);
and U23591 (N_23591,N_23160,N_23104);
or U23592 (N_23592,N_23030,N_23005);
nor U23593 (N_23593,N_23208,N_23119);
nor U23594 (N_23594,N_23362,N_22888);
nor U23595 (N_23595,N_23017,N_22807);
nor U23596 (N_23596,N_22877,N_23234);
nand U23597 (N_23597,N_23045,N_22872);
nor U23598 (N_23598,N_23062,N_23094);
nor U23599 (N_23599,N_22902,N_23235);
nand U23600 (N_23600,N_23229,N_22951);
nand U23601 (N_23601,N_23373,N_23164);
or U23602 (N_23602,N_22829,N_22941);
and U23603 (N_23603,N_23256,N_23238);
or U23604 (N_23604,N_22972,N_23183);
and U23605 (N_23605,N_23302,N_23173);
nor U23606 (N_23606,N_23276,N_23066);
and U23607 (N_23607,N_23212,N_22845);
nor U23608 (N_23608,N_22906,N_22927);
nor U23609 (N_23609,N_23262,N_23270);
nor U23610 (N_23610,N_23093,N_23078);
and U23611 (N_23611,N_23046,N_23240);
nand U23612 (N_23612,N_23068,N_23287);
and U23613 (N_23613,N_23095,N_23351);
nand U23614 (N_23614,N_23016,N_22998);
nor U23615 (N_23615,N_22945,N_23019);
or U23616 (N_23616,N_22903,N_23055);
nand U23617 (N_23617,N_23290,N_22803);
or U23618 (N_23618,N_22886,N_23393);
nand U23619 (N_23619,N_23137,N_22800);
nand U23620 (N_23620,N_23268,N_23372);
nor U23621 (N_23621,N_23027,N_23126);
or U23622 (N_23622,N_23304,N_23162);
nor U23623 (N_23623,N_22854,N_23391);
and U23624 (N_23624,N_22935,N_23301);
nand U23625 (N_23625,N_22815,N_23395);
and U23626 (N_23626,N_23100,N_23377);
and U23627 (N_23627,N_23012,N_22915);
or U23628 (N_23628,N_23219,N_23140);
or U23629 (N_23629,N_23200,N_23336);
nand U23630 (N_23630,N_23375,N_22820);
nor U23631 (N_23631,N_23065,N_23286);
and U23632 (N_23632,N_23051,N_23185);
nor U23633 (N_23633,N_22822,N_22985);
nor U23634 (N_23634,N_23102,N_22989);
nand U23635 (N_23635,N_22860,N_23061);
nor U23636 (N_23636,N_23092,N_23250);
nor U23637 (N_23637,N_23360,N_23156);
nand U23638 (N_23638,N_23248,N_23352);
and U23639 (N_23639,N_23180,N_22851);
or U23640 (N_23640,N_23029,N_23039);
and U23641 (N_23641,N_22930,N_23242);
nand U23642 (N_23642,N_23283,N_23098);
or U23643 (N_23643,N_22981,N_22958);
nor U23644 (N_23644,N_23191,N_23189);
nor U23645 (N_23645,N_23384,N_22882);
and U23646 (N_23646,N_23038,N_23088);
or U23647 (N_23647,N_23111,N_23161);
or U23648 (N_23648,N_22953,N_22832);
nor U23649 (N_23649,N_23365,N_23383);
nor U23650 (N_23650,N_22878,N_22914);
nor U23651 (N_23651,N_23089,N_23398);
and U23652 (N_23652,N_23366,N_23369);
or U23653 (N_23653,N_22931,N_23026);
or U23654 (N_23654,N_22971,N_22957);
nor U23655 (N_23655,N_22839,N_22959);
and U23656 (N_23656,N_22922,N_23335);
nand U23657 (N_23657,N_23150,N_23223);
and U23658 (N_23658,N_23139,N_23136);
nand U23659 (N_23659,N_23043,N_22824);
or U23660 (N_23660,N_22859,N_22899);
nand U23661 (N_23661,N_23225,N_22937);
nand U23662 (N_23662,N_23075,N_23076);
or U23663 (N_23663,N_23385,N_22858);
and U23664 (N_23664,N_23323,N_23294);
nand U23665 (N_23665,N_22897,N_23000);
or U23666 (N_23666,N_23168,N_22997);
or U23667 (N_23667,N_23120,N_23215);
and U23668 (N_23668,N_23135,N_23165);
nor U23669 (N_23669,N_22853,N_23202);
nor U23670 (N_23670,N_23279,N_22838);
or U23671 (N_23671,N_23020,N_22913);
nand U23672 (N_23672,N_22879,N_23274);
and U23673 (N_23673,N_23327,N_23047);
and U23674 (N_23674,N_23146,N_22961);
or U23675 (N_23675,N_23211,N_22964);
xor U23676 (N_23676,N_23186,N_23123);
and U23677 (N_23677,N_23300,N_23188);
or U23678 (N_23678,N_23087,N_23112);
nand U23679 (N_23679,N_23170,N_23249);
nand U23680 (N_23680,N_23217,N_23342);
nor U23681 (N_23681,N_23272,N_22818);
or U23682 (N_23682,N_23226,N_22802);
or U23683 (N_23683,N_22880,N_23008);
or U23684 (N_23684,N_23299,N_23056);
or U23685 (N_23685,N_22834,N_23293);
and U23686 (N_23686,N_23118,N_23155);
nand U23687 (N_23687,N_23315,N_23096);
nor U23688 (N_23688,N_23303,N_23380);
nor U23689 (N_23689,N_23389,N_23378);
nand U23690 (N_23690,N_23318,N_23221);
nand U23691 (N_23691,N_23033,N_23227);
and U23692 (N_23692,N_22881,N_22847);
and U23693 (N_23693,N_23306,N_23081);
and U23694 (N_23694,N_23359,N_23086);
nor U23695 (N_23695,N_23049,N_23271);
and U23696 (N_23696,N_23277,N_23041);
nor U23697 (N_23697,N_22831,N_22887);
nor U23698 (N_23698,N_23163,N_23205);
nand U23699 (N_23699,N_22885,N_23332);
and U23700 (N_23700,N_22830,N_22922);
and U23701 (N_23701,N_23269,N_23373);
nand U23702 (N_23702,N_23362,N_23265);
or U23703 (N_23703,N_23263,N_23286);
nor U23704 (N_23704,N_23091,N_23307);
nand U23705 (N_23705,N_23254,N_23250);
and U23706 (N_23706,N_23383,N_23323);
nor U23707 (N_23707,N_23009,N_22923);
and U23708 (N_23708,N_23100,N_22955);
nor U23709 (N_23709,N_22865,N_23000);
or U23710 (N_23710,N_23386,N_23173);
nor U23711 (N_23711,N_23322,N_23155);
nand U23712 (N_23712,N_23080,N_23306);
and U23713 (N_23713,N_23242,N_23363);
or U23714 (N_23714,N_23334,N_22897);
and U23715 (N_23715,N_23073,N_23396);
nand U23716 (N_23716,N_23256,N_23131);
xor U23717 (N_23717,N_23253,N_23275);
or U23718 (N_23718,N_22873,N_22904);
or U23719 (N_23719,N_23254,N_23299);
and U23720 (N_23720,N_23323,N_22808);
or U23721 (N_23721,N_23060,N_23151);
or U23722 (N_23722,N_23190,N_23288);
and U23723 (N_23723,N_23100,N_23080);
and U23724 (N_23724,N_23092,N_22971);
nand U23725 (N_23725,N_23216,N_23006);
nor U23726 (N_23726,N_23208,N_22925);
or U23727 (N_23727,N_23047,N_22925);
and U23728 (N_23728,N_23186,N_23187);
and U23729 (N_23729,N_23273,N_22822);
nand U23730 (N_23730,N_23164,N_22895);
nand U23731 (N_23731,N_23249,N_23089);
or U23732 (N_23732,N_22838,N_22828);
and U23733 (N_23733,N_22973,N_23160);
nor U23734 (N_23734,N_23377,N_22923);
nor U23735 (N_23735,N_23344,N_23250);
and U23736 (N_23736,N_23093,N_23253);
nand U23737 (N_23737,N_23022,N_23018);
nand U23738 (N_23738,N_23175,N_23207);
or U23739 (N_23739,N_23219,N_23245);
nor U23740 (N_23740,N_23284,N_22866);
and U23741 (N_23741,N_23263,N_23073);
nand U23742 (N_23742,N_23285,N_22960);
nand U23743 (N_23743,N_23301,N_23234);
nor U23744 (N_23744,N_23044,N_22836);
nand U23745 (N_23745,N_23390,N_23353);
or U23746 (N_23746,N_23112,N_23144);
and U23747 (N_23747,N_23163,N_22993);
nor U23748 (N_23748,N_23161,N_23243);
and U23749 (N_23749,N_22960,N_22875);
or U23750 (N_23750,N_23271,N_22859);
nand U23751 (N_23751,N_22876,N_22963);
or U23752 (N_23752,N_23374,N_22802);
nor U23753 (N_23753,N_22969,N_23031);
or U23754 (N_23754,N_23220,N_23060);
nand U23755 (N_23755,N_23259,N_22991);
nand U23756 (N_23756,N_23164,N_23338);
nor U23757 (N_23757,N_23009,N_23283);
or U23758 (N_23758,N_23158,N_23086);
nand U23759 (N_23759,N_23192,N_23242);
and U23760 (N_23760,N_23392,N_23221);
or U23761 (N_23761,N_23077,N_22898);
and U23762 (N_23762,N_23064,N_23232);
nand U23763 (N_23763,N_23378,N_23106);
and U23764 (N_23764,N_23393,N_22897);
or U23765 (N_23765,N_23361,N_22853);
or U23766 (N_23766,N_23099,N_23184);
nor U23767 (N_23767,N_22881,N_23311);
nand U23768 (N_23768,N_23326,N_23075);
and U23769 (N_23769,N_22877,N_23071);
and U23770 (N_23770,N_22884,N_23047);
or U23771 (N_23771,N_23319,N_22955);
nand U23772 (N_23772,N_23132,N_23030);
nand U23773 (N_23773,N_23114,N_22849);
and U23774 (N_23774,N_22842,N_22932);
nand U23775 (N_23775,N_23091,N_23117);
nand U23776 (N_23776,N_23232,N_22883);
nand U23777 (N_23777,N_22895,N_22983);
nor U23778 (N_23778,N_23024,N_23383);
and U23779 (N_23779,N_23087,N_23042);
nor U23780 (N_23780,N_23217,N_22991);
or U23781 (N_23781,N_23348,N_23364);
nand U23782 (N_23782,N_23110,N_23185);
or U23783 (N_23783,N_23289,N_23020);
and U23784 (N_23784,N_22991,N_23204);
nor U23785 (N_23785,N_22993,N_22843);
and U23786 (N_23786,N_23036,N_23215);
nand U23787 (N_23787,N_22989,N_23193);
nand U23788 (N_23788,N_23133,N_23183);
or U23789 (N_23789,N_23394,N_23389);
or U23790 (N_23790,N_23198,N_22913);
and U23791 (N_23791,N_22828,N_23160);
or U23792 (N_23792,N_23180,N_23018);
nor U23793 (N_23793,N_22963,N_22937);
nor U23794 (N_23794,N_23271,N_22851);
nand U23795 (N_23795,N_23275,N_23331);
nand U23796 (N_23796,N_23207,N_23209);
nand U23797 (N_23797,N_22816,N_23013);
nor U23798 (N_23798,N_23056,N_23225);
and U23799 (N_23799,N_23159,N_23359);
nand U23800 (N_23800,N_22982,N_22973);
nor U23801 (N_23801,N_23224,N_22909);
nand U23802 (N_23802,N_23156,N_23319);
or U23803 (N_23803,N_23013,N_22921);
or U23804 (N_23804,N_22879,N_22903);
nand U23805 (N_23805,N_23323,N_23064);
or U23806 (N_23806,N_23184,N_23117);
nand U23807 (N_23807,N_22916,N_22864);
nand U23808 (N_23808,N_22912,N_23006);
nand U23809 (N_23809,N_23388,N_22943);
or U23810 (N_23810,N_23379,N_23037);
nand U23811 (N_23811,N_23151,N_22987);
or U23812 (N_23812,N_22948,N_22893);
and U23813 (N_23813,N_23000,N_22976);
xor U23814 (N_23814,N_22982,N_22800);
and U23815 (N_23815,N_23184,N_23239);
nor U23816 (N_23816,N_23001,N_22884);
and U23817 (N_23817,N_23066,N_23008);
nand U23818 (N_23818,N_23311,N_22885);
xor U23819 (N_23819,N_23259,N_23216);
and U23820 (N_23820,N_22910,N_23180);
or U23821 (N_23821,N_23135,N_22820);
nand U23822 (N_23822,N_23341,N_22903);
and U23823 (N_23823,N_23054,N_22823);
nand U23824 (N_23824,N_23192,N_23236);
nand U23825 (N_23825,N_22819,N_23123);
nand U23826 (N_23826,N_23313,N_23250);
nor U23827 (N_23827,N_23040,N_22834);
and U23828 (N_23828,N_23372,N_22917);
xor U23829 (N_23829,N_23112,N_23275);
or U23830 (N_23830,N_23293,N_22875);
nand U23831 (N_23831,N_22800,N_23058);
or U23832 (N_23832,N_23226,N_23001);
or U23833 (N_23833,N_22999,N_23107);
and U23834 (N_23834,N_23242,N_23377);
and U23835 (N_23835,N_23285,N_23207);
nand U23836 (N_23836,N_23244,N_23131);
nor U23837 (N_23837,N_23023,N_23212);
nand U23838 (N_23838,N_23372,N_23122);
or U23839 (N_23839,N_22837,N_22847);
or U23840 (N_23840,N_23174,N_23167);
nor U23841 (N_23841,N_23069,N_23232);
or U23842 (N_23842,N_23230,N_22997);
and U23843 (N_23843,N_23132,N_23094);
or U23844 (N_23844,N_23213,N_23067);
nand U23845 (N_23845,N_23156,N_23061);
or U23846 (N_23846,N_23335,N_23330);
and U23847 (N_23847,N_22869,N_22936);
or U23848 (N_23848,N_22810,N_23197);
nor U23849 (N_23849,N_23153,N_23333);
nand U23850 (N_23850,N_23114,N_23207);
and U23851 (N_23851,N_23031,N_23178);
and U23852 (N_23852,N_23128,N_22948);
nor U23853 (N_23853,N_23061,N_23391);
nor U23854 (N_23854,N_23028,N_22941);
xor U23855 (N_23855,N_22858,N_22866);
and U23856 (N_23856,N_23349,N_22812);
or U23857 (N_23857,N_23330,N_23336);
nand U23858 (N_23858,N_23133,N_23121);
or U23859 (N_23859,N_22824,N_23191);
or U23860 (N_23860,N_22929,N_22851);
or U23861 (N_23861,N_22859,N_23135);
and U23862 (N_23862,N_23230,N_23248);
and U23863 (N_23863,N_22937,N_23061);
nand U23864 (N_23864,N_23377,N_22969);
nor U23865 (N_23865,N_23130,N_23103);
and U23866 (N_23866,N_22829,N_23072);
nor U23867 (N_23867,N_23307,N_23150);
and U23868 (N_23868,N_23186,N_22840);
and U23869 (N_23869,N_23046,N_22892);
nand U23870 (N_23870,N_23246,N_23049);
and U23871 (N_23871,N_23198,N_22944);
nor U23872 (N_23872,N_23323,N_23137);
nand U23873 (N_23873,N_23326,N_22801);
or U23874 (N_23874,N_22904,N_23243);
xor U23875 (N_23875,N_22891,N_23024);
or U23876 (N_23876,N_22947,N_23176);
nand U23877 (N_23877,N_23254,N_23211);
nor U23878 (N_23878,N_23162,N_23226);
and U23879 (N_23879,N_23260,N_23127);
nand U23880 (N_23880,N_23176,N_23324);
and U23881 (N_23881,N_22958,N_22928);
nor U23882 (N_23882,N_23161,N_23326);
or U23883 (N_23883,N_22977,N_23043);
nor U23884 (N_23884,N_22953,N_23318);
nand U23885 (N_23885,N_22804,N_22824);
nor U23886 (N_23886,N_23055,N_23285);
nor U23887 (N_23887,N_23374,N_22967);
and U23888 (N_23888,N_23296,N_23331);
and U23889 (N_23889,N_22893,N_22822);
nand U23890 (N_23890,N_22891,N_23378);
and U23891 (N_23891,N_23021,N_22909);
nor U23892 (N_23892,N_23119,N_23347);
nor U23893 (N_23893,N_23018,N_22882);
or U23894 (N_23894,N_23237,N_23016);
or U23895 (N_23895,N_22844,N_23113);
and U23896 (N_23896,N_22879,N_23184);
nor U23897 (N_23897,N_23123,N_23201);
or U23898 (N_23898,N_22893,N_22875);
or U23899 (N_23899,N_22832,N_23248);
and U23900 (N_23900,N_22923,N_23213);
nor U23901 (N_23901,N_22957,N_23009);
and U23902 (N_23902,N_23245,N_23194);
and U23903 (N_23903,N_23253,N_23376);
or U23904 (N_23904,N_23369,N_23373);
nand U23905 (N_23905,N_22857,N_22800);
or U23906 (N_23906,N_23081,N_22886);
or U23907 (N_23907,N_22817,N_22905);
nand U23908 (N_23908,N_23194,N_23262);
nand U23909 (N_23909,N_22890,N_23103);
and U23910 (N_23910,N_23089,N_23371);
and U23911 (N_23911,N_23144,N_22887);
nand U23912 (N_23912,N_22822,N_22987);
nand U23913 (N_23913,N_22909,N_23099);
xor U23914 (N_23914,N_23059,N_23280);
and U23915 (N_23915,N_22926,N_23065);
nand U23916 (N_23916,N_23026,N_23116);
and U23917 (N_23917,N_23326,N_23287);
and U23918 (N_23918,N_23284,N_22944);
nand U23919 (N_23919,N_23080,N_23067);
or U23920 (N_23920,N_23236,N_23137);
nor U23921 (N_23921,N_22850,N_23075);
nor U23922 (N_23922,N_22801,N_22852);
and U23923 (N_23923,N_22907,N_23217);
or U23924 (N_23924,N_23367,N_23069);
nand U23925 (N_23925,N_22917,N_23131);
and U23926 (N_23926,N_23242,N_23337);
nor U23927 (N_23927,N_22973,N_22815);
nand U23928 (N_23928,N_23082,N_23219);
nand U23929 (N_23929,N_22860,N_22957);
or U23930 (N_23930,N_23350,N_22863);
or U23931 (N_23931,N_22990,N_23059);
and U23932 (N_23932,N_23354,N_22861);
or U23933 (N_23933,N_22826,N_23334);
or U23934 (N_23934,N_23339,N_22886);
nor U23935 (N_23935,N_23380,N_22955);
and U23936 (N_23936,N_22890,N_23106);
nand U23937 (N_23937,N_23133,N_23278);
or U23938 (N_23938,N_23070,N_23260);
nor U23939 (N_23939,N_23254,N_23105);
or U23940 (N_23940,N_22864,N_22841);
or U23941 (N_23941,N_23067,N_22861);
and U23942 (N_23942,N_23260,N_22846);
and U23943 (N_23943,N_23289,N_22886);
and U23944 (N_23944,N_22853,N_23166);
nor U23945 (N_23945,N_23355,N_22941);
nor U23946 (N_23946,N_23196,N_23076);
nor U23947 (N_23947,N_23158,N_23283);
nor U23948 (N_23948,N_23389,N_23338);
nor U23949 (N_23949,N_22880,N_23186);
nor U23950 (N_23950,N_22832,N_22836);
nor U23951 (N_23951,N_22930,N_23090);
nand U23952 (N_23952,N_23283,N_23120);
and U23953 (N_23953,N_23096,N_23186);
and U23954 (N_23954,N_22868,N_22984);
and U23955 (N_23955,N_23173,N_23265);
nand U23956 (N_23956,N_23274,N_23048);
and U23957 (N_23957,N_23150,N_22895);
and U23958 (N_23958,N_23057,N_23106);
xor U23959 (N_23959,N_23177,N_23142);
and U23960 (N_23960,N_23126,N_23397);
nand U23961 (N_23961,N_23123,N_22925);
nor U23962 (N_23962,N_23155,N_23216);
or U23963 (N_23963,N_22974,N_23321);
and U23964 (N_23964,N_23307,N_22816);
or U23965 (N_23965,N_22837,N_23013);
nand U23966 (N_23966,N_23114,N_22981);
nand U23967 (N_23967,N_23146,N_22827);
or U23968 (N_23968,N_23255,N_23029);
or U23969 (N_23969,N_23038,N_23372);
and U23970 (N_23970,N_23199,N_23046);
or U23971 (N_23971,N_22926,N_22859);
and U23972 (N_23972,N_23232,N_23181);
nor U23973 (N_23973,N_22910,N_23068);
and U23974 (N_23974,N_22918,N_23310);
nor U23975 (N_23975,N_23146,N_23217);
or U23976 (N_23976,N_23246,N_23132);
nand U23977 (N_23977,N_23360,N_23254);
nor U23978 (N_23978,N_22845,N_23028);
and U23979 (N_23979,N_23067,N_23012);
nand U23980 (N_23980,N_22949,N_22992);
and U23981 (N_23981,N_23039,N_22914);
nand U23982 (N_23982,N_23255,N_23105);
and U23983 (N_23983,N_22875,N_22998);
or U23984 (N_23984,N_23238,N_23039);
nor U23985 (N_23985,N_22888,N_22861);
nand U23986 (N_23986,N_23383,N_23304);
and U23987 (N_23987,N_23233,N_22853);
and U23988 (N_23988,N_23128,N_22944);
nand U23989 (N_23989,N_23216,N_23023);
and U23990 (N_23990,N_22847,N_23000);
xor U23991 (N_23991,N_22900,N_22968);
xor U23992 (N_23992,N_22943,N_22951);
nand U23993 (N_23993,N_22911,N_22986);
or U23994 (N_23994,N_23114,N_23082);
and U23995 (N_23995,N_22995,N_22842);
and U23996 (N_23996,N_23205,N_23177);
and U23997 (N_23997,N_23330,N_23185);
or U23998 (N_23998,N_23303,N_22963);
or U23999 (N_23999,N_23107,N_22973);
or U24000 (N_24000,N_23812,N_23536);
or U24001 (N_24001,N_23652,N_23571);
nand U24002 (N_24002,N_23718,N_23809);
or U24003 (N_24003,N_23522,N_23727);
nor U24004 (N_24004,N_23725,N_23649);
nand U24005 (N_24005,N_23963,N_23676);
and U24006 (N_24006,N_23885,N_23816);
or U24007 (N_24007,N_23712,N_23710);
nand U24008 (N_24008,N_23513,N_23547);
or U24009 (N_24009,N_23528,N_23716);
or U24010 (N_24010,N_23577,N_23913);
nor U24011 (N_24011,N_23616,N_23978);
and U24012 (N_24012,N_23987,N_23926);
nand U24013 (N_24013,N_23484,N_23793);
nand U24014 (N_24014,N_23975,N_23824);
nor U24015 (N_24015,N_23455,N_23500);
nand U24016 (N_24016,N_23803,N_23935);
or U24017 (N_24017,N_23944,N_23559);
and U24018 (N_24018,N_23655,N_23554);
nand U24019 (N_24019,N_23686,N_23863);
nand U24020 (N_24020,N_23767,N_23411);
nor U24021 (N_24021,N_23465,N_23674);
xnor U24022 (N_24022,N_23921,N_23900);
nand U24023 (N_24023,N_23423,N_23908);
nor U24024 (N_24024,N_23589,N_23432);
and U24025 (N_24025,N_23949,N_23651);
xnor U24026 (N_24026,N_23928,N_23830);
or U24027 (N_24027,N_23808,N_23731);
or U24028 (N_24028,N_23879,N_23805);
nor U24029 (N_24029,N_23988,N_23499);
and U24030 (N_24030,N_23592,N_23737);
and U24031 (N_24031,N_23877,N_23740);
or U24032 (N_24032,N_23886,N_23779);
and U24033 (N_24033,N_23508,N_23562);
and U24034 (N_24034,N_23498,N_23807);
nor U24035 (N_24035,N_23929,N_23497);
nor U24036 (N_24036,N_23580,N_23504);
and U24037 (N_24037,N_23622,N_23845);
nor U24038 (N_24038,N_23843,N_23736);
or U24039 (N_24039,N_23626,N_23524);
or U24040 (N_24040,N_23704,N_23448);
or U24041 (N_24041,N_23873,N_23797);
nor U24042 (N_24042,N_23694,N_23867);
nor U24043 (N_24043,N_23685,N_23990);
nor U24044 (N_24044,N_23770,N_23532);
or U24045 (N_24045,N_23839,N_23996);
nor U24046 (N_24046,N_23678,N_23550);
nand U24047 (N_24047,N_23695,N_23683);
and U24048 (N_24048,N_23857,N_23855);
xor U24049 (N_24049,N_23438,N_23410);
nand U24050 (N_24050,N_23569,N_23958);
nor U24051 (N_24051,N_23614,N_23478);
and U24052 (N_24052,N_23897,N_23980);
nor U24053 (N_24053,N_23464,N_23720);
nand U24054 (N_24054,N_23822,N_23777);
or U24055 (N_24055,N_23837,N_23623);
and U24056 (N_24056,N_23682,N_23454);
nor U24057 (N_24057,N_23675,N_23881);
nor U24058 (N_24058,N_23565,N_23466);
or U24059 (N_24059,N_23692,N_23766);
and U24060 (N_24060,N_23851,N_23875);
nand U24061 (N_24061,N_23435,N_23653);
nor U24062 (N_24062,N_23968,N_23989);
and U24063 (N_24063,N_23708,N_23880);
nor U24064 (N_24064,N_23775,N_23768);
nand U24065 (N_24065,N_23818,N_23733);
and U24066 (N_24066,N_23788,N_23630);
or U24067 (N_24067,N_23892,N_23742);
nor U24068 (N_24068,N_23890,N_23514);
or U24069 (N_24069,N_23907,N_23756);
or U24070 (N_24070,N_23889,N_23539);
or U24071 (N_24071,N_23611,N_23638);
nor U24072 (N_24072,N_23861,N_23677);
or U24073 (N_24073,N_23858,N_23995);
nand U24074 (N_24074,N_23505,N_23599);
or U24075 (N_24075,N_23888,N_23691);
nor U24076 (N_24076,N_23939,N_23531);
nand U24077 (N_24077,N_23488,N_23525);
nor U24078 (N_24078,N_23546,N_23759);
nand U24079 (N_24079,N_23799,N_23431);
and U24080 (N_24080,N_23463,N_23956);
nand U24081 (N_24081,N_23841,N_23801);
and U24082 (N_24082,N_23673,N_23933);
nor U24083 (N_24083,N_23705,N_23717);
nor U24084 (N_24084,N_23896,N_23869);
nor U24085 (N_24085,N_23934,N_23507);
nor U24086 (N_24086,N_23575,N_23729);
or U24087 (N_24087,N_23456,N_23937);
xnor U24088 (N_24088,N_23671,N_23699);
and U24089 (N_24089,N_23610,N_23631);
nand U24090 (N_24090,N_23428,N_23607);
nand U24091 (N_24091,N_23475,N_23648);
nor U24092 (N_24092,N_23986,N_23998);
nand U24093 (N_24093,N_23574,N_23474);
or U24094 (N_24094,N_23922,N_23954);
nor U24095 (N_24095,N_23615,N_23780);
or U24096 (N_24096,N_23840,N_23621);
or U24097 (N_24097,N_23693,N_23506);
nand U24098 (N_24098,N_23865,N_23723);
nor U24099 (N_24099,N_23483,N_23407);
nand U24100 (N_24100,N_23469,N_23810);
or U24101 (N_24101,N_23821,N_23625);
nor U24102 (N_24102,N_23590,N_23871);
and U24103 (N_24103,N_23608,N_23931);
nand U24104 (N_24104,N_23715,N_23600);
and U24105 (N_24105,N_23602,N_23591);
or U24106 (N_24106,N_23472,N_23519);
xor U24107 (N_24107,N_23859,N_23595);
or U24108 (N_24108,N_23635,N_23834);
and U24109 (N_24109,N_23643,N_23618);
or U24110 (N_24110,N_23534,N_23923);
nor U24111 (N_24111,N_23526,N_23702);
nor U24112 (N_24112,N_23510,N_23650);
nand U24113 (N_24113,N_23434,N_23482);
xnor U24114 (N_24114,N_23751,N_23530);
or U24115 (N_24115,N_23835,N_23919);
nand U24116 (N_24116,N_23771,N_23960);
nand U24117 (N_24117,N_23932,N_23620);
or U24118 (N_24118,N_23870,N_23558);
and U24119 (N_24119,N_23427,N_23952);
and U24120 (N_24120,N_23814,N_23669);
nand U24121 (N_24121,N_23420,N_23884);
nand U24122 (N_24122,N_23874,N_23953);
nor U24123 (N_24123,N_23906,N_23412);
nor U24124 (N_24124,N_23951,N_23785);
nand U24125 (N_24125,N_23860,N_23838);
xnor U24126 (N_24126,N_23493,N_23690);
or U24127 (N_24127,N_23417,N_23862);
or U24128 (N_24128,N_23582,N_23537);
or U24129 (N_24129,N_23452,N_23645);
or U24130 (N_24130,N_23624,N_23772);
nor U24131 (N_24131,N_23430,N_23490);
or U24132 (N_24132,N_23533,N_23647);
and U24133 (N_24133,N_23979,N_23882);
and U24134 (N_24134,N_23656,N_23741);
or U24135 (N_24135,N_23698,N_23509);
nand U24136 (N_24136,N_23627,N_23786);
nor U24137 (N_24137,N_23854,N_23992);
nand U24138 (N_24138,N_23750,N_23480);
or U24139 (N_24139,N_23829,N_23403);
nand U24140 (N_24140,N_23898,N_23981);
nand U24141 (N_24141,N_23902,N_23658);
and U24142 (N_24142,N_23422,N_23557);
nand U24143 (N_24143,N_23872,N_23585);
nand U24144 (N_24144,N_23703,N_23548);
nand U24145 (N_24145,N_23878,N_23802);
and U24146 (N_24146,N_23847,N_23549);
nor U24147 (N_24147,N_23903,N_23588);
or U24148 (N_24148,N_23706,N_23637);
nand U24149 (N_24149,N_23846,N_23660);
and U24150 (N_24150,N_23852,N_23947);
or U24151 (N_24151,N_23689,N_23564);
and U24152 (N_24152,N_23697,N_23665);
or U24153 (N_24153,N_23769,N_23450);
and U24154 (N_24154,N_23713,N_23844);
nor U24155 (N_24155,N_23568,N_23991);
nor U24156 (N_24156,N_23617,N_23666);
and U24157 (N_24157,N_23918,N_23494);
nor U24158 (N_24158,N_23856,N_23468);
nor U24159 (N_24159,N_23762,N_23485);
nand U24160 (N_24160,N_23798,N_23925);
nand U24161 (N_24161,N_23601,N_23603);
and U24162 (N_24162,N_23664,N_23481);
nand U24163 (N_24163,N_23778,N_23982);
and U24164 (N_24164,N_23700,N_23940);
or U24165 (N_24165,N_23680,N_23842);
nor U24166 (N_24166,N_23701,N_23811);
nand U24167 (N_24167,N_23924,N_23942);
and U24168 (N_24168,N_23738,N_23722);
and U24169 (N_24169,N_23535,N_23899);
nor U24170 (N_24170,N_23429,N_23911);
and U24171 (N_24171,N_23609,N_23679);
or U24172 (N_24172,N_23804,N_23632);
or U24173 (N_24173,N_23629,N_23447);
nand U24174 (N_24174,N_23787,N_23901);
nand U24175 (N_24175,N_23439,N_23583);
nand U24176 (N_24176,N_23728,N_23806);
nor U24177 (N_24177,N_23521,N_23781);
and U24178 (N_24178,N_23789,N_23512);
nand U24179 (N_24179,N_23761,N_23795);
nor U24180 (N_24180,N_23409,N_23467);
and U24181 (N_24181,N_23634,N_23572);
nand U24182 (N_24182,N_23753,N_23401);
or U24183 (N_24183,N_23776,N_23819);
or U24184 (N_24184,N_23461,N_23644);
and U24185 (N_24185,N_23477,N_23560);
or U24186 (N_24186,N_23419,N_23628);
and U24187 (N_24187,N_23416,N_23749);
or U24188 (N_24188,N_23985,N_23437);
nor U24189 (N_24189,N_23576,N_23791);
xnor U24190 (N_24190,N_23966,N_23556);
or U24191 (N_24191,N_23764,N_23421);
and U24192 (N_24192,N_23579,N_23408);
and U24193 (N_24193,N_23540,N_23910);
and U24194 (N_24194,N_23544,N_23605);
nor U24195 (N_24195,N_23760,N_23486);
and U24196 (N_24196,N_23983,N_23523);
and U24197 (N_24197,N_23612,N_23894);
and U24198 (N_24198,N_23654,N_23684);
nor U24199 (N_24199,N_23883,N_23646);
or U24200 (N_24200,N_23948,N_23470);
nor U24201 (N_24201,N_23783,N_23520);
nand U24202 (N_24202,N_23492,N_23459);
nor U24203 (N_24203,N_23545,N_23529);
or U24204 (N_24204,N_23440,N_23551);
or U24205 (N_24205,N_23613,N_23709);
and U24206 (N_24206,N_23938,N_23891);
and U24207 (N_24207,N_23657,N_23849);
nor U24208 (N_24208,N_23425,N_23688);
and U24209 (N_24209,N_23578,N_23971);
nand U24210 (N_24210,N_23593,N_23977);
nor U24211 (N_24211,N_23543,N_23441);
and U24212 (N_24212,N_23471,N_23414);
or U24213 (N_24213,N_23792,N_23825);
and U24214 (N_24214,N_23972,N_23426);
and U24215 (N_24215,N_23445,N_23920);
nor U24216 (N_24216,N_23730,N_23502);
nor U24217 (N_24217,N_23604,N_23476);
and U24218 (N_24218,N_23946,N_23827);
or U24219 (N_24219,N_23541,N_23866);
nor U24220 (N_24220,N_23587,N_23823);
xor U24221 (N_24221,N_23436,N_23491);
nor U24222 (N_24222,N_23916,N_23517);
nand U24223 (N_24223,N_23570,N_23744);
and U24224 (N_24224,N_23831,N_23893);
and U24225 (N_24225,N_23959,N_23670);
nand U24226 (N_24226,N_23501,N_23941);
or U24227 (N_24227,N_23681,N_23739);
and U24228 (N_24228,N_23784,N_23999);
nand U24229 (N_24229,N_23487,N_23909);
and U24230 (N_24230,N_23668,N_23553);
or U24231 (N_24231,N_23406,N_23765);
nor U24232 (N_24232,N_23561,N_23443);
nand U24233 (N_24233,N_23790,N_23433);
nor U24234 (N_24234,N_23976,N_23662);
nor U24235 (N_24235,N_23826,N_23489);
nand U24236 (N_24236,N_23997,N_23479);
nand U24237 (N_24237,N_23813,N_23573);
xor U24238 (N_24238,N_23538,N_23763);
nor U24239 (N_24239,N_23415,N_23404);
or U24240 (N_24240,N_23915,N_23917);
and U24241 (N_24241,N_23503,N_23828);
nand U24242 (N_24242,N_23597,N_23950);
nor U24243 (N_24243,N_23967,N_23596);
and U24244 (N_24244,N_23927,N_23796);
and U24245 (N_24245,N_23773,N_23735);
nor U24246 (N_24246,N_23955,N_23418);
nand U24247 (N_24247,N_23453,N_23707);
nor U24248 (N_24248,N_23904,N_23748);
and U24249 (N_24249,N_23800,N_23930);
nand U24250 (N_24250,N_23672,N_23598);
or U24251 (N_24251,N_23758,N_23965);
nand U24252 (N_24252,N_23914,N_23640);
and U24253 (N_24253,N_23659,N_23451);
nand U24254 (N_24254,N_23757,N_23462);
nand U24255 (N_24255,N_23460,N_23444);
and U24256 (N_24256,N_23782,N_23405);
xor U24257 (N_24257,N_23853,N_23721);
or U24258 (N_24258,N_23711,N_23876);
and U24259 (N_24259,N_23974,N_23639);
and U24260 (N_24260,N_23732,N_23957);
nand U24261 (N_24261,N_23794,N_23912);
and U24262 (N_24262,N_23868,N_23518);
nor U24263 (N_24263,N_23400,N_23567);
nand U24264 (N_24264,N_23719,N_23636);
and U24265 (N_24265,N_23815,N_23446);
nand U24266 (N_24266,N_23943,N_23754);
nor U24267 (N_24267,N_23642,N_23973);
or U24268 (N_24268,N_23542,N_23848);
or U24269 (N_24269,N_23936,N_23495);
and U24270 (N_24270,N_23864,N_23850);
or U24271 (N_24271,N_23619,N_23402);
nand U24272 (N_24272,N_23993,N_23726);
or U24273 (N_24273,N_23887,N_23752);
nand U24274 (N_24274,N_23516,N_23641);
or U24275 (N_24275,N_23515,N_23687);
nor U24276 (N_24276,N_23566,N_23442);
nor U24277 (N_24277,N_23961,N_23970);
and U24278 (N_24278,N_23606,N_23745);
nor U24279 (N_24279,N_23836,N_23633);
and U24280 (N_24280,N_23584,N_23555);
and U24281 (N_24281,N_23746,N_23774);
or U24282 (N_24282,N_23449,N_23969);
and U24283 (N_24283,N_23424,N_23511);
nor U24284 (N_24284,N_23994,N_23895);
nor U24285 (N_24285,N_23663,N_23905);
or U24286 (N_24286,N_23984,N_23527);
nand U24287 (N_24287,N_23755,N_23714);
nor U24288 (N_24288,N_23964,N_23747);
xnor U24289 (N_24289,N_23586,N_23581);
and U24290 (N_24290,N_23945,N_23743);
nor U24291 (N_24291,N_23496,N_23696);
nor U24292 (N_24292,N_23832,N_23820);
nor U24293 (N_24293,N_23833,N_23962);
nor U24294 (N_24294,N_23734,N_23594);
and U24295 (N_24295,N_23667,N_23473);
nor U24296 (N_24296,N_23563,N_23724);
xnor U24297 (N_24297,N_23661,N_23457);
nand U24298 (N_24298,N_23817,N_23552);
nor U24299 (N_24299,N_23413,N_23458);
nand U24300 (N_24300,N_23860,N_23953);
nor U24301 (N_24301,N_23637,N_23582);
and U24302 (N_24302,N_23617,N_23601);
and U24303 (N_24303,N_23882,N_23884);
and U24304 (N_24304,N_23780,N_23816);
and U24305 (N_24305,N_23637,N_23614);
and U24306 (N_24306,N_23641,N_23475);
and U24307 (N_24307,N_23455,N_23734);
and U24308 (N_24308,N_23750,N_23449);
nand U24309 (N_24309,N_23917,N_23953);
nor U24310 (N_24310,N_23616,N_23976);
nand U24311 (N_24311,N_23924,N_23932);
xnor U24312 (N_24312,N_23967,N_23655);
nor U24313 (N_24313,N_23499,N_23408);
and U24314 (N_24314,N_23582,N_23575);
nor U24315 (N_24315,N_23587,N_23544);
nand U24316 (N_24316,N_23567,N_23554);
or U24317 (N_24317,N_23573,N_23876);
nand U24318 (N_24318,N_23527,N_23653);
or U24319 (N_24319,N_23599,N_23485);
nand U24320 (N_24320,N_23433,N_23607);
nor U24321 (N_24321,N_23592,N_23824);
and U24322 (N_24322,N_23694,N_23552);
nor U24323 (N_24323,N_23922,N_23906);
nor U24324 (N_24324,N_23602,N_23500);
nor U24325 (N_24325,N_23736,N_23782);
nor U24326 (N_24326,N_23692,N_23716);
nor U24327 (N_24327,N_23768,N_23509);
or U24328 (N_24328,N_23485,N_23406);
nor U24329 (N_24329,N_23971,N_23908);
and U24330 (N_24330,N_23970,N_23655);
and U24331 (N_24331,N_23873,N_23601);
nor U24332 (N_24332,N_23688,N_23672);
or U24333 (N_24333,N_23503,N_23540);
nand U24334 (N_24334,N_23919,N_23976);
and U24335 (N_24335,N_23780,N_23433);
and U24336 (N_24336,N_23933,N_23753);
nor U24337 (N_24337,N_23436,N_23759);
or U24338 (N_24338,N_23674,N_23878);
nor U24339 (N_24339,N_23504,N_23617);
and U24340 (N_24340,N_23944,N_23453);
or U24341 (N_24341,N_23668,N_23686);
or U24342 (N_24342,N_23625,N_23926);
and U24343 (N_24343,N_23705,N_23762);
or U24344 (N_24344,N_23412,N_23723);
and U24345 (N_24345,N_23631,N_23597);
or U24346 (N_24346,N_23434,N_23469);
nand U24347 (N_24347,N_23620,N_23956);
nor U24348 (N_24348,N_23651,N_23845);
or U24349 (N_24349,N_23404,N_23942);
nand U24350 (N_24350,N_23855,N_23436);
and U24351 (N_24351,N_23613,N_23694);
and U24352 (N_24352,N_23482,N_23436);
and U24353 (N_24353,N_23763,N_23592);
and U24354 (N_24354,N_23706,N_23752);
nor U24355 (N_24355,N_23715,N_23949);
nor U24356 (N_24356,N_23843,N_23608);
and U24357 (N_24357,N_23804,N_23762);
or U24358 (N_24358,N_23673,N_23847);
nand U24359 (N_24359,N_23946,N_23480);
and U24360 (N_24360,N_23753,N_23452);
or U24361 (N_24361,N_23554,N_23573);
nor U24362 (N_24362,N_23626,N_23899);
nand U24363 (N_24363,N_23887,N_23840);
and U24364 (N_24364,N_23559,N_23519);
nand U24365 (N_24365,N_23548,N_23649);
or U24366 (N_24366,N_23619,N_23941);
or U24367 (N_24367,N_23689,N_23707);
or U24368 (N_24368,N_23852,N_23915);
nor U24369 (N_24369,N_23932,N_23868);
nand U24370 (N_24370,N_23672,N_23739);
and U24371 (N_24371,N_23705,N_23615);
and U24372 (N_24372,N_23492,N_23483);
and U24373 (N_24373,N_23449,N_23753);
nand U24374 (N_24374,N_23444,N_23614);
nand U24375 (N_24375,N_23550,N_23419);
nand U24376 (N_24376,N_23494,N_23490);
or U24377 (N_24377,N_23557,N_23655);
and U24378 (N_24378,N_23496,N_23816);
or U24379 (N_24379,N_23701,N_23760);
nand U24380 (N_24380,N_23946,N_23706);
nor U24381 (N_24381,N_23652,N_23958);
or U24382 (N_24382,N_23587,N_23530);
nand U24383 (N_24383,N_23751,N_23840);
and U24384 (N_24384,N_23527,N_23575);
or U24385 (N_24385,N_23735,N_23743);
or U24386 (N_24386,N_23550,N_23474);
or U24387 (N_24387,N_23755,N_23454);
nand U24388 (N_24388,N_23706,N_23527);
and U24389 (N_24389,N_23447,N_23605);
nor U24390 (N_24390,N_23899,N_23865);
nor U24391 (N_24391,N_23758,N_23960);
nor U24392 (N_24392,N_23931,N_23706);
nor U24393 (N_24393,N_23754,N_23550);
nor U24394 (N_24394,N_23656,N_23792);
and U24395 (N_24395,N_23666,N_23761);
nand U24396 (N_24396,N_23799,N_23645);
and U24397 (N_24397,N_23729,N_23428);
or U24398 (N_24398,N_23619,N_23686);
and U24399 (N_24399,N_23650,N_23506);
or U24400 (N_24400,N_23848,N_23682);
and U24401 (N_24401,N_23694,N_23408);
nor U24402 (N_24402,N_23958,N_23729);
nor U24403 (N_24403,N_23896,N_23868);
nor U24404 (N_24404,N_23499,N_23473);
or U24405 (N_24405,N_23558,N_23557);
and U24406 (N_24406,N_23918,N_23798);
nand U24407 (N_24407,N_23859,N_23715);
nor U24408 (N_24408,N_23505,N_23444);
nand U24409 (N_24409,N_23420,N_23601);
or U24410 (N_24410,N_23674,N_23409);
xnor U24411 (N_24411,N_23469,N_23647);
and U24412 (N_24412,N_23908,N_23731);
nand U24413 (N_24413,N_23790,N_23905);
nand U24414 (N_24414,N_23841,N_23551);
nand U24415 (N_24415,N_23982,N_23411);
nor U24416 (N_24416,N_23913,N_23601);
and U24417 (N_24417,N_23502,N_23605);
and U24418 (N_24418,N_23446,N_23957);
and U24419 (N_24419,N_23810,N_23776);
or U24420 (N_24420,N_23560,N_23667);
nand U24421 (N_24421,N_23574,N_23769);
or U24422 (N_24422,N_23894,N_23433);
nor U24423 (N_24423,N_23794,N_23722);
or U24424 (N_24424,N_23592,N_23801);
nor U24425 (N_24425,N_23745,N_23712);
nor U24426 (N_24426,N_23533,N_23430);
or U24427 (N_24427,N_23579,N_23470);
nor U24428 (N_24428,N_23506,N_23507);
nor U24429 (N_24429,N_23804,N_23904);
nand U24430 (N_24430,N_23478,N_23767);
nor U24431 (N_24431,N_23429,N_23481);
nor U24432 (N_24432,N_23771,N_23962);
nor U24433 (N_24433,N_23794,N_23877);
and U24434 (N_24434,N_23753,N_23802);
nor U24435 (N_24435,N_23566,N_23602);
nand U24436 (N_24436,N_23601,N_23507);
or U24437 (N_24437,N_23758,N_23948);
and U24438 (N_24438,N_23773,N_23600);
and U24439 (N_24439,N_23408,N_23452);
or U24440 (N_24440,N_23901,N_23538);
nor U24441 (N_24441,N_23710,N_23990);
and U24442 (N_24442,N_23451,N_23414);
nand U24443 (N_24443,N_23515,N_23954);
or U24444 (N_24444,N_23557,N_23908);
xor U24445 (N_24445,N_23773,N_23968);
nand U24446 (N_24446,N_23894,N_23597);
and U24447 (N_24447,N_23551,N_23427);
nand U24448 (N_24448,N_23677,N_23441);
nor U24449 (N_24449,N_23418,N_23769);
nor U24450 (N_24450,N_23911,N_23590);
or U24451 (N_24451,N_23615,N_23783);
or U24452 (N_24452,N_23578,N_23669);
or U24453 (N_24453,N_23889,N_23928);
or U24454 (N_24454,N_23767,N_23640);
and U24455 (N_24455,N_23956,N_23420);
nand U24456 (N_24456,N_23587,N_23675);
nor U24457 (N_24457,N_23808,N_23462);
and U24458 (N_24458,N_23568,N_23598);
and U24459 (N_24459,N_23831,N_23464);
nor U24460 (N_24460,N_23668,N_23679);
nand U24461 (N_24461,N_23818,N_23674);
or U24462 (N_24462,N_23408,N_23411);
or U24463 (N_24463,N_23941,N_23413);
or U24464 (N_24464,N_23732,N_23955);
or U24465 (N_24465,N_23884,N_23725);
and U24466 (N_24466,N_23733,N_23745);
nor U24467 (N_24467,N_23950,N_23542);
nand U24468 (N_24468,N_23846,N_23664);
or U24469 (N_24469,N_23508,N_23742);
nand U24470 (N_24470,N_23629,N_23571);
nand U24471 (N_24471,N_23954,N_23967);
and U24472 (N_24472,N_23548,N_23962);
nand U24473 (N_24473,N_23688,N_23599);
or U24474 (N_24474,N_23553,N_23783);
nor U24475 (N_24475,N_23827,N_23442);
and U24476 (N_24476,N_23978,N_23416);
or U24477 (N_24477,N_23832,N_23649);
and U24478 (N_24478,N_23509,N_23650);
and U24479 (N_24479,N_23776,N_23620);
and U24480 (N_24480,N_23502,N_23908);
or U24481 (N_24481,N_23609,N_23634);
or U24482 (N_24482,N_23893,N_23789);
nor U24483 (N_24483,N_23502,N_23759);
or U24484 (N_24484,N_23467,N_23426);
and U24485 (N_24485,N_23665,N_23940);
nor U24486 (N_24486,N_23999,N_23795);
and U24487 (N_24487,N_23854,N_23477);
or U24488 (N_24488,N_23752,N_23922);
nor U24489 (N_24489,N_23467,N_23549);
xor U24490 (N_24490,N_23464,N_23494);
or U24491 (N_24491,N_23935,N_23959);
and U24492 (N_24492,N_23874,N_23667);
nand U24493 (N_24493,N_23734,N_23616);
and U24494 (N_24494,N_23781,N_23515);
nand U24495 (N_24495,N_23413,N_23470);
nor U24496 (N_24496,N_23743,N_23781);
or U24497 (N_24497,N_23690,N_23594);
nor U24498 (N_24498,N_23496,N_23673);
nor U24499 (N_24499,N_23586,N_23918);
xor U24500 (N_24500,N_23908,N_23737);
nand U24501 (N_24501,N_23626,N_23429);
nand U24502 (N_24502,N_23761,N_23764);
nor U24503 (N_24503,N_23750,N_23918);
nor U24504 (N_24504,N_23717,N_23534);
or U24505 (N_24505,N_23619,N_23577);
and U24506 (N_24506,N_23452,N_23893);
and U24507 (N_24507,N_23738,N_23713);
and U24508 (N_24508,N_23926,N_23557);
xnor U24509 (N_24509,N_23431,N_23735);
or U24510 (N_24510,N_23710,N_23641);
or U24511 (N_24511,N_23971,N_23721);
or U24512 (N_24512,N_23714,N_23431);
or U24513 (N_24513,N_23610,N_23599);
nor U24514 (N_24514,N_23659,N_23429);
and U24515 (N_24515,N_23880,N_23876);
and U24516 (N_24516,N_23919,N_23400);
nand U24517 (N_24517,N_23896,N_23982);
nor U24518 (N_24518,N_23846,N_23880);
or U24519 (N_24519,N_23870,N_23676);
and U24520 (N_24520,N_23551,N_23647);
nand U24521 (N_24521,N_23863,N_23533);
nand U24522 (N_24522,N_23476,N_23413);
nand U24523 (N_24523,N_23825,N_23897);
nand U24524 (N_24524,N_23513,N_23562);
and U24525 (N_24525,N_23455,N_23532);
and U24526 (N_24526,N_23606,N_23418);
or U24527 (N_24527,N_23521,N_23825);
and U24528 (N_24528,N_23745,N_23477);
or U24529 (N_24529,N_23492,N_23696);
nor U24530 (N_24530,N_23746,N_23704);
or U24531 (N_24531,N_23703,N_23457);
or U24532 (N_24532,N_23731,N_23479);
and U24533 (N_24533,N_23906,N_23762);
or U24534 (N_24534,N_23909,N_23629);
and U24535 (N_24535,N_23479,N_23552);
nor U24536 (N_24536,N_23675,N_23510);
and U24537 (N_24537,N_23825,N_23498);
nand U24538 (N_24538,N_23527,N_23494);
or U24539 (N_24539,N_23479,N_23992);
nor U24540 (N_24540,N_23947,N_23452);
or U24541 (N_24541,N_23730,N_23995);
and U24542 (N_24542,N_23601,N_23423);
or U24543 (N_24543,N_23489,N_23714);
nand U24544 (N_24544,N_23740,N_23716);
nor U24545 (N_24545,N_23874,N_23594);
xnor U24546 (N_24546,N_23498,N_23932);
nor U24547 (N_24547,N_23725,N_23663);
nand U24548 (N_24548,N_23960,N_23621);
and U24549 (N_24549,N_23925,N_23534);
nand U24550 (N_24550,N_23962,N_23762);
and U24551 (N_24551,N_23458,N_23581);
and U24552 (N_24552,N_23845,N_23592);
and U24553 (N_24553,N_23550,N_23746);
or U24554 (N_24554,N_23586,N_23832);
nand U24555 (N_24555,N_23948,N_23789);
nor U24556 (N_24556,N_23433,N_23642);
nor U24557 (N_24557,N_23904,N_23619);
nor U24558 (N_24558,N_23899,N_23534);
xor U24559 (N_24559,N_23920,N_23742);
and U24560 (N_24560,N_23946,N_23551);
or U24561 (N_24561,N_23773,N_23591);
and U24562 (N_24562,N_23826,N_23459);
or U24563 (N_24563,N_23616,N_23523);
and U24564 (N_24564,N_23590,N_23913);
and U24565 (N_24565,N_23867,N_23702);
or U24566 (N_24566,N_23846,N_23710);
or U24567 (N_24567,N_23647,N_23750);
nor U24568 (N_24568,N_23797,N_23552);
and U24569 (N_24569,N_23432,N_23805);
nor U24570 (N_24570,N_23981,N_23978);
or U24571 (N_24571,N_23651,N_23434);
and U24572 (N_24572,N_23646,N_23667);
and U24573 (N_24573,N_23479,N_23475);
xnor U24574 (N_24574,N_23688,N_23890);
and U24575 (N_24575,N_23975,N_23557);
nor U24576 (N_24576,N_23670,N_23632);
nand U24577 (N_24577,N_23433,N_23764);
nor U24578 (N_24578,N_23901,N_23839);
or U24579 (N_24579,N_23978,N_23668);
xnor U24580 (N_24580,N_23603,N_23946);
nand U24581 (N_24581,N_23864,N_23921);
or U24582 (N_24582,N_23885,N_23551);
nand U24583 (N_24583,N_23627,N_23628);
xnor U24584 (N_24584,N_23652,N_23867);
or U24585 (N_24585,N_23802,N_23471);
and U24586 (N_24586,N_23613,N_23914);
nand U24587 (N_24587,N_23554,N_23409);
xor U24588 (N_24588,N_23440,N_23596);
nor U24589 (N_24589,N_23736,N_23881);
nor U24590 (N_24590,N_23601,N_23952);
or U24591 (N_24591,N_23801,N_23849);
or U24592 (N_24592,N_23616,N_23712);
and U24593 (N_24593,N_23613,N_23853);
or U24594 (N_24594,N_23764,N_23521);
and U24595 (N_24595,N_23421,N_23557);
or U24596 (N_24596,N_23569,N_23902);
and U24597 (N_24597,N_23711,N_23618);
or U24598 (N_24598,N_23489,N_23968);
and U24599 (N_24599,N_23446,N_23539);
and U24600 (N_24600,N_24034,N_24598);
or U24601 (N_24601,N_24387,N_24329);
nor U24602 (N_24602,N_24545,N_24564);
and U24603 (N_24603,N_24417,N_24193);
or U24604 (N_24604,N_24420,N_24172);
or U24605 (N_24605,N_24526,N_24064);
nor U24606 (N_24606,N_24406,N_24316);
and U24607 (N_24607,N_24393,N_24135);
and U24608 (N_24608,N_24424,N_24546);
nor U24609 (N_24609,N_24415,N_24250);
and U24610 (N_24610,N_24289,N_24475);
nand U24611 (N_24611,N_24037,N_24515);
nand U24612 (N_24612,N_24043,N_24079);
and U24613 (N_24613,N_24256,N_24480);
and U24614 (N_24614,N_24335,N_24108);
or U24615 (N_24615,N_24371,N_24314);
nor U24616 (N_24616,N_24410,N_24328);
xor U24617 (N_24617,N_24435,N_24476);
xnor U24618 (N_24618,N_24072,N_24436);
nand U24619 (N_24619,N_24584,N_24185);
and U24620 (N_24620,N_24042,N_24096);
or U24621 (N_24621,N_24433,N_24082);
nand U24622 (N_24622,N_24426,N_24565);
or U24623 (N_24623,N_24047,N_24211);
or U24624 (N_24624,N_24178,N_24155);
nor U24625 (N_24625,N_24075,N_24296);
nor U24626 (N_24626,N_24137,N_24209);
nand U24627 (N_24627,N_24257,N_24573);
nand U24628 (N_24628,N_24512,N_24310);
nor U24629 (N_24629,N_24380,N_24482);
or U24630 (N_24630,N_24262,N_24378);
nand U24631 (N_24631,N_24241,N_24498);
nor U24632 (N_24632,N_24114,N_24409);
nor U24633 (N_24633,N_24265,N_24572);
nor U24634 (N_24634,N_24014,N_24098);
nand U24635 (N_24635,N_24418,N_24148);
or U24636 (N_24636,N_24493,N_24499);
or U24637 (N_24637,N_24359,N_24210);
nor U24638 (N_24638,N_24394,N_24116);
and U24639 (N_24639,N_24192,N_24497);
and U24640 (N_24640,N_24428,N_24060);
and U24641 (N_24641,N_24284,N_24143);
or U24642 (N_24642,N_24449,N_24260);
or U24643 (N_24643,N_24491,N_24000);
nor U24644 (N_24644,N_24112,N_24529);
nor U24645 (N_24645,N_24208,N_24212);
nor U24646 (N_24646,N_24366,N_24121);
nand U24647 (N_24647,N_24288,N_24432);
nor U24648 (N_24648,N_24590,N_24005);
nand U24649 (N_24649,N_24245,N_24131);
xor U24650 (N_24650,N_24351,N_24347);
or U24651 (N_24651,N_24050,N_24528);
nand U24652 (N_24652,N_24466,N_24510);
or U24653 (N_24653,N_24074,N_24297);
nor U24654 (N_24654,N_24002,N_24307);
xnor U24655 (N_24655,N_24009,N_24223);
nor U24656 (N_24656,N_24575,N_24246);
or U24657 (N_24657,N_24569,N_24157);
or U24658 (N_24658,N_24599,N_24063);
and U24659 (N_24659,N_24562,N_24225);
nor U24660 (N_24660,N_24059,N_24158);
nand U24661 (N_24661,N_24129,N_24336);
or U24662 (N_24662,N_24083,N_24429);
nor U24663 (N_24663,N_24125,N_24281);
or U24664 (N_24664,N_24219,N_24069);
nand U24665 (N_24665,N_24495,N_24502);
nor U24666 (N_24666,N_24003,N_24441);
nand U24667 (N_24667,N_24474,N_24306);
and U24668 (N_24668,N_24358,N_24081);
nor U24669 (N_24669,N_24031,N_24170);
nor U24670 (N_24670,N_24248,N_24560);
or U24671 (N_24671,N_24293,N_24434);
nand U24672 (N_24672,N_24317,N_24205);
nor U24673 (N_24673,N_24383,N_24066);
or U24674 (N_24674,N_24587,N_24097);
nor U24675 (N_24675,N_24056,N_24032);
and U24676 (N_24676,N_24551,N_24127);
nor U24677 (N_24677,N_24396,N_24117);
nor U24678 (N_24678,N_24091,N_24136);
or U24679 (N_24679,N_24045,N_24525);
nand U24680 (N_24680,N_24222,N_24354);
and U24681 (N_24681,N_24197,N_24001);
nor U24682 (N_24682,N_24176,N_24249);
nor U24683 (N_24683,N_24052,N_24278);
and U24684 (N_24684,N_24574,N_24044);
and U24685 (N_24685,N_24240,N_24386);
nor U24686 (N_24686,N_24544,N_24334);
nand U24687 (N_24687,N_24118,N_24518);
and U24688 (N_24688,N_24038,N_24139);
nand U24689 (N_24689,N_24189,N_24486);
nor U24690 (N_24690,N_24258,N_24403);
and U24691 (N_24691,N_24028,N_24054);
nor U24692 (N_24692,N_24227,N_24389);
or U24693 (N_24693,N_24589,N_24533);
nor U24694 (N_24694,N_24431,N_24279);
and U24695 (N_24695,N_24370,N_24315);
nand U24696 (N_24696,N_24239,N_24244);
nand U24697 (N_24697,N_24101,N_24465);
nand U24698 (N_24698,N_24377,N_24319);
and U24699 (N_24699,N_24352,N_24013);
or U24700 (N_24700,N_24492,N_24110);
and U24701 (N_24701,N_24107,N_24100);
nand U24702 (N_24702,N_24517,N_24472);
nand U24703 (N_24703,N_24468,N_24375);
and U24704 (N_24704,N_24015,N_24065);
and U24705 (N_24705,N_24190,N_24488);
nand U24706 (N_24706,N_24531,N_24164);
nand U24707 (N_24707,N_24312,N_24071);
and U24708 (N_24708,N_24221,N_24168);
nand U24709 (N_24709,N_24411,N_24182);
nor U24710 (N_24710,N_24271,N_24459);
and U24711 (N_24711,N_24215,N_24350);
nand U24712 (N_24712,N_24295,N_24057);
nand U24713 (N_24713,N_24326,N_24412);
and U24714 (N_24714,N_24049,N_24563);
and U24715 (N_24715,N_24594,N_24122);
nor U24716 (N_24716,N_24463,N_24452);
nand U24717 (N_24717,N_24408,N_24151);
and U24718 (N_24718,N_24173,N_24445);
nand U24719 (N_24719,N_24365,N_24089);
nor U24720 (N_24720,N_24458,N_24530);
nor U24721 (N_24721,N_24092,N_24161);
or U24722 (N_24722,N_24030,N_24171);
and U24723 (N_24723,N_24035,N_24355);
nand U24724 (N_24724,N_24552,N_24541);
or U24725 (N_24725,N_24274,N_24280);
nor U24726 (N_24726,N_24140,N_24308);
or U24727 (N_24727,N_24156,N_24166);
nand U24728 (N_24728,N_24179,N_24471);
and U24729 (N_24729,N_24067,N_24453);
or U24730 (N_24730,N_24442,N_24134);
or U24731 (N_24731,N_24163,N_24537);
and U24732 (N_24732,N_24341,N_24174);
or U24733 (N_24733,N_24554,N_24291);
nor U24734 (N_24734,N_24070,N_24450);
or U24735 (N_24735,N_24457,N_24305);
and U24736 (N_24736,N_24017,N_24090);
nor U24737 (N_24737,N_24519,N_24285);
xnor U24738 (N_24738,N_24369,N_24467);
nor U24739 (N_24739,N_24019,N_24099);
nor U24740 (N_24740,N_24373,N_24534);
xnor U24741 (N_24741,N_24016,N_24195);
nand U24742 (N_24742,N_24571,N_24421);
nor U24743 (N_24743,N_24404,N_24202);
nand U24744 (N_24744,N_24327,N_24242);
nand U24745 (N_24745,N_24303,N_24253);
and U24746 (N_24746,N_24356,N_24349);
and U24747 (N_24747,N_24267,N_24299);
nand U24748 (N_24748,N_24124,N_24479);
and U24749 (N_24749,N_24368,N_24400);
nor U24750 (N_24750,N_24093,N_24363);
nor U24751 (N_24751,N_24454,N_24141);
and U24752 (N_24752,N_24167,N_24084);
nand U24753 (N_24753,N_24133,N_24150);
nand U24754 (N_24754,N_24346,N_24376);
xor U24755 (N_24755,N_24496,N_24570);
and U24756 (N_24756,N_24321,N_24128);
nand U24757 (N_24757,N_24029,N_24509);
and U24758 (N_24758,N_24183,N_24577);
or U24759 (N_24759,N_24025,N_24055);
nor U24760 (N_24760,N_24204,N_24439);
nor U24761 (N_24761,N_24180,N_24333);
nand U24762 (N_24762,N_24342,N_24105);
or U24763 (N_24763,N_24588,N_24505);
nor U24764 (N_24764,N_24010,N_24582);
nand U24765 (N_24765,N_24490,N_24581);
and U24766 (N_24766,N_24283,N_24177);
and U24767 (N_24767,N_24460,N_24413);
nand U24768 (N_24768,N_24058,N_24027);
nor U24769 (N_24769,N_24233,N_24224);
nand U24770 (N_24770,N_24448,N_24290);
or U24771 (N_24771,N_24535,N_24251);
and U24772 (N_24772,N_24324,N_24191);
nor U24773 (N_24773,N_24543,N_24111);
nor U24774 (N_24774,N_24444,N_24046);
nor U24775 (N_24775,N_24149,N_24181);
and U24776 (N_24776,N_24578,N_24451);
nand U24777 (N_24777,N_24331,N_24423);
or U24778 (N_24778,N_24007,N_24263);
nor U24779 (N_24779,N_24033,N_24048);
or U24780 (N_24780,N_24304,N_24477);
and U24781 (N_24781,N_24184,N_24523);
and U24782 (N_24782,N_24095,N_24362);
nor U24783 (N_24783,N_24254,N_24547);
nand U24784 (N_24784,N_24591,N_24381);
and U24785 (N_24785,N_24576,N_24536);
nand U24786 (N_24786,N_24238,N_24286);
nor U24787 (N_24787,N_24006,N_24123);
nor U24788 (N_24788,N_24159,N_24275);
nand U24789 (N_24789,N_24372,N_24226);
and U24790 (N_24790,N_24469,N_24447);
or U24791 (N_24791,N_24300,N_24504);
nand U24792 (N_24792,N_24332,N_24313);
nor U24793 (N_24793,N_24548,N_24199);
nor U24794 (N_24794,N_24360,N_24217);
nand U24795 (N_24795,N_24119,N_24367);
or U24796 (N_24796,N_24216,N_24395);
and U24797 (N_24797,N_24154,N_24165);
nand U24798 (N_24798,N_24230,N_24340);
xnor U24799 (N_24799,N_24266,N_24527);
nor U24800 (N_24800,N_24113,N_24021);
nand U24801 (N_24801,N_24388,N_24399);
nor U24802 (N_24802,N_24522,N_24478);
and U24803 (N_24803,N_24322,N_24018);
nor U24804 (N_24804,N_24580,N_24489);
or U24805 (N_24805,N_24061,N_24255);
nand U24806 (N_24806,N_24218,N_24264);
nand U24807 (N_24807,N_24085,N_24115);
nor U24808 (N_24808,N_24203,N_24153);
and U24809 (N_24809,N_24142,N_24485);
and U24810 (N_24810,N_24427,N_24595);
or U24811 (N_24811,N_24464,N_24596);
nand U24812 (N_24812,N_24169,N_24446);
nand U24813 (N_24813,N_24273,N_24501);
nand U24814 (N_24814,N_24540,N_24511);
and U24815 (N_24815,N_24542,N_24068);
nor U24816 (N_24816,N_24138,N_24268);
nor U24817 (N_24817,N_24385,N_24298);
and U24818 (N_24818,N_24053,N_24384);
nor U24819 (N_24819,N_24585,N_24419);
or U24820 (N_24820,N_24126,N_24521);
nand U24821 (N_24821,N_24120,N_24024);
nand U24822 (N_24822,N_24022,N_24344);
and U24823 (N_24823,N_24390,N_24220);
or U24824 (N_24824,N_24259,N_24508);
or U24825 (N_24825,N_24102,N_24586);
nor U24826 (N_24826,N_24483,N_24261);
nand U24827 (N_24827,N_24188,N_24455);
and U24828 (N_24828,N_24077,N_24398);
nor U24829 (N_24829,N_24008,N_24311);
nor U24830 (N_24830,N_24235,N_24555);
nand U24831 (N_24831,N_24301,N_24549);
nand U24832 (N_24832,N_24345,N_24041);
and U24833 (N_24833,N_24382,N_24276);
or U24834 (N_24834,N_24086,N_24532);
and U24835 (N_24835,N_24109,N_24361);
nand U24836 (N_24836,N_24330,N_24391);
or U24837 (N_24837,N_24236,N_24407);
and U24838 (N_24838,N_24513,N_24470);
nand U24839 (N_24839,N_24402,N_24144);
nand U24840 (N_24840,N_24556,N_24080);
and U24841 (N_24841,N_24557,N_24397);
and U24842 (N_24842,N_24073,N_24062);
and U24843 (N_24843,N_24323,N_24287);
and U24844 (N_24844,N_24237,N_24430);
nand U24845 (N_24845,N_24405,N_24198);
or U24846 (N_24846,N_24103,N_24196);
or U24847 (N_24847,N_24186,N_24473);
nand U24848 (N_24848,N_24484,N_24229);
nor U24849 (N_24849,N_24437,N_24036);
or U24850 (N_24850,N_24425,N_24130);
and U24851 (N_24851,N_24520,N_24401);
nand U24852 (N_24852,N_24392,N_24214);
or U24853 (N_24853,N_24106,N_24004);
nand U24854 (N_24854,N_24247,N_24160);
nor U24855 (N_24855,N_24078,N_24539);
nor U24856 (N_24856,N_24011,N_24320);
nor U24857 (N_24857,N_24270,N_24023);
and U24858 (N_24858,N_24087,N_24207);
nor U24859 (N_24859,N_24026,N_24012);
and U24860 (N_24860,N_24558,N_24422);
or U24861 (N_24861,N_24132,N_24088);
and U24862 (N_24862,N_24243,N_24364);
nor U24863 (N_24863,N_24302,N_24272);
nor U24864 (N_24864,N_24213,N_24187);
or U24865 (N_24865,N_24353,N_24559);
or U24866 (N_24866,N_24462,N_24456);
and U24867 (N_24867,N_24553,N_24040);
nor U24868 (N_24868,N_24538,N_24294);
and U24869 (N_24869,N_24162,N_24583);
or U24870 (N_24870,N_24194,N_24147);
nand U24871 (N_24871,N_24597,N_24269);
nor U24872 (N_24872,N_24228,N_24379);
nand U24873 (N_24873,N_24200,N_24343);
and U24874 (N_24874,N_24325,N_24374);
and U24875 (N_24875,N_24524,N_24487);
nand U24876 (N_24876,N_24292,N_24567);
xnor U24877 (N_24877,N_24152,N_24566);
and U24878 (N_24878,N_24104,N_24234);
xnor U24879 (N_24879,N_24592,N_24494);
or U24880 (N_24880,N_24145,N_24039);
nand U24881 (N_24881,N_24094,N_24282);
and U24882 (N_24882,N_24593,N_24206);
or U24883 (N_24883,N_24414,N_24506);
and U24884 (N_24884,N_24416,N_24461);
nor U24885 (N_24885,N_24309,N_24568);
and U24886 (N_24886,N_24438,N_24579);
and U24887 (N_24887,N_24503,N_24561);
nand U24888 (N_24888,N_24277,N_24357);
nand U24889 (N_24889,N_24252,N_24440);
nand U24890 (N_24890,N_24550,N_24507);
nand U24891 (N_24891,N_24175,N_24481);
nor U24892 (N_24892,N_24337,N_24051);
nand U24893 (N_24893,N_24516,N_24514);
or U24894 (N_24894,N_24232,N_24231);
nand U24895 (N_24895,N_24201,N_24146);
and U24896 (N_24896,N_24339,N_24076);
and U24897 (N_24897,N_24318,N_24500);
or U24898 (N_24898,N_24020,N_24338);
and U24899 (N_24899,N_24443,N_24348);
and U24900 (N_24900,N_24356,N_24257);
xnor U24901 (N_24901,N_24122,N_24274);
nand U24902 (N_24902,N_24525,N_24544);
nor U24903 (N_24903,N_24106,N_24245);
and U24904 (N_24904,N_24497,N_24362);
and U24905 (N_24905,N_24320,N_24266);
nand U24906 (N_24906,N_24303,N_24538);
nor U24907 (N_24907,N_24131,N_24288);
or U24908 (N_24908,N_24347,N_24096);
and U24909 (N_24909,N_24313,N_24510);
or U24910 (N_24910,N_24141,N_24028);
nand U24911 (N_24911,N_24069,N_24529);
nand U24912 (N_24912,N_24324,N_24334);
nor U24913 (N_24913,N_24154,N_24349);
nand U24914 (N_24914,N_24384,N_24142);
and U24915 (N_24915,N_24560,N_24258);
or U24916 (N_24916,N_24000,N_24334);
or U24917 (N_24917,N_24005,N_24133);
nand U24918 (N_24918,N_24369,N_24076);
nand U24919 (N_24919,N_24307,N_24137);
nand U24920 (N_24920,N_24496,N_24541);
nor U24921 (N_24921,N_24072,N_24552);
or U24922 (N_24922,N_24542,N_24033);
and U24923 (N_24923,N_24435,N_24272);
nor U24924 (N_24924,N_24353,N_24136);
and U24925 (N_24925,N_24486,N_24317);
nor U24926 (N_24926,N_24578,N_24593);
and U24927 (N_24927,N_24300,N_24469);
nor U24928 (N_24928,N_24423,N_24278);
nor U24929 (N_24929,N_24062,N_24255);
or U24930 (N_24930,N_24306,N_24249);
and U24931 (N_24931,N_24299,N_24294);
xnor U24932 (N_24932,N_24018,N_24459);
or U24933 (N_24933,N_24495,N_24122);
nand U24934 (N_24934,N_24187,N_24384);
nor U24935 (N_24935,N_24336,N_24529);
and U24936 (N_24936,N_24102,N_24152);
and U24937 (N_24937,N_24572,N_24577);
and U24938 (N_24938,N_24263,N_24474);
nand U24939 (N_24939,N_24056,N_24567);
nor U24940 (N_24940,N_24303,N_24234);
or U24941 (N_24941,N_24257,N_24407);
or U24942 (N_24942,N_24069,N_24144);
nand U24943 (N_24943,N_24067,N_24471);
and U24944 (N_24944,N_24587,N_24373);
and U24945 (N_24945,N_24409,N_24346);
and U24946 (N_24946,N_24557,N_24598);
nand U24947 (N_24947,N_24417,N_24127);
or U24948 (N_24948,N_24087,N_24394);
nor U24949 (N_24949,N_24018,N_24072);
nand U24950 (N_24950,N_24528,N_24056);
nand U24951 (N_24951,N_24431,N_24306);
or U24952 (N_24952,N_24306,N_24443);
and U24953 (N_24953,N_24185,N_24122);
nor U24954 (N_24954,N_24046,N_24154);
or U24955 (N_24955,N_24214,N_24156);
and U24956 (N_24956,N_24061,N_24514);
and U24957 (N_24957,N_24377,N_24310);
or U24958 (N_24958,N_24353,N_24519);
xnor U24959 (N_24959,N_24171,N_24584);
and U24960 (N_24960,N_24283,N_24184);
or U24961 (N_24961,N_24397,N_24362);
and U24962 (N_24962,N_24024,N_24315);
nand U24963 (N_24963,N_24190,N_24061);
or U24964 (N_24964,N_24269,N_24438);
and U24965 (N_24965,N_24417,N_24552);
nand U24966 (N_24966,N_24109,N_24481);
and U24967 (N_24967,N_24270,N_24067);
nand U24968 (N_24968,N_24130,N_24482);
xnor U24969 (N_24969,N_24294,N_24065);
and U24970 (N_24970,N_24597,N_24069);
or U24971 (N_24971,N_24267,N_24471);
nor U24972 (N_24972,N_24211,N_24251);
or U24973 (N_24973,N_24170,N_24439);
nor U24974 (N_24974,N_24439,N_24554);
nand U24975 (N_24975,N_24087,N_24019);
nor U24976 (N_24976,N_24004,N_24597);
nor U24977 (N_24977,N_24461,N_24457);
nor U24978 (N_24978,N_24459,N_24316);
or U24979 (N_24979,N_24569,N_24017);
nand U24980 (N_24980,N_24089,N_24045);
nand U24981 (N_24981,N_24048,N_24101);
and U24982 (N_24982,N_24075,N_24496);
xor U24983 (N_24983,N_24029,N_24213);
and U24984 (N_24984,N_24597,N_24165);
or U24985 (N_24985,N_24514,N_24112);
nand U24986 (N_24986,N_24554,N_24572);
or U24987 (N_24987,N_24342,N_24000);
nor U24988 (N_24988,N_24182,N_24105);
and U24989 (N_24989,N_24233,N_24164);
nand U24990 (N_24990,N_24374,N_24306);
nand U24991 (N_24991,N_24107,N_24376);
and U24992 (N_24992,N_24429,N_24586);
nand U24993 (N_24993,N_24456,N_24248);
nor U24994 (N_24994,N_24461,N_24156);
nor U24995 (N_24995,N_24572,N_24400);
or U24996 (N_24996,N_24233,N_24575);
nand U24997 (N_24997,N_24179,N_24223);
and U24998 (N_24998,N_24469,N_24499);
or U24999 (N_24999,N_24295,N_24139);
nand U25000 (N_25000,N_24101,N_24283);
or U25001 (N_25001,N_24552,N_24413);
and U25002 (N_25002,N_24404,N_24311);
nor U25003 (N_25003,N_24138,N_24360);
or U25004 (N_25004,N_24266,N_24550);
nand U25005 (N_25005,N_24228,N_24512);
or U25006 (N_25006,N_24245,N_24371);
and U25007 (N_25007,N_24485,N_24052);
nand U25008 (N_25008,N_24558,N_24410);
nor U25009 (N_25009,N_24463,N_24522);
nand U25010 (N_25010,N_24312,N_24478);
and U25011 (N_25011,N_24193,N_24428);
nor U25012 (N_25012,N_24353,N_24317);
nand U25013 (N_25013,N_24250,N_24082);
or U25014 (N_25014,N_24170,N_24033);
and U25015 (N_25015,N_24059,N_24429);
nand U25016 (N_25016,N_24599,N_24364);
and U25017 (N_25017,N_24518,N_24599);
nor U25018 (N_25018,N_24205,N_24184);
nand U25019 (N_25019,N_24184,N_24448);
and U25020 (N_25020,N_24541,N_24558);
and U25021 (N_25021,N_24410,N_24056);
and U25022 (N_25022,N_24503,N_24443);
nor U25023 (N_25023,N_24037,N_24203);
nand U25024 (N_25024,N_24296,N_24240);
nand U25025 (N_25025,N_24212,N_24278);
and U25026 (N_25026,N_24197,N_24485);
nand U25027 (N_25027,N_24592,N_24511);
nor U25028 (N_25028,N_24107,N_24357);
and U25029 (N_25029,N_24194,N_24167);
nor U25030 (N_25030,N_24568,N_24409);
or U25031 (N_25031,N_24479,N_24552);
and U25032 (N_25032,N_24534,N_24331);
nand U25033 (N_25033,N_24564,N_24524);
or U25034 (N_25034,N_24597,N_24050);
and U25035 (N_25035,N_24531,N_24498);
and U25036 (N_25036,N_24312,N_24108);
or U25037 (N_25037,N_24584,N_24002);
or U25038 (N_25038,N_24567,N_24132);
or U25039 (N_25039,N_24125,N_24353);
and U25040 (N_25040,N_24223,N_24212);
and U25041 (N_25041,N_24522,N_24148);
nand U25042 (N_25042,N_24255,N_24523);
and U25043 (N_25043,N_24367,N_24304);
or U25044 (N_25044,N_24472,N_24026);
nor U25045 (N_25045,N_24184,N_24347);
and U25046 (N_25046,N_24162,N_24556);
nand U25047 (N_25047,N_24055,N_24289);
and U25048 (N_25048,N_24504,N_24427);
and U25049 (N_25049,N_24314,N_24036);
and U25050 (N_25050,N_24284,N_24120);
or U25051 (N_25051,N_24171,N_24493);
and U25052 (N_25052,N_24190,N_24351);
and U25053 (N_25053,N_24540,N_24440);
or U25054 (N_25054,N_24389,N_24477);
nor U25055 (N_25055,N_24372,N_24295);
nand U25056 (N_25056,N_24251,N_24511);
nand U25057 (N_25057,N_24154,N_24315);
or U25058 (N_25058,N_24290,N_24366);
or U25059 (N_25059,N_24523,N_24146);
nand U25060 (N_25060,N_24384,N_24568);
or U25061 (N_25061,N_24437,N_24092);
nor U25062 (N_25062,N_24409,N_24250);
or U25063 (N_25063,N_24516,N_24349);
and U25064 (N_25064,N_24465,N_24236);
nand U25065 (N_25065,N_24129,N_24175);
nand U25066 (N_25066,N_24426,N_24468);
or U25067 (N_25067,N_24218,N_24304);
nand U25068 (N_25068,N_24590,N_24499);
nor U25069 (N_25069,N_24324,N_24146);
and U25070 (N_25070,N_24290,N_24167);
and U25071 (N_25071,N_24584,N_24320);
or U25072 (N_25072,N_24079,N_24526);
or U25073 (N_25073,N_24179,N_24279);
and U25074 (N_25074,N_24117,N_24370);
or U25075 (N_25075,N_24566,N_24293);
nor U25076 (N_25076,N_24320,N_24142);
or U25077 (N_25077,N_24584,N_24510);
and U25078 (N_25078,N_24487,N_24526);
or U25079 (N_25079,N_24030,N_24440);
nor U25080 (N_25080,N_24580,N_24099);
and U25081 (N_25081,N_24292,N_24524);
or U25082 (N_25082,N_24149,N_24596);
and U25083 (N_25083,N_24567,N_24424);
or U25084 (N_25084,N_24065,N_24200);
nor U25085 (N_25085,N_24156,N_24239);
nor U25086 (N_25086,N_24390,N_24089);
and U25087 (N_25087,N_24200,N_24453);
nand U25088 (N_25088,N_24203,N_24147);
and U25089 (N_25089,N_24214,N_24024);
and U25090 (N_25090,N_24288,N_24239);
nor U25091 (N_25091,N_24151,N_24098);
or U25092 (N_25092,N_24127,N_24188);
or U25093 (N_25093,N_24020,N_24385);
and U25094 (N_25094,N_24589,N_24195);
or U25095 (N_25095,N_24305,N_24332);
or U25096 (N_25096,N_24129,N_24299);
nor U25097 (N_25097,N_24426,N_24178);
xnor U25098 (N_25098,N_24477,N_24176);
and U25099 (N_25099,N_24140,N_24115);
nand U25100 (N_25100,N_24342,N_24449);
nor U25101 (N_25101,N_24365,N_24383);
nor U25102 (N_25102,N_24553,N_24032);
nor U25103 (N_25103,N_24380,N_24175);
or U25104 (N_25104,N_24507,N_24217);
nand U25105 (N_25105,N_24279,N_24336);
nand U25106 (N_25106,N_24552,N_24122);
nor U25107 (N_25107,N_24341,N_24356);
and U25108 (N_25108,N_24035,N_24447);
nor U25109 (N_25109,N_24458,N_24136);
nand U25110 (N_25110,N_24543,N_24047);
nand U25111 (N_25111,N_24346,N_24474);
nand U25112 (N_25112,N_24151,N_24211);
or U25113 (N_25113,N_24466,N_24414);
xnor U25114 (N_25114,N_24283,N_24442);
nor U25115 (N_25115,N_24000,N_24241);
and U25116 (N_25116,N_24499,N_24246);
or U25117 (N_25117,N_24341,N_24123);
and U25118 (N_25118,N_24162,N_24486);
or U25119 (N_25119,N_24596,N_24307);
and U25120 (N_25120,N_24550,N_24239);
nor U25121 (N_25121,N_24445,N_24587);
or U25122 (N_25122,N_24439,N_24378);
nor U25123 (N_25123,N_24098,N_24313);
nand U25124 (N_25124,N_24167,N_24358);
nand U25125 (N_25125,N_24314,N_24455);
or U25126 (N_25126,N_24490,N_24579);
and U25127 (N_25127,N_24251,N_24099);
or U25128 (N_25128,N_24430,N_24568);
and U25129 (N_25129,N_24395,N_24248);
and U25130 (N_25130,N_24110,N_24159);
or U25131 (N_25131,N_24255,N_24536);
nor U25132 (N_25132,N_24503,N_24384);
nor U25133 (N_25133,N_24454,N_24336);
or U25134 (N_25134,N_24399,N_24174);
nor U25135 (N_25135,N_24291,N_24199);
and U25136 (N_25136,N_24104,N_24282);
or U25137 (N_25137,N_24506,N_24412);
or U25138 (N_25138,N_24278,N_24597);
or U25139 (N_25139,N_24454,N_24244);
nand U25140 (N_25140,N_24500,N_24416);
nand U25141 (N_25141,N_24456,N_24552);
or U25142 (N_25142,N_24542,N_24408);
and U25143 (N_25143,N_24435,N_24414);
nor U25144 (N_25144,N_24006,N_24526);
xnor U25145 (N_25145,N_24001,N_24265);
nand U25146 (N_25146,N_24497,N_24160);
nand U25147 (N_25147,N_24303,N_24039);
nor U25148 (N_25148,N_24021,N_24164);
and U25149 (N_25149,N_24484,N_24525);
or U25150 (N_25150,N_24363,N_24011);
xor U25151 (N_25151,N_24482,N_24543);
and U25152 (N_25152,N_24073,N_24326);
nand U25153 (N_25153,N_24546,N_24058);
and U25154 (N_25154,N_24397,N_24099);
and U25155 (N_25155,N_24415,N_24360);
nand U25156 (N_25156,N_24497,N_24390);
nand U25157 (N_25157,N_24209,N_24524);
nor U25158 (N_25158,N_24216,N_24436);
nand U25159 (N_25159,N_24393,N_24179);
or U25160 (N_25160,N_24573,N_24289);
nor U25161 (N_25161,N_24249,N_24596);
nand U25162 (N_25162,N_24599,N_24047);
and U25163 (N_25163,N_24478,N_24485);
nor U25164 (N_25164,N_24257,N_24460);
nand U25165 (N_25165,N_24580,N_24593);
and U25166 (N_25166,N_24265,N_24531);
and U25167 (N_25167,N_24596,N_24558);
and U25168 (N_25168,N_24216,N_24084);
nand U25169 (N_25169,N_24585,N_24186);
or U25170 (N_25170,N_24346,N_24444);
or U25171 (N_25171,N_24368,N_24146);
nand U25172 (N_25172,N_24013,N_24417);
and U25173 (N_25173,N_24486,N_24243);
and U25174 (N_25174,N_24120,N_24484);
nand U25175 (N_25175,N_24564,N_24483);
nand U25176 (N_25176,N_24181,N_24110);
and U25177 (N_25177,N_24451,N_24553);
or U25178 (N_25178,N_24133,N_24421);
nand U25179 (N_25179,N_24501,N_24561);
nand U25180 (N_25180,N_24255,N_24429);
or U25181 (N_25181,N_24295,N_24589);
or U25182 (N_25182,N_24160,N_24491);
nor U25183 (N_25183,N_24293,N_24015);
nor U25184 (N_25184,N_24407,N_24341);
nand U25185 (N_25185,N_24314,N_24270);
xnor U25186 (N_25186,N_24348,N_24539);
and U25187 (N_25187,N_24491,N_24531);
or U25188 (N_25188,N_24422,N_24171);
nor U25189 (N_25189,N_24328,N_24150);
nand U25190 (N_25190,N_24416,N_24197);
or U25191 (N_25191,N_24495,N_24227);
nor U25192 (N_25192,N_24202,N_24039);
or U25193 (N_25193,N_24590,N_24419);
nand U25194 (N_25194,N_24568,N_24292);
and U25195 (N_25195,N_24014,N_24008);
and U25196 (N_25196,N_24548,N_24486);
nor U25197 (N_25197,N_24532,N_24489);
and U25198 (N_25198,N_24451,N_24388);
xor U25199 (N_25199,N_24532,N_24531);
or U25200 (N_25200,N_25011,N_25023);
and U25201 (N_25201,N_24751,N_24750);
or U25202 (N_25202,N_24827,N_24730);
nand U25203 (N_25203,N_24996,N_24963);
nand U25204 (N_25204,N_24894,N_24653);
and U25205 (N_25205,N_24676,N_24806);
nor U25206 (N_25206,N_24833,N_24947);
nor U25207 (N_25207,N_25134,N_25091);
nand U25208 (N_25208,N_24747,N_25154);
or U25209 (N_25209,N_24640,N_24921);
nor U25210 (N_25210,N_24993,N_24732);
nand U25211 (N_25211,N_25130,N_25178);
and U25212 (N_25212,N_24717,N_24803);
or U25213 (N_25213,N_24712,N_24883);
or U25214 (N_25214,N_25060,N_24656);
nor U25215 (N_25215,N_24753,N_24848);
nor U25216 (N_25216,N_24805,N_25073);
nand U25217 (N_25217,N_24633,N_24807);
nand U25218 (N_25218,N_24831,N_24877);
and U25219 (N_25219,N_25123,N_24605);
xor U25220 (N_25220,N_24892,N_24957);
and U25221 (N_25221,N_24725,N_24649);
or U25222 (N_25222,N_25009,N_24879);
nor U25223 (N_25223,N_24721,N_24861);
or U25224 (N_25224,N_25152,N_24799);
nor U25225 (N_25225,N_24776,N_24985);
nor U25226 (N_25226,N_24847,N_24853);
nor U25227 (N_25227,N_24771,N_25158);
nand U25228 (N_25228,N_24977,N_24933);
or U25229 (N_25229,N_25160,N_24875);
and U25230 (N_25230,N_24792,N_24772);
xor U25231 (N_25231,N_24723,N_24692);
nor U25232 (N_25232,N_24718,N_24797);
nand U25233 (N_25233,N_24997,N_25197);
or U25234 (N_25234,N_24979,N_24959);
and U25235 (N_25235,N_24785,N_25147);
or U25236 (N_25236,N_24742,N_24667);
xnor U25237 (N_25237,N_24924,N_24919);
or U25238 (N_25238,N_25195,N_24694);
nand U25239 (N_25239,N_24913,N_24629);
nand U25240 (N_25240,N_24800,N_24982);
nand U25241 (N_25241,N_24809,N_24974);
or U25242 (N_25242,N_25029,N_24659);
and U25243 (N_25243,N_24720,N_24737);
nor U25244 (N_25244,N_25078,N_24862);
and U25245 (N_25245,N_25128,N_24691);
and U25246 (N_25246,N_24689,N_24960);
nand U25247 (N_25247,N_24697,N_24948);
and U25248 (N_25248,N_25013,N_24849);
and U25249 (N_25249,N_24609,N_25016);
nand U25250 (N_25250,N_24880,N_25108);
nor U25251 (N_25251,N_24731,N_25040);
or U25252 (N_25252,N_24744,N_25105);
nand U25253 (N_25253,N_24650,N_25021);
nor U25254 (N_25254,N_25099,N_24683);
nand U25255 (N_25255,N_25014,N_25174);
nor U25256 (N_25256,N_25120,N_25006);
nand U25257 (N_25257,N_24829,N_25103);
nand U25258 (N_25258,N_24622,N_24876);
or U25259 (N_25259,N_24617,N_24884);
and U25260 (N_25260,N_25156,N_25141);
nand U25261 (N_25261,N_24930,N_24961);
and U25262 (N_25262,N_24976,N_25140);
or U25263 (N_25263,N_25157,N_24782);
nand U25264 (N_25264,N_25176,N_24600);
nand U25265 (N_25265,N_25070,N_24699);
and U25266 (N_25266,N_24991,N_24830);
or U25267 (N_25267,N_24925,N_24821);
and U25268 (N_25268,N_24678,N_25100);
or U25269 (N_25269,N_25098,N_24802);
nand U25270 (N_25270,N_24845,N_24654);
and U25271 (N_25271,N_24855,N_24860);
or U25272 (N_25272,N_24859,N_24670);
nor U25273 (N_25273,N_24666,N_24873);
nor U25274 (N_25274,N_24752,N_25037);
and U25275 (N_25275,N_25090,N_24872);
or U25276 (N_25276,N_24677,N_25024);
nor U25277 (N_25277,N_25121,N_24675);
nor U25278 (N_25278,N_24901,N_25146);
or U25279 (N_25279,N_25093,N_24625);
nand U25280 (N_25280,N_24614,N_24841);
and U25281 (N_25281,N_24701,N_24906);
and U25282 (N_25282,N_25075,N_24920);
xnor U25283 (N_25283,N_25076,N_24887);
nand U25284 (N_25284,N_25065,N_25153);
or U25285 (N_25285,N_25062,N_24754);
nor U25286 (N_25286,N_25113,N_25072);
or U25287 (N_25287,N_24851,N_25196);
or U25288 (N_25288,N_25018,N_24922);
nor U25289 (N_25289,N_24673,N_25032);
or U25290 (N_25290,N_24763,N_25109);
xnor U25291 (N_25291,N_24994,N_24909);
nand U25292 (N_25292,N_24612,N_24623);
xor U25293 (N_25293,N_25087,N_24888);
nand U25294 (N_25294,N_25181,N_24755);
and U25295 (N_25295,N_24973,N_24932);
or U25296 (N_25296,N_25114,N_24988);
or U25297 (N_25297,N_24634,N_24604);
or U25298 (N_25298,N_25119,N_24828);
nor U25299 (N_25299,N_24607,N_24652);
or U25300 (N_25300,N_24905,N_24885);
and U25301 (N_25301,N_24671,N_25044);
nor U25302 (N_25302,N_25097,N_24890);
or U25303 (N_25303,N_24941,N_24635);
or U25304 (N_25304,N_24601,N_24837);
nor U25305 (N_25305,N_25057,N_24722);
and U25306 (N_25306,N_25186,N_25155);
nor U25307 (N_25307,N_25033,N_25169);
nor U25308 (N_25308,N_24900,N_24955);
nor U25309 (N_25309,N_24990,N_25191);
or U25310 (N_25310,N_24825,N_25194);
or U25311 (N_25311,N_25004,N_24910);
or U25312 (N_25312,N_25061,N_24715);
or U25313 (N_25313,N_24672,N_24714);
nor U25314 (N_25314,N_24708,N_24914);
nand U25315 (N_25315,N_24946,N_24681);
or U25316 (N_25316,N_24713,N_24953);
nand U25317 (N_25317,N_25094,N_25170);
nor U25318 (N_25318,N_25054,N_25089);
nor U25319 (N_25319,N_24679,N_25071);
nor U25320 (N_25320,N_24664,N_25110);
nand U25321 (N_25321,N_24962,N_24857);
nand U25322 (N_25322,N_25095,N_24936);
nor U25323 (N_25323,N_25049,N_24937);
nor U25324 (N_25324,N_24639,N_25126);
nor U25325 (N_25325,N_25167,N_24989);
nand U25326 (N_25326,N_24606,N_25081);
nor U25327 (N_25327,N_24696,N_25086);
nor U25328 (N_25328,N_24964,N_25005);
or U25329 (N_25329,N_25159,N_24661);
and U25330 (N_25330,N_24808,N_24967);
nor U25331 (N_25331,N_24608,N_24844);
or U25332 (N_25332,N_25066,N_24711);
or U25333 (N_25333,N_25106,N_24693);
nand U25334 (N_25334,N_24944,N_24647);
and U25335 (N_25335,N_24646,N_24745);
or U25336 (N_25336,N_25038,N_24835);
nand U25337 (N_25337,N_24868,N_24870);
or U25338 (N_25338,N_25111,N_25080);
and U25339 (N_25339,N_24998,N_25028);
and U25340 (N_25340,N_24655,N_24954);
and U25341 (N_25341,N_24854,N_25041);
and U25342 (N_25342,N_25022,N_24628);
nor U25343 (N_25343,N_24773,N_24891);
or U25344 (N_25344,N_24956,N_24775);
nand U25345 (N_25345,N_24603,N_24602);
nor U25346 (N_25346,N_25188,N_25096);
and U25347 (N_25347,N_24728,N_24810);
and U25348 (N_25348,N_24846,N_25177);
nand U25349 (N_25349,N_25118,N_25046);
or U25350 (N_25350,N_25036,N_24889);
nand U25351 (N_25351,N_24762,N_24686);
or U25352 (N_25352,N_24703,N_24770);
or U25353 (N_25353,N_24758,N_25012);
nand U25354 (N_25354,N_24630,N_24878);
nand U25355 (N_25355,N_24719,N_24724);
nor U25356 (N_25356,N_24984,N_25102);
or U25357 (N_25357,N_24726,N_25162);
and U25358 (N_25358,N_24780,N_24789);
and U25359 (N_25359,N_24934,N_24816);
or U25360 (N_25360,N_24978,N_25035);
or U25361 (N_25361,N_24987,N_24980);
nor U25362 (N_25362,N_25043,N_24918);
nand U25363 (N_25363,N_25165,N_25064);
nand U25364 (N_25364,N_24651,N_25107);
or U25365 (N_25365,N_24644,N_24788);
nor U25366 (N_25366,N_24850,N_25161);
or U25367 (N_25367,N_25144,N_24814);
nand U25368 (N_25368,N_24760,N_25132);
nor U25369 (N_25369,N_25131,N_24995);
and U25370 (N_25370,N_24759,N_24903);
and U25371 (N_25371,N_24838,N_24627);
and U25372 (N_25372,N_25164,N_24923);
and U25373 (N_25373,N_24710,N_25112);
nor U25374 (N_25374,N_25179,N_24779);
and U25375 (N_25375,N_25034,N_25166);
or U25376 (N_25376,N_25042,N_24778);
and U25377 (N_25377,N_25008,N_25168);
or U25378 (N_25378,N_24858,N_24611);
nor U25379 (N_25379,N_24869,N_24743);
nand U25380 (N_25380,N_24916,N_24768);
or U25381 (N_25381,N_24663,N_24615);
xnor U25382 (N_25382,N_24702,N_25050);
nor U25383 (N_25383,N_24975,N_25124);
or U25384 (N_25384,N_24610,N_25088);
or U25385 (N_25385,N_25190,N_24929);
nand U25386 (N_25386,N_24902,N_24813);
or U25387 (N_25387,N_24843,N_25025);
nor U25388 (N_25388,N_24740,N_24836);
and U25389 (N_25389,N_24784,N_24842);
nand U25390 (N_25390,N_25051,N_24613);
nand U25391 (N_25391,N_25030,N_24965);
nand U25392 (N_25392,N_25077,N_24815);
or U25393 (N_25393,N_25084,N_24950);
nor U25394 (N_25394,N_25150,N_24817);
or U25395 (N_25395,N_24791,N_24826);
nor U25396 (N_25396,N_24662,N_24939);
nand U25397 (N_25397,N_24709,N_25063);
and U25398 (N_25398,N_24822,N_24787);
nor U25399 (N_25399,N_25129,N_24820);
nor U25400 (N_25400,N_24665,N_24695);
and U25401 (N_25401,N_25010,N_24999);
or U25402 (N_25402,N_24812,N_24966);
xnor U25403 (N_25403,N_24736,N_24790);
and U25404 (N_25404,N_24972,N_24794);
and U25405 (N_25405,N_24866,N_24907);
nor U25406 (N_25406,N_24899,N_25145);
and U25407 (N_25407,N_25003,N_25019);
and U25408 (N_25408,N_25139,N_24777);
nand U25409 (N_25409,N_24971,N_25083);
and U25410 (N_25410,N_24840,N_24637);
or U25411 (N_25411,N_25056,N_25002);
nor U25412 (N_25412,N_25133,N_25039);
nor U25413 (N_25413,N_24832,N_24893);
xor U25414 (N_25414,N_25163,N_24704);
or U25415 (N_25415,N_24911,N_24882);
or U25416 (N_25416,N_25053,N_24917);
or U25417 (N_25417,N_24685,N_24818);
or U25418 (N_25418,N_24735,N_25058);
or U25419 (N_25419,N_24874,N_24738);
nand U25420 (N_25420,N_25116,N_24931);
and U25421 (N_25421,N_24781,N_24690);
or U25422 (N_25422,N_24643,N_24864);
nor U25423 (N_25423,N_24823,N_24886);
or U25424 (N_25424,N_25182,N_24766);
nand U25425 (N_25425,N_24867,N_24616);
xnor U25426 (N_25426,N_24636,N_25185);
nand U25427 (N_25427,N_24926,N_25027);
and U25428 (N_25428,N_24912,N_24648);
nor U25429 (N_25429,N_24700,N_24795);
nor U25430 (N_25430,N_25101,N_24749);
nor U25431 (N_25431,N_25092,N_24660);
and U25432 (N_25432,N_25031,N_24684);
nand U25433 (N_25433,N_25067,N_25082);
or U25434 (N_25434,N_25149,N_24658);
nor U25435 (N_25435,N_25173,N_24970);
nor U25436 (N_25436,N_24927,N_25171);
nand U25437 (N_25437,N_24881,N_25199);
and U25438 (N_25438,N_25175,N_25074);
nor U25439 (N_25439,N_25125,N_24727);
and U25440 (N_25440,N_24992,N_24687);
and U25441 (N_25441,N_24698,N_24949);
or U25442 (N_25442,N_24739,N_24618);
nor U25443 (N_25443,N_24968,N_24638);
or U25444 (N_25444,N_24895,N_24839);
nor U25445 (N_25445,N_25001,N_25104);
nor U25446 (N_25446,N_25189,N_25026);
nand U25447 (N_25447,N_24641,N_24707);
xnor U25448 (N_25448,N_25085,N_25143);
and U25449 (N_25449,N_24705,N_25187);
nand U25450 (N_25450,N_25192,N_24951);
nor U25451 (N_25451,N_25048,N_24945);
or U25452 (N_25452,N_24798,N_25069);
or U25453 (N_25453,N_25137,N_24958);
and U25454 (N_25454,N_24824,N_24631);
and U25455 (N_25455,N_25047,N_24680);
nor U25456 (N_25456,N_24856,N_24834);
or U25457 (N_25457,N_24716,N_24621);
nand U25458 (N_25458,N_24940,N_24915);
nor U25459 (N_25459,N_24619,N_24952);
or U25460 (N_25460,N_25052,N_24688);
nand U25461 (N_25461,N_25079,N_25148);
or U25462 (N_25462,N_24938,N_24969);
or U25463 (N_25463,N_25180,N_25015);
nand U25464 (N_25464,N_24626,N_25059);
and U25465 (N_25465,N_24863,N_24897);
and U25466 (N_25466,N_24748,N_24819);
nor U25467 (N_25467,N_24774,N_25151);
and U25468 (N_25468,N_24632,N_24669);
or U25469 (N_25469,N_24761,N_24642);
nand U25470 (N_25470,N_24811,N_24908);
and U25471 (N_25471,N_24783,N_24786);
nand U25472 (N_25472,N_24733,N_24645);
and U25473 (N_25473,N_25172,N_24741);
xor U25474 (N_25474,N_24756,N_25127);
and U25475 (N_25475,N_25068,N_24981);
nor U25476 (N_25476,N_24801,N_25135);
nand U25477 (N_25477,N_25184,N_24746);
nor U25478 (N_25478,N_25183,N_25142);
and U25479 (N_25479,N_25122,N_24668);
or U25480 (N_25480,N_25020,N_24852);
and U25481 (N_25481,N_24729,N_24943);
nand U25482 (N_25482,N_25117,N_24674);
nor U25483 (N_25483,N_24764,N_24765);
nor U25484 (N_25484,N_24871,N_24935);
and U25485 (N_25485,N_25007,N_24682);
nor U25486 (N_25486,N_24865,N_24620);
and U25487 (N_25487,N_24804,N_24769);
and U25488 (N_25488,N_24904,N_25198);
nand U25489 (N_25489,N_24986,N_24942);
or U25490 (N_25490,N_24896,N_24767);
nand U25491 (N_25491,N_24657,N_24796);
xnor U25492 (N_25492,N_24706,N_24734);
and U25493 (N_25493,N_25138,N_24793);
and U25494 (N_25494,N_24928,N_25055);
xor U25495 (N_25495,N_25115,N_24757);
nor U25496 (N_25496,N_25193,N_25000);
nand U25497 (N_25497,N_25045,N_25017);
or U25498 (N_25498,N_25136,N_24898);
or U25499 (N_25499,N_24983,N_24624);
nand U25500 (N_25500,N_24877,N_24870);
nor U25501 (N_25501,N_24792,N_25182);
nor U25502 (N_25502,N_24860,N_24902);
or U25503 (N_25503,N_24765,N_25152);
and U25504 (N_25504,N_24702,N_25006);
nor U25505 (N_25505,N_25121,N_24800);
nand U25506 (N_25506,N_25064,N_25079);
and U25507 (N_25507,N_24706,N_25063);
nand U25508 (N_25508,N_24738,N_24996);
and U25509 (N_25509,N_25020,N_24716);
nor U25510 (N_25510,N_24892,N_24989);
or U25511 (N_25511,N_24829,N_24932);
and U25512 (N_25512,N_25158,N_24745);
and U25513 (N_25513,N_24900,N_24625);
and U25514 (N_25514,N_25135,N_25198);
nand U25515 (N_25515,N_24669,N_24780);
nand U25516 (N_25516,N_25161,N_24876);
or U25517 (N_25517,N_24639,N_25087);
and U25518 (N_25518,N_24767,N_25014);
nand U25519 (N_25519,N_24615,N_24916);
nand U25520 (N_25520,N_25105,N_24843);
nor U25521 (N_25521,N_24946,N_24772);
nor U25522 (N_25522,N_25127,N_25001);
and U25523 (N_25523,N_25102,N_24633);
nand U25524 (N_25524,N_25033,N_24894);
nand U25525 (N_25525,N_24967,N_24926);
nor U25526 (N_25526,N_24646,N_25070);
or U25527 (N_25527,N_24851,N_24809);
or U25528 (N_25528,N_24670,N_25063);
and U25529 (N_25529,N_24866,N_24707);
and U25530 (N_25530,N_24790,N_24873);
xor U25531 (N_25531,N_24874,N_25093);
nand U25532 (N_25532,N_25022,N_24603);
or U25533 (N_25533,N_24695,N_25062);
and U25534 (N_25534,N_24821,N_24688);
nor U25535 (N_25535,N_25198,N_24704);
and U25536 (N_25536,N_25132,N_25198);
nor U25537 (N_25537,N_25066,N_24912);
and U25538 (N_25538,N_25016,N_24698);
xor U25539 (N_25539,N_25103,N_24937);
and U25540 (N_25540,N_25107,N_24847);
and U25541 (N_25541,N_25134,N_24746);
and U25542 (N_25542,N_24811,N_24864);
nand U25543 (N_25543,N_24764,N_25056);
nor U25544 (N_25544,N_25062,N_24962);
and U25545 (N_25545,N_24919,N_25099);
and U25546 (N_25546,N_25131,N_24880);
nor U25547 (N_25547,N_25168,N_24806);
nand U25548 (N_25548,N_25025,N_24868);
or U25549 (N_25549,N_24917,N_24947);
nand U25550 (N_25550,N_25062,N_24639);
or U25551 (N_25551,N_25052,N_24682);
and U25552 (N_25552,N_24921,N_24697);
and U25553 (N_25553,N_24684,N_24874);
and U25554 (N_25554,N_24843,N_24666);
or U25555 (N_25555,N_25008,N_24803);
or U25556 (N_25556,N_24620,N_24951);
or U25557 (N_25557,N_25039,N_24699);
nor U25558 (N_25558,N_25037,N_25102);
nand U25559 (N_25559,N_25179,N_24767);
nand U25560 (N_25560,N_24953,N_25138);
or U25561 (N_25561,N_24822,N_24845);
or U25562 (N_25562,N_24959,N_24602);
or U25563 (N_25563,N_24930,N_25045);
nor U25564 (N_25564,N_24988,N_24645);
nor U25565 (N_25565,N_24753,N_24892);
or U25566 (N_25566,N_24690,N_25192);
xnor U25567 (N_25567,N_24648,N_24620);
nand U25568 (N_25568,N_25102,N_25191);
and U25569 (N_25569,N_24705,N_24879);
nor U25570 (N_25570,N_25181,N_25182);
nor U25571 (N_25571,N_24633,N_24924);
or U25572 (N_25572,N_24805,N_24632);
or U25573 (N_25573,N_24619,N_25063);
or U25574 (N_25574,N_25085,N_24695);
and U25575 (N_25575,N_24866,N_25154);
or U25576 (N_25576,N_24797,N_24877);
nor U25577 (N_25577,N_24731,N_24667);
or U25578 (N_25578,N_25169,N_24889);
or U25579 (N_25579,N_24613,N_25003);
or U25580 (N_25580,N_24836,N_25177);
and U25581 (N_25581,N_24894,N_25105);
or U25582 (N_25582,N_24619,N_25039);
nand U25583 (N_25583,N_24669,N_24670);
or U25584 (N_25584,N_24805,N_25157);
and U25585 (N_25585,N_24927,N_24983);
nor U25586 (N_25586,N_24812,N_25192);
and U25587 (N_25587,N_25090,N_24783);
and U25588 (N_25588,N_25097,N_24675);
and U25589 (N_25589,N_24981,N_24999);
nor U25590 (N_25590,N_24805,N_24731);
and U25591 (N_25591,N_24623,N_25066);
xnor U25592 (N_25592,N_24715,N_25119);
nand U25593 (N_25593,N_24716,N_24601);
nand U25594 (N_25594,N_25197,N_24986);
nand U25595 (N_25595,N_24829,N_24977);
nand U25596 (N_25596,N_24850,N_25171);
nand U25597 (N_25597,N_24965,N_24877);
and U25598 (N_25598,N_25003,N_24873);
nand U25599 (N_25599,N_24773,N_25058);
nand U25600 (N_25600,N_24654,N_24798);
nand U25601 (N_25601,N_24896,N_24846);
or U25602 (N_25602,N_24635,N_25075);
nor U25603 (N_25603,N_24854,N_24765);
nand U25604 (N_25604,N_24796,N_25057);
nor U25605 (N_25605,N_25183,N_24609);
or U25606 (N_25606,N_25087,N_24949);
or U25607 (N_25607,N_25016,N_24627);
and U25608 (N_25608,N_24976,N_25039);
and U25609 (N_25609,N_24826,N_24986);
or U25610 (N_25610,N_25052,N_24915);
and U25611 (N_25611,N_25161,N_24704);
nor U25612 (N_25612,N_24644,N_25125);
nand U25613 (N_25613,N_24978,N_24920);
and U25614 (N_25614,N_24955,N_25148);
and U25615 (N_25615,N_24731,N_25092);
nor U25616 (N_25616,N_24938,N_24913);
nand U25617 (N_25617,N_24900,N_24603);
and U25618 (N_25618,N_24867,N_24685);
and U25619 (N_25619,N_24660,N_24997);
xnor U25620 (N_25620,N_24778,N_24815);
or U25621 (N_25621,N_24851,N_25159);
nand U25622 (N_25622,N_25161,N_25055);
or U25623 (N_25623,N_25000,N_24602);
nand U25624 (N_25624,N_24611,N_25033);
and U25625 (N_25625,N_25057,N_24786);
and U25626 (N_25626,N_25158,N_24885);
nor U25627 (N_25627,N_24623,N_24693);
nand U25628 (N_25628,N_25155,N_24795);
nand U25629 (N_25629,N_24613,N_25083);
or U25630 (N_25630,N_24631,N_25166);
or U25631 (N_25631,N_24782,N_24959);
and U25632 (N_25632,N_25093,N_25118);
and U25633 (N_25633,N_25078,N_24729);
nand U25634 (N_25634,N_24774,N_24619);
or U25635 (N_25635,N_24841,N_24810);
nand U25636 (N_25636,N_24953,N_24726);
nor U25637 (N_25637,N_25031,N_24617);
and U25638 (N_25638,N_24830,N_24949);
or U25639 (N_25639,N_24744,N_24816);
and U25640 (N_25640,N_24714,N_24827);
nand U25641 (N_25641,N_24960,N_25121);
and U25642 (N_25642,N_25184,N_24718);
or U25643 (N_25643,N_25117,N_24951);
nand U25644 (N_25644,N_24764,N_24833);
or U25645 (N_25645,N_24982,N_25043);
and U25646 (N_25646,N_24870,N_24990);
nand U25647 (N_25647,N_24650,N_24613);
nand U25648 (N_25648,N_24789,N_24952);
or U25649 (N_25649,N_24811,N_25172);
or U25650 (N_25650,N_24626,N_25026);
or U25651 (N_25651,N_25091,N_24645);
or U25652 (N_25652,N_25172,N_24765);
nand U25653 (N_25653,N_25047,N_25033);
or U25654 (N_25654,N_25003,N_24892);
xor U25655 (N_25655,N_24734,N_25069);
and U25656 (N_25656,N_25026,N_24658);
or U25657 (N_25657,N_24601,N_24897);
or U25658 (N_25658,N_24949,N_25173);
nand U25659 (N_25659,N_24816,N_25076);
nand U25660 (N_25660,N_25055,N_24936);
nand U25661 (N_25661,N_24954,N_25049);
nand U25662 (N_25662,N_24700,N_25108);
xnor U25663 (N_25663,N_24822,N_24627);
xor U25664 (N_25664,N_24693,N_24794);
or U25665 (N_25665,N_25039,N_24697);
or U25666 (N_25666,N_25166,N_24726);
nand U25667 (N_25667,N_24697,N_24819);
nor U25668 (N_25668,N_24941,N_24658);
and U25669 (N_25669,N_24980,N_24815);
nand U25670 (N_25670,N_25026,N_25191);
or U25671 (N_25671,N_24905,N_25058);
nand U25672 (N_25672,N_25052,N_25156);
and U25673 (N_25673,N_25153,N_24656);
nand U25674 (N_25674,N_24948,N_24758);
and U25675 (N_25675,N_24759,N_24777);
or U25676 (N_25676,N_25008,N_24966);
nand U25677 (N_25677,N_24797,N_25095);
and U25678 (N_25678,N_24648,N_24903);
nor U25679 (N_25679,N_25042,N_24929);
and U25680 (N_25680,N_24838,N_24955);
nor U25681 (N_25681,N_24683,N_25089);
or U25682 (N_25682,N_24809,N_24865);
nand U25683 (N_25683,N_24857,N_24703);
nor U25684 (N_25684,N_25028,N_25024);
nand U25685 (N_25685,N_24689,N_24909);
nand U25686 (N_25686,N_24773,N_24913);
or U25687 (N_25687,N_24667,N_24727);
or U25688 (N_25688,N_24970,N_24668);
or U25689 (N_25689,N_24823,N_25098);
or U25690 (N_25690,N_25076,N_25130);
nor U25691 (N_25691,N_24896,N_24679);
nor U25692 (N_25692,N_25082,N_25057);
nor U25693 (N_25693,N_24780,N_24966);
and U25694 (N_25694,N_24797,N_25017);
and U25695 (N_25695,N_24674,N_24615);
or U25696 (N_25696,N_24712,N_24634);
nand U25697 (N_25697,N_25160,N_24836);
nand U25698 (N_25698,N_25008,N_24777);
nand U25699 (N_25699,N_25052,N_24722);
and U25700 (N_25700,N_25119,N_24650);
and U25701 (N_25701,N_24826,N_24885);
or U25702 (N_25702,N_25093,N_25196);
nand U25703 (N_25703,N_25095,N_24625);
or U25704 (N_25704,N_24895,N_24748);
and U25705 (N_25705,N_24777,N_25198);
nor U25706 (N_25706,N_24632,N_24741);
nor U25707 (N_25707,N_25106,N_24941);
nor U25708 (N_25708,N_24931,N_24798);
nor U25709 (N_25709,N_25136,N_24912);
and U25710 (N_25710,N_24967,N_24988);
nand U25711 (N_25711,N_25022,N_25117);
or U25712 (N_25712,N_24749,N_24936);
nand U25713 (N_25713,N_24621,N_25033);
and U25714 (N_25714,N_24756,N_24826);
nor U25715 (N_25715,N_24806,N_25173);
and U25716 (N_25716,N_25152,N_25008);
nor U25717 (N_25717,N_24702,N_24862);
and U25718 (N_25718,N_24791,N_25148);
and U25719 (N_25719,N_25110,N_24980);
and U25720 (N_25720,N_24630,N_24756);
or U25721 (N_25721,N_24848,N_24999);
or U25722 (N_25722,N_24891,N_24994);
or U25723 (N_25723,N_24913,N_24908);
nand U25724 (N_25724,N_25161,N_25094);
nor U25725 (N_25725,N_24604,N_25052);
and U25726 (N_25726,N_24777,N_24951);
nand U25727 (N_25727,N_25072,N_24961);
nand U25728 (N_25728,N_24877,N_24715);
nor U25729 (N_25729,N_25076,N_24694);
nand U25730 (N_25730,N_24923,N_25137);
nor U25731 (N_25731,N_24624,N_25026);
nand U25732 (N_25732,N_25039,N_24794);
and U25733 (N_25733,N_24799,N_25083);
nor U25734 (N_25734,N_24615,N_24692);
nand U25735 (N_25735,N_24656,N_24869);
and U25736 (N_25736,N_25117,N_24980);
and U25737 (N_25737,N_24678,N_25199);
and U25738 (N_25738,N_25102,N_24736);
nor U25739 (N_25739,N_24741,N_24700);
nand U25740 (N_25740,N_25095,N_24689);
nor U25741 (N_25741,N_24608,N_24887);
or U25742 (N_25742,N_24701,N_25160);
and U25743 (N_25743,N_24879,N_25066);
nor U25744 (N_25744,N_25117,N_24931);
and U25745 (N_25745,N_24789,N_25057);
and U25746 (N_25746,N_24823,N_25136);
nor U25747 (N_25747,N_24632,N_24681);
nand U25748 (N_25748,N_24897,N_25076);
or U25749 (N_25749,N_24681,N_24967);
or U25750 (N_25750,N_25104,N_24834);
or U25751 (N_25751,N_24989,N_24977);
nand U25752 (N_25752,N_25088,N_25022);
nand U25753 (N_25753,N_24667,N_25071);
nand U25754 (N_25754,N_24992,N_24771);
and U25755 (N_25755,N_24891,N_24763);
or U25756 (N_25756,N_24615,N_25121);
and U25757 (N_25757,N_24968,N_25049);
nor U25758 (N_25758,N_24682,N_25130);
nor U25759 (N_25759,N_24647,N_24865);
or U25760 (N_25760,N_24625,N_24642);
or U25761 (N_25761,N_24739,N_24848);
nor U25762 (N_25762,N_24802,N_24928);
or U25763 (N_25763,N_25082,N_24953);
or U25764 (N_25764,N_24874,N_25196);
nor U25765 (N_25765,N_24725,N_24601);
and U25766 (N_25766,N_24738,N_25082);
nor U25767 (N_25767,N_24689,N_25149);
and U25768 (N_25768,N_24988,N_24699);
or U25769 (N_25769,N_24620,N_24773);
nand U25770 (N_25770,N_24762,N_24943);
nand U25771 (N_25771,N_25161,N_24757);
nand U25772 (N_25772,N_25165,N_25197);
nor U25773 (N_25773,N_24602,N_24754);
nor U25774 (N_25774,N_24799,N_25112);
nand U25775 (N_25775,N_24741,N_24701);
xor U25776 (N_25776,N_25009,N_24689);
or U25777 (N_25777,N_25011,N_24611);
or U25778 (N_25778,N_25047,N_24809);
or U25779 (N_25779,N_24907,N_24931);
nor U25780 (N_25780,N_24919,N_24739);
or U25781 (N_25781,N_24927,N_25150);
or U25782 (N_25782,N_24996,N_25079);
or U25783 (N_25783,N_24774,N_24692);
or U25784 (N_25784,N_25035,N_25087);
nand U25785 (N_25785,N_24623,N_25081);
nand U25786 (N_25786,N_25107,N_24889);
and U25787 (N_25787,N_25189,N_24656);
nand U25788 (N_25788,N_24919,N_25175);
xnor U25789 (N_25789,N_24994,N_24787);
nand U25790 (N_25790,N_24611,N_24714);
nand U25791 (N_25791,N_25040,N_24923);
and U25792 (N_25792,N_25055,N_24733);
nor U25793 (N_25793,N_25079,N_24733);
and U25794 (N_25794,N_24635,N_25055);
or U25795 (N_25795,N_24824,N_24783);
or U25796 (N_25796,N_25066,N_24766);
xnor U25797 (N_25797,N_25150,N_25059);
nand U25798 (N_25798,N_25019,N_24679);
nand U25799 (N_25799,N_25048,N_24654);
or U25800 (N_25800,N_25497,N_25241);
or U25801 (N_25801,N_25778,N_25558);
nand U25802 (N_25802,N_25368,N_25288);
or U25803 (N_25803,N_25271,N_25696);
or U25804 (N_25804,N_25785,N_25638);
nand U25805 (N_25805,N_25701,N_25329);
and U25806 (N_25806,N_25485,N_25431);
nand U25807 (N_25807,N_25756,N_25570);
nor U25808 (N_25808,N_25261,N_25470);
nand U25809 (N_25809,N_25649,N_25416);
xor U25810 (N_25810,N_25510,N_25582);
and U25811 (N_25811,N_25281,N_25730);
nor U25812 (N_25812,N_25568,N_25243);
or U25813 (N_25813,N_25627,N_25611);
nor U25814 (N_25814,N_25695,N_25527);
or U25815 (N_25815,N_25762,N_25466);
and U25816 (N_25816,N_25467,N_25548);
nand U25817 (N_25817,N_25666,N_25704);
nor U25818 (N_25818,N_25700,N_25262);
and U25819 (N_25819,N_25289,N_25215);
nand U25820 (N_25820,N_25463,N_25655);
and U25821 (N_25821,N_25508,N_25745);
or U25822 (N_25822,N_25566,N_25279);
nor U25823 (N_25823,N_25617,N_25505);
xor U25824 (N_25824,N_25488,N_25425);
nand U25825 (N_25825,N_25353,N_25639);
nand U25826 (N_25826,N_25433,N_25320);
nor U25827 (N_25827,N_25385,N_25454);
and U25828 (N_25828,N_25294,N_25712);
or U25829 (N_25829,N_25343,N_25452);
nand U25830 (N_25830,N_25710,N_25274);
nand U25831 (N_25831,N_25217,N_25460);
nand U25832 (N_25832,N_25348,N_25699);
and U25833 (N_25833,N_25253,N_25543);
and U25834 (N_25834,N_25642,N_25647);
or U25835 (N_25835,N_25672,N_25677);
nand U25836 (N_25836,N_25683,N_25438);
nor U25837 (N_25837,N_25352,N_25635);
nor U25838 (N_25838,N_25507,N_25596);
nand U25839 (N_25839,N_25523,N_25761);
nor U25840 (N_25840,N_25685,N_25686);
nand U25841 (N_25841,N_25480,N_25398);
and U25842 (N_25842,N_25207,N_25300);
nor U25843 (N_25843,N_25220,N_25226);
and U25844 (N_25844,N_25235,N_25484);
nand U25845 (N_25845,N_25245,N_25412);
nor U25846 (N_25846,N_25204,N_25489);
and U25847 (N_25847,N_25334,N_25516);
or U25848 (N_25848,N_25268,N_25751);
nor U25849 (N_25849,N_25475,N_25400);
nor U25850 (N_25850,N_25342,N_25278);
nand U25851 (N_25851,N_25621,N_25780);
nand U25852 (N_25852,N_25284,N_25563);
or U25853 (N_25853,N_25509,N_25440);
nand U25854 (N_25854,N_25733,N_25585);
and U25855 (N_25855,N_25572,N_25703);
nand U25856 (N_25856,N_25275,N_25252);
or U25857 (N_25857,N_25238,N_25739);
and U25858 (N_25858,N_25656,N_25628);
and U25859 (N_25859,N_25513,N_25394);
nor U25860 (N_25860,N_25227,N_25589);
xnor U25861 (N_25861,N_25740,N_25673);
and U25862 (N_25862,N_25234,N_25715);
and U25863 (N_25863,N_25346,N_25461);
or U25864 (N_25864,N_25749,N_25758);
nor U25865 (N_25865,N_25541,N_25729);
nand U25866 (N_25866,N_25362,N_25794);
or U25867 (N_25867,N_25328,N_25256);
nor U25868 (N_25868,N_25378,N_25242);
nand U25869 (N_25869,N_25657,N_25308);
or U25870 (N_25870,N_25637,N_25392);
or U25871 (N_25871,N_25280,N_25233);
and U25872 (N_25872,N_25415,N_25623);
and U25873 (N_25873,N_25397,N_25512);
nand U25874 (N_25874,N_25551,N_25318);
and U25875 (N_25875,N_25532,N_25290);
nand U25876 (N_25876,N_25501,N_25727);
nor U25877 (N_25877,N_25239,N_25723);
and U25878 (N_25878,N_25326,N_25203);
nand U25879 (N_25879,N_25456,N_25269);
and U25880 (N_25880,N_25282,N_25283);
nor U25881 (N_25881,N_25725,N_25444);
or U25882 (N_25882,N_25626,N_25769);
and U25883 (N_25883,N_25313,N_25408);
and U25884 (N_25884,N_25607,N_25544);
and U25885 (N_25885,N_25735,N_25767);
or U25886 (N_25886,N_25731,N_25616);
and U25887 (N_25887,N_25371,N_25219);
nand U25888 (N_25888,N_25427,N_25646);
and U25889 (N_25889,N_25266,N_25539);
nor U25890 (N_25890,N_25522,N_25486);
or U25891 (N_25891,N_25298,N_25552);
or U25892 (N_25892,N_25345,N_25779);
nor U25893 (N_25893,N_25535,N_25609);
and U25894 (N_25894,N_25529,N_25306);
and U25895 (N_25895,N_25554,N_25765);
nand U25896 (N_25896,N_25369,N_25212);
nand U25897 (N_25897,N_25303,N_25316);
or U25898 (N_25898,N_25200,N_25618);
or U25899 (N_25899,N_25546,N_25366);
or U25900 (N_25900,N_25511,N_25653);
nor U25901 (N_25901,N_25766,N_25381);
nand U25902 (N_25902,N_25619,N_25521);
or U25903 (N_25903,N_25605,N_25755);
nor U25904 (N_25904,N_25406,N_25747);
nand U25905 (N_25905,N_25395,N_25292);
nor U25906 (N_25906,N_25559,N_25377);
and U25907 (N_25907,N_25561,N_25724);
and U25908 (N_25908,N_25692,N_25314);
and U25909 (N_25909,N_25597,N_25526);
or U25910 (N_25910,N_25569,N_25270);
nand U25911 (N_25911,N_25276,N_25500);
or U25912 (N_25912,N_25545,N_25549);
nor U25913 (N_25913,N_25386,N_25285);
or U25914 (N_25914,N_25413,N_25716);
nand U25915 (N_25915,N_25499,N_25437);
nor U25916 (N_25916,N_25713,N_25250);
or U25917 (N_25917,N_25520,N_25795);
or U25918 (N_25918,N_25721,N_25632);
nand U25919 (N_25919,N_25644,N_25665);
and U25920 (N_25920,N_25711,N_25240);
nor U25921 (N_25921,N_25741,N_25468);
nand U25922 (N_25922,N_25267,N_25670);
nor U25923 (N_25923,N_25319,N_25201);
nor U25924 (N_25924,N_25211,N_25449);
or U25925 (N_25925,N_25594,N_25702);
nor U25926 (N_25926,N_25722,N_25798);
and U25927 (N_25927,N_25379,N_25580);
and U25928 (N_25928,N_25364,N_25593);
nor U25929 (N_25929,N_25560,N_25445);
or U25930 (N_25930,N_25652,N_25325);
or U25931 (N_25931,N_25694,N_25365);
or U25932 (N_25932,N_25236,N_25663);
nand U25933 (N_25933,N_25595,N_25530);
nand U25934 (N_25934,N_25759,N_25356);
and U25935 (N_25935,N_25464,N_25213);
or U25936 (N_25936,N_25671,N_25459);
and U25937 (N_25937,N_25764,N_25732);
nand U25938 (N_25938,N_25455,N_25358);
and U25939 (N_25939,N_25299,N_25697);
or U25940 (N_25940,N_25693,N_25681);
and U25941 (N_25941,N_25717,N_25311);
or U25942 (N_25942,N_25351,N_25407);
or U25943 (N_25943,N_25575,N_25422);
nand U25944 (N_25944,N_25469,N_25772);
nor U25945 (N_25945,N_25206,N_25577);
nand U25946 (N_25946,N_25777,N_25481);
nor U25947 (N_25947,N_25660,N_25676);
and U25948 (N_25948,N_25610,N_25757);
or U25949 (N_25949,N_25327,N_25746);
nand U25950 (N_25950,N_25251,N_25781);
and U25951 (N_25951,N_25442,N_25567);
nor U25952 (N_25952,N_25606,N_25332);
nor U25953 (N_25953,N_25797,N_25230);
nor U25954 (N_25954,N_25424,N_25564);
or U25955 (N_25955,N_25426,N_25341);
or U25956 (N_25956,N_25380,N_25361);
or U25957 (N_25957,N_25375,N_25333);
nand U25958 (N_25958,N_25423,N_25331);
and U25959 (N_25959,N_25783,N_25528);
and U25960 (N_25960,N_25718,N_25542);
nand U25961 (N_25961,N_25232,N_25429);
nand U25962 (N_25962,N_25517,N_25583);
nor U25963 (N_25963,N_25453,N_25349);
and U25964 (N_25964,N_25465,N_25457);
nand U25965 (N_25965,N_25748,N_25750);
nand U25966 (N_25966,N_25436,N_25247);
nor U25967 (N_25967,N_25363,N_25602);
nor U25968 (N_25968,N_25643,N_25390);
nor U25969 (N_25969,N_25726,N_25374);
or U25970 (N_25970,N_25336,N_25293);
and U25971 (N_25971,N_25579,N_25448);
or U25972 (N_25972,N_25624,N_25474);
nor U25973 (N_25973,N_25738,N_25302);
and U25974 (N_25974,N_25492,N_25525);
nand U25975 (N_25975,N_25689,N_25337);
or U25976 (N_25976,N_25791,N_25471);
or U25977 (N_25977,N_25228,N_25387);
nand U25978 (N_25978,N_25418,N_25265);
and U25979 (N_25979,N_25592,N_25335);
nand U25980 (N_25980,N_25793,N_25237);
nor U25981 (N_25981,N_25221,N_25301);
and U25982 (N_25982,N_25691,N_25409);
or U25983 (N_25983,N_25600,N_25209);
nand U25984 (N_25984,N_25744,N_25405);
and U25985 (N_25985,N_25494,N_25340);
and U25986 (N_25986,N_25305,N_25753);
nand U25987 (N_25987,N_25590,N_25477);
or U25988 (N_25988,N_25705,N_25376);
or U25989 (N_25989,N_25678,N_25790);
or U25990 (N_25990,N_25439,N_25555);
nor U25991 (N_25991,N_25519,N_25706);
xor U25992 (N_25992,N_25502,N_25799);
nor U25993 (N_25993,N_25355,N_25402);
and U25994 (N_25994,N_25734,N_25773);
or U25995 (N_25995,N_25556,N_25255);
nor U25996 (N_25996,N_25410,N_25789);
or U25997 (N_25997,N_25222,N_25434);
nand U25998 (N_25998,N_25514,N_25272);
and U25999 (N_25999,N_25728,N_25675);
and U26000 (N_26000,N_25372,N_25630);
nand U26001 (N_26001,N_25441,N_25614);
nand U26002 (N_26002,N_25792,N_25312);
and U26003 (N_26003,N_25506,N_25458);
and U26004 (N_26004,N_25383,N_25622);
nor U26005 (N_26005,N_25651,N_25359);
nor U26006 (N_26006,N_25538,N_25629);
nor U26007 (N_26007,N_25553,N_25659);
nor U26008 (N_26008,N_25478,N_25679);
or U26009 (N_26009,N_25536,N_25518);
or U26010 (N_26010,N_25490,N_25664);
and U26011 (N_26011,N_25771,N_25354);
and U26012 (N_26012,N_25287,N_25350);
xor U26013 (N_26013,N_25736,N_25291);
and U26014 (N_26014,N_25472,N_25752);
and U26015 (N_26015,N_25491,N_25446);
nand U26016 (N_26016,N_25216,N_25373);
and U26017 (N_26017,N_25246,N_25550);
nand U26018 (N_26018,N_25317,N_25263);
and U26019 (N_26019,N_25384,N_25615);
and U26020 (N_26020,N_25401,N_25304);
and U26021 (N_26021,N_25339,N_25260);
and U26022 (N_26022,N_25309,N_25450);
and U26023 (N_26023,N_25286,N_25669);
nand U26024 (N_26024,N_25571,N_25770);
or U26025 (N_26025,N_25613,N_25205);
or U26026 (N_26026,N_25760,N_25248);
nand U26027 (N_26027,N_25487,N_25229);
nor U26028 (N_26028,N_25584,N_25668);
nand U26029 (N_26029,N_25598,N_25708);
nand U26030 (N_26030,N_25462,N_25581);
nand U26031 (N_26031,N_25537,N_25447);
nand U26032 (N_26032,N_25743,N_25432);
nor U26033 (N_26033,N_25620,N_25684);
and U26034 (N_26034,N_25295,N_25565);
and U26035 (N_26035,N_25451,N_25310);
nand U26036 (N_26036,N_25688,N_25367);
nor U26037 (N_26037,N_25557,N_25608);
nor U26038 (N_26038,N_25625,N_25641);
and U26039 (N_26039,N_25709,N_25719);
nand U26040 (N_26040,N_25257,N_25443);
nor U26041 (N_26041,N_25742,N_25210);
or U26042 (N_26042,N_25667,N_25588);
or U26043 (N_26043,N_25404,N_25674);
or U26044 (N_26044,N_25504,N_25591);
and U26045 (N_26045,N_25254,N_25391);
nand U26046 (N_26046,N_25224,N_25495);
nand U26047 (N_26047,N_25421,N_25763);
nand U26048 (N_26048,N_25786,N_25698);
nand U26049 (N_26049,N_25498,N_25493);
or U26050 (N_26050,N_25259,N_25403);
or U26051 (N_26051,N_25399,N_25603);
nand U26052 (N_26052,N_25357,N_25788);
or U26053 (N_26053,N_25574,N_25690);
and U26054 (N_26054,N_25482,N_25389);
and U26055 (N_26055,N_25223,N_25636);
nand U26056 (N_26056,N_25633,N_25393);
or U26057 (N_26057,N_25277,N_25202);
or U26058 (N_26058,N_25540,N_25428);
nor U26059 (N_26059,N_25524,N_25218);
nor U26060 (N_26060,N_25662,N_25338);
or U26061 (N_26061,N_25754,N_25476);
and U26062 (N_26062,N_25782,N_25658);
nor U26063 (N_26063,N_25515,N_25648);
and U26064 (N_26064,N_25347,N_25714);
or U26065 (N_26065,N_25388,N_25214);
or U26066 (N_26066,N_25587,N_25599);
nor U26067 (N_26067,N_25419,N_25562);
and U26068 (N_26068,N_25775,N_25307);
nor U26069 (N_26069,N_25707,N_25586);
or U26070 (N_26070,N_25680,N_25654);
and U26071 (N_26071,N_25370,N_25737);
or U26072 (N_26072,N_25787,N_25547);
nor U26073 (N_26073,N_25612,N_25435);
nor U26074 (N_26074,N_25682,N_25322);
and U26075 (N_26075,N_25344,N_25768);
nand U26076 (N_26076,N_25776,N_25645);
and U26077 (N_26077,N_25796,N_25496);
and U26078 (N_26078,N_25360,N_25650);
nor U26079 (N_26079,N_25258,N_25297);
xor U26080 (N_26080,N_25640,N_25324);
nand U26081 (N_26081,N_25420,N_25417);
or U26082 (N_26082,N_25273,N_25483);
and U26083 (N_26083,N_25784,N_25225);
nor U26084 (N_26084,N_25323,N_25249);
nor U26085 (N_26085,N_25479,N_25315);
xnor U26086 (N_26086,N_25411,N_25604);
nand U26087 (N_26087,N_25396,N_25576);
nor U26088 (N_26088,N_25330,N_25382);
nand U26089 (N_26089,N_25414,N_25503);
and U26090 (N_26090,N_25430,N_25631);
and U26091 (N_26091,N_25774,N_25264);
and U26092 (N_26092,N_25601,N_25321);
and U26093 (N_26093,N_25573,N_25208);
xor U26094 (N_26094,N_25533,N_25296);
nor U26095 (N_26095,N_25473,N_25531);
or U26096 (N_26096,N_25231,N_25687);
nor U26097 (N_26097,N_25578,N_25534);
nor U26098 (N_26098,N_25244,N_25661);
or U26099 (N_26099,N_25720,N_25634);
nand U26100 (N_26100,N_25418,N_25477);
nor U26101 (N_26101,N_25522,N_25510);
and U26102 (N_26102,N_25452,N_25465);
nor U26103 (N_26103,N_25524,N_25231);
or U26104 (N_26104,N_25337,N_25460);
nor U26105 (N_26105,N_25252,N_25479);
or U26106 (N_26106,N_25220,N_25682);
or U26107 (N_26107,N_25618,N_25748);
nor U26108 (N_26108,N_25544,N_25214);
or U26109 (N_26109,N_25311,N_25672);
or U26110 (N_26110,N_25464,N_25301);
nor U26111 (N_26111,N_25711,N_25276);
nand U26112 (N_26112,N_25416,N_25564);
nor U26113 (N_26113,N_25311,N_25567);
and U26114 (N_26114,N_25364,N_25711);
nor U26115 (N_26115,N_25713,N_25636);
nor U26116 (N_26116,N_25421,N_25793);
nand U26117 (N_26117,N_25599,N_25362);
or U26118 (N_26118,N_25569,N_25378);
nor U26119 (N_26119,N_25623,N_25409);
and U26120 (N_26120,N_25305,N_25525);
nor U26121 (N_26121,N_25526,N_25640);
nor U26122 (N_26122,N_25579,N_25223);
or U26123 (N_26123,N_25540,N_25201);
and U26124 (N_26124,N_25688,N_25238);
nor U26125 (N_26125,N_25347,N_25632);
nand U26126 (N_26126,N_25545,N_25538);
nand U26127 (N_26127,N_25661,N_25472);
nor U26128 (N_26128,N_25593,N_25309);
nand U26129 (N_26129,N_25641,N_25391);
nor U26130 (N_26130,N_25617,N_25705);
nand U26131 (N_26131,N_25707,N_25752);
nor U26132 (N_26132,N_25377,N_25437);
and U26133 (N_26133,N_25448,N_25518);
or U26134 (N_26134,N_25257,N_25615);
nor U26135 (N_26135,N_25400,N_25731);
nor U26136 (N_26136,N_25326,N_25579);
or U26137 (N_26137,N_25587,N_25388);
or U26138 (N_26138,N_25322,N_25357);
nand U26139 (N_26139,N_25699,N_25204);
nor U26140 (N_26140,N_25576,N_25601);
nand U26141 (N_26141,N_25520,N_25469);
nand U26142 (N_26142,N_25587,N_25504);
nor U26143 (N_26143,N_25208,N_25545);
or U26144 (N_26144,N_25338,N_25737);
nor U26145 (N_26145,N_25581,N_25740);
or U26146 (N_26146,N_25633,N_25608);
nor U26147 (N_26147,N_25399,N_25223);
or U26148 (N_26148,N_25655,N_25568);
or U26149 (N_26149,N_25341,N_25693);
or U26150 (N_26150,N_25223,N_25493);
and U26151 (N_26151,N_25437,N_25247);
and U26152 (N_26152,N_25586,N_25525);
and U26153 (N_26153,N_25307,N_25753);
and U26154 (N_26154,N_25380,N_25740);
and U26155 (N_26155,N_25363,N_25423);
nor U26156 (N_26156,N_25312,N_25354);
nand U26157 (N_26157,N_25322,N_25475);
nor U26158 (N_26158,N_25652,N_25680);
nand U26159 (N_26159,N_25534,N_25217);
or U26160 (N_26160,N_25401,N_25345);
and U26161 (N_26161,N_25287,N_25263);
and U26162 (N_26162,N_25550,N_25358);
or U26163 (N_26163,N_25517,N_25418);
nor U26164 (N_26164,N_25602,N_25613);
or U26165 (N_26165,N_25545,N_25216);
nand U26166 (N_26166,N_25490,N_25326);
nand U26167 (N_26167,N_25701,N_25276);
nand U26168 (N_26168,N_25651,N_25618);
or U26169 (N_26169,N_25360,N_25228);
nand U26170 (N_26170,N_25706,N_25668);
or U26171 (N_26171,N_25216,N_25411);
nor U26172 (N_26172,N_25496,N_25537);
nor U26173 (N_26173,N_25264,N_25302);
or U26174 (N_26174,N_25437,N_25588);
nand U26175 (N_26175,N_25529,N_25328);
nand U26176 (N_26176,N_25213,N_25584);
or U26177 (N_26177,N_25376,N_25266);
nand U26178 (N_26178,N_25328,N_25400);
or U26179 (N_26179,N_25571,N_25449);
nand U26180 (N_26180,N_25429,N_25537);
and U26181 (N_26181,N_25455,N_25438);
or U26182 (N_26182,N_25436,N_25230);
and U26183 (N_26183,N_25313,N_25798);
and U26184 (N_26184,N_25312,N_25427);
or U26185 (N_26185,N_25511,N_25732);
nor U26186 (N_26186,N_25455,N_25574);
and U26187 (N_26187,N_25770,N_25468);
xnor U26188 (N_26188,N_25794,N_25286);
nor U26189 (N_26189,N_25515,N_25693);
and U26190 (N_26190,N_25242,N_25302);
nor U26191 (N_26191,N_25387,N_25593);
xnor U26192 (N_26192,N_25383,N_25456);
and U26193 (N_26193,N_25313,N_25691);
nand U26194 (N_26194,N_25658,N_25391);
nand U26195 (N_26195,N_25651,N_25354);
xor U26196 (N_26196,N_25474,N_25281);
nor U26197 (N_26197,N_25565,N_25625);
or U26198 (N_26198,N_25309,N_25750);
nor U26199 (N_26199,N_25557,N_25786);
nand U26200 (N_26200,N_25437,N_25677);
nor U26201 (N_26201,N_25556,N_25777);
nand U26202 (N_26202,N_25226,N_25793);
or U26203 (N_26203,N_25568,N_25206);
nand U26204 (N_26204,N_25675,N_25634);
or U26205 (N_26205,N_25537,N_25252);
nand U26206 (N_26206,N_25671,N_25332);
and U26207 (N_26207,N_25681,N_25748);
and U26208 (N_26208,N_25435,N_25319);
nand U26209 (N_26209,N_25300,N_25592);
nor U26210 (N_26210,N_25250,N_25263);
nand U26211 (N_26211,N_25597,N_25209);
or U26212 (N_26212,N_25471,N_25444);
and U26213 (N_26213,N_25227,N_25668);
nor U26214 (N_26214,N_25348,N_25284);
nor U26215 (N_26215,N_25446,N_25560);
xor U26216 (N_26216,N_25437,N_25495);
nor U26217 (N_26217,N_25517,N_25693);
nor U26218 (N_26218,N_25652,N_25385);
and U26219 (N_26219,N_25590,N_25508);
nand U26220 (N_26220,N_25318,N_25205);
and U26221 (N_26221,N_25388,N_25445);
nand U26222 (N_26222,N_25498,N_25745);
and U26223 (N_26223,N_25414,N_25293);
nor U26224 (N_26224,N_25460,N_25750);
nand U26225 (N_26225,N_25790,N_25436);
or U26226 (N_26226,N_25679,N_25533);
nor U26227 (N_26227,N_25430,N_25749);
nand U26228 (N_26228,N_25499,N_25519);
nor U26229 (N_26229,N_25732,N_25792);
nor U26230 (N_26230,N_25588,N_25432);
nor U26231 (N_26231,N_25526,N_25577);
or U26232 (N_26232,N_25785,N_25793);
and U26233 (N_26233,N_25546,N_25617);
or U26234 (N_26234,N_25605,N_25604);
nand U26235 (N_26235,N_25618,N_25764);
and U26236 (N_26236,N_25525,N_25289);
nor U26237 (N_26237,N_25264,N_25720);
and U26238 (N_26238,N_25650,N_25263);
nor U26239 (N_26239,N_25415,N_25725);
nand U26240 (N_26240,N_25449,N_25360);
nor U26241 (N_26241,N_25234,N_25328);
xnor U26242 (N_26242,N_25416,N_25720);
or U26243 (N_26243,N_25389,N_25630);
or U26244 (N_26244,N_25754,N_25500);
nand U26245 (N_26245,N_25465,N_25556);
and U26246 (N_26246,N_25259,N_25374);
and U26247 (N_26247,N_25640,N_25723);
nor U26248 (N_26248,N_25574,N_25425);
and U26249 (N_26249,N_25261,N_25795);
nand U26250 (N_26250,N_25278,N_25501);
and U26251 (N_26251,N_25438,N_25721);
or U26252 (N_26252,N_25544,N_25443);
or U26253 (N_26253,N_25262,N_25663);
nand U26254 (N_26254,N_25679,N_25617);
xor U26255 (N_26255,N_25200,N_25790);
nor U26256 (N_26256,N_25315,N_25634);
or U26257 (N_26257,N_25403,N_25476);
nor U26258 (N_26258,N_25503,N_25776);
or U26259 (N_26259,N_25250,N_25202);
nor U26260 (N_26260,N_25500,N_25548);
xnor U26261 (N_26261,N_25793,N_25495);
or U26262 (N_26262,N_25537,N_25674);
xnor U26263 (N_26263,N_25403,N_25634);
nand U26264 (N_26264,N_25589,N_25278);
nand U26265 (N_26265,N_25731,N_25512);
or U26266 (N_26266,N_25612,N_25540);
nor U26267 (N_26267,N_25522,N_25362);
and U26268 (N_26268,N_25659,N_25740);
nor U26269 (N_26269,N_25721,N_25648);
or U26270 (N_26270,N_25255,N_25561);
and U26271 (N_26271,N_25439,N_25546);
and U26272 (N_26272,N_25257,N_25307);
nor U26273 (N_26273,N_25389,N_25418);
or U26274 (N_26274,N_25653,N_25437);
nor U26275 (N_26275,N_25349,N_25368);
nand U26276 (N_26276,N_25415,N_25481);
and U26277 (N_26277,N_25794,N_25738);
and U26278 (N_26278,N_25660,N_25344);
nor U26279 (N_26279,N_25781,N_25526);
or U26280 (N_26280,N_25223,N_25560);
nor U26281 (N_26281,N_25621,N_25453);
and U26282 (N_26282,N_25628,N_25322);
nor U26283 (N_26283,N_25267,N_25356);
nor U26284 (N_26284,N_25539,N_25653);
nand U26285 (N_26285,N_25278,N_25538);
nand U26286 (N_26286,N_25338,N_25469);
nor U26287 (N_26287,N_25652,N_25646);
or U26288 (N_26288,N_25612,N_25233);
and U26289 (N_26289,N_25633,N_25418);
nor U26290 (N_26290,N_25491,N_25277);
nor U26291 (N_26291,N_25252,N_25687);
nand U26292 (N_26292,N_25393,N_25478);
or U26293 (N_26293,N_25496,N_25467);
or U26294 (N_26294,N_25421,N_25713);
nand U26295 (N_26295,N_25506,N_25234);
or U26296 (N_26296,N_25206,N_25298);
or U26297 (N_26297,N_25654,N_25266);
or U26298 (N_26298,N_25340,N_25625);
nand U26299 (N_26299,N_25511,N_25523);
or U26300 (N_26300,N_25613,N_25665);
and U26301 (N_26301,N_25564,N_25227);
and U26302 (N_26302,N_25754,N_25752);
nor U26303 (N_26303,N_25626,N_25257);
and U26304 (N_26304,N_25794,N_25343);
or U26305 (N_26305,N_25513,N_25346);
or U26306 (N_26306,N_25466,N_25765);
or U26307 (N_26307,N_25287,N_25316);
or U26308 (N_26308,N_25461,N_25632);
nand U26309 (N_26309,N_25280,N_25229);
or U26310 (N_26310,N_25211,N_25371);
and U26311 (N_26311,N_25524,N_25352);
nand U26312 (N_26312,N_25499,N_25526);
and U26313 (N_26313,N_25708,N_25278);
or U26314 (N_26314,N_25320,N_25744);
nor U26315 (N_26315,N_25483,N_25712);
or U26316 (N_26316,N_25770,N_25581);
nand U26317 (N_26317,N_25453,N_25334);
nor U26318 (N_26318,N_25358,N_25747);
and U26319 (N_26319,N_25288,N_25674);
nor U26320 (N_26320,N_25657,N_25355);
or U26321 (N_26321,N_25258,N_25647);
nor U26322 (N_26322,N_25734,N_25697);
nor U26323 (N_26323,N_25686,N_25462);
nand U26324 (N_26324,N_25286,N_25574);
nor U26325 (N_26325,N_25567,N_25710);
nand U26326 (N_26326,N_25709,N_25715);
or U26327 (N_26327,N_25405,N_25545);
or U26328 (N_26328,N_25270,N_25644);
or U26329 (N_26329,N_25444,N_25734);
and U26330 (N_26330,N_25612,N_25751);
and U26331 (N_26331,N_25244,N_25246);
nand U26332 (N_26332,N_25737,N_25378);
and U26333 (N_26333,N_25687,N_25287);
nand U26334 (N_26334,N_25207,N_25291);
nand U26335 (N_26335,N_25299,N_25280);
or U26336 (N_26336,N_25732,N_25490);
and U26337 (N_26337,N_25729,N_25681);
and U26338 (N_26338,N_25759,N_25679);
and U26339 (N_26339,N_25769,N_25503);
or U26340 (N_26340,N_25525,N_25601);
nor U26341 (N_26341,N_25732,N_25643);
nor U26342 (N_26342,N_25735,N_25778);
nand U26343 (N_26343,N_25612,N_25723);
and U26344 (N_26344,N_25577,N_25459);
or U26345 (N_26345,N_25633,N_25250);
or U26346 (N_26346,N_25565,N_25328);
nand U26347 (N_26347,N_25436,N_25474);
or U26348 (N_26348,N_25783,N_25712);
nand U26349 (N_26349,N_25242,N_25584);
and U26350 (N_26350,N_25221,N_25324);
xor U26351 (N_26351,N_25527,N_25520);
nor U26352 (N_26352,N_25683,N_25666);
or U26353 (N_26353,N_25628,N_25285);
nor U26354 (N_26354,N_25526,N_25354);
or U26355 (N_26355,N_25226,N_25740);
xor U26356 (N_26356,N_25663,N_25605);
nor U26357 (N_26357,N_25400,N_25264);
and U26358 (N_26358,N_25273,N_25599);
or U26359 (N_26359,N_25684,N_25599);
nand U26360 (N_26360,N_25329,N_25776);
nor U26361 (N_26361,N_25642,N_25316);
nand U26362 (N_26362,N_25217,N_25643);
nor U26363 (N_26363,N_25205,N_25274);
and U26364 (N_26364,N_25650,N_25497);
and U26365 (N_26365,N_25326,N_25404);
or U26366 (N_26366,N_25238,N_25475);
and U26367 (N_26367,N_25764,N_25412);
nand U26368 (N_26368,N_25234,N_25657);
nor U26369 (N_26369,N_25573,N_25329);
nand U26370 (N_26370,N_25464,N_25669);
nor U26371 (N_26371,N_25534,N_25202);
nand U26372 (N_26372,N_25448,N_25409);
and U26373 (N_26373,N_25301,N_25382);
nand U26374 (N_26374,N_25612,N_25787);
nand U26375 (N_26375,N_25450,N_25233);
or U26376 (N_26376,N_25737,N_25681);
or U26377 (N_26377,N_25237,N_25339);
nor U26378 (N_26378,N_25784,N_25233);
or U26379 (N_26379,N_25719,N_25364);
nand U26380 (N_26380,N_25729,N_25394);
and U26381 (N_26381,N_25653,N_25394);
and U26382 (N_26382,N_25589,N_25345);
nand U26383 (N_26383,N_25718,N_25371);
and U26384 (N_26384,N_25570,N_25695);
and U26385 (N_26385,N_25494,N_25279);
and U26386 (N_26386,N_25312,N_25673);
and U26387 (N_26387,N_25663,N_25425);
and U26388 (N_26388,N_25722,N_25656);
nor U26389 (N_26389,N_25621,N_25637);
and U26390 (N_26390,N_25290,N_25289);
or U26391 (N_26391,N_25393,N_25443);
nor U26392 (N_26392,N_25334,N_25298);
and U26393 (N_26393,N_25260,N_25216);
nor U26394 (N_26394,N_25200,N_25211);
and U26395 (N_26395,N_25424,N_25614);
and U26396 (N_26396,N_25711,N_25438);
nor U26397 (N_26397,N_25290,N_25602);
or U26398 (N_26398,N_25532,N_25235);
nand U26399 (N_26399,N_25786,N_25791);
nor U26400 (N_26400,N_26260,N_26238);
nand U26401 (N_26401,N_26229,N_26006);
nand U26402 (N_26402,N_26291,N_26374);
or U26403 (N_26403,N_25861,N_25885);
nor U26404 (N_26404,N_26340,N_26095);
and U26405 (N_26405,N_25862,N_26258);
or U26406 (N_26406,N_26193,N_26005);
xnor U26407 (N_26407,N_25998,N_26345);
xnor U26408 (N_26408,N_26314,N_25850);
or U26409 (N_26409,N_26011,N_25841);
or U26410 (N_26410,N_26267,N_26104);
nor U26411 (N_26411,N_26353,N_25995);
and U26412 (N_26412,N_26307,N_26155);
nand U26413 (N_26413,N_25991,N_25871);
or U26414 (N_26414,N_25986,N_26173);
and U26415 (N_26415,N_25879,N_25881);
xnor U26416 (N_26416,N_25920,N_25821);
nor U26417 (N_26417,N_26209,N_26244);
and U26418 (N_26418,N_26280,N_26089);
nor U26419 (N_26419,N_26042,N_26248);
or U26420 (N_26420,N_25978,N_25804);
nor U26421 (N_26421,N_26312,N_26182);
nand U26422 (N_26422,N_26008,N_26096);
nand U26423 (N_26423,N_26204,N_26187);
nand U26424 (N_26424,N_26144,N_26360);
nor U26425 (N_26425,N_26088,N_26196);
nor U26426 (N_26426,N_26143,N_26121);
nand U26427 (N_26427,N_26053,N_26166);
and U26428 (N_26428,N_25926,N_26357);
and U26429 (N_26429,N_26253,N_26092);
nand U26430 (N_26430,N_25963,N_26230);
and U26431 (N_26431,N_25810,N_26098);
nand U26432 (N_26432,N_26276,N_25817);
and U26433 (N_26433,N_26156,N_26003);
and U26434 (N_26434,N_25925,N_26079);
nand U26435 (N_26435,N_26086,N_25863);
nor U26436 (N_26436,N_26164,N_25967);
and U26437 (N_26437,N_25945,N_26215);
nand U26438 (N_26438,N_26128,N_26054);
and U26439 (N_26439,N_26059,N_26334);
and U26440 (N_26440,N_26037,N_25917);
nor U26441 (N_26441,N_26183,N_25895);
nor U26442 (N_26442,N_25903,N_26284);
and U26443 (N_26443,N_25875,N_25912);
and U26444 (N_26444,N_26289,N_25883);
and U26445 (N_26445,N_25975,N_26061);
nand U26446 (N_26446,N_26337,N_26002);
nor U26447 (N_26447,N_26336,N_25834);
nor U26448 (N_26448,N_26249,N_26397);
or U26449 (N_26449,N_26222,N_26024);
and U26450 (N_26450,N_26090,N_26243);
nand U26451 (N_26451,N_25909,N_25935);
nand U26452 (N_26452,N_26073,N_25872);
and U26453 (N_26453,N_26110,N_26264);
and U26454 (N_26454,N_25901,N_26081);
nand U26455 (N_26455,N_26069,N_25851);
or U26456 (N_26456,N_26254,N_25959);
and U26457 (N_26457,N_26318,N_26093);
nand U26458 (N_26458,N_25825,N_25980);
and U26459 (N_26459,N_26389,N_25853);
nand U26460 (N_26460,N_26169,N_25882);
or U26461 (N_26461,N_26192,N_26056);
nor U26462 (N_26462,N_25904,N_26298);
or U26463 (N_26463,N_26027,N_26206);
nand U26464 (N_26464,N_25969,N_25809);
nand U26465 (N_26465,N_26064,N_25907);
nor U26466 (N_26466,N_25892,N_26299);
and U26467 (N_26467,N_25974,N_25988);
nand U26468 (N_26468,N_26372,N_26177);
or U26469 (N_26469,N_26235,N_26295);
nor U26470 (N_26470,N_25927,N_26242);
xor U26471 (N_26471,N_25830,N_26210);
or U26472 (N_26472,N_26306,N_26287);
and U26473 (N_26473,N_26102,N_26218);
or U26474 (N_26474,N_26286,N_26065);
nor U26475 (N_26475,N_25921,N_25962);
or U26476 (N_26476,N_26224,N_25824);
xor U26477 (N_26477,N_26203,N_26097);
nand U26478 (N_26478,N_26040,N_25874);
and U26479 (N_26479,N_25865,N_26269);
and U26480 (N_26480,N_26375,N_26111);
or U26481 (N_26481,N_26029,N_25803);
xnor U26482 (N_26482,N_26139,N_25968);
and U26483 (N_26483,N_26329,N_26311);
or U26484 (N_26484,N_26341,N_26259);
nor U26485 (N_26485,N_25994,N_26300);
nor U26486 (N_26486,N_25965,N_25807);
nor U26487 (N_26487,N_25955,N_26068);
or U26488 (N_26488,N_26162,N_26366);
or U26489 (N_26489,N_25835,N_26256);
or U26490 (N_26490,N_26383,N_26189);
nor U26491 (N_26491,N_26220,N_26232);
or U26492 (N_26492,N_26050,N_25939);
and U26493 (N_26493,N_26344,N_26127);
nor U26494 (N_26494,N_26246,N_26045);
and U26495 (N_26495,N_26292,N_25930);
nor U26496 (N_26496,N_26191,N_26154);
nand U26497 (N_26497,N_25948,N_26018);
nand U26498 (N_26498,N_25946,N_26039);
nand U26499 (N_26499,N_26009,N_26172);
nor U26500 (N_26500,N_26138,N_26352);
or U26501 (N_26501,N_26240,N_26161);
and U26502 (N_26502,N_26396,N_26371);
and U26503 (N_26503,N_25977,N_26219);
nand U26504 (N_26504,N_25877,N_26369);
nor U26505 (N_26505,N_26361,N_25828);
nor U26506 (N_26506,N_25818,N_25833);
or U26507 (N_26507,N_26294,N_25934);
nor U26508 (N_26508,N_25944,N_26355);
nand U26509 (N_26509,N_25808,N_25814);
and U26510 (N_26510,N_26058,N_26152);
or U26511 (N_26511,N_25888,N_25849);
xnor U26512 (N_26512,N_26150,N_26350);
nand U26513 (N_26513,N_26216,N_25823);
or U26514 (N_26514,N_25820,N_26207);
nand U26515 (N_26515,N_26010,N_25936);
nor U26516 (N_26516,N_25836,N_25845);
and U26517 (N_26517,N_26308,N_26084);
nor U26518 (N_26518,N_26339,N_26321);
nand U26519 (N_26519,N_26384,N_26025);
nand U26520 (N_26520,N_25916,N_26087);
and U26521 (N_26521,N_26133,N_25982);
or U26522 (N_26522,N_26033,N_26060);
or U26523 (N_26523,N_25816,N_26171);
nor U26524 (N_26524,N_26113,N_26099);
nor U26525 (N_26525,N_25812,N_26380);
and U26526 (N_26526,N_26153,N_26176);
nand U26527 (N_26527,N_25911,N_26062);
nor U26528 (N_26528,N_26019,N_26313);
nand U26529 (N_26529,N_26022,N_25842);
and U26530 (N_26530,N_26226,N_26293);
or U26531 (N_26531,N_26358,N_25932);
nand U26532 (N_26532,N_25899,N_26221);
nand U26533 (N_26533,N_26075,N_26028);
nand U26534 (N_26534,N_26142,N_26195);
nor U26535 (N_26535,N_25940,N_26208);
nand U26536 (N_26536,N_25894,N_26163);
nor U26537 (N_26537,N_25897,N_26119);
nand U26538 (N_26538,N_26145,N_25949);
or U26539 (N_26539,N_26325,N_26198);
or U26540 (N_26540,N_25848,N_26381);
and U26541 (N_26541,N_26034,N_26117);
nand U26542 (N_26542,N_25800,N_26326);
nand U26543 (N_26543,N_26237,N_26082);
and U26544 (N_26544,N_26103,N_26363);
nor U26545 (N_26545,N_26083,N_26250);
nand U26546 (N_26546,N_26275,N_26115);
and U26547 (N_26547,N_26324,N_26342);
or U26548 (N_26548,N_26211,N_25910);
or U26549 (N_26549,N_25964,N_26303);
and U26550 (N_26550,N_26094,N_25838);
and U26551 (N_26551,N_25933,N_26051);
nand U26552 (N_26552,N_26388,N_25870);
nor U26553 (N_26553,N_26035,N_26365);
or U26554 (N_26554,N_26078,N_25905);
or U26555 (N_26555,N_25919,N_26335);
nand U26556 (N_26556,N_26330,N_25958);
xnor U26557 (N_26557,N_26399,N_25873);
or U26558 (N_26558,N_25947,N_26251);
or U26559 (N_26559,N_26016,N_26131);
nand U26560 (N_26560,N_26348,N_25976);
and U26561 (N_26561,N_26323,N_25992);
nor U26562 (N_26562,N_26108,N_26168);
and U26563 (N_26563,N_25999,N_26174);
and U26564 (N_26564,N_26320,N_25996);
nor U26565 (N_26565,N_25854,N_25979);
and U26566 (N_26566,N_26316,N_25900);
nand U26567 (N_26567,N_25966,N_25931);
nor U26568 (N_26568,N_26013,N_26020);
and U26569 (N_26569,N_26200,N_25973);
nand U26570 (N_26570,N_26140,N_26043);
or U26571 (N_26571,N_26199,N_26378);
nor U26572 (N_26572,N_26288,N_25860);
and U26573 (N_26573,N_25913,N_25971);
and U26574 (N_26574,N_25990,N_26181);
nor U26575 (N_26575,N_26227,N_26252);
nor U26576 (N_26576,N_26158,N_26074);
and U26577 (N_26577,N_26109,N_26201);
nand U26578 (N_26578,N_26188,N_26290);
nand U26579 (N_26579,N_26038,N_25839);
or U26580 (N_26580,N_26012,N_25876);
nand U26581 (N_26581,N_26296,N_26283);
and U26582 (N_26582,N_26175,N_26071);
nor U26583 (N_26583,N_26036,N_25884);
nand U26584 (N_26584,N_26202,N_26368);
nor U26585 (N_26585,N_25811,N_26072);
nand U26586 (N_26586,N_26017,N_26046);
nand U26587 (N_26587,N_26387,N_26233);
nor U26588 (N_26588,N_26304,N_26091);
and U26589 (N_26589,N_26266,N_25827);
nor U26590 (N_26590,N_25922,N_25889);
nor U26591 (N_26591,N_26076,N_26376);
nand U26592 (N_26592,N_25829,N_25923);
nand U26593 (N_26593,N_25866,N_25898);
nor U26594 (N_26594,N_26055,N_26373);
nor U26595 (N_26595,N_25918,N_26149);
nor U26596 (N_26596,N_25886,N_26107);
nand U26597 (N_26597,N_26302,N_25981);
nor U26598 (N_26598,N_26070,N_25893);
and U26599 (N_26599,N_26178,N_25985);
nor U26600 (N_26600,N_25890,N_26274);
and U26601 (N_26601,N_25831,N_26123);
and U26602 (N_26602,N_26147,N_25987);
nand U26603 (N_26603,N_25844,N_25813);
and U26604 (N_26604,N_26228,N_25993);
nor U26605 (N_26605,N_25840,N_26067);
or U26606 (N_26606,N_25938,N_26122);
xnor U26607 (N_26607,N_26338,N_25950);
or U26608 (N_26608,N_26052,N_26186);
xnor U26609 (N_26609,N_25954,N_25952);
nand U26610 (N_26610,N_26231,N_25805);
and U26611 (N_26611,N_25822,N_25887);
and U26612 (N_26612,N_26394,N_25857);
nand U26613 (N_26613,N_25984,N_25891);
or U26614 (N_26614,N_26030,N_25819);
nor U26615 (N_26615,N_26031,N_26118);
nand U26616 (N_26616,N_26393,N_26116);
and U26617 (N_26617,N_25880,N_26268);
or U26618 (N_26618,N_26129,N_26063);
nand U26619 (N_26619,N_26023,N_26026);
nand U26620 (N_26620,N_26385,N_25914);
and U26621 (N_26621,N_26212,N_25997);
and U26622 (N_26622,N_25941,N_26362);
and U26623 (N_26623,N_26001,N_26349);
or U26624 (N_26624,N_26124,N_25989);
nor U26625 (N_26625,N_26223,N_26197);
nor U26626 (N_26626,N_26066,N_26379);
nor U26627 (N_26627,N_25972,N_26333);
xnor U26628 (N_26628,N_26382,N_26180);
and U26629 (N_26629,N_26241,N_26356);
and U26630 (N_26630,N_25843,N_26261);
or U26631 (N_26631,N_26134,N_26148);
nor U26632 (N_26632,N_25937,N_26322);
xnor U26633 (N_26633,N_26137,N_26000);
nand U26634 (N_26634,N_26146,N_25951);
and U26635 (N_26635,N_26151,N_26315);
and U26636 (N_26636,N_26395,N_25859);
and U26637 (N_26637,N_26159,N_26167);
nor U26638 (N_26638,N_26190,N_26165);
nand U26639 (N_26639,N_26359,N_26236);
and U26640 (N_26640,N_26347,N_25957);
nand U26641 (N_26641,N_26263,N_26234);
nand U26642 (N_26642,N_26044,N_26057);
nand U26643 (N_26643,N_26112,N_26279);
nor U26644 (N_26644,N_25858,N_26377);
and U26645 (N_26645,N_26317,N_26328);
nor U26646 (N_26646,N_25908,N_25961);
or U26647 (N_26647,N_26213,N_26217);
nor U26648 (N_26648,N_25915,N_26343);
nand U26649 (N_26649,N_26354,N_26157);
and U26650 (N_26650,N_26281,N_26047);
nand U26651 (N_26651,N_25928,N_26239);
nand U26652 (N_26652,N_25801,N_26332);
or U26653 (N_26653,N_25837,N_26136);
nand U26654 (N_26654,N_26309,N_25868);
nand U26655 (N_26655,N_26007,N_26214);
nand U26656 (N_26656,N_26021,N_26106);
and U26657 (N_26657,N_26265,N_26285);
or U26658 (N_26658,N_26398,N_25956);
nor U26659 (N_26659,N_26205,N_26310);
nand U26660 (N_26660,N_25855,N_25832);
or U26661 (N_26661,N_26247,N_26004);
nand U26662 (N_26662,N_25942,N_26390);
nand U26663 (N_26663,N_25856,N_26273);
or U26664 (N_26664,N_26114,N_26270);
nand U26665 (N_26665,N_25929,N_26100);
nand U26666 (N_26666,N_26278,N_25906);
or U26667 (N_26667,N_25983,N_26120);
and U26668 (N_26668,N_26262,N_26364);
nand U26669 (N_26669,N_26367,N_26032);
and U26670 (N_26670,N_26392,N_26282);
and U26671 (N_26671,N_25806,N_26225);
nand U26672 (N_26672,N_25896,N_25960);
nand U26673 (N_26673,N_26130,N_26370);
or U26674 (N_26674,N_26080,N_26185);
or U26675 (N_26675,N_26245,N_25852);
or U26676 (N_26676,N_26048,N_26327);
nand U26677 (N_26677,N_26391,N_25943);
nand U26678 (N_26678,N_26125,N_26272);
nor U26679 (N_26679,N_25847,N_26132);
nand U26680 (N_26680,N_26077,N_25802);
nand U26681 (N_26681,N_26305,N_26386);
xnor U26682 (N_26682,N_26297,N_26346);
nand U26683 (N_26683,N_26277,N_26160);
and U26684 (N_26684,N_26105,N_26085);
and U26685 (N_26685,N_26194,N_26184);
nor U26686 (N_26686,N_26331,N_26014);
or U26687 (N_26687,N_25924,N_26141);
and U26688 (N_26688,N_26041,N_25878);
nor U26689 (N_26689,N_26135,N_26257);
nor U26690 (N_26690,N_26179,N_26126);
and U26691 (N_26691,N_25864,N_25867);
nor U26692 (N_26692,N_25869,N_25953);
nor U26693 (N_26693,N_26271,N_26049);
nand U26694 (N_26694,N_26101,N_26015);
nand U26695 (N_26695,N_26301,N_25846);
or U26696 (N_26696,N_26170,N_25902);
nand U26697 (N_26697,N_25970,N_26319);
or U26698 (N_26698,N_25815,N_25826);
nand U26699 (N_26699,N_26255,N_26351);
nor U26700 (N_26700,N_26081,N_25993);
nor U26701 (N_26701,N_26198,N_26283);
nand U26702 (N_26702,N_25859,N_26187);
and U26703 (N_26703,N_26043,N_26282);
or U26704 (N_26704,N_25967,N_26245);
xor U26705 (N_26705,N_26313,N_26120);
and U26706 (N_26706,N_25873,N_26378);
or U26707 (N_26707,N_26096,N_26388);
nor U26708 (N_26708,N_26279,N_26175);
or U26709 (N_26709,N_25921,N_26320);
and U26710 (N_26710,N_26269,N_26301);
nand U26711 (N_26711,N_25887,N_26287);
and U26712 (N_26712,N_25948,N_26280);
nand U26713 (N_26713,N_26376,N_25908);
and U26714 (N_26714,N_26172,N_25804);
nor U26715 (N_26715,N_26202,N_26144);
and U26716 (N_26716,N_26274,N_26028);
and U26717 (N_26717,N_26326,N_26153);
or U26718 (N_26718,N_25846,N_26353);
nand U26719 (N_26719,N_25993,N_26215);
nor U26720 (N_26720,N_25985,N_26029);
nand U26721 (N_26721,N_26065,N_26280);
or U26722 (N_26722,N_25934,N_25973);
and U26723 (N_26723,N_26352,N_25950);
nor U26724 (N_26724,N_26296,N_25832);
nand U26725 (N_26725,N_26043,N_26223);
nor U26726 (N_26726,N_26254,N_26338);
or U26727 (N_26727,N_25949,N_25948);
nor U26728 (N_26728,N_26357,N_26264);
or U26729 (N_26729,N_26357,N_26309);
and U26730 (N_26730,N_25932,N_26363);
or U26731 (N_26731,N_25840,N_26025);
or U26732 (N_26732,N_26362,N_26150);
nand U26733 (N_26733,N_26124,N_26202);
nand U26734 (N_26734,N_26077,N_26257);
or U26735 (N_26735,N_26133,N_26238);
nand U26736 (N_26736,N_26070,N_25805);
xor U26737 (N_26737,N_26170,N_25811);
nor U26738 (N_26738,N_25938,N_26178);
and U26739 (N_26739,N_26205,N_26124);
nand U26740 (N_26740,N_25912,N_26373);
and U26741 (N_26741,N_25809,N_26107);
and U26742 (N_26742,N_26228,N_26016);
nand U26743 (N_26743,N_25954,N_26371);
and U26744 (N_26744,N_26048,N_26304);
or U26745 (N_26745,N_26196,N_25941);
nand U26746 (N_26746,N_26005,N_25976);
nand U26747 (N_26747,N_25847,N_25968);
and U26748 (N_26748,N_26043,N_25855);
nand U26749 (N_26749,N_25911,N_26018);
nor U26750 (N_26750,N_25946,N_25952);
nand U26751 (N_26751,N_26209,N_25885);
nor U26752 (N_26752,N_25864,N_25819);
and U26753 (N_26753,N_25901,N_26189);
nor U26754 (N_26754,N_26225,N_26014);
and U26755 (N_26755,N_25913,N_26041);
nand U26756 (N_26756,N_26311,N_26153);
nor U26757 (N_26757,N_25885,N_26350);
and U26758 (N_26758,N_25817,N_26201);
nand U26759 (N_26759,N_26164,N_26359);
nand U26760 (N_26760,N_25889,N_25820);
and U26761 (N_26761,N_26118,N_26357);
or U26762 (N_26762,N_25929,N_26130);
or U26763 (N_26763,N_25815,N_26217);
and U26764 (N_26764,N_26138,N_26321);
nand U26765 (N_26765,N_26249,N_26008);
nor U26766 (N_26766,N_26127,N_25887);
nand U26767 (N_26767,N_25976,N_26264);
nor U26768 (N_26768,N_25820,N_26218);
or U26769 (N_26769,N_26192,N_26062);
or U26770 (N_26770,N_26357,N_26221);
and U26771 (N_26771,N_26333,N_26214);
or U26772 (N_26772,N_25823,N_26227);
or U26773 (N_26773,N_26116,N_25801);
nand U26774 (N_26774,N_25913,N_26011);
xor U26775 (N_26775,N_25900,N_26310);
or U26776 (N_26776,N_26183,N_26289);
and U26777 (N_26777,N_25853,N_26148);
and U26778 (N_26778,N_26330,N_26074);
and U26779 (N_26779,N_26336,N_26101);
nor U26780 (N_26780,N_26379,N_26129);
nand U26781 (N_26781,N_25883,N_26226);
nor U26782 (N_26782,N_25929,N_26186);
nand U26783 (N_26783,N_25914,N_25936);
and U26784 (N_26784,N_26234,N_25962);
nor U26785 (N_26785,N_25900,N_26282);
or U26786 (N_26786,N_26265,N_26398);
or U26787 (N_26787,N_26188,N_26289);
or U26788 (N_26788,N_26060,N_26301);
nor U26789 (N_26789,N_26158,N_26398);
nand U26790 (N_26790,N_26147,N_25924);
and U26791 (N_26791,N_26004,N_26190);
nor U26792 (N_26792,N_26178,N_26272);
and U26793 (N_26793,N_25869,N_26174);
nor U26794 (N_26794,N_26331,N_25965);
or U26795 (N_26795,N_26302,N_26379);
or U26796 (N_26796,N_26082,N_26184);
nor U26797 (N_26797,N_25822,N_26033);
nand U26798 (N_26798,N_26335,N_26087);
or U26799 (N_26799,N_26331,N_26183);
nor U26800 (N_26800,N_26118,N_26002);
and U26801 (N_26801,N_26011,N_26118);
nor U26802 (N_26802,N_25839,N_26204);
nand U26803 (N_26803,N_25991,N_25972);
nor U26804 (N_26804,N_26257,N_25989);
nand U26805 (N_26805,N_26235,N_26045);
nor U26806 (N_26806,N_25940,N_26140);
nand U26807 (N_26807,N_26125,N_26380);
or U26808 (N_26808,N_25894,N_26352);
and U26809 (N_26809,N_26195,N_25859);
nor U26810 (N_26810,N_26120,N_26110);
nor U26811 (N_26811,N_25812,N_25959);
nand U26812 (N_26812,N_26254,N_26196);
nor U26813 (N_26813,N_26135,N_26177);
nand U26814 (N_26814,N_25892,N_26347);
nor U26815 (N_26815,N_26343,N_25901);
and U26816 (N_26816,N_26376,N_26096);
nand U26817 (N_26817,N_26263,N_26254);
and U26818 (N_26818,N_25820,N_25910);
and U26819 (N_26819,N_25836,N_26221);
nand U26820 (N_26820,N_26029,N_25957);
and U26821 (N_26821,N_26201,N_26155);
nand U26822 (N_26822,N_25865,N_25942);
and U26823 (N_26823,N_25824,N_25812);
or U26824 (N_26824,N_26300,N_26196);
and U26825 (N_26825,N_26351,N_26115);
nand U26826 (N_26826,N_26195,N_26120);
and U26827 (N_26827,N_25939,N_26344);
nand U26828 (N_26828,N_25977,N_25817);
and U26829 (N_26829,N_26372,N_26238);
nor U26830 (N_26830,N_25846,N_26112);
and U26831 (N_26831,N_26139,N_26106);
and U26832 (N_26832,N_26364,N_25917);
nor U26833 (N_26833,N_25935,N_26371);
nand U26834 (N_26834,N_26399,N_25857);
nor U26835 (N_26835,N_25897,N_26276);
nor U26836 (N_26836,N_26130,N_26291);
or U26837 (N_26837,N_26040,N_26106);
and U26838 (N_26838,N_26180,N_26337);
xor U26839 (N_26839,N_26070,N_26114);
or U26840 (N_26840,N_25837,N_25911);
nor U26841 (N_26841,N_26309,N_26083);
and U26842 (N_26842,N_26256,N_25916);
nor U26843 (N_26843,N_26378,N_26186);
nand U26844 (N_26844,N_25913,N_26167);
and U26845 (N_26845,N_25996,N_26164);
nand U26846 (N_26846,N_26348,N_26232);
nor U26847 (N_26847,N_26038,N_25864);
or U26848 (N_26848,N_26352,N_26306);
or U26849 (N_26849,N_25818,N_25938);
and U26850 (N_26850,N_26347,N_26047);
or U26851 (N_26851,N_25925,N_26385);
nor U26852 (N_26852,N_26270,N_25887);
or U26853 (N_26853,N_26098,N_26127);
nor U26854 (N_26854,N_26194,N_26274);
or U26855 (N_26855,N_25817,N_26081);
nand U26856 (N_26856,N_25917,N_26313);
and U26857 (N_26857,N_26248,N_25945);
or U26858 (N_26858,N_25849,N_25857);
and U26859 (N_26859,N_26322,N_26079);
or U26860 (N_26860,N_26162,N_26012);
or U26861 (N_26861,N_25832,N_26166);
nand U26862 (N_26862,N_25971,N_26092);
nand U26863 (N_26863,N_26184,N_26390);
and U26864 (N_26864,N_26324,N_25927);
nor U26865 (N_26865,N_26190,N_26230);
and U26866 (N_26866,N_25938,N_26088);
and U26867 (N_26867,N_26131,N_26146);
or U26868 (N_26868,N_25847,N_26218);
and U26869 (N_26869,N_25877,N_26050);
nand U26870 (N_26870,N_26387,N_26052);
nor U26871 (N_26871,N_26353,N_26328);
nor U26872 (N_26872,N_25979,N_26303);
nand U26873 (N_26873,N_25988,N_26226);
and U26874 (N_26874,N_26378,N_26132);
nor U26875 (N_26875,N_26111,N_26177);
nand U26876 (N_26876,N_25813,N_25909);
or U26877 (N_26877,N_26205,N_26197);
nand U26878 (N_26878,N_26104,N_25891);
nand U26879 (N_26879,N_26258,N_26106);
nor U26880 (N_26880,N_26040,N_25938);
nand U26881 (N_26881,N_26174,N_25962);
nand U26882 (N_26882,N_26031,N_26335);
nor U26883 (N_26883,N_26371,N_26287);
nor U26884 (N_26884,N_26114,N_25807);
and U26885 (N_26885,N_26378,N_26338);
nor U26886 (N_26886,N_25923,N_25900);
nand U26887 (N_26887,N_25842,N_26346);
and U26888 (N_26888,N_25818,N_26347);
and U26889 (N_26889,N_26375,N_26022);
or U26890 (N_26890,N_25966,N_26220);
nor U26891 (N_26891,N_26112,N_26213);
and U26892 (N_26892,N_26315,N_26316);
and U26893 (N_26893,N_25927,N_26183);
nor U26894 (N_26894,N_25872,N_25868);
nand U26895 (N_26895,N_25958,N_25855);
and U26896 (N_26896,N_26056,N_25978);
or U26897 (N_26897,N_26143,N_26220);
or U26898 (N_26898,N_26298,N_26142);
nor U26899 (N_26899,N_26243,N_25935);
nand U26900 (N_26900,N_25836,N_26164);
nand U26901 (N_26901,N_25925,N_25874);
nor U26902 (N_26902,N_25884,N_26131);
and U26903 (N_26903,N_26285,N_26267);
nand U26904 (N_26904,N_26044,N_26258);
and U26905 (N_26905,N_26188,N_25961);
or U26906 (N_26906,N_26314,N_26290);
nor U26907 (N_26907,N_25906,N_26136);
and U26908 (N_26908,N_26375,N_25865);
and U26909 (N_26909,N_26148,N_26312);
or U26910 (N_26910,N_25875,N_26188);
nor U26911 (N_26911,N_26387,N_26024);
nand U26912 (N_26912,N_26058,N_26283);
nand U26913 (N_26913,N_26320,N_26208);
xor U26914 (N_26914,N_26069,N_26368);
or U26915 (N_26915,N_25887,N_26144);
nand U26916 (N_26916,N_26148,N_25902);
and U26917 (N_26917,N_25943,N_26019);
or U26918 (N_26918,N_26285,N_25855);
and U26919 (N_26919,N_25881,N_25906);
nor U26920 (N_26920,N_25928,N_26041);
or U26921 (N_26921,N_26016,N_26115);
or U26922 (N_26922,N_25866,N_25922);
or U26923 (N_26923,N_25802,N_26391);
or U26924 (N_26924,N_26180,N_25813);
nor U26925 (N_26925,N_26258,N_26388);
or U26926 (N_26926,N_26143,N_26036);
nand U26927 (N_26927,N_26193,N_26210);
or U26928 (N_26928,N_26382,N_26392);
and U26929 (N_26929,N_25827,N_26282);
nand U26930 (N_26930,N_25903,N_25996);
or U26931 (N_26931,N_26308,N_26057);
nand U26932 (N_26932,N_26306,N_25860);
xor U26933 (N_26933,N_26126,N_26275);
and U26934 (N_26934,N_25889,N_26110);
and U26935 (N_26935,N_25975,N_26376);
nand U26936 (N_26936,N_25914,N_26208);
and U26937 (N_26937,N_26296,N_26325);
or U26938 (N_26938,N_26258,N_25868);
or U26939 (N_26939,N_26348,N_26123);
and U26940 (N_26940,N_26171,N_25878);
nor U26941 (N_26941,N_26380,N_26002);
or U26942 (N_26942,N_25996,N_26081);
nand U26943 (N_26943,N_26173,N_25934);
nor U26944 (N_26944,N_26368,N_25945);
nand U26945 (N_26945,N_25984,N_26195);
nor U26946 (N_26946,N_26391,N_26246);
and U26947 (N_26947,N_25985,N_26039);
and U26948 (N_26948,N_26255,N_25979);
nand U26949 (N_26949,N_25994,N_26085);
nor U26950 (N_26950,N_25943,N_26280);
nor U26951 (N_26951,N_25885,N_25868);
nor U26952 (N_26952,N_26021,N_26307);
or U26953 (N_26953,N_26016,N_25966);
nor U26954 (N_26954,N_26137,N_26128);
nor U26955 (N_26955,N_25943,N_26194);
or U26956 (N_26956,N_26273,N_25879);
nor U26957 (N_26957,N_26264,N_25970);
or U26958 (N_26958,N_25984,N_25922);
nor U26959 (N_26959,N_26318,N_26252);
or U26960 (N_26960,N_26009,N_25931);
and U26961 (N_26961,N_25939,N_25843);
nand U26962 (N_26962,N_26207,N_25943);
or U26963 (N_26963,N_26098,N_26155);
and U26964 (N_26964,N_26256,N_25860);
nor U26965 (N_26965,N_26156,N_26274);
or U26966 (N_26966,N_26076,N_26240);
and U26967 (N_26967,N_25866,N_25989);
and U26968 (N_26968,N_26130,N_26105);
nor U26969 (N_26969,N_26130,N_25989);
and U26970 (N_26970,N_26101,N_26320);
nand U26971 (N_26971,N_26192,N_26113);
nand U26972 (N_26972,N_25904,N_26287);
nor U26973 (N_26973,N_26129,N_25999);
nor U26974 (N_26974,N_25999,N_25989);
nand U26975 (N_26975,N_26264,N_26296);
and U26976 (N_26976,N_26186,N_26372);
or U26977 (N_26977,N_25964,N_26221);
and U26978 (N_26978,N_25879,N_26104);
and U26979 (N_26979,N_25831,N_25952);
nand U26980 (N_26980,N_26085,N_26311);
or U26981 (N_26981,N_26384,N_25813);
or U26982 (N_26982,N_25857,N_26092);
nand U26983 (N_26983,N_26371,N_26246);
and U26984 (N_26984,N_26343,N_26141);
and U26985 (N_26985,N_26288,N_26225);
nor U26986 (N_26986,N_26007,N_26382);
nand U26987 (N_26987,N_26017,N_26379);
or U26988 (N_26988,N_26058,N_26267);
nor U26989 (N_26989,N_26095,N_26381);
nand U26990 (N_26990,N_25908,N_26000);
and U26991 (N_26991,N_26182,N_26240);
xor U26992 (N_26992,N_26253,N_26096);
nand U26993 (N_26993,N_26231,N_26370);
and U26994 (N_26994,N_25932,N_26318);
and U26995 (N_26995,N_26348,N_26338);
xnor U26996 (N_26996,N_26204,N_26168);
nand U26997 (N_26997,N_26065,N_25940);
nor U26998 (N_26998,N_26365,N_25937);
nor U26999 (N_26999,N_26302,N_26143);
nand U27000 (N_27000,N_26608,N_26637);
nand U27001 (N_27001,N_26772,N_26931);
and U27002 (N_27002,N_26694,N_26783);
nand U27003 (N_27003,N_26537,N_26746);
nand U27004 (N_27004,N_26603,N_26950);
and U27005 (N_27005,N_26564,N_26526);
or U27006 (N_27006,N_26509,N_26992);
or U27007 (N_27007,N_26575,N_26978);
nand U27008 (N_27008,N_26627,N_26579);
or U27009 (N_27009,N_26623,N_26458);
xnor U27010 (N_27010,N_26493,N_26883);
nand U27011 (N_27011,N_26695,N_26501);
or U27012 (N_27012,N_26704,N_26766);
nor U27013 (N_27013,N_26962,N_26860);
nor U27014 (N_27014,N_26632,N_26634);
nand U27015 (N_27015,N_26787,N_26503);
and U27016 (N_27016,N_26845,N_26409);
or U27017 (N_27017,N_26643,N_26780);
or U27018 (N_27018,N_26825,N_26764);
nand U27019 (N_27019,N_26555,N_26854);
nor U27020 (N_27020,N_26915,N_26818);
nor U27021 (N_27021,N_26817,N_26923);
nand U27022 (N_27022,N_26420,N_26431);
or U27023 (N_27023,N_26686,N_26466);
and U27024 (N_27024,N_26789,N_26943);
nor U27025 (N_27025,N_26903,N_26816);
nor U27026 (N_27026,N_26901,N_26546);
nand U27027 (N_27027,N_26940,N_26538);
or U27028 (N_27028,N_26582,N_26613);
or U27029 (N_27029,N_26678,N_26917);
nor U27030 (N_27030,N_26957,N_26455);
nor U27031 (N_27031,N_26497,N_26664);
nor U27032 (N_27032,N_26451,N_26986);
or U27033 (N_27033,N_26449,N_26658);
and U27034 (N_27034,N_26720,N_26732);
and U27035 (N_27035,N_26887,N_26747);
or U27036 (N_27036,N_26463,N_26697);
or U27037 (N_27037,N_26750,N_26976);
or U27038 (N_27038,N_26610,N_26738);
or U27039 (N_27039,N_26606,N_26562);
nand U27040 (N_27040,N_26857,N_26706);
nand U27041 (N_27041,N_26459,N_26897);
or U27042 (N_27042,N_26598,N_26511);
nor U27043 (N_27043,N_26536,N_26479);
nor U27044 (N_27044,N_26487,N_26784);
and U27045 (N_27045,N_26419,N_26909);
nand U27046 (N_27046,N_26837,N_26760);
nor U27047 (N_27047,N_26997,N_26922);
or U27048 (N_27048,N_26660,N_26970);
or U27049 (N_27049,N_26989,N_26731);
and U27050 (N_27050,N_26871,N_26651);
or U27051 (N_27051,N_26902,N_26592);
and U27052 (N_27052,N_26404,N_26400);
nor U27053 (N_27053,N_26947,N_26440);
xnor U27054 (N_27054,N_26979,N_26771);
nand U27055 (N_27055,N_26645,N_26799);
xnor U27056 (N_27056,N_26937,N_26904);
xor U27057 (N_27057,N_26494,N_26763);
and U27058 (N_27058,N_26891,N_26878);
nand U27059 (N_27059,N_26552,N_26585);
and U27060 (N_27060,N_26462,N_26519);
xor U27061 (N_27061,N_26587,N_26896);
nand U27062 (N_27062,N_26718,N_26846);
nor U27063 (N_27063,N_26406,N_26926);
and U27064 (N_27064,N_26507,N_26952);
nand U27065 (N_27065,N_26499,N_26522);
or U27066 (N_27066,N_26630,N_26412);
and U27067 (N_27067,N_26557,N_26534);
nand U27068 (N_27068,N_26659,N_26864);
or U27069 (N_27069,N_26551,N_26910);
nand U27070 (N_27070,N_26713,N_26468);
and U27071 (N_27071,N_26432,N_26516);
and U27072 (N_27072,N_26452,N_26402);
and U27073 (N_27073,N_26595,N_26828);
nor U27074 (N_27074,N_26542,N_26918);
and U27075 (N_27075,N_26682,N_26850);
or U27076 (N_27076,N_26733,N_26607);
nor U27077 (N_27077,N_26792,N_26527);
or U27078 (N_27078,N_26426,N_26653);
nor U27079 (N_27079,N_26712,N_26584);
nor U27080 (N_27080,N_26528,N_26888);
or U27081 (N_27081,N_26486,N_26473);
and U27082 (N_27082,N_26510,N_26749);
nor U27083 (N_27083,N_26898,N_26863);
or U27084 (N_27084,N_26401,N_26959);
nor U27085 (N_27085,N_26728,N_26958);
nor U27086 (N_27086,N_26570,N_26853);
nor U27087 (N_27087,N_26998,N_26944);
or U27088 (N_27088,N_26841,N_26647);
nor U27089 (N_27089,N_26740,N_26561);
and U27090 (N_27090,N_26965,N_26635);
nor U27091 (N_27091,N_26921,N_26521);
and U27092 (N_27092,N_26422,N_26525);
or U27093 (N_27093,N_26933,N_26788);
nand U27094 (N_27094,N_26960,N_26942);
or U27095 (N_27095,N_26945,N_26985);
and U27096 (N_27096,N_26457,N_26681);
or U27097 (N_27097,N_26470,N_26886);
or U27098 (N_27098,N_26756,N_26672);
and U27099 (N_27099,N_26671,N_26652);
xor U27100 (N_27100,N_26812,N_26905);
nand U27101 (N_27101,N_26482,N_26867);
nand U27102 (N_27102,N_26714,N_26434);
or U27103 (N_27103,N_26725,N_26670);
nand U27104 (N_27104,N_26474,N_26791);
nand U27105 (N_27105,N_26790,N_26796);
nand U27106 (N_27106,N_26924,N_26831);
nand U27107 (N_27107,N_26578,N_26589);
or U27108 (N_27108,N_26549,N_26977);
and U27109 (N_27109,N_26815,N_26934);
nand U27110 (N_27110,N_26530,N_26558);
and U27111 (N_27111,N_26734,N_26702);
or U27112 (N_27112,N_26705,N_26990);
or U27113 (N_27113,N_26775,N_26781);
nand U27114 (N_27114,N_26456,N_26810);
and U27115 (N_27115,N_26410,N_26951);
and U27116 (N_27116,N_26506,N_26644);
and U27117 (N_27117,N_26767,N_26852);
nor U27118 (N_27118,N_26475,N_26491);
or U27119 (N_27119,N_26488,N_26826);
nand U27120 (N_27120,N_26742,N_26648);
nor U27121 (N_27121,N_26829,N_26948);
xor U27122 (N_27122,N_26827,N_26708);
nor U27123 (N_27123,N_26569,N_26877);
and U27124 (N_27124,N_26502,N_26735);
and U27125 (N_27125,N_26498,N_26436);
nand U27126 (N_27126,N_26604,N_26984);
nand U27127 (N_27127,N_26759,N_26531);
and U27128 (N_27128,N_26469,N_26983);
nand U27129 (N_27129,N_26722,N_26638);
nor U27130 (N_27130,N_26515,N_26936);
and U27131 (N_27131,N_26752,N_26885);
or U27132 (N_27132,N_26969,N_26701);
nor U27133 (N_27133,N_26529,N_26851);
nand U27134 (N_27134,N_26471,N_26941);
nor U27135 (N_27135,N_26689,N_26961);
nor U27136 (N_27136,N_26920,N_26566);
and U27137 (N_27137,N_26517,N_26927);
nor U27138 (N_27138,N_26880,N_26698);
or U27139 (N_27139,N_26461,N_26797);
nand U27140 (N_27140,N_26541,N_26744);
or U27141 (N_27141,N_26547,N_26865);
and U27142 (N_27142,N_26571,N_26687);
and U27143 (N_27143,N_26626,N_26559);
xor U27144 (N_27144,N_26593,N_26548);
or U27145 (N_27145,N_26594,N_26999);
nor U27146 (N_27146,N_26963,N_26809);
and U27147 (N_27147,N_26472,N_26618);
nor U27148 (N_27148,N_26971,N_26974);
nor U27149 (N_27149,N_26667,N_26408);
or U27150 (N_27150,N_26615,N_26741);
nor U27151 (N_27151,N_26478,N_26893);
nand U27152 (N_27152,N_26715,N_26862);
and U27153 (N_27153,N_26612,N_26655);
nor U27154 (N_27154,N_26485,N_26730);
or U27155 (N_27155,N_26418,N_26554);
or U27156 (N_27156,N_26576,N_26964);
and U27157 (N_27157,N_26794,N_26691);
nor U27158 (N_27158,N_26504,N_26629);
or U27159 (N_27159,N_26801,N_26512);
nor U27160 (N_27160,N_26609,N_26840);
nand U27161 (N_27161,N_26938,N_26911);
nand U27162 (N_27162,N_26523,N_26813);
or U27163 (N_27163,N_26711,N_26914);
and U27164 (N_27164,N_26811,N_26761);
or U27165 (N_27165,N_26786,N_26447);
nand U27166 (N_27166,N_26916,N_26968);
and U27167 (N_27167,N_26520,N_26777);
nand U27168 (N_27168,N_26617,N_26778);
and U27169 (N_27169,N_26641,N_26876);
nand U27170 (N_27170,N_26873,N_26821);
nand U27171 (N_27171,N_26939,N_26439);
nor U27172 (N_27172,N_26535,N_26484);
xor U27173 (N_27173,N_26858,N_26601);
and U27174 (N_27174,N_26954,N_26673);
or U27175 (N_27175,N_26892,N_26993);
or U27176 (N_27176,N_26636,N_26755);
xnor U27177 (N_27177,N_26518,N_26745);
nor U27178 (N_27178,N_26567,N_26573);
nor U27179 (N_27179,N_26805,N_26707);
xnor U27180 (N_27180,N_26605,N_26727);
or U27181 (N_27181,N_26824,N_26692);
nor U27182 (N_27182,N_26500,N_26913);
and U27183 (N_27183,N_26649,N_26847);
or U27184 (N_27184,N_26429,N_26416);
and U27185 (N_27185,N_26650,N_26631);
and U27186 (N_27186,N_26717,N_26513);
nand U27187 (N_27187,N_26577,N_26413);
and U27188 (N_27188,N_26869,N_26848);
and U27189 (N_27189,N_26748,N_26699);
nand U27190 (N_27190,N_26987,N_26928);
nor U27191 (N_27191,N_26785,N_26590);
nor U27192 (N_27192,N_26804,N_26540);
and U27193 (N_27193,N_26830,N_26640);
nor U27194 (N_27194,N_26953,N_26981);
nand U27195 (N_27195,N_26553,N_26693);
nand U27196 (N_27196,N_26683,N_26996);
and U27197 (N_27197,N_26421,N_26628);
and U27198 (N_27198,N_26820,N_26675);
nor U27199 (N_27199,N_26622,N_26556);
or U27200 (N_27200,N_26688,N_26442);
and U27201 (N_27201,N_26460,N_26435);
and U27202 (N_27202,N_26855,N_26890);
nor U27203 (N_27203,N_26586,N_26879);
or U27204 (N_27204,N_26620,N_26762);
nor U27205 (N_27205,N_26899,N_26550);
and U27206 (N_27206,N_26773,N_26405);
nand U27207 (N_27207,N_26972,N_26476);
nand U27208 (N_27208,N_26543,N_26669);
and U27209 (N_27209,N_26446,N_26441);
nor U27210 (N_27210,N_26430,N_26793);
nor U27211 (N_27211,N_26657,N_26591);
nor U27212 (N_27212,N_26425,N_26754);
nand U27213 (N_27213,N_26737,N_26619);
or U27214 (N_27214,N_26674,N_26870);
nor U27215 (N_27215,N_26490,N_26802);
nor U27216 (N_27216,N_26882,N_26489);
or U27217 (N_27217,N_26800,N_26895);
nor U27218 (N_27218,N_26465,N_26685);
or U27219 (N_27219,N_26616,N_26417);
nor U27220 (N_27220,N_26467,N_26611);
nand U27221 (N_27221,N_26776,N_26665);
nor U27222 (N_27222,N_26625,N_26668);
and U27223 (N_27223,N_26581,N_26819);
nor U27224 (N_27224,N_26690,N_26836);
nand U27225 (N_27225,N_26495,N_26995);
nand U27226 (N_27226,N_26724,N_26900);
nor U27227 (N_27227,N_26803,N_26935);
nor U27228 (N_27228,N_26496,N_26600);
and U27229 (N_27229,N_26729,N_26753);
and U27230 (N_27230,N_26889,N_26843);
nor U27231 (N_27231,N_26574,N_26834);
and U27232 (N_27232,N_26709,N_26700);
nor U27233 (N_27233,N_26765,N_26403);
and U27234 (N_27234,N_26925,N_26443);
nor U27235 (N_27235,N_26842,N_26743);
nor U27236 (N_27236,N_26415,N_26768);
and U27237 (N_27237,N_26838,N_26975);
and U27238 (N_27238,N_26407,N_26454);
and U27239 (N_27239,N_26477,N_26438);
or U27240 (N_27240,N_26894,N_26769);
nor U27241 (N_27241,N_26833,N_26483);
nand U27242 (N_27242,N_26808,N_26532);
or U27243 (N_27243,N_26946,N_26912);
nor U27244 (N_27244,N_26849,N_26423);
and U27245 (N_27245,N_26450,N_26861);
nand U27246 (N_27246,N_26716,N_26624);
nor U27247 (N_27247,N_26654,N_26583);
and U27248 (N_27248,N_26437,N_26994);
or U27249 (N_27249,N_26621,N_26949);
or U27250 (N_27250,N_26684,N_26433);
nand U27251 (N_27251,N_26444,N_26874);
and U27252 (N_27252,N_26982,N_26736);
or U27253 (N_27253,N_26588,N_26774);
nor U27254 (N_27254,N_26696,N_26967);
nor U27255 (N_27255,N_26480,N_26806);
nor U27256 (N_27256,N_26908,N_26560);
or U27257 (N_27257,N_26875,N_26448);
nand U27258 (N_27258,N_26907,N_26524);
and U27259 (N_27259,N_26411,N_26666);
or U27260 (N_27260,N_26703,N_26719);
and U27261 (N_27261,N_26453,N_26661);
or U27262 (N_27262,N_26710,N_26991);
nand U27263 (N_27263,N_26881,N_26544);
nand U27264 (N_27264,N_26424,N_26505);
or U27265 (N_27265,N_26597,N_26872);
and U27266 (N_27266,N_26614,N_26427);
nand U27267 (N_27267,N_26906,N_26642);
nor U27268 (N_27268,N_26966,N_26795);
nand U27269 (N_27269,N_26539,N_26980);
nand U27270 (N_27270,N_26599,N_26835);
and U27271 (N_27271,N_26757,N_26758);
nor U27272 (N_27272,N_26770,N_26866);
and U27273 (N_27273,N_26639,N_26508);
nor U27274 (N_27274,N_26930,N_26751);
nand U27275 (N_27275,N_26677,N_26533);
nand U27276 (N_27276,N_26572,N_26839);
nor U27277 (N_27277,N_26563,N_26602);
nor U27278 (N_27278,N_26988,N_26832);
and U27279 (N_27279,N_26721,N_26823);
nor U27280 (N_27280,N_26856,N_26868);
and U27281 (N_27281,N_26633,N_26428);
and U27282 (N_27282,N_26568,N_26565);
or U27283 (N_27283,N_26723,N_26932);
nand U27284 (N_27284,N_26545,N_26956);
and U27285 (N_27285,N_26662,N_26726);
and U27286 (N_27286,N_26739,N_26859);
and U27287 (N_27287,N_26464,N_26646);
and U27288 (N_27288,N_26663,N_26679);
or U27289 (N_27289,N_26676,N_26844);
nand U27290 (N_27290,N_26884,N_26919);
nor U27291 (N_27291,N_26414,N_26929);
nand U27292 (N_27292,N_26481,N_26445);
xor U27293 (N_27293,N_26656,N_26814);
nand U27294 (N_27294,N_26779,N_26680);
nor U27295 (N_27295,N_26782,N_26973);
nand U27296 (N_27296,N_26822,N_26596);
or U27297 (N_27297,N_26514,N_26955);
or U27298 (N_27298,N_26580,N_26492);
and U27299 (N_27299,N_26807,N_26798);
nand U27300 (N_27300,N_26961,N_26510);
nand U27301 (N_27301,N_26751,N_26463);
and U27302 (N_27302,N_26415,N_26752);
nand U27303 (N_27303,N_26579,N_26706);
nor U27304 (N_27304,N_26558,N_26817);
and U27305 (N_27305,N_26911,N_26629);
nand U27306 (N_27306,N_26430,N_26637);
or U27307 (N_27307,N_26680,N_26593);
nand U27308 (N_27308,N_26417,N_26765);
or U27309 (N_27309,N_26656,N_26541);
or U27310 (N_27310,N_26595,N_26485);
or U27311 (N_27311,N_26672,N_26481);
nand U27312 (N_27312,N_26610,N_26538);
nand U27313 (N_27313,N_26551,N_26553);
or U27314 (N_27314,N_26647,N_26838);
and U27315 (N_27315,N_26943,N_26413);
nor U27316 (N_27316,N_26814,N_26486);
and U27317 (N_27317,N_26802,N_26995);
nand U27318 (N_27318,N_26788,N_26978);
nand U27319 (N_27319,N_26549,N_26889);
or U27320 (N_27320,N_26574,N_26716);
nor U27321 (N_27321,N_26677,N_26692);
or U27322 (N_27322,N_26564,N_26439);
nor U27323 (N_27323,N_26642,N_26766);
nand U27324 (N_27324,N_26604,N_26719);
or U27325 (N_27325,N_26482,N_26973);
or U27326 (N_27326,N_26942,N_26723);
and U27327 (N_27327,N_26815,N_26917);
and U27328 (N_27328,N_26809,N_26563);
xor U27329 (N_27329,N_26531,N_26682);
or U27330 (N_27330,N_26808,N_26971);
nand U27331 (N_27331,N_26876,N_26473);
nor U27332 (N_27332,N_26681,N_26782);
nor U27333 (N_27333,N_26977,N_26763);
nor U27334 (N_27334,N_26685,N_26470);
or U27335 (N_27335,N_26803,N_26815);
nand U27336 (N_27336,N_26635,N_26483);
and U27337 (N_27337,N_26483,N_26859);
nand U27338 (N_27338,N_26495,N_26639);
nand U27339 (N_27339,N_26923,N_26596);
nor U27340 (N_27340,N_26560,N_26746);
and U27341 (N_27341,N_26509,N_26564);
or U27342 (N_27342,N_26632,N_26717);
nand U27343 (N_27343,N_26854,N_26531);
or U27344 (N_27344,N_26556,N_26918);
or U27345 (N_27345,N_26618,N_26776);
nor U27346 (N_27346,N_26405,N_26607);
or U27347 (N_27347,N_26633,N_26984);
or U27348 (N_27348,N_26712,N_26713);
or U27349 (N_27349,N_26712,N_26591);
nand U27350 (N_27350,N_26976,N_26760);
nor U27351 (N_27351,N_26571,N_26553);
nand U27352 (N_27352,N_26420,N_26888);
nand U27353 (N_27353,N_26828,N_26486);
nor U27354 (N_27354,N_26940,N_26481);
and U27355 (N_27355,N_26983,N_26519);
and U27356 (N_27356,N_26466,N_26950);
or U27357 (N_27357,N_26651,N_26951);
nor U27358 (N_27358,N_26934,N_26568);
and U27359 (N_27359,N_26629,N_26714);
nor U27360 (N_27360,N_26507,N_26914);
nor U27361 (N_27361,N_26695,N_26456);
nand U27362 (N_27362,N_26447,N_26628);
or U27363 (N_27363,N_26833,N_26781);
and U27364 (N_27364,N_26808,N_26425);
nor U27365 (N_27365,N_26495,N_26569);
nor U27366 (N_27366,N_26417,N_26689);
nor U27367 (N_27367,N_26979,N_26854);
nor U27368 (N_27368,N_26959,N_26728);
nand U27369 (N_27369,N_26702,N_26466);
nor U27370 (N_27370,N_26431,N_26870);
or U27371 (N_27371,N_26521,N_26665);
and U27372 (N_27372,N_26493,N_26628);
or U27373 (N_27373,N_26492,N_26839);
and U27374 (N_27374,N_26577,N_26491);
and U27375 (N_27375,N_26609,N_26545);
and U27376 (N_27376,N_26855,N_26947);
and U27377 (N_27377,N_26460,N_26975);
and U27378 (N_27378,N_26828,N_26623);
nor U27379 (N_27379,N_26679,N_26685);
or U27380 (N_27380,N_26780,N_26894);
nand U27381 (N_27381,N_26726,N_26883);
nand U27382 (N_27382,N_26639,N_26708);
nand U27383 (N_27383,N_26784,N_26777);
or U27384 (N_27384,N_26497,N_26778);
and U27385 (N_27385,N_26727,N_26405);
nand U27386 (N_27386,N_26802,N_26518);
and U27387 (N_27387,N_26623,N_26456);
and U27388 (N_27388,N_26402,N_26424);
and U27389 (N_27389,N_26999,N_26750);
or U27390 (N_27390,N_26545,N_26409);
or U27391 (N_27391,N_26505,N_26535);
xnor U27392 (N_27392,N_26489,N_26834);
nand U27393 (N_27393,N_26686,N_26897);
or U27394 (N_27394,N_26967,N_26440);
and U27395 (N_27395,N_26838,N_26427);
nand U27396 (N_27396,N_26704,N_26726);
or U27397 (N_27397,N_26726,N_26739);
or U27398 (N_27398,N_26889,N_26691);
nor U27399 (N_27399,N_26764,N_26743);
and U27400 (N_27400,N_26519,N_26809);
and U27401 (N_27401,N_26569,N_26732);
and U27402 (N_27402,N_26741,N_26579);
and U27403 (N_27403,N_26431,N_26560);
nor U27404 (N_27404,N_26826,N_26423);
nor U27405 (N_27405,N_26462,N_26918);
or U27406 (N_27406,N_26783,N_26558);
and U27407 (N_27407,N_26443,N_26524);
nor U27408 (N_27408,N_26777,N_26476);
nor U27409 (N_27409,N_26480,N_26927);
or U27410 (N_27410,N_26661,N_26959);
nand U27411 (N_27411,N_26746,N_26469);
and U27412 (N_27412,N_26542,N_26693);
nor U27413 (N_27413,N_26665,N_26476);
nand U27414 (N_27414,N_26821,N_26704);
and U27415 (N_27415,N_26543,N_26623);
and U27416 (N_27416,N_26633,N_26451);
or U27417 (N_27417,N_26799,N_26691);
nor U27418 (N_27418,N_26887,N_26652);
or U27419 (N_27419,N_26956,N_26895);
nand U27420 (N_27420,N_26795,N_26679);
and U27421 (N_27421,N_26437,N_26557);
nor U27422 (N_27422,N_26583,N_26445);
or U27423 (N_27423,N_26913,N_26541);
or U27424 (N_27424,N_26962,N_26886);
or U27425 (N_27425,N_26526,N_26733);
and U27426 (N_27426,N_26833,N_26680);
nor U27427 (N_27427,N_26847,N_26819);
nand U27428 (N_27428,N_26766,N_26767);
and U27429 (N_27429,N_26762,N_26471);
or U27430 (N_27430,N_26839,N_26827);
nand U27431 (N_27431,N_26631,N_26986);
or U27432 (N_27432,N_26468,N_26561);
nor U27433 (N_27433,N_26699,N_26972);
and U27434 (N_27434,N_26474,N_26632);
nor U27435 (N_27435,N_26463,N_26402);
and U27436 (N_27436,N_26481,N_26789);
nand U27437 (N_27437,N_26617,N_26574);
xnor U27438 (N_27438,N_26985,N_26863);
nand U27439 (N_27439,N_26589,N_26741);
nor U27440 (N_27440,N_26696,N_26853);
or U27441 (N_27441,N_26989,N_26465);
and U27442 (N_27442,N_26511,N_26477);
nand U27443 (N_27443,N_26582,N_26784);
nor U27444 (N_27444,N_26527,N_26562);
nand U27445 (N_27445,N_26607,N_26968);
and U27446 (N_27446,N_26499,N_26400);
nor U27447 (N_27447,N_26903,N_26807);
and U27448 (N_27448,N_26416,N_26524);
nand U27449 (N_27449,N_26540,N_26773);
or U27450 (N_27450,N_26927,N_26746);
or U27451 (N_27451,N_26465,N_26979);
and U27452 (N_27452,N_26569,N_26512);
and U27453 (N_27453,N_26923,N_26705);
nand U27454 (N_27454,N_26866,N_26544);
and U27455 (N_27455,N_26462,N_26588);
and U27456 (N_27456,N_26795,N_26927);
or U27457 (N_27457,N_26713,N_26811);
nand U27458 (N_27458,N_26576,N_26593);
nor U27459 (N_27459,N_26663,N_26977);
and U27460 (N_27460,N_26968,N_26834);
nor U27461 (N_27461,N_26401,N_26688);
nand U27462 (N_27462,N_26496,N_26881);
or U27463 (N_27463,N_26657,N_26887);
nand U27464 (N_27464,N_26670,N_26663);
xnor U27465 (N_27465,N_26745,N_26727);
nor U27466 (N_27466,N_26782,N_26928);
and U27467 (N_27467,N_26620,N_26775);
nand U27468 (N_27468,N_26986,N_26985);
nor U27469 (N_27469,N_26615,N_26442);
nand U27470 (N_27470,N_26803,N_26939);
nand U27471 (N_27471,N_26718,N_26642);
nand U27472 (N_27472,N_26770,N_26441);
or U27473 (N_27473,N_26935,N_26521);
and U27474 (N_27474,N_26907,N_26670);
and U27475 (N_27475,N_26989,N_26466);
or U27476 (N_27476,N_26785,N_26532);
nor U27477 (N_27477,N_26499,N_26787);
or U27478 (N_27478,N_26623,N_26694);
nand U27479 (N_27479,N_26639,N_26802);
or U27480 (N_27480,N_26931,N_26916);
or U27481 (N_27481,N_26502,N_26664);
nor U27482 (N_27482,N_26961,N_26727);
and U27483 (N_27483,N_26611,N_26553);
nor U27484 (N_27484,N_26502,N_26436);
and U27485 (N_27485,N_26926,N_26403);
or U27486 (N_27486,N_26419,N_26862);
nor U27487 (N_27487,N_26679,N_26748);
nor U27488 (N_27488,N_26510,N_26703);
nor U27489 (N_27489,N_26756,N_26534);
nor U27490 (N_27490,N_26837,N_26556);
and U27491 (N_27491,N_26504,N_26924);
xnor U27492 (N_27492,N_26704,N_26463);
nor U27493 (N_27493,N_26677,N_26414);
and U27494 (N_27494,N_26570,N_26708);
nor U27495 (N_27495,N_26771,N_26630);
nand U27496 (N_27496,N_26475,N_26474);
or U27497 (N_27497,N_26930,N_26465);
nand U27498 (N_27498,N_26625,N_26582);
and U27499 (N_27499,N_26789,N_26614);
nand U27500 (N_27500,N_26501,N_26741);
nor U27501 (N_27501,N_26884,N_26897);
nand U27502 (N_27502,N_26841,N_26654);
or U27503 (N_27503,N_26687,N_26499);
nor U27504 (N_27504,N_26430,N_26880);
and U27505 (N_27505,N_26912,N_26461);
nand U27506 (N_27506,N_26713,N_26478);
nor U27507 (N_27507,N_26887,N_26630);
nor U27508 (N_27508,N_26600,N_26887);
nand U27509 (N_27509,N_26534,N_26814);
xnor U27510 (N_27510,N_26744,N_26439);
nand U27511 (N_27511,N_26908,N_26763);
and U27512 (N_27512,N_26433,N_26937);
nor U27513 (N_27513,N_26415,N_26951);
and U27514 (N_27514,N_26527,N_26746);
or U27515 (N_27515,N_26821,N_26459);
nand U27516 (N_27516,N_26861,N_26572);
nor U27517 (N_27517,N_26462,N_26671);
nand U27518 (N_27518,N_26544,N_26614);
and U27519 (N_27519,N_26707,N_26418);
nand U27520 (N_27520,N_26977,N_26865);
or U27521 (N_27521,N_26826,N_26847);
nand U27522 (N_27522,N_26636,N_26493);
and U27523 (N_27523,N_26654,N_26515);
nor U27524 (N_27524,N_26617,N_26739);
nand U27525 (N_27525,N_26547,N_26717);
nor U27526 (N_27526,N_26496,N_26415);
and U27527 (N_27527,N_26634,N_26481);
nand U27528 (N_27528,N_26851,N_26461);
nor U27529 (N_27529,N_26572,N_26946);
nand U27530 (N_27530,N_26619,N_26842);
nand U27531 (N_27531,N_26961,N_26921);
nor U27532 (N_27532,N_26815,N_26674);
or U27533 (N_27533,N_26931,N_26958);
nor U27534 (N_27534,N_26771,N_26668);
nor U27535 (N_27535,N_26450,N_26714);
nand U27536 (N_27536,N_26799,N_26869);
or U27537 (N_27537,N_26612,N_26765);
nor U27538 (N_27538,N_26904,N_26558);
nand U27539 (N_27539,N_26819,N_26622);
nor U27540 (N_27540,N_26805,N_26659);
xor U27541 (N_27541,N_26850,N_26992);
nand U27542 (N_27542,N_26890,N_26769);
and U27543 (N_27543,N_26677,N_26867);
nor U27544 (N_27544,N_26880,N_26461);
and U27545 (N_27545,N_26935,N_26559);
or U27546 (N_27546,N_26672,N_26906);
nand U27547 (N_27547,N_26616,N_26948);
xor U27548 (N_27548,N_26960,N_26613);
nor U27549 (N_27549,N_26800,N_26646);
and U27550 (N_27550,N_26869,N_26647);
nor U27551 (N_27551,N_26889,N_26670);
nor U27552 (N_27552,N_26441,N_26889);
nand U27553 (N_27553,N_26524,N_26478);
or U27554 (N_27554,N_26989,N_26799);
or U27555 (N_27555,N_26565,N_26792);
nor U27556 (N_27556,N_26637,N_26624);
xnor U27557 (N_27557,N_26400,N_26531);
nor U27558 (N_27558,N_26934,N_26957);
nand U27559 (N_27559,N_26576,N_26777);
nor U27560 (N_27560,N_26579,N_26732);
or U27561 (N_27561,N_26974,N_26488);
or U27562 (N_27562,N_26934,N_26758);
or U27563 (N_27563,N_26481,N_26808);
nand U27564 (N_27564,N_26529,N_26891);
nor U27565 (N_27565,N_26876,N_26798);
or U27566 (N_27566,N_26874,N_26968);
nor U27567 (N_27567,N_26472,N_26588);
and U27568 (N_27568,N_26646,N_26772);
nand U27569 (N_27569,N_26651,N_26760);
nand U27570 (N_27570,N_26779,N_26873);
and U27571 (N_27571,N_26975,N_26453);
and U27572 (N_27572,N_26805,N_26522);
or U27573 (N_27573,N_26560,N_26980);
or U27574 (N_27574,N_26590,N_26626);
nand U27575 (N_27575,N_26905,N_26872);
nand U27576 (N_27576,N_26983,N_26891);
xor U27577 (N_27577,N_26859,N_26752);
or U27578 (N_27578,N_26776,N_26492);
and U27579 (N_27579,N_26690,N_26728);
nor U27580 (N_27580,N_26939,N_26936);
or U27581 (N_27581,N_26827,N_26403);
or U27582 (N_27582,N_26491,N_26742);
and U27583 (N_27583,N_26606,N_26779);
nor U27584 (N_27584,N_26955,N_26825);
nor U27585 (N_27585,N_26785,N_26562);
and U27586 (N_27586,N_26753,N_26980);
and U27587 (N_27587,N_26845,N_26834);
nand U27588 (N_27588,N_26720,N_26639);
xnor U27589 (N_27589,N_26777,N_26420);
nand U27590 (N_27590,N_26818,N_26992);
nand U27591 (N_27591,N_26718,N_26913);
nor U27592 (N_27592,N_26413,N_26771);
nor U27593 (N_27593,N_26417,N_26794);
and U27594 (N_27594,N_26600,N_26429);
nor U27595 (N_27595,N_26985,N_26806);
nor U27596 (N_27596,N_26967,N_26851);
xnor U27597 (N_27597,N_26653,N_26681);
and U27598 (N_27598,N_26981,N_26491);
nand U27599 (N_27599,N_26482,N_26504);
nand U27600 (N_27600,N_27488,N_27498);
and U27601 (N_27601,N_27076,N_27565);
or U27602 (N_27602,N_27579,N_27454);
nor U27603 (N_27603,N_27172,N_27094);
or U27604 (N_27604,N_27194,N_27478);
nor U27605 (N_27605,N_27267,N_27244);
or U27606 (N_27606,N_27345,N_27415);
xor U27607 (N_27607,N_27093,N_27066);
nor U27608 (N_27608,N_27239,N_27477);
nor U27609 (N_27609,N_27279,N_27189);
nor U27610 (N_27610,N_27551,N_27596);
nor U27611 (N_27611,N_27143,N_27206);
or U27612 (N_27612,N_27136,N_27504);
or U27613 (N_27613,N_27264,N_27408);
or U27614 (N_27614,N_27395,N_27115);
and U27615 (N_27615,N_27424,N_27035);
nand U27616 (N_27616,N_27423,N_27384);
nor U27617 (N_27617,N_27253,N_27195);
nand U27618 (N_27618,N_27528,N_27274);
and U27619 (N_27619,N_27526,N_27305);
nand U27620 (N_27620,N_27499,N_27221);
nor U27621 (N_27621,N_27460,N_27063);
or U27622 (N_27622,N_27134,N_27226);
or U27623 (N_27623,N_27242,N_27394);
nor U27624 (N_27624,N_27339,N_27398);
xor U27625 (N_27625,N_27150,N_27317);
or U27626 (N_27626,N_27257,N_27450);
and U27627 (N_27627,N_27016,N_27427);
nor U27628 (N_27628,N_27381,N_27315);
nand U27629 (N_27629,N_27467,N_27482);
or U27630 (N_27630,N_27042,N_27179);
nand U27631 (N_27631,N_27263,N_27040);
and U27632 (N_27632,N_27425,N_27410);
or U27633 (N_27633,N_27569,N_27506);
or U27634 (N_27634,N_27089,N_27282);
or U27635 (N_27635,N_27404,N_27533);
or U27636 (N_27636,N_27350,N_27457);
nand U27637 (N_27637,N_27503,N_27186);
or U27638 (N_27638,N_27047,N_27534);
or U27639 (N_27639,N_27046,N_27392);
or U27640 (N_27640,N_27241,N_27210);
nand U27641 (N_27641,N_27366,N_27320);
nor U27642 (N_27642,N_27070,N_27472);
or U27643 (N_27643,N_27535,N_27587);
or U27644 (N_27644,N_27441,N_27309);
and U27645 (N_27645,N_27031,N_27289);
or U27646 (N_27646,N_27388,N_27474);
and U27647 (N_27647,N_27589,N_27111);
nand U27648 (N_27648,N_27081,N_27168);
nand U27649 (N_27649,N_27208,N_27343);
or U27650 (N_27650,N_27352,N_27301);
nand U27651 (N_27651,N_27418,N_27517);
or U27652 (N_27652,N_27481,N_27029);
nor U27653 (N_27653,N_27298,N_27543);
and U27654 (N_27654,N_27167,N_27220);
xnor U27655 (N_27655,N_27399,N_27306);
and U27656 (N_27656,N_27575,N_27269);
nor U27657 (N_27657,N_27536,N_27583);
and U27658 (N_27658,N_27148,N_27018);
and U27659 (N_27659,N_27156,N_27416);
or U27660 (N_27660,N_27494,N_27108);
nand U27661 (N_27661,N_27280,N_27554);
nor U27662 (N_27662,N_27329,N_27211);
nor U27663 (N_27663,N_27538,N_27207);
nand U27664 (N_27664,N_27513,N_27495);
and U27665 (N_27665,N_27281,N_27004);
xor U27666 (N_27666,N_27276,N_27200);
and U27667 (N_27667,N_27285,N_27248);
nand U27668 (N_27668,N_27173,N_27165);
and U27669 (N_27669,N_27458,N_27097);
and U27670 (N_27670,N_27130,N_27434);
and U27671 (N_27671,N_27542,N_27255);
nand U27672 (N_27672,N_27584,N_27344);
or U27673 (N_27673,N_27175,N_27303);
or U27674 (N_27674,N_27419,N_27369);
xnor U27675 (N_27675,N_27116,N_27166);
nand U27676 (N_27676,N_27041,N_27030);
nand U27677 (N_27677,N_27372,N_27044);
and U27678 (N_27678,N_27393,N_27162);
or U27679 (N_27679,N_27591,N_27573);
or U27680 (N_27680,N_27412,N_27247);
nor U27681 (N_27681,N_27377,N_27414);
nand U27682 (N_27682,N_27256,N_27451);
nand U27683 (N_27683,N_27515,N_27155);
nor U27684 (N_27684,N_27530,N_27523);
and U27685 (N_27685,N_27198,N_27260);
nor U27686 (N_27686,N_27297,N_27293);
nor U27687 (N_27687,N_27171,N_27382);
and U27688 (N_27688,N_27012,N_27368);
or U27689 (N_27689,N_27456,N_27176);
nand U27690 (N_27690,N_27120,N_27238);
and U27691 (N_27691,N_27237,N_27592);
nand U27692 (N_27692,N_27100,N_27110);
nor U27693 (N_27693,N_27378,N_27582);
nor U27694 (N_27694,N_27400,N_27578);
nand U27695 (N_27695,N_27421,N_27181);
or U27696 (N_27696,N_27015,N_27502);
or U27697 (N_27697,N_27532,N_27231);
nand U27698 (N_27698,N_27122,N_27401);
and U27699 (N_27699,N_27158,N_27058);
and U27700 (N_27700,N_27205,N_27354);
nand U27701 (N_27701,N_27261,N_27327);
nor U27702 (N_27702,N_27001,N_27054);
or U27703 (N_27703,N_27202,N_27539);
nand U27704 (N_27704,N_27307,N_27213);
nand U27705 (N_27705,N_27489,N_27288);
and U27706 (N_27706,N_27357,N_27483);
or U27707 (N_27707,N_27013,N_27531);
or U27708 (N_27708,N_27347,N_27223);
nor U27709 (N_27709,N_27006,N_27032);
and U27710 (N_27710,N_27585,N_27520);
nor U27711 (N_27711,N_27373,N_27518);
or U27712 (N_27712,N_27364,N_27091);
nand U27713 (N_27713,N_27275,N_27118);
nor U27714 (N_27714,N_27462,N_27199);
xnor U27715 (N_27715,N_27077,N_27152);
and U27716 (N_27716,N_27137,N_27092);
nand U27717 (N_27717,N_27020,N_27335);
or U27718 (N_27718,N_27363,N_27505);
or U27719 (N_27719,N_27568,N_27045);
or U27720 (N_27720,N_27153,N_27028);
or U27721 (N_27721,N_27486,N_27272);
or U27722 (N_27722,N_27529,N_27567);
and U27723 (N_27723,N_27413,N_27246);
nor U27724 (N_27724,N_27430,N_27014);
or U27725 (N_27725,N_27580,N_27227);
nand U27726 (N_27726,N_27034,N_27022);
nor U27727 (N_27727,N_27558,N_27559);
nand U27728 (N_27728,N_27300,N_27487);
nor U27729 (N_27729,N_27426,N_27403);
nand U27730 (N_27730,N_27455,N_27201);
nand U27731 (N_27731,N_27524,N_27552);
nor U27732 (N_27732,N_27062,N_27113);
and U27733 (N_27733,N_27229,N_27109);
nor U27734 (N_27734,N_27129,N_27406);
nand U27735 (N_27735,N_27106,N_27117);
nor U27736 (N_27736,N_27501,N_27316);
or U27737 (N_27737,N_27590,N_27361);
or U27738 (N_27738,N_27114,N_27563);
nor U27739 (N_27739,N_27145,N_27271);
nand U27740 (N_27740,N_27180,N_27519);
nand U27741 (N_27741,N_27544,N_27283);
nor U27742 (N_27742,N_27000,N_27250);
nor U27743 (N_27743,N_27371,N_27052);
and U27744 (N_27744,N_27314,N_27219);
and U27745 (N_27745,N_27490,N_27313);
and U27746 (N_27746,N_27449,N_27429);
or U27747 (N_27747,N_27154,N_27119);
nand U27748 (N_27748,N_27196,N_27164);
nor U27749 (N_27749,N_27353,N_27102);
nor U27750 (N_27750,N_27023,N_27096);
nor U27751 (N_27751,N_27078,N_27508);
nand U27752 (N_27752,N_27026,N_27184);
nor U27753 (N_27753,N_27330,N_27243);
xnor U27754 (N_27754,N_27389,N_27514);
nor U27755 (N_27755,N_27209,N_27473);
and U27756 (N_27756,N_27555,N_27254);
nand U27757 (N_27757,N_27431,N_27376);
nor U27758 (N_27758,N_27038,N_27516);
nor U27759 (N_27759,N_27436,N_27442);
nand U27760 (N_27760,N_27547,N_27411);
or U27761 (N_27761,N_27445,N_27385);
nand U27762 (N_27762,N_27349,N_27095);
nand U27763 (N_27763,N_27358,N_27541);
nand U27764 (N_27764,N_27021,N_27571);
or U27765 (N_27765,N_27079,N_27290);
nand U27766 (N_27766,N_27562,N_27367);
xor U27767 (N_27767,N_27512,N_27295);
nand U27768 (N_27768,N_27010,N_27332);
nand U27769 (N_27769,N_27557,N_27187);
xnor U27770 (N_27770,N_27230,N_27391);
nand U27771 (N_27771,N_27548,N_27598);
and U27772 (N_27772,N_27304,N_27071);
nor U27773 (N_27773,N_27140,N_27333);
nor U27774 (N_27774,N_27127,N_27435);
or U27775 (N_27775,N_27461,N_27005);
nor U27776 (N_27776,N_27566,N_27123);
nand U27777 (N_27777,N_27380,N_27178);
nor U27778 (N_27778,N_27322,N_27121);
nor U27779 (N_27779,N_27310,N_27294);
or U27780 (N_27780,N_27278,N_27024);
nand U27781 (N_27781,N_27439,N_27053);
nor U27782 (N_27782,N_27375,N_27011);
nand U27783 (N_27783,N_27002,N_27074);
and U27784 (N_27784,N_27521,N_27438);
and U27785 (N_27785,N_27234,N_27059);
or U27786 (N_27786,N_27328,N_27417);
nand U27787 (N_27787,N_27139,N_27323);
or U27788 (N_27788,N_27588,N_27204);
and U27789 (N_27789,N_27463,N_27446);
or U27790 (N_27790,N_27193,N_27217);
or U27791 (N_27791,N_27064,N_27510);
nand U27792 (N_27792,N_27480,N_27594);
nand U27793 (N_27793,N_27008,N_27469);
nor U27794 (N_27794,N_27222,N_27550);
or U27795 (N_27795,N_27009,N_27485);
xnor U27796 (N_27796,N_27497,N_27556);
nand U27797 (N_27797,N_27465,N_27577);
and U27798 (N_27798,N_27479,N_27390);
and U27799 (N_27799,N_27067,N_27270);
or U27800 (N_27800,N_27311,N_27496);
nand U27801 (N_27801,N_27225,N_27336);
nand U27802 (N_27802,N_27599,N_27087);
and U27803 (N_27803,N_27007,N_27266);
nor U27804 (N_27804,N_27214,N_27525);
nand U27805 (N_27805,N_27459,N_27075);
nand U27806 (N_27806,N_27387,N_27080);
nand U27807 (N_27807,N_27055,N_27084);
and U27808 (N_27808,N_27287,N_27537);
or U27809 (N_27809,N_27337,N_27043);
nand U27810 (N_27810,N_27561,N_27228);
xnor U27811 (N_27811,N_27192,N_27112);
nor U27812 (N_27812,N_27174,N_27037);
nor U27813 (N_27813,N_27397,N_27105);
nand U27814 (N_27814,N_27493,N_27470);
and U27815 (N_27815,N_27265,N_27099);
or U27816 (N_27816,N_27331,N_27197);
or U27817 (N_27817,N_27017,N_27453);
or U27818 (N_27818,N_27593,N_27432);
or U27819 (N_27819,N_27341,N_27235);
nand U27820 (N_27820,N_27048,N_27149);
nor U27821 (N_27821,N_27348,N_27082);
and U27822 (N_27822,N_27386,N_27507);
nand U27823 (N_27823,N_27259,N_27161);
nand U27824 (N_27824,N_27128,N_27428);
nand U27825 (N_27825,N_27103,N_27284);
and U27826 (N_27826,N_27351,N_27360);
and U27827 (N_27827,N_27564,N_27019);
or U27828 (N_27828,N_27324,N_27232);
and U27829 (N_27829,N_27437,N_27060);
nor U27830 (N_27830,N_27182,N_27597);
or U27831 (N_27831,N_27218,N_27402);
nand U27832 (N_27832,N_27144,N_27422);
nor U27833 (N_27833,N_27586,N_27160);
and U27834 (N_27834,N_27433,N_27346);
nand U27835 (N_27835,N_27069,N_27302);
nor U27836 (N_27836,N_27407,N_27240);
and U27837 (N_27837,N_27342,N_27522);
nor U27838 (N_27838,N_27133,N_27468);
nand U27839 (N_27839,N_27251,N_27101);
or U27840 (N_27840,N_27057,N_27088);
nor U27841 (N_27841,N_27546,N_27545);
and U27842 (N_27842,N_27319,N_27471);
nand U27843 (N_27843,N_27374,N_27065);
nor U27844 (N_27844,N_27056,N_27595);
nor U27845 (N_27845,N_27159,N_27203);
or U27846 (N_27846,N_27448,N_27420);
nor U27847 (N_27847,N_27245,N_27560);
nand U27848 (N_27848,N_27572,N_27258);
or U27849 (N_27849,N_27553,N_27540);
or U27850 (N_27850,N_27039,N_27308);
and U27851 (N_27851,N_27190,N_27447);
nand U27852 (N_27852,N_27334,N_27292);
or U27853 (N_27853,N_27135,N_27355);
nand U27854 (N_27854,N_27085,N_27025);
nor U27855 (N_27855,N_27444,N_27003);
nand U27856 (N_27856,N_27236,N_27291);
nand U27857 (N_27857,N_27409,N_27338);
and U27858 (N_27858,N_27191,N_27252);
and U27859 (N_27859,N_27027,N_27326);
nand U27860 (N_27860,N_27132,N_27475);
or U27861 (N_27861,N_27452,N_27464);
nor U27862 (N_27862,N_27492,N_27147);
and U27863 (N_27863,N_27356,N_27511);
or U27864 (N_27864,N_27359,N_27509);
nand U27865 (N_27865,N_27405,N_27273);
and U27866 (N_27866,N_27170,N_27365);
nor U27867 (N_27867,N_27268,N_27576);
nor U27868 (N_27868,N_27146,N_27296);
or U27869 (N_27869,N_27491,N_27050);
xor U27870 (N_27870,N_27484,N_27383);
or U27871 (N_27871,N_27090,N_27188);
nand U27872 (N_27872,N_27277,N_27466);
or U27873 (N_27873,N_27299,N_27443);
or U27874 (N_27874,N_27224,N_27216);
nor U27875 (N_27875,N_27312,N_27169);
or U27876 (N_27876,N_27125,N_27362);
nor U27877 (N_27877,N_27212,N_27370);
nand U27878 (N_27878,N_27131,N_27138);
and U27879 (N_27879,N_27379,N_27440);
nor U27880 (N_27880,N_27036,N_27157);
or U27881 (N_27881,N_27215,N_27104);
or U27882 (N_27882,N_27325,N_27086);
nor U27883 (N_27883,N_27286,N_27396);
and U27884 (N_27884,N_27318,N_27051);
nor U27885 (N_27885,N_27581,N_27107);
or U27886 (N_27886,N_27177,N_27141);
nor U27887 (N_27887,N_27527,N_27340);
or U27888 (N_27888,N_27072,N_27249);
nor U27889 (N_27889,N_27073,N_27083);
nand U27890 (N_27890,N_27570,N_27233);
and U27891 (N_27891,N_27068,N_27098);
nor U27892 (N_27892,N_27476,N_27124);
nand U27893 (N_27893,N_27500,N_27033);
or U27894 (N_27894,N_27574,N_27151);
or U27895 (N_27895,N_27142,N_27049);
nand U27896 (N_27896,N_27321,N_27262);
or U27897 (N_27897,N_27183,N_27126);
or U27898 (N_27898,N_27163,N_27061);
and U27899 (N_27899,N_27185,N_27549);
nor U27900 (N_27900,N_27504,N_27096);
xor U27901 (N_27901,N_27284,N_27224);
or U27902 (N_27902,N_27005,N_27002);
or U27903 (N_27903,N_27185,N_27592);
and U27904 (N_27904,N_27403,N_27192);
nor U27905 (N_27905,N_27514,N_27065);
or U27906 (N_27906,N_27563,N_27528);
nand U27907 (N_27907,N_27387,N_27465);
nor U27908 (N_27908,N_27216,N_27139);
nand U27909 (N_27909,N_27332,N_27553);
nand U27910 (N_27910,N_27236,N_27055);
nor U27911 (N_27911,N_27470,N_27585);
nor U27912 (N_27912,N_27225,N_27593);
xor U27913 (N_27913,N_27212,N_27310);
xor U27914 (N_27914,N_27357,N_27319);
nor U27915 (N_27915,N_27072,N_27118);
nand U27916 (N_27916,N_27144,N_27339);
nor U27917 (N_27917,N_27013,N_27070);
or U27918 (N_27918,N_27248,N_27287);
and U27919 (N_27919,N_27382,N_27545);
or U27920 (N_27920,N_27162,N_27163);
nor U27921 (N_27921,N_27134,N_27290);
and U27922 (N_27922,N_27366,N_27352);
nor U27923 (N_27923,N_27077,N_27492);
or U27924 (N_27924,N_27440,N_27362);
and U27925 (N_27925,N_27193,N_27117);
and U27926 (N_27926,N_27169,N_27481);
or U27927 (N_27927,N_27272,N_27546);
nand U27928 (N_27928,N_27547,N_27225);
or U27929 (N_27929,N_27143,N_27266);
or U27930 (N_27930,N_27291,N_27010);
and U27931 (N_27931,N_27253,N_27104);
nand U27932 (N_27932,N_27272,N_27315);
nand U27933 (N_27933,N_27052,N_27024);
nor U27934 (N_27934,N_27366,N_27177);
nand U27935 (N_27935,N_27446,N_27028);
or U27936 (N_27936,N_27416,N_27443);
or U27937 (N_27937,N_27380,N_27127);
or U27938 (N_27938,N_27194,N_27021);
nor U27939 (N_27939,N_27530,N_27341);
and U27940 (N_27940,N_27038,N_27387);
nor U27941 (N_27941,N_27552,N_27060);
or U27942 (N_27942,N_27546,N_27174);
nor U27943 (N_27943,N_27122,N_27372);
and U27944 (N_27944,N_27466,N_27241);
nor U27945 (N_27945,N_27342,N_27191);
or U27946 (N_27946,N_27411,N_27057);
and U27947 (N_27947,N_27345,N_27506);
nand U27948 (N_27948,N_27204,N_27178);
nand U27949 (N_27949,N_27292,N_27444);
nor U27950 (N_27950,N_27045,N_27021);
and U27951 (N_27951,N_27256,N_27045);
nand U27952 (N_27952,N_27386,N_27573);
nand U27953 (N_27953,N_27587,N_27585);
and U27954 (N_27954,N_27120,N_27182);
or U27955 (N_27955,N_27363,N_27199);
nand U27956 (N_27956,N_27057,N_27453);
and U27957 (N_27957,N_27139,N_27198);
nand U27958 (N_27958,N_27407,N_27162);
nor U27959 (N_27959,N_27484,N_27018);
nor U27960 (N_27960,N_27032,N_27055);
nor U27961 (N_27961,N_27555,N_27210);
nor U27962 (N_27962,N_27060,N_27438);
and U27963 (N_27963,N_27450,N_27144);
nor U27964 (N_27964,N_27283,N_27576);
or U27965 (N_27965,N_27007,N_27223);
or U27966 (N_27966,N_27270,N_27433);
and U27967 (N_27967,N_27252,N_27515);
or U27968 (N_27968,N_27458,N_27027);
and U27969 (N_27969,N_27127,N_27035);
and U27970 (N_27970,N_27434,N_27503);
nor U27971 (N_27971,N_27317,N_27292);
nor U27972 (N_27972,N_27522,N_27396);
or U27973 (N_27973,N_27132,N_27078);
and U27974 (N_27974,N_27074,N_27052);
and U27975 (N_27975,N_27161,N_27264);
nor U27976 (N_27976,N_27378,N_27097);
and U27977 (N_27977,N_27244,N_27090);
nand U27978 (N_27978,N_27512,N_27151);
nor U27979 (N_27979,N_27366,N_27444);
nor U27980 (N_27980,N_27450,N_27095);
or U27981 (N_27981,N_27390,N_27365);
nand U27982 (N_27982,N_27376,N_27326);
nand U27983 (N_27983,N_27286,N_27108);
nor U27984 (N_27984,N_27036,N_27455);
and U27985 (N_27985,N_27079,N_27018);
nand U27986 (N_27986,N_27306,N_27551);
nor U27987 (N_27987,N_27153,N_27400);
nor U27988 (N_27988,N_27442,N_27544);
or U27989 (N_27989,N_27062,N_27588);
nand U27990 (N_27990,N_27142,N_27341);
or U27991 (N_27991,N_27495,N_27406);
or U27992 (N_27992,N_27173,N_27377);
nand U27993 (N_27993,N_27132,N_27315);
or U27994 (N_27994,N_27045,N_27348);
nand U27995 (N_27995,N_27451,N_27405);
nor U27996 (N_27996,N_27217,N_27592);
or U27997 (N_27997,N_27417,N_27041);
and U27998 (N_27998,N_27005,N_27477);
nor U27999 (N_27999,N_27304,N_27516);
and U28000 (N_28000,N_27199,N_27358);
or U28001 (N_28001,N_27131,N_27573);
and U28002 (N_28002,N_27127,N_27249);
or U28003 (N_28003,N_27056,N_27128);
nand U28004 (N_28004,N_27196,N_27388);
or U28005 (N_28005,N_27009,N_27368);
and U28006 (N_28006,N_27143,N_27120);
nand U28007 (N_28007,N_27098,N_27572);
nor U28008 (N_28008,N_27064,N_27321);
nand U28009 (N_28009,N_27234,N_27339);
nor U28010 (N_28010,N_27429,N_27417);
or U28011 (N_28011,N_27355,N_27513);
nand U28012 (N_28012,N_27559,N_27202);
nand U28013 (N_28013,N_27385,N_27367);
nor U28014 (N_28014,N_27134,N_27429);
nand U28015 (N_28015,N_27324,N_27539);
nand U28016 (N_28016,N_27245,N_27435);
and U28017 (N_28017,N_27582,N_27390);
and U28018 (N_28018,N_27402,N_27356);
nand U28019 (N_28019,N_27395,N_27371);
nor U28020 (N_28020,N_27552,N_27228);
nor U28021 (N_28021,N_27309,N_27164);
nor U28022 (N_28022,N_27079,N_27534);
nand U28023 (N_28023,N_27411,N_27453);
xor U28024 (N_28024,N_27462,N_27192);
nor U28025 (N_28025,N_27128,N_27044);
xor U28026 (N_28026,N_27136,N_27175);
or U28027 (N_28027,N_27338,N_27388);
and U28028 (N_28028,N_27576,N_27396);
nor U28029 (N_28029,N_27569,N_27164);
nor U28030 (N_28030,N_27007,N_27547);
and U28031 (N_28031,N_27478,N_27534);
nor U28032 (N_28032,N_27091,N_27307);
nand U28033 (N_28033,N_27370,N_27378);
nor U28034 (N_28034,N_27352,N_27325);
nor U28035 (N_28035,N_27099,N_27005);
and U28036 (N_28036,N_27354,N_27324);
and U28037 (N_28037,N_27514,N_27490);
xor U28038 (N_28038,N_27440,N_27585);
and U28039 (N_28039,N_27314,N_27178);
or U28040 (N_28040,N_27139,N_27001);
nor U28041 (N_28041,N_27363,N_27388);
and U28042 (N_28042,N_27557,N_27080);
nand U28043 (N_28043,N_27586,N_27061);
or U28044 (N_28044,N_27034,N_27164);
nor U28045 (N_28045,N_27470,N_27065);
nor U28046 (N_28046,N_27550,N_27272);
nor U28047 (N_28047,N_27226,N_27102);
nand U28048 (N_28048,N_27107,N_27058);
nor U28049 (N_28049,N_27572,N_27268);
or U28050 (N_28050,N_27306,N_27135);
xor U28051 (N_28051,N_27179,N_27584);
nand U28052 (N_28052,N_27137,N_27352);
nor U28053 (N_28053,N_27407,N_27054);
and U28054 (N_28054,N_27250,N_27587);
or U28055 (N_28055,N_27189,N_27229);
xor U28056 (N_28056,N_27225,N_27255);
nand U28057 (N_28057,N_27188,N_27540);
nor U28058 (N_28058,N_27548,N_27034);
nor U28059 (N_28059,N_27310,N_27053);
and U28060 (N_28060,N_27248,N_27068);
or U28061 (N_28061,N_27377,N_27310);
nor U28062 (N_28062,N_27353,N_27503);
nor U28063 (N_28063,N_27058,N_27385);
nor U28064 (N_28064,N_27078,N_27238);
or U28065 (N_28065,N_27205,N_27177);
and U28066 (N_28066,N_27512,N_27472);
nand U28067 (N_28067,N_27073,N_27196);
nor U28068 (N_28068,N_27343,N_27182);
or U28069 (N_28069,N_27206,N_27033);
nor U28070 (N_28070,N_27434,N_27077);
or U28071 (N_28071,N_27467,N_27248);
and U28072 (N_28072,N_27304,N_27079);
nor U28073 (N_28073,N_27047,N_27266);
xnor U28074 (N_28074,N_27581,N_27458);
nand U28075 (N_28075,N_27211,N_27085);
xnor U28076 (N_28076,N_27118,N_27453);
and U28077 (N_28077,N_27541,N_27330);
nor U28078 (N_28078,N_27200,N_27573);
and U28079 (N_28079,N_27251,N_27028);
xor U28080 (N_28080,N_27261,N_27541);
nor U28081 (N_28081,N_27461,N_27096);
nand U28082 (N_28082,N_27255,N_27582);
nand U28083 (N_28083,N_27388,N_27021);
nand U28084 (N_28084,N_27242,N_27002);
or U28085 (N_28085,N_27088,N_27422);
or U28086 (N_28086,N_27174,N_27239);
and U28087 (N_28087,N_27236,N_27493);
and U28088 (N_28088,N_27083,N_27415);
nor U28089 (N_28089,N_27273,N_27115);
or U28090 (N_28090,N_27520,N_27416);
nor U28091 (N_28091,N_27115,N_27537);
or U28092 (N_28092,N_27467,N_27414);
nor U28093 (N_28093,N_27414,N_27493);
or U28094 (N_28094,N_27515,N_27402);
nand U28095 (N_28095,N_27384,N_27177);
nand U28096 (N_28096,N_27581,N_27289);
and U28097 (N_28097,N_27140,N_27252);
nand U28098 (N_28098,N_27565,N_27480);
nand U28099 (N_28099,N_27543,N_27140);
nand U28100 (N_28100,N_27338,N_27385);
xnor U28101 (N_28101,N_27395,N_27194);
nor U28102 (N_28102,N_27454,N_27428);
and U28103 (N_28103,N_27399,N_27020);
or U28104 (N_28104,N_27506,N_27237);
xnor U28105 (N_28105,N_27084,N_27334);
nand U28106 (N_28106,N_27184,N_27114);
nor U28107 (N_28107,N_27227,N_27465);
nor U28108 (N_28108,N_27590,N_27473);
and U28109 (N_28109,N_27452,N_27333);
nand U28110 (N_28110,N_27239,N_27238);
and U28111 (N_28111,N_27550,N_27453);
nand U28112 (N_28112,N_27215,N_27442);
nand U28113 (N_28113,N_27109,N_27096);
nor U28114 (N_28114,N_27576,N_27230);
nand U28115 (N_28115,N_27157,N_27005);
nor U28116 (N_28116,N_27455,N_27341);
nand U28117 (N_28117,N_27243,N_27004);
and U28118 (N_28118,N_27353,N_27462);
nand U28119 (N_28119,N_27514,N_27191);
and U28120 (N_28120,N_27193,N_27081);
nand U28121 (N_28121,N_27587,N_27160);
and U28122 (N_28122,N_27567,N_27418);
and U28123 (N_28123,N_27309,N_27392);
and U28124 (N_28124,N_27099,N_27306);
nor U28125 (N_28125,N_27353,N_27423);
nor U28126 (N_28126,N_27047,N_27040);
nand U28127 (N_28127,N_27208,N_27012);
nand U28128 (N_28128,N_27484,N_27357);
nor U28129 (N_28129,N_27243,N_27312);
and U28130 (N_28130,N_27170,N_27162);
nor U28131 (N_28131,N_27455,N_27082);
nand U28132 (N_28132,N_27490,N_27380);
or U28133 (N_28133,N_27554,N_27158);
nand U28134 (N_28134,N_27223,N_27189);
and U28135 (N_28135,N_27166,N_27399);
nor U28136 (N_28136,N_27311,N_27459);
nand U28137 (N_28137,N_27513,N_27019);
or U28138 (N_28138,N_27353,N_27311);
or U28139 (N_28139,N_27397,N_27525);
nand U28140 (N_28140,N_27096,N_27566);
nor U28141 (N_28141,N_27407,N_27329);
and U28142 (N_28142,N_27426,N_27272);
nor U28143 (N_28143,N_27533,N_27515);
nor U28144 (N_28144,N_27331,N_27194);
nor U28145 (N_28145,N_27516,N_27275);
nand U28146 (N_28146,N_27224,N_27091);
nor U28147 (N_28147,N_27342,N_27410);
nor U28148 (N_28148,N_27514,N_27169);
nor U28149 (N_28149,N_27364,N_27538);
and U28150 (N_28150,N_27063,N_27211);
and U28151 (N_28151,N_27528,N_27464);
nor U28152 (N_28152,N_27069,N_27456);
nand U28153 (N_28153,N_27250,N_27109);
or U28154 (N_28154,N_27147,N_27563);
and U28155 (N_28155,N_27457,N_27400);
and U28156 (N_28156,N_27516,N_27105);
and U28157 (N_28157,N_27226,N_27498);
and U28158 (N_28158,N_27250,N_27582);
and U28159 (N_28159,N_27017,N_27350);
or U28160 (N_28160,N_27145,N_27152);
nor U28161 (N_28161,N_27010,N_27129);
or U28162 (N_28162,N_27504,N_27379);
xnor U28163 (N_28163,N_27572,N_27226);
nand U28164 (N_28164,N_27516,N_27522);
nand U28165 (N_28165,N_27060,N_27296);
nand U28166 (N_28166,N_27329,N_27057);
nand U28167 (N_28167,N_27081,N_27191);
nand U28168 (N_28168,N_27104,N_27302);
nand U28169 (N_28169,N_27441,N_27036);
nor U28170 (N_28170,N_27433,N_27220);
and U28171 (N_28171,N_27546,N_27336);
or U28172 (N_28172,N_27509,N_27517);
and U28173 (N_28173,N_27557,N_27272);
nor U28174 (N_28174,N_27306,N_27448);
and U28175 (N_28175,N_27023,N_27340);
or U28176 (N_28176,N_27054,N_27526);
nor U28177 (N_28177,N_27338,N_27286);
nor U28178 (N_28178,N_27034,N_27485);
nand U28179 (N_28179,N_27265,N_27279);
and U28180 (N_28180,N_27451,N_27117);
or U28181 (N_28181,N_27574,N_27596);
nor U28182 (N_28182,N_27144,N_27340);
nand U28183 (N_28183,N_27018,N_27190);
nor U28184 (N_28184,N_27385,N_27562);
nor U28185 (N_28185,N_27368,N_27388);
nor U28186 (N_28186,N_27093,N_27035);
nor U28187 (N_28187,N_27385,N_27509);
or U28188 (N_28188,N_27098,N_27225);
or U28189 (N_28189,N_27262,N_27300);
nand U28190 (N_28190,N_27446,N_27225);
nand U28191 (N_28191,N_27273,N_27509);
nor U28192 (N_28192,N_27340,N_27009);
nand U28193 (N_28193,N_27244,N_27324);
and U28194 (N_28194,N_27552,N_27134);
and U28195 (N_28195,N_27047,N_27537);
nand U28196 (N_28196,N_27115,N_27511);
and U28197 (N_28197,N_27188,N_27216);
nand U28198 (N_28198,N_27543,N_27209);
and U28199 (N_28199,N_27279,N_27197);
and U28200 (N_28200,N_27671,N_28016);
nand U28201 (N_28201,N_28114,N_27680);
and U28202 (N_28202,N_28179,N_27732);
nand U28203 (N_28203,N_28031,N_27602);
nor U28204 (N_28204,N_28046,N_27990);
nor U28205 (N_28205,N_27682,N_28049);
nor U28206 (N_28206,N_27679,N_28177);
nand U28207 (N_28207,N_28175,N_27704);
nand U28208 (N_28208,N_27721,N_27821);
and U28209 (N_28209,N_27952,N_28026);
nor U28210 (N_28210,N_27639,N_28022);
xnor U28211 (N_28211,N_27713,N_28020);
nand U28212 (N_28212,N_27810,N_27861);
and U28213 (N_28213,N_27710,N_28190);
nand U28214 (N_28214,N_28089,N_27853);
nor U28215 (N_28215,N_28075,N_27651);
and U28216 (N_28216,N_28134,N_27731);
or U28217 (N_28217,N_28129,N_27927);
and U28218 (N_28218,N_27768,N_28132);
nand U28219 (N_28219,N_27871,N_28101);
and U28220 (N_28220,N_28193,N_28181);
and U28221 (N_28221,N_27984,N_27706);
nand U28222 (N_28222,N_28055,N_27995);
nand U28223 (N_28223,N_28117,N_27972);
nor U28224 (N_28224,N_27686,N_28113);
nand U28225 (N_28225,N_28010,N_27833);
nor U28226 (N_28226,N_27856,N_27695);
nor U28227 (N_28227,N_28041,N_28009);
and U28228 (N_28228,N_28173,N_28081);
and U28229 (N_28229,N_27608,N_27741);
nand U28230 (N_28230,N_27794,N_28038);
nand U28231 (N_28231,N_27940,N_27791);
nand U28232 (N_28232,N_28032,N_27830);
nor U28233 (N_28233,N_27998,N_27719);
nand U28234 (N_28234,N_28195,N_27699);
nor U28235 (N_28235,N_27735,N_28112);
nand U28236 (N_28236,N_27837,N_27975);
nor U28237 (N_28237,N_27987,N_28052);
nor U28238 (N_28238,N_28199,N_27626);
or U28239 (N_28239,N_28054,N_27764);
nor U28240 (N_28240,N_27920,N_27784);
nand U28241 (N_28241,N_27907,N_28168);
or U28242 (N_28242,N_28150,N_27829);
nor U28243 (N_28243,N_28119,N_27778);
nor U28244 (N_28244,N_28005,N_28169);
nand U28245 (N_28245,N_28084,N_28111);
or U28246 (N_28246,N_28043,N_28183);
nand U28247 (N_28247,N_27634,N_28118);
and U28248 (N_28248,N_27900,N_27958);
or U28249 (N_28249,N_28057,N_27879);
nand U28250 (N_28250,N_27649,N_28069);
nand U28251 (N_28251,N_27672,N_27961);
and U28252 (N_28252,N_28108,N_28187);
xnor U28253 (N_28253,N_27766,N_27727);
and U28254 (N_28254,N_28036,N_27960);
and U28255 (N_28255,N_27733,N_27926);
or U28256 (N_28256,N_27911,N_28191);
and U28257 (N_28257,N_27687,N_27755);
and U28258 (N_28258,N_27798,N_28065);
xor U28259 (N_28259,N_27740,N_28125);
or U28260 (N_28260,N_27802,N_27955);
nand U28261 (N_28261,N_27666,N_28166);
or U28262 (N_28262,N_27771,N_27773);
nand U28263 (N_28263,N_27908,N_27715);
or U28264 (N_28264,N_27889,N_28088);
nand U28265 (N_28265,N_27916,N_28085);
or U28266 (N_28266,N_27752,N_27973);
nor U28267 (N_28267,N_27854,N_27992);
xnor U28268 (N_28268,N_28066,N_27658);
or U28269 (N_28269,N_27693,N_27838);
xnor U28270 (N_28270,N_27997,N_27858);
and U28271 (N_28271,N_27865,N_27758);
or U28272 (N_28272,N_28139,N_27867);
nor U28273 (N_28273,N_27925,N_27759);
nor U28274 (N_28274,N_28171,N_27882);
nand U28275 (N_28275,N_27722,N_27909);
or U28276 (N_28276,N_27941,N_27915);
nor U28277 (N_28277,N_27754,N_27690);
xnor U28278 (N_28278,N_27665,N_27795);
or U28279 (N_28279,N_27967,N_28015);
nand U28280 (N_28280,N_27994,N_27923);
nand U28281 (N_28281,N_27825,N_27828);
or U28282 (N_28282,N_27612,N_27816);
and U28283 (N_28283,N_27930,N_28017);
nand U28284 (N_28284,N_27776,N_27709);
nor U28285 (N_28285,N_28174,N_27790);
or U28286 (N_28286,N_27603,N_27880);
nand U28287 (N_28287,N_27783,N_28182);
or U28288 (N_28288,N_27921,N_27876);
nand U28289 (N_28289,N_28006,N_27656);
and U28290 (N_28290,N_27760,N_27931);
nor U28291 (N_28291,N_28033,N_27614);
nor U28292 (N_28292,N_27866,N_27953);
or U28293 (N_28293,N_28144,N_27730);
or U28294 (N_28294,N_28160,N_27806);
nand U28295 (N_28295,N_27697,N_28023);
nor U28296 (N_28296,N_27692,N_27942);
nand U28297 (N_28297,N_28120,N_27939);
nor U28298 (N_28298,N_27847,N_27616);
and U28299 (N_28299,N_28067,N_27933);
xnor U28300 (N_28300,N_27922,N_28186);
or U28301 (N_28301,N_28061,N_27738);
nand U28302 (N_28302,N_27849,N_28180);
or U28303 (N_28303,N_27875,N_27604);
xor U28304 (N_28304,N_27750,N_27996);
nor U28305 (N_28305,N_27674,N_28126);
and U28306 (N_28306,N_27796,N_28109);
or U28307 (N_28307,N_28077,N_27747);
nand U28308 (N_28308,N_28058,N_28124);
nor U28309 (N_28309,N_27834,N_28042);
and U28310 (N_28310,N_28063,N_28189);
and U28311 (N_28311,N_27648,N_27895);
nor U28312 (N_28312,N_27630,N_27729);
or U28313 (N_28313,N_27696,N_27976);
xor U28314 (N_28314,N_28176,N_28086);
nand U28315 (N_28315,N_27919,N_27661);
nand U28316 (N_28316,N_27846,N_28121);
nor U28317 (N_28317,N_27891,N_27711);
or U28318 (N_28318,N_27888,N_27652);
and U28319 (N_28319,N_27950,N_28098);
and U28320 (N_28320,N_28140,N_28045);
or U28321 (N_28321,N_27971,N_28192);
nand U28322 (N_28322,N_27873,N_27818);
and U28323 (N_28323,N_27782,N_27887);
xor U28324 (N_28324,N_28198,N_28037);
and U28325 (N_28325,N_28083,N_27800);
or U28326 (N_28326,N_28153,N_28155);
or U28327 (N_28327,N_28133,N_27769);
nor U28328 (N_28328,N_28094,N_27787);
and U28329 (N_28329,N_28048,N_27650);
or U28330 (N_28330,N_27848,N_28165);
and U28331 (N_28331,N_27788,N_28019);
nand U28332 (N_28332,N_27611,N_27897);
nor U28333 (N_28333,N_27884,N_28154);
and U28334 (N_28334,N_27844,N_27663);
nor U28335 (N_28335,N_27670,N_27748);
nand U28336 (N_28336,N_27845,N_28012);
nand U28337 (N_28337,N_28095,N_27749);
or U28338 (N_28338,N_28188,N_27803);
and U28339 (N_28339,N_28172,N_27765);
or U28340 (N_28340,N_27944,N_27969);
or U28341 (N_28341,N_28135,N_28073);
and U28342 (N_28342,N_28029,N_28137);
xnor U28343 (N_28343,N_27691,N_27780);
or U28344 (N_28344,N_27763,N_27945);
nor U28345 (N_28345,N_27831,N_27965);
nand U28346 (N_28346,N_27762,N_27645);
nor U28347 (N_28347,N_28024,N_28011);
nand U28348 (N_28348,N_27653,N_27947);
nor U28349 (N_28349,N_28167,N_27757);
nand U28350 (N_28350,N_27986,N_28184);
and U28351 (N_28351,N_27899,N_27989);
or U28352 (N_28352,N_27705,N_27607);
nor U28353 (N_28353,N_27797,N_28161);
or U28354 (N_28354,N_27872,N_28136);
and U28355 (N_28355,N_27936,N_27684);
or U28356 (N_28356,N_28156,N_27781);
nand U28357 (N_28357,N_28064,N_27823);
and U28358 (N_28358,N_27896,N_28130);
nand U28359 (N_28359,N_27770,N_28151);
nor U28360 (N_28360,N_27644,N_27761);
or U28361 (N_28361,N_27647,N_27643);
nor U28362 (N_28362,N_28116,N_27929);
xnor U28363 (N_28363,N_27843,N_27617);
and U28364 (N_28364,N_28002,N_28142);
nand U28365 (N_28365,N_28128,N_27917);
and U28366 (N_28366,N_28122,N_27662);
nor U28367 (N_28367,N_28178,N_28141);
nand U28368 (N_28368,N_27792,N_27898);
or U28369 (N_28369,N_28008,N_27901);
nand U28370 (N_28370,N_27894,N_27957);
nor U28371 (N_28371,N_28027,N_28090);
nor U28372 (N_28372,N_28013,N_27779);
nand U28373 (N_28373,N_27734,N_27840);
xor U28374 (N_28374,N_28001,N_27869);
nand U28375 (N_28375,N_28163,N_27775);
nor U28376 (N_28376,N_27777,N_27789);
nor U28377 (N_28377,N_28053,N_27689);
and U28378 (N_28378,N_27655,N_27677);
or U28379 (N_28379,N_28072,N_27724);
or U28380 (N_28380,N_27736,N_27683);
nor U28381 (N_28381,N_27799,N_28115);
nor U28382 (N_28382,N_27673,N_27903);
and U28383 (N_28383,N_27659,N_28197);
nor U28384 (N_28384,N_27842,N_28143);
nand U28385 (N_28385,N_28105,N_27725);
or U28386 (N_28386,N_28068,N_27720);
or U28387 (N_28387,N_28025,N_27906);
and U28388 (N_28388,N_28076,N_28018);
nand U28389 (N_28389,N_27913,N_28030);
and U28390 (N_28390,N_27943,N_27954);
and U28391 (N_28391,N_27714,N_27669);
nor U28392 (N_28392,N_28104,N_28159);
nor U28393 (N_28393,N_27610,N_28096);
or U28394 (N_28394,N_28091,N_27746);
nand U28395 (N_28395,N_28003,N_27707);
nand U28396 (N_28396,N_27751,N_28050);
nand U28397 (N_28397,N_28147,N_27708);
nand U28398 (N_28398,N_27977,N_27902);
or U28399 (N_28399,N_27657,N_27868);
nor U28400 (N_28400,N_27811,N_28035);
and U28401 (N_28401,N_28127,N_27624);
and U28402 (N_28402,N_28071,N_27964);
nor U28403 (N_28403,N_27855,N_27852);
or U28404 (N_28404,N_27959,N_28152);
and U28405 (N_28405,N_27716,N_27621);
or U28406 (N_28406,N_28007,N_28051);
nor U28407 (N_28407,N_28102,N_27668);
and U28408 (N_28408,N_27827,N_27970);
or U28409 (N_28409,N_28107,N_28044);
or U28410 (N_28410,N_27619,N_27813);
nand U28411 (N_28411,N_27678,N_27851);
nor U28412 (N_28412,N_27822,N_27982);
and U28413 (N_28413,N_27703,N_27966);
and U28414 (N_28414,N_27999,N_28146);
nand U28415 (N_28415,N_28060,N_27937);
and U28416 (N_28416,N_28062,N_27814);
nor U28417 (N_28417,N_27786,N_27935);
and U28418 (N_28418,N_27820,N_28110);
and U28419 (N_28419,N_27974,N_28097);
nand U28420 (N_28420,N_28170,N_27932);
nor U28421 (N_28421,N_28158,N_27642);
nor U28422 (N_28422,N_27817,N_28034);
or U28423 (N_28423,N_27863,N_27744);
nor U28424 (N_28424,N_27743,N_27637);
nand U28425 (N_28425,N_27910,N_27737);
or U28426 (N_28426,N_28123,N_27946);
and U28427 (N_28427,N_27874,N_27885);
and U28428 (N_28428,N_27615,N_27963);
nor U28429 (N_28429,N_28131,N_27841);
and U28430 (N_28430,N_27685,N_28040);
nand U28431 (N_28431,N_27613,N_27681);
nor U28432 (N_28432,N_27633,N_28196);
and U28433 (N_28433,N_27819,N_27636);
nand U28434 (N_28434,N_28099,N_27812);
or U28435 (N_28435,N_27983,N_28082);
nand U28436 (N_28436,N_27606,N_27904);
and U28437 (N_28437,N_27857,N_28059);
nor U28438 (N_28438,N_28194,N_27890);
nor U28439 (N_28439,N_27980,N_28185);
nor U28440 (N_28440,N_27801,N_27859);
and U28441 (N_28441,N_27622,N_28148);
and U28442 (N_28442,N_27667,N_28070);
and U28443 (N_28443,N_27839,N_28078);
or U28444 (N_28444,N_27832,N_27864);
or U28445 (N_28445,N_27892,N_27698);
and U28446 (N_28446,N_27739,N_28021);
and U28447 (N_28447,N_27914,N_27815);
and U28448 (N_28448,N_28162,N_27883);
and U28449 (N_28449,N_27993,N_27676);
and U28450 (N_28450,N_28100,N_27793);
or U28451 (N_28451,N_27878,N_28103);
and U28452 (N_28452,N_28149,N_27951);
nor U28453 (N_28453,N_27893,N_27905);
or U28454 (N_28454,N_28164,N_27772);
or U28455 (N_28455,N_27981,N_27717);
and U28456 (N_28456,N_27767,N_28106);
nor U28457 (N_28457,N_27654,N_27675);
or U28458 (N_28458,N_28092,N_27988);
and U28459 (N_28459,N_28028,N_27948);
nand U28460 (N_28460,N_27627,N_27701);
and U28461 (N_28461,N_28014,N_27640);
nand U28462 (N_28462,N_27809,N_27753);
or U28463 (N_28463,N_27886,N_27660);
nor U28464 (N_28464,N_27646,N_27805);
nand U28465 (N_28465,N_27718,N_28093);
or U28466 (N_28466,N_27712,N_27912);
and U28467 (N_28467,N_27862,N_27991);
and U28468 (N_28468,N_27609,N_27928);
nand U28469 (N_28469,N_27807,N_28080);
and U28470 (N_28470,N_27601,N_27620);
nor U28471 (N_28471,N_27638,N_28056);
nand U28472 (N_28472,N_27625,N_27835);
nand U28473 (N_28473,N_27949,N_27978);
or U28474 (N_28474,N_27618,N_27785);
nand U28475 (N_28475,N_27881,N_28145);
nor U28476 (N_28476,N_27702,N_28087);
nor U28477 (N_28477,N_27924,N_27600);
nand U28478 (N_28478,N_27635,N_27934);
and U28479 (N_28479,N_28039,N_28157);
nor U28480 (N_28480,N_27623,N_27756);
nand U28481 (N_28481,N_27826,N_27938);
or U28482 (N_28482,N_27968,N_28138);
nand U28483 (N_28483,N_27742,N_28074);
nand U28484 (N_28484,N_27700,N_27664);
nand U28485 (N_28485,N_27956,N_28047);
nor U28486 (N_28486,N_27774,N_27918);
nor U28487 (N_28487,N_27962,N_27985);
and U28488 (N_28488,N_27726,N_27728);
nand U28489 (N_28489,N_28004,N_28000);
xnor U28490 (N_28490,N_27629,N_27745);
or U28491 (N_28491,N_27694,N_27688);
and U28492 (N_28492,N_27641,N_27877);
and U28493 (N_28493,N_27824,N_27723);
and U28494 (N_28494,N_27850,N_27860);
nor U28495 (N_28495,N_27808,N_27804);
nand U28496 (N_28496,N_27605,N_27628);
nand U28497 (N_28497,N_27632,N_27870);
and U28498 (N_28498,N_27979,N_27836);
xnor U28499 (N_28499,N_28079,N_27631);
nand U28500 (N_28500,N_27677,N_27814);
and U28501 (N_28501,N_27949,N_27624);
nand U28502 (N_28502,N_27711,N_27899);
nor U28503 (N_28503,N_27758,N_28169);
nand U28504 (N_28504,N_28166,N_27694);
or U28505 (N_28505,N_27966,N_27649);
nor U28506 (N_28506,N_27854,N_27985);
nand U28507 (N_28507,N_28124,N_27806);
and U28508 (N_28508,N_27930,N_27602);
nor U28509 (N_28509,N_27940,N_27967);
and U28510 (N_28510,N_27666,N_28133);
and U28511 (N_28511,N_27927,N_27996);
and U28512 (N_28512,N_28003,N_27914);
or U28513 (N_28513,N_27635,N_27627);
nand U28514 (N_28514,N_27627,N_27922);
nand U28515 (N_28515,N_27860,N_27748);
nor U28516 (N_28516,N_27995,N_27901);
and U28517 (N_28517,N_27921,N_27662);
and U28518 (N_28518,N_27850,N_27986);
or U28519 (N_28519,N_28124,N_28116);
or U28520 (N_28520,N_27809,N_27813);
and U28521 (N_28521,N_28096,N_27782);
or U28522 (N_28522,N_27765,N_27772);
nor U28523 (N_28523,N_27706,N_28029);
or U28524 (N_28524,N_27829,N_28032);
or U28525 (N_28525,N_27783,N_27942);
or U28526 (N_28526,N_27729,N_27865);
nor U28527 (N_28527,N_28088,N_27833);
and U28528 (N_28528,N_27675,N_28121);
nor U28529 (N_28529,N_27818,N_27741);
and U28530 (N_28530,N_27975,N_27672);
and U28531 (N_28531,N_27677,N_28187);
nor U28532 (N_28532,N_27891,N_27861);
nor U28533 (N_28533,N_27960,N_27997);
and U28534 (N_28534,N_27867,N_27659);
or U28535 (N_28535,N_28148,N_27969);
and U28536 (N_28536,N_28167,N_27965);
or U28537 (N_28537,N_27726,N_27886);
nand U28538 (N_28538,N_28155,N_27900);
nand U28539 (N_28539,N_27654,N_27632);
nand U28540 (N_28540,N_27806,N_27628);
nor U28541 (N_28541,N_28099,N_28106);
and U28542 (N_28542,N_27753,N_27723);
and U28543 (N_28543,N_27728,N_27916);
nor U28544 (N_28544,N_27809,N_27940);
nor U28545 (N_28545,N_27743,N_27744);
nand U28546 (N_28546,N_27799,N_27825);
or U28547 (N_28547,N_27817,N_27985);
or U28548 (N_28548,N_28154,N_27858);
xnor U28549 (N_28549,N_27748,N_28117);
and U28550 (N_28550,N_27698,N_27865);
and U28551 (N_28551,N_27691,N_27882);
or U28552 (N_28552,N_27727,N_28062);
or U28553 (N_28553,N_28160,N_28095);
nor U28554 (N_28554,N_28061,N_27861);
nor U28555 (N_28555,N_28040,N_27977);
or U28556 (N_28556,N_27656,N_28098);
nor U28557 (N_28557,N_27622,N_27869);
nand U28558 (N_28558,N_27610,N_27735);
nor U28559 (N_28559,N_28170,N_27966);
nor U28560 (N_28560,N_27701,N_27799);
or U28561 (N_28561,N_27957,N_27908);
and U28562 (N_28562,N_27649,N_28129);
nor U28563 (N_28563,N_28010,N_27954);
xor U28564 (N_28564,N_28198,N_27812);
and U28565 (N_28565,N_27913,N_27615);
and U28566 (N_28566,N_27940,N_27948);
nand U28567 (N_28567,N_28137,N_27684);
and U28568 (N_28568,N_28190,N_27808);
or U28569 (N_28569,N_27793,N_27795);
nor U28570 (N_28570,N_28178,N_27986);
or U28571 (N_28571,N_27650,N_27809);
or U28572 (N_28572,N_28066,N_27772);
nor U28573 (N_28573,N_27659,N_27698);
nor U28574 (N_28574,N_28074,N_27837);
and U28575 (N_28575,N_28149,N_27604);
or U28576 (N_28576,N_27741,N_28064);
nor U28577 (N_28577,N_27673,N_28115);
or U28578 (N_28578,N_27628,N_27894);
nor U28579 (N_28579,N_28031,N_27970);
or U28580 (N_28580,N_27721,N_27843);
and U28581 (N_28581,N_27638,N_27713);
and U28582 (N_28582,N_27806,N_28184);
nand U28583 (N_28583,N_27964,N_27820);
nand U28584 (N_28584,N_28111,N_28026);
or U28585 (N_28585,N_27675,N_28133);
nand U28586 (N_28586,N_27678,N_27944);
nor U28587 (N_28587,N_27754,N_27881);
or U28588 (N_28588,N_27613,N_27869);
and U28589 (N_28589,N_27818,N_28128);
or U28590 (N_28590,N_28075,N_28154);
or U28591 (N_28591,N_28094,N_28005);
or U28592 (N_28592,N_27714,N_28145);
nand U28593 (N_28593,N_27647,N_27985);
and U28594 (N_28594,N_28013,N_27825);
and U28595 (N_28595,N_27913,N_27663);
or U28596 (N_28596,N_28182,N_27823);
nand U28597 (N_28597,N_27816,N_27844);
nand U28598 (N_28598,N_27768,N_27652);
and U28599 (N_28599,N_27794,N_28020);
nand U28600 (N_28600,N_27676,N_27995);
nor U28601 (N_28601,N_27837,N_28138);
and U28602 (N_28602,N_28036,N_27901);
xnor U28603 (N_28603,N_27651,N_27950);
nor U28604 (N_28604,N_28051,N_27698);
and U28605 (N_28605,N_27691,N_28087);
or U28606 (N_28606,N_27798,N_27771);
nand U28607 (N_28607,N_27978,N_27823);
nand U28608 (N_28608,N_27845,N_27927);
nor U28609 (N_28609,N_27862,N_27966);
or U28610 (N_28610,N_28045,N_27819);
and U28611 (N_28611,N_27716,N_28166);
nor U28612 (N_28612,N_28080,N_28098);
or U28613 (N_28613,N_27772,N_27888);
or U28614 (N_28614,N_27616,N_27647);
nand U28615 (N_28615,N_28194,N_28149);
nand U28616 (N_28616,N_27885,N_27689);
or U28617 (N_28617,N_27920,N_27808);
nor U28618 (N_28618,N_27832,N_27610);
or U28619 (N_28619,N_28072,N_28119);
xnor U28620 (N_28620,N_27980,N_27821);
and U28621 (N_28621,N_27751,N_27939);
nor U28622 (N_28622,N_27692,N_27630);
nor U28623 (N_28623,N_28186,N_27667);
nand U28624 (N_28624,N_28125,N_27912);
nand U28625 (N_28625,N_27759,N_27812);
nand U28626 (N_28626,N_27969,N_28046);
or U28627 (N_28627,N_28119,N_27737);
xnor U28628 (N_28628,N_28057,N_27954);
xor U28629 (N_28629,N_28181,N_27860);
nor U28630 (N_28630,N_27909,N_27896);
nor U28631 (N_28631,N_27878,N_27791);
or U28632 (N_28632,N_28122,N_27738);
or U28633 (N_28633,N_27994,N_27908);
and U28634 (N_28634,N_27648,N_27987);
nand U28635 (N_28635,N_27622,N_27842);
and U28636 (N_28636,N_27678,N_27992);
xnor U28637 (N_28637,N_27889,N_27673);
nand U28638 (N_28638,N_28118,N_27826);
and U28639 (N_28639,N_28199,N_27870);
and U28640 (N_28640,N_27910,N_27854);
nor U28641 (N_28641,N_28154,N_28053);
nor U28642 (N_28642,N_27614,N_27916);
or U28643 (N_28643,N_27919,N_27926);
nand U28644 (N_28644,N_28015,N_28047);
nor U28645 (N_28645,N_28012,N_27945);
and U28646 (N_28646,N_27677,N_27619);
and U28647 (N_28647,N_28023,N_28075);
nand U28648 (N_28648,N_27984,N_28024);
and U28649 (N_28649,N_27693,N_27746);
or U28650 (N_28650,N_27823,N_27675);
xor U28651 (N_28651,N_27609,N_28117);
xnor U28652 (N_28652,N_27744,N_27824);
nor U28653 (N_28653,N_27938,N_27939);
and U28654 (N_28654,N_27803,N_27843);
or U28655 (N_28655,N_28069,N_27950);
nand U28656 (N_28656,N_28148,N_27767);
nor U28657 (N_28657,N_27868,N_28150);
nor U28658 (N_28658,N_27870,N_28066);
xor U28659 (N_28659,N_28123,N_28043);
nor U28660 (N_28660,N_27884,N_27839);
or U28661 (N_28661,N_27666,N_28112);
nand U28662 (N_28662,N_28166,N_27663);
nor U28663 (N_28663,N_27633,N_27968);
nand U28664 (N_28664,N_27983,N_27647);
xor U28665 (N_28665,N_27658,N_28137);
xor U28666 (N_28666,N_28155,N_27918);
nand U28667 (N_28667,N_28070,N_27884);
and U28668 (N_28668,N_28001,N_28038);
or U28669 (N_28669,N_27751,N_27744);
nor U28670 (N_28670,N_27994,N_27703);
and U28671 (N_28671,N_27946,N_27955);
and U28672 (N_28672,N_28010,N_28002);
nor U28673 (N_28673,N_27821,N_28184);
or U28674 (N_28674,N_27746,N_27836);
nand U28675 (N_28675,N_27965,N_27791);
and U28676 (N_28676,N_27714,N_27833);
nor U28677 (N_28677,N_28026,N_28172);
and U28678 (N_28678,N_28072,N_27906);
nand U28679 (N_28679,N_27752,N_27735);
nor U28680 (N_28680,N_28041,N_27639);
or U28681 (N_28681,N_27899,N_28020);
nand U28682 (N_28682,N_28128,N_27991);
or U28683 (N_28683,N_27808,N_27759);
or U28684 (N_28684,N_27855,N_28093);
nand U28685 (N_28685,N_27946,N_27926);
nand U28686 (N_28686,N_27801,N_28031);
nor U28687 (N_28687,N_28174,N_27733);
and U28688 (N_28688,N_28124,N_27752);
and U28689 (N_28689,N_27879,N_27927);
or U28690 (N_28690,N_28036,N_27985);
and U28691 (N_28691,N_27840,N_27890);
and U28692 (N_28692,N_27830,N_28159);
and U28693 (N_28693,N_28018,N_27655);
nand U28694 (N_28694,N_27924,N_27751);
and U28695 (N_28695,N_27925,N_28041);
nand U28696 (N_28696,N_27914,N_28079);
nor U28697 (N_28697,N_28120,N_27759);
or U28698 (N_28698,N_28013,N_28194);
nand U28699 (N_28699,N_27971,N_27675);
or U28700 (N_28700,N_27769,N_27956);
and U28701 (N_28701,N_27966,N_28063);
nor U28702 (N_28702,N_27814,N_28044);
nand U28703 (N_28703,N_28130,N_27824);
or U28704 (N_28704,N_28065,N_27913);
or U28705 (N_28705,N_27812,N_27783);
nor U28706 (N_28706,N_27607,N_27746);
nand U28707 (N_28707,N_27887,N_27936);
and U28708 (N_28708,N_27873,N_27673);
nor U28709 (N_28709,N_28001,N_28184);
nand U28710 (N_28710,N_28185,N_27629);
and U28711 (N_28711,N_27806,N_27630);
or U28712 (N_28712,N_27670,N_27759);
xor U28713 (N_28713,N_27842,N_28044);
or U28714 (N_28714,N_28015,N_27990);
nor U28715 (N_28715,N_27967,N_28142);
nor U28716 (N_28716,N_27968,N_27870);
xor U28717 (N_28717,N_28195,N_28031);
nor U28718 (N_28718,N_28156,N_27808);
nor U28719 (N_28719,N_27856,N_27844);
nand U28720 (N_28720,N_27781,N_27779);
xor U28721 (N_28721,N_27933,N_27678);
or U28722 (N_28722,N_28075,N_28019);
nor U28723 (N_28723,N_27825,N_27759);
and U28724 (N_28724,N_28155,N_27922);
or U28725 (N_28725,N_28035,N_27799);
nor U28726 (N_28726,N_27857,N_28160);
nor U28727 (N_28727,N_28038,N_27949);
and U28728 (N_28728,N_27889,N_27978);
or U28729 (N_28729,N_28104,N_28101);
and U28730 (N_28730,N_27870,N_27961);
nand U28731 (N_28731,N_28039,N_28107);
nand U28732 (N_28732,N_27781,N_27726);
nand U28733 (N_28733,N_27647,N_27909);
xnor U28734 (N_28734,N_28190,N_27742);
and U28735 (N_28735,N_27842,N_27994);
nand U28736 (N_28736,N_28183,N_28113);
nor U28737 (N_28737,N_27789,N_27779);
and U28738 (N_28738,N_27806,N_28188);
or U28739 (N_28739,N_28171,N_28075);
and U28740 (N_28740,N_27620,N_27746);
nand U28741 (N_28741,N_28082,N_27634);
nand U28742 (N_28742,N_28154,N_27770);
or U28743 (N_28743,N_28030,N_27711);
nand U28744 (N_28744,N_27939,N_27819);
and U28745 (N_28745,N_28008,N_27690);
or U28746 (N_28746,N_27943,N_27732);
or U28747 (N_28747,N_27836,N_28080);
nand U28748 (N_28748,N_28173,N_27783);
or U28749 (N_28749,N_28185,N_28108);
xor U28750 (N_28750,N_27973,N_27714);
or U28751 (N_28751,N_27820,N_27749);
nor U28752 (N_28752,N_27911,N_28166);
and U28753 (N_28753,N_27915,N_27956);
nor U28754 (N_28754,N_28019,N_27672);
nor U28755 (N_28755,N_27754,N_27745);
and U28756 (N_28756,N_27848,N_27846);
nor U28757 (N_28757,N_27986,N_27637);
nand U28758 (N_28758,N_28155,N_27852);
or U28759 (N_28759,N_27803,N_27888);
and U28760 (N_28760,N_27947,N_28101);
nor U28761 (N_28761,N_28116,N_27664);
or U28762 (N_28762,N_27787,N_28088);
and U28763 (N_28763,N_27866,N_28174);
or U28764 (N_28764,N_28060,N_28107);
or U28765 (N_28765,N_28096,N_27838);
xor U28766 (N_28766,N_28125,N_27899);
nand U28767 (N_28767,N_27621,N_27802);
and U28768 (N_28768,N_27884,N_27791);
xnor U28769 (N_28769,N_27727,N_27904);
nor U28770 (N_28770,N_28059,N_27884);
nand U28771 (N_28771,N_27799,N_27657);
and U28772 (N_28772,N_27768,N_27913);
nor U28773 (N_28773,N_27685,N_28167);
or U28774 (N_28774,N_27992,N_27643);
and U28775 (N_28775,N_27940,N_28008);
nand U28776 (N_28776,N_27935,N_27902);
and U28777 (N_28777,N_27702,N_27715);
nand U28778 (N_28778,N_27660,N_28087);
nand U28779 (N_28779,N_27663,N_27948);
and U28780 (N_28780,N_27857,N_28062);
and U28781 (N_28781,N_27952,N_27737);
and U28782 (N_28782,N_27787,N_27636);
nand U28783 (N_28783,N_27710,N_27655);
or U28784 (N_28784,N_27874,N_28119);
nor U28785 (N_28785,N_27939,N_27946);
nor U28786 (N_28786,N_28108,N_28104);
or U28787 (N_28787,N_27613,N_27983);
nor U28788 (N_28788,N_28166,N_27881);
nand U28789 (N_28789,N_27922,N_27618);
nor U28790 (N_28790,N_27831,N_28186);
nor U28791 (N_28791,N_28002,N_27656);
and U28792 (N_28792,N_27861,N_27812);
and U28793 (N_28793,N_27638,N_27667);
nand U28794 (N_28794,N_27966,N_28033);
and U28795 (N_28795,N_27707,N_28054);
or U28796 (N_28796,N_27644,N_27823);
nor U28797 (N_28797,N_28026,N_27733);
nand U28798 (N_28798,N_27754,N_27917);
or U28799 (N_28799,N_27865,N_27792);
or U28800 (N_28800,N_28376,N_28403);
nor U28801 (N_28801,N_28664,N_28387);
or U28802 (N_28802,N_28570,N_28404);
and U28803 (N_28803,N_28660,N_28600);
nand U28804 (N_28804,N_28236,N_28458);
and U28805 (N_28805,N_28245,N_28340);
nand U28806 (N_28806,N_28279,N_28406);
and U28807 (N_28807,N_28321,N_28456);
or U28808 (N_28808,N_28379,N_28433);
nor U28809 (N_28809,N_28370,N_28506);
nand U28810 (N_28810,N_28790,N_28558);
and U28811 (N_28811,N_28538,N_28218);
nand U28812 (N_28812,N_28276,N_28495);
and U28813 (N_28813,N_28785,N_28281);
or U28814 (N_28814,N_28498,N_28718);
or U28815 (N_28815,N_28644,N_28744);
and U28816 (N_28816,N_28601,N_28647);
or U28817 (N_28817,N_28546,N_28743);
nor U28818 (N_28818,N_28761,N_28714);
nand U28819 (N_28819,N_28623,N_28760);
nor U28820 (N_28820,N_28206,N_28637);
nand U28821 (N_28821,N_28753,N_28727);
nand U28822 (N_28822,N_28528,N_28500);
nand U28823 (N_28823,N_28698,N_28795);
and U28824 (N_28824,N_28662,N_28515);
or U28825 (N_28825,N_28338,N_28695);
and U28826 (N_28826,N_28751,N_28421);
and U28827 (N_28827,N_28369,N_28333);
and U28828 (N_28828,N_28277,N_28490);
and U28829 (N_28829,N_28657,N_28548);
and U28830 (N_28830,N_28510,N_28724);
and U28831 (N_28831,N_28287,N_28661);
and U28832 (N_28832,N_28545,N_28678);
nand U28833 (N_28833,N_28308,N_28642);
or U28834 (N_28834,N_28413,N_28241);
nand U28835 (N_28835,N_28658,N_28351);
and U28836 (N_28836,N_28617,N_28215);
or U28837 (N_28837,N_28450,N_28365);
and U28838 (N_28838,N_28765,N_28687);
nand U28839 (N_28839,N_28447,N_28768);
and U28840 (N_28840,N_28242,N_28706);
and U28841 (N_28841,N_28514,N_28350);
and U28842 (N_28842,N_28475,N_28599);
xnor U28843 (N_28843,N_28460,N_28256);
and U28844 (N_28844,N_28366,N_28257);
and U28845 (N_28845,N_28311,N_28651);
or U28846 (N_28846,N_28282,N_28571);
and U28847 (N_28847,N_28532,N_28253);
or U28848 (N_28848,N_28405,N_28569);
nand U28849 (N_28849,N_28305,N_28411);
or U28850 (N_28850,N_28686,N_28564);
nor U28851 (N_28851,N_28621,N_28221);
and U28852 (N_28852,N_28699,N_28534);
and U28853 (N_28853,N_28396,N_28477);
nand U28854 (N_28854,N_28296,N_28696);
and U28855 (N_28855,N_28508,N_28323);
or U28856 (N_28856,N_28665,N_28512);
nand U28857 (N_28857,N_28233,N_28730);
or U28858 (N_28858,N_28463,N_28552);
nor U28859 (N_28859,N_28622,N_28685);
nand U28860 (N_28860,N_28654,N_28720);
nand U28861 (N_28861,N_28234,N_28434);
nor U28862 (N_28862,N_28742,N_28452);
or U28863 (N_28863,N_28430,N_28373);
nand U28864 (N_28864,N_28371,N_28295);
or U28865 (N_28865,N_28645,N_28399);
xor U28866 (N_28866,N_28384,N_28220);
nor U28867 (N_28867,N_28326,N_28388);
nand U28868 (N_28868,N_28354,N_28337);
nand U28869 (N_28869,N_28381,N_28264);
or U28870 (N_28870,N_28292,N_28580);
nand U28871 (N_28871,N_28205,N_28469);
nand U28872 (N_28872,N_28734,N_28641);
or U28873 (N_28873,N_28501,N_28408);
nand U28874 (N_28874,N_28705,N_28598);
and U28875 (N_28875,N_28536,N_28789);
xnor U28876 (N_28876,N_28520,N_28225);
or U28877 (N_28877,N_28227,N_28736);
nor U28878 (N_28878,N_28527,N_28380);
or U28879 (N_28879,N_28378,N_28291);
or U28880 (N_28880,N_28575,N_28219);
nand U28881 (N_28881,N_28325,N_28222);
or U28882 (N_28882,N_28675,N_28588);
nor U28883 (N_28883,N_28697,N_28497);
and U28884 (N_28884,N_28513,N_28492);
or U28885 (N_28885,N_28486,N_28315);
or U28886 (N_28886,N_28583,N_28269);
nor U28887 (N_28887,N_28625,N_28401);
nand U28888 (N_28888,N_28799,N_28737);
nand U28889 (N_28889,N_28339,N_28267);
or U28890 (N_28890,N_28432,N_28638);
nor U28891 (N_28891,N_28355,N_28721);
nor U28892 (N_28892,N_28713,N_28530);
nor U28893 (N_28893,N_28443,N_28398);
or U28894 (N_28894,N_28607,N_28783);
nor U28895 (N_28895,N_28602,N_28758);
nor U28896 (N_28896,N_28493,N_28455);
xor U28897 (N_28897,N_28347,N_28288);
and U28898 (N_28898,N_28551,N_28274);
nor U28899 (N_28899,N_28395,N_28672);
and U28900 (N_28900,N_28336,N_28481);
or U28901 (N_28901,N_28748,N_28467);
nor U28902 (N_28902,N_28230,N_28313);
and U28903 (N_28903,N_28576,N_28591);
and U28904 (N_28904,N_28511,N_28254);
nor U28905 (N_28905,N_28329,N_28435);
nor U28906 (N_28906,N_28509,N_28352);
nor U28907 (N_28907,N_28409,N_28719);
or U28908 (N_28908,N_28605,N_28632);
or U28909 (N_28909,N_28250,N_28286);
or U28910 (N_28910,N_28441,N_28397);
or U28911 (N_28911,N_28201,N_28478);
or U28912 (N_28912,N_28519,N_28717);
nand U28913 (N_28913,N_28494,N_28423);
nand U28914 (N_28914,N_28555,N_28244);
or U28915 (N_28915,N_28579,N_28786);
xor U28916 (N_28916,N_28611,N_28312);
or U28917 (N_28917,N_28680,N_28792);
nand U28918 (N_28918,N_28301,N_28504);
nor U28919 (N_28919,N_28525,N_28248);
and U28920 (N_28920,N_28547,N_28763);
nor U28921 (N_28921,N_28563,N_28483);
xnor U28922 (N_28922,N_28728,N_28470);
nor U28923 (N_28923,N_28702,N_28585);
and U28924 (N_28924,N_28263,N_28375);
nor U28925 (N_28925,N_28733,N_28335);
nor U28926 (N_28926,N_28344,N_28226);
and U28927 (N_28927,N_28209,N_28780);
nand U28928 (N_28928,N_28668,N_28341);
and U28929 (N_28929,N_28353,N_28415);
nand U28930 (N_28930,N_28297,N_28620);
and U28931 (N_28931,N_28703,N_28723);
or U28932 (N_28932,N_28589,N_28797);
nand U28933 (N_28933,N_28453,N_28302);
nor U28934 (N_28934,N_28412,N_28232);
or U28935 (N_28935,N_28400,N_28283);
and U28936 (N_28936,N_28473,N_28779);
and U28937 (N_28937,N_28771,N_28659);
nor U28938 (N_28938,N_28561,N_28541);
or U28939 (N_28939,N_28386,N_28567);
nor U28940 (N_28940,N_28704,N_28382);
nor U28941 (N_28941,N_28449,N_28422);
nor U28942 (N_28942,N_28584,N_28310);
nand U28943 (N_28943,N_28228,N_28667);
or U28944 (N_28944,N_28499,N_28300);
or U28945 (N_28945,N_28726,N_28476);
nor U28946 (N_28946,N_28457,N_28722);
and U28947 (N_28947,N_28327,N_28796);
or U28948 (N_28948,N_28440,N_28739);
nor U28949 (N_28949,N_28677,N_28787);
nor U28950 (N_28950,N_28488,N_28759);
nand U28951 (N_28951,N_28522,N_28314);
or U28952 (N_28952,N_28682,N_28590);
and U28953 (N_28953,N_28643,N_28770);
and U28954 (N_28954,N_28578,N_28749);
nand U28955 (N_28955,N_28289,N_28633);
nand U28956 (N_28956,N_28710,N_28343);
nor U28957 (N_28957,N_28556,N_28480);
nor U28958 (N_28958,N_28461,N_28445);
nor U28959 (N_28959,N_28772,N_28442);
nand U28960 (N_28960,N_28251,N_28729);
nand U28961 (N_28961,N_28752,N_28479);
and U28962 (N_28962,N_28437,N_28627);
nor U28963 (N_28963,N_28273,N_28210);
nand U28964 (N_28964,N_28526,N_28246);
or U28965 (N_28965,N_28524,N_28656);
nand U28966 (N_28966,N_28419,N_28418);
nor U28967 (N_28967,N_28745,N_28290);
or U28968 (N_28968,N_28725,N_28414);
nand U28969 (N_28969,N_28416,N_28581);
nand U28970 (N_28970,N_28207,N_28505);
and U28971 (N_28971,N_28577,N_28631);
or U28972 (N_28972,N_28554,N_28653);
or U28973 (N_28973,N_28781,N_28565);
nand U28974 (N_28974,N_28775,N_28769);
nor U28975 (N_28975,N_28436,N_28258);
nand U28976 (N_28976,N_28424,N_28293);
nand U28977 (N_28977,N_28630,N_28417);
and U28978 (N_28978,N_28238,N_28328);
and U28979 (N_28979,N_28502,N_28663);
nand U28980 (N_28980,N_28691,N_28701);
or U28981 (N_28981,N_28275,N_28367);
nor U28982 (N_28982,N_28420,N_28700);
nor U28983 (N_28983,N_28217,N_28747);
nand U28984 (N_28984,N_28539,N_28609);
nand U28985 (N_28985,N_28235,N_28200);
nand U28986 (N_28986,N_28392,N_28754);
or U28987 (N_28987,N_28778,N_28793);
or U28988 (N_28988,N_28635,N_28618);
nand U28989 (N_28989,N_28383,N_28431);
or U28990 (N_28990,N_28543,N_28262);
nand U28991 (N_28991,N_28655,N_28229);
and U28992 (N_28992,N_28298,N_28307);
nor U28993 (N_28993,N_28342,N_28410);
xor U28994 (N_28994,N_28582,N_28596);
nor U28995 (N_28995,N_28610,N_28688);
or U28996 (N_28996,N_28639,N_28252);
nand U28997 (N_28997,N_28741,N_28766);
nor U28998 (N_28998,N_28650,N_28331);
or U28999 (N_28999,N_28427,N_28407);
nor U29000 (N_29000,N_28303,N_28626);
or U29001 (N_29001,N_28446,N_28223);
and U29002 (N_29002,N_28224,N_28603);
nand U29003 (N_29003,N_28346,N_28542);
and U29004 (N_29004,N_28648,N_28531);
and U29005 (N_29005,N_28597,N_28683);
nor U29006 (N_29006,N_28604,N_28214);
nand U29007 (N_29007,N_28249,N_28798);
nand U29008 (N_29008,N_28709,N_28272);
nand U29009 (N_29009,N_28390,N_28784);
nor U29010 (N_29010,N_28372,N_28204);
and U29011 (N_29011,N_28472,N_28774);
and U29012 (N_29012,N_28304,N_28360);
and U29013 (N_29013,N_28348,N_28762);
and U29014 (N_29014,N_28776,N_28593);
nor U29015 (N_29015,N_28374,N_28482);
nor U29016 (N_29016,N_28237,N_28389);
nor U29017 (N_29017,N_28491,N_28208);
nand U29018 (N_29018,N_28592,N_28213);
or U29019 (N_29019,N_28791,N_28594);
nand U29020 (N_29020,N_28516,N_28690);
nand U29021 (N_29021,N_28364,N_28299);
nand U29022 (N_29022,N_28271,N_28523);
nand U29023 (N_29023,N_28557,N_28402);
nand U29024 (N_29024,N_28606,N_28629);
nor U29025 (N_29025,N_28268,N_28608);
or U29026 (N_29026,N_28533,N_28612);
nor U29027 (N_29027,N_28624,N_28731);
nor U29028 (N_29028,N_28586,N_28681);
nor U29029 (N_29029,N_28693,N_28465);
or U29030 (N_29030,N_28361,N_28535);
nand U29031 (N_29031,N_28464,N_28777);
nor U29032 (N_29032,N_28270,N_28517);
and U29033 (N_29033,N_28708,N_28451);
and U29034 (N_29034,N_28489,N_28484);
nor U29035 (N_29035,N_28485,N_28572);
and U29036 (N_29036,N_28521,N_28646);
nand U29037 (N_29037,N_28694,N_28711);
or U29038 (N_29038,N_28587,N_28255);
and U29039 (N_29039,N_28507,N_28757);
or U29040 (N_29040,N_28679,N_28294);
nor U29041 (N_29041,N_28550,N_28503);
and U29042 (N_29042,N_28203,N_28319);
or U29043 (N_29043,N_28318,N_28544);
and U29044 (N_29044,N_28385,N_28448);
or U29045 (N_29045,N_28549,N_28767);
nand U29046 (N_29046,N_28559,N_28332);
and U29047 (N_29047,N_28707,N_28362);
nor U29048 (N_29048,N_28560,N_28738);
nor U29049 (N_29049,N_28540,N_28574);
or U29050 (N_29050,N_28356,N_28358);
and U29051 (N_29051,N_28740,N_28496);
nand U29052 (N_29052,N_28712,N_28670);
and U29053 (N_29053,N_28359,N_28750);
or U29054 (N_29054,N_28773,N_28231);
and U29055 (N_29055,N_28278,N_28628);
xor U29056 (N_29056,N_28518,N_28649);
and U29057 (N_29057,N_28334,N_28616);
or U29058 (N_29058,N_28674,N_28756);
nand U29059 (N_29059,N_28466,N_28428);
or U29060 (N_29060,N_28553,N_28474);
and U29061 (N_29061,N_28316,N_28689);
and U29062 (N_29062,N_28322,N_28471);
and U29063 (N_29063,N_28261,N_28614);
nand U29064 (N_29064,N_28345,N_28317);
nand U29065 (N_29065,N_28349,N_28202);
and U29066 (N_29066,N_28652,N_28426);
or U29067 (N_29067,N_28216,N_28468);
and U29068 (N_29068,N_28755,N_28438);
nor U29069 (N_29069,N_28615,N_28243);
or U29070 (N_29070,N_28377,N_28487);
and U29071 (N_29071,N_28746,N_28666);
or U29072 (N_29072,N_28280,N_28247);
nor U29073 (N_29073,N_28259,N_28239);
and U29074 (N_29074,N_28684,N_28454);
nand U29075 (N_29075,N_28459,N_28260);
and U29076 (N_29076,N_28265,N_28330);
nor U29077 (N_29077,N_28562,N_28671);
and U29078 (N_29078,N_28240,N_28595);
or U29079 (N_29079,N_28394,N_28764);
nand U29080 (N_29080,N_28368,N_28794);
and U29081 (N_29081,N_28393,N_28537);
nor U29082 (N_29082,N_28425,N_28285);
or U29083 (N_29083,N_28788,N_28732);
or U29084 (N_29084,N_28391,N_28306);
and U29085 (N_29085,N_28357,N_28444);
nand U29086 (N_29086,N_28619,N_28636);
nor U29087 (N_29087,N_28568,N_28692);
or U29088 (N_29088,N_28566,N_28284);
and U29089 (N_29089,N_28782,N_28529);
nand U29090 (N_29090,N_28363,N_28669);
and U29091 (N_29091,N_28266,N_28613);
or U29092 (N_29092,N_28429,N_28211);
or U29093 (N_29093,N_28439,N_28324);
or U29094 (N_29094,N_28309,N_28716);
or U29095 (N_29095,N_28320,N_28462);
nand U29096 (N_29096,N_28676,N_28634);
nor U29097 (N_29097,N_28640,N_28212);
or U29098 (N_29098,N_28573,N_28673);
and U29099 (N_29099,N_28735,N_28715);
nand U29100 (N_29100,N_28625,N_28431);
and U29101 (N_29101,N_28373,N_28718);
nor U29102 (N_29102,N_28412,N_28530);
nor U29103 (N_29103,N_28624,N_28554);
or U29104 (N_29104,N_28356,N_28289);
or U29105 (N_29105,N_28570,N_28495);
nand U29106 (N_29106,N_28252,N_28705);
nor U29107 (N_29107,N_28719,N_28229);
nor U29108 (N_29108,N_28377,N_28472);
and U29109 (N_29109,N_28702,N_28319);
or U29110 (N_29110,N_28697,N_28590);
nor U29111 (N_29111,N_28376,N_28427);
and U29112 (N_29112,N_28622,N_28207);
or U29113 (N_29113,N_28470,N_28323);
nand U29114 (N_29114,N_28521,N_28686);
nand U29115 (N_29115,N_28312,N_28795);
nand U29116 (N_29116,N_28732,N_28771);
or U29117 (N_29117,N_28508,N_28520);
xor U29118 (N_29118,N_28664,N_28203);
nand U29119 (N_29119,N_28298,N_28447);
nor U29120 (N_29120,N_28617,N_28376);
or U29121 (N_29121,N_28654,N_28504);
or U29122 (N_29122,N_28237,N_28395);
or U29123 (N_29123,N_28459,N_28554);
nor U29124 (N_29124,N_28741,N_28644);
or U29125 (N_29125,N_28381,N_28451);
or U29126 (N_29126,N_28712,N_28506);
nand U29127 (N_29127,N_28449,N_28301);
nor U29128 (N_29128,N_28253,N_28288);
and U29129 (N_29129,N_28271,N_28471);
or U29130 (N_29130,N_28411,N_28463);
nor U29131 (N_29131,N_28227,N_28608);
nand U29132 (N_29132,N_28611,N_28431);
nor U29133 (N_29133,N_28708,N_28325);
nor U29134 (N_29134,N_28221,N_28510);
and U29135 (N_29135,N_28778,N_28252);
or U29136 (N_29136,N_28223,N_28756);
nand U29137 (N_29137,N_28312,N_28213);
and U29138 (N_29138,N_28402,N_28773);
nor U29139 (N_29139,N_28556,N_28607);
nand U29140 (N_29140,N_28577,N_28486);
nor U29141 (N_29141,N_28360,N_28278);
or U29142 (N_29142,N_28748,N_28306);
or U29143 (N_29143,N_28431,N_28341);
and U29144 (N_29144,N_28422,N_28595);
nand U29145 (N_29145,N_28722,N_28582);
nor U29146 (N_29146,N_28505,N_28425);
xnor U29147 (N_29147,N_28501,N_28415);
nand U29148 (N_29148,N_28413,N_28227);
and U29149 (N_29149,N_28477,N_28744);
nor U29150 (N_29150,N_28334,N_28794);
and U29151 (N_29151,N_28606,N_28657);
and U29152 (N_29152,N_28350,N_28620);
nand U29153 (N_29153,N_28708,N_28510);
xnor U29154 (N_29154,N_28703,N_28518);
nor U29155 (N_29155,N_28752,N_28575);
and U29156 (N_29156,N_28504,N_28706);
nor U29157 (N_29157,N_28238,N_28467);
nor U29158 (N_29158,N_28525,N_28670);
xor U29159 (N_29159,N_28536,N_28492);
or U29160 (N_29160,N_28296,N_28343);
or U29161 (N_29161,N_28640,N_28375);
and U29162 (N_29162,N_28488,N_28674);
and U29163 (N_29163,N_28700,N_28374);
nor U29164 (N_29164,N_28247,N_28549);
nand U29165 (N_29165,N_28597,N_28311);
and U29166 (N_29166,N_28411,N_28670);
nand U29167 (N_29167,N_28702,N_28436);
nand U29168 (N_29168,N_28409,N_28332);
nand U29169 (N_29169,N_28649,N_28367);
or U29170 (N_29170,N_28672,N_28662);
or U29171 (N_29171,N_28732,N_28384);
nor U29172 (N_29172,N_28670,N_28709);
nor U29173 (N_29173,N_28399,N_28332);
nor U29174 (N_29174,N_28373,N_28211);
nor U29175 (N_29175,N_28234,N_28419);
or U29176 (N_29176,N_28637,N_28333);
or U29177 (N_29177,N_28468,N_28442);
or U29178 (N_29178,N_28500,N_28483);
nand U29179 (N_29179,N_28338,N_28585);
nand U29180 (N_29180,N_28576,N_28233);
nor U29181 (N_29181,N_28433,N_28279);
xor U29182 (N_29182,N_28220,N_28517);
and U29183 (N_29183,N_28448,N_28522);
nand U29184 (N_29184,N_28411,N_28473);
nand U29185 (N_29185,N_28421,N_28333);
nand U29186 (N_29186,N_28228,N_28578);
nor U29187 (N_29187,N_28744,N_28390);
nand U29188 (N_29188,N_28659,N_28261);
nand U29189 (N_29189,N_28473,N_28496);
nand U29190 (N_29190,N_28746,N_28649);
xor U29191 (N_29191,N_28422,N_28371);
or U29192 (N_29192,N_28256,N_28285);
nand U29193 (N_29193,N_28578,N_28579);
or U29194 (N_29194,N_28341,N_28224);
and U29195 (N_29195,N_28663,N_28799);
nor U29196 (N_29196,N_28581,N_28250);
or U29197 (N_29197,N_28468,N_28501);
or U29198 (N_29198,N_28529,N_28206);
nor U29199 (N_29199,N_28566,N_28658);
or U29200 (N_29200,N_28420,N_28258);
or U29201 (N_29201,N_28703,N_28730);
and U29202 (N_29202,N_28516,N_28312);
nor U29203 (N_29203,N_28592,N_28701);
nand U29204 (N_29204,N_28394,N_28736);
and U29205 (N_29205,N_28429,N_28435);
nor U29206 (N_29206,N_28733,N_28429);
xnor U29207 (N_29207,N_28207,N_28787);
nand U29208 (N_29208,N_28412,N_28629);
and U29209 (N_29209,N_28504,N_28291);
nand U29210 (N_29210,N_28772,N_28678);
nor U29211 (N_29211,N_28298,N_28599);
nor U29212 (N_29212,N_28209,N_28781);
nor U29213 (N_29213,N_28380,N_28620);
nand U29214 (N_29214,N_28728,N_28741);
nand U29215 (N_29215,N_28655,N_28707);
nor U29216 (N_29216,N_28203,N_28792);
and U29217 (N_29217,N_28709,N_28233);
or U29218 (N_29218,N_28733,N_28491);
and U29219 (N_29219,N_28702,N_28581);
or U29220 (N_29220,N_28254,N_28721);
nand U29221 (N_29221,N_28383,N_28421);
and U29222 (N_29222,N_28398,N_28221);
nor U29223 (N_29223,N_28353,N_28715);
and U29224 (N_29224,N_28357,N_28549);
and U29225 (N_29225,N_28322,N_28461);
or U29226 (N_29226,N_28212,N_28228);
nor U29227 (N_29227,N_28438,N_28678);
or U29228 (N_29228,N_28397,N_28342);
and U29229 (N_29229,N_28262,N_28600);
and U29230 (N_29230,N_28700,N_28730);
or U29231 (N_29231,N_28296,N_28387);
or U29232 (N_29232,N_28666,N_28299);
nand U29233 (N_29233,N_28254,N_28256);
or U29234 (N_29234,N_28781,N_28779);
nand U29235 (N_29235,N_28699,N_28594);
nand U29236 (N_29236,N_28300,N_28648);
nand U29237 (N_29237,N_28529,N_28774);
xor U29238 (N_29238,N_28614,N_28293);
nor U29239 (N_29239,N_28744,N_28541);
nand U29240 (N_29240,N_28681,N_28528);
or U29241 (N_29241,N_28778,N_28404);
nor U29242 (N_29242,N_28583,N_28272);
nor U29243 (N_29243,N_28578,N_28297);
nand U29244 (N_29244,N_28522,N_28561);
and U29245 (N_29245,N_28676,N_28596);
or U29246 (N_29246,N_28336,N_28442);
or U29247 (N_29247,N_28230,N_28342);
and U29248 (N_29248,N_28733,N_28374);
nand U29249 (N_29249,N_28417,N_28511);
or U29250 (N_29250,N_28793,N_28443);
nor U29251 (N_29251,N_28436,N_28430);
nor U29252 (N_29252,N_28442,N_28581);
nand U29253 (N_29253,N_28363,N_28410);
and U29254 (N_29254,N_28437,N_28293);
or U29255 (N_29255,N_28699,N_28741);
or U29256 (N_29256,N_28597,N_28611);
nor U29257 (N_29257,N_28443,N_28470);
and U29258 (N_29258,N_28250,N_28698);
nor U29259 (N_29259,N_28388,N_28451);
xor U29260 (N_29260,N_28249,N_28522);
or U29261 (N_29261,N_28388,N_28452);
nor U29262 (N_29262,N_28409,N_28276);
xnor U29263 (N_29263,N_28297,N_28295);
and U29264 (N_29264,N_28550,N_28745);
or U29265 (N_29265,N_28792,N_28507);
or U29266 (N_29266,N_28783,N_28212);
or U29267 (N_29267,N_28688,N_28442);
and U29268 (N_29268,N_28227,N_28429);
or U29269 (N_29269,N_28305,N_28750);
nand U29270 (N_29270,N_28340,N_28444);
nand U29271 (N_29271,N_28344,N_28708);
and U29272 (N_29272,N_28723,N_28508);
nor U29273 (N_29273,N_28542,N_28590);
xor U29274 (N_29274,N_28701,N_28394);
nor U29275 (N_29275,N_28215,N_28323);
or U29276 (N_29276,N_28350,N_28252);
and U29277 (N_29277,N_28772,N_28344);
and U29278 (N_29278,N_28502,N_28504);
or U29279 (N_29279,N_28207,N_28662);
and U29280 (N_29280,N_28640,N_28682);
nor U29281 (N_29281,N_28563,N_28701);
nor U29282 (N_29282,N_28526,N_28620);
or U29283 (N_29283,N_28474,N_28701);
or U29284 (N_29284,N_28426,N_28265);
or U29285 (N_29285,N_28545,N_28264);
and U29286 (N_29286,N_28666,N_28727);
nor U29287 (N_29287,N_28735,N_28455);
and U29288 (N_29288,N_28323,N_28656);
or U29289 (N_29289,N_28530,N_28247);
and U29290 (N_29290,N_28750,N_28351);
and U29291 (N_29291,N_28407,N_28308);
and U29292 (N_29292,N_28284,N_28458);
and U29293 (N_29293,N_28558,N_28601);
or U29294 (N_29294,N_28457,N_28464);
and U29295 (N_29295,N_28774,N_28271);
or U29296 (N_29296,N_28217,N_28451);
nor U29297 (N_29297,N_28202,N_28387);
nand U29298 (N_29298,N_28467,N_28253);
nor U29299 (N_29299,N_28587,N_28428);
nor U29300 (N_29300,N_28575,N_28735);
nor U29301 (N_29301,N_28403,N_28733);
nor U29302 (N_29302,N_28566,N_28334);
or U29303 (N_29303,N_28592,N_28710);
nand U29304 (N_29304,N_28338,N_28464);
or U29305 (N_29305,N_28757,N_28760);
nor U29306 (N_29306,N_28279,N_28665);
and U29307 (N_29307,N_28552,N_28644);
and U29308 (N_29308,N_28352,N_28235);
or U29309 (N_29309,N_28669,N_28756);
and U29310 (N_29310,N_28239,N_28368);
and U29311 (N_29311,N_28335,N_28275);
nand U29312 (N_29312,N_28230,N_28282);
nand U29313 (N_29313,N_28229,N_28454);
or U29314 (N_29314,N_28448,N_28260);
or U29315 (N_29315,N_28620,N_28363);
nor U29316 (N_29316,N_28447,N_28468);
xor U29317 (N_29317,N_28467,N_28519);
or U29318 (N_29318,N_28277,N_28298);
nand U29319 (N_29319,N_28776,N_28545);
nor U29320 (N_29320,N_28285,N_28443);
or U29321 (N_29321,N_28721,N_28540);
or U29322 (N_29322,N_28419,N_28596);
or U29323 (N_29323,N_28659,N_28514);
nand U29324 (N_29324,N_28293,N_28612);
nand U29325 (N_29325,N_28499,N_28784);
nand U29326 (N_29326,N_28646,N_28700);
or U29327 (N_29327,N_28416,N_28541);
nor U29328 (N_29328,N_28572,N_28538);
nor U29329 (N_29329,N_28379,N_28776);
nand U29330 (N_29330,N_28399,N_28610);
or U29331 (N_29331,N_28233,N_28739);
or U29332 (N_29332,N_28506,N_28327);
or U29333 (N_29333,N_28216,N_28439);
nor U29334 (N_29334,N_28760,N_28383);
or U29335 (N_29335,N_28447,N_28712);
nand U29336 (N_29336,N_28205,N_28595);
nand U29337 (N_29337,N_28580,N_28724);
and U29338 (N_29338,N_28332,N_28201);
nand U29339 (N_29339,N_28687,N_28416);
and U29340 (N_29340,N_28364,N_28664);
nor U29341 (N_29341,N_28451,N_28727);
and U29342 (N_29342,N_28700,N_28422);
and U29343 (N_29343,N_28691,N_28325);
nand U29344 (N_29344,N_28757,N_28693);
or U29345 (N_29345,N_28747,N_28639);
nand U29346 (N_29346,N_28736,N_28696);
nor U29347 (N_29347,N_28678,N_28225);
nand U29348 (N_29348,N_28470,N_28545);
nand U29349 (N_29349,N_28678,N_28777);
or U29350 (N_29350,N_28211,N_28691);
nand U29351 (N_29351,N_28255,N_28369);
nor U29352 (N_29352,N_28410,N_28739);
nor U29353 (N_29353,N_28749,N_28547);
nor U29354 (N_29354,N_28516,N_28287);
and U29355 (N_29355,N_28470,N_28400);
nand U29356 (N_29356,N_28570,N_28523);
nand U29357 (N_29357,N_28633,N_28785);
and U29358 (N_29358,N_28577,N_28594);
xor U29359 (N_29359,N_28722,N_28669);
and U29360 (N_29360,N_28757,N_28674);
or U29361 (N_29361,N_28726,N_28797);
nand U29362 (N_29362,N_28224,N_28767);
nand U29363 (N_29363,N_28770,N_28792);
nor U29364 (N_29364,N_28409,N_28670);
or U29365 (N_29365,N_28367,N_28230);
or U29366 (N_29366,N_28499,N_28331);
nor U29367 (N_29367,N_28785,N_28663);
nand U29368 (N_29368,N_28680,N_28328);
and U29369 (N_29369,N_28686,N_28441);
xor U29370 (N_29370,N_28296,N_28247);
nand U29371 (N_29371,N_28491,N_28323);
and U29372 (N_29372,N_28275,N_28622);
nor U29373 (N_29373,N_28348,N_28392);
nor U29374 (N_29374,N_28233,N_28472);
or U29375 (N_29375,N_28696,N_28699);
xnor U29376 (N_29376,N_28428,N_28784);
and U29377 (N_29377,N_28610,N_28253);
nor U29378 (N_29378,N_28649,N_28398);
or U29379 (N_29379,N_28596,N_28680);
nand U29380 (N_29380,N_28554,N_28628);
nand U29381 (N_29381,N_28602,N_28749);
or U29382 (N_29382,N_28740,N_28402);
or U29383 (N_29383,N_28228,N_28519);
and U29384 (N_29384,N_28674,N_28361);
xnor U29385 (N_29385,N_28497,N_28510);
xnor U29386 (N_29386,N_28315,N_28653);
and U29387 (N_29387,N_28284,N_28332);
nand U29388 (N_29388,N_28621,N_28518);
nor U29389 (N_29389,N_28532,N_28297);
or U29390 (N_29390,N_28591,N_28595);
nor U29391 (N_29391,N_28586,N_28351);
or U29392 (N_29392,N_28310,N_28446);
nand U29393 (N_29393,N_28747,N_28283);
or U29394 (N_29394,N_28501,N_28667);
nor U29395 (N_29395,N_28229,N_28479);
nand U29396 (N_29396,N_28551,N_28318);
nand U29397 (N_29397,N_28652,N_28575);
and U29398 (N_29398,N_28773,N_28255);
and U29399 (N_29399,N_28322,N_28544);
nor U29400 (N_29400,N_29029,N_29169);
and U29401 (N_29401,N_28996,N_29046);
nand U29402 (N_29402,N_28862,N_29385);
or U29403 (N_29403,N_29135,N_29311);
nand U29404 (N_29404,N_28885,N_29147);
and U29405 (N_29405,N_29065,N_29032);
or U29406 (N_29406,N_29093,N_29172);
and U29407 (N_29407,N_28886,N_28961);
or U29408 (N_29408,N_29320,N_29001);
and U29409 (N_29409,N_29200,N_29085);
or U29410 (N_29410,N_29387,N_28873);
nor U29411 (N_29411,N_29013,N_28867);
nor U29412 (N_29412,N_29342,N_29055);
nand U29413 (N_29413,N_29313,N_28874);
or U29414 (N_29414,N_29073,N_29347);
nor U29415 (N_29415,N_29116,N_28808);
and U29416 (N_29416,N_29341,N_29136);
nor U29417 (N_29417,N_29301,N_29272);
or U29418 (N_29418,N_28810,N_29047);
nand U29419 (N_29419,N_28868,N_29010);
and U29420 (N_29420,N_29023,N_29294);
nand U29421 (N_29421,N_29042,N_29119);
nand U29422 (N_29422,N_29212,N_29120);
or U29423 (N_29423,N_29143,N_29340);
or U29424 (N_29424,N_29367,N_29397);
and U29425 (N_29425,N_29243,N_29239);
and U29426 (N_29426,N_29148,N_29319);
nand U29427 (N_29427,N_29198,N_29140);
or U29428 (N_29428,N_29356,N_29197);
nand U29429 (N_29429,N_29184,N_29051);
nor U29430 (N_29430,N_29209,N_28872);
nand U29431 (N_29431,N_28849,N_29003);
and U29432 (N_29432,N_29314,N_29078);
nand U29433 (N_29433,N_28954,N_29327);
and U29434 (N_29434,N_28894,N_29063);
nor U29435 (N_29435,N_29205,N_28821);
and U29436 (N_29436,N_29274,N_29287);
nor U29437 (N_29437,N_29052,N_29025);
nor U29438 (N_29438,N_29081,N_28822);
or U29439 (N_29439,N_29258,N_28817);
nor U29440 (N_29440,N_28850,N_29203);
or U29441 (N_29441,N_29333,N_28933);
or U29442 (N_29442,N_29168,N_29237);
or U29443 (N_29443,N_28820,N_28823);
nor U29444 (N_29444,N_29335,N_28999);
nand U29445 (N_29445,N_29157,N_29303);
and U29446 (N_29446,N_28837,N_29176);
or U29447 (N_29447,N_29229,N_29125);
nand U29448 (N_29448,N_29087,N_29286);
nor U29449 (N_29449,N_28920,N_29145);
or U29450 (N_29450,N_29280,N_28847);
or U29451 (N_29451,N_29056,N_29040);
and U29452 (N_29452,N_28912,N_29097);
or U29453 (N_29453,N_29260,N_29088);
nor U29454 (N_29454,N_28935,N_29139);
and U29455 (N_29455,N_29371,N_29373);
nor U29456 (N_29456,N_28898,N_28905);
or U29457 (N_29457,N_29207,N_28835);
or U29458 (N_29458,N_29393,N_29376);
nor U29459 (N_29459,N_29283,N_29045);
nand U29460 (N_29460,N_29338,N_28809);
and U29461 (N_29461,N_29105,N_29251);
nand U29462 (N_29462,N_29284,N_29226);
and U29463 (N_29463,N_29104,N_28976);
nor U29464 (N_29464,N_29219,N_28942);
or U29465 (N_29465,N_29192,N_29043);
xor U29466 (N_29466,N_29038,N_29034);
nand U29467 (N_29467,N_29107,N_29016);
nand U29468 (N_29468,N_28978,N_28969);
and U29469 (N_29469,N_28975,N_29378);
xor U29470 (N_29470,N_29112,N_29066);
and U29471 (N_29471,N_28930,N_29254);
nand U29472 (N_29472,N_28901,N_29354);
nor U29473 (N_29473,N_29196,N_29384);
nor U29474 (N_29474,N_29020,N_28829);
nand U29475 (N_29475,N_28981,N_29372);
nand U29476 (N_29476,N_29344,N_29253);
nand U29477 (N_29477,N_28892,N_29162);
nor U29478 (N_29478,N_29309,N_29129);
or U29479 (N_29479,N_28889,N_28914);
nor U29480 (N_29480,N_28962,N_29185);
nand U29481 (N_29481,N_28923,N_29211);
nor U29482 (N_29482,N_28876,N_28921);
nand U29483 (N_29483,N_28988,N_29221);
and U29484 (N_29484,N_28979,N_29110);
nand U29485 (N_29485,N_28811,N_29059);
nand U29486 (N_29486,N_29270,N_29101);
nand U29487 (N_29487,N_29188,N_29318);
nand U29488 (N_29488,N_29252,N_28986);
and U29489 (N_29489,N_28842,N_29131);
or U29490 (N_29490,N_29095,N_29322);
nand U29491 (N_29491,N_29144,N_29083);
nand U29492 (N_29492,N_29236,N_29193);
nand U29493 (N_29493,N_29127,N_29288);
nor U29494 (N_29494,N_29050,N_29109);
nor U29495 (N_29495,N_29033,N_29346);
nor U29496 (N_29496,N_28993,N_29194);
or U29497 (N_29497,N_29114,N_28927);
and U29498 (N_29498,N_28841,N_28870);
or U29499 (N_29499,N_29111,N_28917);
nand U29500 (N_29500,N_29289,N_29343);
nand U29501 (N_29501,N_29015,N_29302);
nor U29502 (N_29502,N_28989,N_28970);
and U29503 (N_29503,N_29156,N_29262);
or U29504 (N_29504,N_29227,N_29218);
or U29505 (N_29505,N_28906,N_28839);
nand U29506 (N_29506,N_28893,N_29080);
or U29507 (N_29507,N_29382,N_29171);
or U29508 (N_29508,N_28858,N_28866);
nand U29509 (N_29509,N_29255,N_28852);
nor U29510 (N_29510,N_28967,N_28955);
or U29511 (N_29511,N_29024,N_29079);
nand U29512 (N_29512,N_29297,N_29041);
and U29513 (N_29513,N_29021,N_29113);
nand U29514 (N_29514,N_28836,N_29053);
nand U29515 (N_29515,N_29009,N_29357);
and U29516 (N_29516,N_29155,N_29233);
and U29517 (N_29517,N_29293,N_28825);
nor U29518 (N_29518,N_29177,N_28803);
and U29519 (N_29519,N_28851,N_29091);
or U29520 (N_29520,N_28983,N_29228);
and U29521 (N_29521,N_29365,N_29049);
nor U29522 (N_29522,N_28958,N_28884);
nor U29523 (N_29523,N_29395,N_28888);
nand U29524 (N_29524,N_29183,N_28953);
nand U29525 (N_29525,N_29214,N_29012);
and U29526 (N_29526,N_29290,N_28949);
and U29527 (N_29527,N_29123,N_29108);
or U29528 (N_29528,N_29115,N_29000);
or U29529 (N_29529,N_29334,N_29307);
or U29530 (N_29530,N_29216,N_28907);
nand U29531 (N_29531,N_28840,N_29142);
nor U29532 (N_29532,N_28992,N_29077);
or U29533 (N_29533,N_28819,N_28816);
or U29534 (N_29534,N_29208,N_28944);
nor U29535 (N_29535,N_29121,N_28934);
and U29536 (N_29536,N_28990,N_29076);
nor U29537 (N_29537,N_29019,N_28966);
or U29538 (N_29538,N_29030,N_29360);
nor U29539 (N_29539,N_29086,N_28952);
nand U29540 (N_29540,N_29153,N_29035);
or U29541 (N_29541,N_28913,N_28865);
or U29542 (N_29542,N_29008,N_28982);
nand U29543 (N_29543,N_29304,N_29323);
nor U29544 (N_29544,N_28895,N_29225);
nor U29545 (N_29545,N_28972,N_29224);
or U29546 (N_29546,N_28991,N_29231);
nand U29547 (N_29547,N_29339,N_29275);
or U29548 (N_29548,N_28887,N_28924);
or U29549 (N_29549,N_29069,N_29386);
and U29550 (N_29550,N_29150,N_29247);
nand U29551 (N_29551,N_29261,N_29092);
nand U29552 (N_29552,N_28959,N_29256);
nor U29553 (N_29553,N_29285,N_29217);
nor U29554 (N_29554,N_29291,N_29295);
or U29555 (N_29555,N_29223,N_29039);
nand U29556 (N_29556,N_29308,N_28857);
nand U29557 (N_29557,N_28878,N_28916);
or U29558 (N_29558,N_29158,N_28891);
nor U29559 (N_29559,N_28964,N_29004);
or U29560 (N_29560,N_28879,N_29244);
nor U29561 (N_29561,N_29048,N_29186);
nand U29562 (N_29562,N_28883,N_29175);
nand U29563 (N_29563,N_28807,N_29234);
nand U29564 (N_29564,N_29266,N_29054);
or U29565 (N_29565,N_28815,N_29130);
nor U29566 (N_29566,N_29369,N_28998);
nand U29567 (N_29567,N_29267,N_28896);
or U29568 (N_29568,N_29241,N_29324);
nand U29569 (N_29569,N_29392,N_29279);
and U29570 (N_29570,N_28802,N_29232);
nor U29571 (N_29571,N_29202,N_29263);
and U29572 (N_29572,N_29213,N_28931);
nand U29573 (N_29573,N_28801,N_29165);
or U29574 (N_29574,N_29368,N_29161);
or U29575 (N_29575,N_29242,N_29206);
or U29576 (N_29576,N_28985,N_29014);
nor U29577 (N_29577,N_29329,N_29248);
nand U29578 (N_29578,N_28994,N_29364);
or U29579 (N_29579,N_29278,N_28938);
or U29580 (N_29580,N_28956,N_28846);
or U29581 (N_29581,N_28939,N_29160);
nand U29582 (N_29582,N_29174,N_28827);
or U29583 (N_29583,N_28854,N_28824);
nand U29584 (N_29584,N_29068,N_28831);
or U29585 (N_29585,N_28848,N_29235);
nand U29586 (N_29586,N_29190,N_28909);
nand U29587 (N_29587,N_28928,N_29271);
or U29588 (N_29588,N_28936,N_29074);
and U29589 (N_29589,N_29268,N_29179);
or U29590 (N_29590,N_28863,N_28818);
or U29591 (N_29591,N_29399,N_29173);
nand U29592 (N_29592,N_29067,N_29096);
nor U29593 (N_29593,N_29375,N_28864);
or U29594 (N_29594,N_29103,N_29210);
and U29595 (N_29595,N_29022,N_29292);
and U29596 (N_29596,N_28828,N_29006);
nand U29597 (N_29597,N_29383,N_28869);
nor U29598 (N_29598,N_29259,N_29352);
and U29599 (N_29599,N_29027,N_28945);
nor U29600 (N_29600,N_29351,N_29363);
nand U29601 (N_29601,N_29277,N_29305);
nand U29602 (N_29602,N_29379,N_29299);
and U29603 (N_29603,N_29181,N_29321);
nand U29604 (N_29604,N_29037,N_28877);
nand U29605 (N_29605,N_29315,N_29370);
nor U29606 (N_29606,N_29090,N_29276);
and U29607 (N_29607,N_29359,N_28833);
or U29608 (N_29608,N_28908,N_29124);
nand U29609 (N_29609,N_28910,N_28844);
and U29610 (N_29610,N_29220,N_29316);
nand U29611 (N_29611,N_29164,N_29222);
nand U29612 (N_29612,N_28903,N_29170);
nand U29613 (N_29613,N_28843,N_29134);
and U29614 (N_29614,N_28980,N_28919);
or U29615 (N_29615,N_28984,N_29337);
and U29616 (N_29616,N_29132,N_29345);
nand U29617 (N_29617,N_28814,N_29163);
nand U29618 (N_29618,N_29167,N_29374);
nor U29619 (N_29619,N_29326,N_29036);
and U29620 (N_29620,N_28915,N_28918);
and U29621 (N_29621,N_28951,N_29180);
nor U29622 (N_29622,N_28875,N_29099);
nor U29623 (N_29623,N_29366,N_28871);
nor U29624 (N_29624,N_29018,N_29269);
nor U29625 (N_29625,N_28861,N_28890);
nand U29626 (N_29626,N_29350,N_29146);
and U29627 (N_29627,N_29159,N_29058);
and U29628 (N_29628,N_29215,N_29098);
nand U29629 (N_29629,N_29011,N_29298);
and U29630 (N_29630,N_28832,N_29317);
nor U29631 (N_29631,N_28900,N_29355);
and U29632 (N_29632,N_28973,N_28950);
nand U29633 (N_29633,N_28812,N_28881);
or U29634 (N_29634,N_29361,N_29250);
nor U29635 (N_29635,N_28806,N_28940);
and U29636 (N_29636,N_29151,N_29204);
or U29637 (N_29637,N_28859,N_29362);
and U29638 (N_29638,N_29191,N_29389);
or U29639 (N_29639,N_29102,N_28880);
nand U29640 (N_29640,N_29028,N_29187);
nor U29641 (N_29641,N_29031,N_28929);
and U29642 (N_29642,N_29348,N_28804);
or U29643 (N_29643,N_29166,N_28977);
xnor U29644 (N_29644,N_28826,N_29330);
nand U29645 (N_29645,N_29336,N_28995);
nor U29646 (N_29646,N_28960,N_29017);
nor U29647 (N_29647,N_28856,N_29398);
and U29648 (N_29648,N_29118,N_29082);
nor U29649 (N_29649,N_28947,N_29332);
or U29650 (N_29650,N_29089,N_29281);
or U29651 (N_29651,N_29388,N_28926);
nand U29652 (N_29652,N_29353,N_28957);
or U29653 (N_29653,N_29061,N_29312);
nor U29654 (N_29654,N_28965,N_29245);
or U29655 (N_29655,N_28834,N_28813);
or U29656 (N_29656,N_29396,N_29084);
nand U29657 (N_29657,N_28902,N_29182);
or U29658 (N_29658,N_28911,N_29265);
and U29659 (N_29659,N_28922,N_28925);
nand U29660 (N_29660,N_29117,N_28805);
and U29661 (N_29661,N_29189,N_29230);
nand U29662 (N_29662,N_29005,N_29195);
nor U29663 (N_29663,N_29094,N_29381);
or U29664 (N_29664,N_29358,N_29377);
nor U29665 (N_29665,N_29325,N_29257);
or U29666 (N_29666,N_29300,N_29154);
nor U29667 (N_29667,N_29310,N_29044);
nor U29668 (N_29668,N_29390,N_28830);
and U29669 (N_29669,N_29126,N_28882);
or U29670 (N_29670,N_29328,N_28948);
nor U29671 (N_29671,N_29149,N_29273);
nor U29672 (N_29672,N_28838,N_29057);
nand U29673 (N_29673,N_29122,N_29002);
nor U29674 (N_29674,N_29026,N_29201);
xnor U29675 (N_29675,N_29240,N_28974);
nor U29676 (N_29676,N_28800,N_29075);
nand U29677 (N_29677,N_29152,N_29296);
or U29678 (N_29678,N_28971,N_28860);
nand U29679 (N_29679,N_28946,N_29106);
nand U29680 (N_29680,N_29070,N_28899);
nand U29681 (N_29681,N_29178,N_29349);
nand U29682 (N_29682,N_28968,N_29394);
and U29683 (N_29683,N_29007,N_29282);
and U29684 (N_29684,N_28845,N_28855);
xor U29685 (N_29685,N_29137,N_29380);
or U29686 (N_29686,N_29246,N_29141);
and U29687 (N_29687,N_29238,N_29100);
nor U29688 (N_29688,N_29391,N_28943);
nor U29689 (N_29689,N_28897,N_29199);
nand U29690 (N_29690,N_28932,N_28937);
or U29691 (N_29691,N_29060,N_29138);
nand U29692 (N_29692,N_28853,N_28997);
nor U29693 (N_29693,N_29264,N_29306);
nand U29694 (N_29694,N_29128,N_28941);
or U29695 (N_29695,N_29133,N_29064);
and U29696 (N_29696,N_29331,N_28987);
nand U29697 (N_29697,N_28963,N_29071);
nor U29698 (N_29698,N_29249,N_29062);
nor U29699 (N_29699,N_28904,N_29072);
nor U29700 (N_29700,N_29144,N_29113);
and U29701 (N_29701,N_29237,N_29170);
nand U29702 (N_29702,N_28936,N_29343);
xor U29703 (N_29703,N_29257,N_29020);
or U29704 (N_29704,N_28934,N_29366);
or U29705 (N_29705,N_29077,N_28932);
and U29706 (N_29706,N_29186,N_29368);
nor U29707 (N_29707,N_29158,N_29234);
and U29708 (N_29708,N_28939,N_29023);
and U29709 (N_29709,N_28895,N_28814);
nor U29710 (N_29710,N_29173,N_28951);
nand U29711 (N_29711,N_28897,N_29096);
and U29712 (N_29712,N_29168,N_29053);
nand U29713 (N_29713,N_29059,N_29146);
or U29714 (N_29714,N_29397,N_29323);
nand U29715 (N_29715,N_28842,N_28980);
and U29716 (N_29716,N_28946,N_29178);
nor U29717 (N_29717,N_29200,N_29360);
nor U29718 (N_29718,N_28830,N_29362);
nor U29719 (N_29719,N_29323,N_29147);
or U29720 (N_29720,N_29323,N_29064);
and U29721 (N_29721,N_29082,N_29241);
and U29722 (N_29722,N_29329,N_28912);
or U29723 (N_29723,N_29017,N_29214);
and U29724 (N_29724,N_28805,N_29125);
nor U29725 (N_29725,N_28963,N_28827);
nand U29726 (N_29726,N_28859,N_29054);
nor U29727 (N_29727,N_28898,N_29202);
nor U29728 (N_29728,N_29178,N_28975);
nand U29729 (N_29729,N_29097,N_29265);
and U29730 (N_29730,N_29132,N_29271);
nor U29731 (N_29731,N_29247,N_28976);
and U29732 (N_29732,N_28902,N_28815);
and U29733 (N_29733,N_28897,N_29334);
nor U29734 (N_29734,N_29244,N_29399);
nand U29735 (N_29735,N_29097,N_29111);
or U29736 (N_29736,N_29289,N_28999);
nand U29737 (N_29737,N_28924,N_29106);
and U29738 (N_29738,N_29106,N_29086);
nand U29739 (N_29739,N_29260,N_29224);
nand U29740 (N_29740,N_29099,N_29349);
or U29741 (N_29741,N_29194,N_28946);
and U29742 (N_29742,N_29348,N_28908);
xor U29743 (N_29743,N_28862,N_29218);
nor U29744 (N_29744,N_29110,N_28972);
nor U29745 (N_29745,N_29212,N_29023);
nand U29746 (N_29746,N_28824,N_28818);
nor U29747 (N_29747,N_29383,N_28987);
and U29748 (N_29748,N_29190,N_29257);
nor U29749 (N_29749,N_28904,N_29246);
or U29750 (N_29750,N_29391,N_29267);
nor U29751 (N_29751,N_29284,N_29049);
nor U29752 (N_29752,N_29178,N_28923);
or U29753 (N_29753,N_28900,N_29315);
nand U29754 (N_29754,N_29370,N_29107);
nand U29755 (N_29755,N_29151,N_29035);
nand U29756 (N_29756,N_28819,N_28821);
or U29757 (N_29757,N_28862,N_29191);
and U29758 (N_29758,N_29227,N_29095);
and U29759 (N_29759,N_29194,N_29025);
xor U29760 (N_29760,N_29248,N_28912);
nand U29761 (N_29761,N_29320,N_28811);
nor U29762 (N_29762,N_29115,N_28909);
and U29763 (N_29763,N_29016,N_29362);
nor U29764 (N_29764,N_29077,N_28956);
or U29765 (N_29765,N_29120,N_29086);
or U29766 (N_29766,N_29340,N_29394);
and U29767 (N_29767,N_28856,N_29310);
nand U29768 (N_29768,N_28937,N_29071);
and U29769 (N_29769,N_29281,N_28878);
and U29770 (N_29770,N_28825,N_29354);
nor U29771 (N_29771,N_28911,N_29315);
or U29772 (N_29772,N_29181,N_29069);
or U29773 (N_29773,N_29080,N_29089);
nor U29774 (N_29774,N_29138,N_29292);
nor U29775 (N_29775,N_29005,N_29297);
and U29776 (N_29776,N_29379,N_29244);
nor U29777 (N_29777,N_28928,N_29161);
and U29778 (N_29778,N_29155,N_29196);
and U29779 (N_29779,N_28856,N_28883);
and U29780 (N_29780,N_29395,N_29207);
nand U29781 (N_29781,N_29064,N_29060);
or U29782 (N_29782,N_29096,N_28940);
and U29783 (N_29783,N_29143,N_28978);
or U29784 (N_29784,N_28863,N_29036);
nor U29785 (N_29785,N_29070,N_28862);
or U29786 (N_29786,N_28833,N_28984);
and U29787 (N_29787,N_28985,N_29308);
nand U29788 (N_29788,N_29122,N_28938);
nand U29789 (N_29789,N_28963,N_29232);
nor U29790 (N_29790,N_28959,N_29346);
or U29791 (N_29791,N_29383,N_28904);
or U29792 (N_29792,N_28851,N_29354);
or U29793 (N_29793,N_28898,N_28867);
nor U29794 (N_29794,N_29136,N_29013);
nor U29795 (N_29795,N_28837,N_29024);
nand U29796 (N_29796,N_29255,N_28859);
nand U29797 (N_29797,N_28826,N_28969);
nor U29798 (N_29798,N_29102,N_28864);
and U29799 (N_29799,N_29252,N_29320);
nor U29800 (N_29800,N_29343,N_29065);
and U29801 (N_29801,N_29046,N_28864);
nand U29802 (N_29802,N_29004,N_29325);
nand U29803 (N_29803,N_29062,N_29196);
and U29804 (N_29804,N_29004,N_29236);
xnor U29805 (N_29805,N_28839,N_29276);
nor U29806 (N_29806,N_29278,N_29290);
and U29807 (N_29807,N_29117,N_29008);
and U29808 (N_29808,N_29207,N_29224);
nor U29809 (N_29809,N_28982,N_29376);
nor U29810 (N_29810,N_29343,N_29244);
nand U29811 (N_29811,N_28889,N_29231);
and U29812 (N_29812,N_29110,N_29301);
nand U29813 (N_29813,N_29054,N_29115);
nor U29814 (N_29814,N_29320,N_28831);
or U29815 (N_29815,N_29181,N_28937);
or U29816 (N_29816,N_29078,N_29182);
nor U29817 (N_29817,N_28810,N_28829);
or U29818 (N_29818,N_29211,N_29079);
nand U29819 (N_29819,N_28802,N_29314);
nor U29820 (N_29820,N_29344,N_29100);
and U29821 (N_29821,N_28951,N_29396);
or U29822 (N_29822,N_29045,N_29206);
and U29823 (N_29823,N_29352,N_29323);
nand U29824 (N_29824,N_28932,N_28915);
or U29825 (N_29825,N_29317,N_29098);
and U29826 (N_29826,N_28859,N_29029);
nor U29827 (N_29827,N_28960,N_29271);
nand U29828 (N_29828,N_29047,N_28888);
nand U29829 (N_29829,N_29145,N_28831);
or U29830 (N_29830,N_29040,N_29202);
nor U29831 (N_29831,N_29253,N_28936);
nand U29832 (N_29832,N_28971,N_28960);
or U29833 (N_29833,N_29127,N_29267);
and U29834 (N_29834,N_28868,N_29305);
and U29835 (N_29835,N_28883,N_28880);
and U29836 (N_29836,N_29253,N_28900);
xnor U29837 (N_29837,N_29182,N_28987);
or U29838 (N_29838,N_28976,N_29264);
and U29839 (N_29839,N_29136,N_28828);
and U29840 (N_29840,N_28874,N_29121);
nand U29841 (N_29841,N_29193,N_29324);
nand U29842 (N_29842,N_29218,N_29113);
nand U29843 (N_29843,N_29079,N_29265);
nor U29844 (N_29844,N_29218,N_29159);
nand U29845 (N_29845,N_29315,N_29240);
or U29846 (N_29846,N_28931,N_28987);
nand U29847 (N_29847,N_29334,N_29096);
nand U29848 (N_29848,N_29286,N_28994);
nor U29849 (N_29849,N_29298,N_28837);
nor U29850 (N_29850,N_29390,N_29283);
or U29851 (N_29851,N_29011,N_29273);
or U29852 (N_29852,N_29210,N_29330);
nand U29853 (N_29853,N_29348,N_29152);
nor U29854 (N_29854,N_29287,N_28968);
or U29855 (N_29855,N_29132,N_29151);
nand U29856 (N_29856,N_29238,N_28859);
nor U29857 (N_29857,N_28916,N_29148);
and U29858 (N_29858,N_29188,N_29181);
nand U29859 (N_29859,N_29103,N_29285);
nand U29860 (N_29860,N_28823,N_29099);
and U29861 (N_29861,N_29360,N_28829);
nor U29862 (N_29862,N_29041,N_28989);
and U29863 (N_29863,N_28910,N_28906);
or U29864 (N_29864,N_29018,N_29243);
or U29865 (N_29865,N_29365,N_29093);
xnor U29866 (N_29866,N_29038,N_29179);
and U29867 (N_29867,N_28865,N_29346);
and U29868 (N_29868,N_29014,N_29182);
nand U29869 (N_29869,N_28934,N_28980);
nor U29870 (N_29870,N_28977,N_29317);
nand U29871 (N_29871,N_29369,N_28858);
nand U29872 (N_29872,N_29361,N_28827);
nand U29873 (N_29873,N_28835,N_28824);
nor U29874 (N_29874,N_29160,N_29375);
nand U29875 (N_29875,N_28964,N_28885);
nor U29876 (N_29876,N_29309,N_29304);
and U29877 (N_29877,N_29073,N_29159);
nor U29878 (N_29878,N_28895,N_28841);
nor U29879 (N_29879,N_29252,N_29106);
or U29880 (N_29880,N_29392,N_28971);
and U29881 (N_29881,N_28956,N_29287);
nor U29882 (N_29882,N_29216,N_29398);
xor U29883 (N_29883,N_29356,N_29361);
or U29884 (N_29884,N_28931,N_29391);
or U29885 (N_29885,N_28809,N_28958);
nor U29886 (N_29886,N_28969,N_29137);
or U29887 (N_29887,N_29096,N_29232);
nand U29888 (N_29888,N_29256,N_28812);
nand U29889 (N_29889,N_29198,N_29179);
nand U29890 (N_29890,N_29358,N_29365);
nand U29891 (N_29891,N_28844,N_29273);
nand U29892 (N_29892,N_29116,N_29110);
and U29893 (N_29893,N_29050,N_29316);
and U29894 (N_29894,N_29393,N_29395);
or U29895 (N_29895,N_28930,N_29140);
and U29896 (N_29896,N_29097,N_28890);
or U29897 (N_29897,N_28997,N_29294);
or U29898 (N_29898,N_29029,N_28922);
nor U29899 (N_29899,N_28829,N_29333);
xor U29900 (N_29900,N_29100,N_28869);
xnor U29901 (N_29901,N_28987,N_28988);
or U29902 (N_29902,N_29316,N_28980);
nand U29903 (N_29903,N_29357,N_28803);
nand U29904 (N_29904,N_29341,N_29325);
or U29905 (N_29905,N_28921,N_28922);
nand U29906 (N_29906,N_28848,N_28872);
and U29907 (N_29907,N_28856,N_28898);
and U29908 (N_29908,N_29297,N_28815);
nand U29909 (N_29909,N_28955,N_29321);
nor U29910 (N_29910,N_28874,N_28905);
and U29911 (N_29911,N_29153,N_28913);
and U29912 (N_29912,N_29208,N_29357);
or U29913 (N_29913,N_29065,N_29053);
and U29914 (N_29914,N_29110,N_28994);
xor U29915 (N_29915,N_29262,N_28862);
nor U29916 (N_29916,N_29007,N_29106);
or U29917 (N_29917,N_29242,N_29360);
or U29918 (N_29918,N_29206,N_29177);
or U29919 (N_29919,N_29188,N_29019);
nor U29920 (N_29920,N_29304,N_28837);
or U29921 (N_29921,N_28986,N_29284);
and U29922 (N_29922,N_28968,N_29197);
and U29923 (N_29923,N_29320,N_29279);
xor U29924 (N_29924,N_29001,N_29356);
xor U29925 (N_29925,N_28855,N_29299);
nor U29926 (N_29926,N_29169,N_29047);
nor U29927 (N_29927,N_29096,N_28888);
and U29928 (N_29928,N_28845,N_29174);
and U29929 (N_29929,N_29221,N_29127);
or U29930 (N_29930,N_28930,N_29017);
nand U29931 (N_29931,N_28907,N_28869);
nand U29932 (N_29932,N_28835,N_29329);
or U29933 (N_29933,N_28872,N_28843);
or U29934 (N_29934,N_29274,N_28956);
or U29935 (N_29935,N_29272,N_28987);
and U29936 (N_29936,N_28925,N_29004);
nor U29937 (N_29937,N_29178,N_29132);
nand U29938 (N_29938,N_29028,N_29076);
and U29939 (N_29939,N_29101,N_29068);
or U29940 (N_29940,N_29338,N_29222);
or U29941 (N_29941,N_28830,N_29300);
or U29942 (N_29942,N_29297,N_29077);
nand U29943 (N_29943,N_29241,N_28878);
and U29944 (N_29944,N_29351,N_29287);
nand U29945 (N_29945,N_29192,N_29340);
nor U29946 (N_29946,N_29191,N_29232);
nor U29947 (N_29947,N_29262,N_29137);
and U29948 (N_29948,N_29370,N_28857);
nand U29949 (N_29949,N_29329,N_29177);
or U29950 (N_29950,N_29252,N_29243);
and U29951 (N_29951,N_28867,N_28853);
or U29952 (N_29952,N_28974,N_28949);
xnor U29953 (N_29953,N_29390,N_28980);
or U29954 (N_29954,N_28943,N_28937);
or U29955 (N_29955,N_29137,N_28945);
or U29956 (N_29956,N_28963,N_29195);
and U29957 (N_29957,N_28835,N_29058);
nor U29958 (N_29958,N_29276,N_29043);
nand U29959 (N_29959,N_29128,N_29137);
xnor U29960 (N_29960,N_29238,N_29133);
and U29961 (N_29961,N_29315,N_28993);
or U29962 (N_29962,N_29371,N_29245);
and U29963 (N_29963,N_29151,N_29101);
and U29964 (N_29964,N_29257,N_29181);
or U29965 (N_29965,N_29299,N_29343);
nand U29966 (N_29966,N_29153,N_28928);
nor U29967 (N_29967,N_29363,N_28877);
or U29968 (N_29968,N_28993,N_29236);
and U29969 (N_29969,N_29222,N_29280);
and U29970 (N_29970,N_28970,N_29216);
and U29971 (N_29971,N_28817,N_29022);
or U29972 (N_29972,N_28928,N_29174);
nand U29973 (N_29973,N_29232,N_28951);
nor U29974 (N_29974,N_29255,N_29361);
nor U29975 (N_29975,N_28808,N_28835);
or U29976 (N_29976,N_29227,N_28989);
nor U29977 (N_29977,N_29096,N_29269);
or U29978 (N_29978,N_29334,N_29263);
nor U29979 (N_29979,N_28931,N_29239);
nand U29980 (N_29980,N_29027,N_29261);
or U29981 (N_29981,N_29323,N_29026);
or U29982 (N_29982,N_29140,N_29383);
or U29983 (N_29983,N_29240,N_29057);
nand U29984 (N_29984,N_28901,N_29195);
nor U29985 (N_29985,N_28894,N_28982);
nor U29986 (N_29986,N_29344,N_29033);
or U29987 (N_29987,N_29047,N_28979);
and U29988 (N_29988,N_28882,N_29203);
nor U29989 (N_29989,N_29256,N_28973);
and U29990 (N_29990,N_29164,N_29330);
nand U29991 (N_29991,N_28997,N_29214);
or U29992 (N_29992,N_29270,N_29321);
nor U29993 (N_29993,N_29188,N_28948);
nor U29994 (N_29994,N_29357,N_29301);
nor U29995 (N_29995,N_29241,N_29266);
nor U29996 (N_29996,N_29348,N_28955);
xor U29997 (N_29997,N_29191,N_29027);
nor U29998 (N_29998,N_29399,N_29395);
or U29999 (N_29999,N_29098,N_28971);
and UO_0 (O_0,N_29784,N_29756);
or UO_1 (O_1,N_29429,N_29864);
and UO_2 (O_2,N_29506,N_29910);
xnor UO_3 (O_3,N_29854,N_29510);
nor UO_4 (O_4,N_29764,N_29745);
and UO_5 (O_5,N_29741,N_29759);
or UO_6 (O_6,N_29433,N_29403);
and UO_7 (O_7,N_29462,N_29900);
nor UO_8 (O_8,N_29488,N_29856);
nand UO_9 (O_9,N_29762,N_29877);
nand UO_10 (O_10,N_29995,N_29678);
or UO_11 (O_11,N_29752,N_29642);
nand UO_12 (O_12,N_29711,N_29987);
or UO_13 (O_13,N_29643,N_29931);
and UO_14 (O_14,N_29773,N_29966);
nor UO_15 (O_15,N_29958,N_29695);
nand UO_16 (O_16,N_29683,N_29672);
or UO_17 (O_17,N_29645,N_29454);
nor UO_18 (O_18,N_29973,N_29679);
or UO_19 (O_19,N_29845,N_29412);
nor UO_20 (O_20,N_29559,N_29545);
or UO_21 (O_21,N_29727,N_29967);
nand UO_22 (O_22,N_29582,N_29828);
nor UO_23 (O_23,N_29460,N_29792);
or UO_24 (O_24,N_29786,N_29539);
nand UO_25 (O_25,N_29436,N_29708);
or UO_26 (O_26,N_29541,N_29937);
nand UO_27 (O_27,N_29451,N_29810);
nor UO_28 (O_28,N_29661,N_29951);
or UO_29 (O_29,N_29915,N_29467);
xnor UO_30 (O_30,N_29530,N_29984);
or UO_31 (O_31,N_29461,N_29674);
or UO_32 (O_32,N_29558,N_29485);
nor UO_33 (O_33,N_29639,N_29847);
nand UO_34 (O_34,N_29564,N_29840);
nor UO_35 (O_35,N_29832,N_29423);
or UO_36 (O_36,N_29596,N_29556);
or UO_37 (O_37,N_29599,N_29668);
or UO_38 (O_38,N_29540,N_29621);
nand UO_39 (O_39,N_29664,N_29749);
nand UO_40 (O_40,N_29746,N_29822);
and UO_41 (O_41,N_29554,N_29945);
nor UO_42 (O_42,N_29647,N_29535);
and UO_43 (O_43,N_29938,N_29990);
nor UO_44 (O_44,N_29422,N_29921);
or UO_45 (O_45,N_29791,N_29870);
nor UO_46 (O_46,N_29899,N_29496);
and UO_47 (O_47,N_29775,N_29842);
nor UO_48 (O_48,N_29761,N_29821);
or UO_49 (O_49,N_29862,N_29841);
nor UO_50 (O_50,N_29766,N_29774);
nor UO_51 (O_51,N_29769,N_29884);
and UO_52 (O_52,N_29763,N_29489);
and UO_53 (O_53,N_29503,N_29501);
xnor UO_54 (O_54,N_29972,N_29863);
and UO_55 (O_55,N_29872,N_29594);
nor UO_56 (O_56,N_29930,N_29513);
nand UO_57 (O_57,N_29728,N_29913);
or UO_58 (O_58,N_29612,N_29902);
and UO_59 (O_59,N_29524,N_29646);
nor UO_60 (O_60,N_29609,N_29666);
xor UO_61 (O_61,N_29585,N_29904);
and UO_62 (O_62,N_29498,N_29908);
and UO_63 (O_63,N_29450,N_29464);
nand UO_64 (O_64,N_29969,N_29520);
xor UO_65 (O_65,N_29698,N_29697);
and UO_66 (O_66,N_29502,N_29799);
or UO_67 (O_67,N_29754,N_29421);
nand UO_68 (O_68,N_29411,N_29970);
or UO_69 (O_69,N_29947,N_29889);
and UO_70 (O_70,N_29660,N_29523);
or UO_71 (O_71,N_29684,N_29569);
and UO_72 (O_72,N_29525,N_29481);
or UO_73 (O_73,N_29509,N_29744);
nand UO_74 (O_74,N_29576,N_29444);
or UO_75 (O_75,N_29719,N_29875);
or UO_76 (O_76,N_29878,N_29446);
and UO_77 (O_77,N_29976,N_29750);
xor UO_78 (O_78,N_29805,N_29891);
or UO_79 (O_79,N_29824,N_29692);
nand UO_80 (O_80,N_29562,N_29855);
nor UO_81 (O_81,N_29567,N_29964);
nor UO_82 (O_82,N_29626,N_29575);
nor UO_83 (O_83,N_29430,N_29456);
nand UO_84 (O_84,N_29867,N_29514);
or UO_85 (O_85,N_29613,N_29515);
nor UO_86 (O_86,N_29640,N_29425);
and UO_87 (O_87,N_29492,N_29748);
nand UO_88 (O_88,N_29482,N_29505);
nor UO_89 (O_89,N_29998,N_29797);
nand UO_90 (O_90,N_29507,N_29993);
nand UO_91 (O_91,N_29572,N_29529);
and UO_92 (O_92,N_29691,N_29800);
and UO_93 (O_93,N_29758,N_29948);
or UO_94 (O_94,N_29416,N_29755);
and UO_95 (O_95,N_29406,N_29475);
nand UO_96 (O_96,N_29839,N_29893);
nand UO_97 (O_97,N_29537,N_29979);
nor UO_98 (O_98,N_29605,N_29504);
or UO_99 (O_99,N_29953,N_29455);
nor UO_100 (O_100,N_29882,N_29965);
nor UO_101 (O_101,N_29850,N_29952);
nor UO_102 (O_102,N_29490,N_29742);
and UO_103 (O_103,N_29722,N_29592);
nor UO_104 (O_104,N_29486,N_29570);
nor UO_105 (O_105,N_29787,N_29770);
or UO_106 (O_106,N_29608,N_29971);
and UO_107 (O_107,N_29439,N_29637);
nor UO_108 (O_108,N_29852,N_29549);
or UO_109 (O_109,N_29419,N_29468);
and UO_110 (O_110,N_29932,N_29941);
and UO_111 (O_111,N_29400,N_29868);
or UO_112 (O_112,N_29782,N_29603);
and UO_113 (O_113,N_29794,N_29417);
nand UO_114 (O_114,N_29988,N_29413);
or UO_115 (O_115,N_29729,N_29895);
nand UO_116 (O_116,N_29779,N_29473);
xnor UO_117 (O_117,N_29956,N_29491);
and UO_118 (O_118,N_29887,N_29954);
nor UO_119 (O_119,N_29886,N_29543);
nand UO_120 (O_120,N_29624,N_29981);
nand UO_121 (O_121,N_29614,N_29630);
or UO_122 (O_122,N_29793,N_29441);
or UO_123 (O_123,N_29838,N_29577);
nand UO_124 (O_124,N_29844,N_29894);
or UO_125 (O_125,N_29829,N_29607);
nand UO_126 (O_126,N_29696,N_29890);
nand UO_127 (O_127,N_29590,N_29431);
nor UO_128 (O_128,N_29574,N_29531);
nand UO_129 (O_129,N_29669,N_29789);
nor UO_130 (O_130,N_29714,N_29978);
or UO_131 (O_131,N_29848,N_29866);
or UO_132 (O_132,N_29655,N_29943);
or UO_133 (O_133,N_29682,N_29494);
and UO_134 (O_134,N_29709,N_29720);
nor UO_135 (O_135,N_29452,N_29686);
or UO_136 (O_136,N_29476,N_29536);
nand UO_137 (O_137,N_29670,N_29768);
nor UO_138 (O_138,N_29765,N_29725);
and UO_139 (O_139,N_29665,N_29896);
nor UO_140 (O_140,N_29751,N_29857);
or UO_141 (O_141,N_29659,N_29408);
nor UO_142 (O_142,N_29469,N_29817);
or UO_143 (O_143,N_29477,N_29449);
nor UO_144 (O_144,N_29478,N_29808);
or UO_145 (O_145,N_29772,N_29542);
nand UO_146 (O_146,N_29631,N_29892);
nor UO_147 (O_147,N_29432,N_29906);
or UO_148 (O_148,N_29658,N_29671);
nand UO_149 (O_149,N_29493,N_29813);
nor UO_150 (O_150,N_29706,N_29690);
nand UO_151 (O_151,N_29633,N_29760);
and UO_152 (O_152,N_29579,N_29985);
xnor UO_153 (O_153,N_29737,N_29833);
and UO_154 (O_154,N_29560,N_29919);
and UO_155 (O_155,N_29825,N_29940);
nor UO_156 (O_156,N_29726,N_29804);
nor UO_157 (O_157,N_29625,N_29905);
or UO_158 (O_158,N_29410,N_29986);
and UO_159 (O_159,N_29939,N_29914);
and UO_160 (O_160,N_29500,N_29834);
nor UO_161 (O_161,N_29815,N_29611);
nand UO_162 (O_162,N_29546,N_29928);
nor UO_163 (O_163,N_29803,N_29435);
nor UO_164 (O_164,N_29521,N_29566);
xnor UO_165 (O_165,N_29635,N_29694);
nand UO_166 (O_166,N_29801,N_29946);
or UO_167 (O_167,N_29718,N_29811);
and UO_168 (O_168,N_29909,N_29814);
nor UO_169 (O_169,N_29480,N_29533);
or UO_170 (O_170,N_29641,N_29802);
nor UO_171 (O_171,N_29920,N_29616);
or UO_172 (O_172,N_29740,N_29831);
nand UO_173 (O_173,N_29827,N_29547);
nor UO_174 (O_174,N_29903,N_29883);
and UO_175 (O_175,N_29517,N_29795);
or UO_176 (O_176,N_29881,N_29702);
or UO_177 (O_177,N_29897,N_29653);
nor UO_178 (O_178,N_29508,N_29519);
nand UO_179 (O_179,N_29463,N_29552);
nand UO_180 (O_180,N_29876,N_29734);
and UO_181 (O_181,N_29420,N_29681);
nand UO_182 (O_182,N_29442,N_29618);
nand UO_183 (O_183,N_29458,N_29918);
nand UO_184 (O_184,N_29716,N_29898);
or UO_185 (O_185,N_29780,N_29944);
or UO_186 (O_186,N_29601,N_29409);
nor UO_187 (O_187,N_29623,N_29959);
nand UO_188 (O_188,N_29654,N_29414);
and UO_189 (O_189,N_29602,N_29550);
and UO_190 (O_190,N_29604,N_29544);
and UO_191 (O_191,N_29471,N_29551);
xor UO_192 (O_192,N_29942,N_29443);
nand UO_193 (O_193,N_29415,N_29923);
and UO_194 (O_194,N_29687,N_29688);
nor UO_195 (O_195,N_29961,N_29627);
nand UO_196 (O_196,N_29497,N_29648);
nand UO_197 (O_197,N_29700,N_29999);
and UO_198 (O_198,N_29600,N_29879);
nand UO_199 (O_199,N_29578,N_29721);
and UO_200 (O_200,N_29924,N_29538);
or UO_201 (O_201,N_29629,N_29484);
and UO_202 (O_202,N_29796,N_29401);
nand UO_203 (O_203,N_29790,N_29816);
nand UO_204 (O_204,N_29619,N_29968);
and UO_205 (O_205,N_29565,N_29487);
nor UO_206 (O_206,N_29771,N_29818);
and UO_207 (O_207,N_29632,N_29901);
or UO_208 (O_208,N_29717,N_29781);
nand UO_209 (O_209,N_29622,N_29597);
nand UO_210 (O_210,N_29593,N_29997);
or UO_211 (O_211,N_29962,N_29853);
nor UO_212 (O_212,N_29738,N_29526);
and UO_213 (O_213,N_29584,N_29732);
or UO_214 (O_214,N_29823,N_29858);
and UO_215 (O_215,N_29583,N_29638);
nand UO_216 (O_216,N_29836,N_29936);
nor UO_217 (O_217,N_29483,N_29826);
or UO_218 (O_218,N_29849,N_29982);
and UO_219 (O_219,N_29499,N_29662);
or UO_220 (O_220,N_29511,N_29677);
or UO_221 (O_221,N_29447,N_29437);
nor UO_222 (O_222,N_29426,N_29820);
nand UO_223 (O_223,N_29405,N_29991);
nand UO_224 (O_224,N_29812,N_29907);
or UO_225 (O_225,N_29925,N_29470);
nand UO_226 (O_226,N_29620,N_29950);
or UO_227 (O_227,N_29712,N_29534);
nor UO_228 (O_228,N_29563,N_29516);
nand UO_229 (O_229,N_29438,N_29929);
nand UO_230 (O_230,N_29865,N_29587);
xor UO_231 (O_231,N_29788,N_29689);
or UO_232 (O_232,N_29860,N_29707);
or UO_233 (O_233,N_29873,N_29685);
or UO_234 (O_234,N_29739,N_29992);
nand UO_235 (O_235,N_29819,N_29553);
and UO_236 (O_236,N_29977,N_29595);
and UO_237 (O_237,N_29957,N_29851);
and UO_238 (O_238,N_29644,N_29747);
nand UO_239 (O_239,N_29743,N_29778);
and UO_240 (O_240,N_29424,N_29404);
nor UO_241 (O_241,N_29581,N_29636);
and UO_242 (O_242,N_29843,N_29675);
and UO_243 (O_243,N_29809,N_29753);
or UO_244 (O_244,N_29888,N_29912);
and UO_245 (O_245,N_29974,N_29652);
and UO_246 (O_246,N_29407,N_29713);
and UO_247 (O_247,N_29960,N_29785);
and UO_248 (O_248,N_29846,N_29428);
nand UO_249 (O_249,N_29798,N_29680);
or UO_250 (O_250,N_29548,N_29980);
nor UO_251 (O_251,N_29715,N_29457);
nand UO_252 (O_252,N_29983,N_29434);
or UO_253 (O_253,N_29479,N_29649);
or UO_254 (O_254,N_29731,N_29704);
and UO_255 (O_255,N_29927,N_29736);
nor UO_256 (O_256,N_29634,N_29911);
or UO_257 (O_257,N_29589,N_29757);
nor UO_258 (O_258,N_29586,N_29657);
nor UO_259 (O_259,N_29591,N_29573);
nand UO_260 (O_260,N_29518,N_29474);
xnor UO_261 (O_261,N_29667,N_29830);
nand UO_262 (O_262,N_29532,N_29733);
nand UO_263 (O_263,N_29459,N_29528);
nor UO_264 (O_264,N_29628,N_29427);
and UO_265 (O_265,N_29874,N_29861);
nand UO_266 (O_266,N_29933,N_29580);
nand UO_267 (O_267,N_29651,N_29701);
and UO_268 (O_268,N_29955,N_29693);
or UO_269 (O_269,N_29767,N_29935);
or UO_270 (O_270,N_29880,N_29994);
and UO_271 (O_271,N_29656,N_29512);
or UO_272 (O_272,N_29710,N_29522);
or UO_273 (O_273,N_29465,N_29663);
nor UO_274 (O_274,N_29588,N_29871);
and UO_275 (O_275,N_29617,N_29466);
nand UO_276 (O_276,N_29723,N_29571);
or UO_277 (O_277,N_29561,N_29440);
nor UO_278 (O_278,N_29598,N_29934);
and UO_279 (O_279,N_29673,N_29777);
nor UO_280 (O_280,N_29869,N_29926);
and UO_281 (O_281,N_29807,N_29859);
nor UO_282 (O_282,N_29735,N_29922);
nand UO_283 (O_283,N_29650,N_29448);
nand UO_284 (O_284,N_29402,N_29837);
nand UO_285 (O_285,N_29949,N_29835);
nor UO_286 (O_286,N_29557,N_29676);
nor UO_287 (O_287,N_29917,N_29776);
nor UO_288 (O_288,N_29472,N_29527);
and UO_289 (O_289,N_29975,N_29730);
nor UO_290 (O_290,N_29989,N_29606);
and UO_291 (O_291,N_29724,N_29996);
or UO_292 (O_292,N_29555,N_29916);
or UO_293 (O_293,N_29453,N_29963);
nor UO_294 (O_294,N_29806,N_29705);
or UO_295 (O_295,N_29568,N_29610);
and UO_296 (O_296,N_29783,N_29495);
nor UO_297 (O_297,N_29703,N_29418);
nor UO_298 (O_298,N_29885,N_29699);
nor UO_299 (O_299,N_29445,N_29615);
nand UO_300 (O_300,N_29980,N_29465);
and UO_301 (O_301,N_29410,N_29629);
nor UO_302 (O_302,N_29589,N_29900);
or UO_303 (O_303,N_29485,N_29529);
nor UO_304 (O_304,N_29946,N_29906);
or UO_305 (O_305,N_29827,N_29759);
and UO_306 (O_306,N_29908,N_29625);
and UO_307 (O_307,N_29501,N_29456);
nor UO_308 (O_308,N_29468,N_29671);
and UO_309 (O_309,N_29878,N_29517);
nand UO_310 (O_310,N_29599,N_29486);
nor UO_311 (O_311,N_29524,N_29847);
nand UO_312 (O_312,N_29554,N_29542);
and UO_313 (O_313,N_29472,N_29883);
nor UO_314 (O_314,N_29686,N_29438);
and UO_315 (O_315,N_29595,N_29474);
or UO_316 (O_316,N_29534,N_29513);
nor UO_317 (O_317,N_29801,N_29513);
and UO_318 (O_318,N_29494,N_29782);
and UO_319 (O_319,N_29999,N_29510);
nor UO_320 (O_320,N_29995,N_29471);
or UO_321 (O_321,N_29583,N_29893);
or UO_322 (O_322,N_29422,N_29439);
nor UO_323 (O_323,N_29660,N_29431);
or UO_324 (O_324,N_29888,N_29450);
nand UO_325 (O_325,N_29812,N_29966);
and UO_326 (O_326,N_29744,N_29479);
nand UO_327 (O_327,N_29834,N_29857);
or UO_328 (O_328,N_29884,N_29411);
nor UO_329 (O_329,N_29837,N_29548);
or UO_330 (O_330,N_29722,N_29938);
nor UO_331 (O_331,N_29418,N_29925);
and UO_332 (O_332,N_29733,N_29935);
and UO_333 (O_333,N_29893,N_29745);
or UO_334 (O_334,N_29998,N_29484);
nand UO_335 (O_335,N_29555,N_29518);
or UO_336 (O_336,N_29559,N_29952);
nand UO_337 (O_337,N_29715,N_29427);
nand UO_338 (O_338,N_29863,N_29747);
nor UO_339 (O_339,N_29663,N_29519);
nor UO_340 (O_340,N_29782,N_29929);
and UO_341 (O_341,N_29822,N_29673);
or UO_342 (O_342,N_29660,N_29510);
and UO_343 (O_343,N_29746,N_29995);
nor UO_344 (O_344,N_29655,N_29644);
or UO_345 (O_345,N_29857,N_29519);
nand UO_346 (O_346,N_29664,N_29650);
and UO_347 (O_347,N_29772,N_29460);
and UO_348 (O_348,N_29683,N_29843);
and UO_349 (O_349,N_29718,N_29976);
nor UO_350 (O_350,N_29814,N_29521);
and UO_351 (O_351,N_29645,N_29561);
or UO_352 (O_352,N_29976,N_29927);
nand UO_353 (O_353,N_29760,N_29702);
and UO_354 (O_354,N_29929,N_29541);
or UO_355 (O_355,N_29796,N_29893);
xnor UO_356 (O_356,N_29775,N_29494);
nand UO_357 (O_357,N_29695,N_29736);
nor UO_358 (O_358,N_29513,N_29403);
or UO_359 (O_359,N_29886,N_29475);
or UO_360 (O_360,N_29424,N_29416);
or UO_361 (O_361,N_29892,N_29594);
nor UO_362 (O_362,N_29874,N_29891);
nand UO_363 (O_363,N_29467,N_29622);
nor UO_364 (O_364,N_29911,N_29645);
nor UO_365 (O_365,N_29575,N_29739);
and UO_366 (O_366,N_29960,N_29578);
and UO_367 (O_367,N_29422,N_29401);
nand UO_368 (O_368,N_29686,N_29458);
and UO_369 (O_369,N_29699,N_29579);
and UO_370 (O_370,N_29745,N_29809);
or UO_371 (O_371,N_29443,N_29454);
and UO_372 (O_372,N_29707,N_29628);
nor UO_373 (O_373,N_29448,N_29829);
nor UO_374 (O_374,N_29950,N_29949);
nand UO_375 (O_375,N_29950,N_29781);
or UO_376 (O_376,N_29787,N_29913);
nor UO_377 (O_377,N_29484,N_29543);
nand UO_378 (O_378,N_29404,N_29476);
nor UO_379 (O_379,N_29992,N_29708);
nor UO_380 (O_380,N_29965,N_29906);
nor UO_381 (O_381,N_29868,N_29808);
or UO_382 (O_382,N_29601,N_29625);
nand UO_383 (O_383,N_29940,N_29689);
nand UO_384 (O_384,N_29461,N_29592);
nand UO_385 (O_385,N_29658,N_29475);
nand UO_386 (O_386,N_29791,N_29690);
and UO_387 (O_387,N_29492,N_29551);
nor UO_388 (O_388,N_29719,N_29557);
nor UO_389 (O_389,N_29847,N_29990);
nor UO_390 (O_390,N_29561,N_29901);
nor UO_391 (O_391,N_29928,N_29400);
nor UO_392 (O_392,N_29901,N_29494);
nand UO_393 (O_393,N_29481,N_29934);
or UO_394 (O_394,N_29831,N_29589);
or UO_395 (O_395,N_29998,N_29651);
nor UO_396 (O_396,N_29639,N_29938);
nor UO_397 (O_397,N_29607,N_29759);
xor UO_398 (O_398,N_29879,N_29581);
nand UO_399 (O_399,N_29435,N_29945);
or UO_400 (O_400,N_29777,N_29608);
or UO_401 (O_401,N_29744,N_29652);
or UO_402 (O_402,N_29443,N_29552);
nor UO_403 (O_403,N_29901,N_29660);
and UO_404 (O_404,N_29750,N_29638);
xnor UO_405 (O_405,N_29612,N_29952);
and UO_406 (O_406,N_29544,N_29714);
and UO_407 (O_407,N_29855,N_29581);
and UO_408 (O_408,N_29675,N_29920);
nor UO_409 (O_409,N_29803,N_29484);
nand UO_410 (O_410,N_29649,N_29541);
and UO_411 (O_411,N_29890,N_29572);
nor UO_412 (O_412,N_29695,N_29716);
nand UO_413 (O_413,N_29638,N_29888);
nand UO_414 (O_414,N_29690,N_29665);
nand UO_415 (O_415,N_29578,N_29811);
and UO_416 (O_416,N_29416,N_29403);
or UO_417 (O_417,N_29540,N_29726);
nand UO_418 (O_418,N_29445,N_29588);
nor UO_419 (O_419,N_29415,N_29463);
nor UO_420 (O_420,N_29893,N_29966);
or UO_421 (O_421,N_29429,N_29572);
and UO_422 (O_422,N_29903,N_29709);
or UO_423 (O_423,N_29631,N_29697);
or UO_424 (O_424,N_29892,N_29678);
or UO_425 (O_425,N_29574,N_29565);
or UO_426 (O_426,N_29717,N_29540);
or UO_427 (O_427,N_29654,N_29715);
nand UO_428 (O_428,N_29559,N_29829);
and UO_429 (O_429,N_29406,N_29512);
or UO_430 (O_430,N_29722,N_29803);
or UO_431 (O_431,N_29575,N_29649);
and UO_432 (O_432,N_29883,N_29941);
nor UO_433 (O_433,N_29631,N_29545);
and UO_434 (O_434,N_29833,N_29956);
and UO_435 (O_435,N_29972,N_29991);
and UO_436 (O_436,N_29485,N_29817);
and UO_437 (O_437,N_29603,N_29915);
nand UO_438 (O_438,N_29544,N_29790);
nand UO_439 (O_439,N_29641,N_29435);
and UO_440 (O_440,N_29652,N_29617);
nor UO_441 (O_441,N_29928,N_29762);
or UO_442 (O_442,N_29824,N_29509);
xnor UO_443 (O_443,N_29630,N_29483);
and UO_444 (O_444,N_29957,N_29863);
or UO_445 (O_445,N_29785,N_29660);
and UO_446 (O_446,N_29611,N_29732);
or UO_447 (O_447,N_29769,N_29734);
and UO_448 (O_448,N_29711,N_29613);
or UO_449 (O_449,N_29488,N_29596);
or UO_450 (O_450,N_29688,N_29825);
nand UO_451 (O_451,N_29551,N_29445);
nand UO_452 (O_452,N_29676,N_29840);
nor UO_453 (O_453,N_29482,N_29449);
nor UO_454 (O_454,N_29439,N_29614);
or UO_455 (O_455,N_29628,N_29597);
and UO_456 (O_456,N_29824,N_29880);
and UO_457 (O_457,N_29936,N_29580);
nor UO_458 (O_458,N_29475,N_29835);
or UO_459 (O_459,N_29588,N_29510);
or UO_460 (O_460,N_29828,N_29522);
nand UO_461 (O_461,N_29753,N_29573);
nor UO_462 (O_462,N_29799,N_29487);
and UO_463 (O_463,N_29506,N_29626);
and UO_464 (O_464,N_29856,N_29514);
and UO_465 (O_465,N_29528,N_29465);
and UO_466 (O_466,N_29533,N_29951);
or UO_467 (O_467,N_29932,N_29893);
and UO_468 (O_468,N_29578,N_29843);
and UO_469 (O_469,N_29640,N_29960);
or UO_470 (O_470,N_29550,N_29875);
and UO_471 (O_471,N_29938,N_29815);
nor UO_472 (O_472,N_29464,N_29666);
nand UO_473 (O_473,N_29903,N_29835);
nor UO_474 (O_474,N_29419,N_29994);
or UO_475 (O_475,N_29733,N_29916);
nand UO_476 (O_476,N_29629,N_29716);
nand UO_477 (O_477,N_29638,N_29961);
xor UO_478 (O_478,N_29691,N_29838);
or UO_479 (O_479,N_29628,N_29567);
nor UO_480 (O_480,N_29678,N_29538);
or UO_481 (O_481,N_29618,N_29682);
or UO_482 (O_482,N_29550,N_29573);
nor UO_483 (O_483,N_29692,N_29908);
nand UO_484 (O_484,N_29547,N_29937);
or UO_485 (O_485,N_29500,N_29589);
or UO_486 (O_486,N_29991,N_29858);
nand UO_487 (O_487,N_29495,N_29679);
nor UO_488 (O_488,N_29929,N_29776);
or UO_489 (O_489,N_29552,N_29486);
or UO_490 (O_490,N_29951,N_29780);
nand UO_491 (O_491,N_29443,N_29803);
nand UO_492 (O_492,N_29937,N_29879);
and UO_493 (O_493,N_29964,N_29409);
nor UO_494 (O_494,N_29580,N_29891);
and UO_495 (O_495,N_29986,N_29872);
or UO_496 (O_496,N_29447,N_29427);
or UO_497 (O_497,N_29877,N_29495);
and UO_498 (O_498,N_29823,N_29589);
nand UO_499 (O_499,N_29794,N_29595);
and UO_500 (O_500,N_29923,N_29994);
and UO_501 (O_501,N_29708,N_29420);
or UO_502 (O_502,N_29481,N_29939);
or UO_503 (O_503,N_29871,N_29875);
or UO_504 (O_504,N_29755,N_29799);
and UO_505 (O_505,N_29899,N_29808);
nand UO_506 (O_506,N_29711,N_29708);
nor UO_507 (O_507,N_29475,N_29515);
and UO_508 (O_508,N_29530,N_29890);
nor UO_509 (O_509,N_29693,N_29629);
nor UO_510 (O_510,N_29804,N_29879);
nor UO_511 (O_511,N_29542,N_29680);
and UO_512 (O_512,N_29998,N_29868);
or UO_513 (O_513,N_29746,N_29696);
or UO_514 (O_514,N_29779,N_29994);
nor UO_515 (O_515,N_29668,N_29836);
nand UO_516 (O_516,N_29570,N_29578);
or UO_517 (O_517,N_29704,N_29541);
xnor UO_518 (O_518,N_29859,N_29410);
nor UO_519 (O_519,N_29462,N_29970);
nand UO_520 (O_520,N_29476,N_29515);
or UO_521 (O_521,N_29522,N_29922);
nor UO_522 (O_522,N_29444,N_29997);
nor UO_523 (O_523,N_29434,N_29718);
nor UO_524 (O_524,N_29551,N_29411);
or UO_525 (O_525,N_29996,N_29784);
and UO_526 (O_526,N_29872,N_29827);
nand UO_527 (O_527,N_29452,N_29699);
nor UO_528 (O_528,N_29710,N_29433);
and UO_529 (O_529,N_29891,N_29558);
xor UO_530 (O_530,N_29948,N_29462);
nand UO_531 (O_531,N_29938,N_29536);
nor UO_532 (O_532,N_29701,N_29643);
nand UO_533 (O_533,N_29671,N_29678);
and UO_534 (O_534,N_29497,N_29447);
and UO_535 (O_535,N_29541,N_29563);
or UO_536 (O_536,N_29755,N_29626);
and UO_537 (O_537,N_29640,N_29580);
or UO_538 (O_538,N_29910,N_29998);
or UO_539 (O_539,N_29798,N_29534);
nor UO_540 (O_540,N_29681,N_29404);
or UO_541 (O_541,N_29458,N_29596);
nand UO_542 (O_542,N_29443,N_29560);
nand UO_543 (O_543,N_29860,N_29563);
or UO_544 (O_544,N_29937,N_29463);
and UO_545 (O_545,N_29543,N_29889);
or UO_546 (O_546,N_29729,N_29925);
nor UO_547 (O_547,N_29904,N_29417);
nor UO_548 (O_548,N_29758,N_29897);
or UO_549 (O_549,N_29671,N_29861);
or UO_550 (O_550,N_29711,N_29949);
or UO_551 (O_551,N_29618,N_29771);
nor UO_552 (O_552,N_29854,N_29620);
nor UO_553 (O_553,N_29587,N_29682);
xor UO_554 (O_554,N_29689,N_29632);
nand UO_555 (O_555,N_29907,N_29960);
nand UO_556 (O_556,N_29687,N_29652);
or UO_557 (O_557,N_29542,N_29913);
or UO_558 (O_558,N_29722,N_29621);
nor UO_559 (O_559,N_29765,N_29593);
nor UO_560 (O_560,N_29447,N_29935);
nor UO_561 (O_561,N_29998,N_29564);
nor UO_562 (O_562,N_29913,N_29879);
nor UO_563 (O_563,N_29790,N_29796);
nand UO_564 (O_564,N_29426,N_29915);
nand UO_565 (O_565,N_29702,N_29473);
nor UO_566 (O_566,N_29719,N_29432);
nand UO_567 (O_567,N_29483,N_29773);
and UO_568 (O_568,N_29908,N_29675);
nand UO_569 (O_569,N_29965,N_29740);
and UO_570 (O_570,N_29864,N_29401);
or UO_571 (O_571,N_29913,N_29488);
and UO_572 (O_572,N_29588,N_29876);
nand UO_573 (O_573,N_29957,N_29791);
and UO_574 (O_574,N_29752,N_29958);
nor UO_575 (O_575,N_29568,N_29577);
nand UO_576 (O_576,N_29425,N_29893);
or UO_577 (O_577,N_29749,N_29640);
or UO_578 (O_578,N_29554,N_29844);
and UO_579 (O_579,N_29890,N_29702);
nand UO_580 (O_580,N_29876,N_29642);
nor UO_581 (O_581,N_29763,N_29699);
xor UO_582 (O_582,N_29480,N_29990);
and UO_583 (O_583,N_29623,N_29872);
and UO_584 (O_584,N_29849,N_29581);
and UO_585 (O_585,N_29761,N_29577);
or UO_586 (O_586,N_29942,N_29992);
or UO_587 (O_587,N_29696,N_29434);
or UO_588 (O_588,N_29749,N_29539);
nor UO_589 (O_589,N_29524,N_29891);
nand UO_590 (O_590,N_29409,N_29454);
and UO_591 (O_591,N_29653,N_29448);
and UO_592 (O_592,N_29480,N_29758);
nor UO_593 (O_593,N_29957,N_29722);
nor UO_594 (O_594,N_29410,N_29847);
nand UO_595 (O_595,N_29778,N_29458);
nor UO_596 (O_596,N_29771,N_29458);
nand UO_597 (O_597,N_29654,N_29705);
nor UO_598 (O_598,N_29717,N_29688);
and UO_599 (O_599,N_29559,N_29582);
nand UO_600 (O_600,N_29515,N_29763);
and UO_601 (O_601,N_29672,N_29522);
nor UO_602 (O_602,N_29689,N_29536);
nor UO_603 (O_603,N_29673,N_29410);
nand UO_604 (O_604,N_29779,N_29708);
xor UO_605 (O_605,N_29862,N_29693);
nand UO_606 (O_606,N_29482,N_29437);
or UO_607 (O_607,N_29731,N_29850);
or UO_608 (O_608,N_29824,N_29515);
nor UO_609 (O_609,N_29476,N_29800);
or UO_610 (O_610,N_29944,N_29949);
nand UO_611 (O_611,N_29569,N_29631);
and UO_612 (O_612,N_29903,N_29726);
nor UO_613 (O_613,N_29710,N_29606);
nor UO_614 (O_614,N_29946,N_29415);
nor UO_615 (O_615,N_29656,N_29828);
nor UO_616 (O_616,N_29474,N_29802);
or UO_617 (O_617,N_29911,N_29463);
and UO_618 (O_618,N_29457,N_29897);
and UO_619 (O_619,N_29531,N_29685);
nand UO_620 (O_620,N_29788,N_29625);
and UO_621 (O_621,N_29513,N_29445);
and UO_622 (O_622,N_29406,N_29569);
xnor UO_623 (O_623,N_29740,N_29564);
or UO_624 (O_624,N_29760,N_29552);
or UO_625 (O_625,N_29559,N_29943);
or UO_626 (O_626,N_29710,N_29769);
nor UO_627 (O_627,N_29674,N_29976);
nor UO_628 (O_628,N_29945,N_29865);
nor UO_629 (O_629,N_29747,N_29643);
nor UO_630 (O_630,N_29748,N_29683);
xor UO_631 (O_631,N_29520,N_29406);
or UO_632 (O_632,N_29797,N_29512);
nor UO_633 (O_633,N_29564,N_29539);
xor UO_634 (O_634,N_29820,N_29619);
nand UO_635 (O_635,N_29438,N_29655);
and UO_636 (O_636,N_29761,N_29766);
or UO_637 (O_637,N_29857,N_29431);
and UO_638 (O_638,N_29578,N_29895);
and UO_639 (O_639,N_29941,N_29467);
nand UO_640 (O_640,N_29566,N_29911);
and UO_641 (O_641,N_29830,N_29446);
nand UO_642 (O_642,N_29601,N_29975);
or UO_643 (O_643,N_29938,N_29580);
or UO_644 (O_644,N_29648,N_29730);
nor UO_645 (O_645,N_29415,N_29546);
nor UO_646 (O_646,N_29709,N_29576);
and UO_647 (O_647,N_29792,N_29631);
nand UO_648 (O_648,N_29532,N_29843);
nand UO_649 (O_649,N_29729,N_29514);
and UO_650 (O_650,N_29608,N_29536);
nor UO_651 (O_651,N_29959,N_29486);
nor UO_652 (O_652,N_29944,N_29808);
nand UO_653 (O_653,N_29594,N_29489);
or UO_654 (O_654,N_29440,N_29690);
nor UO_655 (O_655,N_29663,N_29718);
and UO_656 (O_656,N_29578,N_29726);
and UO_657 (O_657,N_29584,N_29662);
nand UO_658 (O_658,N_29587,N_29785);
nand UO_659 (O_659,N_29401,N_29997);
or UO_660 (O_660,N_29444,N_29564);
nor UO_661 (O_661,N_29497,N_29817);
and UO_662 (O_662,N_29932,N_29483);
xnor UO_663 (O_663,N_29678,N_29685);
nor UO_664 (O_664,N_29816,N_29758);
and UO_665 (O_665,N_29800,N_29511);
xor UO_666 (O_666,N_29618,N_29868);
nand UO_667 (O_667,N_29828,N_29497);
nand UO_668 (O_668,N_29599,N_29720);
nor UO_669 (O_669,N_29738,N_29581);
and UO_670 (O_670,N_29684,N_29841);
nor UO_671 (O_671,N_29940,N_29577);
or UO_672 (O_672,N_29495,N_29466);
or UO_673 (O_673,N_29832,N_29769);
nor UO_674 (O_674,N_29956,N_29645);
or UO_675 (O_675,N_29524,N_29589);
nand UO_676 (O_676,N_29988,N_29507);
nand UO_677 (O_677,N_29844,N_29874);
nor UO_678 (O_678,N_29452,N_29849);
and UO_679 (O_679,N_29647,N_29975);
nor UO_680 (O_680,N_29666,N_29719);
nand UO_681 (O_681,N_29894,N_29593);
and UO_682 (O_682,N_29717,N_29759);
nor UO_683 (O_683,N_29734,N_29847);
or UO_684 (O_684,N_29780,N_29994);
and UO_685 (O_685,N_29748,N_29446);
and UO_686 (O_686,N_29793,N_29934);
or UO_687 (O_687,N_29793,N_29944);
xor UO_688 (O_688,N_29686,N_29987);
nor UO_689 (O_689,N_29415,N_29695);
nand UO_690 (O_690,N_29458,N_29483);
or UO_691 (O_691,N_29979,N_29618);
nor UO_692 (O_692,N_29639,N_29727);
and UO_693 (O_693,N_29536,N_29430);
or UO_694 (O_694,N_29627,N_29897);
nor UO_695 (O_695,N_29685,N_29766);
and UO_696 (O_696,N_29528,N_29629);
nor UO_697 (O_697,N_29856,N_29795);
nor UO_698 (O_698,N_29975,N_29565);
nor UO_699 (O_699,N_29455,N_29784);
nor UO_700 (O_700,N_29971,N_29733);
and UO_701 (O_701,N_29671,N_29912);
and UO_702 (O_702,N_29981,N_29581);
nor UO_703 (O_703,N_29588,N_29490);
or UO_704 (O_704,N_29901,N_29404);
or UO_705 (O_705,N_29562,N_29649);
or UO_706 (O_706,N_29457,N_29976);
nand UO_707 (O_707,N_29551,N_29953);
nand UO_708 (O_708,N_29944,N_29604);
and UO_709 (O_709,N_29695,N_29641);
nor UO_710 (O_710,N_29464,N_29959);
nand UO_711 (O_711,N_29543,N_29743);
nand UO_712 (O_712,N_29462,N_29989);
and UO_713 (O_713,N_29906,N_29407);
nor UO_714 (O_714,N_29844,N_29776);
and UO_715 (O_715,N_29811,N_29476);
nor UO_716 (O_716,N_29568,N_29642);
nor UO_717 (O_717,N_29912,N_29507);
or UO_718 (O_718,N_29549,N_29920);
nand UO_719 (O_719,N_29791,N_29478);
or UO_720 (O_720,N_29406,N_29461);
nand UO_721 (O_721,N_29987,N_29452);
or UO_722 (O_722,N_29599,N_29690);
and UO_723 (O_723,N_29574,N_29792);
xnor UO_724 (O_724,N_29903,N_29776);
or UO_725 (O_725,N_29664,N_29727);
xnor UO_726 (O_726,N_29970,N_29415);
nor UO_727 (O_727,N_29482,N_29688);
and UO_728 (O_728,N_29424,N_29456);
nand UO_729 (O_729,N_29714,N_29606);
xnor UO_730 (O_730,N_29613,N_29701);
and UO_731 (O_731,N_29895,N_29613);
or UO_732 (O_732,N_29730,N_29800);
xor UO_733 (O_733,N_29472,N_29703);
nor UO_734 (O_734,N_29920,N_29570);
and UO_735 (O_735,N_29553,N_29563);
and UO_736 (O_736,N_29661,N_29578);
nand UO_737 (O_737,N_29491,N_29639);
nor UO_738 (O_738,N_29630,N_29861);
and UO_739 (O_739,N_29857,N_29901);
nand UO_740 (O_740,N_29499,N_29654);
or UO_741 (O_741,N_29977,N_29484);
nand UO_742 (O_742,N_29574,N_29738);
nor UO_743 (O_743,N_29531,N_29774);
nand UO_744 (O_744,N_29604,N_29449);
and UO_745 (O_745,N_29546,N_29816);
or UO_746 (O_746,N_29541,N_29849);
nor UO_747 (O_747,N_29760,N_29406);
and UO_748 (O_748,N_29506,N_29854);
nor UO_749 (O_749,N_29407,N_29598);
nor UO_750 (O_750,N_29685,N_29872);
xnor UO_751 (O_751,N_29924,N_29914);
nor UO_752 (O_752,N_29491,N_29941);
or UO_753 (O_753,N_29548,N_29943);
and UO_754 (O_754,N_29841,N_29471);
and UO_755 (O_755,N_29726,N_29587);
nor UO_756 (O_756,N_29429,N_29849);
or UO_757 (O_757,N_29667,N_29767);
nor UO_758 (O_758,N_29885,N_29547);
nand UO_759 (O_759,N_29468,N_29934);
or UO_760 (O_760,N_29512,N_29493);
nor UO_761 (O_761,N_29919,N_29641);
nor UO_762 (O_762,N_29862,N_29976);
or UO_763 (O_763,N_29932,N_29831);
and UO_764 (O_764,N_29496,N_29663);
or UO_765 (O_765,N_29703,N_29616);
nor UO_766 (O_766,N_29577,N_29765);
and UO_767 (O_767,N_29956,N_29957);
nand UO_768 (O_768,N_29851,N_29603);
and UO_769 (O_769,N_29825,N_29913);
and UO_770 (O_770,N_29840,N_29624);
or UO_771 (O_771,N_29583,N_29873);
nor UO_772 (O_772,N_29469,N_29670);
nand UO_773 (O_773,N_29517,N_29748);
nor UO_774 (O_774,N_29421,N_29970);
nor UO_775 (O_775,N_29847,N_29864);
nor UO_776 (O_776,N_29478,N_29831);
xnor UO_777 (O_777,N_29689,N_29576);
nor UO_778 (O_778,N_29720,N_29989);
and UO_779 (O_779,N_29840,N_29436);
or UO_780 (O_780,N_29920,N_29745);
nand UO_781 (O_781,N_29967,N_29507);
nand UO_782 (O_782,N_29820,N_29551);
nand UO_783 (O_783,N_29913,N_29463);
or UO_784 (O_784,N_29960,N_29903);
nor UO_785 (O_785,N_29608,N_29867);
nor UO_786 (O_786,N_29852,N_29797);
and UO_787 (O_787,N_29990,N_29856);
xnor UO_788 (O_788,N_29665,N_29902);
nor UO_789 (O_789,N_29598,N_29559);
nand UO_790 (O_790,N_29924,N_29963);
nand UO_791 (O_791,N_29938,N_29690);
or UO_792 (O_792,N_29707,N_29572);
xor UO_793 (O_793,N_29826,N_29498);
nor UO_794 (O_794,N_29534,N_29555);
nor UO_795 (O_795,N_29717,N_29621);
or UO_796 (O_796,N_29712,N_29592);
or UO_797 (O_797,N_29739,N_29940);
nor UO_798 (O_798,N_29788,N_29431);
nor UO_799 (O_799,N_29821,N_29830);
nand UO_800 (O_800,N_29501,N_29885);
or UO_801 (O_801,N_29665,N_29456);
and UO_802 (O_802,N_29897,N_29900);
and UO_803 (O_803,N_29759,N_29528);
nor UO_804 (O_804,N_29672,N_29801);
nor UO_805 (O_805,N_29501,N_29849);
and UO_806 (O_806,N_29658,N_29606);
nor UO_807 (O_807,N_29946,N_29760);
nor UO_808 (O_808,N_29810,N_29978);
nor UO_809 (O_809,N_29908,N_29948);
and UO_810 (O_810,N_29746,N_29974);
nor UO_811 (O_811,N_29472,N_29960);
and UO_812 (O_812,N_29822,N_29561);
and UO_813 (O_813,N_29762,N_29482);
nor UO_814 (O_814,N_29749,N_29915);
nand UO_815 (O_815,N_29733,N_29518);
and UO_816 (O_816,N_29813,N_29868);
nor UO_817 (O_817,N_29830,N_29805);
or UO_818 (O_818,N_29621,N_29829);
nor UO_819 (O_819,N_29703,N_29676);
nand UO_820 (O_820,N_29750,N_29995);
and UO_821 (O_821,N_29895,N_29701);
nand UO_822 (O_822,N_29926,N_29747);
nor UO_823 (O_823,N_29861,N_29744);
nor UO_824 (O_824,N_29996,N_29612);
nor UO_825 (O_825,N_29950,N_29751);
nor UO_826 (O_826,N_29738,N_29557);
nand UO_827 (O_827,N_29714,N_29683);
or UO_828 (O_828,N_29950,N_29739);
nor UO_829 (O_829,N_29939,N_29538);
or UO_830 (O_830,N_29777,N_29810);
or UO_831 (O_831,N_29719,N_29999);
and UO_832 (O_832,N_29864,N_29638);
nor UO_833 (O_833,N_29621,N_29973);
or UO_834 (O_834,N_29781,N_29922);
nand UO_835 (O_835,N_29733,N_29536);
nand UO_836 (O_836,N_29563,N_29888);
and UO_837 (O_837,N_29719,N_29767);
or UO_838 (O_838,N_29687,N_29993);
and UO_839 (O_839,N_29959,N_29964);
xnor UO_840 (O_840,N_29668,N_29483);
or UO_841 (O_841,N_29619,N_29540);
nand UO_842 (O_842,N_29588,N_29784);
nor UO_843 (O_843,N_29707,N_29960);
nor UO_844 (O_844,N_29619,N_29774);
and UO_845 (O_845,N_29593,N_29930);
nand UO_846 (O_846,N_29929,N_29653);
xnor UO_847 (O_847,N_29934,N_29584);
nor UO_848 (O_848,N_29898,N_29792);
or UO_849 (O_849,N_29419,N_29418);
nor UO_850 (O_850,N_29816,N_29523);
or UO_851 (O_851,N_29861,N_29522);
nor UO_852 (O_852,N_29697,N_29486);
nor UO_853 (O_853,N_29576,N_29919);
nand UO_854 (O_854,N_29969,N_29476);
nor UO_855 (O_855,N_29852,N_29407);
nand UO_856 (O_856,N_29413,N_29495);
nor UO_857 (O_857,N_29902,N_29846);
nor UO_858 (O_858,N_29716,N_29636);
nor UO_859 (O_859,N_29993,N_29422);
nor UO_860 (O_860,N_29525,N_29922);
or UO_861 (O_861,N_29995,N_29459);
nand UO_862 (O_862,N_29709,N_29951);
nand UO_863 (O_863,N_29866,N_29946);
and UO_864 (O_864,N_29747,N_29701);
and UO_865 (O_865,N_29487,N_29421);
or UO_866 (O_866,N_29960,N_29920);
and UO_867 (O_867,N_29691,N_29854);
and UO_868 (O_868,N_29661,N_29543);
or UO_869 (O_869,N_29758,N_29813);
nor UO_870 (O_870,N_29674,N_29910);
nand UO_871 (O_871,N_29777,N_29721);
nand UO_872 (O_872,N_29793,N_29938);
and UO_873 (O_873,N_29845,N_29407);
nand UO_874 (O_874,N_29540,N_29880);
or UO_875 (O_875,N_29445,N_29460);
nor UO_876 (O_876,N_29832,N_29555);
or UO_877 (O_877,N_29436,N_29825);
and UO_878 (O_878,N_29453,N_29829);
and UO_879 (O_879,N_29628,N_29485);
nor UO_880 (O_880,N_29725,N_29832);
and UO_881 (O_881,N_29521,N_29958);
nand UO_882 (O_882,N_29924,N_29463);
or UO_883 (O_883,N_29637,N_29499);
xnor UO_884 (O_884,N_29616,N_29673);
or UO_885 (O_885,N_29789,N_29402);
and UO_886 (O_886,N_29991,N_29707);
nor UO_887 (O_887,N_29989,N_29412);
and UO_888 (O_888,N_29593,N_29937);
or UO_889 (O_889,N_29666,N_29427);
nand UO_890 (O_890,N_29543,N_29958);
nor UO_891 (O_891,N_29486,N_29896);
nor UO_892 (O_892,N_29626,N_29683);
and UO_893 (O_893,N_29843,N_29556);
nand UO_894 (O_894,N_29438,N_29612);
and UO_895 (O_895,N_29843,N_29416);
and UO_896 (O_896,N_29914,N_29652);
and UO_897 (O_897,N_29584,N_29514);
xor UO_898 (O_898,N_29478,N_29531);
nor UO_899 (O_899,N_29798,N_29922);
nand UO_900 (O_900,N_29576,N_29771);
nor UO_901 (O_901,N_29546,N_29835);
or UO_902 (O_902,N_29907,N_29880);
nand UO_903 (O_903,N_29969,N_29664);
or UO_904 (O_904,N_29765,N_29597);
nor UO_905 (O_905,N_29556,N_29988);
nor UO_906 (O_906,N_29632,N_29699);
or UO_907 (O_907,N_29473,N_29554);
or UO_908 (O_908,N_29576,N_29692);
nor UO_909 (O_909,N_29885,N_29764);
nand UO_910 (O_910,N_29947,N_29459);
nor UO_911 (O_911,N_29755,N_29538);
and UO_912 (O_912,N_29586,N_29493);
xnor UO_913 (O_913,N_29513,N_29507);
and UO_914 (O_914,N_29718,N_29659);
nor UO_915 (O_915,N_29594,N_29865);
nor UO_916 (O_916,N_29645,N_29703);
nand UO_917 (O_917,N_29688,N_29531);
nand UO_918 (O_918,N_29649,N_29914);
and UO_919 (O_919,N_29434,N_29639);
or UO_920 (O_920,N_29911,N_29635);
nor UO_921 (O_921,N_29652,N_29542);
or UO_922 (O_922,N_29740,N_29717);
and UO_923 (O_923,N_29513,N_29795);
or UO_924 (O_924,N_29471,N_29528);
or UO_925 (O_925,N_29866,N_29656);
nand UO_926 (O_926,N_29779,N_29658);
nor UO_927 (O_927,N_29958,N_29846);
nor UO_928 (O_928,N_29467,N_29641);
or UO_929 (O_929,N_29674,N_29697);
nand UO_930 (O_930,N_29867,N_29795);
nor UO_931 (O_931,N_29640,N_29539);
and UO_932 (O_932,N_29551,N_29947);
and UO_933 (O_933,N_29510,N_29749);
nand UO_934 (O_934,N_29767,N_29933);
and UO_935 (O_935,N_29525,N_29676);
nand UO_936 (O_936,N_29935,N_29968);
nand UO_937 (O_937,N_29710,N_29734);
or UO_938 (O_938,N_29850,N_29683);
or UO_939 (O_939,N_29789,N_29449);
and UO_940 (O_940,N_29754,N_29686);
or UO_941 (O_941,N_29928,N_29449);
xor UO_942 (O_942,N_29465,N_29985);
nand UO_943 (O_943,N_29585,N_29754);
or UO_944 (O_944,N_29779,N_29564);
and UO_945 (O_945,N_29551,N_29733);
and UO_946 (O_946,N_29953,N_29425);
and UO_947 (O_947,N_29602,N_29647);
or UO_948 (O_948,N_29942,N_29978);
nand UO_949 (O_949,N_29989,N_29509);
nand UO_950 (O_950,N_29606,N_29430);
nand UO_951 (O_951,N_29696,N_29885);
nand UO_952 (O_952,N_29433,N_29512);
nand UO_953 (O_953,N_29513,N_29883);
nor UO_954 (O_954,N_29647,N_29732);
nand UO_955 (O_955,N_29811,N_29450);
and UO_956 (O_956,N_29432,N_29769);
nor UO_957 (O_957,N_29822,N_29562);
nor UO_958 (O_958,N_29631,N_29859);
and UO_959 (O_959,N_29771,N_29420);
nor UO_960 (O_960,N_29457,N_29522);
nor UO_961 (O_961,N_29504,N_29637);
or UO_962 (O_962,N_29709,N_29413);
nand UO_963 (O_963,N_29461,N_29875);
or UO_964 (O_964,N_29863,N_29602);
or UO_965 (O_965,N_29889,N_29508);
nor UO_966 (O_966,N_29617,N_29642);
nand UO_967 (O_967,N_29799,N_29683);
and UO_968 (O_968,N_29727,N_29826);
nor UO_969 (O_969,N_29440,N_29969);
and UO_970 (O_970,N_29657,N_29471);
nand UO_971 (O_971,N_29686,N_29824);
nor UO_972 (O_972,N_29633,N_29996);
nor UO_973 (O_973,N_29575,N_29543);
nand UO_974 (O_974,N_29520,N_29831);
nand UO_975 (O_975,N_29927,N_29426);
nor UO_976 (O_976,N_29443,N_29785);
nor UO_977 (O_977,N_29810,N_29962);
nor UO_978 (O_978,N_29905,N_29968);
and UO_979 (O_979,N_29749,N_29863);
and UO_980 (O_980,N_29758,N_29560);
nor UO_981 (O_981,N_29591,N_29881);
nor UO_982 (O_982,N_29842,N_29686);
and UO_983 (O_983,N_29787,N_29864);
or UO_984 (O_984,N_29797,N_29587);
or UO_985 (O_985,N_29985,N_29521);
or UO_986 (O_986,N_29732,N_29578);
nand UO_987 (O_987,N_29661,N_29415);
or UO_988 (O_988,N_29874,N_29683);
or UO_989 (O_989,N_29864,N_29678);
nand UO_990 (O_990,N_29627,N_29947);
or UO_991 (O_991,N_29854,N_29623);
and UO_992 (O_992,N_29688,N_29990);
and UO_993 (O_993,N_29551,N_29827);
xnor UO_994 (O_994,N_29885,N_29474);
and UO_995 (O_995,N_29787,N_29498);
and UO_996 (O_996,N_29646,N_29490);
and UO_997 (O_997,N_29606,N_29499);
and UO_998 (O_998,N_29643,N_29684);
and UO_999 (O_999,N_29460,N_29577);
or UO_1000 (O_1000,N_29432,N_29822);
and UO_1001 (O_1001,N_29526,N_29891);
nand UO_1002 (O_1002,N_29819,N_29671);
nand UO_1003 (O_1003,N_29604,N_29907);
nor UO_1004 (O_1004,N_29400,N_29960);
and UO_1005 (O_1005,N_29606,N_29818);
and UO_1006 (O_1006,N_29505,N_29934);
nand UO_1007 (O_1007,N_29486,N_29607);
nand UO_1008 (O_1008,N_29884,N_29753);
or UO_1009 (O_1009,N_29641,N_29838);
nor UO_1010 (O_1010,N_29636,N_29834);
or UO_1011 (O_1011,N_29539,N_29644);
or UO_1012 (O_1012,N_29625,N_29626);
or UO_1013 (O_1013,N_29793,N_29807);
xnor UO_1014 (O_1014,N_29558,N_29567);
nor UO_1015 (O_1015,N_29552,N_29530);
and UO_1016 (O_1016,N_29544,N_29856);
nand UO_1017 (O_1017,N_29431,N_29411);
nand UO_1018 (O_1018,N_29538,N_29821);
nand UO_1019 (O_1019,N_29444,N_29932);
nand UO_1020 (O_1020,N_29905,N_29840);
nand UO_1021 (O_1021,N_29844,N_29712);
nor UO_1022 (O_1022,N_29733,N_29779);
nor UO_1023 (O_1023,N_29486,N_29880);
nor UO_1024 (O_1024,N_29667,N_29413);
and UO_1025 (O_1025,N_29696,N_29851);
or UO_1026 (O_1026,N_29614,N_29576);
xnor UO_1027 (O_1027,N_29691,N_29527);
nor UO_1028 (O_1028,N_29923,N_29896);
nand UO_1029 (O_1029,N_29651,N_29632);
or UO_1030 (O_1030,N_29968,N_29525);
nor UO_1031 (O_1031,N_29489,N_29687);
and UO_1032 (O_1032,N_29923,N_29487);
nand UO_1033 (O_1033,N_29770,N_29651);
nor UO_1034 (O_1034,N_29827,N_29788);
nor UO_1035 (O_1035,N_29861,N_29907);
nand UO_1036 (O_1036,N_29778,N_29683);
nand UO_1037 (O_1037,N_29770,N_29758);
or UO_1038 (O_1038,N_29935,N_29741);
nor UO_1039 (O_1039,N_29521,N_29689);
nand UO_1040 (O_1040,N_29731,N_29629);
nor UO_1041 (O_1041,N_29628,N_29878);
nor UO_1042 (O_1042,N_29818,N_29682);
nand UO_1043 (O_1043,N_29880,N_29429);
nand UO_1044 (O_1044,N_29929,N_29414);
nand UO_1045 (O_1045,N_29720,N_29611);
nand UO_1046 (O_1046,N_29508,N_29523);
nor UO_1047 (O_1047,N_29638,N_29427);
nor UO_1048 (O_1048,N_29443,N_29684);
nor UO_1049 (O_1049,N_29736,N_29844);
nor UO_1050 (O_1050,N_29435,N_29727);
nand UO_1051 (O_1051,N_29869,N_29658);
nor UO_1052 (O_1052,N_29532,N_29741);
nand UO_1053 (O_1053,N_29648,N_29637);
nor UO_1054 (O_1054,N_29611,N_29752);
nand UO_1055 (O_1055,N_29514,N_29573);
xor UO_1056 (O_1056,N_29947,N_29982);
and UO_1057 (O_1057,N_29995,N_29918);
and UO_1058 (O_1058,N_29907,N_29917);
nor UO_1059 (O_1059,N_29703,N_29915);
xnor UO_1060 (O_1060,N_29835,N_29930);
nand UO_1061 (O_1061,N_29841,N_29983);
nor UO_1062 (O_1062,N_29479,N_29929);
nor UO_1063 (O_1063,N_29704,N_29996);
nor UO_1064 (O_1064,N_29425,N_29572);
or UO_1065 (O_1065,N_29664,N_29673);
nand UO_1066 (O_1066,N_29980,N_29836);
nor UO_1067 (O_1067,N_29693,N_29474);
or UO_1068 (O_1068,N_29480,N_29682);
and UO_1069 (O_1069,N_29827,N_29649);
xor UO_1070 (O_1070,N_29549,N_29659);
and UO_1071 (O_1071,N_29694,N_29732);
and UO_1072 (O_1072,N_29704,N_29665);
nor UO_1073 (O_1073,N_29756,N_29571);
xnor UO_1074 (O_1074,N_29438,N_29724);
nor UO_1075 (O_1075,N_29776,N_29881);
or UO_1076 (O_1076,N_29691,N_29496);
and UO_1077 (O_1077,N_29454,N_29552);
and UO_1078 (O_1078,N_29909,N_29777);
nor UO_1079 (O_1079,N_29847,N_29839);
nor UO_1080 (O_1080,N_29995,N_29705);
nor UO_1081 (O_1081,N_29600,N_29619);
nand UO_1082 (O_1082,N_29997,N_29498);
or UO_1083 (O_1083,N_29762,N_29607);
nor UO_1084 (O_1084,N_29512,N_29593);
nand UO_1085 (O_1085,N_29691,N_29877);
or UO_1086 (O_1086,N_29625,N_29561);
nand UO_1087 (O_1087,N_29849,N_29700);
nand UO_1088 (O_1088,N_29601,N_29979);
and UO_1089 (O_1089,N_29430,N_29722);
nand UO_1090 (O_1090,N_29870,N_29765);
nor UO_1091 (O_1091,N_29544,N_29662);
nor UO_1092 (O_1092,N_29555,N_29734);
and UO_1093 (O_1093,N_29692,N_29408);
or UO_1094 (O_1094,N_29580,N_29514);
and UO_1095 (O_1095,N_29859,N_29884);
nand UO_1096 (O_1096,N_29979,N_29459);
and UO_1097 (O_1097,N_29996,N_29507);
nor UO_1098 (O_1098,N_29622,N_29916);
nand UO_1099 (O_1099,N_29430,N_29444);
nand UO_1100 (O_1100,N_29949,N_29843);
or UO_1101 (O_1101,N_29963,N_29791);
and UO_1102 (O_1102,N_29542,N_29937);
nor UO_1103 (O_1103,N_29906,N_29554);
nor UO_1104 (O_1104,N_29779,N_29442);
or UO_1105 (O_1105,N_29876,N_29960);
nand UO_1106 (O_1106,N_29869,N_29833);
nand UO_1107 (O_1107,N_29728,N_29597);
or UO_1108 (O_1108,N_29850,N_29450);
nand UO_1109 (O_1109,N_29636,N_29915);
nor UO_1110 (O_1110,N_29974,N_29657);
nor UO_1111 (O_1111,N_29492,N_29796);
nand UO_1112 (O_1112,N_29569,N_29933);
or UO_1113 (O_1113,N_29723,N_29481);
nor UO_1114 (O_1114,N_29509,N_29695);
xnor UO_1115 (O_1115,N_29614,N_29664);
and UO_1116 (O_1116,N_29821,N_29798);
nand UO_1117 (O_1117,N_29441,N_29827);
and UO_1118 (O_1118,N_29840,N_29719);
and UO_1119 (O_1119,N_29807,N_29908);
nand UO_1120 (O_1120,N_29989,N_29499);
and UO_1121 (O_1121,N_29662,N_29753);
and UO_1122 (O_1122,N_29886,N_29542);
or UO_1123 (O_1123,N_29800,N_29686);
nand UO_1124 (O_1124,N_29899,N_29863);
or UO_1125 (O_1125,N_29627,N_29938);
nor UO_1126 (O_1126,N_29879,N_29724);
xnor UO_1127 (O_1127,N_29926,N_29889);
or UO_1128 (O_1128,N_29989,N_29823);
or UO_1129 (O_1129,N_29698,N_29735);
or UO_1130 (O_1130,N_29489,N_29898);
and UO_1131 (O_1131,N_29863,N_29830);
and UO_1132 (O_1132,N_29497,N_29487);
nor UO_1133 (O_1133,N_29525,N_29669);
and UO_1134 (O_1134,N_29818,N_29914);
nand UO_1135 (O_1135,N_29575,N_29680);
nand UO_1136 (O_1136,N_29882,N_29755);
nor UO_1137 (O_1137,N_29570,N_29893);
nor UO_1138 (O_1138,N_29985,N_29699);
and UO_1139 (O_1139,N_29866,N_29682);
and UO_1140 (O_1140,N_29992,N_29804);
and UO_1141 (O_1141,N_29480,N_29665);
nand UO_1142 (O_1142,N_29432,N_29580);
and UO_1143 (O_1143,N_29552,N_29895);
or UO_1144 (O_1144,N_29415,N_29980);
nor UO_1145 (O_1145,N_29531,N_29957);
nand UO_1146 (O_1146,N_29490,N_29560);
or UO_1147 (O_1147,N_29552,N_29784);
xor UO_1148 (O_1148,N_29732,N_29588);
or UO_1149 (O_1149,N_29417,N_29889);
nand UO_1150 (O_1150,N_29413,N_29662);
nor UO_1151 (O_1151,N_29554,N_29442);
or UO_1152 (O_1152,N_29782,N_29706);
or UO_1153 (O_1153,N_29954,N_29537);
or UO_1154 (O_1154,N_29564,N_29775);
or UO_1155 (O_1155,N_29647,N_29576);
or UO_1156 (O_1156,N_29839,N_29853);
nand UO_1157 (O_1157,N_29672,N_29713);
and UO_1158 (O_1158,N_29598,N_29915);
nor UO_1159 (O_1159,N_29694,N_29703);
and UO_1160 (O_1160,N_29626,N_29848);
nor UO_1161 (O_1161,N_29815,N_29450);
and UO_1162 (O_1162,N_29628,N_29624);
and UO_1163 (O_1163,N_29899,N_29628);
nand UO_1164 (O_1164,N_29863,N_29664);
nor UO_1165 (O_1165,N_29481,N_29664);
and UO_1166 (O_1166,N_29435,N_29449);
nor UO_1167 (O_1167,N_29797,N_29491);
nor UO_1168 (O_1168,N_29923,N_29929);
and UO_1169 (O_1169,N_29455,N_29977);
and UO_1170 (O_1170,N_29679,N_29796);
nand UO_1171 (O_1171,N_29533,N_29493);
nand UO_1172 (O_1172,N_29999,N_29907);
nand UO_1173 (O_1173,N_29786,N_29909);
and UO_1174 (O_1174,N_29759,N_29649);
nor UO_1175 (O_1175,N_29412,N_29775);
nand UO_1176 (O_1176,N_29774,N_29750);
nor UO_1177 (O_1177,N_29750,N_29981);
and UO_1178 (O_1178,N_29461,N_29827);
or UO_1179 (O_1179,N_29714,N_29638);
or UO_1180 (O_1180,N_29883,N_29673);
and UO_1181 (O_1181,N_29637,N_29716);
or UO_1182 (O_1182,N_29943,N_29732);
or UO_1183 (O_1183,N_29957,N_29570);
nand UO_1184 (O_1184,N_29899,N_29925);
or UO_1185 (O_1185,N_29648,N_29729);
and UO_1186 (O_1186,N_29434,N_29998);
and UO_1187 (O_1187,N_29937,N_29617);
nor UO_1188 (O_1188,N_29915,N_29631);
nand UO_1189 (O_1189,N_29793,N_29751);
nand UO_1190 (O_1190,N_29710,N_29735);
nor UO_1191 (O_1191,N_29416,N_29526);
nor UO_1192 (O_1192,N_29668,N_29723);
nand UO_1193 (O_1193,N_29402,N_29810);
xor UO_1194 (O_1194,N_29913,N_29797);
or UO_1195 (O_1195,N_29584,N_29827);
and UO_1196 (O_1196,N_29683,N_29548);
or UO_1197 (O_1197,N_29703,N_29796);
or UO_1198 (O_1198,N_29509,N_29558);
or UO_1199 (O_1199,N_29839,N_29515);
nand UO_1200 (O_1200,N_29826,N_29691);
nand UO_1201 (O_1201,N_29808,N_29867);
or UO_1202 (O_1202,N_29902,N_29747);
nand UO_1203 (O_1203,N_29414,N_29460);
and UO_1204 (O_1204,N_29549,N_29587);
nor UO_1205 (O_1205,N_29451,N_29916);
or UO_1206 (O_1206,N_29782,N_29658);
nor UO_1207 (O_1207,N_29675,N_29863);
or UO_1208 (O_1208,N_29767,N_29803);
nand UO_1209 (O_1209,N_29500,N_29625);
nor UO_1210 (O_1210,N_29937,N_29497);
and UO_1211 (O_1211,N_29642,N_29756);
nand UO_1212 (O_1212,N_29780,N_29441);
or UO_1213 (O_1213,N_29429,N_29568);
nor UO_1214 (O_1214,N_29415,N_29657);
nand UO_1215 (O_1215,N_29439,N_29459);
and UO_1216 (O_1216,N_29786,N_29478);
nand UO_1217 (O_1217,N_29688,N_29959);
nor UO_1218 (O_1218,N_29812,N_29813);
nor UO_1219 (O_1219,N_29463,N_29447);
nand UO_1220 (O_1220,N_29465,N_29468);
nor UO_1221 (O_1221,N_29552,N_29614);
and UO_1222 (O_1222,N_29436,N_29729);
nand UO_1223 (O_1223,N_29659,N_29618);
or UO_1224 (O_1224,N_29637,N_29798);
or UO_1225 (O_1225,N_29966,N_29599);
nor UO_1226 (O_1226,N_29848,N_29507);
and UO_1227 (O_1227,N_29875,N_29902);
and UO_1228 (O_1228,N_29631,N_29882);
nand UO_1229 (O_1229,N_29921,N_29932);
and UO_1230 (O_1230,N_29463,N_29859);
nor UO_1231 (O_1231,N_29466,N_29696);
or UO_1232 (O_1232,N_29470,N_29487);
nor UO_1233 (O_1233,N_29606,N_29517);
and UO_1234 (O_1234,N_29907,N_29770);
nor UO_1235 (O_1235,N_29798,N_29937);
or UO_1236 (O_1236,N_29837,N_29655);
and UO_1237 (O_1237,N_29436,N_29742);
or UO_1238 (O_1238,N_29641,N_29869);
or UO_1239 (O_1239,N_29514,N_29884);
or UO_1240 (O_1240,N_29530,N_29749);
and UO_1241 (O_1241,N_29476,N_29730);
nand UO_1242 (O_1242,N_29934,N_29888);
and UO_1243 (O_1243,N_29549,N_29851);
and UO_1244 (O_1244,N_29414,N_29784);
nor UO_1245 (O_1245,N_29875,N_29823);
nand UO_1246 (O_1246,N_29679,N_29862);
or UO_1247 (O_1247,N_29649,N_29836);
nand UO_1248 (O_1248,N_29982,N_29889);
nand UO_1249 (O_1249,N_29787,N_29960);
nor UO_1250 (O_1250,N_29637,N_29938);
nand UO_1251 (O_1251,N_29580,N_29472);
or UO_1252 (O_1252,N_29827,N_29715);
or UO_1253 (O_1253,N_29576,N_29816);
or UO_1254 (O_1254,N_29540,N_29404);
and UO_1255 (O_1255,N_29900,N_29859);
nor UO_1256 (O_1256,N_29436,N_29683);
or UO_1257 (O_1257,N_29799,N_29435);
nor UO_1258 (O_1258,N_29718,N_29672);
nor UO_1259 (O_1259,N_29628,N_29494);
or UO_1260 (O_1260,N_29472,N_29464);
or UO_1261 (O_1261,N_29956,N_29671);
and UO_1262 (O_1262,N_29655,N_29590);
or UO_1263 (O_1263,N_29778,N_29848);
nor UO_1264 (O_1264,N_29442,N_29508);
and UO_1265 (O_1265,N_29992,N_29588);
or UO_1266 (O_1266,N_29907,N_29879);
or UO_1267 (O_1267,N_29533,N_29816);
nand UO_1268 (O_1268,N_29915,N_29817);
or UO_1269 (O_1269,N_29566,N_29862);
nor UO_1270 (O_1270,N_29890,N_29707);
nand UO_1271 (O_1271,N_29913,N_29513);
nand UO_1272 (O_1272,N_29607,N_29889);
nor UO_1273 (O_1273,N_29908,N_29463);
or UO_1274 (O_1274,N_29948,N_29994);
or UO_1275 (O_1275,N_29704,N_29983);
or UO_1276 (O_1276,N_29944,N_29694);
and UO_1277 (O_1277,N_29697,N_29965);
nand UO_1278 (O_1278,N_29930,N_29718);
and UO_1279 (O_1279,N_29680,N_29693);
nand UO_1280 (O_1280,N_29518,N_29472);
or UO_1281 (O_1281,N_29841,N_29731);
nor UO_1282 (O_1282,N_29553,N_29822);
and UO_1283 (O_1283,N_29927,N_29678);
or UO_1284 (O_1284,N_29844,N_29585);
and UO_1285 (O_1285,N_29604,N_29916);
nor UO_1286 (O_1286,N_29520,N_29764);
nor UO_1287 (O_1287,N_29997,N_29952);
nand UO_1288 (O_1288,N_29530,N_29669);
nand UO_1289 (O_1289,N_29576,N_29700);
nand UO_1290 (O_1290,N_29583,N_29591);
nand UO_1291 (O_1291,N_29753,N_29626);
or UO_1292 (O_1292,N_29621,N_29479);
and UO_1293 (O_1293,N_29597,N_29731);
nor UO_1294 (O_1294,N_29640,N_29598);
or UO_1295 (O_1295,N_29569,N_29959);
and UO_1296 (O_1296,N_29880,N_29410);
and UO_1297 (O_1297,N_29770,N_29764);
nand UO_1298 (O_1298,N_29664,N_29898);
or UO_1299 (O_1299,N_29458,N_29782);
and UO_1300 (O_1300,N_29633,N_29982);
nor UO_1301 (O_1301,N_29683,N_29936);
or UO_1302 (O_1302,N_29428,N_29971);
or UO_1303 (O_1303,N_29921,N_29618);
nand UO_1304 (O_1304,N_29780,N_29621);
nand UO_1305 (O_1305,N_29921,N_29978);
and UO_1306 (O_1306,N_29455,N_29651);
and UO_1307 (O_1307,N_29983,N_29873);
and UO_1308 (O_1308,N_29657,N_29928);
and UO_1309 (O_1309,N_29526,N_29505);
nand UO_1310 (O_1310,N_29808,N_29619);
and UO_1311 (O_1311,N_29877,N_29755);
nand UO_1312 (O_1312,N_29440,N_29962);
or UO_1313 (O_1313,N_29598,N_29498);
nor UO_1314 (O_1314,N_29651,N_29858);
and UO_1315 (O_1315,N_29901,N_29881);
and UO_1316 (O_1316,N_29899,N_29763);
or UO_1317 (O_1317,N_29575,N_29530);
or UO_1318 (O_1318,N_29792,N_29939);
and UO_1319 (O_1319,N_29527,N_29791);
or UO_1320 (O_1320,N_29660,N_29757);
nor UO_1321 (O_1321,N_29584,N_29419);
and UO_1322 (O_1322,N_29432,N_29497);
or UO_1323 (O_1323,N_29521,N_29979);
or UO_1324 (O_1324,N_29983,N_29488);
xnor UO_1325 (O_1325,N_29648,N_29557);
nand UO_1326 (O_1326,N_29549,N_29450);
xnor UO_1327 (O_1327,N_29966,N_29972);
nor UO_1328 (O_1328,N_29794,N_29879);
or UO_1329 (O_1329,N_29798,N_29830);
or UO_1330 (O_1330,N_29684,N_29587);
nor UO_1331 (O_1331,N_29564,N_29572);
xor UO_1332 (O_1332,N_29662,N_29575);
and UO_1333 (O_1333,N_29966,N_29580);
or UO_1334 (O_1334,N_29604,N_29724);
xor UO_1335 (O_1335,N_29790,N_29921);
nor UO_1336 (O_1336,N_29748,N_29456);
nor UO_1337 (O_1337,N_29999,N_29678);
and UO_1338 (O_1338,N_29433,N_29954);
nand UO_1339 (O_1339,N_29935,N_29563);
nand UO_1340 (O_1340,N_29706,N_29625);
nor UO_1341 (O_1341,N_29473,N_29679);
nand UO_1342 (O_1342,N_29594,N_29826);
nand UO_1343 (O_1343,N_29547,N_29916);
nand UO_1344 (O_1344,N_29776,N_29524);
xor UO_1345 (O_1345,N_29678,N_29591);
nor UO_1346 (O_1346,N_29754,N_29620);
nand UO_1347 (O_1347,N_29515,N_29845);
nand UO_1348 (O_1348,N_29862,N_29584);
or UO_1349 (O_1349,N_29809,N_29608);
and UO_1350 (O_1350,N_29818,N_29535);
and UO_1351 (O_1351,N_29727,N_29762);
nand UO_1352 (O_1352,N_29785,N_29841);
and UO_1353 (O_1353,N_29440,N_29479);
nand UO_1354 (O_1354,N_29925,N_29413);
or UO_1355 (O_1355,N_29693,N_29782);
nor UO_1356 (O_1356,N_29738,N_29913);
and UO_1357 (O_1357,N_29446,N_29490);
nor UO_1358 (O_1358,N_29557,N_29998);
nor UO_1359 (O_1359,N_29526,N_29847);
nor UO_1360 (O_1360,N_29774,N_29853);
nand UO_1361 (O_1361,N_29443,N_29650);
nand UO_1362 (O_1362,N_29440,N_29431);
xnor UO_1363 (O_1363,N_29977,N_29567);
and UO_1364 (O_1364,N_29443,N_29431);
nor UO_1365 (O_1365,N_29950,N_29597);
nand UO_1366 (O_1366,N_29552,N_29489);
or UO_1367 (O_1367,N_29999,N_29635);
or UO_1368 (O_1368,N_29983,N_29741);
nor UO_1369 (O_1369,N_29652,N_29831);
or UO_1370 (O_1370,N_29893,N_29632);
or UO_1371 (O_1371,N_29745,N_29521);
and UO_1372 (O_1372,N_29761,N_29801);
nand UO_1373 (O_1373,N_29794,N_29418);
nand UO_1374 (O_1374,N_29630,N_29491);
or UO_1375 (O_1375,N_29672,N_29632);
nand UO_1376 (O_1376,N_29640,N_29639);
and UO_1377 (O_1377,N_29898,N_29468);
and UO_1378 (O_1378,N_29770,N_29763);
and UO_1379 (O_1379,N_29847,N_29998);
or UO_1380 (O_1380,N_29825,N_29883);
nor UO_1381 (O_1381,N_29919,N_29905);
or UO_1382 (O_1382,N_29525,N_29556);
nor UO_1383 (O_1383,N_29977,N_29514);
and UO_1384 (O_1384,N_29749,N_29499);
or UO_1385 (O_1385,N_29639,N_29661);
or UO_1386 (O_1386,N_29785,N_29488);
or UO_1387 (O_1387,N_29641,N_29962);
nor UO_1388 (O_1388,N_29913,N_29755);
nand UO_1389 (O_1389,N_29567,N_29474);
and UO_1390 (O_1390,N_29593,N_29922);
or UO_1391 (O_1391,N_29895,N_29414);
nand UO_1392 (O_1392,N_29740,N_29828);
nor UO_1393 (O_1393,N_29902,N_29807);
nor UO_1394 (O_1394,N_29731,N_29596);
xor UO_1395 (O_1395,N_29977,N_29720);
nand UO_1396 (O_1396,N_29743,N_29582);
nor UO_1397 (O_1397,N_29801,N_29993);
xor UO_1398 (O_1398,N_29412,N_29518);
or UO_1399 (O_1399,N_29440,N_29998);
nor UO_1400 (O_1400,N_29893,N_29788);
and UO_1401 (O_1401,N_29617,N_29579);
and UO_1402 (O_1402,N_29412,N_29960);
nand UO_1403 (O_1403,N_29610,N_29961);
nor UO_1404 (O_1404,N_29783,N_29768);
nand UO_1405 (O_1405,N_29887,N_29854);
nor UO_1406 (O_1406,N_29800,N_29906);
nand UO_1407 (O_1407,N_29531,N_29619);
nand UO_1408 (O_1408,N_29630,N_29850);
and UO_1409 (O_1409,N_29824,N_29558);
and UO_1410 (O_1410,N_29900,N_29668);
nand UO_1411 (O_1411,N_29913,N_29823);
or UO_1412 (O_1412,N_29762,N_29725);
and UO_1413 (O_1413,N_29740,N_29582);
xnor UO_1414 (O_1414,N_29964,N_29668);
or UO_1415 (O_1415,N_29412,N_29819);
nand UO_1416 (O_1416,N_29432,N_29443);
nand UO_1417 (O_1417,N_29861,N_29704);
and UO_1418 (O_1418,N_29863,N_29499);
nand UO_1419 (O_1419,N_29790,N_29538);
or UO_1420 (O_1420,N_29579,N_29882);
nor UO_1421 (O_1421,N_29654,N_29508);
nor UO_1422 (O_1422,N_29428,N_29605);
or UO_1423 (O_1423,N_29785,N_29820);
or UO_1424 (O_1424,N_29903,N_29632);
or UO_1425 (O_1425,N_29927,N_29714);
nor UO_1426 (O_1426,N_29510,N_29457);
nor UO_1427 (O_1427,N_29854,N_29798);
and UO_1428 (O_1428,N_29668,N_29505);
and UO_1429 (O_1429,N_29518,N_29856);
nor UO_1430 (O_1430,N_29532,N_29664);
nor UO_1431 (O_1431,N_29985,N_29476);
nand UO_1432 (O_1432,N_29621,N_29617);
and UO_1433 (O_1433,N_29541,N_29527);
or UO_1434 (O_1434,N_29735,N_29688);
nor UO_1435 (O_1435,N_29989,N_29874);
nand UO_1436 (O_1436,N_29773,N_29564);
or UO_1437 (O_1437,N_29689,N_29962);
nand UO_1438 (O_1438,N_29565,N_29883);
and UO_1439 (O_1439,N_29602,N_29687);
and UO_1440 (O_1440,N_29804,N_29906);
nand UO_1441 (O_1441,N_29436,N_29801);
and UO_1442 (O_1442,N_29980,N_29759);
nand UO_1443 (O_1443,N_29860,N_29930);
nand UO_1444 (O_1444,N_29594,N_29967);
nor UO_1445 (O_1445,N_29720,N_29822);
or UO_1446 (O_1446,N_29940,N_29523);
and UO_1447 (O_1447,N_29928,N_29577);
or UO_1448 (O_1448,N_29730,N_29671);
nor UO_1449 (O_1449,N_29509,N_29533);
nand UO_1450 (O_1450,N_29760,N_29871);
nor UO_1451 (O_1451,N_29744,N_29621);
nor UO_1452 (O_1452,N_29462,N_29861);
and UO_1453 (O_1453,N_29833,N_29758);
nand UO_1454 (O_1454,N_29900,N_29917);
and UO_1455 (O_1455,N_29484,N_29899);
nor UO_1456 (O_1456,N_29995,N_29680);
nand UO_1457 (O_1457,N_29579,N_29485);
or UO_1458 (O_1458,N_29840,N_29640);
nor UO_1459 (O_1459,N_29467,N_29767);
and UO_1460 (O_1460,N_29705,N_29443);
nand UO_1461 (O_1461,N_29643,N_29504);
or UO_1462 (O_1462,N_29576,N_29518);
and UO_1463 (O_1463,N_29407,N_29404);
nor UO_1464 (O_1464,N_29570,N_29702);
or UO_1465 (O_1465,N_29953,N_29802);
nand UO_1466 (O_1466,N_29760,N_29561);
nand UO_1467 (O_1467,N_29899,N_29746);
nor UO_1468 (O_1468,N_29549,N_29420);
and UO_1469 (O_1469,N_29930,N_29732);
and UO_1470 (O_1470,N_29487,N_29560);
xor UO_1471 (O_1471,N_29950,N_29512);
nor UO_1472 (O_1472,N_29792,N_29715);
and UO_1473 (O_1473,N_29549,N_29454);
and UO_1474 (O_1474,N_29400,N_29693);
nand UO_1475 (O_1475,N_29448,N_29973);
and UO_1476 (O_1476,N_29993,N_29829);
nand UO_1477 (O_1477,N_29687,N_29908);
or UO_1478 (O_1478,N_29726,N_29737);
and UO_1479 (O_1479,N_29586,N_29545);
nor UO_1480 (O_1480,N_29635,N_29708);
and UO_1481 (O_1481,N_29506,N_29615);
nand UO_1482 (O_1482,N_29792,N_29695);
and UO_1483 (O_1483,N_29950,N_29740);
nand UO_1484 (O_1484,N_29574,N_29594);
or UO_1485 (O_1485,N_29866,N_29467);
or UO_1486 (O_1486,N_29522,N_29743);
or UO_1487 (O_1487,N_29991,N_29419);
nand UO_1488 (O_1488,N_29784,N_29720);
nor UO_1489 (O_1489,N_29854,N_29414);
nor UO_1490 (O_1490,N_29872,N_29523);
or UO_1491 (O_1491,N_29643,N_29977);
nor UO_1492 (O_1492,N_29774,N_29891);
and UO_1493 (O_1493,N_29507,N_29677);
or UO_1494 (O_1494,N_29587,N_29493);
or UO_1495 (O_1495,N_29924,N_29904);
nand UO_1496 (O_1496,N_29550,N_29611);
and UO_1497 (O_1497,N_29598,N_29964);
nand UO_1498 (O_1498,N_29534,N_29783);
and UO_1499 (O_1499,N_29400,N_29635);
nor UO_1500 (O_1500,N_29705,N_29837);
nor UO_1501 (O_1501,N_29665,N_29702);
or UO_1502 (O_1502,N_29430,N_29630);
xnor UO_1503 (O_1503,N_29519,N_29547);
xnor UO_1504 (O_1504,N_29548,N_29741);
nor UO_1505 (O_1505,N_29983,N_29677);
and UO_1506 (O_1506,N_29815,N_29816);
nor UO_1507 (O_1507,N_29734,N_29949);
or UO_1508 (O_1508,N_29693,N_29855);
or UO_1509 (O_1509,N_29775,N_29974);
and UO_1510 (O_1510,N_29679,N_29765);
or UO_1511 (O_1511,N_29952,N_29896);
nor UO_1512 (O_1512,N_29736,N_29566);
or UO_1513 (O_1513,N_29452,N_29454);
nor UO_1514 (O_1514,N_29623,N_29862);
nand UO_1515 (O_1515,N_29595,N_29823);
xor UO_1516 (O_1516,N_29905,N_29470);
and UO_1517 (O_1517,N_29432,N_29585);
and UO_1518 (O_1518,N_29638,N_29987);
nand UO_1519 (O_1519,N_29406,N_29428);
and UO_1520 (O_1520,N_29921,N_29592);
and UO_1521 (O_1521,N_29811,N_29848);
or UO_1522 (O_1522,N_29491,N_29817);
nand UO_1523 (O_1523,N_29730,N_29788);
nand UO_1524 (O_1524,N_29613,N_29689);
and UO_1525 (O_1525,N_29452,N_29767);
nand UO_1526 (O_1526,N_29466,N_29488);
or UO_1527 (O_1527,N_29401,N_29513);
and UO_1528 (O_1528,N_29901,N_29878);
nor UO_1529 (O_1529,N_29797,N_29590);
or UO_1530 (O_1530,N_29710,N_29781);
and UO_1531 (O_1531,N_29917,N_29532);
nand UO_1532 (O_1532,N_29949,N_29424);
nand UO_1533 (O_1533,N_29969,N_29780);
or UO_1534 (O_1534,N_29417,N_29463);
nor UO_1535 (O_1535,N_29772,N_29739);
nand UO_1536 (O_1536,N_29911,N_29564);
nor UO_1537 (O_1537,N_29493,N_29781);
nand UO_1538 (O_1538,N_29434,N_29811);
and UO_1539 (O_1539,N_29542,N_29468);
nor UO_1540 (O_1540,N_29734,N_29869);
nor UO_1541 (O_1541,N_29796,N_29691);
xor UO_1542 (O_1542,N_29866,N_29677);
nor UO_1543 (O_1543,N_29507,N_29675);
nor UO_1544 (O_1544,N_29852,N_29765);
nand UO_1545 (O_1545,N_29659,N_29991);
or UO_1546 (O_1546,N_29465,N_29687);
or UO_1547 (O_1547,N_29898,N_29982);
nand UO_1548 (O_1548,N_29528,N_29449);
or UO_1549 (O_1549,N_29985,N_29848);
nor UO_1550 (O_1550,N_29408,N_29987);
and UO_1551 (O_1551,N_29510,N_29567);
nor UO_1552 (O_1552,N_29837,N_29946);
xnor UO_1553 (O_1553,N_29417,N_29800);
nand UO_1554 (O_1554,N_29499,N_29803);
or UO_1555 (O_1555,N_29507,N_29632);
nor UO_1556 (O_1556,N_29878,N_29681);
nand UO_1557 (O_1557,N_29955,N_29838);
and UO_1558 (O_1558,N_29705,N_29476);
nor UO_1559 (O_1559,N_29701,N_29906);
xnor UO_1560 (O_1560,N_29468,N_29600);
nand UO_1561 (O_1561,N_29753,N_29768);
and UO_1562 (O_1562,N_29960,N_29421);
and UO_1563 (O_1563,N_29740,N_29975);
or UO_1564 (O_1564,N_29439,N_29456);
and UO_1565 (O_1565,N_29779,N_29586);
or UO_1566 (O_1566,N_29733,N_29662);
nor UO_1567 (O_1567,N_29867,N_29688);
nand UO_1568 (O_1568,N_29787,N_29584);
or UO_1569 (O_1569,N_29657,N_29617);
or UO_1570 (O_1570,N_29447,N_29595);
nor UO_1571 (O_1571,N_29535,N_29581);
and UO_1572 (O_1572,N_29691,N_29603);
nor UO_1573 (O_1573,N_29441,N_29642);
nor UO_1574 (O_1574,N_29909,N_29870);
or UO_1575 (O_1575,N_29792,N_29692);
and UO_1576 (O_1576,N_29707,N_29609);
nor UO_1577 (O_1577,N_29470,N_29892);
nand UO_1578 (O_1578,N_29473,N_29904);
or UO_1579 (O_1579,N_29610,N_29683);
or UO_1580 (O_1580,N_29918,N_29491);
and UO_1581 (O_1581,N_29622,N_29477);
nor UO_1582 (O_1582,N_29805,N_29572);
and UO_1583 (O_1583,N_29656,N_29519);
nand UO_1584 (O_1584,N_29466,N_29555);
and UO_1585 (O_1585,N_29611,N_29675);
and UO_1586 (O_1586,N_29784,N_29682);
and UO_1587 (O_1587,N_29437,N_29653);
and UO_1588 (O_1588,N_29502,N_29564);
nor UO_1589 (O_1589,N_29997,N_29682);
or UO_1590 (O_1590,N_29743,N_29715);
or UO_1591 (O_1591,N_29840,N_29627);
and UO_1592 (O_1592,N_29872,N_29858);
nor UO_1593 (O_1593,N_29508,N_29977);
nand UO_1594 (O_1594,N_29596,N_29667);
or UO_1595 (O_1595,N_29484,N_29940);
nor UO_1596 (O_1596,N_29746,N_29933);
xor UO_1597 (O_1597,N_29531,N_29818);
nand UO_1598 (O_1598,N_29951,N_29539);
nand UO_1599 (O_1599,N_29713,N_29911);
nand UO_1600 (O_1600,N_29636,N_29997);
nand UO_1601 (O_1601,N_29506,N_29597);
and UO_1602 (O_1602,N_29897,N_29655);
or UO_1603 (O_1603,N_29498,N_29406);
nor UO_1604 (O_1604,N_29447,N_29981);
and UO_1605 (O_1605,N_29608,N_29836);
or UO_1606 (O_1606,N_29977,N_29933);
and UO_1607 (O_1607,N_29775,N_29557);
nand UO_1608 (O_1608,N_29662,N_29923);
nor UO_1609 (O_1609,N_29651,N_29897);
or UO_1610 (O_1610,N_29568,N_29643);
nor UO_1611 (O_1611,N_29717,N_29444);
or UO_1612 (O_1612,N_29799,N_29885);
and UO_1613 (O_1613,N_29803,N_29985);
nand UO_1614 (O_1614,N_29760,N_29764);
or UO_1615 (O_1615,N_29412,N_29918);
nand UO_1616 (O_1616,N_29952,N_29774);
nand UO_1617 (O_1617,N_29464,N_29421);
nand UO_1618 (O_1618,N_29558,N_29468);
nand UO_1619 (O_1619,N_29510,N_29943);
or UO_1620 (O_1620,N_29920,N_29969);
or UO_1621 (O_1621,N_29849,N_29404);
nand UO_1622 (O_1622,N_29414,N_29951);
or UO_1623 (O_1623,N_29629,N_29584);
xor UO_1624 (O_1624,N_29747,N_29767);
and UO_1625 (O_1625,N_29715,N_29458);
and UO_1626 (O_1626,N_29631,N_29507);
or UO_1627 (O_1627,N_29463,N_29736);
nor UO_1628 (O_1628,N_29778,N_29959);
nor UO_1629 (O_1629,N_29887,N_29414);
nor UO_1630 (O_1630,N_29487,N_29716);
and UO_1631 (O_1631,N_29499,N_29781);
nor UO_1632 (O_1632,N_29864,N_29580);
and UO_1633 (O_1633,N_29707,N_29535);
nand UO_1634 (O_1634,N_29940,N_29671);
nor UO_1635 (O_1635,N_29724,N_29768);
or UO_1636 (O_1636,N_29581,N_29490);
and UO_1637 (O_1637,N_29808,N_29438);
nand UO_1638 (O_1638,N_29975,N_29738);
or UO_1639 (O_1639,N_29705,N_29719);
and UO_1640 (O_1640,N_29991,N_29971);
nor UO_1641 (O_1641,N_29701,N_29957);
and UO_1642 (O_1642,N_29751,N_29993);
or UO_1643 (O_1643,N_29681,N_29445);
nor UO_1644 (O_1644,N_29723,N_29407);
and UO_1645 (O_1645,N_29765,N_29605);
or UO_1646 (O_1646,N_29547,N_29906);
nand UO_1647 (O_1647,N_29462,N_29690);
and UO_1648 (O_1648,N_29567,N_29413);
nand UO_1649 (O_1649,N_29444,N_29710);
nor UO_1650 (O_1650,N_29776,N_29402);
and UO_1651 (O_1651,N_29751,N_29960);
and UO_1652 (O_1652,N_29643,N_29891);
or UO_1653 (O_1653,N_29912,N_29882);
xnor UO_1654 (O_1654,N_29650,N_29980);
and UO_1655 (O_1655,N_29862,N_29969);
nor UO_1656 (O_1656,N_29976,N_29468);
nand UO_1657 (O_1657,N_29879,N_29694);
nor UO_1658 (O_1658,N_29459,N_29677);
nand UO_1659 (O_1659,N_29614,N_29679);
or UO_1660 (O_1660,N_29780,N_29485);
nor UO_1661 (O_1661,N_29818,N_29415);
nand UO_1662 (O_1662,N_29420,N_29809);
or UO_1663 (O_1663,N_29594,N_29841);
nor UO_1664 (O_1664,N_29496,N_29941);
and UO_1665 (O_1665,N_29640,N_29439);
nand UO_1666 (O_1666,N_29705,N_29698);
or UO_1667 (O_1667,N_29784,N_29607);
nor UO_1668 (O_1668,N_29628,N_29589);
or UO_1669 (O_1669,N_29518,N_29843);
and UO_1670 (O_1670,N_29604,N_29446);
or UO_1671 (O_1671,N_29676,N_29672);
nand UO_1672 (O_1672,N_29706,N_29865);
or UO_1673 (O_1673,N_29690,N_29724);
nor UO_1674 (O_1674,N_29461,N_29515);
nand UO_1675 (O_1675,N_29629,N_29433);
nand UO_1676 (O_1676,N_29627,N_29659);
and UO_1677 (O_1677,N_29999,N_29743);
and UO_1678 (O_1678,N_29733,N_29986);
and UO_1679 (O_1679,N_29605,N_29783);
nor UO_1680 (O_1680,N_29694,N_29480);
or UO_1681 (O_1681,N_29410,N_29769);
nand UO_1682 (O_1682,N_29846,N_29780);
nor UO_1683 (O_1683,N_29705,N_29623);
and UO_1684 (O_1684,N_29522,N_29903);
nor UO_1685 (O_1685,N_29559,N_29760);
nand UO_1686 (O_1686,N_29613,N_29759);
nand UO_1687 (O_1687,N_29883,N_29483);
and UO_1688 (O_1688,N_29481,N_29496);
xnor UO_1689 (O_1689,N_29492,N_29400);
nor UO_1690 (O_1690,N_29562,N_29870);
and UO_1691 (O_1691,N_29502,N_29478);
nand UO_1692 (O_1692,N_29769,N_29457);
xor UO_1693 (O_1693,N_29914,N_29544);
or UO_1694 (O_1694,N_29778,N_29667);
nand UO_1695 (O_1695,N_29843,N_29979);
nand UO_1696 (O_1696,N_29423,N_29524);
or UO_1697 (O_1697,N_29733,N_29495);
nor UO_1698 (O_1698,N_29442,N_29713);
or UO_1699 (O_1699,N_29598,N_29724);
and UO_1700 (O_1700,N_29502,N_29905);
or UO_1701 (O_1701,N_29715,N_29493);
nand UO_1702 (O_1702,N_29802,N_29876);
or UO_1703 (O_1703,N_29809,N_29826);
and UO_1704 (O_1704,N_29409,N_29971);
nand UO_1705 (O_1705,N_29938,N_29500);
nor UO_1706 (O_1706,N_29972,N_29424);
or UO_1707 (O_1707,N_29849,N_29899);
nor UO_1708 (O_1708,N_29465,N_29943);
nand UO_1709 (O_1709,N_29940,N_29679);
nand UO_1710 (O_1710,N_29425,N_29614);
and UO_1711 (O_1711,N_29579,N_29636);
nor UO_1712 (O_1712,N_29685,N_29464);
or UO_1713 (O_1713,N_29751,N_29538);
or UO_1714 (O_1714,N_29598,N_29818);
or UO_1715 (O_1715,N_29471,N_29575);
nor UO_1716 (O_1716,N_29849,N_29870);
nor UO_1717 (O_1717,N_29848,N_29992);
and UO_1718 (O_1718,N_29871,N_29900);
nand UO_1719 (O_1719,N_29557,N_29617);
and UO_1720 (O_1720,N_29731,N_29560);
nor UO_1721 (O_1721,N_29794,N_29689);
and UO_1722 (O_1722,N_29502,N_29711);
or UO_1723 (O_1723,N_29869,N_29679);
nor UO_1724 (O_1724,N_29966,N_29643);
or UO_1725 (O_1725,N_29431,N_29518);
nand UO_1726 (O_1726,N_29762,N_29905);
nor UO_1727 (O_1727,N_29775,N_29621);
or UO_1728 (O_1728,N_29739,N_29781);
nand UO_1729 (O_1729,N_29445,N_29885);
nor UO_1730 (O_1730,N_29783,N_29521);
and UO_1731 (O_1731,N_29513,N_29899);
nand UO_1732 (O_1732,N_29888,N_29910);
and UO_1733 (O_1733,N_29566,N_29660);
or UO_1734 (O_1734,N_29583,N_29507);
or UO_1735 (O_1735,N_29647,N_29608);
or UO_1736 (O_1736,N_29717,N_29583);
xor UO_1737 (O_1737,N_29512,N_29983);
nand UO_1738 (O_1738,N_29943,N_29503);
nor UO_1739 (O_1739,N_29487,N_29434);
or UO_1740 (O_1740,N_29964,N_29430);
nand UO_1741 (O_1741,N_29646,N_29876);
or UO_1742 (O_1742,N_29820,N_29929);
and UO_1743 (O_1743,N_29711,N_29909);
nand UO_1744 (O_1744,N_29460,N_29630);
nand UO_1745 (O_1745,N_29913,N_29501);
nand UO_1746 (O_1746,N_29908,N_29701);
nor UO_1747 (O_1747,N_29904,N_29478);
and UO_1748 (O_1748,N_29567,N_29786);
and UO_1749 (O_1749,N_29824,N_29683);
xnor UO_1750 (O_1750,N_29859,N_29512);
nand UO_1751 (O_1751,N_29898,N_29576);
nand UO_1752 (O_1752,N_29642,N_29686);
nand UO_1753 (O_1753,N_29591,N_29960);
nand UO_1754 (O_1754,N_29688,N_29658);
nand UO_1755 (O_1755,N_29660,N_29948);
nand UO_1756 (O_1756,N_29873,N_29531);
nand UO_1757 (O_1757,N_29978,N_29531);
xor UO_1758 (O_1758,N_29604,N_29612);
nand UO_1759 (O_1759,N_29934,N_29679);
and UO_1760 (O_1760,N_29565,N_29979);
nor UO_1761 (O_1761,N_29945,N_29857);
or UO_1762 (O_1762,N_29475,N_29620);
nor UO_1763 (O_1763,N_29772,N_29421);
and UO_1764 (O_1764,N_29598,N_29924);
or UO_1765 (O_1765,N_29444,N_29569);
or UO_1766 (O_1766,N_29766,N_29403);
or UO_1767 (O_1767,N_29988,N_29715);
and UO_1768 (O_1768,N_29909,N_29704);
nand UO_1769 (O_1769,N_29807,N_29897);
nor UO_1770 (O_1770,N_29546,N_29726);
and UO_1771 (O_1771,N_29562,N_29436);
nor UO_1772 (O_1772,N_29791,N_29444);
xnor UO_1773 (O_1773,N_29959,N_29751);
and UO_1774 (O_1774,N_29599,N_29667);
nand UO_1775 (O_1775,N_29579,N_29462);
and UO_1776 (O_1776,N_29400,N_29500);
nand UO_1777 (O_1777,N_29618,N_29708);
nand UO_1778 (O_1778,N_29697,N_29607);
nor UO_1779 (O_1779,N_29866,N_29511);
or UO_1780 (O_1780,N_29783,N_29837);
or UO_1781 (O_1781,N_29541,N_29401);
and UO_1782 (O_1782,N_29852,N_29521);
and UO_1783 (O_1783,N_29560,N_29495);
or UO_1784 (O_1784,N_29614,N_29845);
nor UO_1785 (O_1785,N_29989,N_29617);
nor UO_1786 (O_1786,N_29502,N_29470);
or UO_1787 (O_1787,N_29511,N_29954);
or UO_1788 (O_1788,N_29493,N_29611);
or UO_1789 (O_1789,N_29939,N_29953);
nor UO_1790 (O_1790,N_29573,N_29919);
nor UO_1791 (O_1791,N_29915,N_29726);
nand UO_1792 (O_1792,N_29415,N_29457);
nor UO_1793 (O_1793,N_29630,N_29572);
nand UO_1794 (O_1794,N_29718,N_29668);
or UO_1795 (O_1795,N_29634,N_29435);
and UO_1796 (O_1796,N_29660,N_29655);
and UO_1797 (O_1797,N_29412,N_29668);
and UO_1798 (O_1798,N_29624,N_29494);
and UO_1799 (O_1799,N_29578,N_29451);
or UO_1800 (O_1800,N_29992,N_29510);
and UO_1801 (O_1801,N_29705,N_29886);
nor UO_1802 (O_1802,N_29621,N_29859);
nand UO_1803 (O_1803,N_29660,N_29864);
nor UO_1804 (O_1804,N_29961,N_29863);
nor UO_1805 (O_1805,N_29849,N_29938);
or UO_1806 (O_1806,N_29927,N_29638);
xor UO_1807 (O_1807,N_29844,N_29482);
nand UO_1808 (O_1808,N_29596,N_29896);
and UO_1809 (O_1809,N_29444,N_29651);
or UO_1810 (O_1810,N_29443,N_29799);
or UO_1811 (O_1811,N_29534,N_29786);
nand UO_1812 (O_1812,N_29505,N_29904);
and UO_1813 (O_1813,N_29996,N_29591);
nand UO_1814 (O_1814,N_29831,N_29684);
and UO_1815 (O_1815,N_29776,N_29841);
nor UO_1816 (O_1816,N_29816,N_29930);
nand UO_1817 (O_1817,N_29528,N_29870);
nor UO_1818 (O_1818,N_29414,N_29849);
or UO_1819 (O_1819,N_29832,N_29548);
or UO_1820 (O_1820,N_29790,N_29869);
nor UO_1821 (O_1821,N_29729,N_29528);
or UO_1822 (O_1822,N_29493,N_29941);
and UO_1823 (O_1823,N_29640,N_29471);
nor UO_1824 (O_1824,N_29746,N_29845);
nor UO_1825 (O_1825,N_29534,N_29618);
nand UO_1826 (O_1826,N_29408,N_29690);
or UO_1827 (O_1827,N_29660,N_29954);
nor UO_1828 (O_1828,N_29732,N_29521);
and UO_1829 (O_1829,N_29685,N_29706);
nand UO_1830 (O_1830,N_29833,N_29430);
or UO_1831 (O_1831,N_29542,N_29974);
and UO_1832 (O_1832,N_29821,N_29753);
nand UO_1833 (O_1833,N_29749,N_29413);
nand UO_1834 (O_1834,N_29839,N_29595);
nor UO_1835 (O_1835,N_29401,N_29565);
or UO_1836 (O_1836,N_29772,N_29933);
nand UO_1837 (O_1837,N_29478,N_29851);
nor UO_1838 (O_1838,N_29480,N_29753);
or UO_1839 (O_1839,N_29872,N_29728);
or UO_1840 (O_1840,N_29985,N_29896);
and UO_1841 (O_1841,N_29743,N_29807);
nand UO_1842 (O_1842,N_29892,N_29506);
xor UO_1843 (O_1843,N_29691,N_29959);
or UO_1844 (O_1844,N_29434,N_29518);
or UO_1845 (O_1845,N_29584,N_29476);
nor UO_1846 (O_1846,N_29705,N_29815);
or UO_1847 (O_1847,N_29826,N_29597);
nor UO_1848 (O_1848,N_29550,N_29693);
and UO_1849 (O_1849,N_29610,N_29500);
or UO_1850 (O_1850,N_29718,N_29933);
or UO_1851 (O_1851,N_29626,N_29684);
and UO_1852 (O_1852,N_29674,N_29706);
or UO_1853 (O_1853,N_29601,N_29463);
nor UO_1854 (O_1854,N_29654,N_29951);
or UO_1855 (O_1855,N_29577,N_29603);
and UO_1856 (O_1856,N_29805,N_29900);
and UO_1857 (O_1857,N_29449,N_29486);
and UO_1858 (O_1858,N_29537,N_29880);
or UO_1859 (O_1859,N_29718,N_29401);
nor UO_1860 (O_1860,N_29473,N_29770);
nand UO_1861 (O_1861,N_29424,N_29674);
nor UO_1862 (O_1862,N_29912,N_29725);
xor UO_1863 (O_1863,N_29813,N_29802);
and UO_1864 (O_1864,N_29707,N_29636);
or UO_1865 (O_1865,N_29468,N_29642);
or UO_1866 (O_1866,N_29840,N_29805);
and UO_1867 (O_1867,N_29751,N_29749);
and UO_1868 (O_1868,N_29532,N_29801);
and UO_1869 (O_1869,N_29426,N_29566);
nand UO_1870 (O_1870,N_29467,N_29832);
or UO_1871 (O_1871,N_29919,N_29808);
or UO_1872 (O_1872,N_29646,N_29694);
and UO_1873 (O_1873,N_29477,N_29878);
nor UO_1874 (O_1874,N_29901,N_29859);
or UO_1875 (O_1875,N_29454,N_29728);
nor UO_1876 (O_1876,N_29952,N_29866);
and UO_1877 (O_1877,N_29799,N_29607);
and UO_1878 (O_1878,N_29988,N_29519);
nand UO_1879 (O_1879,N_29575,N_29726);
and UO_1880 (O_1880,N_29597,N_29966);
and UO_1881 (O_1881,N_29554,N_29609);
xnor UO_1882 (O_1882,N_29413,N_29879);
and UO_1883 (O_1883,N_29999,N_29804);
or UO_1884 (O_1884,N_29658,N_29401);
or UO_1885 (O_1885,N_29982,N_29712);
nand UO_1886 (O_1886,N_29599,N_29708);
and UO_1887 (O_1887,N_29404,N_29756);
nand UO_1888 (O_1888,N_29628,N_29818);
nand UO_1889 (O_1889,N_29431,N_29773);
and UO_1890 (O_1890,N_29585,N_29613);
xor UO_1891 (O_1891,N_29698,N_29640);
nand UO_1892 (O_1892,N_29819,N_29954);
or UO_1893 (O_1893,N_29569,N_29834);
and UO_1894 (O_1894,N_29971,N_29776);
and UO_1895 (O_1895,N_29723,N_29956);
nor UO_1896 (O_1896,N_29835,N_29653);
or UO_1897 (O_1897,N_29636,N_29584);
and UO_1898 (O_1898,N_29666,N_29855);
nand UO_1899 (O_1899,N_29636,N_29478);
nand UO_1900 (O_1900,N_29491,N_29869);
or UO_1901 (O_1901,N_29666,N_29727);
nor UO_1902 (O_1902,N_29407,N_29846);
nand UO_1903 (O_1903,N_29963,N_29459);
nand UO_1904 (O_1904,N_29719,N_29789);
nand UO_1905 (O_1905,N_29678,N_29436);
and UO_1906 (O_1906,N_29750,N_29801);
nor UO_1907 (O_1907,N_29538,N_29915);
or UO_1908 (O_1908,N_29627,N_29423);
or UO_1909 (O_1909,N_29764,N_29411);
or UO_1910 (O_1910,N_29874,N_29798);
and UO_1911 (O_1911,N_29570,N_29776);
or UO_1912 (O_1912,N_29924,N_29978);
nand UO_1913 (O_1913,N_29530,N_29839);
nand UO_1914 (O_1914,N_29402,N_29411);
nor UO_1915 (O_1915,N_29759,N_29416);
nand UO_1916 (O_1916,N_29828,N_29503);
nor UO_1917 (O_1917,N_29892,N_29465);
nand UO_1918 (O_1918,N_29885,N_29407);
and UO_1919 (O_1919,N_29827,N_29618);
nor UO_1920 (O_1920,N_29656,N_29548);
and UO_1921 (O_1921,N_29546,N_29568);
nor UO_1922 (O_1922,N_29888,N_29732);
and UO_1923 (O_1923,N_29487,N_29808);
or UO_1924 (O_1924,N_29663,N_29607);
nor UO_1925 (O_1925,N_29733,N_29670);
nand UO_1926 (O_1926,N_29678,N_29492);
nor UO_1927 (O_1927,N_29912,N_29812);
xor UO_1928 (O_1928,N_29740,N_29858);
nand UO_1929 (O_1929,N_29640,N_29911);
nor UO_1930 (O_1930,N_29493,N_29856);
or UO_1931 (O_1931,N_29801,N_29470);
or UO_1932 (O_1932,N_29886,N_29655);
nor UO_1933 (O_1933,N_29849,N_29532);
nor UO_1934 (O_1934,N_29447,N_29890);
or UO_1935 (O_1935,N_29802,N_29486);
and UO_1936 (O_1936,N_29420,N_29656);
and UO_1937 (O_1937,N_29930,N_29700);
nand UO_1938 (O_1938,N_29828,N_29573);
nand UO_1939 (O_1939,N_29465,N_29539);
nor UO_1940 (O_1940,N_29856,N_29629);
nor UO_1941 (O_1941,N_29565,N_29648);
nand UO_1942 (O_1942,N_29734,N_29634);
and UO_1943 (O_1943,N_29702,N_29806);
or UO_1944 (O_1944,N_29587,N_29884);
and UO_1945 (O_1945,N_29567,N_29650);
nand UO_1946 (O_1946,N_29798,N_29446);
and UO_1947 (O_1947,N_29919,N_29475);
and UO_1948 (O_1948,N_29703,N_29885);
xor UO_1949 (O_1949,N_29721,N_29795);
xor UO_1950 (O_1950,N_29976,N_29411);
nand UO_1951 (O_1951,N_29716,N_29556);
nand UO_1952 (O_1952,N_29898,N_29698);
xor UO_1953 (O_1953,N_29882,N_29806);
or UO_1954 (O_1954,N_29839,N_29562);
nor UO_1955 (O_1955,N_29489,N_29577);
and UO_1956 (O_1956,N_29594,N_29905);
nor UO_1957 (O_1957,N_29732,N_29772);
nand UO_1958 (O_1958,N_29489,N_29678);
and UO_1959 (O_1959,N_29791,N_29694);
nand UO_1960 (O_1960,N_29764,N_29582);
nor UO_1961 (O_1961,N_29971,N_29474);
nor UO_1962 (O_1962,N_29989,N_29402);
nand UO_1963 (O_1963,N_29638,N_29692);
nor UO_1964 (O_1964,N_29403,N_29597);
or UO_1965 (O_1965,N_29694,N_29644);
and UO_1966 (O_1966,N_29512,N_29755);
nand UO_1967 (O_1967,N_29618,N_29596);
and UO_1968 (O_1968,N_29771,N_29597);
and UO_1969 (O_1969,N_29499,N_29457);
nand UO_1970 (O_1970,N_29460,N_29534);
nor UO_1971 (O_1971,N_29439,N_29429);
and UO_1972 (O_1972,N_29500,N_29819);
or UO_1973 (O_1973,N_29400,N_29454);
and UO_1974 (O_1974,N_29464,N_29499);
and UO_1975 (O_1975,N_29676,N_29463);
or UO_1976 (O_1976,N_29561,N_29535);
nor UO_1977 (O_1977,N_29961,N_29570);
nand UO_1978 (O_1978,N_29545,N_29759);
nand UO_1979 (O_1979,N_29821,N_29416);
nand UO_1980 (O_1980,N_29991,N_29564);
nand UO_1981 (O_1981,N_29635,N_29866);
nand UO_1982 (O_1982,N_29672,N_29521);
or UO_1983 (O_1983,N_29752,N_29908);
and UO_1984 (O_1984,N_29705,N_29861);
or UO_1985 (O_1985,N_29411,N_29714);
xor UO_1986 (O_1986,N_29658,N_29662);
nand UO_1987 (O_1987,N_29548,N_29436);
and UO_1988 (O_1988,N_29646,N_29904);
or UO_1989 (O_1989,N_29681,N_29922);
and UO_1990 (O_1990,N_29855,N_29843);
and UO_1991 (O_1991,N_29750,N_29676);
nor UO_1992 (O_1992,N_29974,N_29637);
and UO_1993 (O_1993,N_29857,N_29867);
nor UO_1994 (O_1994,N_29941,N_29994);
or UO_1995 (O_1995,N_29485,N_29421);
nand UO_1996 (O_1996,N_29571,N_29507);
nand UO_1997 (O_1997,N_29505,N_29909);
or UO_1998 (O_1998,N_29753,N_29490);
and UO_1999 (O_1999,N_29531,N_29867);
or UO_2000 (O_2000,N_29630,N_29740);
nor UO_2001 (O_2001,N_29982,N_29859);
nor UO_2002 (O_2002,N_29565,N_29623);
nor UO_2003 (O_2003,N_29644,N_29653);
or UO_2004 (O_2004,N_29644,N_29673);
nand UO_2005 (O_2005,N_29980,N_29704);
nor UO_2006 (O_2006,N_29894,N_29868);
or UO_2007 (O_2007,N_29877,N_29743);
nand UO_2008 (O_2008,N_29953,N_29423);
and UO_2009 (O_2009,N_29485,N_29486);
and UO_2010 (O_2010,N_29811,N_29859);
nand UO_2011 (O_2011,N_29887,N_29413);
nor UO_2012 (O_2012,N_29849,N_29597);
nand UO_2013 (O_2013,N_29508,N_29591);
nand UO_2014 (O_2014,N_29940,N_29876);
nor UO_2015 (O_2015,N_29787,N_29638);
and UO_2016 (O_2016,N_29729,N_29800);
nor UO_2017 (O_2017,N_29502,N_29716);
and UO_2018 (O_2018,N_29531,N_29838);
and UO_2019 (O_2019,N_29602,N_29716);
nor UO_2020 (O_2020,N_29753,N_29529);
nor UO_2021 (O_2021,N_29666,N_29816);
nand UO_2022 (O_2022,N_29723,N_29515);
nor UO_2023 (O_2023,N_29585,N_29405);
nor UO_2024 (O_2024,N_29633,N_29673);
or UO_2025 (O_2025,N_29901,N_29824);
nor UO_2026 (O_2026,N_29877,N_29405);
xor UO_2027 (O_2027,N_29818,N_29666);
and UO_2028 (O_2028,N_29977,N_29414);
or UO_2029 (O_2029,N_29659,N_29405);
nor UO_2030 (O_2030,N_29451,N_29459);
nor UO_2031 (O_2031,N_29511,N_29544);
or UO_2032 (O_2032,N_29854,N_29600);
nor UO_2033 (O_2033,N_29981,N_29666);
nor UO_2034 (O_2034,N_29862,N_29674);
nor UO_2035 (O_2035,N_29785,N_29663);
nand UO_2036 (O_2036,N_29846,N_29804);
nor UO_2037 (O_2037,N_29856,N_29887);
nor UO_2038 (O_2038,N_29982,N_29605);
nand UO_2039 (O_2039,N_29473,N_29816);
nand UO_2040 (O_2040,N_29729,N_29839);
nand UO_2041 (O_2041,N_29683,N_29818);
or UO_2042 (O_2042,N_29962,N_29677);
nor UO_2043 (O_2043,N_29611,N_29523);
nand UO_2044 (O_2044,N_29481,N_29550);
or UO_2045 (O_2045,N_29792,N_29642);
nor UO_2046 (O_2046,N_29452,N_29725);
and UO_2047 (O_2047,N_29485,N_29934);
nor UO_2048 (O_2048,N_29433,N_29523);
nor UO_2049 (O_2049,N_29859,N_29780);
or UO_2050 (O_2050,N_29443,N_29940);
nor UO_2051 (O_2051,N_29836,N_29986);
and UO_2052 (O_2052,N_29836,N_29742);
nor UO_2053 (O_2053,N_29627,N_29885);
nor UO_2054 (O_2054,N_29507,N_29800);
and UO_2055 (O_2055,N_29663,N_29683);
nand UO_2056 (O_2056,N_29534,N_29812);
or UO_2057 (O_2057,N_29576,N_29770);
nor UO_2058 (O_2058,N_29545,N_29903);
nand UO_2059 (O_2059,N_29687,N_29647);
or UO_2060 (O_2060,N_29593,N_29980);
and UO_2061 (O_2061,N_29633,N_29900);
and UO_2062 (O_2062,N_29628,N_29516);
and UO_2063 (O_2063,N_29884,N_29949);
nand UO_2064 (O_2064,N_29504,N_29666);
nor UO_2065 (O_2065,N_29420,N_29573);
nand UO_2066 (O_2066,N_29768,N_29565);
and UO_2067 (O_2067,N_29548,N_29977);
or UO_2068 (O_2068,N_29657,N_29768);
or UO_2069 (O_2069,N_29742,N_29883);
and UO_2070 (O_2070,N_29512,N_29617);
or UO_2071 (O_2071,N_29705,N_29514);
and UO_2072 (O_2072,N_29692,N_29634);
nor UO_2073 (O_2073,N_29801,N_29700);
nor UO_2074 (O_2074,N_29409,N_29417);
and UO_2075 (O_2075,N_29596,N_29878);
or UO_2076 (O_2076,N_29758,N_29455);
or UO_2077 (O_2077,N_29782,N_29754);
nor UO_2078 (O_2078,N_29700,N_29855);
nor UO_2079 (O_2079,N_29492,N_29831);
and UO_2080 (O_2080,N_29511,N_29817);
nand UO_2081 (O_2081,N_29435,N_29683);
nor UO_2082 (O_2082,N_29658,N_29548);
or UO_2083 (O_2083,N_29430,N_29681);
and UO_2084 (O_2084,N_29822,N_29491);
nand UO_2085 (O_2085,N_29952,N_29695);
nor UO_2086 (O_2086,N_29696,N_29409);
xor UO_2087 (O_2087,N_29408,N_29721);
nand UO_2088 (O_2088,N_29664,N_29625);
and UO_2089 (O_2089,N_29418,N_29443);
or UO_2090 (O_2090,N_29565,N_29753);
and UO_2091 (O_2091,N_29500,N_29442);
and UO_2092 (O_2092,N_29686,N_29467);
nor UO_2093 (O_2093,N_29672,N_29850);
nor UO_2094 (O_2094,N_29610,N_29753);
and UO_2095 (O_2095,N_29966,N_29450);
nand UO_2096 (O_2096,N_29570,N_29697);
nor UO_2097 (O_2097,N_29608,N_29533);
nor UO_2098 (O_2098,N_29764,N_29503);
and UO_2099 (O_2099,N_29978,N_29848);
nor UO_2100 (O_2100,N_29927,N_29640);
xnor UO_2101 (O_2101,N_29994,N_29621);
or UO_2102 (O_2102,N_29828,N_29476);
or UO_2103 (O_2103,N_29521,N_29938);
nor UO_2104 (O_2104,N_29454,N_29725);
and UO_2105 (O_2105,N_29981,N_29953);
or UO_2106 (O_2106,N_29828,N_29634);
nor UO_2107 (O_2107,N_29545,N_29990);
nor UO_2108 (O_2108,N_29868,N_29960);
and UO_2109 (O_2109,N_29677,N_29794);
and UO_2110 (O_2110,N_29897,N_29581);
nand UO_2111 (O_2111,N_29945,N_29992);
and UO_2112 (O_2112,N_29982,N_29698);
or UO_2113 (O_2113,N_29753,N_29684);
and UO_2114 (O_2114,N_29791,N_29402);
xor UO_2115 (O_2115,N_29494,N_29467);
and UO_2116 (O_2116,N_29574,N_29589);
or UO_2117 (O_2117,N_29943,N_29853);
nand UO_2118 (O_2118,N_29646,N_29967);
nand UO_2119 (O_2119,N_29792,N_29910);
nand UO_2120 (O_2120,N_29593,N_29767);
nand UO_2121 (O_2121,N_29699,N_29702);
nor UO_2122 (O_2122,N_29713,N_29793);
nor UO_2123 (O_2123,N_29928,N_29800);
nand UO_2124 (O_2124,N_29811,N_29727);
nand UO_2125 (O_2125,N_29980,N_29524);
or UO_2126 (O_2126,N_29929,N_29443);
nor UO_2127 (O_2127,N_29446,N_29953);
nand UO_2128 (O_2128,N_29988,N_29996);
nand UO_2129 (O_2129,N_29465,N_29635);
and UO_2130 (O_2130,N_29857,N_29580);
nor UO_2131 (O_2131,N_29833,N_29528);
nor UO_2132 (O_2132,N_29914,N_29411);
xnor UO_2133 (O_2133,N_29809,N_29756);
nor UO_2134 (O_2134,N_29693,N_29419);
nor UO_2135 (O_2135,N_29474,N_29903);
nand UO_2136 (O_2136,N_29893,N_29872);
nor UO_2137 (O_2137,N_29465,N_29851);
nand UO_2138 (O_2138,N_29596,N_29601);
and UO_2139 (O_2139,N_29654,N_29984);
or UO_2140 (O_2140,N_29400,N_29713);
nand UO_2141 (O_2141,N_29863,N_29755);
and UO_2142 (O_2142,N_29803,N_29480);
or UO_2143 (O_2143,N_29425,N_29430);
nor UO_2144 (O_2144,N_29717,N_29454);
nand UO_2145 (O_2145,N_29489,N_29979);
and UO_2146 (O_2146,N_29934,N_29971);
nand UO_2147 (O_2147,N_29851,N_29492);
and UO_2148 (O_2148,N_29476,N_29419);
xnor UO_2149 (O_2149,N_29756,N_29726);
or UO_2150 (O_2150,N_29622,N_29889);
nor UO_2151 (O_2151,N_29954,N_29408);
and UO_2152 (O_2152,N_29603,N_29608);
nand UO_2153 (O_2153,N_29408,N_29678);
or UO_2154 (O_2154,N_29590,N_29576);
nand UO_2155 (O_2155,N_29933,N_29406);
nor UO_2156 (O_2156,N_29764,N_29445);
and UO_2157 (O_2157,N_29900,N_29916);
nand UO_2158 (O_2158,N_29953,N_29688);
nand UO_2159 (O_2159,N_29803,N_29607);
nand UO_2160 (O_2160,N_29822,N_29507);
nor UO_2161 (O_2161,N_29740,N_29594);
and UO_2162 (O_2162,N_29685,N_29855);
nand UO_2163 (O_2163,N_29951,N_29833);
or UO_2164 (O_2164,N_29566,N_29538);
and UO_2165 (O_2165,N_29603,N_29973);
and UO_2166 (O_2166,N_29495,N_29840);
and UO_2167 (O_2167,N_29908,N_29578);
nand UO_2168 (O_2168,N_29840,N_29936);
and UO_2169 (O_2169,N_29635,N_29410);
and UO_2170 (O_2170,N_29818,N_29939);
and UO_2171 (O_2171,N_29752,N_29418);
nor UO_2172 (O_2172,N_29524,N_29599);
or UO_2173 (O_2173,N_29421,N_29962);
nor UO_2174 (O_2174,N_29530,N_29610);
nand UO_2175 (O_2175,N_29685,N_29676);
and UO_2176 (O_2176,N_29908,N_29635);
and UO_2177 (O_2177,N_29753,N_29696);
nor UO_2178 (O_2178,N_29899,N_29675);
nand UO_2179 (O_2179,N_29649,N_29985);
xor UO_2180 (O_2180,N_29654,N_29405);
and UO_2181 (O_2181,N_29766,N_29844);
nor UO_2182 (O_2182,N_29473,N_29942);
nor UO_2183 (O_2183,N_29849,N_29787);
nor UO_2184 (O_2184,N_29406,N_29616);
nor UO_2185 (O_2185,N_29831,N_29915);
nand UO_2186 (O_2186,N_29533,N_29516);
nor UO_2187 (O_2187,N_29511,N_29939);
nor UO_2188 (O_2188,N_29918,N_29512);
nor UO_2189 (O_2189,N_29722,N_29582);
nor UO_2190 (O_2190,N_29838,N_29489);
and UO_2191 (O_2191,N_29925,N_29555);
nand UO_2192 (O_2192,N_29519,N_29511);
nand UO_2193 (O_2193,N_29913,N_29672);
nor UO_2194 (O_2194,N_29866,N_29520);
and UO_2195 (O_2195,N_29804,N_29559);
xnor UO_2196 (O_2196,N_29974,N_29778);
nand UO_2197 (O_2197,N_29626,N_29411);
or UO_2198 (O_2198,N_29678,N_29993);
and UO_2199 (O_2199,N_29413,N_29756);
and UO_2200 (O_2200,N_29465,N_29671);
and UO_2201 (O_2201,N_29929,N_29622);
nand UO_2202 (O_2202,N_29535,N_29713);
and UO_2203 (O_2203,N_29769,N_29645);
and UO_2204 (O_2204,N_29545,N_29707);
or UO_2205 (O_2205,N_29850,N_29999);
nand UO_2206 (O_2206,N_29920,N_29921);
nand UO_2207 (O_2207,N_29857,N_29633);
nand UO_2208 (O_2208,N_29484,N_29840);
or UO_2209 (O_2209,N_29810,N_29676);
or UO_2210 (O_2210,N_29512,N_29820);
or UO_2211 (O_2211,N_29647,N_29968);
nand UO_2212 (O_2212,N_29993,N_29581);
and UO_2213 (O_2213,N_29951,N_29818);
nor UO_2214 (O_2214,N_29810,N_29444);
and UO_2215 (O_2215,N_29988,N_29576);
nand UO_2216 (O_2216,N_29722,N_29573);
or UO_2217 (O_2217,N_29772,N_29790);
nand UO_2218 (O_2218,N_29870,N_29995);
or UO_2219 (O_2219,N_29508,N_29854);
nor UO_2220 (O_2220,N_29702,N_29499);
nand UO_2221 (O_2221,N_29642,N_29636);
nand UO_2222 (O_2222,N_29605,N_29514);
and UO_2223 (O_2223,N_29650,N_29912);
and UO_2224 (O_2224,N_29655,N_29836);
nand UO_2225 (O_2225,N_29715,N_29856);
and UO_2226 (O_2226,N_29884,N_29797);
nor UO_2227 (O_2227,N_29918,N_29450);
or UO_2228 (O_2228,N_29854,N_29805);
nor UO_2229 (O_2229,N_29561,N_29795);
or UO_2230 (O_2230,N_29553,N_29640);
or UO_2231 (O_2231,N_29803,N_29682);
or UO_2232 (O_2232,N_29548,N_29461);
or UO_2233 (O_2233,N_29948,N_29609);
and UO_2234 (O_2234,N_29706,N_29799);
or UO_2235 (O_2235,N_29461,N_29457);
nand UO_2236 (O_2236,N_29558,N_29602);
xnor UO_2237 (O_2237,N_29697,N_29478);
nor UO_2238 (O_2238,N_29731,N_29868);
or UO_2239 (O_2239,N_29664,N_29918);
and UO_2240 (O_2240,N_29627,N_29549);
and UO_2241 (O_2241,N_29461,N_29947);
or UO_2242 (O_2242,N_29981,N_29920);
or UO_2243 (O_2243,N_29434,N_29553);
xnor UO_2244 (O_2244,N_29762,N_29755);
xnor UO_2245 (O_2245,N_29805,N_29451);
or UO_2246 (O_2246,N_29837,N_29971);
nand UO_2247 (O_2247,N_29868,N_29836);
and UO_2248 (O_2248,N_29878,N_29920);
and UO_2249 (O_2249,N_29510,N_29923);
and UO_2250 (O_2250,N_29569,N_29866);
or UO_2251 (O_2251,N_29862,N_29602);
or UO_2252 (O_2252,N_29486,N_29834);
nor UO_2253 (O_2253,N_29649,N_29887);
nand UO_2254 (O_2254,N_29615,N_29610);
or UO_2255 (O_2255,N_29840,N_29769);
nor UO_2256 (O_2256,N_29761,N_29697);
nand UO_2257 (O_2257,N_29641,N_29649);
and UO_2258 (O_2258,N_29540,N_29554);
or UO_2259 (O_2259,N_29814,N_29538);
and UO_2260 (O_2260,N_29920,N_29709);
or UO_2261 (O_2261,N_29749,N_29709);
and UO_2262 (O_2262,N_29818,N_29480);
nor UO_2263 (O_2263,N_29529,N_29716);
or UO_2264 (O_2264,N_29685,N_29561);
or UO_2265 (O_2265,N_29716,N_29430);
nor UO_2266 (O_2266,N_29817,N_29696);
nand UO_2267 (O_2267,N_29811,N_29813);
nor UO_2268 (O_2268,N_29895,N_29456);
nor UO_2269 (O_2269,N_29593,N_29993);
xnor UO_2270 (O_2270,N_29513,N_29798);
and UO_2271 (O_2271,N_29947,N_29689);
and UO_2272 (O_2272,N_29927,N_29406);
and UO_2273 (O_2273,N_29465,N_29804);
or UO_2274 (O_2274,N_29471,N_29904);
nor UO_2275 (O_2275,N_29427,N_29632);
nor UO_2276 (O_2276,N_29661,N_29742);
and UO_2277 (O_2277,N_29716,N_29933);
xor UO_2278 (O_2278,N_29437,N_29502);
nor UO_2279 (O_2279,N_29927,N_29786);
or UO_2280 (O_2280,N_29809,N_29805);
nand UO_2281 (O_2281,N_29475,N_29854);
and UO_2282 (O_2282,N_29679,N_29590);
nor UO_2283 (O_2283,N_29713,N_29883);
or UO_2284 (O_2284,N_29905,N_29736);
or UO_2285 (O_2285,N_29754,N_29568);
nor UO_2286 (O_2286,N_29758,N_29671);
nand UO_2287 (O_2287,N_29739,N_29831);
nor UO_2288 (O_2288,N_29580,N_29453);
or UO_2289 (O_2289,N_29899,N_29796);
or UO_2290 (O_2290,N_29801,N_29885);
or UO_2291 (O_2291,N_29874,N_29977);
or UO_2292 (O_2292,N_29586,N_29780);
nand UO_2293 (O_2293,N_29795,N_29892);
nor UO_2294 (O_2294,N_29973,N_29794);
or UO_2295 (O_2295,N_29586,N_29643);
nor UO_2296 (O_2296,N_29539,N_29801);
nand UO_2297 (O_2297,N_29858,N_29729);
and UO_2298 (O_2298,N_29668,N_29839);
and UO_2299 (O_2299,N_29851,N_29533);
nand UO_2300 (O_2300,N_29973,N_29777);
and UO_2301 (O_2301,N_29978,N_29872);
or UO_2302 (O_2302,N_29623,N_29510);
or UO_2303 (O_2303,N_29862,N_29512);
nand UO_2304 (O_2304,N_29721,N_29697);
and UO_2305 (O_2305,N_29595,N_29986);
nand UO_2306 (O_2306,N_29449,N_29633);
nor UO_2307 (O_2307,N_29615,N_29635);
nor UO_2308 (O_2308,N_29953,N_29740);
nand UO_2309 (O_2309,N_29827,N_29452);
or UO_2310 (O_2310,N_29636,N_29646);
nor UO_2311 (O_2311,N_29452,N_29978);
nand UO_2312 (O_2312,N_29863,N_29978);
nor UO_2313 (O_2313,N_29608,N_29542);
nand UO_2314 (O_2314,N_29998,N_29740);
nand UO_2315 (O_2315,N_29738,N_29944);
or UO_2316 (O_2316,N_29597,N_29706);
or UO_2317 (O_2317,N_29929,N_29891);
nand UO_2318 (O_2318,N_29874,N_29431);
and UO_2319 (O_2319,N_29512,N_29961);
nor UO_2320 (O_2320,N_29537,N_29422);
or UO_2321 (O_2321,N_29705,N_29647);
or UO_2322 (O_2322,N_29569,N_29621);
and UO_2323 (O_2323,N_29993,N_29942);
nand UO_2324 (O_2324,N_29943,N_29992);
nor UO_2325 (O_2325,N_29488,N_29787);
nand UO_2326 (O_2326,N_29978,N_29773);
or UO_2327 (O_2327,N_29781,N_29582);
or UO_2328 (O_2328,N_29918,N_29808);
nand UO_2329 (O_2329,N_29486,N_29496);
nor UO_2330 (O_2330,N_29851,N_29436);
or UO_2331 (O_2331,N_29713,N_29402);
or UO_2332 (O_2332,N_29412,N_29596);
or UO_2333 (O_2333,N_29882,N_29481);
or UO_2334 (O_2334,N_29521,N_29849);
nor UO_2335 (O_2335,N_29412,N_29479);
nor UO_2336 (O_2336,N_29963,N_29654);
nor UO_2337 (O_2337,N_29466,N_29675);
nor UO_2338 (O_2338,N_29850,N_29929);
or UO_2339 (O_2339,N_29982,N_29512);
nand UO_2340 (O_2340,N_29963,N_29447);
nor UO_2341 (O_2341,N_29614,N_29581);
and UO_2342 (O_2342,N_29735,N_29530);
or UO_2343 (O_2343,N_29705,N_29594);
xor UO_2344 (O_2344,N_29944,N_29943);
and UO_2345 (O_2345,N_29444,N_29679);
nand UO_2346 (O_2346,N_29466,N_29886);
and UO_2347 (O_2347,N_29839,N_29401);
or UO_2348 (O_2348,N_29692,N_29968);
nor UO_2349 (O_2349,N_29413,N_29926);
or UO_2350 (O_2350,N_29709,N_29959);
nor UO_2351 (O_2351,N_29605,N_29792);
or UO_2352 (O_2352,N_29481,N_29754);
and UO_2353 (O_2353,N_29512,N_29737);
nand UO_2354 (O_2354,N_29688,N_29414);
xnor UO_2355 (O_2355,N_29621,N_29438);
nand UO_2356 (O_2356,N_29490,N_29412);
nor UO_2357 (O_2357,N_29908,N_29678);
or UO_2358 (O_2358,N_29851,N_29461);
nand UO_2359 (O_2359,N_29775,N_29460);
nand UO_2360 (O_2360,N_29757,N_29789);
nand UO_2361 (O_2361,N_29569,N_29489);
or UO_2362 (O_2362,N_29577,N_29644);
nand UO_2363 (O_2363,N_29795,N_29568);
nor UO_2364 (O_2364,N_29774,N_29856);
nand UO_2365 (O_2365,N_29494,N_29979);
or UO_2366 (O_2366,N_29584,N_29970);
nand UO_2367 (O_2367,N_29565,N_29985);
nor UO_2368 (O_2368,N_29594,N_29734);
nor UO_2369 (O_2369,N_29986,N_29902);
or UO_2370 (O_2370,N_29792,N_29816);
or UO_2371 (O_2371,N_29561,N_29898);
nand UO_2372 (O_2372,N_29744,N_29943);
and UO_2373 (O_2373,N_29772,N_29689);
and UO_2374 (O_2374,N_29570,N_29617);
or UO_2375 (O_2375,N_29406,N_29485);
and UO_2376 (O_2376,N_29703,N_29850);
or UO_2377 (O_2377,N_29939,N_29743);
or UO_2378 (O_2378,N_29652,N_29935);
and UO_2379 (O_2379,N_29673,N_29831);
or UO_2380 (O_2380,N_29975,N_29426);
nor UO_2381 (O_2381,N_29742,N_29640);
xnor UO_2382 (O_2382,N_29722,N_29947);
nand UO_2383 (O_2383,N_29532,N_29606);
nand UO_2384 (O_2384,N_29882,N_29568);
and UO_2385 (O_2385,N_29686,N_29451);
and UO_2386 (O_2386,N_29479,N_29696);
or UO_2387 (O_2387,N_29470,N_29917);
nor UO_2388 (O_2388,N_29507,N_29989);
and UO_2389 (O_2389,N_29544,N_29640);
xor UO_2390 (O_2390,N_29907,N_29449);
nand UO_2391 (O_2391,N_29724,N_29537);
or UO_2392 (O_2392,N_29948,N_29997);
or UO_2393 (O_2393,N_29997,N_29899);
nor UO_2394 (O_2394,N_29785,N_29480);
or UO_2395 (O_2395,N_29864,N_29688);
nand UO_2396 (O_2396,N_29537,N_29768);
or UO_2397 (O_2397,N_29692,N_29945);
or UO_2398 (O_2398,N_29469,N_29658);
or UO_2399 (O_2399,N_29411,N_29913);
and UO_2400 (O_2400,N_29820,N_29815);
or UO_2401 (O_2401,N_29726,N_29584);
nor UO_2402 (O_2402,N_29672,N_29422);
nand UO_2403 (O_2403,N_29845,N_29457);
nor UO_2404 (O_2404,N_29798,N_29617);
nand UO_2405 (O_2405,N_29706,N_29475);
or UO_2406 (O_2406,N_29723,N_29894);
nand UO_2407 (O_2407,N_29659,N_29720);
and UO_2408 (O_2408,N_29471,N_29793);
nor UO_2409 (O_2409,N_29819,N_29715);
and UO_2410 (O_2410,N_29672,N_29998);
nand UO_2411 (O_2411,N_29847,N_29821);
or UO_2412 (O_2412,N_29992,N_29740);
nand UO_2413 (O_2413,N_29891,N_29903);
nand UO_2414 (O_2414,N_29737,N_29532);
nand UO_2415 (O_2415,N_29624,N_29596);
or UO_2416 (O_2416,N_29686,N_29493);
nor UO_2417 (O_2417,N_29562,N_29485);
nand UO_2418 (O_2418,N_29850,N_29650);
and UO_2419 (O_2419,N_29581,N_29629);
nand UO_2420 (O_2420,N_29982,N_29564);
nand UO_2421 (O_2421,N_29714,N_29967);
nand UO_2422 (O_2422,N_29748,N_29933);
nor UO_2423 (O_2423,N_29445,N_29424);
or UO_2424 (O_2424,N_29981,N_29587);
nand UO_2425 (O_2425,N_29953,N_29577);
or UO_2426 (O_2426,N_29570,N_29651);
and UO_2427 (O_2427,N_29923,N_29951);
nor UO_2428 (O_2428,N_29927,N_29547);
nor UO_2429 (O_2429,N_29743,N_29721);
nor UO_2430 (O_2430,N_29792,N_29772);
and UO_2431 (O_2431,N_29559,N_29691);
nand UO_2432 (O_2432,N_29594,N_29915);
and UO_2433 (O_2433,N_29641,N_29891);
or UO_2434 (O_2434,N_29513,N_29696);
nand UO_2435 (O_2435,N_29591,N_29692);
xnor UO_2436 (O_2436,N_29535,N_29487);
or UO_2437 (O_2437,N_29986,N_29848);
or UO_2438 (O_2438,N_29824,N_29755);
and UO_2439 (O_2439,N_29899,N_29505);
nor UO_2440 (O_2440,N_29930,N_29657);
nor UO_2441 (O_2441,N_29729,N_29807);
nand UO_2442 (O_2442,N_29827,N_29628);
nor UO_2443 (O_2443,N_29530,N_29905);
or UO_2444 (O_2444,N_29793,N_29791);
or UO_2445 (O_2445,N_29926,N_29961);
nand UO_2446 (O_2446,N_29529,N_29543);
or UO_2447 (O_2447,N_29824,N_29449);
or UO_2448 (O_2448,N_29565,N_29627);
nor UO_2449 (O_2449,N_29549,N_29750);
or UO_2450 (O_2450,N_29526,N_29694);
nor UO_2451 (O_2451,N_29552,N_29763);
nor UO_2452 (O_2452,N_29441,N_29506);
xor UO_2453 (O_2453,N_29613,N_29527);
or UO_2454 (O_2454,N_29501,N_29504);
or UO_2455 (O_2455,N_29994,N_29630);
nor UO_2456 (O_2456,N_29986,N_29679);
and UO_2457 (O_2457,N_29810,N_29819);
nor UO_2458 (O_2458,N_29972,N_29403);
or UO_2459 (O_2459,N_29626,N_29905);
nand UO_2460 (O_2460,N_29518,N_29421);
and UO_2461 (O_2461,N_29553,N_29432);
and UO_2462 (O_2462,N_29486,N_29487);
or UO_2463 (O_2463,N_29895,N_29957);
nor UO_2464 (O_2464,N_29727,N_29763);
and UO_2465 (O_2465,N_29663,N_29889);
xor UO_2466 (O_2466,N_29907,N_29877);
and UO_2467 (O_2467,N_29594,N_29818);
and UO_2468 (O_2468,N_29618,N_29467);
and UO_2469 (O_2469,N_29988,N_29918);
or UO_2470 (O_2470,N_29956,N_29661);
or UO_2471 (O_2471,N_29585,N_29664);
nor UO_2472 (O_2472,N_29843,N_29768);
and UO_2473 (O_2473,N_29802,N_29901);
nor UO_2474 (O_2474,N_29969,N_29612);
nand UO_2475 (O_2475,N_29729,N_29923);
nand UO_2476 (O_2476,N_29519,N_29852);
and UO_2477 (O_2477,N_29583,N_29804);
and UO_2478 (O_2478,N_29512,N_29865);
nand UO_2479 (O_2479,N_29518,N_29812);
nor UO_2480 (O_2480,N_29628,N_29555);
nand UO_2481 (O_2481,N_29622,N_29661);
nand UO_2482 (O_2482,N_29929,N_29405);
and UO_2483 (O_2483,N_29601,N_29949);
nor UO_2484 (O_2484,N_29962,N_29764);
or UO_2485 (O_2485,N_29772,N_29679);
nor UO_2486 (O_2486,N_29476,N_29657);
xnor UO_2487 (O_2487,N_29819,N_29879);
nor UO_2488 (O_2488,N_29881,N_29845);
nor UO_2489 (O_2489,N_29454,N_29898);
or UO_2490 (O_2490,N_29990,N_29907);
nand UO_2491 (O_2491,N_29685,N_29562);
or UO_2492 (O_2492,N_29425,N_29612);
nand UO_2493 (O_2493,N_29927,N_29743);
nand UO_2494 (O_2494,N_29884,N_29625);
or UO_2495 (O_2495,N_29888,N_29718);
and UO_2496 (O_2496,N_29457,N_29745);
nand UO_2497 (O_2497,N_29861,N_29912);
nand UO_2498 (O_2498,N_29914,N_29624);
or UO_2499 (O_2499,N_29855,N_29510);
nor UO_2500 (O_2500,N_29853,N_29935);
nand UO_2501 (O_2501,N_29570,N_29467);
and UO_2502 (O_2502,N_29877,N_29542);
and UO_2503 (O_2503,N_29679,N_29705);
and UO_2504 (O_2504,N_29968,N_29655);
nor UO_2505 (O_2505,N_29482,N_29653);
nor UO_2506 (O_2506,N_29914,N_29534);
and UO_2507 (O_2507,N_29738,N_29947);
nor UO_2508 (O_2508,N_29547,N_29471);
nand UO_2509 (O_2509,N_29674,N_29490);
or UO_2510 (O_2510,N_29743,N_29889);
or UO_2511 (O_2511,N_29568,N_29800);
nor UO_2512 (O_2512,N_29426,N_29729);
nor UO_2513 (O_2513,N_29693,N_29819);
and UO_2514 (O_2514,N_29646,N_29419);
and UO_2515 (O_2515,N_29743,N_29573);
nor UO_2516 (O_2516,N_29563,N_29410);
nand UO_2517 (O_2517,N_29436,N_29933);
nand UO_2518 (O_2518,N_29561,N_29693);
or UO_2519 (O_2519,N_29471,N_29818);
and UO_2520 (O_2520,N_29452,N_29491);
or UO_2521 (O_2521,N_29484,N_29812);
nand UO_2522 (O_2522,N_29536,N_29417);
nor UO_2523 (O_2523,N_29668,N_29938);
or UO_2524 (O_2524,N_29926,N_29441);
and UO_2525 (O_2525,N_29564,N_29631);
nand UO_2526 (O_2526,N_29723,N_29445);
or UO_2527 (O_2527,N_29622,N_29648);
nand UO_2528 (O_2528,N_29531,N_29762);
or UO_2529 (O_2529,N_29881,N_29900);
or UO_2530 (O_2530,N_29848,N_29801);
or UO_2531 (O_2531,N_29673,N_29596);
or UO_2532 (O_2532,N_29433,N_29681);
and UO_2533 (O_2533,N_29874,N_29526);
or UO_2534 (O_2534,N_29670,N_29589);
nand UO_2535 (O_2535,N_29570,N_29848);
nand UO_2536 (O_2536,N_29949,N_29794);
and UO_2537 (O_2537,N_29904,N_29927);
or UO_2538 (O_2538,N_29986,N_29541);
or UO_2539 (O_2539,N_29959,N_29582);
nor UO_2540 (O_2540,N_29983,N_29571);
and UO_2541 (O_2541,N_29466,N_29494);
nor UO_2542 (O_2542,N_29618,N_29635);
nor UO_2543 (O_2543,N_29567,N_29477);
or UO_2544 (O_2544,N_29435,N_29800);
and UO_2545 (O_2545,N_29506,N_29512);
nor UO_2546 (O_2546,N_29474,N_29524);
nor UO_2547 (O_2547,N_29407,N_29466);
and UO_2548 (O_2548,N_29731,N_29925);
nand UO_2549 (O_2549,N_29674,N_29517);
nand UO_2550 (O_2550,N_29930,N_29953);
or UO_2551 (O_2551,N_29926,N_29891);
nand UO_2552 (O_2552,N_29631,N_29890);
or UO_2553 (O_2553,N_29624,N_29756);
nor UO_2554 (O_2554,N_29477,N_29776);
and UO_2555 (O_2555,N_29873,N_29855);
and UO_2556 (O_2556,N_29605,N_29567);
or UO_2557 (O_2557,N_29424,N_29615);
nor UO_2558 (O_2558,N_29551,N_29617);
nor UO_2559 (O_2559,N_29483,N_29626);
or UO_2560 (O_2560,N_29818,N_29499);
and UO_2561 (O_2561,N_29573,N_29598);
and UO_2562 (O_2562,N_29879,N_29690);
nand UO_2563 (O_2563,N_29966,N_29725);
and UO_2564 (O_2564,N_29953,N_29562);
nand UO_2565 (O_2565,N_29612,N_29719);
nand UO_2566 (O_2566,N_29894,N_29708);
nand UO_2567 (O_2567,N_29469,N_29405);
nand UO_2568 (O_2568,N_29523,N_29898);
nor UO_2569 (O_2569,N_29767,N_29976);
or UO_2570 (O_2570,N_29953,N_29420);
or UO_2571 (O_2571,N_29447,N_29800);
nor UO_2572 (O_2572,N_29765,N_29656);
nor UO_2573 (O_2573,N_29507,N_29778);
nand UO_2574 (O_2574,N_29919,N_29453);
and UO_2575 (O_2575,N_29804,N_29678);
nand UO_2576 (O_2576,N_29538,N_29516);
or UO_2577 (O_2577,N_29572,N_29742);
or UO_2578 (O_2578,N_29516,N_29949);
or UO_2579 (O_2579,N_29893,N_29704);
or UO_2580 (O_2580,N_29553,N_29510);
and UO_2581 (O_2581,N_29590,N_29535);
or UO_2582 (O_2582,N_29873,N_29403);
or UO_2583 (O_2583,N_29632,N_29922);
nand UO_2584 (O_2584,N_29970,N_29932);
or UO_2585 (O_2585,N_29866,N_29674);
and UO_2586 (O_2586,N_29848,N_29837);
or UO_2587 (O_2587,N_29410,N_29402);
and UO_2588 (O_2588,N_29897,N_29987);
and UO_2589 (O_2589,N_29560,N_29956);
and UO_2590 (O_2590,N_29732,N_29853);
or UO_2591 (O_2591,N_29770,N_29685);
or UO_2592 (O_2592,N_29521,N_29715);
nor UO_2593 (O_2593,N_29765,N_29818);
and UO_2594 (O_2594,N_29981,N_29601);
and UO_2595 (O_2595,N_29798,N_29564);
nand UO_2596 (O_2596,N_29877,N_29982);
and UO_2597 (O_2597,N_29738,N_29532);
nor UO_2598 (O_2598,N_29791,N_29569);
and UO_2599 (O_2599,N_29658,N_29613);
nor UO_2600 (O_2600,N_29615,N_29476);
nor UO_2601 (O_2601,N_29465,N_29843);
nand UO_2602 (O_2602,N_29989,N_29978);
or UO_2603 (O_2603,N_29954,N_29642);
or UO_2604 (O_2604,N_29702,N_29444);
nand UO_2605 (O_2605,N_29995,N_29674);
or UO_2606 (O_2606,N_29706,N_29717);
or UO_2607 (O_2607,N_29984,N_29785);
or UO_2608 (O_2608,N_29985,N_29921);
nor UO_2609 (O_2609,N_29599,N_29601);
nand UO_2610 (O_2610,N_29712,N_29680);
and UO_2611 (O_2611,N_29996,N_29970);
nor UO_2612 (O_2612,N_29730,N_29751);
nor UO_2613 (O_2613,N_29858,N_29577);
or UO_2614 (O_2614,N_29959,N_29889);
nand UO_2615 (O_2615,N_29466,N_29728);
and UO_2616 (O_2616,N_29791,N_29918);
and UO_2617 (O_2617,N_29741,N_29591);
nand UO_2618 (O_2618,N_29489,N_29869);
nor UO_2619 (O_2619,N_29639,N_29569);
nand UO_2620 (O_2620,N_29982,N_29503);
nand UO_2621 (O_2621,N_29525,N_29739);
or UO_2622 (O_2622,N_29619,N_29421);
and UO_2623 (O_2623,N_29679,N_29463);
or UO_2624 (O_2624,N_29952,N_29996);
and UO_2625 (O_2625,N_29984,N_29705);
nand UO_2626 (O_2626,N_29710,N_29424);
and UO_2627 (O_2627,N_29599,N_29933);
or UO_2628 (O_2628,N_29583,N_29601);
or UO_2629 (O_2629,N_29880,N_29732);
or UO_2630 (O_2630,N_29827,N_29528);
nor UO_2631 (O_2631,N_29577,N_29815);
nand UO_2632 (O_2632,N_29686,N_29990);
and UO_2633 (O_2633,N_29585,N_29944);
nand UO_2634 (O_2634,N_29948,N_29831);
nand UO_2635 (O_2635,N_29801,N_29811);
nor UO_2636 (O_2636,N_29716,N_29500);
and UO_2637 (O_2637,N_29933,N_29952);
or UO_2638 (O_2638,N_29553,N_29823);
nand UO_2639 (O_2639,N_29999,N_29685);
and UO_2640 (O_2640,N_29473,N_29767);
nand UO_2641 (O_2641,N_29777,N_29413);
nand UO_2642 (O_2642,N_29502,N_29866);
nor UO_2643 (O_2643,N_29820,N_29582);
nor UO_2644 (O_2644,N_29492,N_29547);
or UO_2645 (O_2645,N_29597,N_29958);
or UO_2646 (O_2646,N_29594,N_29809);
nor UO_2647 (O_2647,N_29649,N_29875);
and UO_2648 (O_2648,N_29596,N_29641);
and UO_2649 (O_2649,N_29499,N_29671);
or UO_2650 (O_2650,N_29649,N_29726);
or UO_2651 (O_2651,N_29913,N_29715);
or UO_2652 (O_2652,N_29467,N_29584);
and UO_2653 (O_2653,N_29707,N_29848);
and UO_2654 (O_2654,N_29401,N_29664);
or UO_2655 (O_2655,N_29635,N_29895);
and UO_2656 (O_2656,N_29584,N_29600);
nor UO_2657 (O_2657,N_29890,N_29442);
xnor UO_2658 (O_2658,N_29756,N_29676);
or UO_2659 (O_2659,N_29757,N_29976);
and UO_2660 (O_2660,N_29714,N_29424);
or UO_2661 (O_2661,N_29973,N_29718);
and UO_2662 (O_2662,N_29881,N_29899);
and UO_2663 (O_2663,N_29776,N_29666);
and UO_2664 (O_2664,N_29414,N_29893);
nor UO_2665 (O_2665,N_29823,N_29466);
and UO_2666 (O_2666,N_29827,N_29457);
or UO_2667 (O_2667,N_29475,N_29469);
and UO_2668 (O_2668,N_29827,N_29973);
or UO_2669 (O_2669,N_29905,N_29843);
xor UO_2670 (O_2670,N_29815,N_29974);
nor UO_2671 (O_2671,N_29882,N_29732);
and UO_2672 (O_2672,N_29577,N_29445);
nand UO_2673 (O_2673,N_29874,N_29827);
nand UO_2674 (O_2674,N_29693,N_29463);
or UO_2675 (O_2675,N_29475,N_29983);
or UO_2676 (O_2676,N_29978,N_29528);
nand UO_2677 (O_2677,N_29425,N_29400);
xnor UO_2678 (O_2678,N_29780,N_29749);
nand UO_2679 (O_2679,N_29408,N_29785);
nand UO_2680 (O_2680,N_29447,N_29682);
nand UO_2681 (O_2681,N_29755,N_29820);
nand UO_2682 (O_2682,N_29613,N_29596);
or UO_2683 (O_2683,N_29465,N_29720);
nor UO_2684 (O_2684,N_29516,N_29736);
nand UO_2685 (O_2685,N_29618,N_29996);
nand UO_2686 (O_2686,N_29822,N_29454);
nand UO_2687 (O_2687,N_29872,N_29863);
or UO_2688 (O_2688,N_29908,N_29428);
nand UO_2689 (O_2689,N_29670,N_29835);
nand UO_2690 (O_2690,N_29617,N_29820);
nor UO_2691 (O_2691,N_29431,N_29883);
nand UO_2692 (O_2692,N_29914,N_29451);
nand UO_2693 (O_2693,N_29820,N_29663);
nor UO_2694 (O_2694,N_29633,N_29623);
nor UO_2695 (O_2695,N_29855,N_29681);
or UO_2696 (O_2696,N_29704,N_29755);
nand UO_2697 (O_2697,N_29687,N_29965);
and UO_2698 (O_2698,N_29428,N_29981);
nor UO_2699 (O_2699,N_29966,N_29614);
nor UO_2700 (O_2700,N_29823,N_29402);
and UO_2701 (O_2701,N_29452,N_29586);
nor UO_2702 (O_2702,N_29536,N_29641);
nor UO_2703 (O_2703,N_29997,N_29764);
or UO_2704 (O_2704,N_29796,N_29674);
nor UO_2705 (O_2705,N_29689,N_29473);
and UO_2706 (O_2706,N_29717,N_29549);
nor UO_2707 (O_2707,N_29799,N_29904);
or UO_2708 (O_2708,N_29454,N_29500);
nor UO_2709 (O_2709,N_29749,N_29902);
nor UO_2710 (O_2710,N_29534,N_29543);
nand UO_2711 (O_2711,N_29883,N_29503);
xor UO_2712 (O_2712,N_29888,N_29717);
or UO_2713 (O_2713,N_29989,N_29830);
or UO_2714 (O_2714,N_29662,N_29616);
nor UO_2715 (O_2715,N_29911,N_29930);
nor UO_2716 (O_2716,N_29587,N_29524);
and UO_2717 (O_2717,N_29760,N_29986);
nand UO_2718 (O_2718,N_29793,N_29858);
nand UO_2719 (O_2719,N_29914,N_29540);
nand UO_2720 (O_2720,N_29602,N_29539);
and UO_2721 (O_2721,N_29940,N_29847);
nor UO_2722 (O_2722,N_29772,N_29894);
and UO_2723 (O_2723,N_29845,N_29630);
nor UO_2724 (O_2724,N_29642,N_29595);
nor UO_2725 (O_2725,N_29989,N_29898);
nand UO_2726 (O_2726,N_29913,N_29678);
and UO_2727 (O_2727,N_29810,N_29797);
xor UO_2728 (O_2728,N_29996,N_29542);
or UO_2729 (O_2729,N_29463,N_29719);
or UO_2730 (O_2730,N_29484,N_29965);
nand UO_2731 (O_2731,N_29956,N_29886);
nor UO_2732 (O_2732,N_29988,N_29664);
nor UO_2733 (O_2733,N_29606,N_29440);
nand UO_2734 (O_2734,N_29658,N_29628);
and UO_2735 (O_2735,N_29426,N_29766);
nand UO_2736 (O_2736,N_29883,N_29897);
or UO_2737 (O_2737,N_29956,N_29730);
nor UO_2738 (O_2738,N_29972,N_29788);
or UO_2739 (O_2739,N_29606,N_29634);
nand UO_2740 (O_2740,N_29734,N_29983);
or UO_2741 (O_2741,N_29419,N_29536);
or UO_2742 (O_2742,N_29590,N_29430);
and UO_2743 (O_2743,N_29911,N_29978);
nor UO_2744 (O_2744,N_29418,N_29786);
nand UO_2745 (O_2745,N_29732,N_29404);
or UO_2746 (O_2746,N_29401,N_29902);
or UO_2747 (O_2747,N_29509,N_29687);
nor UO_2748 (O_2748,N_29406,N_29456);
nor UO_2749 (O_2749,N_29521,N_29468);
or UO_2750 (O_2750,N_29824,N_29459);
or UO_2751 (O_2751,N_29887,N_29771);
nor UO_2752 (O_2752,N_29576,N_29902);
nor UO_2753 (O_2753,N_29985,N_29746);
nand UO_2754 (O_2754,N_29650,N_29510);
and UO_2755 (O_2755,N_29915,N_29504);
and UO_2756 (O_2756,N_29438,N_29829);
or UO_2757 (O_2757,N_29974,N_29488);
nand UO_2758 (O_2758,N_29443,N_29943);
or UO_2759 (O_2759,N_29527,N_29433);
nand UO_2760 (O_2760,N_29511,N_29600);
and UO_2761 (O_2761,N_29482,N_29859);
or UO_2762 (O_2762,N_29433,N_29871);
and UO_2763 (O_2763,N_29602,N_29919);
nand UO_2764 (O_2764,N_29495,N_29827);
or UO_2765 (O_2765,N_29481,N_29591);
and UO_2766 (O_2766,N_29821,N_29634);
or UO_2767 (O_2767,N_29424,N_29582);
nand UO_2768 (O_2768,N_29920,N_29661);
or UO_2769 (O_2769,N_29534,N_29648);
nor UO_2770 (O_2770,N_29417,N_29691);
nand UO_2771 (O_2771,N_29727,N_29492);
and UO_2772 (O_2772,N_29793,N_29660);
or UO_2773 (O_2773,N_29745,N_29655);
nand UO_2774 (O_2774,N_29656,N_29687);
nand UO_2775 (O_2775,N_29503,N_29782);
nor UO_2776 (O_2776,N_29606,N_29902);
nor UO_2777 (O_2777,N_29620,N_29640);
nor UO_2778 (O_2778,N_29820,N_29457);
nor UO_2779 (O_2779,N_29665,N_29619);
or UO_2780 (O_2780,N_29483,N_29491);
nor UO_2781 (O_2781,N_29581,N_29763);
or UO_2782 (O_2782,N_29415,N_29711);
nand UO_2783 (O_2783,N_29720,N_29467);
and UO_2784 (O_2784,N_29953,N_29592);
nor UO_2785 (O_2785,N_29491,N_29414);
and UO_2786 (O_2786,N_29493,N_29823);
nand UO_2787 (O_2787,N_29416,N_29492);
or UO_2788 (O_2788,N_29816,N_29653);
or UO_2789 (O_2789,N_29424,N_29756);
nor UO_2790 (O_2790,N_29791,N_29602);
nor UO_2791 (O_2791,N_29944,N_29670);
and UO_2792 (O_2792,N_29892,N_29734);
nand UO_2793 (O_2793,N_29545,N_29864);
or UO_2794 (O_2794,N_29526,N_29612);
or UO_2795 (O_2795,N_29953,N_29843);
and UO_2796 (O_2796,N_29803,N_29560);
nand UO_2797 (O_2797,N_29403,N_29845);
nor UO_2798 (O_2798,N_29834,N_29814);
or UO_2799 (O_2799,N_29932,N_29628);
and UO_2800 (O_2800,N_29836,N_29458);
nand UO_2801 (O_2801,N_29831,N_29412);
or UO_2802 (O_2802,N_29588,N_29993);
nand UO_2803 (O_2803,N_29841,N_29629);
or UO_2804 (O_2804,N_29907,N_29782);
nor UO_2805 (O_2805,N_29687,N_29423);
nor UO_2806 (O_2806,N_29737,N_29666);
or UO_2807 (O_2807,N_29642,N_29509);
nand UO_2808 (O_2808,N_29692,N_29547);
nor UO_2809 (O_2809,N_29916,N_29748);
and UO_2810 (O_2810,N_29993,N_29963);
and UO_2811 (O_2811,N_29868,N_29781);
or UO_2812 (O_2812,N_29515,N_29780);
and UO_2813 (O_2813,N_29524,N_29578);
nand UO_2814 (O_2814,N_29855,N_29461);
nand UO_2815 (O_2815,N_29464,N_29412);
nor UO_2816 (O_2816,N_29450,N_29821);
nor UO_2817 (O_2817,N_29776,N_29995);
nand UO_2818 (O_2818,N_29506,N_29431);
or UO_2819 (O_2819,N_29452,N_29762);
and UO_2820 (O_2820,N_29851,N_29774);
and UO_2821 (O_2821,N_29556,N_29578);
nand UO_2822 (O_2822,N_29676,N_29963);
nand UO_2823 (O_2823,N_29534,N_29811);
or UO_2824 (O_2824,N_29904,N_29901);
nor UO_2825 (O_2825,N_29824,N_29819);
or UO_2826 (O_2826,N_29586,N_29618);
or UO_2827 (O_2827,N_29503,N_29776);
and UO_2828 (O_2828,N_29821,N_29521);
or UO_2829 (O_2829,N_29603,N_29468);
nor UO_2830 (O_2830,N_29727,N_29498);
nor UO_2831 (O_2831,N_29901,N_29806);
and UO_2832 (O_2832,N_29894,N_29943);
nand UO_2833 (O_2833,N_29988,N_29607);
and UO_2834 (O_2834,N_29716,N_29560);
or UO_2835 (O_2835,N_29637,N_29755);
and UO_2836 (O_2836,N_29466,N_29650);
nand UO_2837 (O_2837,N_29400,N_29553);
and UO_2838 (O_2838,N_29572,N_29723);
nor UO_2839 (O_2839,N_29443,N_29863);
nor UO_2840 (O_2840,N_29473,N_29477);
nor UO_2841 (O_2841,N_29962,N_29715);
nor UO_2842 (O_2842,N_29531,N_29665);
nand UO_2843 (O_2843,N_29493,N_29590);
and UO_2844 (O_2844,N_29424,N_29767);
nor UO_2845 (O_2845,N_29834,N_29505);
and UO_2846 (O_2846,N_29975,N_29440);
or UO_2847 (O_2847,N_29983,N_29524);
and UO_2848 (O_2848,N_29470,N_29461);
and UO_2849 (O_2849,N_29741,N_29646);
nand UO_2850 (O_2850,N_29456,N_29449);
or UO_2851 (O_2851,N_29627,N_29481);
or UO_2852 (O_2852,N_29634,N_29936);
or UO_2853 (O_2853,N_29936,N_29960);
nand UO_2854 (O_2854,N_29807,N_29440);
nand UO_2855 (O_2855,N_29660,N_29697);
and UO_2856 (O_2856,N_29640,N_29839);
and UO_2857 (O_2857,N_29884,N_29451);
nand UO_2858 (O_2858,N_29408,N_29796);
and UO_2859 (O_2859,N_29859,N_29485);
nand UO_2860 (O_2860,N_29829,N_29477);
and UO_2861 (O_2861,N_29495,N_29759);
nand UO_2862 (O_2862,N_29757,N_29579);
and UO_2863 (O_2863,N_29770,N_29625);
nand UO_2864 (O_2864,N_29948,N_29717);
nor UO_2865 (O_2865,N_29593,N_29683);
and UO_2866 (O_2866,N_29812,N_29664);
or UO_2867 (O_2867,N_29874,N_29920);
or UO_2868 (O_2868,N_29708,N_29488);
or UO_2869 (O_2869,N_29642,N_29412);
nand UO_2870 (O_2870,N_29718,N_29892);
and UO_2871 (O_2871,N_29601,N_29653);
and UO_2872 (O_2872,N_29971,N_29673);
nor UO_2873 (O_2873,N_29908,N_29413);
nor UO_2874 (O_2874,N_29933,N_29869);
nand UO_2875 (O_2875,N_29981,N_29897);
and UO_2876 (O_2876,N_29899,N_29559);
nand UO_2877 (O_2877,N_29436,N_29907);
nor UO_2878 (O_2878,N_29464,N_29698);
or UO_2879 (O_2879,N_29551,N_29750);
nand UO_2880 (O_2880,N_29700,N_29729);
and UO_2881 (O_2881,N_29986,N_29895);
nor UO_2882 (O_2882,N_29783,N_29590);
nand UO_2883 (O_2883,N_29987,N_29920);
nor UO_2884 (O_2884,N_29930,N_29805);
and UO_2885 (O_2885,N_29605,N_29609);
or UO_2886 (O_2886,N_29547,N_29628);
or UO_2887 (O_2887,N_29867,N_29550);
or UO_2888 (O_2888,N_29408,N_29609);
nor UO_2889 (O_2889,N_29443,N_29413);
xor UO_2890 (O_2890,N_29481,N_29715);
or UO_2891 (O_2891,N_29742,N_29653);
or UO_2892 (O_2892,N_29735,N_29559);
or UO_2893 (O_2893,N_29813,N_29959);
nand UO_2894 (O_2894,N_29763,N_29786);
nand UO_2895 (O_2895,N_29869,N_29514);
or UO_2896 (O_2896,N_29401,N_29856);
and UO_2897 (O_2897,N_29707,N_29932);
nand UO_2898 (O_2898,N_29440,N_29700);
and UO_2899 (O_2899,N_29474,N_29714);
or UO_2900 (O_2900,N_29570,N_29989);
and UO_2901 (O_2901,N_29803,N_29784);
nand UO_2902 (O_2902,N_29734,N_29852);
nor UO_2903 (O_2903,N_29982,N_29886);
or UO_2904 (O_2904,N_29822,N_29756);
xor UO_2905 (O_2905,N_29731,N_29486);
and UO_2906 (O_2906,N_29972,N_29699);
and UO_2907 (O_2907,N_29736,N_29988);
and UO_2908 (O_2908,N_29639,N_29685);
and UO_2909 (O_2909,N_29474,N_29642);
and UO_2910 (O_2910,N_29687,N_29994);
xnor UO_2911 (O_2911,N_29439,N_29739);
and UO_2912 (O_2912,N_29777,N_29718);
nand UO_2913 (O_2913,N_29455,N_29845);
and UO_2914 (O_2914,N_29709,N_29668);
and UO_2915 (O_2915,N_29695,N_29585);
nand UO_2916 (O_2916,N_29779,N_29896);
and UO_2917 (O_2917,N_29640,N_29974);
or UO_2918 (O_2918,N_29625,N_29650);
or UO_2919 (O_2919,N_29941,N_29888);
or UO_2920 (O_2920,N_29657,N_29524);
or UO_2921 (O_2921,N_29759,N_29926);
nor UO_2922 (O_2922,N_29986,N_29766);
nand UO_2923 (O_2923,N_29662,N_29830);
and UO_2924 (O_2924,N_29752,N_29639);
nand UO_2925 (O_2925,N_29648,N_29925);
nand UO_2926 (O_2926,N_29833,N_29680);
nand UO_2927 (O_2927,N_29493,N_29514);
nor UO_2928 (O_2928,N_29714,N_29614);
or UO_2929 (O_2929,N_29876,N_29778);
and UO_2930 (O_2930,N_29780,N_29826);
and UO_2931 (O_2931,N_29622,N_29513);
and UO_2932 (O_2932,N_29850,N_29932);
and UO_2933 (O_2933,N_29868,N_29575);
or UO_2934 (O_2934,N_29849,N_29484);
nor UO_2935 (O_2935,N_29859,N_29978);
nand UO_2936 (O_2936,N_29855,N_29589);
or UO_2937 (O_2937,N_29930,N_29508);
nand UO_2938 (O_2938,N_29918,N_29511);
or UO_2939 (O_2939,N_29638,N_29554);
and UO_2940 (O_2940,N_29504,N_29429);
nand UO_2941 (O_2941,N_29583,N_29752);
or UO_2942 (O_2942,N_29883,N_29863);
or UO_2943 (O_2943,N_29789,N_29544);
nand UO_2944 (O_2944,N_29442,N_29824);
and UO_2945 (O_2945,N_29562,N_29926);
nor UO_2946 (O_2946,N_29637,N_29765);
nand UO_2947 (O_2947,N_29404,N_29449);
or UO_2948 (O_2948,N_29725,N_29939);
and UO_2949 (O_2949,N_29490,N_29960);
and UO_2950 (O_2950,N_29459,N_29592);
nor UO_2951 (O_2951,N_29536,N_29827);
nor UO_2952 (O_2952,N_29722,N_29567);
or UO_2953 (O_2953,N_29832,N_29808);
xor UO_2954 (O_2954,N_29426,N_29611);
xor UO_2955 (O_2955,N_29558,N_29685);
or UO_2956 (O_2956,N_29632,N_29765);
nand UO_2957 (O_2957,N_29938,N_29465);
xor UO_2958 (O_2958,N_29917,N_29915);
and UO_2959 (O_2959,N_29502,N_29492);
nand UO_2960 (O_2960,N_29806,N_29721);
and UO_2961 (O_2961,N_29862,N_29683);
or UO_2962 (O_2962,N_29694,N_29613);
nor UO_2963 (O_2963,N_29478,N_29968);
nor UO_2964 (O_2964,N_29440,N_29706);
or UO_2965 (O_2965,N_29799,N_29917);
or UO_2966 (O_2966,N_29484,N_29963);
nand UO_2967 (O_2967,N_29401,N_29874);
xor UO_2968 (O_2968,N_29987,N_29510);
nor UO_2969 (O_2969,N_29558,N_29710);
nand UO_2970 (O_2970,N_29872,N_29689);
nor UO_2971 (O_2971,N_29816,N_29401);
or UO_2972 (O_2972,N_29664,N_29954);
nand UO_2973 (O_2973,N_29449,N_29886);
and UO_2974 (O_2974,N_29458,N_29822);
and UO_2975 (O_2975,N_29583,N_29566);
nor UO_2976 (O_2976,N_29524,N_29618);
or UO_2977 (O_2977,N_29932,N_29729);
and UO_2978 (O_2978,N_29576,N_29545);
nor UO_2979 (O_2979,N_29468,N_29776);
or UO_2980 (O_2980,N_29663,N_29998);
nand UO_2981 (O_2981,N_29871,N_29515);
nand UO_2982 (O_2982,N_29969,N_29747);
or UO_2983 (O_2983,N_29596,N_29789);
and UO_2984 (O_2984,N_29833,N_29836);
nor UO_2985 (O_2985,N_29827,N_29917);
nand UO_2986 (O_2986,N_29624,N_29831);
nor UO_2987 (O_2987,N_29986,N_29487);
and UO_2988 (O_2988,N_29660,N_29810);
nand UO_2989 (O_2989,N_29436,N_29995);
nand UO_2990 (O_2990,N_29644,N_29407);
or UO_2991 (O_2991,N_29580,N_29730);
nor UO_2992 (O_2992,N_29505,N_29551);
and UO_2993 (O_2993,N_29672,N_29601);
nor UO_2994 (O_2994,N_29799,N_29843);
nor UO_2995 (O_2995,N_29839,N_29912);
nand UO_2996 (O_2996,N_29635,N_29657);
or UO_2997 (O_2997,N_29434,N_29986);
nand UO_2998 (O_2998,N_29992,N_29908);
nor UO_2999 (O_2999,N_29867,N_29672);
and UO_3000 (O_3000,N_29898,N_29666);
nor UO_3001 (O_3001,N_29608,N_29556);
or UO_3002 (O_3002,N_29956,N_29825);
and UO_3003 (O_3003,N_29718,N_29708);
nand UO_3004 (O_3004,N_29907,N_29558);
xor UO_3005 (O_3005,N_29442,N_29455);
and UO_3006 (O_3006,N_29434,N_29879);
nor UO_3007 (O_3007,N_29723,N_29957);
nand UO_3008 (O_3008,N_29472,N_29591);
and UO_3009 (O_3009,N_29493,N_29906);
nand UO_3010 (O_3010,N_29998,N_29681);
nand UO_3011 (O_3011,N_29768,N_29493);
or UO_3012 (O_3012,N_29497,N_29796);
and UO_3013 (O_3013,N_29528,N_29918);
and UO_3014 (O_3014,N_29716,N_29982);
nand UO_3015 (O_3015,N_29682,N_29914);
xor UO_3016 (O_3016,N_29447,N_29420);
or UO_3017 (O_3017,N_29590,N_29922);
and UO_3018 (O_3018,N_29492,N_29836);
or UO_3019 (O_3019,N_29667,N_29665);
and UO_3020 (O_3020,N_29692,N_29582);
or UO_3021 (O_3021,N_29618,N_29994);
nand UO_3022 (O_3022,N_29690,N_29881);
nand UO_3023 (O_3023,N_29850,N_29613);
and UO_3024 (O_3024,N_29772,N_29617);
or UO_3025 (O_3025,N_29627,N_29750);
nand UO_3026 (O_3026,N_29752,N_29481);
and UO_3027 (O_3027,N_29552,N_29631);
or UO_3028 (O_3028,N_29456,N_29850);
nor UO_3029 (O_3029,N_29682,N_29567);
nor UO_3030 (O_3030,N_29585,N_29722);
or UO_3031 (O_3031,N_29755,N_29905);
or UO_3032 (O_3032,N_29990,N_29663);
or UO_3033 (O_3033,N_29941,N_29472);
nand UO_3034 (O_3034,N_29712,N_29955);
or UO_3035 (O_3035,N_29739,N_29608);
nand UO_3036 (O_3036,N_29946,N_29811);
nand UO_3037 (O_3037,N_29728,N_29518);
nor UO_3038 (O_3038,N_29556,N_29704);
or UO_3039 (O_3039,N_29670,N_29838);
or UO_3040 (O_3040,N_29830,N_29698);
nor UO_3041 (O_3041,N_29682,N_29452);
nor UO_3042 (O_3042,N_29825,N_29707);
nor UO_3043 (O_3043,N_29933,N_29699);
or UO_3044 (O_3044,N_29589,N_29830);
nor UO_3045 (O_3045,N_29470,N_29705);
nand UO_3046 (O_3046,N_29412,N_29997);
and UO_3047 (O_3047,N_29919,N_29985);
nand UO_3048 (O_3048,N_29414,N_29990);
nor UO_3049 (O_3049,N_29795,N_29789);
nand UO_3050 (O_3050,N_29580,N_29694);
or UO_3051 (O_3051,N_29764,N_29584);
nor UO_3052 (O_3052,N_29893,N_29950);
and UO_3053 (O_3053,N_29529,N_29727);
nand UO_3054 (O_3054,N_29430,N_29583);
and UO_3055 (O_3055,N_29745,N_29683);
and UO_3056 (O_3056,N_29578,N_29828);
and UO_3057 (O_3057,N_29640,N_29814);
nand UO_3058 (O_3058,N_29558,N_29568);
nand UO_3059 (O_3059,N_29990,N_29987);
nand UO_3060 (O_3060,N_29497,N_29888);
nor UO_3061 (O_3061,N_29597,N_29524);
nand UO_3062 (O_3062,N_29839,N_29573);
nor UO_3063 (O_3063,N_29537,N_29486);
or UO_3064 (O_3064,N_29623,N_29829);
nand UO_3065 (O_3065,N_29901,N_29722);
nor UO_3066 (O_3066,N_29873,N_29679);
nor UO_3067 (O_3067,N_29501,N_29728);
nand UO_3068 (O_3068,N_29842,N_29482);
nand UO_3069 (O_3069,N_29607,N_29513);
nand UO_3070 (O_3070,N_29920,N_29739);
and UO_3071 (O_3071,N_29699,N_29988);
nand UO_3072 (O_3072,N_29699,N_29968);
nand UO_3073 (O_3073,N_29708,N_29548);
nor UO_3074 (O_3074,N_29598,N_29716);
nor UO_3075 (O_3075,N_29443,N_29882);
nand UO_3076 (O_3076,N_29856,N_29742);
or UO_3077 (O_3077,N_29787,N_29758);
nand UO_3078 (O_3078,N_29590,N_29472);
and UO_3079 (O_3079,N_29594,N_29746);
nor UO_3080 (O_3080,N_29928,N_29477);
and UO_3081 (O_3081,N_29655,N_29961);
or UO_3082 (O_3082,N_29467,N_29452);
and UO_3083 (O_3083,N_29746,N_29712);
and UO_3084 (O_3084,N_29771,N_29847);
xor UO_3085 (O_3085,N_29938,N_29609);
nor UO_3086 (O_3086,N_29427,N_29750);
and UO_3087 (O_3087,N_29515,N_29516);
nor UO_3088 (O_3088,N_29470,N_29653);
nor UO_3089 (O_3089,N_29816,N_29616);
and UO_3090 (O_3090,N_29650,N_29590);
nand UO_3091 (O_3091,N_29965,N_29984);
and UO_3092 (O_3092,N_29581,N_29551);
or UO_3093 (O_3093,N_29467,N_29446);
and UO_3094 (O_3094,N_29921,N_29814);
nand UO_3095 (O_3095,N_29713,N_29929);
nand UO_3096 (O_3096,N_29659,N_29995);
nor UO_3097 (O_3097,N_29915,N_29820);
xor UO_3098 (O_3098,N_29950,N_29757);
nor UO_3099 (O_3099,N_29686,N_29625);
and UO_3100 (O_3100,N_29770,N_29996);
nand UO_3101 (O_3101,N_29439,N_29866);
nor UO_3102 (O_3102,N_29535,N_29528);
or UO_3103 (O_3103,N_29964,N_29819);
or UO_3104 (O_3104,N_29631,N_29423);
or UO_3105 (O_3105,N_29572,N_29699);
or UO_3106 (O_3106,N_29696,N_29536);
nand UO_3107 (O_3107,N_29729,N_29978);
and UO_3108 (O_3108,N_29902,N_29962);
nor UO_3109 (O_3109,N_29762,N_29994);
and UO_3110 (O_3110,N_29698,N_29535);
xnor UO_3111 (O_3111,N_29645,N_29535);
or UO_3112 (O_3112,N_29863,N_29678);
xnor UO_3113 (O_3113,N_29775,N_29463);
nand UO_3114 (O_3114,N_29713,N_29740);
or UO_3115 (O_3115,N_29736,N_29761);
nand UO_3116 (O_3116,N_29542,N_29826);
nand UO_3117 (O_3117,N_29673,N_29618);
or UO_3118 (O_3118,N_29857,N_29838);
nand UO_3119 (O_3119,N_29695,N_29755);
or UO_3120 (O_3120,N_29753,N_29457);
nand UO_3121 (O_3121,N_29744,N_29928);
nand UO_3122 (O_3122,N_29421,N_29661);
or UO_3123 (O_3123,N_29583,N_29687);
or UO_3124 (O_3124,N_29689,N_29724);
or UO_3125 (O_3125,N_29526,N_29969);
and UO_3126 (O_3126,N_29401,N_29478);
or UO_3127 (O_3127,N_29898,N_29762);
nand UO_3128 (O_3128,N_29405,N_29700);
or UO_3129 (O_3129,N_29567,N_29698);
and UO_3130 (O_3130,N_29494,N_29905);
xor UO_3131 (O_3131,N_29864,N_29818);
and UO_3132 (O_3132,N_29766,N_29728);
nor UO_3133 (O_3133,N_29584,N_29816);
xor UO_3134 (O_3134,N_29503,N_29588);
nand UO_3135 (O_3135,N_29581,N_29643);
nor UO_3136 (O_3136,N_29456,N_29685);
nand UO_3137 (O_3137,N_29585,N_29727);
and UO_3138 (O_3138,N_29861,N_29679);
nor UO_3139 (O_3139,N_29759,N_29556);
or UO_3140 (O_3140,N_29776,N_29422);
and UO_3141 (O_3141,N_29987,N_29560);
nand UO_3142 (O_3142,N_29862,N_29621);
nor UO_3143 (O_3143,N_29620,N_29900);
nor UO_3144 (O_3144,N_29679,N_29918);
or UO_3145 (O_3145,N_29951,N_29792);
nand UO_3146 (O_3146,N_29576,N_29570);
and UO_3147 (O_3147,N_29781,N_29557);
nand UO_3148 (O_3148,N_29615,N_29662);
or UO_3149 (O_3149,N_29468,N_29447);
or UO_3150 (O_3150,N_29596,N_29493);
xnor UO_3151 (O_3151,N_29607,N_29507);
xor UO_3152 (O_3152,N_29813,N_29957);
and UO_3153 (O_3153,N_29635,N_29785);
or UO_3154 (O_3154,N_29837,N_29634);
nand UO_3155 (O_3155,N_29423,N_29883);
or UO_3156 (O_3156,N_29662,N_29828);
and UO_3157 (O_3157,N_29622,N_29562);
nor UO_3158 (O_3158,N_29461,N_29643);
and UO_3159 (O_3159,N_29463,N_29921);
or UO_3160 (O_3160,N_29935,N_29930);
and UO_3161 (O_3161,N_29432,N_29979);
and UO_3162 (O_3162,N_29913,N_29990);
nor UO_3163 (O_3163,N_29599,N_29534);
nor UO_3164 (O_3164,N_29443,N_29437);
and UO_3165 (O_3165,N_29772,N_29752);
and UO_3166 (O_3166,N_29649,N_29606);
nand UO_3167 (O_3167,N_29480,N_29547);
nor UO_3168 (O_3168,N_29943,N_29795);
xor UO_3169 (O_3169,N_29581,N_29852);
nand UO_3170 (O_3170,N_29688,N_29814);
xor UO_3171 (O_3171,N_29944,N_29816);
or UO_3172 (O_3172,N_29733,N_29796);
and UO_3173 (O_3173,N_29838,N_29997);
nand UO_3174 (O_3174,N_29556,N_29528);
and UO_3175 (O_3175,N_29540,N_29553);
xor UO_3176 (O_3176,N_29438,N_29944);
or UO_3177 (O_3177,N_29777,N_29820);
nand UO_3178 (O_3178,N_29649,N_29951);
nand UO_3179 (O_3179,N_29736,N_29967);
xor UO_3180 (O_3180,N_29625,N_29559);
and UO_3181 (O_3181,N_29510,N_29794);
nand UO_3182 (O_3182,N_29547,N_29640);
and UO_3183 (O_3183,N_29556,N_29938);
nand UO_3184 (O_3184,N_29834,N_29696);
nand UO_3185 (O_3185,N_29910,N_29986);
or UO_3186 (O_3186,N_29533,N_29527);
or UO_3187 (O_3187,N_29669,N_29438);
xnor UO_3188 (O_3188,N_29827,N_29935);
or UO_3189 (O_3189,N_29740,N_29628);
or UO_3190 (O_3190,N_29535,N_29796);
and UO_3191 (O_3191,N_29901,N_29683);
nand UO_3192 (O_3192,N_29864,N_29779);
and UO_3193 (O_3193,N_29732,N_29525);
and UO_3194 (O_3194,N_29933,N_29464);
or UO_3195 (O_3195,N_29525,N_29815);
nand UO_3196 (O_3196,N_29604,N_29810);
and UO_3197 (O_3197,N_29919,N_29955);
nand UO_3198 (O_3198,N_29402,N_29414);
and UO_3199 (O_3199,N_29909,N_29935);
nand UO_3200 (O_3200,N_29799,N_29510);
and UO_3201 (O_3201,N_29672,N_29795);
nand UO_3202 (O_3202,N_29916,N_29636);
and UO_3203 (O_3203,N_29916,N_29843);
or UO_3204 (O_3204,N_29968,N_29963);
or UO_3205 (O_3205,N_29797,N_29445);
and UO_3206 (O_3206,N_29931,N_29967);
nand UO_3207 (O_3207,N_29983,N_29451);
nor UO_3208 (O_3208,N_29542,N_29779);
and UO_3209 (O_3209,N_29747,N_29614);
and UO_3210 (O_3210,N_29683,N_29492);
or UO_3211 (O_3211,N_29873,N_29697);
and UO_3212 (O_3212,N_29560,N_29671);
and UO_3213 (O_3213,N_29434,N_29600);
and UO_3214 (O_3214,N_29988,N_29433);
nor UO_3215 (O_3215,N_29974,N_29620);
or UO_3216 (O_3216,N_29499,N_29527);
or UO_3217 (O_3217,N_29903,N_29558);
or UO_3218 (O_3218,N_29630,N_29890);
and UO_3219 (O_3219,N_29517,N_29503);
nor UO_3220 (O_3220,N_29826,N_29714);
or UO_3221 (O_3221,N_29828,N_29529);
or UO_3222 (O_3222,N_29591,N_29400);
nor UO_3223 (O_3223,N_29889,N_29893);
nor UO_3224 (O_3224,N_29506,N_29656);
nand UO_3225 (O_3225,N_29492,N_29451);
or UO_3226 (O_3226,N_29970,N_29920);
or UO_3227 (O_3227,N_29449,N_29411);
nor UO_3228 (O_3228,N_29855,N_29807);
and UO_3229 (O_3229,N_29485,N_29498);
or UO_3230 (O_3230,N_29449,N_29628);
and UO_3231 (O_3231,N_29628,N_29575);
and UO_3232 (O_3232,N_29920,N_29978);
and UO_3233 (O_3233,N_29990,N_29492);
or UO_3234 (O_3234,N_29961,N_29603);
and UO_3235 (O_3235,N_29433,N_29728);
nor UO_3236 (O_3236,N_29630,N_29809);
or UO_3237 (O_3237,N_29738,N_29560);
and UO_3238 (O_3238,N_29413,N_29569);
and UO_3239 (O_3239,N_29628,N_29869);
nor UO_3240 (O_3240,N_29850,N_29859);
or UO_3241 (O_3241,N_29826,N_29794);
and UO_3242 (O_3242,N_29708,N_29913);
and UO_3243 (O_3243,N_29450,N_29532);
nor UO_3244 (O_3244,N_29618,N_29447);
nor UO_3245 (O_3245,N_29580,N_29964);
and UO_3246 (O_3246,N_29621,N_29615);
nand UO_3247 (O_3247,N_29744,N_29487);
or UO_3248 (O_3248,N_29891,N_29701);
and UO_3249 (O_3249,N_29992,N_29934);
and UO_3250 (O_3250,N_29619,N_29845);
nand UO_3251 (O_3251,N_29610,N_29949);
nor UO_3252 (O_3252,N_29916,N_29548);
or UO_3253 (O_3253,N_29556,N_29621);
and UO_3254 (O_3254,N_29654,N_29793);
xnor UO_3255 (O_3255,N_29713,N_29981);
and UO_3256 (O_3256,N_29744,N_29842);
nor UO_3257 (O_3257,N_29469,N_29442);
nor UO_3258 (O_3258,N_29951,N_29835);
nand UO_3259 (O_3259,N_29625,N_29508);
nor UO_3260 (O_3260,N_29954,N_29559);
nand UO_3261 (O_3261,N_29931,N_29666);
or UO_3262 (O_3262,N_29772,N_29969);
or UO_3263 (O_3263,N_29582,N_29757);
nor UO_3264 (O_3264,N_29732,N_29582);
or UO_3265 (O_3265,N_29842,N_29539);
and UO_3266 (O_3266,N_29847,N_29884);
nand UO_3267 (O_3267,N_29718,N_29484);
nand UO_3268 (O_3268,N_29523,N_29507);
nand UO_3269 (O_3269,N_29970,N_29618);
nor UO_3270 (O_3270,N_29922,N_29400);
or UO_3271 (O_3271,N_29990,N_29440);
or UO_3272 (O_3272,N_29435,N_29526);
and UO_3273 (O_3273,N_29633,N_29580);
and UO_3274 (O_3274,N_29804,N_29848);
or UO_3275 (O_3275,N_29779,N_29874);
and UO_3276 (O_3276,N_29460,N_29761);
nand UO_3277 (O_3277,N_29766,N_29936);
and UO_3278 (O_3278,N_29902,N_29869);
and UO_3279 (O_3279,N_29866,N_29441);
nand UO_3280 (O_3280,N_29708,N_29868);
nor UO_3281 (O_3281,N_29427,N_29837);
or UO_3282 (O_3282,N_29500,N_29419);
or UO_3283 (O_3283,N_29772,N_29798);
or UO_3284 (O_3284,N_29755,N_29624);
nor UO_3285 (O_3285,N_29446,N_29964);
nor UO_3286 (O_3286,N_29553,N_29747);
nand UO_3287 (O_3287,N_29830,N_29964);
nand UO_3288 (O_3288,N_29427,N_29421);
nand UO_3289 (O_3289,N_29536,N_29722);
and UO_3290 (O_3290,N_29988,N_29454);
nand UO_3291 (O_3291,N_29511,N_29842);
and UO_3292 (O_3292,N_29782,N_29914);
nor UO_3293 (O_3293,N_29865,N_29537);
nor UO_3294 (O_3294,N_29841,N_29451);
nand UO_3295 (O_3295,N_29445,N_29586);
or UO_3296 (O_3296,N_29727,N_29452);
nand UO_3297 (O_3297,N_29527,N_29474);
and UO_3298 (O_3298,N_29942,N_29542);
and UO_3299 (O_3299,N_29899,N_29988);
and UO_3300 (O_3300,N_29957,N_29642);
or UO_3301 (O_3301,N_29595,N_29441);
and UO_3302 (O_3302,N_29797,N_29872);
nor UO_3303 (O_3303,N_29974,N_29480);
nor UO_3304 (O_3304,N_29552,N_29998);
or UO_3305 (O_3305,N_29780,N_29885);
and UO_3306 (O_3306,N_29997,N_29895);
or UO_3307 (O_3307,N_29910,N_29761);
and UO_3308 (O_3308,N_29454,N_29511);
and UO_3309 (O_3309,N_29674,N_29532);
and UO_3310 (O_3310,N_29451,N_29838);
or UO_3311 (O_3311,N_29739,N_29960);
nor UO_3312 (O_3312,N_29934,N_29799);
or UO_3313 (O_3313,N_29778,N_29826);
and UO_3314 (O_3314,N_29666,N_29625);
nor UO_3315 (O_3315,N_29552,N_29549);
nor UO_3316 (O_3316,N_29587,N_29844);
and UO_3317 (O_3317,N_29659,N_29643);
or UO_3318 (O_3318,N_29657,N_29828);
nor UO_3319 (O_3319,N_29842,N_29898);
or UO_3320 (O_3320,N_29959,N_29992);
or UO_3321 (O_3321,N_29720,N_29848);
or UO_3322 (O_3322,N_29546,N_29432);
nand UO_3323 (O_3323,N_29635,N_29529);
nand UO_3324 (O_3324,N_29976,N_29845);
nor UO_3325 (O_3325,N_29804,N_29651);
nor UO_3326 (O_3326,N_29766,N_29744);
nor UO_3327 (O_3327,N_29982,N_29443);
nand UO_3328 (O_3328,N_29445,N_29575);
and UO_3329 (O_3329,N_29664,N_29687);
or UO_3330 (O_3330,N_29460,N_29495);
or UO_3331 (O_3331,N_29915,N_29643);
nor UO_3332 (O_3332,N_29609,N_29966);
nand UO_3333 (O_3333,N_29498,N_29487);
nand UO_3334 (O_3334,N_29618,N_29575);
and UO_3335 (O_3335,N_29445,N_29912);
and UO_3336 (O_3336,N_29975,N_29631);
nand UO_3337 (O_3337,N_29772,N_29556);
nor UO_3338 (O_3338,N_29433,N_29647);
and UO_3339 (O_3339,N_29570,N_29861);
nor UO_3340 (O_3340,N_29954,N_29864);
nand UO_3341 (O_3341,N_29850,N_29597);
nand UO_3342 (O_3342,N_29627,N_29746);
nor UO_3343 (O_3343,N_29464,N_29865);
nor UO_3344 (O_3344,N_29807,N_29962);
nand UO_3345 (O_3345,N_29698,N_29964);
and UO_3346 (O_3346,N_29728,N_29695);
and UO_3347 (O_3347,N_29517,N_29507);
nor UO_3348 (O_3348,N_29945,N_29631);
and UO_3349 (O_3349,N_29548,N_29966);
or UO_3350 (O_3350,N_29538,N_29923);
xnor UO_3351 (O_3351,N_29400,N_29594);
or UO_3352 (O_3352,N_29958,N_29711);
nand UO_3353 (O_3353,N_29635,N_29974);
and UO_3354 (O_3354,N_29692,N_29414);
and UO_3355 (O_3355,N_29805,N_29733);
or UO_3356 (O_3356,N_29812,N_29867);
and UO_3357 (O_3357,N_29807,N_29492);
nor UO_3358 (O_3358,N_29746,N_29699);
or UO_3359 (O_3359,N_29735,N_29613);
nor UO_3360 (O_3360,N_29480,N_29541);
nor UO_3361 (O_3361,N_29537,N_29658);
nor UO_3362 (O_3362,N_29924,N_29683);
nand UO_3363 (O_3363,N_29650,N_29691);
and UO_3364 (O_3364,N_29820,N_29657);
or UO_3365 (O_3365,N_29747,N_29575);
nor UO_3366 (O_3366,N_29488,N_29546);
nand UO_3367 (O_3367,N_29741,N_29727);
nand UO_3368 (O_3368,N_29830,N_29750);
and UO_3369 (O_3369,N_29728,N_29923);
nor UO_3370 (O_3370,N_29608,N_29868);
xor UO_3371 (O_3371,N_29469,N_29925);
xnor UO_3372 (O_3372,N_29560,N_29917);
nor UO_3373 (O_3373,N_29439,N_29897);
or UO_3374 (O_3374,N_29966,N_29654);
and UO_3375 (O_3375,N_29731,N_29756);
or UO_3376 (O_3376,N_29842,N_29549);
and UO_3377 (O_3377,N_29861,N_29703);
nand UO_3378 (O_3378,N_29557,N_29549);
or UO_3379 (O_3379,N_29452,N_29599);
or UO_3380 (O_3380,N_29837,N_29895);
nor UO_3381 (O_3381,N_29827,N_29688);
and UO_3382 (O_3382,N_29578,N_29449);
nor UO_3383 (O_3383,N_29943,N_29932);
nand UO_3384 (O_3384,N_29402,N_29694);
or UO_3385 (O_3385,N_29897,N_29511);
or UO_3386 (O_3386,N_29550,N_29830);
and UO_3387 (O_3387,N_29984,N_29465);
nor UO_3388 (O_3388,N_29641,N_29607);
nor UO_3389 (O_3389,N_29752,N_29890);
nand UO_3390 (O_3390,N_29782,N_29447);
nor UO_3391 (O_3391,N_29477,N_29797);
and UO_3392 (O_3392,N_29888,N_29629);
and UO_3393 (O_3393,N_29577,N_29759);
or UO_3394 (O_3394,N_29685,N_29448);
and UO_3395 (O_3395,N_29835,N_29571);
or UO_3396 (O_3396,N_29768,N_29947);
nand UO_3397 (O_3397,N_29635,N_29885);
nor UO_3398 (O_3398,N_29897,N_29738);
nor UO_3399 (O_3399,N_29408,N_29861);
or UO_3400 (O_3400,N_29872,N_29836);
nand UO_3401 (O_3401,N_29652,N_29905);
nor UO_3402 (O_3402,N_29764,N_29706);
nand UO_3403 (O_3403,N_29524,N_29655);
and UO_3404 (O_3404,N_29548,N_29681);
and UO_3405 (O_3405,N_29496,N_29826);
and UO_3406 (O_3406,N_29667,N_29931);
nor UO_3407 (O_3407,N_29866,N_29973);
nor UO_3408 (O_3408,N_29406,N_29826);
or UO_3409 (O_3409,N_29956,N_29757);
nor UO_3410 (O_3410,N_29617,N_29630);
and UO_3411 (O_3411,N_29852,N_29491);
nand UO_3412 (O_3412,N_29527,N_29964);
nand UO_3413 (O_3413,N_29657,N_29781);
and UO_3414 (O_3414,N_29637,N_29762);
nand UO_3415 (O_3415,N_29682,N_29958);
nor UO_3416 (O_3416,N_29654,N_29829);
and UO_3417 (O_3417,N_29805,N_29477);
nor UO_3418 (O_3418,N_29778,N_29764);
or UO_3419 (O_3419,N_29604,N_29968);
and UO_3420 (O_3420,N_29885,N_29542);
and UO_3421 (O_3421,N_29450,N_29407);
and UO_3422 (O_3422,N_29838,N_29871);
nand UO_3423 (O_3423,N_29944,N_29712);
or UO_3424 (O_3424,N_29646,N_29914);
or UO_3425 (O_3425,N_29508,N_29683);
xor UO_3426 (O_3426,N_29524,N_29691);
or UO_3427 (O_3427,N_29778,N_29467);
nand UO_3428 (O_3428,N_29600,N_29750);
nand UO_3429 (O_3429,N_29635,N_29581);
nand UO_3430 (O_3430,N_29525,N_29677);
or UO_3431 (O_3431,N_29697,N_29762);
nand UO_3432 (O_3432,N_29983,N_29454);
and UO_3433 (O_3433,N_29530,N_29641);
and UO_3434 (O_3434,N_29878,N_29772);
nand UO_3435 (O_3435,N_29424,N_29966);
nand UO_3436 (O_3436,N_29625,N_29670);
and UO_3437 (O_3437,N_29880,N_29555);
nand UO_3438 (O_3438,N_29700,N_29778);
nor UO_3439 (O_3439,N_29585,N_29469);
and UO_3440 (O_3440,N_29746,N_29805);
nor UO_3441 (O_3441,N_29465,N_29503);
nand UO_3442 (O_3442,N_29528,N_29448);
or UO_3443 (O_3443,N_29475,N_29563);
nor UO_3444 (O_3444,N_29864,N_29453);
and UO_3445 (O_3445,N_29893,N_29470);
or UO_3446 (O_3446,N_29461,N_29960);
nor UO_3447 (O_3447,N_29504,N_29701);
nand UO_3448 (O_3448,N_29490,N_29471);
nor UO_3449 (O_3449,N_29733,N_29550);
nor UO_3450 (O_3450,N_29880,N_29989);
or UO_3451 (O_3451,N_29978,N_29759);
nand UO_3452 (O_3452,N_29933,N_29490);
nor UO_3453 (O_3453,N_29877,N_29448);
nand UO_3454 (O_3454,N_29734,N_29655);
or UO_3455 (O_3455,N_29765,N_29859);
nor UO_3456 (O_3456,N_29845,N_29568);
and UO_3457 (O_3457,N_29854,N_29958);
nor UO_3458 (O_3458,N_29427,N_29464);
nand UO_3459 (O_3459,N_29462,N_29795);
and UO_3460 (O_3460,N_29799,N_29716);
and UO_3461 (O_3461,N_29468,N_29812);
or UO_3462 (O_3462,N_29469,N_29666);
or UO_3463 (O_3463,N_29835,N_29943);
nor UO_3464 (O_3464,N_29600,N_29757);
and UO_3465 (O_3465,N_29867,N_29584);
or UO_3466 (O_3466,N_29531,N_29794);
and UO_3467 (O_3467,N_29492,N_29641);
nor UO_3468 (O_3468,N_29689,N_29430);
nand UO_3469 (O_3469,N_29660,N_29690);
and UO_3470 (O_3470,N_29945,N_29916);
and UO_3471 (O_3471,N_29711,N_29887);
nand UO_3472 (O_3472,N_29599,N_29660);
or UO_3473 (O_3473,N_29753,N_29847);
nand UO_3474 (O_3474,N_29775,N_29548);
or UO_3475 (O_3475,N_29605,N_29614);
or UO_3476 (O_3476,N_29450,N_29681);
or UO_3477 (O_3477,N_29610,N_29622);
and UO_3478 (O_3478,N_29537,N_29673);
xor UO_3479 (O_3479,N_29591,N_29784);
and UO_3480 (O_3480,N_29747,N_29560);
and UO_3481 (O_3481,N_29809,N_29641);
or UO_3482 (O_3482,N_29737,N_29504);
nor UO_3483 (O_3483,N_29634,N_29679);
nor UO_3484 (O_3484,N_29468,N_29597);
nand UO_3485 (O_3485,N_29432,N_29453);
and UO_3486 (O_3486,N_29605,N_29512);
or UO_3487 (O_3487,N_29753,N_29745);
and UO_3488 (O_3488,N_29753,N_29477);
and UO_3489 (O_3489,N_29846,N_29977);
and UO_3490 (O_3490,N_29408,N_29774);
and UO_3491 (O_3491,N_29825,N_29407);
nor UO_3492 (O_3492,N_29962,N_29498);
nor UO_3493 (O_3493,N_29448,N_29660);
or UO_3494 (O_3494,N_29686,N_29882);
or UO_3495 (O_3495,N_29683,N_29571);
nor UO_3496 (O_3496,N_29439,N_29702);
nand UO_3497 (O_3497,N_29754,N_29760);
nor UO_3498 (O_3498,N_29865,N_29458);
nor UO_3499 (O_3499,N_29410,N_29470);
endmodule