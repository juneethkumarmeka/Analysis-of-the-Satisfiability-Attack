module basic_750_5000_1000_5_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_258,In_365);
nor U1 (N_1,In_264,In_160);
and U2 (N_2,In_461,In_534);
or U3 (N_3,In_293,In_496);
or U4 (N_4,In_104,In_46);
and U5 (N_5,In_121,In_243);
and U6 (N_6,In_512,In_54);
and U7 (N_7,In_370,In_149);
xor U8 (N_8,In_682,In_84);
nand U9 (N_9,In_234,In_256);
nand U10 (N_10,In_635,In_519);
or U11 (N_11,In_51,In_316);
or U12 (N_12,In_313,In_333);
and U13 (N_13,In_450,In_436);
or U14 (N_14,In_688,In_631);
nor U15 (N_15,In_69,In_398);
and U16 (N_16,In_570,In_699);
nand U17 (N_17,In_711,In_408);
or U18 (N_18,In_576,In_574);
nor U19 (N_19,In_20,In_210);
or U20 (N_20,In_40,In_696);
nand U21 (N_21,In_678,In_384);
and U22 (N_22,In_233,In_77);
nand U23 (N_23,In_579,In_113);
and U24 (N_24,In_493,In_75);
or U25 (N_25,In_589,In_251);
nand U26 (N_26,In_561,In_383);
nor U27 (N_27,In_319,In_608);
xor U28 (N_28,In_118,In_217);
and U29 (N_29,In_394,In_713);
or U30 (N_30,In_128,In_137);
xor U31 (N_31,In_470,In_301);
or U32 (N_32,In_86,In_404);
nor U33 (N_33,In_577,In_261);
nand U34 (N_34,In_98,In_689);
and U35 (N_35,In_308,In_562);
and U36 (N_36,In_24,In_541);
or U37 (N_37,In_721,In_226);
nor U38 (N_38,In_397,In_103);
nand U39 (N_39,In_247,In_277);
and U40 (N_40,In_71,In_532);
and U41 (N_41,In_648,In_215);
nand U42 (N_42,In_654,In_416);
nor U43 (N_43,In_553,In_652);
or U44 (N_44,In_677,In_203);
nor U45 (N_45,In_419,In_194);
nand U46 (N_46,In_503,In_68);
nand U47 (N_47,In_428,In_510);
nand U48 (N_48,In_411,In_235);
or U49 (N_49,In_422,In_427);
nor U50 (N_50,In_460,In_19);
or U51 (N_51,In_260,In_584);
nor U52 (N_52,In_191,In_708);
nor U53 (N_53,In_209,In_352);
nor U54 (N_54,In_35,In_535);
nand U55 (N_55,In_403,In_701);
nand U56 (N_56,In_401,In_431);
or U57 (N_57,In_318,In_244);
nor U58 (N_58,In_178,In_249);
xnor U59 (N_59,In_747,In_520);
nand U60 (N_60,In_691,In_311);
and U61 (N_61,In_458,In_294);
or U62 (N_62,In_9,In_624);
or U63 (N_63,In_373,In_325);
or U64 (N_64,In_399,In_729);
nor U65 (N_65,In_697,In_495);
nor U66 (N_66,In_491,In_192);
nor U67 (N_67,In_615,In_22);
nor U68 (N_68,In_374,In_471);
and U69 (N_69,In_257,In_58);
or U70 (N_70,In_281,In_7);
nor U71 (N_71,In_400,In_671);
and U72 (N_72,In_332,In_492);
xnor U73 (N_73,In_15,In_546);
or U74 (N_74,In_368,In_594);
nor U75 (N_75,In_48,In_307);
or U76 (N_76,In_57,In_129);
nor U77 (N_77,In_228,In_551);
nor U78 (N_78,In_600,In_369);
nor U79 (N_79,In_120,In_457);
nand U80 (N_80,In_274,In_164);
and U81 (N_81,In_517,In_93);
and U82 (N_82,In_662,In_564);
nand U83 (N_83,In_59,In_356);
or U84 (N_84,In_557,In_273);
nand U85 (N_85,In_593,In_702);
or U86 (N_86,In_549,In_425);
xor U87 (N_87,In_296,In_645);
xor U88 (N_88,In_444,In_315);
and U89 (N_89,In_92,In_720);
nor U90 (N_90,In_693,In_611);
and U91 (N_91,In_82,In_483);
or U92 (N_92,In_28,In_441);
nand U93 (N_93,In_38,In_353);
and U94 (N_94,In_230,In_245);
or U95 (N_95,In_237,In_133);
nor U96 (N_96,In_464,In_272);
nor U97 (N_97,In_622,In_321);
nand U98 (N_98,In_110,In_350);
nor U99 (N_99,In_379,In_467);
nor U100 (N_100,In_67,In_544);
and U101 (N_101,In_547,In_629);
and U102 (N_102,In_604,In_34);
nor U103 (N_103,In_423,In_288);
and U104 (N_104,In_651,In_170);
and U105 (N_105,In_539,In_533);
nor U106 (N_106,In_222,In_214);
nand U107 (N_107,In_679,In_744);
and U108 (N_108,In_16,In_672);
and U109 (N_109,In_43,In_636);
nand U110 (N_110,In_601,In_649);
nor U111 (N_111,In_198,In_717);
nand U112 (N_112,In_418,In_537);
and U113 (N_113,In_465,In_502);
and U114 (N_114,In_466,In_481);
nor U115 (N_115,In_530,In_36);
nor U116 (N_116,In_227,In_734);
and U117 (N_117,In_163,In_56);
nor U118 (N_118,In_710,In_115);
and U119 (N_119,In_151,In_168);
nand U120 (N_120,In_50,In_681);
nor U121 (N_121,In_5,In_507);
nand U122 (N_122,In_367,In_33);
or U123 (N_123,In_206,In_501);
nand U124 (N_124,In_80,In_433);
or U125 (N_125,In_437,In_569);
nor U126 (N_126,In_730,In_27);
nand U127 (N_127,In_52,In_141);
nand U128 (N_128,In_154,In_632);
nor U129 (N_129,In_606,In_447);
nor U130 (N_130,In_346,In_182);
nor U131 (N_131,In_148,In_452);
or U132 (N_132,In_665,In_638);
nand U133 (N_133,In_336,In_363);
or U134 (N_134,In_341,In_78);
nand U135 (N_135,In_402,In_79);
nand U136 (N_136,In_468,In_190);
or U137 (N_137,In_498,In_11);
nor U138 (N_138,In_617,In_565);
or U139 (N_139,In_676,In_47);
and U140 (N_140,In_463,In_89);
or U141 (N_141,In_337,In_236);
or U142 (N_142,In_375,In_131);
and U143 (N_143,In_386,In_359);
and U144 (N_144,In_60,In_279);
nor U145 (N_145,In_738,In_349);
nand U146 (N_146,In_12,In_516);
or U147 (N_147,In_372,In_511);
nor U148 (N_148,In_737,In_630);
nand U149 (N_149,In_625,In_587);
nor U150 (N_150,In_73,In_176);
and U151 (N_151,In_263,In_66);
or U152 (N_152,In_240,In_265);
and U153 (N_153,In_613,In_207);
nor U154 (N_154,In_515,In_508);
and U155 (N_155,In_591,In_159);
nor U156 (N_156,In_116,In_647);
nor U157 (N_157,In_18,In_83);
and U158 (N_158,In_195,In_312);
and U159 (N_159,In_527,In_255);
nor U160 (N_160,In_199,In_304);
and U161 (N_161,In_142,In_582);
and U162 (N_162,In_477,In_575);
nand U163 (N_163,In_396,In_513);
and U164 (N_164,In_497,In_571);
nand U165 (N_165,In_581,In_3);
nor U166 (N_166,In_266,In_438);
nor U167 (N_167,In_588,In_742);
and U168 (N_168,In_595,In_123);
nand U169 (N_169,In_674,In_642);
nor U170 (N_170,In_414,In_271);
nor U171 (N_171,In_443,In_719);
nand U172 (N_172,In_31,In_543);
nand U173 (N_173,In_153,In_224);
nor U174 (N_174,In_446,In_268);
or U175 (N_175,In_152,In_572);
and U176 (N_176,In_101,In_165);
or U177 (N_177,In_320,In_690);
nor U178 (N_178,In_76,In_392);
or U179 (N_179,In_698,In_108);
or U180 (N_180,In_482,In_391);
xnor U181 (N_181,In_220,In_716);
or U182 (N_182,In_405,In_692);
nand U183 (N_183,In_25,In_590);
nand U184 (N_184,In_567,In_727);
nand U185 (N_185,In_655,In_669);
or U186 (N_186,In_749,In_90);
nor U187 (N_187,In_454,In_340);
or U188 (N_188,In_695,In_70);
and U189 (N_189,In_139,In_620);
and U190 (N_190,In_687,In_322);
nand U191 (N_191,In_552,In_596);
nor U192 (N_192,In_259,In_189);
or U193 (N_193,In_521,In_23);
nand U194 (N_194,In_732,In_150);
nor U195 (N_195,In_653,In_156);
or U196 (N_196,In_739,In_700);
or U197 (N_197,In_107,In_122);
and U198 (N_198,In_167,In_105);
and U199 (N_199,In_718,In_683);
or U200 (N_200,In_395,In_639);
and U201 (N_201,In_646,In_410);
and U202 (N_202,In_500,In_586);
or U203 (N_203,In_81,In_169);
or U204 (N_204,In_354,In_360);
nand U205 (N_205,In_218,In_585);
or U206 (N_206,In_278,In_284);
nor U207 (N_207,In_602,In_30);
and U208 (N_208,In_314,In_455);
or U209 (N_209,In_451,In_573);
nand U210 (N_210,In_117,In_280);
nor U211 (N_211,In_309,In_724);
nor U212 (N_212,In_1,In_469);
or U213 (N_213,In_420,In_327);
or U214 (N_214,In_37,In_177);
nor U215 (N_215,In_74,In_221);
nand U216 (N_216,In_72,In_343);
nor U217 (N_217,In_14,In_184);
or U218 (N_218,In_705,In_283);
and U219 (N_219,In_173,In_556);
or U220 (N_220,In_714,In_554);
nand U221 (N_221,In_299,In_248);
nor U222 (N_222,In_559,In_435);
xor U223 (N_223,In_49,In_479);
and U224 (N_224,In_204,In_621);
nand U225 (N_225,In_489,In_715);
xnor U226 (N_226,In_41,In_342);
and U227 (N_227,In_310,In_641);
nor U228 (N_228,In_685,In_439);
nand U229 (N_229,In_740,In_487);
and U230 (N_230,In_253,In_509);
and U231 (N_231,In_526,In_112);
and U232 (N_232,In_607,In_331);
and U233 (N_233,In_506,In_667);
nor U234 (N_234,In_389,In_550);
and U235 (N_235,In_643,In_453);
xor U236 (N_236,In_324,In_114);
nand U237 (N_237,In_95,In_96);
nand U238 (N_238,In_171,In_225);
xor U239 (N_239,In_135,In_388);
nor U240 (N_240,In_476,In_475);
or U241 (N_241,In_426,In_640);
nor U242 (N_242,In_741,In_205);
or U243 (N_243,In_140,In_65);
nand U244 (N_244,In_614,In_229);
and U245 (N_245,In_499,In_295);
nor U246 (N_246,In_147,In_548);
and U247 (N_247,In_578,In_109);
or U248 (N_248,In_175,In_523);
or U249 (N_249,In_155,In_219);
nand U250 (N_250,In_282,In_100);
and U251 (N_251,In_241,In_650);
and U252 (N_252,In_657,In_166);
nor U253 (N_253,In_538,In_459);
and U254 (N_254,In_663,In_659);
or U255 (N_255,In_335,In_361);
and U256 (N_256,In_364,In_64);
and U257 (N_257,In_239,In_597);
or U258 (N_258,In_449,In_474);
xnor U259 (N_259,In_382,In_242);
or U260 (N_260,In_473,In_130);
or U261 (N_261,In_136,In_8);
nor U262 (N_262,In_186,In_406);
nand U263 (N_263,In_627,In_270);
xor U264 (N_264,In_85,In_119);
nand U265 (N_265,In_393,In_656);
and U266 (N_266,In_4,In_598);
nand U267 (N_267,In_275,In_421);
and U268 (N_268,In_670,In_185);
nand U269 (N_269,In_612,In_42);
and U270 (N_270,In_134,In_728);
or U271 (N_271,In_603,In_703);
nor U272 (N_272,In_32,In_53);
nand U273 (N_273,In_99,In_26);
nor U274 (N_274,In_525,In_633);
and U275 (N_275,In_102,In_726);
nor U276 (N_276,In_390,In_358);
or U277 (N_277,In_658,In_555);
and U278 (N_278,In_528,In_94);
and U279 (N_279,In_376,In_306);
or U280 (N_280,In_387,In_545);
xor U281 (N_281,In_348,In_267);
nand U282 (N_282,In_485,In_157);
nand U283 (N_283,In_490,In_748);
or U284 (N_284,In_430,In_680);
nor U285 (N_285,In_39,In_540);
nor U286 (N_286,In_432,In_733);
nor U287 (N_287,In_712,In_704);
nand U288 (N_288,In_329,In_292);
nand U289 (N_289,In_429,In_456);
and U290 (N_290,In_45,In_434);
nand U291 (N_291,In_366,In_664);
and U292 (N_292,In_626,In_6);
and U293 (N_293,In_518,In_323);
or U294 (N_294,In_480,In_686);
nor U295 (N_295,In_254,In_605);
nand U296 (N_296,In_202,In_305);
nor U297 (N_297,In_180,In_531);
nor U298 (N_298,In_143,In_87);
nand U299 (N_299,In_328,In_347);
nand U300 (N_300,In_462,In_478);
and U301 (N_301,In_303,In_623);
or U302 (N_302,In_196,In_610);
nor U303 (N_303,In_560,In_529);
nand U304 (N_304,In_644,In_731);
and U305 (N_305,In_317,In_326);
nor U306 (N_306,In_232,In_29);
and U307 (N_307,In_484,In_371);
nand U308 (N_308,In_412,In_2);
nand U309 (N_309,In_592,In_504);
nor U310 (N_310,In_351,In_287);
or U311 (N_311,In_145,In_183);
and U312 (N_312,In_558,In_424);
nand U313 (N_313,In_673,In_61);
nor U314 (N_314,In_694,In_124);
nand U315 (N_315,In_599,In_514);
and U316 (N_316,In_125,In_111);
or U317 (N_317,In_618,In_409);
or U318 (N_318,In_377,In_0);
nand U319 (N_319,In_297,In_486);
nor U320 (N_320,In_44,In_725);
and U321 (N_321,In_339,In_661);
or U322 (N_322,In_106,In_262);
nor U323 (N_323,In_378,In_407);
nor U324 (N_324,In_174,In_138);
or U325 (N_325,In_583,In_448);
nand U326 (N_326,In_213,In_187);
and U327 (N_327,In_637,In_21);
nor U328 (N_328,In_634,In_211);
or U329 (N_329,In_505,In_357);
or U330 (N_330,In_162,In_238);
nand U331 (N_331,In_488,In_385);
and U332 (N_332,In_179,In_381);
and U333 (N_333,In_362,In_298);
and U334 (N_334,In_417,In_181);
nor U335 (N_335,In_146,In_246);
and U336 (N_336,In_127,In_619);
and U337 (N_337,In_628,In_290);
and U338 (N_338,In_524,In_722);
or U339 (N_339,In_252,In_97);
nand U340 (N_340,In_10,In_522);
nor U341 (N_341,In_743,In_666);
or U342 (N_342,In_91,In_269);
or U343 (N_343,In_355,In_285);
nand U344 (N_344,In_709,In_132);
and U345 (N_345,In_668,In_338);
xnor U346 (N_346,In_291,In_276);
xnor U347 (N_347,In_494,In_200);
and U348 (N_348,In_442,In_563);
nor U349 (N_349,In_300,In_62);
nor U350 (N_350,In_566,In_334);
and U351 (N_351,In_17,In_330);
and U352 (N_352,In_723,In_212);
nand U353 (N_353,In_568,In_440);
nor U354 (N_354,In_286,In_542);
nor U355 (N_355,In_158,In_161);
or U356 (N_356,In_188,In_55);
nand U357 (N_357,In_445,In_735);
and U358 (N_358,In_684,In_344);
nand U359 (N_359,In_289,In_197);
nor U360 (N_360,In_144,In_250);
nand U361 (N_361,In_675,In_415);
nor U362 (N_362,In_380,In_223);
nor U363 (N_363,In_707,In_745);
nand U364 (N_364,In_126,In_231);
or U365 (N_365,In_193,In_413);
and U366 (N_366,In_746,In_88);
nand U367 (N_367,In_13,In_302);
or U368 (N_368,In_609,In_580);
nor U369 (N_369,In_616,In_736);
nor U370 (N_370,In_63,In_536);
nor U371 (N_371,In_201,In_660);
nor U372 (N_372,In_706,In_472);
or U373 (N_373,In_216,In_208);
nor U374 (N_374,In_345,In_172);
and U375 (N_375,In_281,In_335);
and U376 (N_376,In_576,In_500);
or U377 (N_377,In_15,In_39);
or U378 (N_378,In_44,In_339);
nand U379 (N_379,In_292,In_331);
or U380 (N_380,In_134,In_596);
nor U381 (N_381,In_619,In_6);
and U382 (N_382,In_211,In_500);
and U383 (N_383,In_350,In_563);
nand U384 (N_384,In_28,In_207);
nand U385 (N_385,In_275,In_104);
nand U386 (N_386,In_223,In_623);
nor U387 (N_387,In_270,In_411);
and U388 (N_388,In_183,In_569);
or U389 (N_389,In_478,In_530);
or U390 (N_390,In_596,In_481);
nor U391 (N_391,In_185,In_746);
or U392 (N_392,In_34,In_204);
nand U393 (N_393,In_427,In_508);
and U394 (N_394,In_496,In_714);
and U395 (N_395,In_613,In_266);
nand U396 (N_396,In_175,In_637);
nor U397 (N_397,In_645,In_416);
or U398 (N_398,In_288,In_51);
nor U399 (N_399,In_471,In_301);
nor U400 (N_400,In_322,In_494);
nand U401 (N_401,In_38,In_476);
nor U402 (N_402,In_217,In_458);
or U403 (N_403,In_53,In_395);
and U404 (N_404,In_600,In_3);
or U405 (N_405,In_532,In_14);
or U406 (N_406,In_664,In_314);
and U407 (N_407,In_174,In_109);
or U408 (N_408,In_105,In_570);
nand U409 (N_409,In_682,In_260);
or U410 (N_410,In_2,In_257);
or U411 (N_411,In_630,In_98);
nand U412 (N_412,In_596,In_184);
and U413 (N_413,In_208,In_127);
nor U414 (N_414,In_459,In_96);
nor U415 (N_415,In_49,In_418);
or U416 (N_416,In_734,In_115);
or U417 (N_417,In_249,In_30);
or U418 (N_418,In_406,In_324);
and U419 (N_419,In_67,In_430);
and U420 (N_420,In_238,In_641);
nand U421 (N_421,In_594,In_339);
and U422 (N_422,In_443,In_262);
nand U423 (N_423,In_81,In_99);
and U424 (N_424,In_190,In_347);
xor U425 (N_425,In_25,In_106);
and U426 (N_426,In_14,In_715);
nor U427 (N_427,In_577,In_87);
nor U428 (N_428,In_466,In_450);
nand U429 (N_429,In_707,In_604);
or U430 (N_430,In_544,In_274);
nand U431 (N_431,In_439,In_744);
nand U432 (N_432,In_335,In_357);
nand U433 (N_433,In_435,In_726);
or U434 (N_434,In_513,In_545);
or U435 (N_435,In_321,In_710);
or U436 (N_436,In_563,In_55);
nor U437 (N_437,In_95,In_399);
or U438 (N_438,In_520,In_321);
nor U439 (N_439,In_645,In_412);
and U440 (N_440,In_591,In_345);
nor U441 (N_441,In_168,In_77);
or U442 (N_442,In_619,In_332);
nand U443 (N_443,In_225,In_52);
nand U444 (N_444,In_504,In_631);
or U445 (N_445,In_601,In_683);
nor U446 (N_446,In_218,In_470);
or U447 (N_447,In_232,In_159);
nand U448 (N_448,In_506,In_455);
or U449 (N_449,In_361,In_587);
nand U450 (N_450,In_402,In_543);
or U451 (N_451,In_504,In_351);
nor U452 (N_452,In_82,In_436);
nand U453 (N_453,In_536,In_565);
or U454 (N_454,In_136,In_587);
nand U455 (N_455,In_410,In_440);
nand U456 (N_456,In_399,In_697);
nand U457 (N_457,In_96,In_392);
and U458 (N_458,In_177,In_732);
nor U459 (N_459,In_565,In_169);
nand U460 (N_460,In_575,In_343);
nand U461 (N_461,In_72,In_722);
and U462 (N_462,In_401,In_429);
or U463 (N_463,In_262,In_412);
nand U464 (N_464,In_485,In_474);
nand U465 (N_465,In_157,In_679);
or U466 (N_466,In_23,In_469);
or U467 (N_467,In_43,In_532);
and U468 (N_468,In_473,In_506);
nand U469 (N_469,In_239,In_29);
and U470 (N_470,In_452,In_496);
nor U471 (N_471,In_432,In_201);
nor U472 (N_472,In_616,In_664);
xor U473 (N_473,In_384,In_666);
nor U474 (N_474,In_96,In_299);
and U475 (N_475,In_298,In_51);
nor U476 (N_476,In_367,In_188);
nand U477 (N_477,In_539,In_405);
and U478 (N_478,In_259,In_587);
and U479 (N_479,In_212,In_389);
nand U480 (N_480,In_377,In_18);
and U481 (N_481,In_420,In_286);
or U482 (N_482,In_253,In_562);
nand U483 (N_483,In_263,In_351);
nor U484 (N_484,In_437,In_189);
nand U485 (N_485,In_332,In_165);
and U486 (N_486,In_127,In_87);
nor U487 (N_487,In_398,In_237);
and U488 (N_488,In_171,In_567);
or U489 (N_489,In_35,In_541);
and U490 (N_490,In_707,In_527);
or U491 (N_491,In_136,In_541);
and U492 (N_492,In_669,In_230);
nor U493 (N_493,In_135,In_740);
nand U494 (N_494,In_111,In_11);
or U495 (N_495,In_483,In_24);
or U496 (N_496,In_740,In_23);
and U497 (N_497,In_63,In_318);
nand U498 (N_498,In_33,In_380);
or U499 (N_499,In_175,In_568);
and U500 (N_500,In_411,In_172);
nor U501 (N_501,In_97,In_419);
or U502 (N_502,In_632,In_680);
and U503 (N_503,In_215,In_371);
and U504 (N_504,In_270,In_477);
or U505 (N_505,In_58,In_54);
nor U506 (N_506,In_122,In_472);
or U507 (N_507,In_274,In_429);
and U508 (N_508,In_691,In_267);
xnor U509 (N_509,In_681,In_633);
and U510 (N_510,In_563,In_677);
or U511 (N_511,In_562,In_581);
or U512 (N_512,In_221,In_349);
and U513 (N_513,In_504,In_253);
nand U514 (N_514,In_680,In_479);
nor U515 (N_515,In_104,In_261);
nand U516 (N_516,In_197,In_413);
nor U517 (N_517,In_108,In_42);
or U518 (N_518,In_294,In_599);
nand U519 (N_519,In_120,In_240);
nor U520 (N_520,In_26,In_539);
nor U521 (N_521,In_492,In_146);
nand U522 (N_522,In_403,In_0);
nor U523 (N_523,In_494,In_260);
or U524 (N_524,In_55,In_66);
nor U525 (N_525,In_69,In_453);
or U526 (N_526,In_720,In_5);
or U527 (N_527,In_326,In_312);
or U528 (N_528,In_273,In_148);
nor U529 (N_529,In_146,In_479);
or U530 (N_530,In_479,In_249);
nand U531 (N_531,In_690,In_651);
nand U532 (N_532,In_626,In_71);
nand U533 (N_533,In_577,In_154);
and U534 (N_534,In_593,In_668);
and U535 (N_535,In_199,In_10);
or U536 (N_536,In_122,In_633);
or U537 (N_537,In_49,In_39);
nand U538 (N_538,In_165,In_457);
and U539 (N_539,In_427,In_30);
xnor U540 (N_540,In_269,In_12);
and U541 (N_541,In_187,In_174);
and U542 (N_542,In_281,In_638);
nand U543 (N_543,In_468,In_598);
nor U544 (N_544,In_25,In_434);
or U545 (N_545,In_138,In_604);
nand U546 (N_546,In_476,In_378);
nor U547 (N_547,In_641,In_121);
and U548 (N_548,In_331,In_125);
nor U549 (N_549,In_473,In_244);
nor U550 (N_550,In_594,In_379);
nor U551 (N_551,In_185,In_580);
or U552 (N_552,In_676,In_598);
and U553 (N_553,In_445,In_344);
and U554 (N_554,In_363,In_344);
or U555 (N_555,In_741,In_261);
or U556 (N_556,In_27,In_253);
nor U557 (N_557,In_125,In_399);
and U558 (N_558,In_487,In_76);
nor U559 (N_559,In_309,In_344);
or U560 (N_560,In_504,In_67);
or U561 (N_561,In_338,In_327);
nand U562 (N_562,In_510,In_60);
nand U563 (N_563,In_480,In_82);
nand U564 (N_564,In_265,In_326);
nor U565 (N_565,In_211,In_44);
or U566 (N_566,In_628,In_746);
and U567 (N_567,In_712,In_348);
or U568 (N_568,In_713,In_489);
nand U569 (N_569,In_4,In_123);
and U570 (N_570,In_623,In_452);
nand U571 (N_571,In_355,In_564);
nor U572 (N_572,In_530,In_275);
or U573 (N_573,In_276,In_378);
nand U574 (N_574,In_204,In_268);
or U575 (N_575,In_693,In_659);
nand U576 (N_576,In_272,In_60);
nand U577 (N_577,In_154,In_546);
and U578 (N_578,In_553,In_196);
or U579 (N_579,In_171,In_164);
nand U580 (N_580,In_652,In_608);
or U581 (N_581,In_548,In_167);
and U582 (N_582,In_358,In_628);
nor U583 (N_583,In_155,In_665);
nor U584 (N_584,In_656,In_714);
nand U585 (N_585,In_160,In_252);
nand U586 (N_586,In_367,In_267);
nor U587 (N_587,In_536,In_299);
nand U588 (N_588,In_209,In_600);
or U589 (N_589,In_499,In_550);
nand U590 (N_590,In_603,In_246);
or U591 (N_591,In_679,In_387);
or U592 (N_592,In_703,In_577);
and U593 (N_593,In_19,In_165);
nand U594 (N_594,In_14,In_300);
and U595 (N_595,In_656,In_373);
and U596 (N_596,In_615,In_666);
nor U597 (N_597,In_167,In_605);
and U598 (N_598,In_47,In_182);
nand U599 (N_599,In_266,In_701);
or U600 (N_600,In_292,In_702);
or U601 (N_601,In_396,In_350);
nor U602 (N_602,In_18,In_8);
nand U603 (N_603,In_365,In_168);
and U604 (N_604,In_366,In_399);
nor U605 (N_605,In_309,In_647);
and U606 (N_606,In_339,In_546);
and U607 (N_607,In_63,In_614);
nand U608 (N_608,In_502,In_654);
and U609 (N_609,In_476,In_281);
or U610 (N_610,In_258,In_382);
and U611 (N_611,In_94,In_33);
and U612 (N_612,In_355,In_626);
or U613 (N_613,In_663,In_323);
or U614 (N_614,In_126,In_139);
nor U615 (N_615,In_152,In_129);
and U616 (N_616,In_212,In_296);
nor U617 (N_617,In_328,In_312);
nor U618 (N_618,In_355,In_562);
and U619 (N_619,In_322,In_82);
and U620 (N_620,In_157,In_59);
nor U621 (N_621,In_540,In_285);
or U622 (N_622,In_482,In_656);
and U623 (N_623,In_677,In_674);
and U624 (N_624,In_485,In_427);
nor U625 (N_625,In_148,In_324);
nand U626 (N_626,In_159,In_366);
or U627 (N_627,In_81,In_140);
and U628 (N_628,In_12,In_735);
or U629 (N_629,In_73,In_308);
nand U630 (N_630,In_436,In_272);
nor U631 (N_631,In_71,In_623);
or U632 (N_632,In_456,In_150);
or U633 (N_633,In_502,In_551);
nor U634 (N_634,In_576,In_327);
nor U635 (N_635,In_214,In_283);
nand U636 (N_636,In_581,In_10);
or U637 (N_637,In_314,In_722);
xor U638 (N_638,In_383,In_686);
xnor U639 (N_639,In_733,In_141);
nor U640 (N_640,In_258,In_473);
nor U641 (N_641,In_304,In_495);
or U642 (N_642,In_524,In_291);
nor U643 (N_643,In_592,In_203);
nor U644 (N_644,In_327,In_351);
or U645 (N_645,In_478,In_725);
nand U646 (N_646,In_288,In_147);
and U647 (N_647,In_584,In_210);
or U648 (N_648,In_696,In_735);
or U649 (N_649,In_313,In_520);
xor U650 (N_650,In_220,In_67);
and U651 (N_651,In_351,In_738);
nand U652 (N_652,In_464,In_75);
and U653 (N_653,In_592,In_475);
nand U654 (N_654,In_293,In_5);
nand U655 (N_655,In_189,In_11);
nand U656 (N_656,In_31,In_542);
or U657 (N_657,In_420,In_591);
nand U658 (N_658,In_576,In_376);
and U659 (N_659,In_459,In_619);
nor U660 (N_660,In_390,In_25);
nand U661 (N_661,In_453,In_203);
nand U662 (N_662,In_379,In_334);
and U663 (N_663,In_299,In_231);
nand U664 (N_664,In_21,In_130);
nor U665 (N_665,In_454,In_257);
nand U666 (N_666,In_613,In_514);
and U667 (N_667,In_223,In_78);
and U668 (N_668,In_468,In_548);
or U669 (N_669,In_467,In_449);
and U670 (N_670,In_126,In_502);
nand U671 (N_671,In_25,In_192);
nand U672 (N_672,In_303,In_390);
or U673 (N_673,In_97,In_326);
and U674 (N_674,In_193,In_401);
nor U675 (N_675,In_528,In_651);
nor U676 (N_676,In_661,In_334);
xor U677 (N_677,In_387,In_478);
nand U678 (N_678,In_510,In_113);
nor U679 (N_679,In_571,In_731);
nor U680 (N_680,In_614,In_442);
nand U681 (N_681,In_454,In_183);
nor U682 (N_682,In_231,In_311);
or U683 (N_683,In_367,In_475);
xnor U684 (N_684,In_378,In_488);
nand U685 (N_685,In_397,In_211);
nand U686 (N_686,In_423,In_338);
nor U687 (N_687,In_520,In_146);
nor U688 (N_688,In_628,In_321);
nor U689 (N_689,In_543,In_8);
nor U690 (N_690,In_307,In_33);
or U691 (N_691,In_434,In_380);
and U692 (N_692,In_488,In_468);
or U693 (N_693,In_385,In_293);
or U694 (N_694,In_32,In_290);
nor U695 (N_695,In_244,In_31);
and U696 (N_696,In_199,In_352);
nand U697 (N_697,In_465,In_332);
and U698 (N_698,In_318,In_356);
or U699 (N_699,In_379,In_76);
xor U700 (N_700,In_261,In_437);
nand U701 (N_701,In_403,In_411);
and U702 (N_702,In_211,In_252);
or U703 (N_703,In_383,In_231);
nor U704 (N_704,In_746,In_75);
or U705 (N_705,In_549,In_620);
nand U706 (N_706,In_197,In_492);
nor U707 (N_707,In_27,In_206);
nor U708 (N_708,In_152,In_638);
nor U709 (N_709,In_648,In_85);
and U710 (N_710,In_405,In_364);
nand U711 (N_711,In_221,In_319);
nand U712 (N_712,In_276,In_351);
or U713 (N_713,In_629,In_140);
or U714 (N_714,In_731,In_189);
or U715 (N_715,In_592,In_429);
nand U716 (N_716,In_0,In_158);
and U717 (N_717,In_449,In_78);
or U718 (N_718,In_255,In_691);
and U719 (N_719,In_633,In_84);
and U720 (N_720,In_456,In_57);
or U721 (N_721,In_198,In_53);
or U722 (N_722,In_617,In_71);
and U723 (N_723,In_388,In_121);
nor U724 (N_724,In_416,In_95);
nor U725 (N_725,In_121,In_430);
nor U726 (N_726,In_638,In_746);
and U727 (N_727,In_60,In_88);
or U728 (N_728,In_609,In_205);
and U729 (N_729,In_22,In_114);
or U730 (N_730,In_275,In_59);
nand U731 (N_731,In_549,In_496);
nand U732 (N_732,In_521,In_252);
or U733 (N_733,In_436,In_602);
and U734 (N_734,In_496,In_573);
and U735 (N_735,In_501,In_456);
nand U736 (N_736,In_685,In_467);
or U737 (N_737,In_728,In_6);
or U738 (N_738,In_165,In_716);
and U739 (N_739,In_706,In_714);
nor U740 (N_740,In_58,In_330);
nand U741 (N_741,In_695,In_454);
and U742 (N_742,In_449,In_504);
and U743 (N_743,In_259,In_127);
nor U744 (N_744,In_313,In_659);
nand U745 (N_745,In_414,In_224);
or U746 (N_746,In_710,In_643);
or U747 (N_747,In_332,In_166);
nor U748 (N_748,In_465,In_225);
nand U749 (N_749,In_397,In_214);
or U750 (N_750,In_186,In_184);
nand U751 (N_751,In_305,In_629);
nor U752 (N_752,In_707,In_363);
nand U753 (N_753,In_442,In_536);
nand U754 (N_754,In_284,In_426);
nand U755 (N_755,In_568,In_287);
or U756 (N_756,In_443,In_5);
nor U757 (N_757,In_423,In_398);
nor U758 (N_758,In_264,In_16);
nor U759 (N_759,In_740,In_720);
and U760 (N_760,In_623,In_578);
and U761 (N_761,In_233,In_544);
xor U762 (N_762,In_318,In_90);
nor U763 (N_763,In_503,In_419);
and U764 (N_764,In_625,In_685);
and U765 (N_765,In_629,In_554);
and U766 (N_766,In_387,In_92);
nand U767 (N_767,In_315,In_280);
nor U768 (N_768,In_370,In_733);
or U769 (N_769,In_82,In_698);
xor U770 (N_770,In_33,In_558);
and U771 (N_771,In_579,In_535);
nand U772 (N_772,In_575,In_486);
and U773 (N_773,In_309,In_326);
or U774 (N_774,In_269,In_109);
nand U775 (N_775,In_225,In_137);
nor U776 (N_776,In_548,In_39);
nor U777 (N_777,In_605,In_562);
nand U778 (N_778,In_245,In_107);
nor U779 (N_779,In_713,In_578);
and U780 (N_780,In_407,In_687);
nand U781 (N_781,In_108,In_162);
or U782 (N_782,In_521,In_253);
nor U783 (N_783,In_447,In_77);
and U784 (N_784,In_23,In_212);
and U785 (N_785,In_546,In_107);
nor U786 (N_786,In_639,In_601);
nor U787 (N_787,In_290,In_6);
nor U788 (N_788,In_273,In_666);
and U789 (N_789,In_484,In_649);
nand U790 (N_790,In_90,In_395);
nor U791 (N_791,In_207,In_143);
nor U792 (N_792,In_635,In_423);
or U793 (N_793,In_647,In_419);
or U794 (N_794,In_351,In_665);
and U795 (N_795,In_0,In_458);
nand U796 (N_796,In_14,In_709);
nand U797 (N_797,In_733,In_573);
nand U798 (N_798,In_277,In_734);
nand U799 (N_799,In_617,In_153);
nor U800 (N_800,In_337,In_456);
xnor U801 (N_801,In_618,In_421);
nor U802 (N_802,In_548,In_234);
nand U803 (N_803,In_656,In_553);
or U804 (N_804,In_226,In_264);
and U805 (N_805,In_486,In_349);
or U806 (N_806,In_27,In_628);
or U807 (N_807,In_378,In_483);
or U808 (N_808,In_68,In_307);
or U809 (N_809,In_408,In_684);
and U810 (N_810,In_679,In_296);
or U811 (N_811,In_686,In_31);
nand U812 (N_812,In_136,In_657);
xnor U813 (N_813,In_150,In_253);
nand U814 (N_814,In_284,In_200);
nor U815 (N_815,In_740,In_577);
nor U816 (N_816,In_44,In_299);
or U817 (N_817,In_12,In_648);
or U818 (N_818,In_367,In_296);
nand U819 (N_819,In_67,In_382);
and U820 (N_820,In_249,In_521);
or U821 (N_821,In_427,In_207);
and U822 (N_822,In_611,In_603);
and U823 (N_823,In_106,In_0);
or U824 (N_824,In_417,In_738);
and U825 (N_825,In_422,In_19);
or U826 (N_826,In_95,In_53);
nor U827 (N_827,In_506,In_435);
nor U828 (N_828,In_41,In_90);
nand U829 (N_829,In_542,In_268);
nand U830 (N_830,In_688,In_426);
nand U831 (N_831,In_261,In_246);
and U832 (N_832,In_734,In_345);
xor U833 (N_833,In_408,In_215);
and U834 (N_834,In_108,In_260);
nor U835 (N_835,In_604,In_346);
or U836 (N_836,In_704,In_648);
nor U837 (N_837,In_518,In_395);
nand U838 (N_838,In_623,In_688);
or U839 (N_839,In_253,In_104);
or U840 (N_840,In_345,In_211);
nand U841 (N_841,In_45,In_264);
and U842 (N_842,In_509,In_460);
nor U843 (N_843,In_585,In_471);
or U844 (N_844,In_641,In_660);
or U845 (N_845,In_242,In_310);
nand U846 (N_846,In_276,In_341);
nand U847 (N_847,In_478,In_243);
nand U848 (N_848,In_646,In_684);
or U849 (N_849,In_441,In_568);
nand U850 (N_850,In_634,In_11);
or U851 (N_851,In_251,In_46);
nand U852 (N_852,In_565,In_174);
or U853 (N_853,In_732,In_155);
nor U854 (N_854,In_137,In_325);
nand U855 (N_855,In_236,In_325);
or U856 (N_856,In_45,In_514);
and U857 (N_857,In_40,In_673);
and U858 (N_858,In_114,In_450);
nand U859 (N_859,In_501,In_363);
nor U860 (N_860,In_5,In_749);
and U861 (N_861,In_394,In_507);
and U862 (N_862,In_484,In_604);
or U863 (N_863,In_178,In_322);
nor U864 (N_864,In_618,In_370);
or U865 (N_865,In_105,In_48);
and U866 (N_866,In_515,In_239);
nand U867 (N_867,In_716,In_61);
and U868 (N_868,In_645,In_486);
or U869 (N_869,In_708,In_187);
or U870 (N_870,In_240,In_443);
nand U871 (N_871,In_358,In_182);
nand U872 (N_872,In_444,In_229);
or U873 (N_873,In_396,In_225);
nand U874 (N_874,In_608,In_262);
nor U875 (N_875,In_153,In_450);
nand U876 (N_876,In_280,In_738);
or U877 (N_877,In_85,In_734);
or U878 (N_878,In_521,In_62);
nor U879 (N_879,In_6,In_235);
and U880 (N_880,In_288,In_182);
nor U881 (N_881,In_441,In_156);
nand U882 (N_882,In_499,In_692);
nand U883 (N_883,In_447,In_246);
or U884 (N_884,In_411,In_323);
nor U885 (N_885,In_475,In_527);
and U886 (N_886,In_85,In_625);
nor U887 (N_887,In_249,In_365);
nand U888 (N_888,In_544,In_549);
and U889 (N_889,In_536,In_735);
or U890 (N_890,In_350,In_585);
or U891 (N_891,In_141,In_673);
nor U892 (N_892,In_381,In_578);
and U893 (N_893,In_544,In_223);
and U894 (N_894,In_364,In_207);
nand U895 (N_895,In_453,In_154);
and U896 (N_896,In_648,In_631);
and U897 (N_897,In_523,In_1);
nand U898 (N_898,In_241,In_289);
and U899 (N_899,In_500,In_473);
or U900 (N_900,In_281,In_255);
nand U901 (N_901,In_56,In_641);
or U902 (N_902,In_587,In_271);
nand U903 (N_903,In_645,In_316);
and U904 (N_904,In_87,In_184);
nand U905 (N_905,In_716,In_614);
and U906 (N_906,In_121,In_368);
and U907 (N_907,In_304,In_169);
nor U908 (N_908,In_660,In_227);
nand U909 (N_909,In_743,In_534);
and U910 (N_910,In_234,In_361);
xor U911 (N_911,In_658,In_396);
and U912 (N_912,In_259,In_456);
and U913 (N_913,In_488,In_373);
nor U914 (N_914,In_149,In_423);
nand U915 (N_915,In_49,In_175);
nor U916 (N_916,In_589,In_442);
or U917 (N_917,In_488,In_333);
nand U918 (N_918,In_344,In_605);
or U919 (N_919,In_479,In_749);
nor U920 (N_920,In_540,In_717);
or U921 (N_921,In_203,In_460);
nor U922 (N_922,In_618,In_325);
nor U923 (N_923,In_435,In_183);
nand U924 (N_924,In_350,In_493);
or U925 (N_925,In_456,In_710);
nor U926 (N_926,In_376,In_520);
xor U927 (N_927,In_677,In_154);
nand U928 (N_928,In_718,In_507);
nor U929 (N_929,In_9,In_35);
nand U930 (N_930,In_40,In_741);
nor U931 (N_931,In_47,In_635);
or U932 (N_932,In_247,In_221);
and U933 (N_933,In_746,In_356);
or U934 (N_934,In_109,In_429);
nor U935 (N_935,In_171,In_97);
or U936 (N_936,In_257,In_370);
and U937 (N_937,In_711,In_200);
and U938 (N_938,In_222,In_743);
nand U939 (N_939,In_738,In_670);
or U940 (N_940,In_486,In_284);
and U941 (N_941,In_396,In_85);
nand U942 (N_942,In_684,In_596);
or U943 (N_943,In_237,In_180);
nand U944 (N_944,In_263,In_280);
or U945 (N_945,In_572,In_206);
nor U946 (N_946,In_287,In_721);
nand U947 (N_947,In_711,In_304);
nand U948 (N_948,In_169,In_274);
and U949 (N_949,In_655,In_557);
nand U950 (N_950,In_295,In_214);
and U951 (N_951,In_509,In_414);
or U952 (N_952,In_304,In_76);
nor U953 (N_953,In_631,In_417);
or U954 (N_954,In_570,In_246);
or U955 (N_955,In_418,In_208);
nand U956 (N_956,In_449,In_415);
nor U957 (N_957,In_259,In_441);
or U958 (N_958,In_615,In_227);
nor U959 (N_959,In_294,In_38);
and U960 (N_960,In_301,In_310);
or U961 (N_961,In_747,In_575);
and U962 (N_962,In_267,In_244);
and U963 (N_963,In_353,In_565);
or U964 (N_964,In_289,In_219);
and U965 (N_965,In_591,In_418);
nand U966 (N_966,In_467,In_411);
or U967 (N_967,In_151,In_595);
or U968 (N_968,In_700,In_453);
or U969 (N_969,In_644,In_664);
or U970 (N_970,In_364,In_0);
or U971 (N_971,In_227,In_708);
nor U972 (N_972,In_429,In_643);
nor U973 (N_973,In_700,In_277);
nand U974 (N_974,In_385,In_160);
nand U975 (N_975,In_529,In_589);
or U976 (N_976,In_538,In_634);
and U977 (N_977,In_445,In_254);
xor U978 (N_978,In_187,In_324);
or U979 (N_979,In_588,In_568);
and U980 (N_980,In_188,In_596);
or U981 (N_981,In_115,In_249);
or U982 (N_982,In_94,In_99);
nand U983 (N_983,In_401,In_491);
nand U984 (N_984,In_682,In_622);
or U985 (N_985,In_448,In_169);
nor U986 (N_986,In_67,In_243);
nor U987 (N_987,In_685,In_344);
nand U988 (N_988,In_527,In_452);
nor U989 (N_989,In_692,In_733);
nor U990 (N_990,In_731,In_364);
nand U991 (N_991,In_145,In_638);
and U992 (N_992,In_231,In_355);
nor U993 (N_993,In_455,In_229);
nor U994 (N_994,In_422,In_489);
and U995 (N_995,In_245,In_636);
or U996 (N_996,In_431,In_287);
and U997 (N_997,In_46,In_210);
and U998 (N_998,In_483,In_549);
and U999 (N_999,In_665,In_444);
nor U1000 (N_1000,N_193,N_243);
or U1001 (N_1001,N_276,N_20);
or U1002 (N_1002,N_523,N_562);
nand U1003 (N_1003,N_524,N_568);
and U1004 (N_1004,N_679,N_170);
or U1005 (N_1005,N_355,N_596);
or U1006 (N_1006,N_39,N_196);
nand U1007 (N_1007,N_538,N_379);
nand U1008 (N_1008,N_438,N_471);
or U1009 (N_1009,N_201,N_483);
nor U1010 (N_1010,N_18,N_305);
nor U1011 (N_1011,N_927,N_966);
nand U1012 (N_1012,N_179,N_768);
nand U1013 (N_1013,N_142,N_623);
nand U1014 (N_1014,N_628,N_751);
nand U1015 (N_1015,N_718,N_332);
xor U1016 (N_1016,N_990,N_485);
nor U1017 (N_1017,N_235,N_865);
nor U1018 (N_1018,N_463,N_534);
nor U1019 (N_1019,N_748,N_656);
nor U1020 (N_1020,N_869,N_51);
or U1021 (N_1021,N_260,N_694);
nand U1022 (N_1022,N_324,N_896);
and U1023 (N_1023,N_863,N_653);
nor U1024 (N_1024,N_610,N_849);
or U1025 (N_1025,N_635,N_868);
and U1026 (N_1026,N_116,N_644);
nor U1027 (N_1027,N_77,N_648);
and U1028 (N_1028,N_634,N_950);
nor U1029 (N_1029,N_25,N_108);
nand U1030 (N_1030,N_331,N_970);
nor U1031 (N_1031,N_111,N_346);
nand U1032 (N_1032,N_21,N_289);
or U1033 (N_1033,N_167,N_78);
or U1034 (N_1034,N_241,N_302);
or U1035 (N_1035,N_301,N_754);
xnor U1036 (N_1036,N_758,N_282);
nand U1037 (N_1037,N_627,N_238);
and U1038 (N_1038,N_360,N_531);
and U1039 (N_1039,N_873,N_808);
nand U1040 (N_1040,N_707,N_138);
and U1041 (N_1041,N_382,N_5);
or U1042 (N_1042,N_746,N_233);
nand U1043 (N_1043,N_573,N_174);
nor U1044 (N_1044,N_685,N_861);
nand U1045 (N_1045,N_587,N_398);
or U1046 (N_1046,N_197,N_969);
or U1047 (N_1047,N_456,N_124);
nand U1048 (N_1048,N_971,N_749);
nor U1049 (N_1049,N_689,N_383);
or U1050 (N_1050,N_242,N_986);
or U1051 (N_1051,N_390,N_487);
xnor U1052 (N_1052,N_886,N_350);
or U1053 (N_1053,N_684,N_900);
nor U1054 (N_1054,N_821,N_697);
xor U1055 (N_1055,N_838,N_774);
nor U1056 (N_1056,N_424,N_829);
nor U1057 (N_1057,N_10,N_572);
nor U1058 (N_1058,N_31,N_513);
or U1059 (N_1059,N_56,N_545);
or U1060 (N_1060,N_431,N_52);
nand U1061 (N_1061,N_614,N_95);
and U1062 (N_1062,N_140,N_472);
nand U1063 (N_1063,N_102,N_269);
and U1064 (N_1064,N_207,N_100);
and U1065 (N_1065,N_680,N_586);
xor U1066 (N_1066,N_294,N_361);
and U1067 (N_1067,N_367,N_191);
nand U1068 (N_1068,N_760,N_880);
or U1069 (N_1069,N_901,N_629);
or U1070 (N_1070,N_581,N_957);
nand U1071 (N_1071,N_19,N_80);
or U1072 (N_1072,N_622,N_267);
or U1073 (N_1073,N_359,N_908);
nor U1074 (N_1074,N_701,N_521);
and U1075 (N_1075,N_882,N_212);
or U1076 (N_1076,N_642,N_668);
and U1077 (N_1077,N_387,N_700);
or U1078 (N_1078,N_507,N_248);
nand U1079 (N_1079,N_539,N_834);
and U1080 (N_1080,N_351,N_410);
nor U1081 (N_1081,N_29,N_226);
nand U1082 (N_1082,N_724,N_625);
nand U1083 (N_1083,N_293,N_532);
and U1084 (N_1084,N_613,N_744);
nand U1085 (N_1085,N_696,N_322);
or U1086 (N_1086,N_951,N_512);
nand U1087 (N_1087,N_291,N_203);
xnor U1088 (N_1088,N_711,N_736);
or U1089 (N_1089,N_32,N_344);
and U1090 (N_1090,N_63,N_921);
or U1091 (N_1091,N_475,N_376);
and U1092 (N_1092,N_666,N_851);
nor U1093 (N_1093,N_594,N_582);
and U1094 (N_1094,N_395,N_989);
and U1095 (N_1095,N_27,N_283);
nor U1096 (N_1096,N_255,N_339);
and U1097 (N_1097,N_418,N_998);
and U1098 (N_1098,N_576,N_725);
and U1099 (N_1099,N_476,N_103);
nor U1100 (N_1100,N_541,N_416);
nor U1101 (N_1101,N_415,N_738);
xor U1102 (N_1102,N_369,N_45);
nand U1103 (N_1103,N_13,N_447);
or U1104 (N_1104,N_854,N_683);
and U1105 (N_1105,N_178,N_617);
or U1106 (N_1106,N_780,N_953);
and U1107 (N_1107,N_765,N_200);
nor U1108 (N_1108,N_514,N_783);
nor U1109 (N_1109,N_368,N_540);
nand U1110 (N_1110,N_828,N_917);
nand U1111 (N_1111,N_944,N_57);
or U1112 (N_1112,N_631,N_352);
or U1113 (N_1113,N_239,N_673);
nor U1114 (N_1114,N_505,N_954);
or U1115 (N_1115,N_776,N_816);
nor U1116 (N_1116,N_402,N_584);
and U1117 (N_1117,N_389,N_589);
nor U1118 (N_1118,N_598,N_775);
and U1119 (N_1119,N_552,N_354);
or U1120 (N_1120,N_872,N_947);
nand U1121 (N_1121,N_396,N_399);
or U1122 (N_1122,N_37,N_364);
or U1123 (N_1123,N_356,N_48);
and U1124 (N_1124,N_606,N_640);
nand U1125 (N_1125,N_789,N_669);
and U1126 (N_1126,N_934,N_47);
nor U1127 (N_1127,N_187,N_727);
or U1128 (N_1128,N_114,N_244);
or U1129 (N_1129,N_722,N_348);
and U1130 (N_1130,N_68,N_777);
or U1131 (N_1131,N_563,N_842);
or U1132 (N_1132,N_34,N_4);
nand U1133 (N_1133,N_215,N_509);
nand U1134 (N_1134,N_559,N_61);
nor U1135 (N_1135,N_518,N_793);
and U1136 (N_1136,N_962,N_906);
nor U1137 (N_1137,N_588,N_575);
nor U1138 (N_1138,N_604,N_251);
nand U1139 (N_1139,N_608,N_533);
nand U1140 (N_1140,N_79,N_979);
nor U1141 (N_1141,N_366,N_690);
and U1142 (N_1142,N_747,N_705);
nor U1143 (N_1143,N_188,N_150);
or U1144 (N_1144,N_159,N_151);
nor U1145 (N_1145,N_117,N_497);
and U1146 (N_1146,N_90,N_478);
nand U1147 (N_1147,N_15,N_510);
nand U1148 (N_1148,N_184,N_600);
nor U1149 (N_1149,N_959,N_153);
nor U1150 (N_1150,N_319,N_227);
or U1151 (N_1151,N_826,N_413);
or U1152 (N_1152,N_23,N_479);
and U1153 (N_1153,N_494,N_411);
and U1154 (N_1154,N_466,N_208);
nor U1155 (N_1155,N_155,N_905);
and U1156 (N_1156,N_490,N_735);
nor U1157 (N_1157,N_249,N_246);
nand U1158 (N_1158,N_902,N_770);
nor U1159 (N_1159,N_406,N_473);
nor U1160 (N_1160,N_730,N_655);
and U1161 (N_1161,N_618,N_72);
nand U1162 (N_1162,N_468,N_46);
nor U1163 (N_1163,N_189,N_595);
and U1164 (N_1164,N_601,N_785);
or U1165 (N_1165,N_554,N_3);
and U1166 (N_1166,N_247,N_22);
nand U1167 (N_1167,N_611,N_43);
and U1168 (N_1168,N_85,N_183);
nor U1169 (N_1169,N_871,N_856);
and U1170 (N_1170,N_528,N_603);
nand U1171 (N_1171,N_41,N_542);
nor U1172 (N_1172,N_340,N_42);
nand U1173 (N_1173,N_591,N_374);
or U1174 (N_1174,N_796,N_753);
or U1175 (N_1175,N_277,N_459);
nor U1176 (N_1176,N_194,N_980);
and U1177 (N_1177,N_663,N_984);
or U1178 (N_1178,N_657,N_632);
nand U1179 (N_1179,N_977,N_337);
nand U1180 (N_1180,N_213,N_890);
nor U1181 (N_1181,N_136,N_253);
and U1182 (N_1182,N_312,N_144);
or U1183 (N_1183,N_134,N_687);
xnor U1184 (N_1184,N_240,N_417);
or U1185 (N_1185,N_887,N_470);
and U1186 (N_1186,N_93,N_574);
and U1187 (N_1187,N_225,N_66);
and U1188 (N_1188,N_38,N_59);
nor U1189 (N_1189,N_802,N_119);
nor U1190 (N_1190,N_723,N_445);
nand U1191 (N_1191,N_385,N_916);
nand U1192 (N_1192,N_809,N_897);
and U1193 (N_1193,N_940,N_561);
and U1194 (N_1194,N_73,N_742);
nand U1195 (N_1195,N_862,N_421);
nor U1196 (N_1196,N_557,N_65);
nor U1197 (N_1197,N_797,N_630);
nor U1198 (N_1198,N_806,N_949);
and U1199 (N_1199,N_743,N_892);
nor U1200 (N_1200,N_499,N_616);
and U1201 (N_1201,N_222,N_373);
and U1202 (N_1202,N_717,N_437);
nor U1203 (N_1203,N_316,N_578);
or U1204 (N_1204,N_372,N_67);
or U1205 (N_1205,N_162,N_24);
and U1206 (N_1206,N_825,N_974);
and U1207 (N_1207,N_257,N_11);
nor U1208 (N_1208,N_434,N_76);
nor U1209 (N_1209,N_2,N_822);
or U1210 (N_1210,N_885,N_791);
nand U1211 (N_1211,N_937,N_948);
nand U1212 (N_1212,N_771,N_288);
or U1213 (N_1213,N_903,N_120);
xor U1214 (N_1214,N_146,N_202);
and U1215 (N_1215,N_993,N_784);
nor U1216 (N_1216,N_699,N_508);
or U1217 (N_1217,N_536,N_677);
or U1218 (N_1218,N_731,N_81);
or U1219 (N_1219,N_206,N_981);
nor U1220 (N_1220,N_565,N_988);
and U1221 (N_1221,N_664,N_40);
and U1222 (N_1222,N_995,N_752);
nand U1223 (N_1223,N_217,N_703);
nand U1224 (N_1224,N_318,N_778);
nor U1225 (N_1225,N_493,N_650);
nor U1226 (N_1226,N_488,N_156);
nand U1227 (N_1227,N_945,N_726);
or U1228 (N_1228,N_946,N_972);
xnor U1229 (N_1229,N_939,N_409);
xnor U1230 (N_1230,N_830,N_320);
and U1231 (N_1231,N_549,N_516);
nand U1232 (N_1232,N_583,N_133);
or U1233 (N_1233,N_172,N_708);
nor U1234 (N_1234,N_363,N_992);
nand U1235 (N_1235,N_190,N_30);
or U1236 (N_1236,N_489,N_109);
and U1237 (N_1237,N_914,N_527);
nand U1238 (N_1238,N_506,N_607);
nor U1239 (N_1239,N_866,N_918);
xnor U1240 (N_1240,N_553,N_615);
nand U1241 (N_1241,N_919,N_262);
nand U1242 (N_1242,N_772,N_263);
nor U1243 (N_1243,N_425,N_501);
and U1244 (N_1244,N_333,N_145);
nor U1245 (N_1245,N_295,N_272);
and U1246 (N_1246,N_280,N_204);
or U1247 (N_1247,N_137,N_706);
and U1248 (N_1248,N_535,N_186);
and U1249 (N_1249,N_526,N_769);
or U1250 (N_1250,N_807,N_341);
nor U1251 (N_1251,N_127,N_804);
or U1252 (N_1252,N_786,N_870);
nand U1253 (N_1253,N_97,N_938);
and U1254 (N_1254,N_139,N_739);
nor U1255 (N_1255,N_449,N_198);
and U1256 (N_1256,N_439,N_28);
or U1257 (N_1257,N_646,N_864);
xor U1258 (N_1258,N_328,N_813);
nand U1259 (N_1259,N_234,N_123);
or U1260 (N_1260,N_349,N_429);
and U1261 (N_1261,N_712,N_795);
nand U1262 (N_1262,N_308,N_296);
nor U1263 (N_1263,N_560,N_814);
or U1264 (N_1264,N_313,N_375);
nand U1265 (N_1265,N_790,N_237);
or U1266 (N_1266,N_530,N_147);
nor U1267 (N_1267,N_199,N_336);
nand U1268 (N_1268,N_729,N_104);
nor U1269 (N_1269,N_460,N_928);
nor U1270 (N_1270,N_118,N_857);
and U1271 (N_1271,N_968,N_762);
and U1272 (N_1272,N_486,N_693);
or U1273 (N_1273,N_256,N_462);
nor U1274 (N_1274,N_143,N_185);
and U1275 (N_1275,N_546,N_405);
nand U1276 (N_1276,N_290,N_781);
nor U1277 (N_1277,N_404,N_287);
nor U1278 (N_1278,N_106,N_394);
nor U1279 (N_1279,N_641,N_511);
nor U1280 (N_1280,N_91,N_519);
and U1281 (N_1281,N_278,N_585);
nor U1282 (N_1282,N_850,N_570);
nor U1283 (N_1283,N_209,N_126);
and U1284 (N_1284,N_580,N_297);
and U1285 (N_1285,N_88,N_888);
or U1286 (N_1286,N_740,N_9);
and U1287 (N_1287,N_721,N_250);
nor U1288 (N_1288,N_205,N_430);
or U1289 (N_1289,N_231,N_266);
nor U1290 (N_1290,N_577,N_216);
and U1291 (N_1291,N_325,N_17);
and U1292 (N_1292,N_180,N_401);
nand U1293 (N_1293,N_403,N_858);
and U1294 (N_1294,N_999,N_377);
or U1295 (N_1295,N_883,N_569);
nor U1296 (N_1296,N_105,N_965);
nor U1297 (N_1297,N_329,N_924);
and U1298 (N_1298,N_285,N_321);
or U1299 (N_1299,N_495,N_113);
nand U1300 (N_1300,N_309,N_443);
nand U1301 (N_1301,N_812,N_675);
and U1302 (N_1302,N_943,N_579);
nor U1303 (N_1303,N_60,N_845);
or U1304 (N_1304,N_121,N_681);
and U1305 (N_1305,N_877,N_14);
and U1306 (N_1306,N_913,N_691);
xor U1307 (N_1307,N_852,N_889);
or U1308 (N_1308,N_952,N_602);
or U1309 (N_1309,N_875,N_62);
nand U1310 (N_1310,N_818,N_92);
and U1311 (N_1311,N_94,N_16);
nor U1312 (N_1312,N_408,N_192);
and U1313 (N_1313,N_33,N_164);
or U1314 (N_1314,N_884,N_0);
nand U1315 (N_1315,N_750,N_555);
nor U1316 (N_1316,N_274,N_550);
nand U1317 (N_1317,N_314,N_496);
nand U1318 (N_1318,N_638,N_860);
or U1319 (N_1319,N_457,N_135);
nor U1320 (N_1320,N_347,N_440);
or U1321 (N_1321,N_220,N_978);
nand U1322 (N_1322,N_358,N_279);
nand U1323 (N_1323,N_982,N_678);
nand U1324 (N_1324,N_976,N_393);
nand U1325 (N_1325,N_381,N_338);
or U1326 (N_1326,N_837,N_757);
nand U1327 (N_1327,N_529,N_129);
nand U1328 (N_1328,N_941,N_805);
or U1329 (N_1329,N_265,N_773);
and U1330 (N_1330,N_654,N_543);
xor U1331 (N_1331,N_444,N_702);
nor U1332 (N_1332,N_442,N_715);
or U1333 (N_1333,N_853,N_741);
or U1334 (N_1334,N_682,N_141);
nand U1335 (N_1335,N_958,N_788);
or U1336 (N_1336,N_386,N_365);
nand U1337 (N_1337,N_652,N_716);
and U1338 (N_1338,N_166,N_647);
or U1339 (N_1339,N_258,N_912);
nand U1340 (N_1340,N_175,N_75);
nor U1341 (N_1341,N_502,N_874);
or U1342 (N_1342,N_898,N_633);
nand U1343 (N_1343,N_453,N_879);
and U1344 (N_1344,N_930,N_639);
or U1345 (N_1345,N_910,N_467);
and U1346 (N_1346,N_933,N_426);
nand U1347 (N_1347,N_304,N_315);
nor U1348 (N_1348,N_651,N_7);
nand U1349 (N_1349,N_847,N_171);
xor U1350 (N_1350,N_665,N_317);
or U1351 (N_1351,N_298,N_492);
or U1352 (N_1352,N_484,N_597);
nand U1353 (N_1353,N_480,N_667);
nor U1354 (N_1354,N_955,N_400);
and U1355 (N_1355,N_259,N_74);
xor U1356 (N_1356,N_967,N_210);
and U1357 (N_1357,N_12,N_450);
and U1358 (N_1358,N_799,N_500);
nor U1359 (N_1359,N_44,N_84);
nor U1360 (N_1360,N_517,N_271);
nand U1361 (N_1361,N_148,N_840);
nor U1362 (N_1362,N_660,N_929);
or U1363 (N_1363,N_662,N_626);
and U1364 (N_1364,N_688,N_964);
or U1365 (N_1365,N_551,N_286);
and U1366 (N_1366,N_782,N_823);
nor U1367 (N_1367,N_334,N_923);
nor U1368 (N_1368,N_803,N_335);
nor U1369 (N_1369,N_1,N_704);
and U1370 (N_1370,N_268,N_556);
nor U1371 (N_1371,N_894,N_419);
nand U1372 (N_1372,N_154,N_636);
or U1373 (N_1373,N_71,N_881);
nor U1374 (N_1374,N_307,N_110);
or U1375 (N_1375,N_759,N_236);
xnor U1376 (N_1376,N_831,N_427);
nand U1377 (N_1377,N_219,N_177);
or U1378 (N_1378,N_342,N_841);
xnor U1379 (N_1379,N_451,N_122);
nand U1380 (N_1380,N_391,N_994);
and U1381 (N_1381,N_714,N_566);
nor U1382 (N_1382,N_925,N_547);
nand U1383 (N_1383,N_522,N_281);
and U1384 (N_1384,N_899,N_264);
or U1385 (N_1385,N_713,N_709);
nand U1386 (N_1386,N_132,N_414);
nand U1387 (N_1387,N_407,N_452);
and U1388 (N_1388,N_261,N_798);
nor U1389 (N_1389,N_537,N_676);
nor U1390 (N_1390,N_130,N_36);
nand U1391 (N_1391,N_520,N_35);
nand U1392 (N_1392,N_270,N_695);
and U1393 (N_1393,N_620,N_801);
and U1394 (N_1394,N_432,N_935);
nand U1395 (N_1395,N_50,N_833);
nor U1396 (N_1396,N_6,N_380);
and U1397 (N_1397,N_756,N_371);
nor U1398 (N_1398,N_810,N_820);
nor U1399 (N_1399,N_397,N_284);
and U1400 (N_1400,N_131,N_671);
or U1401 (N_1401,N_378,N_904);
nor U1402 (N_1402,N_211,N_152);
and U1403 (N_1403,N_661,N_792);
nor U1404 (N_1404,N_448,N_911);
nor U1405 (N_1405,N_327,N_973);
nand U1406 (N_1406,N_223,N_839);
or U1407 (N_1407,N_168,N_128);
and U1408 (N_1408,N_876,N_26);
or U1409 (N_1409,N_745,N_454);
or U1410 (N_1410,N_991,N_229);
and U1411 (N_1411,N_895,N_732);
or U1412 (N_1412,N_461,N_619);
and U1413 (N_1413,N_323,N_498);
nor U1414 (N_1414,N_214,N_544);
nor U1415 (N_1415,N_173,N_558);
nor U1416 (N_1416,N_181,N_228);
or U1417 (N_1417,N_564,N_548);
nor U1418 (N_1418,N_624,N_221);
nor U1419 (N_1419,N_158,N_983);
and U1420 (N_1420,N_252,N_423);
nand U1421 (N_1421,N_609,N_464);
nor U1422 (N_1422,N_867,N_844);
nand U1423 (N_1423,N_326,N_859);
and U1424 (N_1424,N_766,N_275);
nand U1425 (N_1425,N_422,N_370);
or U1426 (N_1426,N_182,N_8);
nand U1427 (N_1427,N_515,N_477);
and U1428 (N_1428,N_420,N_891);
nand U1429 (N_1429,N_996,N_357);
nor U1430 (N_1430,N_843,N_720);
or U1431 (N_1431,N_245,N_89);
nor U1432 (N_1432,N_737,N_761);
nor U1433 (N_1433,N_686,N_755);
xor U1434 (N_1434,N_125,N_157);
and U1435 (N_1435,N_300,N_292);
xor U1436 (N_1436,N_310,N_592);
and U1437 (N_1437,N_306,N_392);
nor U1438 (N_1438,N_525,N_160);
nand U1439 (N_1439,N_674,N_932);
or U1440 (N_1440,N_412,N_794);
or U1441 (N_1441,N_637,N_98);
xor U1442 (N_1442,N_353,N_571);
nor U1443 (N_1443,N_956,N_719);
nand U1444 (N_1444,N_303,N_931);
or U1445 (N_1445,N_99,N_824);
nor U1446 (N_1446,N_311,N_176);
nand U1447 (N_1447,N_474,N_230);
or U1448 (N_1448,N_107,N_504);
nand U1449 (N_1449,N_593,N_330);
or U1450 (N_1450,N_428,N_907);
or U1451 (N_1451,N_161,N_817);
nand U1452 (N_1452,N_915,N_779);
nand U1453 (N_1453,N_49,N_458);
nor U1454 (N_1454,N_698,N_54);
nor U1455 (N_1455,N_658,N_469);
nand U1456 (N_1456,N_58,N_224);
or U1457 (N_1457,N_848,N_643);
nand U1458 (N_1458,N_819,N_362);
and U1459 (N_1459,N_942,N_82);
nor U1460 (N_1460,N_670,N_149);
nor U1461 (N_1461,N_112,N_273);
nor U1462 (N_1462,N_388,N_299);
and U1463 (N_1463,N_893,N_961);
nor U1464 (N_1464,N_465,N_53);
nand U1465 (N_1465,N_195,N_835);
nor U1466 (N_1466,N_433,N_481);
and U1467 (N_1467,N_590,N_909);
nand U1468 (N_1468,N_503,N_672);
nor U1469 (N_1469,N_764,N_163);
nor U1470 (N_1470,N_69,N_491);
nor U1471 (N_1471,N_254,N_343);
or U1472 (N_1472,N_878,N_734);
nand U1473 (N_1473,N_441,N_815);
nand U1474 (N_1474,N_811,N_997);
and U1475 (N_1475,N_55,N_64);
or U1476 (N_1476,N_936,N_728);
nand U1477 (N_1477,N_70,N_922);
or U1478 (N_1478,N_83,N_649);
nor U1479 (N_1479,N_165,N_987);
or U1480 (N_1480,N_232,N_169);
or U1481 (N_1481,N_920,N_787);
or U1482 (N_1482,N_960,N_384);
or U1483 (N_1483,N_96,N_621);
or U1484 (N_1484,N_846,N_827);
nand U1485 (N_1485,N_87,N_659);
xnor U1486 (N_1486,N_436,N_733);
nand U1487 (N_1487,N_855,N_612);
nor U1488 (N_1488,N_763,N_86);
and U1489 (N_1489,N_218,N_767);
and U1490 (N_1490,N_482,N_985);
or U1491 (N_1491,N_975,N_963);
or U1492 (N_1492,N_836,N_692);
nand U1493 (N_1493,N_710,N_800);
and U1494 (N_1494,N_645,N_926);
nand U1495 (N_1495,N_115,N_435);
or U1496 (N_1496,N_567,N_101);
nand U1497 (N_1497,N_605,N_446);
nor U1498 (N_1498,N_345,N_832);
and U1499 (N_1499,N_455,N_599);
xnor U1500 (N_1500,N_723,N_86);
nor U1501 (N_1501,N_106,N_30);
xnor U1502 (N_1502,N_455,N_731);
or U1503 (N_1503,N_986,N_477);
nand U1504 (N_1504,N_998,N_159);
or U1505 (N_1505,N_573,N_255);
nand U1506 (N_1506,N_306,N_633);
xnor U1507 (N_1507,N_590,N_289);
or U1508 (N_1508,N_556,N_410);
nor U1509 (N_1509,N_126,N_362);
and U1510 (N_1510,N_393,N_52);
nor U1511 (N_1511,N_32,N_490);
nor U1512 (N_1512,N_870,N_662);
and U1513 (N_1513,N_825,N_306);
and U1514 (N_1514,N_620,N_784);
nor U1515 (N_1515,N_387,N_601);
nand U1516 (N_1516,N_547,N_182);
and U1517 (N_1517,N_45,N_207);
nor U1518 (N_1518,N_861,N_284);
and U1519 (N_1519,N_854,N_237);
or U1520 (N_1520,N_169,N_929);
nor U1521 (N_1521,N_315,N_697);
and U1522 (N_1522,N_954,N_111);
nand U1523 (N_1523,N_680,N_536);
nand U1524 (N_1524,N_927,N_315);
and U1525 (N_1525,N_807,N_384);
and U1526 (N_1526,N_678,N_800);
or U1527 (N_1527,N_242,N_744);
nand U1528 (N_1528,N_127,N_343);
or U1529 (N_1529,N_326,N_466);
or U1530 (N_1530,N_265,N_672);
or U1531 (N_1531,N_105,N_348);
or U1532 (N_1532,N_197,N_918);
nor U1533 (N_1533,N_0,N_398);
nor U1534 (N_1534,N_860,N_351);
and U1535 (N_1535,N_849,N_181);
and U1536 (N_1536,N_269,N_501);
nand U1537 (N_1537,N_232,N_762);
nor U1538 (N_1538,N_209,N_998);
nor U1539 (N_1539,N_204,N_292);
nor U1540 (N_1540,N_16,N_917);
nand U1541 (N_1541,N_760,N_898);
xor U1542 (N_1542,N_167,N_149);
nand U1543 (N_1543,N_595,N_281);
nor U1544 (N_1544,N_31,N_128);
or U1545 (N_1545,N_497,N_302);
nand U1546 (N_1546,N_750,N_393);
nor U1547 (N_1547,N_897,N_996);
or U1548 (N_1548,N_743,N_827);
nand U1549 (N_1549,N_287,N_785);
and U1550 (N_1550,N_12,N_457);
nor U1551 (N_1551,N_13,N_779);
or U1552 (N_1552,N_313,N_226);
nand U1553 (N_1553,N_261,N_61);
nor U1554 (N_1554,N_810,N_382);
or U1555 (N_1555,N_579,N_803);
nand U1556 (N_1556,N_98,N_552);
nor U1557 (N_1557,N_547,N_331);
nor U1558 (N_1558,N_912,N_866);
nand U1559 (N_1559,N_557,N_830);
nand U1560 (N_1560,N_195,N_752);
nand U1561 (N_1561,N_845,N_522);
or U1562 (N_1562,N_462,N_630);
or U1563 (N_1563,N_132,N_456);
nand U1564 (N_1564,N_329,N_936);
nor U1565 (N_1565,N_597,N_929);
or U1566 (N_1566,N_969,N_425);
nand U1567 (N_1567,N_623,N_854);
and U1568 (N_1568,N_700,N_476);
nor U1569 (N_1569,N_524,N_170);
or U1570 (N_1570,N_311,N_897);
nand U1571 (N_1571,N_154,N_707);
and U1572 (N_1572,N_284,N_569);
nor U1573 (N_1573,N_284,N_64);
nand U1574 (N_1574,N_718,N_347);
xor U1575 (N_1575,N_122,N_112);
nor U1576 (N_1576,N_162,N_877);
or U1577 (N_1577,N_381,N_628);
and U1578 (N_1578,N_214,N_95);
or U1579 (N_1579,N_396,N_618);
nor U1580 (N_1580,N_850,N_772);
and U1581 (N_1581,N_180,N_20);
nor U1582 (N_1582,N_283,N_112);
or U1583 (N_1583,N_132,N_794);
or U1584 (N_1584,N_829,N_858);
nand U1585 (N_1585,N_577,N_549);
or U1586 (N_1586,N_703,N_653);
nand U1587 (N_1587,N_292,N_537);
nor U1588 (N_1588,N_629,N_648);
or U1589 (N_1589,N_60,N_391);
nand U1590 (N_1590,N_906,N_634);
nor U1591 (N_1591,N_611,N_989);
nor U1592 (N_1592,N_219,N_53);
and U1593 (N_1593,N_709,N_200);
and U1594 (N_1594,N_964,N_237);
nor U1595 (N_1595,N_327,N_87);
or U1596 (N_1596,N_625,N_886);
or U1597 (N_1597,N_621,N_757);
or U1598 (N_1598,N_489,N_425);
or U1599 (N_1599,N_809,N_330);
or U1600 (N_1600,N_55,N_257);
or U1601 (N_1601,N_893,N_782);
and U1602 (N_1602,N_280,N_312);
nand U1603 (N_1603,N_347,N_138);
nand U1604 (N_1604,N_432,N_650);
or U1605 (N_1605,N_35,N_498);
nor U1606 (N_1606,N_402,N_231);
nor U1607 (N_1607,N_360,N_267);
nor U1608 (N_1608,N_317,N_425);
nor U1609 (N_1609,N_381,N_907);
nand U1610 (N_1610,N_323,N_952);
or U1611 (N_1611,N_20,N_571);
or U1612 (N_1612,N_192,N_786);
nor U1613 (N_1613,N_808,N_307);
and U1614 (N_1614,N_4,N_244);
nor U1615 (N_1615,N_614,N_223);
nor U1616 (N_1616,N_848,N_739);
nand U1617 (N_1617,N_763,N_741);
nor U1618 (N_1618,N_842,N_83);
and U1619 (N_1619,N_432,N_325);
nand U1620 (N_1620,N_141,N_85);
and U1621 (N_1621,N_657,N_448);
and U1622 (N_1622,N_574,N_287);
or U1623 (N_1623,N_675,N_35);
or U1624 (N_1624,N_243,N_830);
nand U1625 (N_1625,N_52,N_197);
and U1626 (N_1626,N_648,N_504);
and U1627 (N_1627,N_209,N_843);
or U1628 (N_1628,N_367,N_462);
or U1629 (N_1629,N_176,N_31);
and U1630 (N_1630,N_299,N_356);
or U1631 (N_1631,N_956,N_637);
nor U1632 (N_1632,N_906,N_807);
or U1633 (N_1633,N_542,N_175);
xnor U1634 (N_1634,N_870,N_242);
nor U1635 (N_1635,N_138,N_799);
or U1636 (N_1636,N_460,N_911);
and U1637 (N_1637,N_605,N_828);
nor U1638 (N_1638,N_468,N_619);
or U1639 (N_1639,N_536,N_678);
or U1640 (N_1640,N_662,N_544);
nor U1641 (N_1641,N_68,N_849);
and U1642 (N_1642,N_33,N_385);
or U1643 (N_1643,N_522,N_590);
or U1644 (N_1644,N_530,N_25);
or U1645 (N_1645,N_0,N_144);
and U1646 (N_1646,N_929,N_655);
nand U1647 (N_1647,N_999,N_455);
nor U1648 (N_1648,N_513,N_915);
or U1649 (N_1649,N_478,N_578);
or U1650 (N_1650,N_521,N_783);
nand U1651 (N_1651,N_523,N_707);
or U1652 (N_1652,N_850,N_530);
or U1653 (N_1653,N_841,N_239);
nand U1654 (N_1654,N_925,N_785);
nor U1655 (N_1655,N_733,N_970);
nor U1656 (N_1656,N_489,N_856);
or U1657 (N_1657,N_157,N_365);
nor U1658 (N_1658,N_980,N_584);
nor U1659 (N_1659,N_76,N_598);
nand U1660 (N_1660,N_760,N_177);
xor U1661 (N_1661,N_316,N_174);
nand U1662 (N_1662,N_146,N_889);
nor U1663 (N_1663,N_386,N_779);
or U1664 (N_1664,N_169,N_178);
nand U1665 (N_1665,N_624,N_414);
xor U1666 (N_1666,N_17,N_320);
or U1667 (N_1667,N_203,N_917);
and U1668 (N_1668,N_313,N_234);
and U1669 (N_1669,N_48,N_901);
and U1670 (N_1670,N_20,N_782);
or U1671 (N_1671,N_325,N_981);
nand U1672 (N_1672,N_195,N_873);
or U1673 (N_1673,N_9,N_701);
and U1674 (N_1674,N_584,N_73);
xor U1675 (N_1675,N_41,N_5);
nand U1676 (N_1676,N_208,N_649);
nand U1677 (N_1677,N_457,N_171);
xnor U1678 (N_1678,N_43,N_193);
or U1679 (N_1679,N_160,N_953);
nand U1680 (N_1680,N_712,N_744);
and U1681 (N_1681,N_30,N_81);
and U1682 (N_1682,N_847,N_313);
or U1683 (N_1683,N_462,N_135);
and U1684 (N_1684,N_712,N_214);
or U1685 (N_1685,N_543,N_727);
nor U1686 (N_1686,N_270,N_775);
and U1687 (N_1687,N_867,N_557);
or U1688 (N_1688,N_472,N_806);
or U1689 (N_1689,N_357,N_943);
nand U1690 (N_1690,N_657,N_112);
nand U1691 (N_1691,N_874,N_685);
or U1692 (N_1692,N_140,N_602);
and U1693 (N_1693,N_657,N_191);
or U1694 (N_1694,N_736,N_778);
or U1695 (N_1695,N_858,N_32);
or U1696 (N_1696,N_920,N_935);
xor U1697 (N_1697,N_715,N_573);
nor U1698 (N_1698,N_158,N_751);
nor U1699 (N_1699,N_4,N_827);
nor U1700 (N_1700,N_774,N_351);
nand U1701 (N_1701,N_130,N_411);
nand U1702 (N_1702,N_957,N_95);
or U1703 (N_1703,N_361,N_114);
nor U1704 (N_1704,N_710,N_659);
and U1705 (N_1705,N_531,N_622);
and U1706 (N_1706,N_482,N_672);
nand U1707 (N_1707,N_650,N_565);
nand U1708 (N_1708,N_419,N_238);
and U1709 (N_1709,N_120,N_294);
or U1710 (N_1710,N_191,N_764);
nor U1711 (N_1711,N_907,N_175);
nand U1712 (N_1712,N_564,N_270);
and U1713 (N_1713,N_54,N_953);
and U1714 (N_1714,N_133,N_387);
nand U1715 (N_1715,N_802,N_128);
nor U1716 (N_1716,N_289,N_929);
nand U1717 (N_1717,N_994,N_534);
and U1718 (N_1718,N_502,N_376);
or U1719 (N_1719,N_617,N_603);
nor U1720 (N_1720,N_786,N_776);
nand U1721 (N_1721,N_605,N_994);
nor U1722 (N_1722,N_206,N_309);
nand U1723 (N_1723,N_650,N_879);
and U1724 (N_1724,N_766,N_287);
xnor U1725 (N_1725,N_628,N_647);
and U1726 (N_1726,N_401,N_136);
and U1727 (N_1727,N_853,N_950);
and U1728 (N_1728,N_783,N_535);
and U1729 (N_1729,N_55,N_119);
nor U1730 (N_1730,N_691,N_94);
or U1731 (N_1731,N_475,N_625);
nand U1732 (N_1732,N_569,N_958);
nor U1733 (N_1733,N_337,N_290);
or U1734 (N_1734,N_923,N_592);
nor U1735 (N_1735,N_56,N_684);
and U1736 (N_1736,N_172,N_159);
nand U1737 (N_1737,N_908,N_61);
nand U1738 (N_1738,N_338,N_745);
nand U1739 (N_1739,N_425,N_849);
and U1740 (N_1740,N_556,N_129);
or U1741 (N_1741,N_612,N_886);
nand U1742 (N_1742,N_263,N_539);
or U1743 (N_1743,N_173,N_764);
nand U1744 (N_1744,N_248,N_200);
or U1745 (N_1745,N_639,N_141);
and U1746 (N_1746,N_45,N_488);
nor U1747 (N_1747,N_671,N_273);
and U1748 (N_1748,N_608,N_496);
nor U1749 (N_1749,N_747,N_228);
and U1750 (N_1750,N_594,N_499);
and U1751 (N_1751,N_860,N_625);
or U1752 (N_1752,N_812,N_311);
nor U1753 (N_1753,N_456,N_537);
or U1754 (N_1754,N_707,N_6);
or U1755 (N_1755,N_309,N_537);
and U1756 (N_1756,N_476,N_851);
and U1757 (N_1757,N_632,N_818);
nor U1758 (N_1758,N_620,N_483);
nor U1759 (N_1759,N_246,N_176);
nand U1760 (N_1760,N_618,N_188);
nand U1761 (N_1761,N_318,N_352);
xnor U1762 (N_1762,N_890,N_867);
or U1763 (N_1763,N_201,N_612);
nand U1764 (N_1764,N_715,N_355);
or U1765 (N_1765,N_615,N_822);
nor U1766 (N_1766,N_796,N_85);
and U1767 (N_1767,N_645,N_15);
nor U1768 (N_1768,N_845,N_984);
nor U1769 (N_1769,N_920,N_899);
nand U1770 (N_1770,N_198,N_784);
nor U1771 (N_1771,N_892,N_151);
or U1772 (N_1772,N_139,N_250);
xnor U1773 (N_1773,N_54,N_228);
nor U1774 (N_1774,N_185,N_306);
or U1775 (N_1775,N_176,N_679);
or U1776 (N_1776,N_233,N_427);
nor U1777 (N_1777,N_315,N_205);
and U1778 (N_1778,N_34,N_948);
nor U1779 (N_1779,N_411,N_910);
and U1780 (N_1780,N_778,N_267);
nor U1781 (N_1781,N_110,N_977);
nand U1782 (N_1782,N_208,N_853);
nor U1783 (N_1783,N_632,N_426);
nor U1784 (N_1784,N_47,N_616);
or U1785 (N_1785,N_349,N_174);
nand U1786 (N_1786,N_853,N_8);
nand U1787 (N_1787,N_67,N_195);
nor U1788 (N_1788,N_53,N_213);
and U1789 (N_1789,N_596,N_898);
nand U1790 (N_1790,N_472,N_765);
nand U1791 (N_1791,N_485,N_957);
nor U1792 (N_1792,N_655,N_750);
and U1793 (N_1793,N_333,N_51);
nor U1794 (N_1794,N_423,N_333);
nand U1795 (N_1795,N_347,N_592);
and U1796 (N_1796,N_91,N_195);
nand U1797 (N_1797,N_873,N_59);
nor U1798 (N_1798,N_295,N_94);
nand U1799 (N_1799,N_803,N_190);
nor U1800 (N_1800,N_992,N_458);
nor U1801 (N_1801,N_598,N_316);
or U1802 (N_1802,N_907,N_946);
and U1803 (N_1803,N_278,N_299);
nand U1804 (N_1804,N_586,N_732);
and U1805 (N_1805,N_905,N_147);
and U1806 (N_1806,N_310,N_766);
nor U1807 (N_1807,N_388,N_458);
nand U1808 (N_1808,N_467,N_897);
or U1809 (N_1809,N_331,N_445);
or U1810 (N_1810,N_106,N_607);
nor U1811 (N_1811,N_255,N_835);
nand U1812 (N_1812,N_293,N_107);
nor U1813 (N_1813,N_553,N_960);
nand U1814 (N_1814,N_475,N_864);
and U1815 (N_1815,N_828,N_604);
or U1816 (N_1816,N_630,N_452);
nand U1817 (N_1817,N_689,N_659);
or U1818 (N_1818,N_195,N_956);
or U1819 (N_1819,N_636,N_936);
or U1820 (N_1820,N_583,N_24);
or U1821 (N_1821,N_278,N_608);
nor U1822 (N_1822,N_387,N_389);
or U1823 (N_1823,N_875,N_928);
xnor U1824 (N_1824,N_659,N_735);
nor U1825 (N_1825,N_444,N_862);
nand U1826 (N_1826,N_467,N_17);
xnor U1827 (N_1827,N_29,N_908);
nor U1828 (N_1828,N_496,N_315);
nor U1829 (N_1829,N_135,N_756);
nor U1830 (N_1830,N_194,N_563);
nor U1831 (N_1831,N_926,N_670);
and U1832 (N_1832,N_749,N_244);
nor U1833 (N_1833,N_626,N_996);
nor U1834 (N_1834,N_232,N_968);
nand U1835 (N_1835,N_129,N_439);
and U1836 (N_1836,N_539,N_315);
nor U1837 (N_1837,N_549,N_183);
nand U1838 (N_1838,N_136,N_180);
nor U1839 (N_1839,N_826,N_844);
nor U1840 (N_1840,N_752,N_653);
nand U1841 (N_1841,N_861,N_519);
and U1842 (N_1842,N_876,N_614);
or U1843 (N_1843,N_965,N_738);
nor U1844 (N_1844,N_517,N_11);
nor U1845 (N_1845,N_380,N_294);
nand U1846 (N_1846,N_137,N_432);
nand U1847 (N_1847,N_507,N_301);
nor U1848 (N_1848,N_293,N_976);
nor U1849 (N_1849,N_780,N_827);
nor U1850 (N_1850,N_489,N_528);
nand U1851 (N_1851,N_305,N_975);
and U1852 (N_1852,N_932,N_870);
nand U1853 (N_1853,N_465,N_549);
or U1854 (N_1854,N_706,N_757);
nor U1855 (N_1855,N_348,N_174);
and U1856 (N_1856,N_384,N_451);
xor U1857 (N_1857,N_891,N_699);
nor U1858 (N_1858,N_46,N_162);
nor U1859 (N_1859,N_505,N_844);
nor U1860 (N_1860,N_287,N_225);
nor U1861 (N_1861,N_131,N_650);
or U1862 (N_1862,N_43,N_246);
or U1863 (N_1863,N_676,N_526);
nor U1864 (N_1864,N_53,N_941);
xor U1865 (N_1865,N_433,N_516);
and U1866 (N_1866,N_747,N_687);
and U1867 (N_1867,N_311,N_700);
nor U1868 (N_1868,N_683,N_875);
or U1869 (N_1869,N_382,N_206);
nand U1870 (N_1870,N_800,N_62);
nor U1871 (N_1871,N_19,N_609);
and U1872 (N_1872,N_36,N_423);
nor U1873 (N_1873,N_10,N_895);
nor U1874 (N_1874,N_678,N_825);
nor U1875 (N_1875,N_627,N_592);
nor U1876 (N_1876,N_578,N_100);
and U1877 (N_1877,N_377,N_492);
nand U1878 (N_1878,N_160,N_648);
and U1879 (N_1879,N_555,N_783);
nand U1880 (N_1880,N_516,N_550);
or U1881 (N_1881,N_532,N_989);
or U1882 (N_1882,N_318,N_962);
nand U1883 (N_1883,N_104,N_34);
nor U1884 (N_1884,N_216,N_637);
or U1885 (N_1885,N_586,N_403);
or U1886 (N_1886,N_570,N_522);
nor U1887 (N_1887,N_108,N_435);
nand U1888 (N_1888,N_226,N_156);
or U1889 (N_1889,N_271,N_192);
and U1890 (N_1890,N_600,N_813);
or U1891 (N_1891,N_996,N_669);
nor U1892 (N_1892,N_213,N_197);
and U1893 (N_1893,N_517,N_418);
and U1894 (N_1894,N_486,N_83);
nor U1895 (N_1895,N_386,N_815);
or U1896 (N_1896,N_316,N_929);
xnor U1897 (N_1897,N_362,N_31);
nand U1898 (N_1898,N_458,N_623);
or U1899 (N_1899,N_762,N_278);
nand U1900 (N_1900,N_305,N_270);
nor U1901 (N_1901,N_65,N_817);
nand U1902 (N_1902,N_235,N_641);
nor U1903 (N_1903,N_468,N_283);
nand U1904 (N_1904,N_271,N_783);
nand U1905 (N_1905,N_948,N_683);
and U1906 (N_1906,N_113,N_5);
and U1907 (N_1907,N_926,N_174);
or U1908 (N_1908,N_477,N_200);
nand U1909 (N_1909,N_871,N_130);
nand U1910 (N_1910,N_137,N_978);
and U1911 (N_1911,N_669,N_810);
nor U1912 (N_1912,N_365,N_687);
or U1913 (N_1913,N_24,N_882);
nand U1914 (N_1914,N_919,N_980);
nor U1915 (N_1915,N_456,N_608);
nor U1916 (N_1916,N_573,N_350);
nand U1917 (N_1917,N_393,N_617);
nor U1918 (N_1918,N_448,N_41);
or U1919 (N_1919,N_28,N_587);
nand U1920 (N_1920,N_872,N_615);
or U1921 (N_1921,N_913,N_195);
xnor U1922 (N_1922,N_631,N_116);
nand U1923 (N_1923,N_128,N_736);
nor U1924 (N_1924,N_9,N_856);
and U1925 (N_1925,N_697,N_43);
nand U1926 (N_1926,N_519,N_969);
or U1927 (N_1927,N_46,N_419);
nand U1928 (N_1928,N_528,N_693);
nand U1929 (N_1929,N_216,N_743);
nor U1930 (N_1930,N_586,N_448);
or U1931 (N_1931,N_383,N_400);
and U1932 (N_1932,N_235,N_916);
or U1933 (N_1933,N_852,N_109);
nor U1934 (N_1934,N_951,N_430);
nand U1935 (N_1935,N_317,N_396);
xnor U1936 (N_1936,N_703,N_132);
or U1937 (N_1937,N_96,N_411);
and U1938 (N_1938,N_80,N_727);
or U1939 (N_1939,N_853,N_190);
nor U1940 (N_1940,N_80,N_795);
and U1941 (N_1941,N_15,N_202);
or U1942 (N_1942,N_220,N_859);
and U1943 (N_1943,N_680,N_413);
or U1944 (N_1944,N_998,N_593);
or U1945 (N_1945,N_55,N_886);
nor U1946 (N_1946,N_188,N_291);
or U1947 (N_1947,N_879,N_608);
and U1948 (N_1948,N_225,N_88);
nand U1949 (N_1949,N_850,N_741);
nor U1950 (N_1950,N_237,N_6);
nand U1951 (N_1951,N_64,N_106);
xor U1952 (N_1952,N_659,N_993);
nor U1953 (N_1953,N_765,N_694);
nand U1954 (N_1954,N_157,N_100);
and U1955 (N_1955,N_548,N_953);
nor U1956 (N_1956,N_554,N_819);
nand U1957 (N_1957,N_114,N_86);
or U1958 (N_1958,N_980,N_734);
nand U1959 (N_1959,N_474,N_92);
or U1960 (N_1960,N_56,N_707);
and U1961 (N_1961,N_841,N_937);
nand U1962 (N_1962,N_401,N_559);
nor U1963 (N_1963,N_573,N_849);
nor U1964 (N_1964,N_845,N_99);
nor U1965 (N_1965,N_840,N_905);
nor U1966 (N_1966,N_534,N_540);
and U1967 (N_1967,N_959,N_23);
nand U1968 (N_1968,N_546,N_205);
nor U1969 (N_1969,N_119,N_931);
and U1970 (N_1970,N_658,N_935);
or U1971 (N_1971,N_693,N_272);
nor U1972 (N_1972,N_37,N_82);
xnor U1973 (N_1973,N_246,N_184);
nand U1974 (N_1974,N_796,N_229);
nand U1975 (N_1975,N_92,N_86);
nor U1976 (N_1976,N_353,N_550);
or U1977 (N_1977,N_260,N_141);
nor U1978 (N_1978,N_503,N_144);
or U1979 (N_1979,N_576,N_816);
or U1980 (N_1980,N_667,N_56);
nor U1981 (N_1981,N_421,N_604);
and U1982 (N_1982,N_149,N_298);
nor U1983 (N_1983,N_104,N_721);
nor U1984 (N_1984,N_175,N_566);
nand U1985 (N_1985,N_127,N_168);
nand U1986 (N_1986,N_343,N_730);
nand U1987 (N_1987,N_313,N_359);
and U1988 (N_1988,N_225,N_521);
or U1989 (N_1989,N_492,N_508);
nor U1990 (N_1990,N_271,N_460);
nand U1991 (N_1991,N_491,N_576);
or U1992 (N_1992,N_394,N_410);
nand U1993 (N_1993,N_863,N_39);
or U1994 (N_1994,N_604,N_152);
or U1995 (N_1995,N_993,N_46);
or U1996 (N_1996,N_982,N_381);
or U1997 (N_1997,N_945,N_569);
nor U1998 (N_1998,N_82,N_218);
nand U1999 (N_1999,N_878,N_516);
or U2000 (N_2000,N_1883,N_1189);
nor U2001 (N_2001,N_1692,N_1718);
and U2002 (N_2002,N_1657,N_1285);
or U2003 (N_2003,N_1422,N_1691);
nor U2004 (N_2004,N_1620,N_1311);
nand U2005 (N_2005,N_1017,N_1713);
nand U2006 (N_2006,N_1769,N_1605);
xor U2007 (N_2007,N_1645,N_1284);
or U2008 (N_2008,N_1612,N_1671);
xor U2009 (N_2009,N_1837,N_1503);
nor U2010 (N_2010,N_1524,N_1611);
nand U2011 (N_2011,N_1350,N_1370);
and U2012 (N_2012,N_1707,N_1548);
nor U2013 (N_2013,N_1720,N_1979);
nor U2014 (N_2014,N_1439,N_1549);
nor U2015 (N_2015,N_1468,N_1745);
nor U2016 (N_2016,N_1403,N_1555);
or U2017 (N_2017,N_1194,N_1289);
and U2018 (N_2018,N_1033,N_1537);
nand U2019 (N_2019,N_1283,N_1462);
nor U2020 (N_2020,N_1497,N_1102);
nor U2021 (N_2021,N_1067,N_1173);
and U2022 (N_2022,N_1743,N_1025);
nand U2023 (N_2023,N_1118,N_1268);
nor U2024 (N_2024,N_1434,N_1132);
nand U2025 (N_2025,N_1272,N_1911);
nand U2026 (N_2026,N_1469,N_1869);
nor U2027 (N_2027,N_1914,N_1801);
nor U2028 (N_2028,N_1894,N_1353);
nor U2029 (N_2029,N_1809,N_1633);
nor U2030 (N_2030,N_1738,N_1898);
nor U2031 (N_2031,N_1701,N_1001);
nand U2032 (N_2032,N_1091,N_1912);
xor U2033 (N_2033,N_1129,N_1617);
nor U2034 (N_2034,N_1952,N_1197);
nor U2035 (N_2035,N_1337,N_1995);
and U2036 (N_2036,N_1184,N_1502);
nand U2037 (N_2037,N_1448,N_1359);
or U2038 (N_2038,N_1774,N_1926);
xor U2039 (N_2039,N_1103,N_1310);
and U2040 (N_2040,N_1160,N_1742);
and U2041 (N_2041,N_1881,N_1843);
or U2042 (N_2042,N_1205,N_1977);
or U2043 (N_2043,N_1968,N_1538);
nor U2044 (N_2044,N_1217,N_1246);
and U2045 (N_2045,N_1980,N_1759);
or U2046 (N_2046,N_1652,N_1375);
or U2047 (N_2047,N_1624,N_1647);
or U2048 (N_2048,N_1013,N_1009);
nor U2049 (N_2049,N_1083,N_1142);
or U2050 (N_2050,N_1356,N_1232);
and U2051 (N_2051,N_1860,N_1642);
nor U2052 (N_2052,N_1279,N_1243);
nor U2053 (N_2053,N_1240,N_1037);
nor U2054 (N_2054,N_1585,N_1404);
and U2055 (N_2055,N_1423,N_1460);
nand U2056 (N_2056,N_1807,N_1248);
nor U2057 (N_2057,N_1724,N_1589);
or U2058 (N_2058,N_1999,N_1676);
or U2059 (N_2059,N_1047,N_1886);
and U2060 (N_2060,N_1494,N_1966);
and U2061 (N_2061,N_1821,N_1044);
or U2062 (N_2062,N_1454,N_1544);
and U2063 (N_2063,N_1314,N_1293);
and U2064 (N_2064,N_1580,N_1507);
or U2065 (N_2065,N_1426,N_1579);
nand U2066 (N_2066,N_1378,N_1270);
or U2067 (N_2067,N_1292,N_1955);
nand U2068 (N_2068,N_1074,N_1204);
and U2069 (N_2069,N_1573,N_1783);
and U2070 (N_2070,N_1053,N_1073);
or U2071 (N_2071,N_1148,N_1690);
and U2072 (N_2072,N_1405,N_1927);
xor U2073 (N_2073,N_1361,N_1334);
or U2074 (N_2074,N_1020,N_1233);
or U2075 (N_2075,N_1062,N_1574);
nor U2076 (N_2076,N_1785,N_1962);
or U2077 (N_2077,N_1365,N_1298);
nor U2078 (N_2078,N_1068,N_1790);
and U2079 (N_2079,N_1629,N_1986);
and U2080 (N_2080,N_1997,N_1249);
or U2081 (N_2081,N_1301,N_1722);
and U2082 (N_2082,N_1851,N_1302);
nand U2083 (N_2083,N_1297,N_1491);
nor U2084 (N_2084,N_1026,N_1152);
or U2085 (N_2085,N_1793,N_1918);
nand U2086 (N_2086,N_1971,N_1552);
or U2087 (N_2087,N_1873,N_1377);
and U2088 (N_2088,N_1147,N_1055);
nand U2089 (N_2089,N_1256,N_1296);
or U2090 (N_2090,N_1655,N_1907);
and U2091 (N_2091,N_1614,N_1588);
nand U2092 (N_2092,N_1784,N_1901);
and U2093 (N_2093,N_1364,N_1495);
nor U2094 (N_2094,N_1562,N_1402);
nand U2095 (N_2095,N_1482,N_1581);
nand U2096 (N_2096,N_1467,N_1957);
nor U2097 (N_2097,N_1667,N_1688);
nor U2098 (N_2098,N_1938,N_1014);
and U2099 (N_2099,N_1778,N_1648);
and U2100 (N_2100,N_1711,N_1450);
nor U2101 (N_2101,N_1835,N_1027);
nand U2102 (N_2102,N_1115,N_1127);
nand U2103 (N_2103,N_1369,N_1440);
and U2104 (N_2104,N_1678,N_1162);
nand U2105 (N_2105,N_1829,N_1700);
and U2106 (N_2106,N_1568,N_1034);
nand U2107 (N_2107,N_1521,N_1376);
or U2108 (N_2108,N_1695,N_1400);
or U2109 (N_2109,N_1312,N_1386);
or U2110 (N_2110,N_1139,N_1125);
nand U2111 (N_2111,N_1438,N_1739);
nand U2112 (N_2112,N_1193,N_1474);
and U2113 (N_2113,N_1882,N_1327);
or U2114 (N_2114,N_1429,N_1456);
nor U2115 (N_2115,N_1185,N_1346);
and U2116 (N_2116,N_1960,N_1109);
or U2117 (N_2117,N_1158,N_1308);
or U2118 (N_2118,N_1399,N_1550);
and U2119 (N_2119,N_1866,N_1824);
and U2120 (N_2120,N_1687,N_1650);
nand U2121 (N_2121,N_1668,N_1081);
nor U2122 (N_2122,N_1244,N_1061);
nand U2123 (N_2123,N_1355,N_1523);
or U2124 (N_2124,N_1983,N_1628);
nor U2125 (N_2125,N_1511,N_1090);
or U2126 (N_2126,N_1181,N_1577);
nand U2127 (N_2127,N_1373,N_1332);
nand U2128 (N_2128,N_1059,N_1318);
nand U2129 (N_2129,N_1638,N_1409);
nand U2130 (N_2130,N_1681,N_1984);
nand U2131 (N_2131,N_1566,N_1848);
nand U2132 (N_2132,N_1572,N_1519);
or U2133 (N_2133,N_1985,N_1763);
nor U2134 (N_2134,N_1374,N_1392);
nand U2135 (N_2135,N_1413,N_1196);
and U2136 (N_2136,N_1871,N_1209);
and U2137 (N_2137,N_1343,N_1388);
and U2138 (N_2138,N_1042,N_1922);
nand U2139 (N_2139,N_1828,N_1049);
nand U2140 (N_2140,N_1056,N_1563);
nor U2141 (N_2141,N_1818,N_1590);
or U2142 (N_2142,N_1751,N_1215);
or U2143 (N_2143,N_1557,N_1512);
nor U2144 (N_2144,N_1251,N_1300);
nand U2145 (N_2145,N_1282,N_1823);
or U2146 (N_2146,N_1206,N_1682);
or U2147 (N_2147,N_1876,N_1096);
nand U2148 (N_2148,N_1664,N_1561);
and U2149 (N_2149,N_1444,N_1547);
nor U2150 (N_2150,N_1211,N_1260);
or U2151 (N_2151,N_1570,N_1075);
and U2152 (N_2152,N_1459,N_1177);
and U2153 (N_2153,N_1263,N_1822);
nand U2154 (N_2154,N_1227,N_1637);
nor U2155 (N_2155,N_1223,N_1208);
nor U2156 (N_2156,N_1916,N_1202);
or U2157 (N_2157,N_1191,N_1554);
and U2158 (N_2158,N_1385,N_1508);
nand U2159 (N_2159,N_1281,N_1295);
or U2160 (N_2160,N_1693,N_1065);
nand U2161 (N_2161,N_1838,N_1273);
nand U2162 (N_2162,N_1335,N_1172);
nand U2163 (N_2163,N_1221,N_1461);
nor U2164 (N_2164,N_1551,N_1736);
xor U2165 (N_2165,N_1754,N_1305);
nor U2166 (N_2166,N_1731,N_1996);
and U2167 (N_2167,N_1245,N_1225);
or U2168 (N_2168,N_1266,N_1760);
or U2169 (N_2169,N_1775,N_1872);
nor U2170 (N_2170,N_1780,N_1321);
nand U2171 (N_2171,N_1900,N_1133);
and U2172 (N_2172,N_1286,N_1051);
and U2173 (N_2173,N_1174,N_1683);
nor U2174 (N_2174,N_1594,N_1452);
or U2175 (N_2175,N_1154,N_1203);
nand U2176 (N_2176,N_1060,N_1261);
nand U2177 (N_2177,N_1150,N_1728);
and U2178 (N_2178,N_1372,N_1704);
nor U2179 (N_2179,N_1137,N_1913);
or U2180 (N_2180,N_1600,N_1316);
nand U2181 (N_2181,N_1956,N_1744);
or U2182 (N_2182,N_1277,N_1239);
or U2183 (N_2183,N_1694,N_1564);
and U2184 (N_2184,N_1915,N_1702);
nor U2185 (N_2185,N_1903,N_1716);
or U2186 (N_2186,N_1290,N_1319);
nand U2187 (N_2187,N_1597,N_1367);
nor U2188 (N_2188,N_1254,N_1043);
or U2189 (N_2189,N_1924,N_1639);
nor U2190 (N_2190,N_1443,N_1510);
nand U2191 (N_2191,N_1826,N_1380);
or U2192 (N_2192,N_1234,N_1499);
nand U2193 (N_2193,N_1608,N_1868);
and U2194 (N_2194,N_1680,N_1477);
and U2195 (N_2195,N_1358,N_1861);
or U2196 (N_2196,N_1219,N_1362);
or U2197 (N_2197,N_1097,N_1411);
nor U2198 (N_2198,N_1333,N_1387);
or U2199 (N_2199,N_1635,N_1906);
nor U2200 (N_2200,N_1085,N_1967);
and U2201 (N_2201,N_1640,N_1057);
and U2202 (N_2202,N_1170,N_1231);
or U2203 (N_2203,N_1076,N_1427);
nor U2204 (N_2204,N_1974,N_1418);
nand U2205 (N_2205,N_1602,N_1220);
nor U2206 (N_2206,N_1982,N_1472);
nor U2207 (N_2207,N_1330,N_1630);
nor U2208 (N_2208,N_1788,N_1844);
and U2209 (N_2209,N_1727,N_1946);
and U2210 (N_2210,N_1099,N_1948);
and U2211 (N_2211,N_1803,N_1522);
and U2212 (N_2212,N_1253,N_1994);
nand U2213 (N_2213,N_1393,N_1379);
and U2214 (N_2214,N_1156,N_1007);
and U2215 (N_2215,N_1601,N_1464);
nor U2216 (N_2216,N_1978,N_1766);
or U2217 (N_2217,N_1309,N_1972);
and U2218 (N_2218,N_1752,N_1070);
nand U2219 (N_2219,N_1627,N_1490);
nand U2220 (N_2220,N_1041,N_1351);
nor U2221 (N_2221,N_1593,N_1271);
and U2222 (N_2222,N_1529,N_1420);
and U2223 (N_2223,N_1395,N_1965);
and U2224 (N_2224,N_1241,N_1679);
nor U2225 (N_2225,N_1038,N_1756);
nand U2226 (N_2226,N_1275,N_1484);
nor U2227 (N_2227,N_1578,N_1862);
or U2228 (N_2228,N_1749,N_1094);
and U2229 (N_2229,N_1762,N_1770);
nor U2230 (N_2230,N_1063,N_1035);
nor U2231 (N_2231,N_1110,N_1684);
nand U2232 (N_2232,N_1870,N_1735);
and U2233 (N_2233,N_1794,N_1709);
and U2234 (N_2234,N_1322,N_1294);
nand U2235 (N_2235,N_1659,N_1149);
nand U2236 (N_2236,N_1326,N_1931);
and U2237 (N_2237,N_1307,N_1222);
and U2238 (N_2238,N_1849,N_1665);
nor U2239 (N_2239,N_1004,N_1626);
xor U2240 (N_2240,N_1415,N_1888);
nand U2241 (N_2241,N_1610,N_1224);
or U2242 (N_2242,N_1981,N_1534);
or U2243 (N_2243,N_1576,N_1928);
xor U2244 (N_2244,N_1079,N_1772);
or U2245 (N_2245,N_1368,N_1252);
or U2246 (N_2246,N_1939,N_1964);
and U2247 (N_2247,N_1182,N_1940);
nand U2248 (N_2248,N_1942,N_1636);
nor U2249 (N_2249,N_1506,N_1816);
nor U2250 (N_2250,N_1814,N_1710);
nor U2251 (N_2251,N_1453,N_1853);
or U2252 (N_2252,N_1930,N_1800);
and U2253 (N_2253,N_1567,N_1480);
nand U2254 (N_2254,N_1781,N_1287);
and U2255 (N_2255,N_1539,N_1991);
nand U2256 (N_2256,N_1151,N_1012);
or U2257 (N_2257,N_1514,N_1541);
nor U2258 (N_2258,N_1155,N_1135);
or U2259 (N_2259,N_1228,N_1808);
nor U2260 (N_2260,N_1841,N_1317);
and U2261 (N_2261,N_1501,N_1168);
and U2262 (N_2262,N_1002,N_1804);
nor U2263 (N_2263,N_1712,N_1806);
or U2264 (N_2264,N_1777,N_1157);
or U2265 (N_2265,N_1666,N_1451);
or U2266 (N_2266,N_1825,N_1998);
and U2267 (N_2267,N_1389,N_1210);
or U2268 (N_2268,N_1836,N_1117);
nand U2269 (N_2269,N_1341,N_1264);
xnor U2270 (N_2270,N_1891,N_1737);
or U2271 (N_2271,N_1144,N_1131);
nor U2272 (N_2272,N_1487,N_1839);
and U2273 (N_2273,N_1779,N_1120);
nand U2274 (N_2274,N_1791,N_1315);
nand U2275 (N_2275,N_1757,N_1407);
or U2276 (N_2276,N_1530,N_1116);
nand U2277 (N_2277,N_1865,N_1328);
or U2278 (N_2278,N_1675,N_1893);
nor U2279 (N_2279,N_1925,N_1080);
and U2280 (N_2280,N_1758,N_1190);
nand U2281 (N_2281,N_1431,N_1164);
nor U2282 (N_2282,N_1280,N_1899);
nand U2283 (N_2283,N_1923,N_1255);
nand U2284 (N_2284,N_1787,N_1516);
or U2285 (N_2285,N_1492,N_1797);
or U2286 (N_2286,N_1463,N_1112);
or U2287 (N_2287,N_1662,N_1815);
and U2288 (N_2288,N_1045,N_1943);
nand U2289 (N_2289,N_1908,N_1618);
nor U2290 (N_2290,N_1006,N_1428);
or U2291 (N_2291,N_1599,N_1218);
nand U2292 (N_2292,N_1072,N_1140);
or U2293 (N_2293,N_1352,N_1746);
nor U2294 (N_2294,N_1706,N_1768);
or U2295 (N_2295,N_1344,N_1119);
and U2296 (N_2296,N_1107,N_1104);
and U2297 (N_2297,N_1944,N_1274);
nor U2298 (N_2298,N_1771,N_1340);
or U2299 (N_2299,N_1625,N_1734);
and U2300 (N_2300,N_1613,N_1799);
and U2301 (N_2301,N_1394,N_1767);
or U2302 (N_2302,N_1186,N_1969);
or U2303 (N_2303,N_1349,N_1656);
nand U2304 (N_2304,N_1481,N_1108);
and U2305 (N_2305,N_1864,N_1226);
nand U2306 (N_2306,N_1646,N_1748);
nor U2307 (N_2307,N_1859,N_1412);
and U2308 (N_2308,N_1488,N_1895);
or U2309 (N_2309,N_1747,N_1010);
nor U2310 (N_2310,N_1291,N_1050);
nor U2311 (N_2311,N_1817,N_1992);
nor U2312 (N_2312,N_1820,N_1171);
xnor U2313 (N_2313,N_1089,N_1698);
or U2314 (N_2314,N_1382,N_1179);
nand U2315 (N_2315,N_1932,N_1528);
nand U2316 (N_2316,N_1532,N_1575);
or U2317 (N_2317,N_1213,N_1854);
nor U2318 (N_2318,N_1313,N_1054);
and U2319 (N_2319,N_1634,N_1084);
nand U2320 (N_2320,N_1792,N_1988);
and U2321 (N_2321,N_1878,N_1471);
nor U2322 (N_2322,N_1212,N_1163);
and U2323 (N_2323,N_1904,N_1660);
or U2324 (N_2324,N_1465,N_1052);
and U2325 (N_2325,N_1850,N_1141);
nor U2326 (N_2326,N_1449,N_1011);
and U2327 (N_2327,N_1658,N_1505);
and U2328 (N_2328,N_1195,N_1805);
and U2329 (N_2329,N_1145,N_1029);
nand U2330 (N_2330,N_1338,N_1559);
nor U2331 (N_2331,N_1919,N_1008);
nand U2332 (N_2332,N_1390,N_1238);
nor U2333 (N_2333,N_1832,N_1410);
nor U2334 (N_2334,N_1531,N_1858);
and U2335 (N_2335,N_1653,N_1686);
or U2336 (N_2336,N_1398,N_1421);
nand U2337 (N_2337,N_1262,N_1733);
and U2338 (N_2338,N_1437,N_1381);
or U2339 (N_2339,N_1833,N_1875);
and U2340 (N_2340,N_1740,N_1885);
nand U2341 (N_2341,N_1436,N_1455);
or U2342 (N_2342,N_1533,N_1857);
or U2343 (N_2343,N_1348,N_1920);
nor U2344 (N_2344,N_1087,N_1371);
nand U2345 (N_2345,N_1265,N_1242);
or U2346 (N_2346,N_1959,N_1237);
nand U2347 (N_2347,N_1098,N_1458);
and U2348 (N_2348,N_1632,N_1216);
and U2349 (N_2349,N_1867,N_1100);
nor U2350 (N_2350,N_1546,N_1954);
and U2351 (N_2351,N_1542,N_1391);
nor U2352 (N_2352,N_1320,N_1603);
nor U2353 (N_2353,N_1031,N_1961);
nand U2354 (N_2354,N_1470,N_1199);
or U2355 (N_2355,N_1071,N_1136);
nor U2356 (N_2356,N_1124,N_1855);
nand U2357 (N_2357,N_1018,N_1200);
nand U2358 (N_2358,N_1121,N_1649);
nor U2359 (N_2359,N_1587,N_1419);
and U2360 (N_2360,N_1021,N_1432);
nor U2361 (N_2361,N_1786,N_1897);
nand U2362 (N_2362,N_1884,N_1130);
or U2363 (N_2363,N_1478,N_1619);
xor U2364 (N_2364,N_1933,N_1354);
nor U2365 (N_2365,N_1595,N_1408);
nand U2366 (N_2366,N_1235,N_1685);
nand U2367 (N_2367,N_1976,N_1299);
or U2368 (N_2368,N_1723,N_1750);
nor U2369 (N_2369,N_1761,N_1384);
xnor U2370 (N_2370,N_1526,N_1143);
and U2371 (N_2371,N_1661,N_1910);
nand U2372 (N_2372,N_1058,N_1414);
or U2373 (N_2373,N_1937,N_1621);
nor U2374 (N_2374,N_1066,N_1105);
and U2375 (N_2375,N_1159,N_1331);
and U2376 (N_2376,N_1834,N_1446);
nand U2377 (N_2377,N_1796,N_1257);
nand U2378 (N_2378,N_1306,N_1896);
nand U2379 (N_2379,N_1669,N_1069);
nor U2380 (N_2380,N_1479,N_1902);
or U2381 (N_2381,N_1674,N_1543);
nand U2382 (N_2382,N_1324,N_1250);
nor U2383 (N_2383,N_1880,N_1717);
and U2384 (N_2384,N_1565,N_1517);
or U2385 (N_2385,N_1134,N_1126);
nor U2386 (N_2386,N_1032,N_1417);
nor U2387 (N_2387,N_1934,N_1123);
nand U2388 (N_2388,N_1023,N_1167);
or U2389 (N_2389,N_1178,N_1879);
nor U2390 (N_2390,N_1106,N_1342);
nand U2391 (N_2391,N_1445,N_1236);
or U2392 (N_2392,N_1486,N_1622);
xnor U2393 (N_2393,N_1229,N_1852);
or U2394 (N_2394,N_1498,N_1259);
and U2395 (N_2395,N_1776,N_1989);
nor U2396 (N_2396,N_1697,N_1582);
or U2397 (N_2397,N_1874,N_1040);
nand U2398 (N_2398,N_1592,N_1963);
or U2399 (N_2399,N_1987,N_1782);
or U2400 (N_2400,N_1558,N_1303);
and U2401 (N_2401,N_1831,N_1586);
or U2402 (N_2402,N_1113,N_1651);
or U2403 (N_2403,N_1515,N_1146);
nand U2404 (N_2404,N_1863,N_1730);
or U2405 (N_2405,N_1773,N_1525);
or U2406 (N_2406,N_1088,N_1175);
and U2407 (N_2407,N_1201,N_1345);
nor U2408 (N_2408,N_1905,N_1489);
and U2409 (N_2409,N_1813,N_1092);
or U2410 (N_2410,N_1111,N_1721);
nor U2411 (N_2411,N_1935,N_1247);
or U2412 (N_2412,N_1949,N_1188);
nand U2413 (N_2413,N_1329,N_1323);
and U2414 (N_2414,N_1811,N_1500);
nand U2415 (N_2415,N_1689,N_1036);
nor U2416 (N_2416,N_1527,N_1483);
or U2417 (N_2417,N_1513,N_1670);
or U2418 (N_2418,N_1540,N_1015);
nor U2419 (N_2419,N_1114,N_1192);
nand U2420 (N_2420,N_1161,N_1267);
nor U2421 (N_2421,N_1936,N_1509);
nor U2422 (N_2422,N_1441,N_1401);
and U2423 (N_2423,N_1030,N_1973);
nor U2424 (N_2424,N_1048,N_1819);
nand U2425 (N_2425,N_1609,N_1416);
nor U2426 (N_2426,N_1641,N_1003);
nand U2427 (N_2427,N_1396,N_1466);
nor U2428 (N_2428,N_1269,N_1755);
or U2429 (N_2429,N_1654,N_1258);
and U2430 (N_2430,N_1536,N_1571);
nand U2431 (N_2431,N_1729,N_1475);
nand U2432 (N_2432,N_1000,N_1725);
nor U2433 (N_2433,N_1024,N_1556);
or U2434 (N_2434,N_1433,N_1699);
or U2435 (N_2435,N_1214,N_1278);
and U2436 (N_2436,N_1169,N_1122);
and U2437 (N_2437,N_1447,N_1086);
nand U2438 (N_2438,N_1128,N_1082);
nand U2439 (N_2439,N_1518,N_1046);
nand U2440 (N_2440,N_1892,N_1138);
nand U2441 (N_2441,N_1604,N_1719);
nand U2442 (N_2442,N_1795,N_1677);
nor U2443 (N_2443,N_1424,N_1696);
or U2444 (N_2444,N_1016,N_1802);
nand U2445 (N_2445,N_1715,N_1039);
nand U2446 (N_2446,N_1183,N_1741);
nor U2447 (N_2447,N_1606,N_1929);
nand U2448 (N_2448,N_1714,N_1703);
nor U2449 (N_2449,N_1553,N_1990);
and U2450 (N_2450,N_1945,N_1789);
or U2451 (N_2451,N_1975,N_1366);
or U2452 (N_2452,N_1847,N_1753);
nand U2453 (N_2453,N_1877,N_1764);
or U2454 (N_2454,N_1917,N_1705);
or U2455 (N_2455,N_1485,N_1643);
and U2456 (N_2456,N_1363,N_1947);
nor U2457 (N_2457,N_1383,N_1078);
nand U2458 (N_2458,N_1663,N_1856);
nor U2459 (N_2459,N_1187,N_1325);
nor U2460 (N_2460,N_1845,N_1028);
nand U2461 (N_2461,N_1623,N_1993);
nor U2462 (N_2462,N_1631,N_1535);
and U2463 (N_2463,N_1584,N_1176);
or U2464 (N_2464,N_1230,N_1909);
or U2465 (N_2465,N_1615,N_1276);
nor U2466 (N_2466,N_1504,N_1953);
nor U2467 (N_2467,N_1493,N_1810);
and U2468 (N_2468,N_1095,N_1798);
or U2469 (N_2469,N_1921,N_1591);
or U2470 (N_2470,N_1476,N_1198);
nor U2471 (N_2471,N_1569,N_1457);
nor U2472 (N_2472,N_1339,N_1890);
nand U2473 (N_2473,N_1732,N_1101);
and U2474 (N_2474,N_1425,N_1827);
nand U2475 (N_2475,N_1397,N_1166);
or U2476 (N_2476,N_1093,N_1598);
nand U2477 (N_2477,N_1889,N_1840);
nor U2478 (N_2478,N_1941,N_1673);
nand U2479 (N_2479,N_1644,N_1812);
nor U2480 (N_2480,N_1288,N_1022);
xnor U2481 (N_2481,N_1830,N_1545);
nand U2482 (N_2482,N_1951,N_1520);
or U2483 (N_2483,N_1406,N_1970);
and U2484 (N_2484,N_1207,N_1165);
and U2485 (N_2485,N_1596,N_1496);
and U2486 (N_2486,N_1950,N_1442);
or U2487 (N_2487,N_1153,N_1607);
nor U2488 (N_2488,N_1672,N_1430);
nor U2489 (N_2489,N_1347,N_1473);
and U2490 (N_2490,N_1765,N_1616);
and U2491 (N_2491,N_1726,N_1077);
nor U2492 (N_2492,N_1360,N_1304);
or U2493 (N_2493,N_1846,N_1064);
and U2494 (N_2494,N_1180,N_1336);
nand U2495 (N_2495,N_1435,N_1842);
xor U2496 (N_2496,N_1005,N_1357);
or U2497 (N_2497,N_1583,N_1019);
and U2498 (N_2498,N_1560,N_1958);
nand U2499 (N_2499,N_1887,N_1708);
or U2500 (N_2500,N_1205,N_1153);
nor U2501 (N_2501,N_1022,N_1998);
nor U2502 (N_2502,N_1141,N_1704);
or U2503 (N_2503,N_1610,N_1024);
nand U2504 (N_2504,N_1986,N_1030);
and U2505 (N_2505,N_1336,N_1956);
and U2506 (N_2506,N_1024,N_1793);
nor U2507 (N_2507,N_1134,N_1051);
nor U2508 (N_2508,N_1676,N_1608);
and U2509 (N_2509,N_1157,N_1227);
xnor U2510 (N_2510,N_1719,N_1073);
and U2511 (N_2511,N_1411,N_1165);
xnor U2512 (N_2512,N_1852,N_1452);
nor U2513 (N_2513,N_1512,N_1662);
or U2514 (N_2514,N_1135,N_1111);
nor U2515 (N_2515,N_1080,N_1405);
and U2516 (N_2516,N_1190,N_1750);
xor U2517 (N_2517,N_1940,N_1191);
and U2518 (N_2518,N_1827,N_1024);
nand U2519 (N_2519,N_1481,N_1199);
or U2520 (N_2520,N_1379,N_1079);
and U2521 (N_2521,N_1473,N_1130);
nand U2522 (N_2522,N_1679,N_1203);
nor U2523 (N_2523,N_1669,N_1698);
nor U2524 (N_2524,N_1488,N_1687);
and U2525 (N_2525,N_1587,N_1404);
nor U2526 (N_2526,N_1232,N_1224);
or U2527 (N_2527,N_1490,N_1870);
nand U2528 (N_2528,N_1579,N_1538);
or U2529 (N_2529,N_1547,N_1086);
nand U2530 (N_2530,N_1898,N_1605);
and U2531 (N_2531,N_1972,N_1809);
or U2532 (N_2532,N_1103,N_1987);
nor U2533 (N_2533,N_1622,N_1011);
or U2534 (N_2534,N_1446,N_1942);
nand U2535 (N_2535,N_1365,N_1375);
and U2536 (N_2536,N_1128,N_1631);
and U2537 (N_2537,N_1464,N_1157);
and U2538 (N_2538,N_1061,N_1310);
nand U2539 (N_2539,N_1846,N_1244);
nand U2540 (N_2540,N_1002,N_1661);
nand U2541 (N_2541,N_1154,N_1414);
and U2542 (N_2542,N_1812,N_1114);
and U2543 (N_2543,N_1858,N_1662);
or U2544 (N_2544,N_1938,N_1519);
nand U2545 (N_2545,N_1428,N_1912);
or U2546 (N_2546,N_1675,N_1338);
nor U2547 (N_2547,N_1298,N_1125);
or U2548 (N_2548,N_1375,N_1713);
nand U2549 (N_2549,N_1773,N_1541);
and U2550 (N_2550,N_1926,N_1133);
or U2551 (N_2551,N_1763,N_1468);
nand U2552 (N_2552,N_1405,N_1971);
and U2553 (N_2553,N_1314,N_1908);
nand U2554 (N_2554,N_1729,N_1693);
xor U2555 (N_2555,N_1919,N_1662);
nor U2556 (N_2556,N_1348,N_1604);
nand U2557 (N_2557,N_1986,N_1213);
nand U2558 (N_2558,N_1683,N_1237);
nor U2559 (N_2559,N_1732,N_1771);
or U2560 (N_2560,N_1386,N_1910);
nand U2561 (N_2561,N_1550,N_1987);
or U2562 (N_2562,N_1403,N_1050);
nor U2563 (N_2563,N_1556,N_1052);
or U2564 (N_2564,N_1451,N_1473);
or U2565 (N_2565,N_1612,N_1942);
nand U2566 (N_2566,N_1146,N_1640);
nor U2567 (N_2567,N_1454,N_1431);
or U2568 (N_2568,N_1098,N_1414);
nor U2569 (N_2569,N_1774,N_1581);
and U2570 (N_2570,N_1593,N_1858);
nor U2571 (N_2571,N_1086,N_1554);
or U2572 (N_2572,N_1039,N_1755);
and U2573 (N_2573,N_1052,N_1639);
and U2574 (N_2574,N_1178,N_1414);
nor U2575 (N_2575,N_1201,N_1200);
or U2576 (N_2576,N_1989,N_1373);
nand U2577 (N_2577,N_1378,N_1029);
and U2578 (N_2578,N_1469,N_1295);
and U2579 (N_2579,N_1496,N_1626);
and U2580 (N_2580,N_1513,N_1162);
nand U2581 (N_2581,N_1559,N_1851);
nand U2582 (N_2582,N_1111,N_1646);
nor U2583 (N_2583,N_1965,N_1556);
xor U2584 (N_2584,N_1582,N_1328);
nor U2585 (N_2585,N_1210,N_1816);
xnor U2586 (N_2586,N_1710,N_1612);
nor U2587 (N_2587,N_1558,N_1164);
nand U2588 (N_2588,N_1113,N_1272);
or U2589 (N_2589,N_1582,N_1473);
nor U2590 (N_2590,N_1966,N_1838);
or U2591 (N_2591,N_1748,N_1642);
nand U2592 (N_2592,N_1678,N_1029);
or U2593 (N_2593,N_1033,N_1679);
and U2594 (N_2594,N_1678,N_1557);
nor U2595 (N_2595,N_1480,N_1266);
nand U2596 (N_2596,N_1135,N_1881);
nor U2597 (N_2597,N_1329,N_1594);
nor U2598 (N_2598,N_1427,N_1718);
nand U2599 (N_2599,N_1165,N_1406);
nand U2600 (N_2600,N_1669,N_1297);
and U2601 (N_2601,N_1035,N_1371);
and U2602 (N_2602,N_1119,N_1660);
nor U2603 (N_2603,N_1401,N_1315);
or U2604 (N_2604,N_1446,N_1111);
nand U2605 (N_2605,N_1975,N_1480);
or U2606 (N_2606,N_1821,N_1697);
nor U2607 (N_2607,N_1866,N_1538);
and U2608 (N_2608,N_1063,N_1736);
nor U2609 (N_2609,N_1811,N_1519);
nor U2610 (N_2610,N_1908,N_1060);
nor U2611 (N_2611,N_1248,N_1909);
or U2612 (N_2612,N_1840,N_1710);
nand U2613 (N_2613,N_1628,N_1070);
nand U2614 (N_2614,N_1962,N_1571);
nand U2615 (N_2615,N_1220,N_1382);
or U2616 (N_2616,N_1925,N_1027);
or U2617 (N_2617,N_1870,N_1711);
and U2618 (N_2618,N_1994,N_1611);
nand U2619 (N_2619,N_1699,N_1792);
nand U2620 (N_2620,N_1216,N_1776);
or U2621 (N_2621,N_1072,N_1337);
and U2622 (N_2622,N_1560,N_1752);
and U2623 (N_2623,N_1454,N_1356);
nand U2624 (N_2624,N_1991,N_1400);
or U2625 (N_2625,N_1377,N_1875);
nand U2626 (N_2626,N_1188,N_1696);
or U2627 (N_2627,N_1877,N_1204);
nand U2628 (N_2628,N_1104,N_1761);
or U2629 (N_2629,N_1023,N_1238);
nor U2630 (N_2630,N_1847,N_1033);
or U2631 (N_2631,N_1794,N_1336);
nand U2632 (N_2632,N_1537,N_1222);
or U2633 (N_2633,N_1122,N_1343);
or U2634 (N_2634,N_1461,N_1020);
or U2635 (N_2635,N_1796,N_1732);
or U2636 (N_2636,N_1318,N_1810);
nand U2637 (N_2637,N_1422,N_1245);
nand U2638 (N_2638,N_1620,N_1052);
nor U2639 (N_2639,N_1408,N_1929);
and U2640 (N_2640,N_1361,N_1670);
nand U2641 (N_2641,N_1665,N_1043);
or U2642 (N_2642,N_1460,N_1895);
and U2643 (N_2643,N_1865,N_1467);
nand U2644 (N_2644,N_1151,N_1297);
or U2645 (N_2645,N_1395,N_1121);
or U2646 (N_2646,N_1493,N_1540);
nor U2647 (N_2647,N_1179,N_1438);
and U2648 (N_2648,N_1948,N_1859);
or U2649 (N_2649,N_1239,N_1387);
or U2650 (N_2650,N_1323,N_1599);
nand U2651 (N_2651,N_1183,N_1951);
nand U2652 (N_2652,N_1566,N_1478);
and U2653 (N_2653,N_1674,N_1878);
and U2654 (N_2654,N_1534,N_1529);
nand U2655 (N_2655,N_1687,N_1953);
nand U2656 (N_2656,N_1779,N_1427);
and U2657 (N_2657,N_1119,N_1245);
xor U2658 (N_2658,N_1396,N_1287);
nor U2659 (N_2659,N_1891,N_1331);
nand U2660 (N_2660,N_1960,N_1929);
nor U2661 (N_2661,N_1163,N_1304);
nand U2662 (N_2662,N_1787,N_1561);
and U2663 (N_2663,N_1948,N_1375);
nor U2664 (N_2664,N_1394,N_1689);
nand U2665 (N_2665,N_1860,N_1611);
nor U2666 (N_2666,N_1299,N_1918);
nor U2667 (N_2667,N_1068,N_1905);
nand U2668 (N_2668,N_1214,N_1514);
nor U2669 (N_2669,N_1156,N_1571);
xnor U2670 (N_2670,N_1241,N_1006);
nor U2671 (N_2671,N_1578,N_1964);
and U2672 (N_2672,N_1220,N_1919);
nor U2673 (N_2673,N_1885,N_1670);
or U2674 (N_2674,N_1458,N_1185);
or U2675 (N_2675,N_1957,N_1882);
nor U2676 (N_2676,N_1296,N_1615);
nor U2677 (N_2677,N_1661,N_1238);
and U2678 (N_2678,N_1150,N_1286);
nand U2679 (N_2679,N_1855,N_1754);
or U2680 (N_2680,N_1618,N_1176);
nor U2681 (N_2681,N_1427,N_1573);
and U2682 (N_2682,N_1477,N_1719);
nand U2683 (N_2683,N_1847,N_1538);
or U2684 (N_2684,N_1846,N_1530);
and U2685 (N_2685,N_1961,N_1098);
nand U2686 (N_2686,N_1952,N_1721);
or U2687 (N_2687,N_1999,N_1162);
or U2688 (N_2688,N_1289,N_1659);
or U2689 (N_2689,N_1534,N_1207);
nor U2690 (N_2690,N_1373,N_1053);
nand U2691 (N_2691,N_1088,N_1261);
and U2692 (N_2692,N_1927,N_1907);
nor U2693 (N_2693,N_1575,N_1849);
and U2694 (N_2694,N_1159,N_1904);
xor U2695 (N_2695,N_1417,N_1582);
xnor U2696 (N_2696,N_1743,N_1221);
nand U2697 (N_2697,N_1453,N_1259);
xor U2698 (N_2698,N_1222,N_1373);
nand U2699 (N_2699,N_1255,N_1746);
nand U2700 (N_2700,N_1354,N_1612);
nand U2701 (N_2701,N_1140,N_1937);
nand U2702 (N_2702,N_1125,N_1387);
nand U2703 (N_2703,N_1993,N_1556);
nand U2704 (N_2704,N_1024,N_1091);
nand U2705 (N_2705,N_1496,N_1729);
or U2706 (N_2706,N_1965,N_1711);
or U2707 (N_2707,N_1973,N_1706);
nand U2708 (N_2708,N_1885,N_1437);
nand U2709 (N_2709,N_1582,N_1306);
nand U2710 (N_2710,N_1721,N_1235);
or U2711 (N_2711,N_1971,N_1233);
or U2712 (N_2712,N_1506,N_1307);
nand U2713 (N_2713,N_1770,N_1424);
or U2714 (N_2714,N_1371,N_1626);
or U2715 (N_2715,N_1227,N_1368);
nor U2716 (N_2716,N_1196,N_1072);
and U2717 (N_2717,N_1767,N_1751);
nor U2718 (N_2718,N_1908,N_1972);
nand U2719 (N_2719,N_1235,N_1529);
nand U2720 (N_2720,N_1775,N_1628);
or U2721 (N_2721,N_1647,N_1292);
xnor U2722 (N_2722,N_1151,N_1005);
nand U2723 (N_2723,N_1031,N_1073);
and U2724 (N_2724,N_1600,N_1285);
or U2725 (N_2725,N_1590,N_1757);
nand U2726 (N_2726,N_1824,N_1669);
nor U2727 (N_2727,N_1244,N_1397);
nand U2728 (N_2728,N_1937,N_1563);
nor U2729 (N_2729,N_1071,N_1835);
or U2730 (N_2730,N_1194,N_1451);
nand U2731 (N_2731,N_1946,N_1811);
nand U2732 (N_2732,N_1115,N_1238);
or U2733 (N_2733,N_1781,N_1610);
nand U2734 (N_2734,N_1989,N_1526);
and U2735 (N_2735,N_1370,N_1118);
nand U2736 (N_2736,N_1440,N_1447);
nor U2737 (N_2737,N_1768,N_1611);
or U2738 (N_2738,N_1005,N_1934);
nor U2739 (N_2739,N_1566,N_1327);
nand U2740 (N_2740,N_1492,N_1122);
nand U2741 (N_2741,N_1894,N_1443);
and U2742 (N_2742,N_1546,N_1733);
nor U2743 (N_2743,N_1610,N_1426);
and U2744 (N_2744,N_1716,N_1314);
nor U2745 (N_2745,N_1679,N_1472);
xor U2746 (N_2746,N_1028,N_1452);
and U2747 (N_2747,N_1096,N_1845);
or U2748 (N_2748,N_1328,N_1985);
nor U2749 (N_2749,N_1402,N_1013);
or U2750 (N_2750,N_1214,N_1264);
and U2751 (N_2751,N_1399,N_1484);
and U2752 (N_2752,N_1100,N_1835);
nand U2753 (N_2753,N_1723,N_1367);
nor U2754 (N_2754,N_1066,N_1465);
and U2755 (N_2755,N_1373,N_1915);
nor U2756 (N_2756,N_1171,N_1152);
nand U2757 (N_2757,N_1466,N_1242);
and U2758 (N_2758,N_1950,N_1620);
or U2759 (N_2759,N_1270,N_1869);
nor U2760 (N_2760,N_1119,N_1856);
nand U2761 (N_2761,N_1329,N_1580);
or U2762 (N_2762,N_1827,N_1610);
nor U2763 (N_2763,N_1343,N_1449);
or U2764 (N_2764,N_1338,N_1321);
or U2765 (N_2765,N_1017,N_1610);
and U2766 (N_2766,N_1112,N_1532);
and U2767 (N_2767,N_1827,N_1007);
nand U2768 (N_2768,N_1423,N_1162);
xor U2769 (N_2769,N_1133,N_1123);
nor U2770 (N_2770,N_1711,N_1837);
or U2771 (N_2771,N_1508,N_1278);
nand U2772 (N_2772,N_1519,N_1994);
or U2773 (N_2773,N_1116,N_1947);
or U2774 (N_2774,N_1888,N_1934);
nor U2775 (N_2775,N_1459,N_1354);
nand U2776 (N_2776,N_1856,N_1887);
and U2777 (N_2777,N_1938,N_1530);
nand U2778 (N_2778,N_1525,N_1357);
nor U2779 (N_2779,N_1012,N_1140);
nor U2780 (N_2780,N_1324,N_1273);
nor U2781 (N_2781,N_1157,N_1590);
nand U2782 (N_2782,N_1131,N_1219);
and U2783 (N_2783,N_1495,N_1104);
nand U2784 (N_2784,N_1781,N_1613);
and U2785 (N_2785,N_1816,N_1897);
and U2786 (N_2786,N_1844,N_1660);
or U2787 (N_2787,N_1919,N_1615);
and U2788 (N_2788,N_1308,N_1476);
or U2789 (N_2789,N_1330,N_1777);
nand U2790 (N_2790,N_1492,N_1449);
nand U2791 (N_2791,N_1684,N_1884);
nand U2792 (N_2792,N_1681,N_1762);
and U2793 (N_2793,N_1195,N_1400);
and U2794 (N_2794,N_1967,N_1645);
and U2795 (N_2795,N_1994,N_1714);
or U2796 (N_2796,N_1142,N_1638);
nand U2797 (N_2797,N_1480,N_1555);
nand U2798 (N_2798,N_1142,N_1357);
nor U2799 (N_2799,N_1154,N_1349);
or U2800 (N_2800,N_1174,N_1260);
nor U2801 (N_2801,N_1300,N_1215);
or U2802 (N_2802,N_1618,N_1815);
nand U2803 (N_2803,N_1490,N_1973);
and U2804 (N_2804,N_1679,N_1734);
and U2805 (N_2805,N_1826,N_1123);
and U2806 (N_2806,N_1931,N_1253);
nor U2807 (N_2807,N_1370,N_1629);
nor U2808 (N_2808,N_1935,N_1328);
nor U2809 (N_2809,N_1316,N_1978);
nand U2810 (N_2810,N_1102,N_1785);
and U2811 (N_2811,N_1876,N_1187);
or U2812 (N_2812,N_1222,N_1469);
nor U2813 (N_2813,N_1830,N_1877);
nor U2814 (N_2814,N_1200,N_1407);
and U2815 (N_2815,N_1234,N_1934);
and U2816 (N_2816,N_1038,N_1666);
nand U2817 (N_2817,N_1480,N_1896);
nand U2818 (N_2818,N_1576,N_1089);
nor U2819 (N_2819,N_1461,N_1374);
or U2820 (N_2820,N_1000,N_1929);
nor U2821 (N_2821,N_1181,N_1800);
nand U2822 (N_2822,N_1393,N_1917);
or U2823 (N_2823,N_1825,N_1156);
and U2824 (N_2824,N_1273,N_1128);
and U2825 (N_2825,N_1033,N_1803);
xnor U2826 (N_2826,N_1641,N_1522);
nor U2827 (N_2827,N_1647,N_1019);
nor U2828 (N_2828,N_1560,N_1721);
nor U2829 (N_2829,N_1232,N_1947);
nand U2830 (N_2830,N_1333,N_1691);
or U2831 (N_2831,N_1674,N_1179);
and U2832 (N_2832,N_1408,N_1666);
and U2833 (N_2833,N_1303,N_1842);
nor U2834 (N_2834,N_1767,N_1057);
or U2835 (N_2835,N_1374,N_1604);
or U2836 (N_2836,N_1606,N_1402);
nand U2837 (N_2837,N_1319,N_1177);
or U2838 (N_2838,N_1986,N_1630);
or U2839 (N_2839,N_1638,N_1071);
and U2840 (N_2840,N_1280,N_1956);
and U2841 (N_2841,N_1054,N_1731);
nand U2842 (N_2842,N_1648,N_1157);
nor U2843 (N_2843,N_1121,N_1365);
and U2844 (N_2844,N_1033,N_1387);
and U2845 (N_2845,N_1127,N_1290);
nor U2846 (N_2846,N_1250,N_1054);
and U2847 (N_2847,N_1974,N_1044);
and U2848 (N_2848,N_1933,N_1719);
or U2849 (N_2849,N_1178,N_1939);
or U2850 (N_2850,N_1627,N_1297);
and U2851 (N_2851,N_1691,N_1199);
or U2852 (N_2852,N_1417,N_1051);
or U2853 (N_2853,N_1762,N_1826);
or U2854 (N_2854,N_1652,N_1703);
nor U2855 (N_2855,N_1696,N_1549);
nand U2856 (N_2856,N_1033,N_1981);
nand U2857 (N_2857,N_1580,N_1181);
xor U2858 (N_2858,N_1362,N_1204);
or U2859 (N_2859,N_1747,N_1860);
or U2860 (N_2860,N_1047,N_1541);
nand U2861 (N_2861,N_1199,N_1587);
or U2862 (N_2862,N_1023,N_1128);
nand U2863 (N_2863,N_1077,N_1873);
and U2864 (N_2864,N_1355,N_1941);
and U2865 (N_2865,N_1270,N_1986);
or U2866 (N_2866,N_1688,N_1398);
nand U2867 (N_2867,N_1536,N_1007);
or U2868 (N_2868,N_1327,N_1483);
nand U2869 (N_2869,N_1105,N_1192);
or U2870 (N_2870,N_1159,N_1574);
or U2871 (N_2871,N_1099,N_1369);
or U2872 (N_2872,N_1762,N_1299);
nand U2873 (N_2873,N_1894,N_1545);
nor U2874 (N_2874,N_1356,N_1275);
and U2875 (N_2875,N_1119,N_1298);
nor U2876 (N_2876,N_1629,N_1674);
and U2877 (N_2877,N_1830,N_1529);
and U2878 (N_2878,N_1258,N_1678);
or U2879 (N_2879,N_1133,N_1843);
nor U2880 (N_2880,N_1726,N_1890);
and U2881 (N_2881,N_1631,N_1996);
and U2882 (N_2882,N_1103,N_1827);
and U2883 (N_2883,N_1887,N_1007);
nor U2884 (N_2884,N_1814,N_1669);
or U2885 (N_2885,N_1913,N_1833);
nand U2886 (N_2886,N_1745,N_1735);
and U2887 (N_2887,N_1495,N_1252);
and U2888 (N_2888,N_1178,N_1753);
nor U2889 (N_2889,N_1565,N_1769);
or U2890 (N_2890,N_1454,N_1904);
nand U2891 (N_2891,N_1130,N_1284);
xnor U2892 (N_2892,N_1469,N_1176);
nand U2893 (N_2893,N_1658,N_1022);
or U2894 (N_2894,N_1373,N_1344);
nand U2895 (N_2895,N_1702,N_1978);
or U2896 (N_2896,N_1711,N_1019);
nand U2897 (N_2897,N_1714,N_1221);
or U2898 (N_2898,N_1315,N_1668);
or U2899 (N_2899,N_1579,N_1103);
or U2900 (N_2900,N_1637,N_1383);
nor U2901 (N_2901,N_1037,N_1802);
or U2902 (N_2902,N_1610,N_1912);
nand U2903 (N_2903,N_1388,N_1970);
nor U2904 (N_2904,N_1289,N_1087);
and U2905 (N_2905,N_1196,N_1783);
or U2906 (N_2906,N_1770,N_1804);
and U2907 (N_2907,N_1227,N_1158);
nand U2908 (N_2908,N_1885,N_1714);
nor U2909 (N_2909,N_1878,N_1469);
nor U2910 (N_2910,N_1829,N_1669);
and U2911 (N_2911,N_1173,N_1468);
or U2912 (N_2912,N_1651,N_1595);
or U2913 (N_2913,N_1217,N_1271);
nor U2914 (N_2914,N_1241,N_1526);
and U2915 (N_2915,N_1454,N_1208);
and U2916 (N_2916,N_1881,N_1400);
xnor U2917 (N_2917,N_1069,N_1817);
nor U2918 (N_2918,N_1538,N_1834);
nor U2919 (N_2919,N_1967,N_1011);
and U2920 (N_2920,N_1776,N_1305);
nand U2921 (N_2921,N_1748,N_1613);
or U2922 (N_2922,N_1616,N_1959);
nor U2923 (N_2923,N_1621,N_1689);
or U2924 (N_2924,N_1858,N_1775);
and U2925 (N_2925,N_1453,N_1672);
and U2926 (N_2926,N_1732,N_1261);
and U2927 (N_2927,N_1758,N_1200);
or U2928 (N_2928,N_1624,N_1301);
or U2929 (N_2929,N_1770,N_1030);
nor U2930 (N_2930,N_1576,N_1969);
or U2931 (N_2931,N_1609,N_1339);
nor U2932 (N_2932,N_1061,N_1487);
and U2933 (N_2933,N_1889,N_1387);
nor U2934 (N_2934,N_1474,N_1323);
or U2935 (N_2935,N_1922,N_1349);
nor U2936 (N_2936,N_1592,N_1206);
or U2937 (N_2937,N_1006,N_1269);
nor U2938 (N_2938,N_1052,N_1601);
xor U2939 (N_2939,N_1642,N_1017);
nor U2940 (N_2940,N_1444,N_1023);
nor U2941 (N_2941,N_1409,N_1772);
and U2942 (N_2942,N_1943,N_1809);
and U2943 (N_2943,N_1508,N_1494);
and U2944 (N_2944,N_1647,N_1757);
nand U2945 (N_2945,N_1529,N_1415);
nor U2946 (N_2946,N_1249,N_1120);
and U2947 (N_2947,N_1941,N_1720);
and U2948 (N_2948,N_1426,N_1977);
and U2949 (N_2949,N_1095,N_1475);
nor U2950 (N_2950,N_1589,N_1050);
and U2951 (N_2951,N_1400,N_1418);
and U2952 (N_2952,N_1214,N_1298);
nand U2953 (N_2953,N_1851,N_1420);
or U2954 (N_2954,N_1189,N_1396);
nor U2955 (N_2955,N_1720,N_1752);
nand U2956 (N_2956,N_1851,N_1211);
xor U2957 (N_2957,N_1605,N_1627);
nand U2958 (N_2958,N_1530,N_1453);
nand U2959 (N_2959,N_1765,N_1527);
and U2960 (N_2960,N_1004,N_1597);
or U2961 (N_2961,N_1465,N_1459);
and U2962 (N_2962,N_1747,N_1651);
nand U2963 (N_2963,N_1882,N_1642);
nor U2964 (N_2964,N_1834,N_1387);
and U2965 (N_2965,N_1355,N_1281);
and U2966 (N_2966,N_1987,N_1386);
nand U2967 (N_2967,N_1697,N_1667);
nand U2968 (N_2968,N_1568,N_1508);
and U2969 (N_2969,N_1030,N_1758);
or U2970 (N_2970,N_1742,N_1126);
nand U2971 (N_2971,N_1537,N_1715);
and U2972 (N_2972,N_1883,N_1462);
nand U2973 (N_2973,N_1501,N_1610);
nand U2974 (N_2974,N_1617,N_1816);
and U2975 (N_2975,N_1541,N_1925);
nor U2976 (N_2976,N_1132,N_1645);
and U2977 (N_2977,N_1368,N_1750);
and U2978 (N_2978,N_1455,N_1056);
nor U2979 (N_2979,N_1158,N_1459);
nor U2980 (N_2980,N_1464,N_1626);
nand U2981 (N_2981,N_1422,N_1085);
and U2982 (N_2982,N_1394,N_1931);
nor U2983 (N_2983,N_1307,N_1705);
nor U2984 (N_2984,N_1578,N_1567);
nand U2985 (N_2985,N_1066,N_1224);
nor U2986 (N_2986,N_1859,N_1675);
or U2987 (N_2987,N_1961,N_1661);
or U2988 (N_2988,N_1840,N_1449);
nor U2989 (N_2989,N_1994,N_1089);
nor U2990 (N_2990,N_1573,N_1624);
or U2991 (N_2991,N_1765,N_1374);
nor U2992 (N_2992,N_1427,N_1132);
xnor U2993 (N_2993,N_1309,N_1743);
nand U2994 (N_2994,N_1487,N_1536);
or U2995 (N_2995,N_1634,N_1010);
nor U2996 (N_2996,N_1660,N_1883);
or U2997 (N_2997,N_1036,N_1043);
nor U2998 (N_2998,N_1176,N_1214);
or U2999 (N_2999,N_1473,N_1718);
nand U3000 (N_3000,N_2456,N_2063);
or U3001 (N_3001,N_2373,N_2277);
nand U3002 (N_3002,N_2648,N_2255);
nand U3003 (N_3003,N_2442,N_2678);
or U3004 (N_3004,N_2332,N_2553);
nor U3005 (N_3005,N_2288,N_2961);
nand U3006 (N_3006,N_2409,N_2374);
nor U3007 (N_3007,N_2851,N_2148);
and U3008 (N_3008,N_2355,N_2054);
nand U3009 (N_3009,N_2938,N_2386);
nor U3010 (N_3010,N_2976,N_2833);
nand U3011 (N_3011,N_2715,N_2001);
xnor U3012 (N_3012,N_2852,N_2778);
or U3013 (N_3013,N_2311,N_2835);
nor U3014 (N_3014,N_2837,N_2800);
and U3015 (N_3015,N_2999,N_2017);
and U3016 (N_3016,N_2049,N_2330);
nor U3017 (N_3017,N_2586,N_2843);
nand U3018 (N_3018,N_2081,N_2686);
and U3019 (N_3019,N_2875,N_2031);
nor U3020 (N_3020,N_2703,N_2015);
nand U3021 (N_3021,N_2014,N_2224);
nand U3022 (N_3022,N_2137,N_2593);
nor U3023 (N_3023,N_2873,N_2499);
and U3024 (N_3024,N_2067,N_2289);
nor U3025 (N_3025,N_2050,N_2786);
nand U3026 (N_3026,N_2170,N_2423);
xnor U3027 (N_3027,N_2662,N_2676);
nand U3028 (N_3028,N_2810,N_2395);
or U3029 (N_3029,N_2460,N_2735);
or U3030 (N_3030,N_2186,N_2155);
or U3031 (N_3031,N_2482,N_2193);
nand U3032 (N_3032,N_2472,N_2891);
and U3033 (N_3033,N_2839,N_2298);
or U3034 (N_3034,N_2190,N_2044);
or U3035 (N_3035,N_2559,N_2942);
or U3036 (N_3036,N_2093,N_2181);
or U3037 (N_3037,N_2591,N_2751);
nor U3038 (N_3038,N_2731,N_2579);
nor U3039 (N_3039,N_2892,N_2799);
nand U3040 (N_3040,N_2932,N_2016);
and U3041 (N_3041,N_2514,N_2466);
and U3042 (N_3042,N_2422,N_2790);
nand U3043 (N_3043,N_2085,N_2232);
nand U3044 (N_3044,N_2398,N_2635);
and U3045 (N_3045,N_2139,N_2073);
or U3046 (N_3046,N_2366,N_2037);
and U3047 (N_3047,N_2177,N_2485);
or U3048 (N_3048,N_2578,N_2996);
nor U3049 (N_3049,N_2838,N_2457);
nor U3050 (N_3050,N_2397,N_2997);
nor U3051 (N_3051,N_2526,N_2825);
nor U3052 (N_3052,N_2087,N_2071);
nor U3053 (N_3053,N_2147,N_2216);
or U3054 (N_3054,N_2122,N_2237);
nand U3055 (N_3055,N_2534,N_2967);
and U3056 (N_3056,N_2639,N_2069);
or U3057 (N_3057,N_2502,N_2336);
or U3058 (N_3058,N_2141,N_2744);
nand U3059 (N_3059,N_2506,N_2279);
and U3060 (N_3060,N_2757,N_2107);
nand U3061 (N_3061,N_2441,N_2354);
or U3062 (N_3062,N_2072,N_2674);
nor U3063 (N_3063,N_2035,N_2975);
nor U3064 (N_3064,N_2937,N_2401);
nand U3065 (N_3065,N_2117,N_2536);
or U3066 (N_3066,N_2769,N_2617);
xnor U3067 (N_3067,N_2042,N_2483);
and U3068 (N_3068,N_2859,N_2969);
or U3069 (N_3069,N_2416,N_2740);
nand U3070 (N_3070,N_2248,N_2023);
or U3071 (N_3071,N_2161,N_2732);
and U3072 (N_3072,N_2677,N_2914);
or U3073 (N_3073,N_2913,N_2840);
or U3074 (N_3074,N_2105,N_2078);
and U3075 (N_3075,N_2251,N_2325);
or U3076 (N_3076,N_2135,N_2206);
and U3077 (N_3077,N_2595,N_2100);
or U3078 (N_3078,N_2813,N_2971);
nor U3079 (N_3079,N_2758,N_2296);
and U3080 (N_3080,N_2712,N_2909);
or U3081 (N_3081,N_2588,N_2644);
nand U3082 (N_3082,N_2259,N_2104);
nand U3083 (N_3083,N_2622,N_2737);
nor U3084 (N_3084,N_2831,N_2657);
nor U3085 (N_3085,N_2267,N_2434);
and U3086 (N_3086,N_2538,N_2749);
and U3087 (N_3087,N_2973,N_2106);
and U3088 (N_3088,N_2565,N_2558);
or U3089 (N_3089,N_2360,N_2992);
nand U3090 (N_3090,N_2609,N_2201);
nand U3091 (N_3091,N_2675,N_2022);
or U3092 (N_3092,N_2064,N_2086);
nor U3093 (N_3093,N_2128,N_2817);
nand U3094 (N_3094,N_2488,N_2291);
nor U3095 (N_3095,N_2858,N_2082);
and U3096 (N_3096,N_2214,N_2504);
or U3097 (N_3097,N_2763,N_2556);
and U3098 (N_3098,N_2908,N_2124);
nand U3099 (N_3099,N_2865,N_2174);
nand U3100 (N_3100,N_2853,N_2295);
nand U3101 (N_3101,N_2682,N_2818);
or U3102 (N_3102,N_2263,N_2467);
nor U3103 (N_3103,N_2782,N_2789);
nor U3104 (N_3104,N_2464,N_2238);
and U3105 (N_3105,N_2356,N_2946);
or U3106 (N_3106,N_2119,N_2702);
nor U3107 (N_3107,N_2221,N_2358);
nand U3108 (N_3108,N_2560,N_2977);
and U3109 (N_3109,N_2529,N_2690);
nor U3110 (N_3110,N_2681,N_2884);
nand U3111 (N_3111,N_2965,N_2191);
nand U3112 (N_3112,N_2384,N_2555);
nand U3113 (N_3113,N_2144,N_2256);
nor U3114 (N_3114,N_2792,N_2981);
nand U3115 (N_3115,N_2739,N_2099);
nand U3116 (N_3116,N_2003,N_2796);
nor U3117 (N_3117,N_2222,N_2955);
nand U3118 (N_3118,N_2521,N_2889);
and U3119 (N_3119,N_2604,N_2945);
or U3120 (N_3120,N_2804,N_2006);
nand U3121 (N_3121,N_2077,N_2590);
nor U3122 (N_3122,N_2315,N_2807);
or U3123 (N_3123,N_2797,N_2663);
nor U3124 (N_3124,N_2376,N_2623);
nor U3125 (N_3125,N_2653,N_2306);
or U3126 (N_3126,N_2949,N_2684);
or U3127 (N_3127,N_2794,N_2723);
and U3128 (N_3128,N_2138,N_2727);
xor U3129 (N_3129,N_2820,N_2448);
xnor U3130 (N_3130,N_2661,N_2136);
nor U3131 (N_3131,N_2822,N_2115);
or U3132 (N_3132,N_2664,N_2948);
or U3133 (N_3133,N_2246,N_2869);
and U3134 (N_3134,N_2930,N_2343);
nor U3135 (N_3135,N_2519,N_2030);
or U3136 (N_3136,N_2926,N_2683);
nand U3137 (N_3137,N_2540,N_2882);
nor U3138 (N_3138,N_2369,N_2584);
nand U3139 (N_3139,N_2812,N_2305);
nor U3140 (N_3140,N_2525,N_2610);
nor U3141 (N_3141,N_2152,N_2211);
and U3142 (N_3142,N_2435,N_2647);
and U3143 (N_3143,N_2987,N_2912);
or U3144 (N_3144,N_2929,N_2140);
nand U3145 (N_3145,N_2862,N_2509);
nand U3146 (N_3146,N_2057,N_2951);
and U3147 (N_3147,N_2405,N_2984);
or U3148 (N_3148,N_2847,N_2611);
nand U3149 (N_3149,N_2012,N_2189);
nor U3150 (N_3150,N_2312,N_2826);
nand U3151 (N_3151,N_2258,N_2752);
and U3152 (N_3152,N_2013,N_2780);
or U3153 (N_3153,N_2308,N_2156);
nand U3154 (N_3154,N_2024,N_2208);
or U3155 (N_3155,N_2824,N_2922);
nand U3156 (N_3156,N_2539,N_2243);
or U3157 (N_3157,N_2303,N_2787);
nand U3158 (N_3158,N_2645,N_2530);
nand U3159 (N_3159,N_2413,N_2785);
or U3160 (N_3160,N_2299,N_2041);
xnor U3161 (N_3161,N_2449,N_2445);
nand U3162 (N_3162,N_2349,N_2959);
and U3163 (N_3163,N_2979,N_2532);
nor U3164 (N_3164,N_2020,N_2097);
and U3165 (N_3165,N_2387,N_2272);
and U3166 (N_3166,N_2480,N_2692);
and U3167 (N_3167,N_2439,N_2229);
nor U3168 (N_3168,N_2285,N_2444);
nor U3169 (N_3169,N_2890,N_2348);
and U3170 (N_3170,N_2130,N_2005);
nand U3171 (N_3171,N_2867,N_2187);
and U3172 (N_3172,N_2832,N_2425);
nor U3173 (N_3173,N_2666,N_2885);
or U3174 (N_3174,N_2742,N_2252);
or U3175 (N_3175,N_2950,N_2471);
and U3176 (N_3176,N_2700,N_2283);
and U3177 (N_3177,N_2379,N_2755);
and U3178 (N_3178,N_2596,N_2173);
and U3179 (N_3179,N_2705,N_2513);
and U3180 (N_3180,N_2944,N_2562);
and U3181 (N_3181,N_2043,N_2178);
nand U3182 (N_3182,N_2748,N_2845);
or U3183 (N_3183,N_2209,N_2324);
or U3184 (N_3184,N_2581,N_2383);
or U3185 (N_3185,N_2364,N_2627);
nand U3186 (N_3186,N_2307,N_2956);
or U3187 (N_3187,N_2327,N_2096);
or U3188 (N_3188,N_2432,N_2300);
nand U3189 (N_3189,N_2265,N_2510);
or U3190 (N_3190,N_2320,N_2402);
and U3191 (N_3191,N_2098,N_2322);
nor U3192 (N_3192,N_2347,N_2109);
and U3193 (N_3193,N_2192,N_2293);
or U3194 (N_3194,N_2989,N_2494);
nor U3195 (N_3195,N_2032,N_2458);
and U3196 (N_3196,N_2074,N_2353);
and U3197 (N_3197,N_2533,N_2271);
nand U3198 (N_3198,N_2228,N_2543);
or U3199 (N_3199,N_2378,N_2110);
nand U3200 (N_3200,N_2428,N_2365);
and U3201 (N_3201,N_2507,N_2011);
nor U3202 (N_3202,N_2287,N_2166);
and U3203 (N_3203,N_2694,N_2916);
and U3204 (N_3204,N_2795,N_2297);
and U3205 (N_3205,N_2991,N_2410);
and U3206 (N_3206,N_2180,N_2046);
nand U3207 (N_3207,N_2709,N_2550);
nor U3208 (N_3208,N_2185,N_2931);
or U3209 (N_3209,N_2933,N_2842);
nor U3210 (N_3210,N_2339,N_2814);
nand U3211 (N_3211,N_2462,N_2415);
nor U3212 (N_3212,N_2094,N_2004);
nor U3213 (N_3213,N_2698,N_2326);
or U3214 (N_3214,N_2768,N_2990);
nor U3215 (N_3215,N_2809,N_2433);
or U3216 (N_3216,N_2895,N_2985);
and U3217 (N_3217,N_2284,N_2888);
and U3218 (N_3218,N_2952,N_2253);
or U3219 (N_3219,N_2566,N_2220);
and U3220 (N_3220,N_2631,N_2132);
and U3221 (N_3221,N_2158,N_2417);
nand U3222 (N_3222,N_2823,N_2045);
nor U3223 (N_3223,N_2947,N_2879);
and U3224 (N_3224,N_2145,N_2338);
nand U3225 (N_3225,N_2655,N_2651);
nand U3226 (N_3226,N_2090,N_2620);
nor U3227 (N_3227,N_2188,N_2427);
and U3228 (N_3228,N_2350,N_2134);
nor U3229 (N_3229,N_2501,N_2034);
or U3230 (N_3230,N_2028,N_2587);
or U3231 (N_3231,N_2828,N_2515);
nand U3232 (N_3232,N_2000,N_2870);
nand U3233 (N_3233,N_2547,N_2375);
nand U3234 (N_3234,N_2286,N_2025);
or U3235 (N_3235,N_2669,N_2541);
nor U3236 (N_3236,N_2414,N_2598);
nor U3237 (N_3237,N_2125,N_2247);
nor U3238 (N_3238,N_2245,N_2738);
or U3239 (N_3239,N_2928,N_2318);
and U3240 (N_3240,N_2710,N_2239);
nand U3241 (N_3241,N_2537,N_2450);
and U3242 (N_3242,N_2089,N_2871);
xnor U3243 (N_3243,N_2592,N_2704);
nor U3244 (N_3244,N_2771,N_2759);
or U3245 (N_3245,N_2774,N_2146);
or U3246 (N_3246,N_2223,N_2168);
or U3247 (N_3247,N_2699,N_2418);
nand U3248 (N_3248,N_2524,N_2461);
nor U3249 (N_3249,N_2359,N_2629);
nand U3250 (N_3250,N_2493,N_2010);
nand U3251 (N_3251,N_2717,N_2301);
and U3252 (N_3252,N_2554,N_2009);
or U3253 (N_3253,N_2390,N_2898);
nor U3254 (N_3254,N_2688,N_2172);
or U3255 (N_3255,N_2061,N_2345);
nand U3256 (N_3256,N_2150,N_2470);
or U3257 (N_3257,N_2491,N_2159);
and U3258 (N_3258,N_2827,N_2630);
and U3259 (N_3259,N_2380,N_2207);
or U3260 (N_3260,N_2492,N_2056);
nand U3261 (N_3261,N_2679,N_2528);
or U3262 (N_3262,N_2169,N_2029);
and U3263 (N_3263,N_2557,N_2954);
nor U3264 (N_3264,N_2143,N_2517);
or U3265 (N_3265,N_2924,N_2021);
nor U3266 (N_3266,N_2872,N_2563);
and U3267 (N_3267,N_2603,N_2811);
nor U3268 (N_3268,N_2070,N_2841);
nand U3269 (N_3269,N_2943,N_2235);
nand U3270 (N_3270,N_2478,N_2652);
nor U3271 (N_3271,N_2575,N_2511);
or U3272 (N_3272,N_2430,N_2079);
or U3273 (N_3273,N_2716,N_2408);
nor U3274 (N_3274,N_2254,N_2725);
nand U3275 (N_3275,N_2846,N_2545);
or U3276 (N_3276,N_2850,N_2278);
or U3277 (N_3277,N_2876,N_2970);
or U3278 (N_3278,N_2665,N_2608);
nand U3279 (N_3279,N_2936,N_2120);
nor U3280 (N_3280,N_2261,N_2420);
or U3281 (N_3281,N_2062,N_2018);
nor U3282 (N_3282,N_2570,N_2002);
nand U3283 (N_3283,N_2199,N_2121);
and U3284 (N_3284,N_2446,N_2400);
or U3285 (N_3285,N_2151,N_2750);
or U3286 (N_3286,N_2549,N_2512);
or U3287 (N_3287,N_2249,N_2861);
nand U3288 (N_3288,N_2231,N_2476);
nand U3289 (N_3289,N_2329,N_2495);
nor U3290 (N_3290,N_2624,N_2227);
and U3291 (N_3291,N_2399,N_2197);
nor U3292 (N_3292,N_2689,N_2368);
xor U3293 (N_3293,N_2244,N_2920);
nand U3294 (N_3294,N_2806,N_2372);
or U3295 (N_3295,N_2571,N_2815);
and U3296 (N_3296,N_2982,N_2585);
nand U3297 (N_3297,N_2848,N_2864);
nor U3298 (N_3298,N_2048,N_2334);
nand U3299 (N_3299,N_2801,N_2691);
and U3300 (N_3300,N_2076,N_2724);
nor U3301 (N_3301,N_2773,N_2654);
and U3302 (N_3302,N_2719,N_2743);
nand U3303 (N_3303,N_2335,N_2520);
or U3304 (N_3304,N_2443,N_2276);
or U3305 (N_3305,N_2438,N_2791);
or U3306 (N_3306,N_2607,N_2998);
and U3307 (N_3307,N_2344,N_2883);
nor U3308 (N_3308,N_2941,N_2381);
and U3309 (N_3309,N_2706,N_2426);
and U3310 (N_3310,N_2972,N_2849);
and U3311 (N_3311,N_2068,N_2756);
and U3312 (N_3312,N_2357,N_2963);
and U3313 (N_3313,N_2396,N_2685);
nor U3314 (N_3314,N_2204,N_2129);
and U3315 (N_3315,N_2091,N_2784);
and U3316 (N_3316,N_2370,N_2116);
xor U3317 (N_3317,N_2918,N_2382);
nor U3318 (N_3318,N_2745,N_2798);
and U3319 (N_3319,N_2707,N_2060);
and U3320 (N_3320,N_2126,N_2899);
and U3321 (N_3321,N_2900,N_2233);
or U3322 (N_3322,N_2361,N_2781);
nand U3323 (N_3323,N_2213,N_2726);
nor U3324 (N_3324,N_2182,N_2280);
and U3325 (N_3325,N_2101,N_2160);
or U3326 (N_3326,N_2551,N_2477);
xnor U3327 (N_3327,N_2114,N_2874);
and U3328 (N_3328,N_2219,N_2292);
nor U3329 (N_3329,N_2452,N_2646);
and U3330 (N_3330,N_2266,N_2194);
and U3331 (N_3331,N_2741,N_2108);
or U3332 (N_3332,N_2393,N_2616);
and U3333 (N_3333,N_2388,N_2896);
or U3334 (N_3334,N_2816,N_2092);
nor U3335 (N_3335,N_2680,N_2281);
nand U3336 (N_3336,N_2331,N_2634);
nand U3337 (N_3337,N_2564,N_2978);
or U3338 (N_3338,N_2866,N_2055);
and U3339 (N_3339,N_2403,N_2764);
and U3340 (N_3340,N_2671,N_2226);
and U3341 (N_3341,N_2176,N_2275);
or U3342 (N_3342,N_2118,N_2019);
or U3343 (N_3343,N_2260,N_2437);
nor U3344 (N_3344,N_2516,N_2974);
nor U3345 (N_3345,N_2660,N_2760);
nor U3346 (N_3346,N_2459,N_2039);
and U3347 (N_3347,N_2167,N_2650);
nor U3348 (N_3348,N_2638,N_2567);
and U3349 (N_3349,N_2316,N_2241);
nand U3350 (N_3350,N_2910,N_2465);
or U3351 (N_3351,N_2917,N_2496);
or U3352 (N_3352,N_2632,N_2656);
nor U3353 (N_3353,N_2641,N_2600);
or U3354 (N_3354,N_2202,N_2886);
xnor U3355 (N_3355,N_2153,N_2589);
or U3356 (N_3356,N_2200,N_2636);
or U3357 (N_3357,N_2487,N_2195);
or U3358 (N_3358,N_2649,N_2988);
nand U3359 (N_3359,N_2095,N_2854);
or U3360 (N_3360,N_2033,N_2819);
nand U3361 (N_3361,N_2407,N_2489);
or U3362 (N_3362,N_2730,N_2340);
and U3363 (N_3363,N_2940,N_2788);
and U3364 (N_3364,N_2154,N_2337);
nand U3365 (N_3365,N_2040,N_2421);
nand U3366 (N_3366,N_2614,N_2980);
nand U3367 (N_3367,N_2203,N_2844);
nor U3368 (N_3368,N_2569,N_2602);
or U3369 (N_3369,N_2860,N_2583);
and U3370 (N_3370,N_2803,N_2429);
nor U3371 (N_3371,N_2453,N_2323);
xor U3372 (N_3372,N_2994,N_2775);
nor U3373 (N_3373,N_2572,N_2412);
and U3374 (N_3374,N_2346,N_2310);
nor U3375 (N_3375,N_2268,N_2294);
nand U3376 (N_3376,N_2230,N_2080);
and U3377 (N_3377,N_2568,N_2451);
or U3378 (N_3378,N_2594,N_2389);
and U3379 (N_3379,N_2905,N_2953);
or U3380 (N_3380,N_2834,N_2038);
and U3381 (N_3381,N_2927,N_2102);
and U3382 (N_3382,N_2149,N_2915);
and U3383 (N_3383,N_2454,N_2321);
or U3384 (N_3384,N_2576,N_2317);
and U3385 (N_3385,N_2436,N_2274);
nor U3386 (N_3386,N_2469,N_2907);
xnor U3387 (N_3387,N_2342,N_2262);
and U3388 (N_3388,N_2212,N_2269);
nor U3389 (N_3389,N_2314,N_2103);
xor U3390 (N_3390,N_2903,N_2793);
nand U3391 (N_3391,N_2720,N_2234);
nor U3392 (N_3392,N_2242,N_2642);
or U3393 (N_3393,N_2830,N_2779);
nor U3394 (N_3394,N_2290,N_2618);
or U3395 (N_3395,N_2754,N_2887);
and U3396 (N_3396,N_2508,N_2475);
and U3397 (N_3397,N_2198,N_2966);
nand U3398 (N_3398,N_2766,N_2419);
or U3399 (N_3399,N_2385,N_2687);
or U3400 (N_3400,N_2761,N_2184);
or U3401 (N_3401,N_2697,N_2729);
nand U3402 (N_3402,N_2264,N_2746);
nand U3403 (N_3403,N_2058,N_2597);
and U3404 (N_3404,N_2580,N_2767);
nor U3405 (N_3405,N_2552,N_2696);
nor U3406 (N_3406,N_2670,N_2765);
nand U3407 (N_3407,N_2855,N_2500);
or U3408 (N_3408,N_2431,N_2701);
nand U3409 (N_3409,N_2829,N_2599);
nand U3410 (N_3410,N_2490,N_2394);
nor U3411 (N_3411,N_2047,N_2574);
nor U3412 (N_3412,N_2821,N_2406);
or U3413 (N_3413,N_2721,N_2210);
xor U3414 (N_3414,N_2911,N_2171);
nor U3415 (N_3415,N_2225,N_2309);
nor U3416 (N_3416,N_2411,N_2051);
or U3417 (N_3417,N_2066,N_2919);
nand U3418 (N_3418,N_2612,N_2205);
and U3419 (N_3419,N_2783,N_2217);
nand U3420 (N_3420,N_2133,N_2333);
nor U3421 (N_3421,N_2906,N_2633);
nand U3422 (N_3422,N_2548,N_2625);
or U3423 (N_3423,N_2363,N_2440);
nand U3424 (N_3424,N_2711,N_2362);
xnor U3425 (N_3425,N_2934,N_2313);
and U3426 (N_3426,N_2179,N_2083);
nand U3427 (N_3427,N_2236,N_2960);
nor U3428 (N_3428,N_2628,N_2527);
or U3429 (N_3429,N_2218,N_2486);
and U3430 (N_3430,N_2542,N_2753);
and U3431 (N_3431,N_2772,N_2673);
or U3432 (N_3432,N_2868,N_2957);
or U3433 (N_3433,N_2498,N_2111);
and U3434 (N_3434,N_2481,N_2695);
nand U3435 (N_3435,N_2718,N_2052);
nor U3436 (N_3436,N_2606,N_2518);
and U3437 (N_3437,N_2923,N_2036);
nor U3438 (N_3438,N_2007,N_2112);
or U3439 (N_3439,N_2546,N_2157);
or U3440 (N_3440,N_2881,N_2164);
nor U3441 (N_3441,N_2352,N_2626);
xnor U3442 (N_3442,N_2165,N_2659);
nand U3443 (N_3443,N_2708,N_2802);
and U3444 (N_3444,N_2505,N_2319);
nor U3445 (N_3445,N_2503,N_2939);
or U3446 (N_3446,N_2474,N_2544);
and U3447 (N_3447,N_2672,N_2113);
nand U3448 (N_3448,N_2270,N_2777);
nor U3449 (N_3449,N_2601,N_2282);
nor U3450 (N_3450,N_2728,N_2668);
or U3451 (N_3451,N_2484,N_2273);
or U3452 (N_3452,N_2523,N_2183);
and U3453 (N_3453,N_2531,N_2131);
or U3454 (N_3454,N_2605,N_2535);
xnor U3455 (N_3455,N_2175,N_2993);
nor U3456 (N_3456,N_2084,N_2734);
nor U3457 (N_3457,N_2857,N_2667);
and U3458 (N_3458,N_2658,N_2561);
or U3459 (N_3459,N_2075,N_2962);
nand U3460 (N_3460,N_2733,N_2302);
nor U3461 (N_3461,N_2776,N_2897);
or U3462 (N_3462,N_2613,N_2479);
or U3463 (N_3463,N_2747,N_2856);
nand U3464 (N_3464,N_2722,N_2964);
nand U3465 (N_3465,N_2473,N_2162);
nand U3466 (N_3466,N_2770,N_2925);
nor U3467 (N_3467,N_2880,N_2059);
nand U3468 (N_3468,N_2065,N_2983);
nand U3469 (N_3469,N_2304,N_2582);
or U3470 (N_3470,N_2455,N_2377);
or U3471 (N_3471,N_2736,N_2878);
or U3472 (N_3472,N_2714,N_2901);
or U3473 (N_3473,N_2424,N_2935);
or U3474 (N_3474,N_2026,N_2637);
or U3475 (N_3475,N_2693,N_2391);
nand U3476 (N_3476,N_2894,N_2497);
xnor U3477 (N_3477,N_2215,N_2573);
nand U3478 (N_3478,N_2008,N_2088);
nand U3479 (N_3479,N_2902,N_2522);
and U3480 (N_3480,N_2196,N_2836);
nor U3481 (N_3481,N_2328,N_2762);
or U3482 (N_3482,N_2351,N_2123);
and U3483 (N_3483,N_2643,N_2619);
and U3484 (N_3484,N_2250,N_2257);
nor U3485 (N_3485,N_2404,N_2163);
and U3486 (N_3486,N_2863,N_2463);
nand U3487 (N_3487,N_2053,N_2640);
nand U3488 (N_3488,N_2615,N_2921);
nor U3489 (N_3489,N_2877,N_2027);
nand U3490 (N_3490,N_2127,N_2968);
nand U3491 (N_3491,N_2808,N_2447);
and U3492 (N_3492,N_2893,N_2805);
and U3493 (N_3493,N_2986,N_2958);
and U3494 (N_3494,N_2713,N_2240);
and U3495 (N_3495,N_2341,N_2142);
or U3496 (N_3496,N_2621,N_2367);
or U3497 (N_3497,N_2371,N_2904);
or U3498 (N_3498,N_2392,N_2995);
nand U3499 (N_3499,N_2468,N_2577);
nand U3500 (N_3500,N_2952,N_2301);
and U3501 (N_3501,N_2377,N_2808);
nand U3502 (N_3502,N_2443,N_2307);
or U3503 (N_3503,N_2225,N_2457);
nand U3504 (N_3504,N_2428,N_2929);
nor U3505 (N_3505,N_2102,N_2244);
nor U3506 (N_3506,N_2058,N_2107);
nand U3507 (N_3507,N_2003,N_2493);
and U3508 (N_3508,N_2717,N_2894);
or U3509 (N_3509,N_2380,N_2362);
nor U3510 (N_3510,N_2474,N_2576);
nand U3511 (N_3511,N_2148,N_2584);
nor U3512 (N_3512,N_2727,N_2522);
and U3513 (N_3513,N_2564,N_2537);
or U3514 (N_3514,N_2084,N_2188);
nor U3515 (N_3515,N_2176,N_2436);
nor U3516 (N_3516,N_2132,N_2731);
nor U3517 (N_3517,N_2603,N_2855);
nand U3518 (N_3518,N_2727,N_2965);
or U3519 (N_3519,N_2261,N_2254);
nand U3520 (N_3520,N_2586,N_2279);
or U3521 (N_3521,N_2071,N_2063);
nand U3522 (N_3522,N_2991,N_2343);
nor U3523 (N_3523,N_2196,N_2441);
or U3524 (N_3524,N_2356,N_2949);
nand U3525 (N_3525,N_2070,N_2274);
and U3526 (N_3526,N_2849,N_2123);
nand U3527 (N_3527,N_2321,N_2743);
nor U3528 (N_3528,N_2555,N_2338);
or U3529 (N_3529,N_2567,N_2860);
nor U3530 (N_3530,N_2411,N_2916);
nand U3531 (N_3531,N_2801,N_2043);
nor U3532 (N_3532,N_2219,N_2689);
and U3533 (N_3533,N_2110,N_2910);
and U3534 (N_3534,N_2345,N_2402);
nor U3535 (N_3535,N_2688,N_2864);
and U3536 (N_3536,N_2764,N_2760);
and U3537 (N_3537,N_2372,N_2229);
and U3538 (N_3538,N_2354,N_2816);
nand U3539 (N_3539,N_2058,N_2020);
or U3540 (N_3540,N_2688,N_2556);
or U3541 (N_3541,N_2981,N_2013);
or U3542 (N_3542,N_2758,N_2813);
nor U3543 (N_3543,N_2589,N_2289);
and U3544 (N_3544,N_2920,N_2629);
nand U3545 (N_3545,N_2792,N_2677);
nand U3546 (N_3546,N_2365,N_2882);
and U3547 (N_3547,N_2319,N_2664);
nand U3548 (N_3548,N_2481,N_2290);
nand U3549 (N_3549,N_2157,N_2604);
and U3550 (N_3550,N_2500,N_2133);
nand U3551 (N_3551,N_2138,N_2443);
and U3552 (N_3552,N_2697,N_2906);
and U3553 (N_3553,N_2807,N_2092);
or U3554 (N_3554,N_2844,N_2658);
and U3555 (N_3555,N_2488,N_2612);
nand U3556 (N_3556,N_2491,N_2664);
nor U3557 (N_3557,N_2710,N_2734);
nand U3558 (N_3558,N_2453,N_2001);
or U3559 (N_3559,N_2586,N_2564);
or U3560 (N_3560,N_2335,N_2020);
nand U3561 (N_3561,N_2684,N_2023);
or U3562 (N_3562,N_2877,N_2308);
nor U3563 (N_3563,N_2110,N_2633);
nand U3564 (N_3564,N_2005,N_2919);
or U3565 (N_3565,N_2080,N_2333);
and U3566 (N_3566,N_2349,N_2563);
and U3567 (N_3567,N_2859,N_2445);
nor U3568 (N_3568,N_2065,N_2564);
nand U3569 (N_3569,N_2769,N_2678);
nand U3570 (N_3570,N_2950,N_2915);
nand U3571 (N_3571,N_2136,N_2091);
nand U3572 (N_3572,N_2690,N_2695);
nand U3573 (N_3573,N_2313,N_2861);
nor U3574 (N_3574,N_2758,N_2080);
nand U3575 (N_3575,N_2829,N_2422);
and U3576 (N_3576,N_2176,N_2288);
or U3577 (N_3577,N_2280,N_2922);
nor U3578 (N_3578,N_2679,N_2688);
nor U3579 (N_3579,N_2055,N_2838);
or U3580 (N_3580,N_2972,N_2722);
nand U3581 (N_3581,N_2373,N_2041);
nor U3582 (N_3582,N_2581,N_2016);
nand U3583 (N_3583,N_2007,N_2635);
nand U3584 (N_3584,N_2767,N_2101);
and U3585 (N_3585,N_2793,N_2909);
or U3586 (N_3586,N_2368,N_2117);
nor U3587 (N_3587,N_2660,N_2240);
nand U3588 (N_3588,N_2703,N_2203);
and U3589 (N_3589,N_2085,N_2498);
nor U3590 (N_3590,N_2936,N_2815);
nand U3591 (N_3591,N_2722,N_2046);
or U3592 (N_3592,N_2112,N_2917);
and U3593 (N_3593,N_2583,N_2861);
nand U3594 (N_3594,N_2297,N_2561);
and U3595 (N_3595,N_2712,N_2087);
xnor U3596 (N_3596,N_2325,N_2710);
and U3597 (N_3597,N_2036,N_2048);
nand U3598 (N_3598,N_2310,N_2048);
or U3599 (N_3599,N_2894,N_2865);
nand U3600 (N_3600,N_2063,N_2238);
and U3601 (N_3601,N_2638,N_2672);
xor U3602 (N_3602,N_2843,N_2323);
nand U3603 (N_3603,N_2512,N_2503);
and U3604 (N_3604,N_2196,N_2115);
and U3605 (N_3605,N_2166,N_2176);
nor U3606 (N_3606,N_2301,N_2012);
nor U3607 (N_3607,N_2349,N_2234);
and U3608 (N_3608,N_2135,N_2872);
and U3609 (N_3609,N_2757,N_2560);
and U3610 (N_3610,N_2076,N_2569);
and U3611 (N_3611,N_2737,N_2609);
or U3612 (N_3612,N_2733,N_2219);
and U3613 (N_3613,N_2057,N_2125);
or U3614 (N_3614,N_2048,N_2806);
and U3615 (N_3615,N_2164,N_2574);
or U3616 (N_3616,N_2794,N_2380);
nor U3617 (N_3617,N_2814,N_2346);
and U3618 (N_3618,N_2717,N_2427);
or U3619 (N_3619,N_2041,N_2673);
nand U3620 (N_3620,N_2029,N_2585);
nor U3621 (N_3621,N_2288,N_2202);
nor U3622 (N_3622,N_2095,N_2842);
nand U3623 (N_3623,N_2104,N_2825);
nand U3624 (N_3624,N_2870,N_2749);
nand U3625 (N_3625,N_2788,N_2748);
nand U3626 (N_3626,N_2897,N_2973);
nor U3627 (N_3627,N_2374,N_2032);
nor U3628 (N_3628,N_2099,N_2790);
or U3629 (N_3629,N_2810,N_2411);
nor U3630 (N_3630,N_2179,N_2135);
or U3631 (N_3631,N_2798,N_2528);
and U3632 (N_3632,N_2502,N_2511);
and U3633 (N_3633,N_2994,N_2903);
xor U3634 (N_3634,N_2724,N_2523);
and U3635 (N_3635,N_2590,N_2705);
and U3636 (N_3636,N_2846,N_2524);
nand U3637 (N_3637,N_2253,N_2314);
nand U3638 (N_3638,N_2728,N_2125);
or U3639 (N_3639,N_2229,N_2664);
or U3640 (N_3640,N_2791,N_2223);
or U3641 (N_3641,N_2674,N_2144);
or U3642 (N_3642,N_2287,N_2817);
xor U3643 (N_3643,N_2987,N_2310);
xor U3644 (N_3644,N_2543,N_2380);
or U3645 (N_3645,N_2367,N_2628);
and U3646 (N_3646,N_2416,N_2425);
or U3647 (N_3647,N_2191,N_2212);
or U3648 (N_3648,N_2356,N_2323);
nor U3649 (N_3649,N_2794,N_2616);
nand U3650 (N_3650,N_2703,N_2484);
nand U3651 (N_3651,N_2396,N_2717);
and U3652 (N_3652,N_2536,N_2578);
nor U3653 (N_3653,N_2239,N_2152);
nor U3654 (N_3654,N_2081,N_2480);
or U3655 (N_3655,N_2587,N_2346);
or U3656 (N_3656,N_2051,N_2125);
or U3657 (N_3657,N_2132,N_2916);
nor U3658 (N_3658,N_2536,N_2543);
and U3659 (N_3659,N_2987,N_2323);
or U3660 (N_3660,N_2619,N_2628);
nor U3661 (N_3661,N_2936,N_2382);
or U3662 (N_3662,N_2462,N_2723);
and U3663 (N_3663,N_2673,N_2354);
nand U3664 (N_3664,N_2175,N_2263);
xnor U3665 (N_3665,N_2519,N_2711);
nand U3666 (N_3666,N_2522,N_2038);
nand U3667 (N_3667,N_2650,N_2310);
nor U3668 (N_3668,N_2186,N_2826);
or U3669 (N_3669,N_2601,N_2750);
and U3670 (N_3670,N_2837,N_2706);
or U3671 (N_3671,N_2436,N_2029);
nand U3672 (N_3672,N_2427,N_2750);
or U3673 (N_3673,N_2356,N_2843);
nand U3674 (N_3674,N_2356,N_2854);
and U3675 (N_3675,N_2126,N_2471);
nand U3676 (N_3676,N_2957,N_2545);
nand U3677 (N_3677,N_2940,N_2502);
nand U3678 (N_3678,N_2105,N_2859);
and U3679 (N_3679,N_2288,N_2274);
nand U3680 (N_3680,N_2755,N_2641);
and U3681 (N_3681,N_2221,N_2387);
nor U3682 (N_3682,N_2591,N_2483);
nor U3683 (N_3683,N_2352,N_2785);
and U3684 (N_3684,N_2072,N_2779);
nand U3685 (N_3685,N_2333,N_2918);
xor U3686 (N_3686,N_2227,N_2939);
nor U3687 (N_3687,N_2285,N_2513);
and U3688 (N_3688,N_2613,N_2171);
nor U3689 (N_3689,N_2470,N_2909);
nor U3690 (N_3690,N_2650,N_2357);
or U3691 (N_3691,N_2345,N_2800);
and U3692 (N_3692,N_2340,N_2277);
or U3693 (N_3693,N_2903,N_2019);
and U3694 (N_3694,N_2139,N_2639);
nor U3695 (N_3695,N_2412,N_2005);
nor U3696 (N_3696,N_2820,N_2351);
or U3697 (N_3697,N_2687,N_2413);
or U3698 (N_3698,N_2901,N_2984);
nand U3699 (N_3699,N_2488,N_2181);
nand U3700 (N_3700,N_2690,N_2777);
nor U3701 (N_3701,N_2919,N_2147);
or U3702 (N_3702,N_2608,N_2179);
and U3703 (N_3703,N_2513,N_2700);
xor U3704 (N_3704,N_2418,N_2112);
nand U3705 (N_3705,N_2002,N_2415);
or U3706 (N_3706,N_2610,N_2581);
and U3707 (N_3707,N_2026,N_2446);
nand U3708 (N_3708,N_2591,N_2047);
or U3709 (N_3709,N_2724,N_2372);
nand U3710 (N_3710,N_2733,N_2040);
nand U3711 (N_3711,N_2427,N_2040);
nand U3712 (N_3712,N_2248,N_2426);
nor U3713 (N_3713,N_2774,N_2974);
and U3714 (N_3714,N_2290,N_2980);
or U3715 (N_3715,N_2082,N_2468);
and U3716 (N_3716,N_2203,N_2233);
nor U3717 (N_3717,N_2034,N_2888);
nor U3718 (N_3718,N_2881,N_2637);
nor U3719 (N_3719,N_2732,N_2416);
nand U3720 (N_3720,N_2832,N_2444);
xor U3721 (N_3721,N_2376,N_2457);
or U3722 (N_3722,N_2343,N_2631);
and U3723 (N_3723,N_2803,N_2495);
nand U3724 (N_3724,N_2989,N_2672);
nor U3725 (N_3725,N_2953,N_2654);
and U3726 (N_3726,N_2789,N_2488);
and U3727 (N_3727,N_2358,N_2727);
and U3728 (N_3728,N_2056,N_2741);
nand U3729 (N_3729,N_2545,N_2316);
or U3730 (N_3730,N_2203,N_2491);
and U3731 (N_3731,N_2656,N_2320);
and U3732 (N_3732,N_2619,N_2320);
nand U3733 (N_3733,N_2532,N_2137);
nor U3734 (N_3734,N_2349,N_2628);
and U3735 (N_3735,N_2285,N_2999);
nand U3736 (N_3736,N_2685,N_2035);
nor U3737 (N_3737,N_2668,N_2278);
or U3738 (N_3738,N_2908,N_2377);
and U3739 (N_3739,N_2605,N_2359);
and U3740 (N_3740,N_2121,N_2714);
or U3741 (N_3741,N_2169,N_2901);
and U3742 (N_3742,N_2940,N_2203);
and U3743 (N_3743,N_2046,N_2979);
nor U3744 (N_3744,N_2538,N_2086);
nand U3745 (N_3745,N_2042,N_2587);
and U3746 (N_3746,N_2797,N_2679);
nand U3747 (N_3747,N_2702,N_2643);
nor U3748 (N_3748,N_2816,N_2796);
and U3749 (N_3749,N_2297,N_2787);
and U3750 (N_3750,N_2164,N_2180);
nor U3751 (N_3751,N_2430,N_2013);
xnor U3752 (N_3752,N_2334,N_2911);
and U3753 (N_3753,N_2716,N_2871);
and U3754 (N_3754,N_2620,N_2965);
nand U3755 (N_3755,N_2470,N_2760);
nor U3756 (N_3756,N_2403,N_2728);
nor U3757 (N_3757,N_2181,N_2411);
nand U3758 (N_3758,N_2717,N_2498);
or U3759 (N_3759,N_2611,N_2864);
nor U3760 (N_3760,N_2143,N_2492);
nor U3761 (N_3761,N_2089,N_2091);
nor U3762 (N_3762,N_2105,N_2655);
nor U3763 (N_3763,N_2558,N_2036);
and U3764 (N_3764,N_2941,N_2616);
nor U3765 (N_3765,N_2618,N_2451);
nand U3766 (N_3766,N_2498,N_2935);
and U3767 (N_3767,N_2567,N_2475);
or U3768 (N_3768,N_2141,N_2401);
nand U3769 (N_3769,N_2787,N_2453);
nor U3770 (N_3770,N_2676,N_2590);
and U3771 (N_3771,N_2470,N_2902);
nor U3772 (N_3772,N_2127,N_2431);
nor U3773 (N_3773,N_2030,N_2259);
or U3774 (N_3774,N_2569,N_2493);
nor U3775 (N_3775,N_2406,N_2423);
and U3776 (N_3776,N_2416,N_2097);
nor U3777 (N_3777,N_2835,N_2356);
nor U3778 (N_3778,N_2777,N_2781);
and U3779 (N_3779,N_2602,N_2404);
or U3780 (N_3780,N_2998,N_2366);
and U3781 (N_3781,N_2966,N_2405);
and U3782 (N_3782,N_2272,N_2640);
xor U3783 (N_3783,N_2452,N_2778);
or U3784 (N_3784,N_2133,N_2586);
nor U3785 (N_3785,N_2228,N_2969);
nand U3786 (N_3786,N_2024,N_2003);
nand U3787 (N_3787,N_2694,N_2527);
xor U3788 (N_3788,N_2201,N_2742);
and U3789 (N_3789,N_2146,N_2943);
and U3790 (N_3790,N_2847,N_2727);
or U3791 (N_3791,N_2979,N_2628);
and U3792 (N_3792,N_2679,N_2196);
xnor U3793 (N_3793,N_2202,N_2652);
nor U3794 (N_3794,N_2024,N_2749);
nor U3795 (N_3795,N_2299,N_2133);
or U3796 (N_3796,N_2278,N_2136);
or U3797 (N_3797,N_2196,N_2022);
nand U3798 (N_3798,N_2958,N_2888);
and U3799 (N_3799,N_2570,N_2496);
or U3800 (N_3800,N_2826,N_2997);
and U3801 (N_3801,N_2740,N_2805);
nand U3802 (N_3802,N_2025,N_2303);
or U3803 (N_3803,N_2698,N_2363);
nand U3804 (N_3804,N_2128,N_2746);
nor U3805 (N_3805,N_2000,N_2287);
nand U3806 (N_3806,N_2376,N_2145);
nand U3807 (N_3807,N_2523,N_2595);
nor U3808 (N_3808,N_2547,N_2088);
and U3809 (N_3809,N_2617,N_2559);
nand U3810 (N_3810,N_2919,N_2329);
nor U3811 (N_3811,N_2472,N_2595);
nand U3812 (N_3812,N_2728,N_2193);
nor U3813 (N_3813,N_2567,N_2522);
nand U3814 (N_3814,N_2687,N_2608);
or U3815 (N_3815,N_2304,N_2898);
nor U3816 (N_3816,N_2464,N_2294);
nand U3817 (N_3817,N_2108,N_2747);
or U3818 (N_3818,N_2015,N_2444);
nor U3819 (N_3819,N_2199,N_2866);
nand U3820 (N_3820,N_2745,N_2957);
or U3821 (N_3821,N_2694,N_2400);
or U3822 (N_3822,N_2208,N_2813);
nand U3823 (N_3823,N_2273,N_2859);
nand U3824 (N_3824,N_2849,N_2071);
or U3825 (N_3825,N_2172,N_2246);
nand U3826 (N_3826,N_2121,N_2946);
or U3827 (N_3827,N_2555,N_2289);
or U3828 (N_3828,N_2196,N_2776);
nor U3829 (N_3829,N_2279,N_2879);
or U3830 (N_3830,N_2683,N_2918);
nor U3831 (N_3831,N_2673,N_2470);
and U3832 (N_3832,N_2807,N_2759);
nor U3833 (N_3833,N_2571,N_2130);
or U3834 (N_3834,N_2945,N_2210);
and U3835 (N_3835,N_2555,N_2281);
or U3836 (N_3836,N_2995,N_2359);
nand U3837 (N_3837,N_2403,N_2099);
and U3838 (N_3838,N_2707,N_2551);
nand U3839 (N_3839,N_2103,N_2941);
nor U3840 (N_3840,N_2359,N_2969);
or U3841 (N_3841,N_2947,N_2705);
and U3842 (N_3842,N_2155,N_2475);
or U3843 (N_3843,N_2782,N_2572);
nand U3844 (N_3844,N_2636,N_2072);
and U3845 (N_3845,N_2249,N_2919);
or U3846 (N_3846,N_2092,N_2789);
or U3847 (N_3847,N_2007,N_2201);
nand U3848 (N_3848,N_2766,N_2810);
nor U3849 (N_3849,N_2900,N_2686);
nor U3850 (N_3850,N_2027,N_2494);
nand U3851 (N_3851,N_2684,N_2327);
nor U3852 (N_3852,N_2566,N_2504);
nand U3853 (N_3853,N_2055,N_2242);
or U3854 (N_3854,N_2758,N_2997);
or U3855 (N_3855,N_2498,N_2695);
or U3856 (N_3856,N_2724,N_2530);
nor U3857 (N_3857,N_2293,N_2296);
or U3858 (N_3858,N_2983,N_2382);
or U3859 (N_3859,N_2880,N_2836);
xnor U3860 (N_3860,N_2065,N_2615);
nor U3861 (N_3861,N_2628,N_2872);
nand U3862 (N_3862,N_2071,N_2445);
nand U3863 (N_3863,N_2633,N_2621);
nor U3864 (N_3864,N_2989,N_2542);
and U3865 (N_3865,N_2026,N_2898);
and U3866 (N_3866,N_2789,N_2297);
nand U3867 (N_3867,N_2248,N_2419);
or U3868 (N_3868,N_2113,N_2407);
nor U3869 (N_3869,N_2320,N_2463);
and U3870 (N_3870,N_2381,N_2569);
nor U3871 (N_3871,N_2968,N_2756);
or U3872 (N_3872,N_2162,N_2953);
nor U3873 (N_3873,N_2869,N_2123);
and U3874 (N_3874,N_2284,N_2542);
nand U3875 (N_3875,N_2504,N_2267);
nor U3876 (N_3876,N_2627,N_2468);
nor U3877 (N_3877,N_2322,N_2702);
nor U3878 (N_3878,N_2142,N_2537);
nand U3879 (N_3879,N_2850,N_2422);
or U3880 (N_3880,N_2748,N_2309);
or U3881 (N_3881,N_2265,N_2021);
nand U3882 (N_3882,N_2968,N_2272);
nand U3883 (N_3883,N_2348,N_2789);
or U3884 (N_3884,N_2911,N_2280);
nor U3885 (N_3885,N_2864,N_2158);
nor U3886 (N_3886,N_2306,N_2855);
nor U3887 (N_3887,N_2309,N_2317);
nand U3888 (N_3888,N_2109,N_2578);
and U3889 (N_3889,N_2924,N_2041);
nor U3890 (N_3890,N_2403,N_2082);
or U3891 (N_3891,N_2585,N_2721);
nor U3892 (N_3892,N_2486,N_2749);
or U3893 (N_3893,N_2085,N_2901);
or U3894 (N_3894,N_2536,N_2561);
nor U3895 (N_3895,N_2611,N_2743);
and U3896 (N_3896,N_2569,N_2829);
or U3897 (N_3897,N_2628,N_2017);
nor U3898 (N_3898,N_2884,N_2795);
or U3899 (N_3899,N_2459,N_2655);
nand U3900 (N_3900,N_2523,N_2941);
and U3901 (N_3901,N_2207,N_2403);
nand U3902 (N_3902,N_2008,N_2491);
nor U3903 (N_3903,N_2064,N_2560);
xor U3904 (N_3904,N_2456,N_2727);
or U3905 (N_3905,N_2389,N_2496);
nor U3906 (N_3906,N_2709,N_2896);
nor U3907 (N_3907,N_2146,N_2714);
or U3908 (N_3908,N_2035,N_2101);
xnor U3909 (N_3909,N_2905,N_2346);
nor U3910 (N_3910,N_2441,N_2545);
nand U3911 (N_3911,N_2550,N_2649);
and U3912 (N_3912,N_2480,N_2117);
nor U3913 (N_3913,N_2391,N_2153);
and U3914 (N_3914,N_2650,N_2581);
nor U3915 (N_3915,N_2759,N_2618);
nand U3916 (N_3916,N_2032,N_2291);
nor U3917 (N_3917,N_2721,N_2523);
nor U3918 (N_3918,N_2960,N_2398);
and U3919 (N_3919,N_2341,N_2796);
or U3920 (N_3920,N_2207,N_2328);
and U3921 (N_3921,N_2984,N_2526);
and U3922 (N_3922,N_2545,N_2765);
and U3923 (N_3923,N_2970,N_2128);
nor U3924 (N_3924,N_2457,N_2783);
and U3925 (N_3925,N_2485,N_2059);
and U3926 (N_3926,N_2628,N_2041);
and U3927 (N_3927,N_2861,N_2169);
or U3928 (N_3928,N_2918,N_2201);
nor U3929 (N_3929,N_2202,N_2074);
nand U3930 (N_3930,N_2016,N_2026);
nand U3931 (N_3931,N_2882,N_2061);
and U3932 (N_3932,N_2734,N_2513);
nor U3933 (N_3933,N_2585,N_2901);
nand U3934 (N_3934,N_2061,N_2229);
or U3935 (N_3935,N_2097,N_2746);
xor U3936 (N_3936,N_2943,N_2427);
and U3937 (N_3937,N_2335,N_2700);
nor U3938 (N_3938,N_2032,N_2528);
nor U3939 (N_3939,N_2630,N_2573);
or U3940 (N_3940,N_2805,N_2191);
and U3941 (N_3941,N_2137,N_2406);
nor U3942 (N_3942,N_2571,N_2905);
nor U3943 (N_3943,N_2273,N_2048);
and U3944 (N_3944,N_2255,N_2098);
nor U3945 (N_3945,N_2166,N_2292);
and U3946 (N_3946,N_2491,N_2253);
or U3947 (N_3947,N_2337,N_2702);
and U3948 (N_3948,N_2175,N_2480);
nand U3949 (N_3949,N_2830,N_2332);
and U3950 (N_3950,N_2646,N_2580);
nand U3951 (N_3951,N_2063,N_2590);
or U3952 (N_3952,N_2329,N_2441);
nand U3953 (N_3953,N_2271,N_2837);
and U3954 (N_3954,N_2500,N_2155);
and U3955 (N_3955,N_2211,N_2632);
nor U3956 (N_3956,N_2644,N_2545);
nor U3957 (N_3957,N_2346,N_2138);
or U3958 (N_3958,N_2077,N_2299);
and U3959 (N_3959,N_2474,N_2410);
or U3960 (N_3960,N_2643,N_2824);
and U3961 (N_3961,N_2753,N_2628);
nand U3962 (N_3962,N_2652,N_2176);
xnor U3963 (N_3963,N_2541,N_2881);
nor U3964 (N_3964,N_2528,N_2882);
nand U3965 (N_3965,N_2667,N_2991);
and U3966 (N_3966,N_2641,N_2506);
and U3967 (N_3967,N_2249,N_2761);
nand U3968 (N_3968,N_2595,N_2496);
nor U3969 (N_3969,N_2524,N_2178);
or U3970 (N_3970,N_2661,N_2003);
nand U3971 (N_3971,N_2323,N_2009);
nand U3972 (N_3972,N_2942,N_2239);
nor U3973 (N_3973,N_2445,N_2602);
or U3974 (N_3974,N_2696,N_2467);
or U3975 (N_3975,N_2190,N_2994);
or U3976 (N_3976,N_2140,N_2080);
nand U3977 (N_3977,N_2773,N_2138);
or U3978 (N_3978,N_2533,N_2342);
nor U3979 (N_3979,N_2124,N_2630);
nand U3980 (N_3980,N_2808,N_2306);
nor U3981 (N_3981,N_2082,N_2531);
nand U3982 (N_3982,N_2054,N_2462);
or U3983 (N_3983,N_2469,N_2113);
or U3984 (N_3984,N_2660,N_2532);
nand U3985 (N_3985,N_2988,N_2842);
nor U3986 (N_3986,N_2080,N_2277);
nand U3987 (N_3987,N_2127,N_2392);
nor U3988 (N_3988,N_2535,N_2736);
or U3989 (N_3989,N_2546,N_2047);
nor U3990 (N_3990,N_2967,N_2364);
nor U3991 (N_3991,N_2086,N_2883);
and U3992 (N_3992,N_2113,N_2574);
or U3993 (N_3993,N_2108,N_2540);
or U3994 (N_3994,N_2875,N_2428);
nand U3995 (N_3995,N_2631,N_2958);
nand U3996 (N_3996,N_2707,N_2247);
or U3997 (N_3997,N_2520,N_2333);
nand U3998 (N_3998,N_2083,N_2100);
and U3999 (N_3999,N_2736,N_2452);
nor U4000 (N_4000,N_3082,N_3584);
or U4001 (N_4001,N_3164,N_3068);
nor U4002 (N_4002,N_3863,N_3104);
and U4003 (N_4003,N_3828,N_3382);
and U4004 (N_4004,N_3227,N_3081);
nor U4005 (N_4005,N_3024,N_3542);
and U4006 (N_4006,N_3557,N_3942);
or U4007 (N_4007,N_3918,N_3262);
nand U4008 (N_4008,N_3532,N_3142);
or U4009 (N_4009,N_3848,N_3258);
nand U4010 (N_4010,N_3075,N_3499);
nand U4011 (N_4011,N_3716,N_3079);
or U4012 (N_4012,N_3965,N_3560);
nand U4013 (N_4013,N_3526,N_3897);
nand U4014 (N_4014,N_3673,N_3363);
and U4015 (N_4015,N_3140,N_3087);
and U4016 (N_4016,N_3598,N_3761);
nand U4017 (N_4017,N_3251,N_3369);
nor U4018 (N_4018,N_3066,N_3564);
and U4019 (N_4019,N_3127,N_3627);
or U4020 (N_4020,N_3888,N_3775);
and U4021 (N_4021,N_3026,N_3281);
and U4022 (N_4022,N_3805,N_3267);
or U4023 (N_4023,N_3120,N_3961);
and U4024 (N_4024,N_3959,N_3744);
or U4025 (N_4025,N_3602,N_3195);
and U4026 (N_4026,N_3751,N_3536);
or U4027 (N_4027,N_3869,N_3652);
nand U4028 (N_4028,N_3752,N_3852);
or U4029 (N_4029,N_3022,N_3807);
nand U4030 (N_4030,N_3137,N_3404);
nand U4031 (N_4031,N_3785,N_3015);
and U4032 (N_4032,N_3853,N_3994);
or U4033 (N_4033,N_3777,N_3397);
nor U4034 (N_4034,N_3946,N_3872);
or U4035 (N_4035,N_3097,N_3972);
nor U4036 (N_4036,N_3044,N_3829);
or U4037 (N_4037,N_3934,N_3403);
or U4038 (N_4038,N_3974,N_3571);
and U4039 (N_4039,N_3992,N_3616);
nand U4040 (N_4040,N_3979,N_3161);
nor U4041 (N_4041,N_3389,N_3481);
or U4042 (N_4042,N_3284,N_3914);
and U4043 (N_4043,N_3924,N_3008);
or U4044 (N_4044,N_3638,N_3701);
nand U4045 (N_4045,N_3130,N_3333);
and U4046 (N_4046,N_3632,N_3462);
or U4047 (N_4047,N_3117,N_3865);
or U4048 (N_4048,N_3190,N_3506);
nand U4049 (N_4049,N_3297,N_3147);
and U4050 (N_4050,N_3430,N_3029);
or U4051 (N_4051,N_3092,N_3327);
and U4052 (N_4052,N_3825,N_3471);
or U4053 (N_4053,N_3786,N_3816);
nor U4054 (N_4054,N_3017,N_3387);
nand U4055 (N_4055,N_3248,N_3574);
nor U4056 (N_4056,N_3131,N_3727);
nand U4057 (N_4057,N_3112,N_3407);
nor U4058 (N_4058,N_3183,N_3824);
and U4059 (N_4059,N_3051,N_3064);
or U4060 (N_4060,N_3344,N_3294);
or U4061 (N_4061,N_3319,N_3362);
nor U4062 (N_4062,N_3796,N_3266);
nor U4063 (N_4063,N_3189,N_3629);
nand U4064 (N_4064,N_3903,N_3108);
or U4065 (N_4065,N_3312,N_3425);
nand U4066 (N_4066,N_3156,N_3039);
or U4067 (N_4067,N_3572,N_3678);
or U4068 (N_4068,N_3640,N_3601);
or U4069 (N_4069,N_3057,N_3392);
and U4070 (N_4070,N_3717,N_3095);
xor U4071 (N_4071,N_3702,N_3093);
nor U4072 (N_4072,N_3525,N_3646);
or U4073 (N_4073,N_3551,N_3929);
and U4074 (N_4074,N_3904,N_3366);
nand U4075 (N_4075,N_3191,N_3573);
and U4076 (N_4076,N_3122,N_3106);
nor U4077 (N_4077,N_3171,N_3799);
or U4078 (N_4078,N_3792,N_3485);
or U4079 (N_4079,N_3444,N_3880);
and U4080 (N_4080,N_3845,N_3222);
nor U4081 (N_4081,N_3693,N_3207);
and U4082 (N_4082,N_3957,N_3042);
or U4083 (N_4083,N_3358,N_3614);
and U4084 (N_4084,N_3505,N_3388);
nor U4085 (N_4085,N_3976,N_3413);
nor U4086 (N_4086,N_3831,N_3107);
or U4087 (N_4087,N_3596,N_3530);
or U4088 (N_4088,N_3018,N_3758);
nor U4089 (N_4089,N_3835,N_3055);
and U4090 (N_4090,N_3232,N_3722);
or U4091 (N_4091,N_3545,N_3298);
nand U4092 (N_4092,N_3442,N_3472);
and U4093 (N_4093,N_3901,N_3375);
nand U4094 (N_4094,N_3780,N_3768);
and U4095 (N_4095,N_3591,N_3743);
or U4096 (N_4096,N_3886,N_3401);
nand U4097 (N_4097,N_3815,N_3205);
or U4098 (N_4098,N_3760,N_3228);
nand U4099 (N_4099,N_3521,N_3136);
nand U4100 (N_4100,N_3151,N_3820);
xnor U4101 (N_4101,N_3109,N_3912);
nand U4102 (N_4102,N_3309,N_3857);
or U4103 (N_4103,N_3062,N_3927);
or U4104 (N_4104,N_3502,N_3335);
nand U4105 (N_4105,N_3535,N_3479);
nand U4106 (N_4106,N_3487,N_3050);
nand U4107 (N_4107,N_3726,N_3488);
or U4108 (N_4108,N_3233,N_3797);
nor U4109 (N_4109,N_3494,N_3742);
nand U4110 (N_4110,N_3482,N_3150);
or U4111 (N_4111,N_3517,N_3184);
or U4112 (N_4112,N_3223,N_3843);
xnor U4113 (N_4113,N_3316,N_3113);
or U4114 (N_4114,N_3791,N_3416);
nor U4115 (N_4115,N_3982,N_3723);
and U4116 (N_4116,N_3453,N_3971);
and U4117 (N_4117,N_3168,N_3625);
nor U4118 (N_4118,N_3178,N_3619);
nand U4119 (N_4119,N_3774,N_3356);
and U4120 (N_4120,N_3623,N_3299);
and U4121 (N_4121,N_3840,N_3892);
nand U4122 (N_4122,N_3862,N_3450);
and U4123 (N_4123,N_3883,N_3443);
or U4124 (N_4124,N_3783,N_3320);
nor U4125 (N_4125,N_3999,N_3846);
or U4126 (N_4126,N_3214,N_3967);
nor U4127 (N_4127,N_3111,N_3659);
and U4128 (N_4128,N_3304,N_3507);
nor U4129 (N_4129,N_3653,N_3311);
and U4130 (N_4130,N_3477,N_3833);
nand U4131 (N_4131,N_3360,N_3514);
nor U4132 (N_4132,N_3578,N_3940);
or U4133 (N_4133,N_3059,N_3098);
and U4134 (N_4134,N_3036,N_3595);
nor U4135 (N_4135,N_3696,N_3370);
or U4136 (N_4136,N_3473,N_3782);
nand U4137 (N_4137,N_3361,N_3391);
nand U4138 (N_4138,N_3870,N_3812);
xnor U4139 (N_4139,N_3539,N_3615);
nor U4140 (N_4140,N_3426,N_3308);
nor U4141 (N_4141,N_3047,N_3428);
or U4142 (N_4142,N_3396,N_3588);
nand U4143 (N_4143,N_3695,N_3121);
nand U4144 (N_4144,N_3464,N_3476);
nor U4145 (N_4145,N_3516,N_3466);
and U4146 (N_4146,N_3867,N_3329);
xnor U4147 (N_4147,N_3295,N_3496);
nand U4148 (N_4148,N_3019,N_3737);
or U4149 (N_4149,N_3674,N_3963);
or U4150 (N_4150,N_3341,N_3420);
nand U4151 (N_4151,N_3322,N_3088);
or U4152 (N_4152,N_3235,N_3714);
nor U4153 (N_4153,N_3977,N_3424);
nor U4154 (N_4154,N_3665,N_3247);
nand U4155 (N_4155,N_3861,N_3409);
nor U4156 (N_4156,N_3239,N_3484);
and U4157 (N_4157,N_3923,N_3594);
and U4158 (N_4158,N_3276,N_3257);
nand U4159 (N_4159,N_3630,N_3114);
nor U4160 (N_4160,N_3949,N_3454);
or U4161 (N_4161,N_3991,N_3528);
and U4162 (N_4162,N_3345,N_3032);
xnor U4163 (N_4163,N_3084,N_3234);
nand U4164 (N_4164,N_3860,N_3342);
or U4165 (N_4165,N_3238,N_3990);
or U4166 (N_4166,N_3993,N_3328);
and U4167 (N_4167,N_3283,N_3152);
nand U4168 (N_4168,N_3633,N_3978);
xnor U4169 (N_4169,N_3670,N_3255);
or U4170 (N_4170,N_3745,N_3209);
and U4171 (N_4171,N_3446,N_3937);
or U4172 (N_4172,N_3023,N_3162);
nor U4173 (N_4173,N_3213,N_3034);
nand U4174 (N_4174,N_3944,N_3278);
nand U4175 (N_4175,N_3393,N_3667);
or U4176 (N_4176,N_3686,N_3682);
nor U4177 (N_4177,N_3445,N_3187);
or U4178 (N_4178,N_3756,N_3802);
or U4179 (N_4179,N_3984,N_3259);
or U4180 (N_4180,N_3395,N_3719);
nand U4181 (N_4181,N_3604,N_3520);
and U4182 (N_4182,N_3415,N_3608);
and U4183 (N_4183,N_3414,N_3938);
nand U4184 (N_4184,N_3793,N_3182);
or U4185 (N_4185,N_3538,N_3699);
or U4186 (N_4186,N_3568,N_3750);
nor U4187 (N_4187,N_3609,N_3202);
and U4188 (N_4188,N_3800,N_3324);
or U4189 (N_4189,N_3406,N_3885);
and U4190 (N_4190,N_3720,N_3175);
nand U4191 (N_4191,N_3011,N_3724);
and U4192 (N_4192,N_3180,N_3533);
and U4193 (N_4193,N_3738,N_3249);
and U4194 (N_4194,N_3637,N_3710);
nor U4195 (N_4195,N_3624,N_3198);
nand U4196 (N_4196,N_3170,N_3256);
and U4197 (N_4197,N_3555,N_3367);
or U4198 (N_4198,N_3922,N_3149);
or U4199 (N_4199,N_3491,N_3157);
nor U4200 (N_4200,N_3292,N_3166);
and U4201 (N_4201,N_3353,N_3123);
nand U4202 (N_4202,N_3983,N_3754);
nor U4203 (N_4203,N_3225,N_3325);
nor U4204 (N_4204,N_3374,N_3787);
nor U4205 (N_4205,N_3091,N_3436);
xnor U4206 (N_4206,N_3570,N_3958);
or U4207 (N_4207,N_3070,N_3053);
nand U4208 (N_4208,N_3250,N_3153);
nand U4209 (N_4209,N_3220,N_3005);
nand U4210 (N_4210,N_3203,N_3432);
or U4211 (N_4211,N_3734,N_3729);
or U4212 (N_4212,N_3480,N_3069);
or U4213 (N_4213,N_3048,N_3129);
or U4214 (N_4214,N_3199,N_3192);
nand U4215 (N_4215,N_3077,N_3890);
xor U4216 (N_4216,N_3989,N_3340);
or U4217 (N_4217,N_3119,N_3871);
and U4218 (N_4218,N_3321,N_3508);
nor U4219 (N_4219,N_3952,N_3931);
nand U4220 (N_4220,N_3240,N_3749);
nand U4221 (N_4221,N_3001,N_3354);
and U4222 (N_4222,N_3613,N_3125);
nor U4223 (N_4223,N_3713,N_3881);
or U4224 (N_4224,N_3478,N_3830);
nor U4225 (N_4225,N_3177,N_3384);
and U4226 (N_4226,N_3819,N_3817);
nor U4227 (N_4227,N_3731,N_3925);
nand U4228 (N_4228,N_3173,N_3408);
nand U4229 (N_4229,N_3296,N_3575);
and U4230 (N_4230,N_3705,N_3894);
nand U4231 (N_4231,N_3617,N_3146);
or U4232 (N_4232,N_3083,N_3417);
or U4233 (N_4233,N_3589,N_3201);
nand U4234 (N_4234,N_3306,N_3216);
nand U4235 (N_4235,N_3736,N_3000);
or U4236 (N_4236,N_3174,N_3995);
nor U4237 (N_4237,N_3429,N_3467);
or U4238 (N_4238,N_3567,N_3941);
nor U4239 (N_4239,N_3926,N_3154);
or U4240 (N_4240,N_3801,N_3987);
xor U4241 (N_4241,N_3461,N_3621);
or U4242 (N_4242,N_3933,N_3103);
or U4243 (N_4243,N_3460,N_3663);
or U4244 (N_4244,N_3126,N_3025);
nand U4245 (N_4245,N_3463,N_3854);
or U4246 (N_4246,N_3597,N_3563);
and U4247 (N_4247,N_3732,N_3725);
nor U4248 (N_4248,N_3757,N_3014);
and U4249 (N_4249,N_3307,N_3317);
and U4250 (N_4250,N_3269,N_3020);
or U4251 (N_4251,N_3030,N_3287);
or U4252 (N_4252,N_3285,N_3910);
and U4253 (N_4253,N_3735,N_3855);
and U4254 (N_4254,N_3357,N_3373);
nor U4255 (N_4255,N_3179,N_3962);
nor U4256 (N_4256,N_3410,N_3512);
nor U4257 (N_4257,N_3781,N_3090);
nor U4258 (N_4258,N_3145,N_3007);
or U4259 (N_4259,N_3882,N_3851);
and U4260 (N_4260,N_3676,N_3385);
and U4261 (N_4261,N_3489,N_3847);
nor U4262 (N_4262,N_3712,N_3501);
or U4263 (N_4263,N_3263,N_3898);
and U4264 (N_4264,N_3753,N_3788);
nand U4265 (N_4265,N_3224,N_3599);
or U4266 (N_4266,N_3981,N_3132);
or U4267 (N_4267,N_3116,N_3503);
nand U4268 (N_4268,N_3932,N_3708);
or U4269 (N_4269,N_3813,N_3822);
or U4270 (N_4270,N_3899,N_3764);
and U4271 (N_4271,N_3160,N_3352);
and U4272 (N_4272,N_3773,N_3035);
xnor U4273 (N_4273,N_3905,N_3540);
and U4274 (N_4274,N_3553,N_3515);
nor U4275 (N_4275,N_3649,N_3155);
nand U4276 (N_4276,N_3537,N_3080);
nand U4277 (N_4277,N_3118,N_3832);
nor U4278 (N_4278,N_3767,N_3347);
nand U4279 (N_4279,N_3778,N_3900);
or U4280 (N_4280,N_3138,N_3271);
or U4281 (N_4281,N_3916,N_3559);
nor U4282 (N_4282,N_3423,N_3094);
nor U4283 (N_4283,N_3422,N_3243);
or U4284 (N_4284,N_3628,N_3133);
and U4285 (N_4285,N_3163,N_3065);
or U4286 (N_4286,N_3074,N_3550);
nor U4287 (N_4287,N_3661,N_3226);
nand U4288 (N_4288,N_3275,N_3606);
and U4289 (N_4289,N_3336,N_3685);
nor U4290 (N_4290,N_3427,N_3704);
nor U4291 (N_4291,N_3864,N_3691);
nand U4292 (N_4292,N_3809,N_3844);
nand U4293 (N_4293,N_3330,N_3185);
and U4294 (N_4294,N_3592,N_3664);
and U4295 (N_4295,N_3197,N_3626);
or U4296 (N_4296,N_3763,N_3798);
and U4297 (N_4297,N_3451,N_3887);
and U4298 (N_4298,N_3966,N_3556);
or U4299 (N_4299,N_3264,N_3486);
nand U4300 (N_4300,N_3431,N_3762);
or U4301 (N_4301,N_3896,N_3056);
nand U4302 (N_4302,N_3215,N_3908);
and U4303 (N_4303,N_3351,N_3365);
xnor U4304 (N_4304,N_3402,N_3859);
nor U4305 (N_4305,N_3611,N_3920);
nor U4306 (N_4306,N_3364,N_3135);
nand U4307 (N_4307,N_3688,N_3245);
nor U4308 (N_4308,N_3172,N_3493);
and U4309 (N_4309,N_3622,N_3811);
nor U4310 (N_4310,N_3144,N_3343);
or U4311 (N_4311,N_3577,N_3902);
and U4312 (N_4312,N_3953,N_3804);
and U4313 (N_4313,N_3237,N_3468);
nor U4314 (N_4314,N_3043,N_3648);
nand U4315 (N_4315,N_3045,N_3288);
and U4316 (N_4316,N_3434,N_3980);
or U4317 (N_4317,N_3518,N_3086);
and U4318 (N_4318,N_3159,N_3509);
nand U4319 (N_4319,N_3740,N_3253);
and U4320 (N_4320,N_3128,N_3677);
nor U4321 (N_4321,N_3527,N_3876);
nor U4322 (N_4322,N_3437,N_3277);
or U4323 (N_4323,N_3465,N_3850);
or U4324 (N_4324,N_3511,N_3891);
nor U4325 (N_4325,N_3523,N_3378);
and U4326 (N_4326,N_3741,N_3513);
nand U4327 (N_4327,N_3348,N_3105);
nand U4328 (N_4328,N_3302,N_3755);
or U4329 (N_4329,N_3634,N_3280);
and U4330 (N_4330,N_3110,N_3519);
nand U4331 (N_4331,N_3274,N_3418);
nand U4332 (N_4332,N_3955,N_3672);
nor U4333 (N_4333,N_3221,N_3930);
nand U4334 (N_4334,N_3593,N_3359);
and U4335 (N_4335,N_3085,N_3167);
nor U4336 (N_4336,N_3658,N_3818);
nand U4337 (N_4337,N_3300,N_3866);
nand U4338 (N_4338,N_3260,N_3707);
nand U4339 (N_4339,N_3823,N_3165);
nand U4340 (N_4340,N_3656,N_3002);
nor U4341 (N_4341,N_3689,N_3548);
nand U4342 (N_4342,N_3405,N_3718);
nand U4343 (N_4343,N_3419,N_3289);
nand U4344 (N_4344,N_3371,N_3242);
nor U4345 (N_4345,N_3875,N_3784);
nand U4346 (N_4346,N_3917,N_3236);
xnor U4347 (N_4347,N_3552,N_3706);
or U4348 (N_4348,N_3618,N_3690);
nand U4349 (N_4349,N_3099,N_3579);
nand U4350 (N_4350,N_3058,N_3006);
nor U4351 (N_4351,N_3470,N_3858);
nor U4352 (N_4352,N_3033,N_3500);
or U4353 (N_4353,N_3457,N_3377);
or U4354 (N_4354,N_3889,N_3906);
or U4355 (N_4355,N_3700,N_3772);
and U4356 (N_4356,N_3169,N_3040);
nor U4357 (N_4357,N_3124,N_3698);
nand U4358 (N_4358,N_3318,N_3497);
nor U4359 (N_4359,N_3038,N_3435);
or U4360 (N_4360,N_3534,N_3586);
nor U4361 (N_4361,N_3810,N_3349);
and U4362 (N_4362,N_3469,N_3270);
and U4363 (N_4363,N_3683,N_3176);
or U4364 (N_4364,N_3948,N_3490);
and U4365 (N_4365,N_3433,N_3368);
or U4366 (N_4366,N_3394,N_3975);
nand U4367 (N_4367,N_3635,N_3438);
and U4368 (N_4368,N_3071,N_3458);
or U4369 (N_4369,N_3522,N_3096);
or U4370 (N_4370,N_3636,N_3181);
or U4371 (N_4371,N_3590,N_3049);
and U4372 (N_4372,N_3390,N_3355);
or U4373 (N_4373,N_3739,N_3669);
and U4374 (N_4374,N_3709,N_3651);
nor U4375 (N_4375,N_3746,N_3607);
nand U4376 (N_4376,N_3254,N_3655);
and U4377 (N_4377,N_3016,N_3838);
xor U4378 (N_4378,N_3076,N_3794);
nand U4379 (N_4379,N_3581,N_3246);
nand U4380 (N_4380,N_3412,N_3668);
nand U4381 (N_4381,N_3439,N_3985);
or U4382 (N_4382,N_3583,N_3013);
nor U4383 (N_4383,N_3721,N_3067);
and U4384 (N_4384,N_3346,N_3680);
nand U4385 (N_4385,N_3576,N_3562);
or U4386 (N_4386,N_3301,N_3654);
nor U4387 (N_4387,N_3675,N_3272);
and U4388 (N_4388,N_3544,N_3662);
nand U4389 (N_4389,N_3943,N_3046);
nor U4390 (N_4390,N_3186,N_3582);
and U4391 (N_4391,N_3600,N_3379);
xnor U4392 (N_4392,N_3954,N_3200);
and U4393 (N_4393,N_3028,N_3687);
nand U4394 (N_4394,N_3986,N_3078);
nor U4395 (N_4395,N_3449,N_3448);
and U4396 (N_4396,N_3970,N_3960);
nor U4397 (N_4397,N_3836,N_3265);
nor U4398 (N_4398,N_3808,N_3456);
nand U4399 (N_4399,N_3268,N_3733);
and U4400 (N_4400,N_3657,N_3947);
and U4401 (N_4401,N_3210,N_3935);
nor U4402 (N_4402,N_3334,N_3290);
or U4403 (N_4403,N_3196,N_3218);
nor U4404 (N_4404,N_3204,N_3303);
nand U4405 (N_4405,N_3305,N_3475);
nand U4406 (N_4406,N_3230,N_3660);
nor U4407 (N_4407,N_3945,N_3291);
nor U4408 (N_4408,N_3561,N_3997);
xor U4409 (N_4409,N_3968,N_3398);
nor U4410 (N_4410,N_3921,N_3459);
nor U4411 (N_4411,N_3679,N_3206);
nand U4412 (N_4412,N_3928,N_3790);
and U4413 (N_4413,N_3645,N_3073);
nor U4414 (N_4414,N_3060,N_3194);
nand U4415 (N_4415,N_3711,N_3323);
nor U4416 (N_4416,N_3770,N_3331);
nor U4417 (N_4417,N_3964,N_3728);
nand U4418 (N_4418,N_3010,N_3061);
nor U4419 (N_4419,N_3795,N_3730);
or U4420 (N_4420,N_3747,N_3337);
and U4421 (N_4421,N_3776,N_3212);
or U4422 (N_4422,N_3543,N_3605);
and U4423 (N_4423,N_3549,N_3681);
nor U4424 (N_4424,N_3694,N_3610);
and U4425 (N_4425,N_3766,N_3031);
nand U4426 (N_4426,N_3769,N_3143);
nor U4427 (N_4427,N_3231,N_3644);
nor U4428 (N_4428,N_3666,N_3834);
or U4429 (N_4429,N_3158,N_3849);
nor U4430 (N_4430,N_3547,N_3969);
nor U4431 (N_4431,N_3217,N_3447);
nand U4432 (N_4432,N_3188,N_3498);
or U4433 (N_4433,N_3376,N_3244);
nor U4434 (N_4434,N_3141,N_3495);
or U4435 (N_4435,N_3671,N_3383);
nand U4436 (N_4436,N_3771,N_3827);
xnor U4437 (N_4437,N_3102,N_3936);
nor U4438 (N_4438,N_3381,N_3803);
nand U4439 (N_4439,N_3541,N_3569);
or U4440 (N_4440,N_3874,N_3504);
nor U4441 (N_4441,N_3715,N_3372);
nand U4442 (N_4442,N_3759,N_3684);
and U4443 (N_4443,N_3492,N_3919);
nor U4444 (N_4444,N_3139,N_3839);
nor U4445 (N_4445,N_3315,N_3988);
nor U4446 (N_4446,N_3452,N_3440);
nand U4447 (N_4447,N_3814,N_3286);
nand U4448 (N_4448,N_3293,N_3421);
or U4449 (N_4449,N_3211,N_3524);
and U4450 (N_4450,N_3338,N_3063);
nor U4451 (N_4451,N_3765,N_3585);
or U4452 (N_4452,N_3241,N_3620);
or U4453 (N_4453,N_3208,N_3907);
nand U4454 (N_4454,N_3021,N_3821);
or U4455 (N_4455,N_3950,N_3339);
or U4456 (N_4456,N_3193,N_3603);
nor U4457 (N_4457,N_3261,N_3350);
nand U4458 (N_4458,N_3273,N_3411);
nand U4459 (N_4459,N_3399,N_3998);
nor U4460 (N_4460,N_3779,N_3400);
nand U4461 (N_4461,N_3806,N_3054);
nor U4462 (N_4462,N_3893,N_3529);
or U4463 (N_4463,N_3219,N_3612);
nand U4464 (N_4464,N_3027,N_3546);
nor U4465 (N_4465,N_3554,N_3641);
or U4466 (N_4466,N_3282,N_3279);
or U4467 (N_4467,N_3326,N_3332);
and U4468 (N_4468,N_3837,N_3386);
nor U4469 (N_4469,N_3915,N_3483);
and U4470 (N_4470,N_3868,N_3842);
and U4471 (N_4471,N_3692,N_3939);
or U4472 (N_4472,N_3134,N_3229);
or U4473 (N_4473,N_3650,N_3089);
or U4474 (N_4474,N_3996,N_3115);
or U4475 (N_4475,N_3558,N_3531);
nand U4476 (N_4476,N_3041,N_3911);
nand U4477 (N_4477,N_3009,N_3703);
xnor U4478 (N_4478,N_3100,N_3313);
or U4479 (N_4479,N_3631,N_3884);
or U4480 (N_4480,N_3580,N_3973);
or U4481 (N_4481,N_3913,N_3587);
nand U4482 (N_4482,N_3380,N_3951);
nand U4483 (N_4483,N_3639,N_3441);
or U4484 (N_4484,N_3566,N_3643);
or U4485 (N_4485,N_3003,N_3841);
nand U4486 (N_4486,N_3856,N_3878);
and U4487 (N_4487,N_3909,N_3877);
xor U4488 (N_4488,N_3148,N_3101);
or U4489 (N_4489,N_3642,N_3310);
or U4490 (N_4490,N_3879,N_3873);
nor U4491 (N_4491,N_3826,N_3072);
and U4492 (N_4492,N_3510,N_3037);
or U4493 (N_4493,N_3895,N_3474);
nor U4494 (N_4494,N_3314,N_3697);
nor U4495 (N_4495,N_3252,N_3565);
nand U4496 (N_4496,N_3012,N_3956);
and U4497 (N_4497,N_3647,N_3052);
or U4498 (N_4498,N_3789,N_3455);
and U4499 (N_4499,N_3748,N_3004);
or U4500 (N_4500,N_3976,N_3626);
nand U4501 (N_4501,N_3147,N_3285);
nand U4502 (N_4502,N_3024,N_3089);
nor U4503 (N_4503,N_3775,N_3577);
and U4504 (N_4504,N_3142,N_3389);
or U4505 (N_4505,N_3984,N_3095);
nor U4506 (N_4506,N_3521,N_3441);
nand U4507 (N_4507,N_3806,N_3837);
or U4508 (N_4508,N_3346,N_3517);
nand U4509 (N_4509,N_3226,N_3394);
nand U4510 (N_4510,N_3703,N_3019);
or U4511 (N_4511,N_3049,N_3810);
or U4512 (N_4512,N_3729,N_3977);
xor U4513 (N_4513,N_3215,N_3108);
nand U4514 (N_4514,N_3729,N_3573);
nand U4515 (N_4515,N_3803,N_3048);
and U4516 (N_4516,N_3521,N_3772);
and U4517 (N_4517,N_3627,N_3738);
nor U4518 (N_4518,N_3209,N_3854);
or U4519 (N_4519,N_3712,N_3636);
xor U4520 (N_4520,N_3924,N_3142);
or U4521 (N_4521,N_3161,N_3378);
or U4522 (N_4522,N_3918,N_3395);
and U4523 (N_4523,N_3358,N_3078);
and U4524 (N_4524,N_3495,N_3839);
nand U4525 (N_4525,N_3854,N_3117);
nor U4526 (N_4526,N_3558,N_3765);
and U4527 (N_4527,N_3131,N_3262);
or U4528 (N_4528,N_3588,N_3106);
nor U4529 (N_4529,N_3459,N_3302);
xor U4530 (N_4530,N_3324,N_3933);
or U4531 (N_4531,N_3701,N_3089);
nand U4532 (N_4532,N_3387,N_3757);
and U4533 (N_4533,N_3040,N_3600);
and U4534 (N_4534,N_3598,N_3805);
or U4535 (N_4535,N_3337,N_3472);
or U4536 (N_4536,N_3778,N_3375);
nor U4537 (N_4537,N_3775,N_3349);
or U4538 (N_4538,N_3662,N_3444);
or U4539 (N_4539,N_3600,N_3586);
and U4540 (N_4540,N_3514,N_3626);
nor U4541 (N_4541,N_3892,N_3556);
nand U4542 (N_4542,N_3846,N_3490);
nor U4543 (N_4543,N_3484,N_3936);
nand U4544 (N_4544,N_3034,N_3953);
nand U4545 (N_4545,N_3069,N_3321);
nor U4546 (N_4546,N_3235,N_3319);
and U4547 (N_4547,N_3142,N_3148);
or U4548 (N_4548,N_3640,N_3566);
and U4549 (N_4549,N_3920,N_3394);
and U4550 (N_4550,N_3736,N_3453);
nand U4551 (N_4551,N_3878,N_3255);
nand U4552 (N_4552,N_3963,N_3640);
nand U4553 (N_4553,N_3534,N_3594);
nand U4554 (N_4554,N_3327,N_3276);
nor U4555 (N_4555,N_3310,N_3208);
nor U4556 (N_4556,N_3006,N_3691);
nor U4557 (N_4557,N_3458,N_3924);
nor U4558 (N_4558,N_3106,N_3892);
and U4559 (N_4559,N_3437,N_3155);
and U4560 (N_4560,N_3868,N_3584);
and U4561 (N_4561,N_3868,N_3132);
xor U4562 (N_4562,N_3666,N_3807);
and U4563 (N_4563,N_3856,N_3591);
nor U4564 (N_4564,N_3111,N_3169);
xnor U4565 (N_4565,N_3840,N_3782);
nor U4566 (N_4566,N_3859,N_3832);
nand U4567 (N_4567,N_3214,N_3577);
xor U4568 (N_4568,N_3595,N_3335);
or U4569 (N_4569,N_3483,N_3129);
nor U4570 (N_4570,N_3556,N_3814);
or U4571 (N_4571,N_3008,N_3485);
or U4572 (N_4572,N_3829,N_3924);
nand U4573 (N_4573,N_3908,N_3760);
nor U4574 (N_4574,N_3344,N_3504);
or U4575 (N_4575,N_3383,N_3535);
and U4576 (N_4576,N_3062,N_3429);
nand U4577 (N_4577,N_3659,N_3619);
nand U4578 (N_4578,N_3949,N_3737);
and U4579 (N_4579,N_3160,N_3340);
nor U4580 (N_4580,N_3051,N_3778);
or U4581 (N_4581,N_3018,N_3968);
or U4582 (N_4582,N_3842,N_3311);
and U4583 (N_4583,N_3171,N_3835);
or U4584 (N_4584,N_3414,N_3410);
nor U4585 (N_4585,N_3534,N_3577);
nor U4586 (N_4586,N_3278,N_3448);
nand U4587 (N_4587,N_3254,N_3115);
xor U4588 (N_4588,N_3388,N_3066);
nor U4589 (N_4589,N_3262,N_3052);
nand U4590 (N_4590,N_3464,N_3784);
nor U4591 (N_4591,N_3900,N_3822);
nand U4592 (N_4592,N_3383,N_3903);
nor U4593 (N_4593,N_3672,N_3614);
and U4594 (N_4594,N_3901,N_3066);
and U4595 (N_4595,N_3325,N_3816);
nand U4596 (N_4596,N_3506,N_3684);
xnor U4597 (N_4597,N_3214,N_3730);
and U4598 (N_4598,N_3981,N_3599);
and U4599 (N_4599,N_3162,N_3918);
or U4600 (N_4600,N_3681,N_3302);
nand U4601 (N_4601,N_3715,N_3862);
nor U4602 (N_4602,N_3498,N_3960);
or U4603 (N_4603,N_3311,N_3830);
nand U4604 (N_4604,N_3705,N_3580);
nand U4605 (N_4605,N_3422,N_3830);
and U4606 (N_4606,N_3495,N_3254);
nand U4607 (N_4607,N_3026,N_3804);
nor U4608 (N_4608,N_3523,N_3998);
nand U4609 (N_4609,N_3544,N_3323);
nand U4610 (N_4610,N_3724,N_3080);
or U4611 (N_4611,N_3061,N_3229);
nand U4612 (N_4612,N_3242,N_3730);
or U4613 (N_4613,N_3148,N_3392);
nand U4614 (N_4614,N_3293,N_3284);
nor U4615 (N_4615,N_3631,N_3210);
nor U4616 (N_4616,N_3239,N_3944);
or U4617 (N_4617,N_3880,N_3674);
or U4618 (N_4618,N_3891,N_3968);
and U4619 (N_4619,N_3269,N_3326);
nor U4620 (N_4620,N_3240,N_3174);
or U4621 (N_4621,N_3714,N_3656);
nand U4622 (N_4622,N_3253,N_3169);
or U4623 (N_4623,N_3929,N_3202);
nand U4624 (N_4624,N_3100,N_3232);
and U4625 (N_4625,N_3859,N_3616);
nand U4626 (N_4626,N_3525,N_3272);
nand U4627 (N_4627,N_3764,N_3802);
nor U4628 (N_4628,N_3783,N_3679);
or U4629 (N_4629,N_3886,N_3156);
nand U4630 (N_4630,N_3707,N_3182);
and U4631 (N_4631,N_3498,N_3720);
nor U4632 (N_4632,N_3419,N_3973);
nand U4633 (N_4633,N_3082,N_3674);
and U4634 (N_4634,N_3835,N_3287);
nand U4635 (N_4635,N_3420,N_3209);
nand U4636 (N_4636,N_3168,N_3194);
nand U4637 (N_4637,N_3045,N_3573);
nand U4638 (N_4638,N_3643,N_3484);
or U4639 (N_4639,N_3962,N_3682);
nand U4640 (N_4640,N_3250,N_3699);
and U4641 (N_4641,N_3744,N_3167);
or U4642 (N_4642,N_3327,N_3981);
nand U4643 (N_4643,N_3940,N_3170);
nor U4644 (N_4644,N_3607,N_3878);
and U4645 (N_4645,N_3117,N_3767);
nand U4646 (N_4646,N_3884,N_3759);
and U4647 (N_4647,N_3811,N_3411);
or U4648 (N_4648,N_3545,N_3819);
and U4649 (N_4649,N_3089,N_3375);
or U4650 (N_4650,N_3441,N_3134);
or U4651 (N_4651,N_3844,N_3089);
nor U4652 (N_4652,N_3011,N_3187);
and U4653 (N_4653,N_3287,N_3408);
and U4654 (N_4654,N_3828,N_3774);
and U4655 (N_4655,N_3662,N_3149);
nor U4656 (N_4656,N_3945,N_3264);
xnor U4657 (N_4657,N_3723,N_3565);
and U4658 (N_4658,N_3702,N_3572);
nor U4659 (N_4659,N_3255,N_3175);
and U4660 (N_4660,N_3127,N_3737);
nand U4661 (N_4661,N_3475,N_3820);
and U4662 (N_4662,N_3683,N_3380);
xnor U4663 (N_4663,N_3310,N_3341);
nand U4664 (N_4664,N_3527,N_3912);
nor U4665 (N_4665,N_3488,N_3100);
nand U4666 (N_4666,N_3519,N_3946);
nor U4667 (N_4667,N_3860,N_3421);
and U4668 (N_4668,N_3642,N_3874);
or U4669 (N_4669,N_3761,N_3544);
nor U4670 (N_4670,N_3148,N_3902);
and U4671 (N_4671,N_3546,N_3071);
and U4672 (N_4672,N_3814,N_3995);
nor U4673 (N_4673,N_3372,N_3308);
and U4674 (N_4674,N_3364,N_3889);
and U4675 (N_4675,N_3854,N_3495);
and U4676 (N_4676,N_3670,N_3323);
nor U4677 (N_4677,N_3906,N_3771);
or U4678 (N_4678,N_3369,N_3076);
and U4679 (N_4679,N_3748,N_3287);
nor U4680 (N_4680,N_3312,N_3678);
and U4681 (N_4681,N_3441,N_3956);
and U4682 (N_4682,N_3937,N_3448);
nor U4683 (N_4683,N_3862,N_3664);
nor U4684 (N_4684,N_3117,N_3798);
nor U4685 (N_4685,N_3509,N_3472);
nand U4686 (N_4686,N_3070,N_3938);
xor U4687 (N_4687,N_3485,N_3971);
or U4688 (N_4688,N_3847,N_3863);
nor U4689 (N_4689,N_3957,N_3216);
nand U4690 (N_4690,N_3079,N_3341);
nor U4691 (N_4691,N_3732,N_3184);
and U4692 (N_4692,N_3372,N_3656);
xnor U4693 (N_4693,N_3777,N_3436);
or U4694 (N_4694,N_3437,N_3125);
nand U4695 (N_4695,N_3900,N_3931);
nand U4696 (N_4696,N_3405,N_3116);
or U4697 (N_4697,N_3622,N_3000);
nand U4698 (N_4698,N_3744,N_3671);
and U4699 (N_4699,N_3227,N_3636);
and U4700 (N_4700,N_3425,N_3019);
or U4701 (N_4701,N_3927,N_3267);
or U4702 (N_4702,N_3935,N_3286);
or U4703 (N_4703,N_3312,N_3245);
nand U4704 (N_4704,N_3078,N_3329);
xnor U4705 (N_4705,N_3977,N_3726);
and U4706 (N_4706,N_3301,N_3581);
nor U4707 (N_4707,N_3136,N_3434);
and U4708 (N_4708,N_3498,N_3512);
nand U4709 (N_4709,N_3045,N_3627);
or U4710 (N_4710,N_3251,N_3259);
nor U4711 (N_4711,N_3451,N_3370);
and U4712 (N_4712,N_3323,N_3586);
or U4713 (N_4713,N_3128,N_3841);
or U4714 (N_4714,N_3711,N_3824);
or U4715 (N_4715,N_3067,N_3616);
or U4716 (N_4716,N_3374,N_3879);
nand U4717 (N_4717,N_3671,N_3422);
nor U4718 (N_4718,N_3093,N_3296);
xnor U4719 (N_4719,N_3089,N_3811);
and U4720 (N_4720,N_3805,N_3120);
and U4721 (N_4721,N_3071,N_3053);
and U4722 (N_4722,N_3601,N_3913);
nor U4723 (N_4723,N_3940,N_3030);
xnor U4724 (N_4724,N_3034,N_3158);
and U4725 (N_4725,N_3245,N_3668);
or U4726 (N_4726,N_3192,N_3550);
or U4727 (N_4727,N_3386,N_3324);
and U4728 (N_4728,N_3662,N_3884);
and U4729 (N_4729,N_3054,N_3829);
nor U4730 (N_4730,N_3130,N_3696);
nor U4731 (N_4731,N_3872,N_3856);
or U4732 (N_4732,N_3884,N_3693);
or U4733 (N_4733,N_3866,N_3325);
nand U4734 (N_4734,N_3946,N_3525);
and U4735 (N_4735,N_3864,N_3227);
or U4736 (N_4736,N_3872,N_3169);
and U4737 (N_4737,N_3559,N_3029);
nand U4738 (N_4738,N_3842,N_3956);
or U4739 (N_4739,N_3729,N_3180);
xnor U4740 (N_4740,N_3322,N_3728);
or U4741 (N_4741,N_3359,N_3996);
nand U4742 (N_4742,N_3043,N_3320);
nor U4743 (N_4743,N_3141,N_3577);
or U4744 (N_4744,N_3810,N_3859);
and U4745 (N_4745,N_3345,N_3001);
nor U4746 (N_4746,N_3040,N_3326);
or U4747 (N_4747,N_3283,N_3662);
or U4748 (N_4748,N_3453,N_3319);
nand U4749 (N_4749,N_3151,N_3482);
or U4750 (N_4750,N_3166,N_3150);
nand U4751 (N_4751,N_3221,N_3289);
or U4752 (N_4752,N_3453,N_3428);
nor U4753 (N_4753,N_3812,N_3215);
and U4754 (N_4754,N_3710,N_3514);
nand U4755 (N_4755,N_3973,N_3993);
or U4756 (N_4756,N_3599,N_3370);
and U4757 (N_4757,N_3631,N_3195);
and U4758 (N_4758,N_3254,N_3275);
nand U4759 (N_4759,N_3789,N_3308);
nor U4760 (N_4760,N_3410,N_3347);
and U4761 (N_4761,N_3748,N_3615);
xnor U4762 (N_4762,N_3118,N_3827);
nand U4763 (N_4763,N_3896,N_3538);
and U4764 (N_4764,N_3127,N_3664);
nor U4765 (N_4765,N_3550,N_3235);
nand U4766 (N_4766,N_3001,N_3051);
nand U4767 (N_4767,N_3777,N_3701);
or U4768 (N_4768,N_3126,N_3553);
and U4769 (N_4769,N_3268,N_3238);
and U4770 (N_4770,N_3545,N_3501);
nand U4771 (N_4771,N_3871,N_3003);
nand U4772 (N_4772,N_3554,N_3031);
nor U4773 (N_4773,N_3931,N_3277);
and U4774 (N_4774,N_3857,N_3139);
nand U4775 (N_4775,N_3265,N_3508);
nand U4776 (N_4776,N_3495,N_3866);
nand U4777 (N_4777,N_3444,N_3617);
nand U4778 (N_4778,N_3188,N_3949);
nand U4779 (N_4779,N_3027,N_3994);
nor U4780 (N_4780,N_3394,N_3962);
or U4781 (N_4781,N_3754,N_3151);
nor U4782 (N_4782,N_3275,N_3045);
nand U4783 (N_4783,N_3194,N_3926);
nor U4784 (N_4784,N_3903,N_3713);
and U4785 (N_4785,N_3660,N_3972);
or U4786 (N_4786,N_3583,N_3381);
nand U4787 (N_4787,N_3354,N_3049);
or U4788 (N_4788,N_3358,N_3098);
xor U4789 (N_4789,N_3771,N_3391);
nand U4790 (N_4790,N_3317,N_3103);
nor U4791 (N_4791,N_3116,N_3303);
nand U4792 (N_4792,N_3614,N_3587);
and U4793 (N_4793,N_3417,N_3318);
nand U4794 (N_4794,N_3393,N_3226);
or U4795 (N_4795,N_3410,N_3365);
and U4796 (N_4796,N_3541,N_3223);
nor U4797 (N_4797,N_3934,N_3374);
nand U4798 (N_4798,N_3949,N_3860);
nor U4799 (N_4799,N_3305,N_3783);
nand U4800 (N_4800,N_3533,N_3112);
nor U4801 (N_4801,N_3764,N_3583);
nor U4802 (N_4802,N_3726,N_3994);
or U4803 (N_4803,N_3176,N_3055);
and U4804 (N_4804,N_3046,N_3119);
nand U4805 (N_4805,N_3925,N_3716);
or U4806 (N_4806,N_3056,N_3733);
and U4807 (N_4807,N_3830,N_3903);
and U4808 (N_4808,N_3924,N_3765);
nor U4809 (N_4809,N_3148,N_3693);
xor U4810 (N_4810,N_3495,N_3361);
nand U4811 (N_4811,N_3125,N_3428);
nand U4812 (N_4812,N_3914,N_3564);
or U4813 (N_4813,N_3449,N_3350);
nor U4814 (N_4814,N_3489,N_3239);
nor U4815 (N_4815,N_3597,N_3370);
or U4816 (N_4816,N_3867,N_3761);
nor U4817 (N_4817,N_3472,N_3160);
or U4818 (N_4818,N_3125,N_3596);
nor U4819 (N_4819,N_3959,N_3593);
nor U4820 (N_4820,N_3252,N_3373);
and U4821 (N_4821,N_3183,N_3903);
nand U4822 (N_4822,N_3659,N_3497);
or U4823 (N_4823,N_3849,N_3511);
and U4824 (N_4824,N_3881,N_3927);
or U4825 (N_4825,N_3434,N_3873);
nand U4826 (N_4826,N_3874,N_3950);
nand U4827 (N_4827,N_3757,N_3949);
and U4828 (N_4828,N_3842,N_3402);
or U4829 (N_4829,N_3208,N_3618);
or U4830 (N_4830,N_3801,N_3220);
or U4831 (N_4831,N_3998,N_3728);
nor U4832 (N_4832,N_3675,N_3242);
and U4833 (N_4833,N_3473,N_3852);
or U4834 (N_4834,N_3272,N_3519);
nor U4835 (N_4835,N_3937,N_3295);
nor U4836 (N_4836,N_3854,N_3961);
nand U4837 (N_4837,N_3996,N_3132);
nor U4838 (N_4838,N_3966,N_3941);
and U4839 (N_4839,N_3832,N_3769);
nor U4840 (N_4840,N_3901,N_3948);
or U4841 (N_4841,N_3382,N_3336);
nor U4842 (N_4842,N_3168,N_3488);
nand U4843 (N_4843,N_3326,N_3840);
nand U4844 (N_4844,N_3035,N_3020);
or U4845 (N_4845,N_3179,N_3650);
nor U4846 (N_4846,N_3029,N_3903);
nand U4847 (N_4847,N_3853,N_3430);
and U4848 (N_4848,N_3716,N_3360);
nand U4849 (N_4849,N_3693,N_3322);
nor U4850 (N_4850,N_3728,N_3489);
nor U4851 (N_4851,N_3040,N_3413);
nor U4852 (N_4852,N_3317,N_3206);
nand U4853 (N_4853,N_3299,N_3132);
or U4854 (N_4854,N_3231,N_3104);
nand U4855 (N_4855,N_3826,N_3116);
and U4856 (N_4856,N_3715,N_3770);
or U4857 (N_4857,N_3489,N_3380);
and U4858 (N_4858,N_3302,N_3639);
or U4859 (N_4859,N_3864,N_3375);
and U4860 (N_4860,N_3467,N_3243);
and U4861 (N_4861,N_3200,N_3588);
and U4862 (N_4862,N_3833,N_3361);
or U4863 (N_4863,N_3399,N_3876);
nor U4864 (N_4864,N_3793,N_3531);
and U4865 (N_4865,N_3264,N_3256);
nand U4866 (N_4866,N_3532,N_3725);
nor U4867 (N_4867,N_3277,N_3920);
nand U4868 (N_4868,N_3068,N_3134);
or U4869 (N_4869,N_3617,N_3299);
nand U4870 (N_4870,N_3356,N_3756);
nand U4871 (N_4871,N_3562,N_3190);
xor U4872 (N_4872,N_3930,N_3691);
or U4873 (N_4873,N_3955,N_3059);
nor U4874 (N_4874,N_3200,N_3829);
or U4875 (N_4875,N_3500,N_3627);
nor U4876 (N_4876,N_3413,N_3082);
nand U4877 (N_4877,N_3985,N_3521);
or U4878 (N_4878,N_3716,N_3456);
nor U4879 (N_4879,N_3611,N_3941);
and U4880 (N_4880,N_3550,N_3631);
nand U4881 (N_4881,N_3666,N_3824);
and U4882 (N_4882,N_3256,N_3315);
xor U4883 (N_4883,N_3086,N_3530);
nor U4884 (N_4884,N_3927,N_3003);
and U4885 (N_4885,N_3208,N_3670);
nand U4886 (N_4886,N_3534,N_3049);
or U4887 (N_4887,N_3836,N_3413);
or U4888 (N_4888,N_3874,N_3581);
and U4889 (N_4889,N_3049,N_3393);
and U4890 (N_4890,N_3018,N_3974);
or U4891 (N_4891,N_3387,N_3806);
or U4892 (N_4892,N_3679,N_3041);
nand U4893 (N_4893,N_3601,N_3308);
nand U4894 (N_4894,N_3632,N_3322);
nor U4895 (N_4895,N_3690,N_3650);
nand U4896 (N_4896,N_3967,N_3977);
and U4897 (N_4897,N_3581,N_3519);
nor U4898 (N_4898,N_3008,N_3492);
nand U4899 (N_4899,N_3142,N_3639);
and U4900 (N_4900,N_3959,N_3675);
nor U4901 (N_4901,N_3380,N_3406);
and U4902 (N_4902,N_3579,N_3030);
nand U4903 (N_4903,N_3501,N_3176);
or U4904 (N_4904,N_3500,N_3387);
xor U4905 (N_4905,N_3495,N_3481);
nand U4906 (N_4906,N_3700,N_3809);
nand U4907 (N_4907,N_3308,N_3343);
nand U4908 (N_4908,N_3275,N_3041);
nor U4909 (N_4909,N_3924,N_3996);
or U4910 (N_4910,N_3755,N_3227);
nand U4911 (N_4911,N_3565,N_3039);
and U4912 (N_4912,N_3179,N_3374);
and U4913 (N_4913,N_3100,N_3109);
and U4914 (N_4914,N_3060,N_3197);
and U4915 (N_4915,N_3251,N_3548);
or U4916 (N_4916,N_3358,N_3010);
nor U4917 (N_4917,N_3903,N_3659);
or U4918 (N_4918,N_3224,N_3654);
nand U4919 (N_4919,N_3085,N_3155);
nor U4920 (N_4920,N_3613,N_3380);
and U4921 (N_4921,N_3298,N_3870);
and U4922 (N_4922,N_3919,N_3431);
nand U4923 (N_4923,N_3439,N_3444);
nor U4924 (N_4924,N_3959,N_3425);
or U4925 (N_4925,N_3793,N_3138);
or U4926 (N_4926,N_3612,N_3321);
xnor U4927 (N_4927,N_3991,N_3592);
nand U4928 (N_4928,N_3548,N_3303);
or U4929 (N_4929,N_3173,N_3973);
or U4930 (N_4930,N_3069,N_3986);
and U4931 (N_4931,N_3237,N_3126);
nand U4932 (N_4932,N_3411,N_3930);
nand U4933 (N_4933,N_3080,N_3341);
and U4934 (N_4934,N_3219,N_3129);
nor U4935 (N_4935,N_3142,N_3216);
nand U4936 (N_4936,N_3797,N_3582);
nor U4937 (N_4937,N_3828,N_3994);
or U4938 (N_4938,N_3596,N_3009);
nor U4939 (N_4939,N_3892,N_3510);
or U4940 (N_4940,N_3906,N_3877);
nor U4941 (N_4941,N_3660,N_3952);
nand U4942 (N_4942,N_3575,N_3862);
and U4943 (N_4943,N_3635,N_3550);
nor U4944 (N_4944,N_3000,N_3430);
or U4945 (N_4945,N_3194,N_3733);
and U4946 (N_4946,N_3388,N_3559);
nor U4947 (N_4947,N_3634,N_3737);
nor U4948 (N_4948,N_3663,N_3314);
nand U4949 (N_4949,N_3828,N_3459);
nor U4950 (N_4950,N_3949,N_3550);
or U4951 (N_4951,N_3633,N_3812);
or U4952 (N_4952,N_3154,N_3596);
and U4953 (N_4953,N_3818,N_3247);
nand U4954 (N_4954,N_3888,N_3993);
nand U4955 (N_4955,N_3550,N_3268);
xor U4956 (N_4956,N_3265,N_3540);
nor U4957 (N_4957,N_3644,N_3097);
nand U4958 (N_4958,N_3966,N_3068);
nand U4959 (N_4959,N_3294,N_3700);
or U4960 (N_4960,N_3749,N_3367);
and U4961 (N_4961,N_3772,N_3651);
nor U4962 (N_4962,N_3126,N_3886);
nand U4963 (N_4963,N_3173,N_3549);
nor U4964 (N_4964,N_3084,N_3902);
or U4965 (N_4965,N_3678,N_3894);
nor U4966 (N_4966,N_3526,N_3464);
and U4967 (N_4967,N_3496,N_3848);
or U4968 (N_4968,N_3740,N_3422);
nand U4969 (N_4969,N_3228,N_3007);
or U4970 (N_4970,N_3136,N_3781);
nand U4971 (N_4971,N_3417,N_3142);
xnor U4972 (N_4972,N_3583,N_3063);
and U4973 (N_4973,N_3188,N_3061);
nand U4974 (N_4974,N_3625,N_3869);
or U4975 (N_4975,N_3844,N_3822);
or U4976 (N_4976,N_3791,N_3213);
nor U4977 (N_4977,N_3102,N_3947);
and U4978 (N_4978,N_3276,N_3355);
nand U4979 (N_4979,N_3328,N_3583);
nor U4980 (N_4980,N_3489,N_3037);
or U4981 (N_4981,N_3446,N_3681);
nor U4982 (N_4982,N_3875,N_3793);
or U4983 (N_4983,N_3376,N_3690);
nand U4984 (N_4984,N_3316,N_3310);
nor U4985 (N_4985,N_3662,N_3741);
nor U4986 (N_4986,N_3923,N_3862);
and U4987 (N_4987,N_3002,N_3351);
nand U4988 (N_4988,N_3646,N_3627);
nand U4989 (N_4989,N_3048,N_3092);
or U4990 (N_4990,N_3548,N_3414);
and U4991 (N_4991,N_3770,N_3389);
nand U4992 (N_4992,N_3256,N_3358);
nand U4993 (N_4993,N_3950,N_3585);
nand U4994 (N_4994,N_3128,N_3035);
xor U4995 (N_4995,N_3714,N_3641);
nand U4996 (N_4996,N_3157,N_3792);
and U4997 (N_4997,N_3925,N_3759);
and U4998 (N_4998,N_3942,N_3610);
or U4999 (N_4999,N_3515,N_3654);
and UO_0 (O_0,N_4040,N_4615);
or UO_1 (O_1,N_4970,N_4343);
or UO_2 (O_2,N_4293,N_4902);
nand UO_3 (O_3,N_4377,N_4887);
nor UO_4 (O_4,N_4808,N_4512);
or UO_5 (O_5,N_4550,N_4637);
xor UO_6 (O_6,N_4553,N_4028);
nand UO_7 (O_7,N_4969,N_4723);
nor UO_8 (O_8,N_4500,N_4708);
or UO_9 (O_9,N_4230,N_4510);
nand UO_10 (O_10,N_4242,N_4009);
nand UO_11 (O_11,N_4146,N_4411);
and UO_12 (O_12,N_4036,N_4365);
nor UO_13 (O_13,N_4698,N_4088);
nand UO_14 (O_14,N_4720,N_4050);
nor UO_15 (O_15,N_4047,N_4699);
nor UO_16 (O_16,N_4710,N_4061);
or UO_17 (O_17,N_4484,N_4246);
nor UO_18 (O_18,N_4844,N_4697);
nor UO_19 (O_19,N_4070,N_4972);
or UO_20 (O_20,N_4630,N_4481);
nor UO_21 (O_21,N_4520,N_4645);
and UO_22 (O_22,N_4412,N_4558);
nor UO_23 (O_23,N_4296,N_4547);
nor UO_24 (O_24,N_4650,N_4864);
nor UO_25 (O_25,N_4700,N_4261);
or UO_26 (O_26,N_4252,N_4342);
and UO_27 (O_27,N_4049,N_4153);
and UO_28 (O_28,N_4718,N_4393);
or UO_29 (O_29,N_4672,N_4578);
or UO_30 (O_30,N_4865,N_4118);
or UO_31 (O_31,N_4385,N_4599);
and UO_32 (O_32,N_4874,N_4013);
and UO_33 (O_33,N_4323,N_4875);
and UO_34 (O_34,N_4920,N_4636);
and UO_35 (O_35,N_4077,N_4125);
xnor UO_36 (O_36,N_4607,N_4420);
nor UO_37 (O_37,N_4286,N_4360);
nand UO_38 (O_38,N_4499,N_4800);
and UO_39 (O_39,N_4458,N_4563);
or UO_40 (O_40,N_4670,N_4171);
or UO_41 (O_41,N_4582,N_4777);
nand UO_42 (O_42,N_4952,N_4614);
or UO_43 (O_43,N_4454,N_4932);
nor UO_44 (O_44,N_4368,N_4811);
nand UO_45 (O_45,N_4965,N_4443);
and UO_46 (O_46,N_4221,N_4735);
nand UO_47 (O_47,N_4459,N_4095);
nor UO_48 (O_48,N_4580,N_4870);
nor UO_49 (O_49,N_4325,N_4148);
nor UO_50 (O_50,N_4472,N_4364);
and UO_51 (O_51,N_4527,N_4189);
nand UO_52 (O_52,N_4593,N_4946);
or UO_53 (O_53,N_4192,N_4098);
and UO_54 (O_54,N_4428,N_4622);
or UO_55 (O_55,N_4348,N_4923);
nand UO_56 (O_56,N_4339,N_4260);
or UO_57 (O_57,N_4725,N_4626);
and UO_58 (O_58,N_4623,N_4683);
nor UO_59 (O_59,N_4618,N_4659);
or UO_60 (O_60,N_4890,N_4301);
and UO_61 (O_61,N_4244,N_4982);
or UO_62 (O_62,N_4926,N_4141);
nand UO_63 (O_63,N_4498,N_4689);
and UO_64 (O_64,N_4959,N_4138);
or UO_65 (O_65,N_4109,N_4503);
xor UO_66 (O_66,N_4702,N_4953);
or UO_67 (O_67,N_4210,N_4713);
or UO_68 (O_68,N_4265,N_4566);
nor UO_69 (O_69,N_4812,N_4737);
nand UO_70 (O_70,N_4934,N_4302);
or UO_71 (O_71,N_4247,N_4372);
and UO_72 (O_72,N_4251,N_4485);
nor UO_73 (O_73,N_4577,N_4313);
or UO_74 (O_74,N_4331,N_4541);
and UO_75 (O_75,N_4426,N_4091);
and UO_76 (O_76,N_4936,N_4943);
xor UO_77 (O_77,N_4401,N_4778);
or UO_78 (O_78,N_4204,N_4392);
nand UO_79 (O_79,N_4971,N_4815);
nor UO_80 (O_80,N_4439,N_4931);
and UO_81 (O_81,N_4271,N_4745);
nor UO_82 (O_82,N_4404,N_4722);
or UO_83 (O_83,N_4306,N_4046);
nand UO_84 (O_84,N_4966,N_4363);
or UO_85 (O_85,N_4494,N_4334);
nand UO_86 (O_86,N_4740,N_4475);
or UO_87 (O_87,N_4048,N_4522);
or UO_88 (O_88,N_4562,N_4862);
nand UO_89 (O_89,N_4387,N_4226);
xnor UO_90 (O_90,N_4609,N_4664);
and UO_91 (O_91,N_4341,N_4430);
nand UO_92 (O_92,N_4906,N_4585);
or UO_93 (O_93,N_4129,N_4976);
or UO_94 (O_94,N_4273,N_4060);
or UO_95 (O_95,N_4398,N_4985);
nand UO_96 (O_96,N_4587,N_4476);
and UO_97 (O_97,N_4792,N_4422);
and UO_98 (O_98,N_4017,N_4573);
nor UO_99 (O_99,N_4405,N_4782);
nand UO_100 (O_100,N_4933,N_4355);
and UO_101 (O_101,N_4384,N_4108);
xnor UO_102 (O_102,N_4993,N_4187);
or UO_103 (O_103,N_4871,N_4043);
and UO_104 (O_104,N_4324,N_4771);
or UO_105 (O_105,N_4660,N_4806);
nand UO_106 (O_106,N_4680,N_4513);
and UO_107 (O_107,N_4116,N_4432);
nor UO_108 (O_108,N_4287,N_4071);
nor UO_109 (O_109,N_4790,N_4904);
nor UO_110 (O_110,N_4268,N_4648);
or UO_111 (O_111,N_4408,N_4880);
or UO_112 (O_112,N_4996,N_4855);
nor UO_113 (O_113,N_4829,N_4546);
or UO_114 (O_114,N_4739,N_4606);
and UO_115 (O_115,N_4295,N_4222);
nand UO_116 (O_116,N_4554,N_4589);
nor UO_117 (O_117,N_4556,N_4386);
and UO_118 (O_118,N_4278,N_4282);
or UO_119 (O_119,N_4051,N_4724);
and UO_120 (O_120,N_4037,N_4687);
nor UO_121 (O_121,N_4575,N_4721);
nor UO_122 (O_122,N_4107,N_4243);
or UO_123 (O_123,N_4135,N_4219);
and UO_124 (O_124,N_4470,N_4004);
and UO_125 (O_125,N_4516,N_4111);
nor UO_126 (O_126,N_4941,N_4315);
or UO_127 (O_127,N_4610,N_4696);
xor UO_128 (O_128,N_4590,N_4403);
nand UO_129 (O_129,N_4717,N_4235);
or UO_130 (O_130,N_4007,N_4317);
nor UO_131 (O_131,N_4850,N_4440);
nand UO_132 (O_132,N_4072,N_4658);
and UO_133 (O_133,N_4240,N_4830);
nand UO_134 (O_134,N_4529,N_4509);
and UO_135 (O_135,N_4504,N_4781);
nor UO_136 (O_136,N_4973,N_4804);
and UO_137 (O_137,N_4845,N_4897);
or UO_138 (O_138,N_4955,N_4126);
nor UO_139 (O_139,N_4102,N_4545);
nand UO_140 (O_140,N_4258,N_4370);
and UO_141 (O_141,N_4526,N_4873);
nor UO_142 (O_142,N_4608,N_4292);
or UO_143 (O_143,N_4951,N_4842);
and UO_144 (O_144,N_4093,N_4540);
xnor UO_145 (O_145,N_4501,N_4528);
or UO_146 (O_146,N_4914,N_4813);
nand UO_147 (O_147,N_4876,N_4863);
nand UO_148 (O_148,N_4568,N_4130);
nand UO_149 (O_149,N_4011,N_4229);
nor UO_150 (O_150,N_4930,N_4935);
and UO_151 (O_151,N_4831,N_4676);
nand UO_152 (O_152,N_4827,N_4044);
xor UO_153 (O_153,N_4947,N_4677);
and UO_154 (O_154,N_4335,N_4746);
nand UO_155 (O_155,N_4802,N_4534);
nor UO_156 (O_156,N_4054,N_4445);
nand UO_157 (O_157,N_4330,N_4021);
or UO_158 (O_158,N_4714,N_4162);
nand UO_159 (O_159,N_4473,N_4086);
and UO_160 (O_160,N_4045,N_4239);
and UO_161 (O_161,N_4888,N_4869);
nand UO_162 (O_162,N_4631,N_4789);
nand UO_163 (O_163,N_4949,N_4073);
nor UO_164 (O_164,N_4068,N_4311);
nand UO_165 (O_165,N_4167,N_4020);
nand UO_166 (O_166,N_4349,N_4327);
and UO_167 (O_167,N_4787,N_4391);
and UO_168 (O_168,N_4431,N_4447);
and UO_169 (O_169,N_4469,N_4760);
nand UO_170 (O_170,N_4892,N_4390);
xnor UO_171 (O_171,N_4465,N_4764);
and UO_172 (O_172,N_4157,N_4195);
nand UO_173 (O_173,N_4267,N_4922);
nor UO_174 (O_174,N_4078,N_4921);
nand UO_175 (O_175,N_4160,N_4279);
nand UO_176 (O_176,N_4193,N_4795);
and UO_177 (O_177,N_4780,N_4127);
nor UO_178 (O_178,N_4826,N_4063);
and UO_179 (O_179,N_4927,N_4997);
or UO_180 (O_180,N_4816,N_4288);
nand UO_181 (O_181,N_4087,N_4200);
nand UO_182 (O_182,N_4438,N_4375);
nand UO_183 (O_183,N_4492,N_4304);
or UO_184 (O_184,N_4491,N_4081);
and UO_185 (O_185,N_4767,N_4706);
nand UO_186 (O_186,N_4164,N_4567);
or UO_187 (O_187,N_4053,N_4451);
and UO_188 (O_188,N_4859,N_4214);
nand UO_189 (O_189,N_4297,N_4346);
nand UO_190 (O_190,N_4264,N_4238);
nor UO_191 (O_191,N_4685,N_4537);
nor UO_192 (O_192,N_4216,N_4307);
and UO_193 (O_193,N_4332,N_4168);
and UO_194 (O_194,N_4150,N_4209);
or UO_195 (O_195,N_4885,N_4818);
and UO_196 (O_196,N_4241,N_4511);
and UO_197 (O_197,N_4784,N_4640);
or UO_198 (O_198,N_4478,N_4326);
nor UO_199 (O_199,N_4359,N_4662);
nor UO_200 (O_200,N_4877,N_4693);
nand UO_201 (O_201,N_4170,N_4211);
nor UO_202 (O_202,N_4741,N_4409);
nor UO_203 (O_203,N_4223,N_4066);
nor UO_204 (O_204,N_4480,N_4726);
and UO_205 (O_205,N_4381,N_4423);
nor UO_206 (O_206,N_4860,N_4096);
and UO_207 (O_207,N_4199,N_4684);
xor UO_208 (O_208,N_4538,N_4218);
nand UO_209 (O_209,N_4518,N_4309);
and UO_210 (O_210,N_4569,N_4205);
nand UO_211 (O_211,N_4514,N_4110);
nand UO_212 (O_212,N_4821,N_4548);
and UO_213 (O_213,N_4539,N_4035);
and UO_214 (O_214,N_4176,N_4316);
and UO_215 (O_215,N_4992,N_4245);
or UO_216 (O_216,N_4433,N_4891);
nor UO_217 (O_217,N_4136,N_4747);
and UO_218 (O_218,N_4612,N_4198);
or UO_219 (O_219,N_4291,N_4604);
or UO_220 (O_220,N_4207,N_4029);
and UO_221 (O_221,N_4103,N_4151);
and UO_222 (O_222,N_4801,N_4979);
nand UO_223 (O_223,N_4559,N_4186);
and UO_224 (O_224,N_4727,N_4889);
nor UO_225 (O_225,N_4983,N_4668);
and UO_226 (O_226,N_4506,N_4924);
or UO_227 (O_227,N_4272,N_4981);
nor UO_228 (O_228,N_4376,N_4532);
nor UO_229 (O_229,N_4446,N_4824);
nand UO_230 (O_230,N_4603,N_4768);
nand UO_231 (O_231,N_4113,N_4344);
nor UO_232 (O_232,N_4001,N_4651);
nand UO_233 (O_233,N_4259,N_4014);
nor UO_234 (O_234,N_4633,N_4990);
or UO_235 (O_235,N_4467,N_4793);
and UO_236 (O_236,N_4655,N_4803);
and UO_237 (O_237,N_4154,N_4119);
nor UO_238 (O_238,N_4595,N_4033);
nand UO_239 (O_239,N_4833,N_4641);
and UO_240 (O_240,N_4773,N_4799);
nand UO_241 (O_241,N_4228,N_4975);
or UO_242 (O_242,N_4038,N_4544);
nor UO_243 (O_243,N_4042,N_4034);
and UO_244 (O_244,N_4089,N_4517);
and UO_245 (O_245,N_4570,N_4303);
nor UO_246 (O_246,N_4715,N_4663);
and UO_247 (O_247,N_4406,N_4591);
or UO_248 (O_248,N_4611,N_4366);
or UO_249 (O_249,N_4661,N_4101);
or UO_250 (O_250,N_4435,N_4237);
nor UO_251 (O_251,N_4085,N_4234);
nor UO_252 (O_252,N_4843,N_4769);
nand UO_253 (O_253,N_4441,N_4709);
nor UO_254 (O_254,N_4958,N_4691);
nor UO_255 (O_255,N_4716,N_4300);
or UO_256 (O_256,N_4882,N_4175);
or UO_257 (O_257,N_4779,N_4620);
xnor UO_258 (O_258,N_4586,N_4531);
nand UO_259 (O_259,N_4122,N_4657);
nand UO_260 (O_260,N_4350,N_4841);
nand UO_261 (O_261,N_4883,N_4156);
or UO_262 (O_262,N_4878,N_4502);
nand UO_263 (O_263,N_4704,N_4253);
nor UO_264 (O_264,N_4820,N_4182);
nor UO_265 (O_265,N_4950,N_4188);
or UO_266 (O_266,N_4421,N_4627);
and UO_267 (O_267,N_4208,N_4576);
nor UO_268 (O_268,N_4774,N_4196);
nor UO_269 (O_269,N_4968,N_4565);
xor UO_270 (O_270,N_4786,N_4015);
and UO_271 (O_271,N_4908,N_4319);
nor UO_272 (O_272,N_4525,N_4450);
nand UO_273 (O_273,N_4916,N_4561);
or UO_274 (O_274,N_4463,N_4290);
and UO_275 (O_275,N_4628,N_4099);
nor UO_276 (O_276,N_4688,N_4999);
or UO_277 (O_277,N_4083,N_4312);
and UO_278 (O_278,N_4400,N_4356);
nor UO_279 (O_279,N_4197,N_4819);
nand UO_280 (O_280,N_4962,N_4928);
or UO_281 (O_281,N_4896,N_4314);
nand UO_282 (O_282,N_4457,N_4579);
nor UO_283 (O_283,N_4158,N_4254);
and UO_284 (O_284,N_4039,N_4329);
or UO_285 (O_285,N_4665,N_4759);
or UO_286 (O_286,N_4879,N_4468);
nor UO_287 (O_287,N_4437,N_4605);
xnor UO_288 (O_288,N_4255,N_4770);
nor UO_289 (O_289,N_4429,N_4624);
xor UO_290 (O_290,N_4551,N_4944);
nand UO_291 (O_291,N_4248,N_4763);
nor UO_292 (O_292,N_4079,N_4213);
nor UO_293 (O_293,N_4643,N_4361);
or UO_294 (O_294,N_4281,N_4191);
nor UO_295 (O_295,N_4601,N_4417);
and UO_296 (O_296,N_4388,N_4847);
nor UO_297 (O_297,N_4012,N_4675);
nand UO_298 (O_298,N_4839,N_4027);
or UO_299 (O_299,N_4909,N_4353);
nand UO_300 (O_300,N_4285,N_4497);
nand UO_301 (O_301,N_4505,N_4690);
nand UO_302 (O_302,N_4978,N_4681);
or UO_303 (O_303,N_4294,N_4711);
nor UO_304 (O_304,N_4893,N_4838);
xor UO_305 (O_305,N_4378,N_4989);
nor UO_306 (O_306,N_4915,N_4456);
and UO_307 (O_307,N_4519,N_4383);
nand UO_308 (O_308,N_4466,N_4058);
and UO_309 (O_309,N_4785,N_4694);
and UO_310 (O_310,N_4963,N_4508);
or UO_311 (O_311,N_4277,N_4772);
and UO_312 (O_312,N_4369,N_4798);
nor UO_313 (O_313,N_4132,N_4629);
or UO_314 (O_314,N_4903,N_4552);
or UO_315 (O_315,N_4600,N_4881);
nor UO_316 (O_316,N_4791,N_4427);
and UO_317 (O_317,N_4674,N_4367);
and UO_318 (O_318,N_4823,N_4318);
or UO_319 (O_319,N_4809,N_4479);
and UO_320 (O_320,N_4743,N_4455);
nor UO_321 (O_321,N_4399,N_4362);
and UO_322 (O_322,N_4765,N_4166);
nor UO_323 (O_323,N_4987,N_4067);
or UO_324 (O_324,N_4460,N_4488);
or UO_325 (O_325,N_4828,N_4337);
nand UO_326 (O_326,N_4834,N_4185);
nand UO_327 (O_327,N_4305,N_4143);
nand UO_328 (O_328,N_4080,N_4805);
or UO_329 (O_329,N_4910,N_4075);
or UO_330 (O_330,N_4733,N_4283);
nand UO_331 (O_331,N_4919,N_4002);
or UO_332 (O_332,N_4752,N_4231);
or UO_333 (O_333,N_4140,N_4671);
nand UO_334 (O_334,N_4775,N_4464);
and UO_335 (O_335,N_4825,N_4742);
nand UO_336 (O_336,N_4280,N_4835);
and UO_337 (O_337,N_4128,N_4515);
or UO_338 (O_338,N_4407,N_4382);
and UO_339 (O_339,N_4137,N_4703);
or UO_340 (O_340,N_4112,N_4986);
or UO_341 (O_341,N_4345,N_4899);
nand UO_342 (O_342,N_4617,N_4227);
or UO_343 (O_343,N_4938,N_4165);
or UO_344 (O_344,N_4434,N_4794);
and UO_345 (O_345,N_4616,N_4380);
nor UO_346 (O_346,N_4194,N_4535);
or UO_347 (O_347,N_4416,N_4052);
nor UO_348 (O_348,N_4555,N_4867);
and UO_349 (O_349,N_4172,N_4788);
or UO_350 (O_350,N_4692,N_4560);
nor UO_351 (O_351,N_4852,N_4495);
nand UO_352 (O_352,N_4588,N_4059);
or UO_353 (O_353,N_4490,N_4179);
and UO_354 (O_354,N_4647,N_4145);
nand UO_355 (O_355,N_4003,N_4964);
nand UO_356 (O_356,N_4948,N_4276);
nor UO_357 (O_357,N_4796,N_4410);
or UO_358 (O_358,N_4649,N_4738);
or UO_359 (O_359,N_4321,N_4937);
nor UO_360 (O_360,N_4415,N_4957);
or UO_361 (O_361,N_4635,N_4761);
and UO_362 (O_362,N_4462,N_4507);
and UO_363 (O_363,N_4905,N_4220);
nand UO_364 (O_364,N_4594,N_4263);
nand UO_365 (O_365,N_4065,N_4482);
nor UO_366 (O_366,N_4984,N_4667);
xnor UO_367 (O_367,N_4901,N_4977);
and UO_368 (O_368,N_4861,N_4728);
nor UO_369 (O_369,N_4489,N_4853);
and UO_370 (O_370,N_4144,N_4016);
nand UO_371 (O_371,N_4705,N_4487);
and UO_372 (O_372,N_4120,N_4666);
nor UO_373 (O_373,N_4632,N_4105);
nor UO_374 (O_374,N_4925,N_4991);
and UO_375 (O_375,N_4275,N_4719);
or UO_376 (O_376,N_4215,N_4602);
or UO_377 (O_377,N_4121,N_4756);
nand UO_378 (O_378,N_4249,N_4308);
and UO_379 (O_379,N_4269,N_4736);
nand UO_380 (O_380,N_4496,N_4621);
or UO_381 (O_381,N_4413,N_4453);
and UO_382 (O_382,N_4751,N_4217);
and UO_383 (O_383,N_4449,N_4338);
nor UO_384 (O_384,N_4596,N_4074);
nor UO_385 (O_385,N_4695,N_4858);
or UO_386 (O_386,N_4524,N_4754);
or UO_387 (O_387,N_4357,N_4006);
nor UO_388 (O_388,N_4114,N_4954);
nand UO_389 (O_389,N_4030,N_4884);
nor UO_390 (O_390,N_4340,N_4474);
and UO_391 (O_391,N_4783,N_4837);
nand UO_392 (O_392,N_4082,N_4177);
nor UO_393 (O_393,N_4100,N_4523);
and UO_394 (O_394,N_4753,N_4678);
nor UO_395 (O_395,N_4572,N_4232);
and UO_396 (O_396,N_4142,N_4533);
and UO_397 (O_397,N_4868,N_4483);
and UO_398 (O_398,N_4521,N_4270);
xnor UO_399 (O_399,N_4945,N_4486);
and UO_400 (O_400,N_4758,N_4730);
and UO_401 (O_401,N_4748,N_4419);
and UO_402 (O_402,N_4912,N_4000);
or UO_403 (O_403,N_4998,N_4159);
nand UO_404 (O_404,N_4206,N_4995);
and UO_405 (O_405,N_4549,N_4682);
or UO_406 (O_406,N_4084,N_4092);
nor UO_407 (O_407,N_4619,N_4298);
nand UO_408 (O_408,N_4994,N_4032);
nand UO_409 (O_409,N_4939,N_4250);
nand UO_410 (O_410,N_4701,N_4396);
and UO_411 (O_411,N_4583,N_4652);
nor UO_412 (O_412,N_4886,N_4822);
and UO_413 (O_413,N_4898,N_4849);
or UO_414 (O_414,N_4094,N_4056);
nand UO_415 (O_415,N_4807,N_4389);
and UO_416 (O_416,N_4322,N_4639);
or UO_417 (O_417,N_4180,N_4418);
and UO_418 (O_418,N_4351,N_4333);
nor UO_419 (O_419,N_4810,N_4203);
or UO_420 (O_420,N_4022,N_4394);
or UO_421 (O_421,N_4832,N_4018);
xnor UO_422 (O_422,N_4872,N_4673);
and UO_423 (O_423,N_4117,N_4584);
and UO_424 (O_424,N_4461,N_4106);
or UO_425 (O_425,N_4289,N_4131);
nand UO_426 (O_426,N_4425,N_4262);
nor UO_427 (O_427,N_4988,N_4266);
xnor UO_428 (O_428,N_4436,N_4707);
nand UO_429 (O_429,N_4076,N_4062);
nor UO_430 (O_430,N_4530,N_4183);
or UO_431 (O_431,N_4940,N_4477);
nand UO_432 (O_432,N_4644,N_4894);
or UO_433 (O_433,N_4642,N_4542);
nor UO_434 (O_434,N_4634,N_4956);
and UO_435 (O_435,N_4379,N_4395);
nand UO_436 (O_436,N_4900,N_4592);
or UO_437 (O_437,N_4471,N_4744);
or UO_438 (O_438,N_4762,N_4201);
nor UO_439 (O_439,N_4638,N_4625);
nand UO_440 (O_440,N_4336,N_4010);
or UO_441 (O_441,N_4797,N_4967);
nand UO_442 (O_442,N_4654,N_4749);
nor UO_443 (O_443,N_4581,N_4373);
xnor UO_444 (O_444,N_4139,N_4907);
nand UO_445 (O_445,N_4731,N_4895);
and UO_446 (O_446,N_4836,N_4233);
or UO_447 (O_447,N_4557,N_4090);
or UO_448 (O_448,N_4866,N_4854);
or UO_449 (O_449,N_4299,N_4358);
nor UO_450 (O_450,N_4817,N_4814);
or UO_451 (O_451,N_4181,N_4184);
and UO_452 (O_452,N_4848,N_4023);
nor UO_453 (O_453,N_4851,N_4202);
nor UO_454 (O_454,N_4960,N_4115);
and UO_455 (O_455,N_4911,N_4917);
nand UO_456 (O_456,N_4354,N_4152);
and UO_457 (O_457,N_4757,N_4173);
nand UO_458 (O_458,N_4147,N_4161);
and UO_459 (O_459,N_4005,N_4224);
nor UO_460 (O_460,N_4442,N_4155);
nand UO_461 (O_461,N_4124,N_4024);
nor UO_462 (O_462,N_4310,N_4913);
and UO_463 (O_463,N_4980,N_4055);
and UO_464 (O_464,N_4918,N_4444);
and UO_465 (O_465,N_4493,N_4031);
nor UO_466 (O_466,N_4846,N_4008);
nor UO_467 (O_467,N_4750,N_4571);
or UO_468 (O_468,N_4653,N_4178);
or UO_469 (O_469,N_4574,N_4840);
nand UO_470 (O_470,N_4057,N_4656);
nor UO_471 (O_471,N_4734,N_4679);
or UO_472 (O_472,N_4856,N_4274);
or UO_473 (O_473,N_4414,N_4212);
or UO_474 (O_474,N_4134,N_4766);
nor UO_475 (O_475,N_4543,N_4169);
nor UO_476 (O_476,N_4133,N_4328);
and UO_477 (O_477,N_4857,N_4104);
or UO_478 (O_478,N_4097,N_4961);
nand UO_479 (O_479,N_4402,N_4598);
nand UO_480 (O_480,N_4564,N_4712);
nand UO_481 (O_481,N_4163,N_4729);
nand UO_482 (O_482,N_4174,N_4320);
nor UO_483 (O_483,N_4597,N_4041);
or UO_484 (O_484,N_4019,N_4025);
nand UO_485 (O_485,N_4236,N_4347);
nand UO_486 (O_486,N_4397,N_4424);
and UO_487 (O_487,N_4929,N_4732);
nand UO_488 (O_488,N_4257,N_4190);
nor UO_489 (O_489,N_4776,N_4448);
nand UO_490 (O_490,N_4669,N_4284);
nand UO_491 (O_491,N_4123,N_4149);
nand UO_492 (O_492,N_4536,N_4374);
or UO_493 (O_493,N_4452,N_4064);
or UO_494 (O_494,N_4352,N_4613);
and UO_495 (O_495,N_4974,N_4686);
and UO_496 (O_496,N_4026,N_4942);
nor UO_497 (O_497,N_4069,N_4371);
nor UO_498 (O_498,N_4646,N_4256);
or UO_499 (O_499,N_4225,N_4755);
and UO_500 (O_500,N_4337,N_4703);
and UO_501 (O_501,N_4817,N_4689);
and UO_502 (O_502,N_4344,N_4985);
or UO_503 (O_503,N_4122,N_4382);
and UO_504 (O_504,N_4869,N_4078);
and UO_505 (O_505,N_4696,N_4615);
or UO_506 (O_506,N_4619,N_4415);
nand UO_507 (O_507,N_4173,N_4706);
nand UO_508 (O_508,N_4860,N_4145);
or UO_509 (O_509,N_4929,N_4820);
nand UO_510 (O_510,N_4898,N_4434);
nor UO_511 (O_511,N_4829,N_4086);
and UO_512 (O_512,N_4400,N_4276);
xnor UO_513 (O_513,N_4872,N_4568);
nor UO_514 (O_514,N_4606,N_4570);
nor UO_515 (O_515,N_4630,N_4669);
or UO_516 (O_516,N_4773,N_4190);
nor UO_517 (O_517,N_4542,N_4324);
or UO_518 (O_518,N_4076,N_4135);
nand UO_519 (O_519,N_4687,N_4312);
and UO_520 (O_520,N_4099,N_4068);
and UO_521 (O_521,N_4882,N_4422);
nand UO_522 (O_522,N_4990,N_4050);
nand UO_523 (O_523,N_4208,N_4486);
or UO_524 (O_524,N_4661,N_4173);
and UO_525 (O_525,N_4710,N_4099);
or UO_526 (O_526,N_4074,N_4252);
and UO_527 (O_527,N_4847,N_4379);
nor UO_528 (O_528,N_4665,N_4694);
nor UO_529 (O_529,N_4530,N_4665);
nand UO_530 (O_530,N_4880,N_4218);
nor UO_531 (O_531,N_4100,N_4672);
and UO_532 (O_532,N_4407,N_4594);
and UO_533 (O_533,N_4398,N_4735);
or UO_534 (O_534,N_4251,N_4533);
and UO_535 (O_535,N_4509,N_4252);
nor UO_536 (O_536,N_4150,N_4060);
nand UO_537 (O_537,N_4188,N_4463);
and UO_538 (O_538,N_4915,N_4440);
nor UO_539 (O_539,N_4354,N_4201);
nand UO_540 (O_540,N_4966,N_4250);
nor UO_541 (O_541,N_4977,N_4446);
and UO_542 (O_542,N_4111,N_4684);
or UO_543 (O_543,N_4513,N_4033);
nor UO_544 (O_544,N_4302,N_4615);
nor UO_545 (O_545,N_4715,N_4496);
or UO_546 (O_546,N_4656,N_4119);
nor UO_547 (O_547,N_4634,N_4241);
nor UO_548 (O_548,N_4948,N_4886);
and UO_549 (O_549,N_4686,N_4917);
nand UO_550 (O_550,N_4199,N_4308);
or UO_551 (O_551,N_4134,N_4439);
or UO_552 (O_552,N_4929,N_4523);
and UO_553 (O_553,N_4094,N_4510);
nor UO_554 (O_554,N_4331,N_4928);
xnor UO_555 (O_555,N_4727,N_4459);
and UO_556 (O_556,N_4304,N_4115);
nand UO_557 (O_557,N_4723,N_4059);
and UO_558 (O_558,N_4533,N_4559);
and UO_559 (O_559,N_4915,N_4627);
nand UO_560 (O_560,N_4891,N_4936);
nor UO_561 (O_561,N_4296,N_4465);
xor UO_562 (O_562,N_4827,N_4597);
nor UO_563 (O_563,N_4450,N_4527);
and UO_564 (O_564,N_4810,N_4224);
and UO_565 (O_565,N_4887,N_4767);
or UO_566 (O_566,N_4101,N_4773);
or UO_567 (O_567,N_4111,N_4453);
xnor UO_568 (O_568,N_4505,N_4538);
and UO_569 (O_569,N_4261,N_4352);
and UO_570 (O_570,N_4897,N_4123);
or UO_571 (O_571,N_4099,N_4784);
nor UO_572 (O_572,N_4501,N_4707);
or UO_573 (O_573,N_4775,N_4893);
nand UO_574 (O_574,N_4096,N_4745);
nor UO_575 (O_575,N_4706,N_4081);
and UO_576 (O_576,N_4141,N_4339);
and UO_577 (O_577,N_4288,N_4312);
nand UO_578 (O_578,N_4168,N_4577);
or UO_579 (O_579,N_4919,N_4594);
nand UO_580 (O_580,N_4812,N_4562);
nand UO_581 (O_581,N_4391,N_4993);
nand UO_582 (O_582,N_4331,N_4662);
nor UO_583 (O_583,N_4043,N_4884);
or UO_584 (O_584,N_4903,N_4784);
or UO_585 (O_585,N_4486,N_4986);
nand UO_586 (O_586,N_4678,N_4751);
and UO_587 (O_587,N_4557,N_4114);
nand UO_588 (O_588,N_4752,N_4787);
nand UO_589 (O_589,N_4695,N_4636);
and UO_590 (O_590,N_4397,N_4174);
or UO_591 (O_591,N_4418,N_4561);
nand UO_592 (O_592,N_4305,N_4231);
nand UO_593 (O_593,N_4947,N_4161);
or UO_594 (O_594,N_4181,N_4968);
nand UO_595 (O_595,N_4112,N_4852);
or UO_596 (O_596,N_4881,N_4963);
or UO_597 (O_597,N_4497,N_4045);
nor UO_598 (O_598,N_4865,N_4945);
or UO_599 (O_599,N_4177,N_4792);
or UO_600 (O_600,N_4160,N_4044);
or UO_601 (O_601,N_4200,N_4995);
nand UO_602 (O_602,N_4255,N_4765);
and UO_603 (O_603,N_4243,N_4891);
or UO_604 (O_604,N_4605,N_4091);
nor UO_605 (O_605,N_4804,N_4261);
nand UO_606 (O_606,N_4837,N_4241);
nand UO_607 (O_607,N_4021,N_4389);
nor UO_608 (O_608,N_4781,N_4672);
or UO_609 (O_609,N_4546,N_4528);
and UO_610 (O_610,N_4563,N_4515);
and UO_611 (O_611,N_4903,N_4882);
or UO_612 (O_612,N_4380,N_4561);
nand UO_613 (O_613,N_4217,N_4605);
or UO_614 (O_614,N_4526,N_4446);
nand UO_615 (O_615,N_4939,N_4297);
nand UO_616 (O_616,N_4963,N_4901);
or UO_617 (O_617,N_4200,N_4073);
and UO_618 (O_618,N_4972,N_4140);
nor UO_619 (O_619,N_4108,N_4308);
nand UO_620 (O_620,N_4894,N_4873);
and UO_621 (O_621,N_4935,N_4155);
nand UO_622 (O_622,N_4241,N_4505);
and UO_623 (O_623,N_4024,N_4383);
or UO_624 (O_624,N_4890,N_4882);
nand UO_625 (O_625,N_4885,N_4004);
and UO_626 (O_626,N_4748,N_4782);
nor UO_627 (O_627,N_4758,N_4842);
nor UO_628 (O_628,N_4181,N_4717);
xor UO_629 (O_629,N_4066,N_4528);
nor UO_630 (O_630,N_4668,N_4548);
or UO_631 (O_631,N_4794,N_4961);
and UO_632 (O_632,N_4320,N_4619);
nand UO_633 (O_633,N_4303,N_4446);
or UO_634 (O_634,N_4610,N_4379);
nor UO_635 (O_635,N_4859,N_4496);
or UO_636 (O_636,N_4922,N_4107);
nand UO_637 (O_637,N_4619,N_4072);
nand UO_638 (O_638,N_4848,N_4729);
or UO_639 (O_639,N_4789,N_4225);
and UO_640 (O_640,N_4560,N_4818);
nand UO_641 (O_641,N_4664,N_4607);
and UO_642 (O_642,N_4911,N_4243);
or UO_643 (O_643,N_4180,N_4850);
nand UO_644 (O_644,N_4416,N_4227);
and UO_645 (O_645,N_4956,N_4246);
and UO_646 (O_646,N_4599,N_4936);
and UO_647 (O_647,N_4785,N_4959);
or UO_648 (O_648,N_4815,N_4047);
nor UO_649 (O_649,N_4445,N_4189);
or UO_650 (O_650,N_4637,N_4954);
and UO_651 (O_651,N_4433,N_4967);
nand UO_652 (O_652,N_4222,N_4249);
nand UO_653 (O_653,N_4143,N_4815);
and UO_654 (O_654,N_4917,N_4523);
and UO_655 (O_655,N_4238,N_4231);
nand UO_656 (O_656,N_4412,N_4647);
nand UO_657 (O_657,N_4545,N_4155);
nand UO_658 (O_658,N_4075,N_4279);
and UO_659 (O_659,N_4835,N_4130);
nor UO_660 (O_660,N_4910,N_4904);
nor UO_661 (O_661,N_4666,N_4556);
nand UO_662 (O_662,N_4850,N_4540);
or UO_663 (O_663,N_4072,N_4818);
or UO_664 (O_664,N_4543,N_4251);
nor UO_665 (O_665,N_4563,N_4859);
and UO_666 (O_666,N_4237,N_4383);
and UO_667 (O_667,N_4432,N_4716);
or UO_668 (O_668,N_4308,N_4785);
or UO_669 (O_669,N_4212,N_4374);
nor UO_670 (O_670,N_4067,N_4671);
nor UO_671 (O_671,N_4442,N_4865);
nand UO_672 (O_672,N_4703,N_4065);
or UO_673 (O_673,N_4801,N_4547);
and UO_674 (O_674,N_4011,N_4029);
and UO_675 (O_675,N_4845,N_4665);
and UO_676 (O_676,N_4824,N_4132);
and UO_677 (O_677,N_4246,N_4296);
nor UO_678 (O_678,N_4993,N_4627);
or UO_679 (O_679,N_4880,N_4613);
or UO_680 (O_680,N_4570,N_4378);
nand UO_681 (O_681,N_4818,N_4311);
or UO_682 (O_682,N_4766,N_4747);
or UO_683 (O_683,N_4987,N_4357);
nor UO_684 (O_684,N_4078,N_4204);
and UO_685 (O_685,N_4153,N_4116);
nand UO_686 (O_686,N_4356,N_4518);
and UO_687 (O_687,N_4259,N_4499);
nor UO_688 (O_688,N_4663,N_4546);
and UO_689 (O_689,N_4325,N_4412);
or UO_690 (O_690,N_4494,N_4250);
xnor UO_691 (O_691,N_4631,N_4522);
or UO_692 (O_692,N_4616,N_4756);
and UO_693 (O_693,N_4348,N_4849);
nand UO_694 (O_694,N_4071,N_4330);
or UO_695 (O_695,N_4498,N_4670);
and UO_696 (O_696,N_4955,N_4605);
or UO_697 (O_697,N_4118,N_4668);
nor UO_698 (O_698,N_4483,N_4415);
and UO_699 (O_699,N_4319,N_4952);
or UO_700 (O_700,N_4775,N_4876);
nor UO_701 (O_701,N_4652,N_4759);
nand UO_702 (O_702,N_4500,N_4985);
or UO_703 (O_703,N_4700,N_4815);
nand UO_704 (O_704,N_4448,N_4576);
nand UO_705 (O_705,N_4950,N_4378);
nor UO_706 (O_706,N_4455,N_4827);
and UO_707 (O_707,N_4954,N_4359);
nor UO_708 (O_708,N_4841,N_4544);
and UO_709 (O_709,N_4170,N_4202);
nand UO_710 (O_710,N_4365,N_4360);
nand UO_711 (O_711,N_4549,N_4505);
and UO_712 (O_712,N_4365,N_4562);
nor UO_713 (O_713,N_4246,N_4561);
nor UO_714 (O_714,N_4390,N_4453);
and UO_715 (O_715,N_4752,N_4983);
or UO_716 (O_716,N_4100,N_4530);
and UO_717 (O_717,N_4770,N_4215);
or UO_718 (O_718,N_4232,N_4018);
or UO_719 (O_719,N_4525,N_4443);
nor UO_720 (O_720,N_4712,N_4783);
or UO_721 (O_721,N_4097,N_4195);
nand UO_722 (O_722,N_4794,N_4278);
nand UO_723 (O_723,N_4177,N_4759);
and UO_724 (O_724,N_4838,N_4494);
nand UO_725 (O_725,N_4688,N_4458);
nor UO_726 (O_726,N_4657,N_4687);
or UO_727 (O_727,N_4769,N_4399);
or UO_728 (O_728,N_4139,N_4865);
and UO_729 (O_729,N_4644,N_4330);
nor UO_730 (O_730,N_4742,N_4251);
and UO_731 (O_731,N_4135,N_4928);
or UO_732 (O_732,N_4230,N_4094);
nor UO_733 (O_733,N_4117,N_4316);
or UO_734 (O_734,N_4720,N_4078);
nand UO_735 (O_735,N_4010,N_4307);
and UO_736 (O_736,N_4967,N_4354);
and UO_737 (O_737,N_4850,N_4862);
or UO_738 (O_738,N_4131,N_4704);
nand UO_739 (O_739,N_4555,N_4442);
and UO_740 (O_740,N_4197,N_4851);
and UO_741 (O_741,N_4011,N_4848);
nor UO_742 (O_742,N_4289,N_4444);
nand UO_743 (O_743,N_4356,N_4974);
nand UO_744 (O_744,N_4596,N_4611);
nor UO_745 (O_745,N_4204,N_4005);
and UO_746 (O_746,N_4618,N_4034);
and UO_747 (O_747,N_4475,N_4800);
or UO_748 (O_748,N_4093,N_4547);
nand UO_749 (O_749,N_4391,N_4656);
nand UO_750 (O_750,N_4749,N_4033);
and UO_751 (O_751,N_4640,N_4347);
or UO_752 (O_752,N_4035,N_4438);
nand UO_753 (O_753,N_4350,N_4221);
nor UO_754 (O_754,N_4331,N_4377);
and UO_755 (O_755,N_4563,N_4297);
or UO_756 (O_756,N_4121,N_4366);
or UO_757 (O_757,N_4389,N_4289);
nand UO_758 (O_758,N_4667,N_4747);
nor UO_759 (O_759,N_4571,N_4784);
or UO_760 (O_760,N_4192,N_4002);
and UO_761 (O_761,N_4808,N_4053);
nor UO_762 (O_762,N_4040,N_4598);
nand UO_763 (O_763,N_4719,N_4749);
and UO_764 (O_764,N_4191,N_4247);
nor UO_765 (O_765,N_4893,N_4907);
nor UO_766 (O_766,N_4198,N_4201);
and UO_767 (O_767,N_4159,N_4757);
nor UO_768 (O_768,N_4035,N_4014);
nand UO_769 (O_769,N_4619,N_4673);
nor UO_770 (O_770,N_4264,N_4720);
or UO_771 (O_771,N_4285,N_4044);
and UO_772 (O_772,N_4076,N_4698);
or UO_773 (O_773,N_4520,N_4813);
and UO_774 (O_774,N_4049,N_4960);
and UO_775 (O_775,N_4556,N_4849);
or UO_776 (O_776,N_4274,N_4450);
and UO_777 (O_777,N_4781,N_4805);
and UO_778 (O_778,N_4204,N_4036);
nor UO_779 (O_779,N_4028,N_4116);
nor UO_780 (O_780,N_4855,N_4282);
or UO_781 (O_781,N_4929,N_4498);
nand UO_782 (O_782,N_4618,N_4292);
nor UO_783 (O_783,N_4238,N_4498);
and UO_784 (O_784,N_4346,N_4636);
nand UO_785 (O_785,N_4435,N_4195);
or UO_786 (O_786,N_4915,N_4295);
or UO_787 (O_787,N_4262,N_4417);
nand UO_788 (O_788,N_4562,N_4360);
nor UO_789 (O_789,N_4246,N_4679);
nor UO_790 (O_790,N_4702,N_4223);
or UO_791 (O_791,N_4936,N_4528);
nand UO_792 (O_792,N_4042,N_4585);
and UO_793 (O_793,N_4994,N_4031);
nor UO_794 (O_794,N_4641,N_4937);
or UO_795 (O_795,N_4920,N_4672);
or UO_796 (O_796,N_4178,N_4292);
nand UO_797 (O_797,N_4923,N_4839);
or UO_798 (O_798,N_4757,N_4777);
nand UO_799 (O_799,N_4116,N_4533);
and UO_800 (O_800,N_4915,N_4976);
and UO_801 (O_801,N_4403,N_4631);
and UO_802 (O_802,N_4383,N_4874);
or UO_803 (O_803,N_4171,N_4557);
nand UO_804 (O_804,N_4945,N_4844);
and UO_805 (O_805,N_4290,N_4836);
and UO_806 (O_806,N_4728,N_4286);
and UO_807 (O_807,N_4398,N_4019);
nor UO_808 (O_808,N_4636,N_4018);
nor UO_809 (O_809,N_4224,N_4420);
nand UO_810 (O_810,N_4433,N_4807);
nand UO_811 (O_811,N_4338,N_4109);
nand UO_812 (O_812,N_4704,N_4463);
or UO_813 (O_813,N_4635,N_4266);
nand UO_814 (O_814,N_4695,N_4334);
nand UO_815 (O_815,N_4911,N_4616);
nand UO_816 (O_816,N_4313,N_4402);
xnor UO_817 (O_817,N_4949,N_4929);
and UO_818 (O_818,N_4376,N_4136);
and UO_819 (O_819,N_4097,N_4711);
nand UO_820 (O_820,N_4394,N_4141);
nor UO_821 (O_821,N_4005,N_4261);
and UO_822 (O_822,N_4776,N_4660);
nor UO_823 (O_823,N_4132,N_4713);
and UO_824 (O_824,N_4906,N_4133);
nor UO_825 (O_825,N_4839,N_4650);
and UO_826 (O_826,N_4750,N_4558);
nor UO_827 (O_827,N_4412,N_4818);
nand UO_828 (O_828,N_4526,N_4935);
and UO_829 (O_829,N_4425,N_4389);
and UO_830 (O_830,N_4413,N_4756);
or UO_831 (O_831,N_4735,N_4023);
nor UO_832 (O_832,N_4325,N_4130);
nor UO_833 (O_833,N_4020,N_4073);
and UO_834 (O_834,N_4328,N_4154);
nand UO_835 (O_835,N_4984,N_4750);
xor UO_836 (O_836,N_4694,N_4137);
and UO_837 (O_837,N_4050,N_4904);
or UO_838 (O_838,N_4520,N_4421);
or UO_839 (O_839,N_4574,N_4152);
nand UO_840 (O_840,N_4202,N_4024);
or UO_841 (O_841,N_4378,N_4219);
and UO_842 (O_842,N_4099,N_4874);
nand UO_843 (O_843,N_4330,N_4520);
nor UO_844 (O_844,N_4737,N_4062);
nor UO_845 (O_845,N_4933,N_4854);
nor UO_846 (O_846,N_4527,N_4342);
nor UO_847 (O_847,N_4244,N_4991);
or UO_848 (O_848,N_4920,N_4153);
or UO_849 (O_849,N_4349,N_4250);
nor UO_850 (O_850,N_4259,N_4803);
and UO_851 (O_851,N_4498,N_4504);
nand UO_852 (O_852,N_4543,N_4333);
and UO_853 (O_853,N_4448,N_4147);
nand UO_854 (O_854,N_4465,N_4895);
and UO_855 (O_855,N_4889,N_4720);
or UO_856 (O_856,N_4147,N_4356);
nor UO_857 (O_857,N_4554,N_4385);
nor UO_858 (O_858,N_4653,N_4490);
or UO_859 (O_859,N_4438,N_4554);
or UO_860 (O_860,N_4300,N_4495);
nor UO_861 (O_861,N_4560,N_4811);
nand UO_862 (O_862,N_4696,N_4893);
or UO_863 (O_863,N_4645,N_4326);
nand UO_864 (O_864,N_4745,N_4656);
and UO_865 (O_865,N_4107,N_4499);
or UO_866 (O_866,N_4087,N_4932);
nand UO_867 (O_867,N_4364,N_4959);
nor UO_868 (O_868,N_4461,N_4258);
nand UO_869 (O_869,N_4012,N_4991);
and UO_870 (O_870,N_4705,N_4106);
nor UO_871 (O_871,N_4535,N_4861);
and UO_872 (O_872,N_4081,N_4278);
nand UO_873 (O_873,N_4701,N_4780);
nand UO_874 (O_874,N_4777,N_4262);
or UO_875 (O_875,N_4973,N_4520);
and UO_876 (O_876,N_4731,N_4673);
nor UO_877 (O_877,N_4458,N_4151);
and UO_878 (O_878,N_4175,N_4744);
or UO_879 (O_879,N_4763,N_4767);
or UO_880 (O_880,N_4624,N_4392);
and UO_881 (O_881,N_4688,N_4368);
nand UO_882 (O_882,N_4026,N_4355);
and UO_883 (O_883,N_4835,N_4890);
and UO_884 (O_884,N_4692,N_4245);
nor UO_885 (O_885,N_4214,N_4392);
or UO_886 (O_886,N_4329,N_4647);
nand UO_887 (O_887,N_4491,N_4187);
or UO_888 (O_888,N_4976,N_4100);
or UO_889 (O_889,N_4730,N_4332);
nand UO_890 (O_890,N_4355,N_4052);
or UO_891 (O_891,N_4188,N_4441);
or UO_892 (O_892,N_4467,N_4301);
nor UO_893 (O_893,N_4619,N_4896);
xor UO_894 (O_894,N_4632,N_4452);
and UO_895 (O_895,N_4118,N_4250);
and UO_896 (O_896,N_4667,N_4636);
or UO_897 (O_897,N_4230,N_4339);
or UO_898 (O_898,N_4710,N_4996);
or UO_899 (O_899,N_4595,N_4825);
nor UO_900 (O_900,N_4457,N_4791);
and UO_901 (O_901,N_4881,N_4860);
or UO_902 (O_902,N_4915,N_4222);
nand UO_903 (O_903,N_4422,N_4610);
xnor UO_904 (O_904,N_4149,N_4714);
nand UO_905 (O_905,N_4057,N_4959);
nor UO_906 (O_906,N_4915,N_4130);
or UO_907 (O_907,N_4282,N_4540);
nand UO_908 (O_908,N_4706,N_4452);
and UO_909 (O_909,N_4532,N_4324);
nor UO_910 (O_910,N_4613,N_4969);
or UO_911 (O_911,N_4541,N_4076);
or UO_912 (O_912,N_4400,N_4196);
nand UO_913 (O_913,N_4594,N_4803);
nor UO_914 (O_914,N_4646,N_4073);
nor UO_915 (O_915,N_4520,N_4260);
or UO_916 (O_916,N_4267,N_4921);
or UO_917 (O_917,N_4713,N_4202);
nor UO_918 (O_918,N_4991,N_4214);
nor UO_919 (O_919,N_4316,N_4255);
and UO_920 (O_920,N_4994,N_4212);
nor UO_921 (O_921,N_4137,N_4733);
and UO_922 (O_922,N_4412,N_4754);
nor UO_923 (O_923,N_4940,N_4606);
nand UO_924 (O_924,N_4523,N_4361);
or UO_925 (O_925,N_4647,N_4709);
nor UO_926 (O_926,N_4328,N_4943);
nand UO_927 (O_927,N_4774,N_4689);
xor UO_928 (O_928,N_4585,N_4415);
or UO_929 (O_929,N_4698,N_4301);
nand UO_930 (O_930,N_4359,N_4817);
or UO_931 (O_931,N_4214,N_4587);
and UO_932 (O_932,N_4447,N_4288);
nor UO_933 (O_933,N_4227,N_4829);
and UO_934 (O_934,N_4899,N_4544);
nor UO_935 (O_935,N_4736,N_4839);
or UO_936 (O_936,N_4701,N_4809);
nor UO_937 (O_937,N_4160,N_4798);
nor UO_938 (O_938,N_4787,N_4527);
nor UO_939 (O_939,N_4722,N_4000);
nor UO_940 (O_940,N_4376,N_4750);
nand UO_941 (O_941,N_4315,N_4365);
xor UO_942 (O_942,N_4084,N_4625);
nand UO_943 (O_943,N_4140,N_4044);
and UO_944 (O_944,N_4402,N_4700);
or UO_945 (O_945,N_4598,N_4138);
and UO_946 (O_946,N_4495,N_4039);
nor UO_947 (O_947,N_4073,N_4419);
and UO_948 (O_948,N_4963,N_4155);
nor UO_949 (O_949,N_4448,N_4322);
nor UO_950 (O_950,N_4812,N_4575);
or UO_951 (O_951,N_4243,N_4716);
and UO_952 (O_952,N_4745,N_4689);
nor UO_953 (O_953,N_4284,N_4216);
or UO_954 (O_954,N_4792,N_4265);
nor UO_955 (O_955,N_4395,N_4400);
and UO_956 (O_956,N_4593,N_4223);
nand UO_957 (O_957,N_4880,N_4453);
nand UO_958 (O_958,N_4912,N_4461);
or UO_959 (O_959,N_4804,N_4920);
nand UO_960 (O_960,N_4201,N_4462);
and UO_961 (O_961,N_4453,N_4320);
and UO_962 (O_962,N_4607,N_4088);
or UO_963 (O_963,N_4214,N_4338);
nor UO_964 (O_964,N_4443,N_4170);
nand UO_965 (O_965,N_4901,N_4778);
nor UO_966 (O_966,N_4177,N_4033);
or UO_967 (O_967,N_4651,N_4071);
nand UO_968 (O_968,N_4993,N_4645);
nand UO_969 (O_969,N_4191,N_4832);
nand UO_970 (O_970,N_4131,N_4133);
or UO_971 (O_971,N_4346,N_4854);
xnor UO_972 (O_972,N_4966,N_4057);
nand UO_973 (O_973,N_4295,N_4914);
nand UO_974 (O_974,N_4487,N_4145);
and UO_975 (O_975,N_4126,N_4491);
nor UO_976 (O_976,N_4146,N_4548);
nor UO_977 (O_977,N_4968,N_4637);
and UO_978 (O_978,N_4511,N_4606);
nand UO_979 (O_979,N_4632,N_4504);
or UO_980 (O_980,N_4172,N_4993);
and UO_981 (O_981,N_4096,N_4874);
or UO_982 (O_982,N_4717,N_4959);
and UO_983 (O_983,N_4556,N_4425);
and UO_984 (O_984,N_4706,N_4354);
and UO_985 (O_985,N_4374,N_4369);
or UO_986 (O_986,N_4936,N_4457);
and UO_987 (O_987,N_4663,N_4667);
or UO_988 (O_988,N_4142,N_4837);
nand UO_989 (O_989,N_4250,N_4645);
or UO_990 (O_990,N_4099,N_4579);
xnor UO_991 (O_991,N_4445,N_4954);
or UO_992 (O_992,N_4253,N_4931);
nand UO_993 (O_993,N_4243,N_4974);
nand UO_994 (O_994,N_4284,N_4677);
or UO_995 (O_995,N_4097,N_4601);
nor UO_996 (O_996,N_4685,N_4741);
and UO_997 (O_997,N_4630,N_4759);
and UO_998 (O_998,N_4175,N_4035);
and UO_999 (O_999,N_4164,N_4100);
endmodule