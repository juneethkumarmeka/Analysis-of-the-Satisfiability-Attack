module basic_750_5000_1000_10_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_624,In_267);
nor U1 (N_1,In_316,In_633);
nor U2 (N_2,In_742,In_606);
and U3 (N_3,In_257,In_336);
and U4 (N_4,In_740,In_48);
nor U5 (N_5,In_642,In_673);
nor U6 (N_6,In_436,In_576);
or U7 (N_7,In_17,In_268);
or U8 (N_8,In_362,In_437);
and U9 (N_9,In_583,In_253);
and U10 (N_10,In_621,In_128);
and U11 (N_11,In_631,In_489);
and U12 (N_12,In_275,In_456);
and U13 (N_13,In_557,In_52);
nand U14 (N_14,In_38,In_263);
xnor U15 (N_15,In_523,In_526);
nand U16 (N_16,In_169,In_78);
nor U17 (N_17,In_208,In_47);
and U18 (N_18,In_385,In_634);
or U19 (N_19,In_415,In_543);
nor U20 (N_20,In_508,In_668);
nand U21 (N_21,In_704,In_441);
nand U22 (N_22,In_544,In_206);
or U23 (N_23,In_195,In_708);
nor U24 (N_24,In_251,In_635);
nand U25 (N_25,In_231,In_524);
nor U26 (N_26,In_393,In_172);
or U27 (N_27,In_693,In_479);
and U28 (N_28,In_644,In_687);
nor U29 (N_29,In_111,In_61);
or U30 (N_30,In_739,In_616);
nor U31 (N_31,In_665,In_310);
nor U32 (N_32,In_395,In_112);
nand U33 (N_33,In_501,In_605);
and U34 (N_34,In_540,In_422);
or U35 (N_35,In_281,In_125);
xor U36 (N_36,In_658,In_555);
nor U37 (N_37,In_329,In_375);
and U38 (N_38,In_389,In_137);
or U39 (N_39,In_748,In_141);
and U40 (N_40,In_712,In_399);
nand U41 (N_41,In_554,In_403);
or U42 (N_42,In_553,In_718);
or U43 (N_43,In_37,In_243);
or U44 (N_44,In_659,In_235);
nor U45 (N_45,In_200,In_716);
nor U46 (N_46,In_44,In_250);
or U47 (N_47,In_204,In_438);
or U48 (N_48,In_154,In_143);
and U49 (N_49,In_379,In_130);
nand U50 (N_50,In_333,In_353);
nand U51 (N_51,In_449,In_57);
xnor U52 (N_52,In_474,In_499);
or U53 (N_53,In_7,In_63);
nand U54 (N_54,In_99,In_215);
or U55 (N_55,In_435,In_498);
or U56 (N_56,In_378,In_160);
or U57 (N_57,In_686,In_21);
nor U58 (N_58,In_105,In_535);
nor U59 (N_59,In_211,In_387);
and U60 (N_60,In_706,In_170);
xnor U61 (N_61,In_695,In_715);
nor U62 (N_62,In_68,In_346);
nand U63 (N_63,In_370,In_343);
nor U64 (N_64,In_28,In_601);
nand U65 (N_65,In_439,In_326);
and U66 (N_66,In_561,In_542);
and U67 (N_67,In_571,In_420);
and U68 (N_68,In_547,In_424);
or U69 (N_69,In_724,In_549);
or U70 (N_70,In_480,In_197);
nor U71 (N_71,In_150,In_233);
nor U72 (N_72,In_529,In_669);
and U73 (N_73,In_296,In_405);
nand U74 (N_74,In_666,In_640);
or U75 (N_75,In_124,In_131);
nand U76 (N_76,In_505,In_140);
nand U77 (N_77,In_155,In_569);
or U78 (N_78,In_737,In_183);
nand U79 (N_79,In_692,In_232);
nand U80 (N_80,In_443,In_367);
or U81 (N_81,In_303,In_174);
nand U82 (N_82,In_476,In_248);
and U83 (N_83,In_432,In_565);
or U84 (N_84,In_168,In_444);
or U85 (N_85,In_397,In_525);
nand U86 (N_86,In_51,In_638);
nor U87 (N_87,In_264,In_455);
or U88 (N_88,In_556,In_203);
nand U89 (N_89,In_110,In_34);
or U90 (N_90,In_593,In_579);
nor U91 (N_91,In_87,In_54);
and U92 (N_92,In_611,In_194);
nand U93 (N_93,In_468,In_56);
or U94 (N_94,In_539,In_163);
and U95 (N_95,In_664,In_186);
and U96 (N_96,In_361,In_573);
nor U97 (N_97,In_746,In_613);
nor U98 (N_98,In_357,In_351);
nand U99 (N_99,In_671,In_698);
nand U100 (N_100,In_500,In_300);
nand U101 (N_101,In_401,In_323);
and U102 (N_102,In_152,In_494);
or U103 (N_103,In_207,In_162);
nand U104 (N_104,In_711,In_428);
nor U105 (N_105,In_491,In_483);
nor U106 (N_106,In_373,In_591);
and U107 (N_107,In_701,In_62);
nor U108 (N_108,In_185,In_452);
xor U109 (N_109,In_83,In_356);
nor U110 (N_110,In_466,In_190);
and U111 (N_111,In_315,In_587);
and U112 (N_112,In_299,In_371);
nand U113 (N_113,In_278,In_199);
or U114 (N_114,In_222,In_426);
or U115 (N_115,In_696,In_84);
and U116 (N_116,In_702,In_509);
nand U117 (N_117,In_728,In_16);
or U118 (N_118,In_358,In_77);
or U119 (N_119,In_512,In_283);
nor U120 (N_120,In_259,In_396);
nor U121 (N_121,In_100,In_433);
nor U122 (N_122,In_503,In_91);
and U123 (N_123,In_89,In_147);
nand U124 (N_124,In_285,In_596);
and U125 (N_125,In_214,In_637);
nor U126 (N_126,In_327,In_306);
or U127 (N_127,In_372,In_74);
nand U128 (N_128,In_590,In_685);
nor U129 (N_129,In_492,In_562);
or U130 (N_130,In_42,In_679);
or U131 (N_131,In_180,In_697);
or U132 (N_132,In_691,In_18);
or U133 (N_133,In_550,In_722);
nand U134 (N_134,In_10,In_221);
or U135 (N_135,In_677,In_462);
and U136 (N_136,In_284,In_646);
nor U137 (N_137,In_50,In_309);
or U138 (N_138,In_689,In_465);
and U139 (N_139,In_442,In_682);
or U140 (N_140,In_114,In_652);
or U141 (N_141,In_240,In_481);
nor U142 (N_142,In_382,In_597);
nor U143 (N_143,In_572,In_538);
nand U144 (N_144,In_325,In_518);
nand U145 (N_145,In_398,In_626);
and U146 (N_146,In_409,In_528);
nand U147 (N_147,In_717,In_72);
nand U148 (N_148,In_317,In_408);
and U149 (N_149,In_600,In_680);
and U150 (N_150,In_651,In_617);
or U151 (N_151,In_36,In_119);
nor U152 (N_152,In_581,In_604);
or U153 (N_153,In_703,In_560);
and U154 (N_154,In_541,In_344);
nor U155 (N_155,In_400,In_135);
xor U156 (N_156,In_330,In_678);
and U157 (N_157,In_212,In_53);
or U158 (N_158,In_447,In_81);
nand U159 (N_159,In_582,In_741);
nor U160 (N_160,In_477,In_238);
and U161 (N_161,In_318,In_532);
nor U162 (N_162,In_217,In_256);
nand U163 (N_163,In_192,In_493);
or U164 (N_164,In_531,In_406);
or U165 (N_165,In_98,In_674);
or U166 (N_166,In_586,In_216);
and U167 (N_167,In_255,In_730);
nand U168 (N_168,In_577,In_165);
nand U169 (N_169,In_339,In_453);
or U170 (N_170,In_291,In_287);
or U171 (N_171,In_134,In_348);
or U172 (N_172,In_609,In_470);
nor U173 (N_173,In_608,In_429);
or U174 (N_174,In_49,In_520);
and U175 (N_175,In_460,In_311);
nand U176 (N_176,In_308,In_102);
and U177 (N_177,In_90,In_510);
or U178 (N_178,In_193,In_384);
nand U179 (N_179,In_210,In_632);
nand U180 (N_180,In_603,In_79);
nor U181 (N_181,In_589,In_101);
nand U182 (N_182,In_258,In_271);
and U183 (N_183,In_32,In_412);
or U184 (N_184,In_521,In_226);
or U185 (N_185,In_707,In_220);
nand U186 (N_186,In_104,In_684);
or U187 (N_187,In_198,In_352);
or U188 (N_188,In_534,In_46);
nor U189 (N_189,In_623,In_417);
and U190 (N_190,In_8,In_80);
or U191 (N_191,In_506,In_584);
nand U192 (N_192,In_558,In_118);
and U193 (N_193,In_239,In_502);
nand U194 (N_194,In_388,In_260);
nand U195 (N_195,In_519,In_545);
nand U196 (N_196,In_187,In_302);
or U197 (N_197,In_146,In_656);
nor U198 (N_198,In_725,In_568);
nor U199 (N_199,In_120,In_138);
nand U200 (N_200,In_566,In_218);
xor U201 (N_201,In_76,In_418);
nor U202 (N_202,In_627,In_341);
nand U203 (N_203,In_657,In_672);
nand U204 (N_204,In_106,In_450);
xnor U205 (N_205,In_368,In_288);
nand U206 (N_206,In_594,In_223);
nor U207 (N_207,In_683,In_592);
and U208 (N_208,In_133,In_35);
nor U209 (N_209,In_363,In_364);
and U210 (N_210,In_340,In_15);
nor U211 (N_211,In_485,In_289);
or U212 (N_212,In_619,In_338);
nor U213 (N_213,In_33,In_570);
and U214 (N_214,In_421,In_45);
nand U215 (N_215,In_234,In_365);
nand U216 (N_216,In_127,In_228);
and U217 (N_217,In_445,In_670);
xor U218 (N_218,In_129,In_376);
nor U219 (N_219,In_144,In_244);
and U220 (N_220,In_14,In_237);
nand U221 (N_221,In_270,In_297);
or U222 (N_222,In_73,In_515);
nor U223 (N_223,In_64,In_643);
nor U224 (N_224,In_705,In_731);
nor U225 (N_225,In_85,In_86);
nor U226 (N_226,In_490,In_459);
and U227 (N_227,In_171,In_121);
nand U228 (N_228,In_298,In_688);
or U229 (N_229,In_337,In_69);
nor U230 (N_230,In_136,In_176);
or U231 (N_231,In_334,In_20);
xnor U232 (N_232,In_205,In_551);
or U233 (N_233,In_294,In_213);
and U234 (N_234,In_369,In_265);
nand U235 (N_235,In_736,In_43);
xor U236 (N_236,In_331,In_55);
nor U237 (N_237,In_132,In_249);
nand U238 (N_238,In_486,In_552);
or U239 (N_239,In_25,In_23);
nand U240 (N_240,In_109,In_404);
and U241 (N_241,In_161,In_738);
or U242 (N_242,In_97,In_578);
and U243 (N_243,In_636,In_639);
nand U244 (N_244,In_391,In_292);
and U245 (N_245,In_290,In_495);
nand U246 (N_246,In_457,In_40);
or U247 (N_247,In_423,In_377);
nor U248 (N_248,In_332,In_522);
and U249 (N_249,In_354,In_647);
or U250 (N_250,In_546,In_747);
xor U251 (N_251,In_484,In_2);
and U252 (N_252,In_312,In_31);
nor U253 (N_253,In_575,In_178);
nor U254 (N_254,In_246,In_660);
nor U255 (N_255,In_663,In_3);
nand U256 (N_256,In_487,In_179);
or U257 (N_257,In_175,In_173);
nor U258 (N_258,In_342,In_448);
nor U259 (N_259,In_390,In_650);
nand U260 (N_260,In_4,In_286);
and U261 (N_261,In_430,In_191);
nor U262 (N_262,In_392,In_735);
and U263 (N_263,In_721,In_530);
or U264 (N_264,In_92,In_458);
or U265 (N_265,In_407,In_598);
or U266 (N_266,In_293,In_280);
or U267 (N_267,In_675,In_383);
nor U268 (N_268,In_321,In_734);
or U269 (N_269,In_236,In_66);
nand U270 (N_270,In_366,In_167);
or U271 (N_271,In_700,In_497);
nor U272 (N_272,In_75,In_641);
xor U273 (N_273,In_599,In_322);
nand U274 (N_274,In_661,In_126);
nand U275 (N_275,In_59,In_727);
or U276 (N_276,In_27,In_559);
and U277 (N_277,In_282,In_649);
and U278 (N_278,In_196,In_305);
or U279 (N_279,In_574,In_122);
or U280 (N_280,In_142,In_709);
and U281 (N_281,In_622,In_504);
and U282 (N_282,In_227,In_720);
and U283 (N_283,In_517,In_607);
nor U284 (N_284,In_602,In_60);
or U285 (N_285,In_723,In_304);
nor U286 (N_286,In_30,In_710);
or U287 (N_287,In_272,In_151);
or U288 (N_288,In_88,In_148);
nor U289 (N_289,In_247,In_9);
or U290 (N_290,In_225,In_472);
or U291 (N_291,In_714,In_24);
or U292 (N_292,In_82,In_269);
or U293 (N_293,In_694,In_419);
or U294 (N_294,In_655,In_645);
or U295 (N_295,In_473,In_380);
or U296 (N_296,In_533,In_230);
nor U297 (N_297,In_625,In_95);
nor U298 (N_298,In_413,In_116);
nor U299 (N_299,In_252,In_158);
or U300 (N_300,In_732,In_229);
and U301 (N_301,In_699,In_301);
or U302 (N_302,In_65,In_202);
nand U303 (N_303,In_482,In_359);
nor U304 (N_304,In_729,In_471);
or U305 (N_305,In_648,In_70);
nor U306 (N_306,In_690,In_653);
nor U307 (N_307,In_629,In_266);
and U308 (N_308,In_411,In_713);
and U309 (N_309,In_527,In_360);
or U310 (N_310,In_580,In_12);
nand U311 (N_311,In_307,In_745);
or U312 (N_312,In_184,In_113);
or U313 (N_313,In_676,In_274);
or U314 (N_314,In_431,In_454);
and U315 (N_315,In_743,In_262);
nand U316 (N_316,In_618,In_219);
and U317 (N_317,In_414,In_209);
and U318 (N_318,In_164,In_628);
nand U319 (N_319,In_595,In_451);
and U320 (N_320,In_277,In_328);
or U321 (N_321,In_475,In_614);
xor U322 (N_322,In_350,In_177);
nor U323 (N_323,In_564,In_145);
and U324 (N_324,In_585,In_157);
xnor U325 (N_325,In_39,In_123);
nor U326 (N_326,In_67,In_276);
or U327 (N_327,In_427,In_615);
xor U328 (N_328,In_513,In_0);
nor U329 (N_329,In_386,In_548);
nand U330 (N_330,In_115,In_347);
nand U331 (N_331,In_654,In_224);
and U332 (N_332,In_463,In_159);
nand U333 (N_333,In_567,In_719);
nand U334 (N_334,In_425,In_726);
nor U335 (N_335,In_612,In_467);
or U336 (N_336,In_261,In_13);
nand U337 (N_337,In_516,In_349);
or U338 (N_338,In_324,In_313);
or U339 (N_339,In_588,In_254);
nor U340 (N_340,In_107,In_5);
or U341 (N_341,In_749,In_96);
nor U342 (N_342,In_71,In_189);
and U343 (N_343,In_563,In_314);
nand U344 (N_344,In_153,In_488);
nor U345 (N_345,In_11,In_279);
or U346 (N_346,In_58,In_434);
and U347 (N_347,In_41,In_507);
nor U348 (N_348,In_103,In_335);
and U349 (N_349,In_667,In_345);
nand U350 (N_350,In_355,In_610);
and U351 (N_351,In_241,In_394);
and U352 (N_352,In_410,In_681);
xor U353 (N_353,In_182,In_117);
nor U354 (N_354,In_464,In_511);
or U355 (N_355,In_245,In_108);
nand U356 (N_356,In_93,In_22);
and U357 (N_357,In_242,In_374);
and U358 (N_358,In_295,In_166);
xnor U359 (N_359,In_733,In_156);
and U360 (N_360,In_537,In_620);
nor U361 (N_361,In_19,In_402);
or U362 (N_362,In_514,In_496);
nor U363 (N_363,In_536,In_201);
and U364 (N_364,In_26,In_744);
nor U365 (N_365,In_478,In_1);
nor U366 (N_366,In_188,In_469);
nor U367 (N_367,In_319,In_416);
nand U368 (N_368,In_6,In_149);
and U369 (N_369,In_94,In_139);
and U370 (N_370,In_320,In_440);
or U371 (N_371,In_181,In_446);
and U372 (N_372,In_461,In_29);
nor U373 (N_373,In_630,In_381);
and U374 (N_374,In_273,In_662);
or U375 (N_375,In_85,In_577);
and U376 (N_376,In_89,In_192);
or U377 (N_377,In_538,In_528);
or U378 (N_378,In_491,In_716);
and U379 (N_379,In_271,In_155);
and U380 (N_380,In_363,In_236);
nand U381 (N_381,In_736,In_35);
nor U382 (N_382,In_346,In_171);
nand U383 (N_383,In_317,In_370);
or U384 (N_384,In_205,In_493);
and U385 (N_385,In_267,In_56);
and U386 (N_386,In_119,In_603);
nor U387 (N_387,In_686,In_9);
or U388 (N_388,In_84,In_308);
nand U389 (N_389,In_517,In_188);
nand U390 (N_390,In_504,In_339);
and U391 (N_391,In_584,In_696);
nand U392 (N_392,In_510,In_606);
or U393 (N_393,In_341,In_210);
nor U394 (N_394,In_266,In_689);
and U395 (N_395,In_210,In_596);
xnor U396 (N_396,In_657,In_399);
nand U397 (N_397,In_265,In_440);
and U398 (N_398,In_323,In_264);
or U399 (N_399,In_408,In_102);
and U400 (N_400,In_89,In_370);
nand U401 (N_401,In_334,In_678);
nand U402 (N_402,In_687,In_500);
nor U403 (N_403,In_401,In_291);
or U404 (N_404,In_362,In_517);
nand U405 (N_405,In_293,In_502);
nor U406 (N_406,In_338,In_428);
and U407 (N_407,In_695,In_490);
nand U408 (N_408,In_311,In_572);
nand U409 (N_409,In_636,In_78);
nand U410 (N_410,In_417,In_136);
nor U411 (N_411,In_482,In_665);
nand U412 (N_412,In_542,In_356);
nor U413 (N_413,In_222,In_407);
nand U414 (N_414,In_432,In_10);
nor U415 (N_415,In_569,In_414);
or U416 (N_416,In_483,In_180);
and U417 (N_417,In_678,In_108);
and U418 (N_418,In_448,In_137);
nand U419 (N_419,In_455,In_340);
and U420 (N_420,In_663,In_535);
and U421 (N_421,In_678,In_105);
and U422 (N_422,In_532,In_159);
nor U423 (N_423,In_287,In_86);
or U424 (N_424,In_528,In_147);
nor U425 (N_425,In_82,In_425);
nand U426 (N_426,In_168,In_300);
or U427 (N_427,In_338,In_292);
and U428 (N_428,In_280,In_18);
xor U429 (N_429,In_642,In_446);
and U430 (N_430,In_628,In_163);
nand U431 (N_431,In_84,In_713);
nand U432 (N_432,In_279,In_487);
nor U433 (N_433,In_121,In_25);
nand U434 (N_434,In_560,In_206);
nand U435 (N_435,In_533,In_503);
nor U436 (N_436,In_406,In_181);
and U437 (N_437,In_625,In_562);
or U438 (N_438,In_650,In_663);
nand U439 (N_439,In_469,In_562);
nand U440 (N_440,In_245,In_698);
nor U441 (N_441,In_432,In_639);
nor U442 (N_442,In_176,In_15);
nor U443 (N_443,In_16,In_478);
xnor U444 (N_444,In_112,In_96);
nand U445 (N_445,In_368,In_439);
or U446 (N_446,In_212,In_127);
nand U447 (N_447,In_516,In_325);
nand U448 (N_448,In_435,In_436);
or U449 (N_449,In_439,In_693);
or U450 (N_450,In_215,In_448);
or U451 (N_451,In_399,In_744);
and U452 (N_452,In_553,In_112);
nor U453 (N_453,In_425,In_274);
nor U454 (N_454,In_185,In_525);
and U455 (N_455,In_648,In_348);
nand U456 (N_456,In_199,In_234);
and U457 (N_457,In_72,In_80);
and U458 (N_458,In_448,In_577);
and U459 (N_459,In_437,In_373);
nand U460 (N_460,In_111,In_566);
nor U461 (N_461,In_263,In_118);
nand U462 (N_462,In_122,In_589);
nor U463 (N_463,In_505,In_489);
nor U464 (N_464,In_463,In_200);
and U465 (N_465,In_228,In_60);
nor U466 (N_466,In_583,In_709);
and U467 (N_467,In_127,In_306);
and U468 (N_468,In_168,In_708);
nand U469 (N_469,In_103,In_220);
and U470 (N_470,In_49,In_362);
nand U471 (N_471,In_718,In_196);
and U472 (N_472,In_571,In_749);
nand U473 (N_473,In_567,In_6);
nand U474 (N_474,In_51,In_627);
and U475 (N_475,In_181,In_187);
nor U476 (N_476,In_454,In_599);
or U477 (N_477,In_160,In_264);
nor U478 (N_478,In_720,In_131);
nor U479 (N_479,In_477,In_95);
or U480 (N_480,In_540,In_157);
nor U481 (N_481,In_77,In_676);
xor U482 (N_482,In_449,In_111);
xnor U483 (N_483,In_91,In_386);
nand U484 (N_484,In_265,In_382);
nor U485 (N_485,In_565,In_740);
xor U486 (N_486,In_463,In_697);
or U487 (N_487,In_379,In_340);
and U488 (N_488,In_455,In_714);
nand U489 (N_489,In_633,In_705);
nor U490 (N_490,In_132,In_181);
nand U491 (N_491,In_255,In_454);
nor U492 (N_492,In_536,In_63);
nor U493 (N_493,In_213,In_652);
or U494 (N_494,In_254,In_359);
nor U495 (N_495,In_357,In_83);
or U496 (N_496,In_93,In_250);
nand U497 (N_497,In_504,In_625);
nand U498 (N_498,In_206,In_51);
nor U499 (N_499,In_172,In_23);
and U500 (N_500,N_415,N_225);
nand U501 (N_501,N_214,N_103);
and U502 (N_502,N_108,N_483);
and U503 (N_503,N_399,N_482);
nor U504 (N_504,N_292,N_0);
nor U505 (N_505,N_142,N_55);
or U506 (N_506,N_72,N_394);
nand U507 (N_507,N_141,N_280);
and U508 (N_508,N_379,N_139);
nand U509 (N_509,N_322,N_97);
nand U510 (N_510,N_429,N_365);
or U511 (N_511,N_318,N_132);
nor U512 (N_512,N_347,N_244);
and U513 (N_513,N_77,N_145);
nand U514 (N_514,N_282,N_8);
nand U515 (N_515,N_431,N_408);
or U516 (N_516,N_1,N_271);
and U517 (N_517,N_478,N_239);
xor U518 (N_518,N_422,N_126);
and U519 (N_519,N_276,N_200);
nor U520 (N_520,N_81,N_363);
nand U521 (N_521,N_310,N_265);
nand U522 (N_522,N_87,N_261);
and U523 (N_523,N_411,N_376);
nand U524 (N_524,N_30,N_341);
or U525 (N_525,N_140,N_161);
or U526 (N_526,N_75,N_168);
and U527 (N_527,N_488,N_116);
and U528 (N_528,N_304,N_333);
nor U529 (N_529,N_66,N_306);
or U530 (N_530,N_20,N_86);
nand U531 (N_531,N_180,N_237);
or U532 (N_532,N_136,N_451);
nand U533 (N_533,N_383,N_85);
and U534 (N_534,N_144,N_95);
or U535 (N_535,N_315,N_209);
nor U536 (N_536,N_38,N_238);
and U537 (N_537,N_91,N_442);
nor U538 (N_538,N_236,N_264);
or U539 (N_539,N_491,N_308);
nor U540 (N_540,N_187,N_455);
nor U541 (N_541,N_36,N_395);
nand U542 (N_542,N_406,N_332);
or U543 (N_543,N_459,N_252);
nor U544 (N_544,N_39,N_270);
and U545 (N_545,N_346,N_42);
nor U546 (N_546,N_45,N_21);
or U547 (N_547,N_336,N_405);
nor U548 (N_548,N_438,N_288);
nor U549 (N_549,N_243,N_289);
nor U550 (N_550,N_471,N_106);
or U551 (N_551,N_47,N_358);
nor U552 (N_552,N_190,N_249);
or U553 (N_553,N_465,N_217);
nand U554 (N_554,N_98,N_389);
and U555 (N_555,N_207,N_246);
and U556 (N_556,N_477,N_247);
and U557 (N_557,N_344,N_109);
or U558 (N_558,N_211,N_165);
nand U559 (N_559,N_170,N_498);
nor U560 (N_560,N_469,N_114);
nand U561 (N_561,N_7,N_96);
nor U562 (N_562,N_460,N_281);
or U563 (N_563,N_226,N_256);
nand U564 (N_564,N_125,N_414);
nand U565 (N_565,N_294,N_423);
nor U566 (N_566,N_439,N_386);
nand U567 (N_567,N_354,N_10);
xnor U568 (N_568,N_495,N_392);
xnor U569 (N_569,N_120,N_11);
nand U570 (N_570,N_195,N_361);
or U571 (N_571,N_413,N_221);
xor U572 (N_572,N_100,N_84);
nor U573 (N_573,N_14,N_489);
xnor U574 (N_574,N_291,N_172);
and U575 (N_575,N_430,N_324);
nand U576 (N_576,N_157,N_260);
or U577 (N_577,N_240,N_44);
or U578 (N_578,N_352,N_94);
or U579 (N_579,N_60,N_150);
xnor U580 (N_580,N_343,N_51);
nor U581 (N_581,N_296,N_2);
and U582 (N_582,N_378,N_49);
nand U583 (N_583,N_257,N_421);
or U584 (N_584,N_335,N_104);
and U585 (N_585,N_267,N_130);
or U586 (N_586,N_171,N_162);
or U587 (N_587,N_339,N_334);
nand U588 (N_588,N_462,N_362);
or U589 (N_589,N_436,N_184);
or U590 (N_590,N_115,N_48);
nand U591 (N_591,N_191,N_192);
nand U592 (N_592,N_416,N_305);
or U593 (N_593,N_353,N_326);
and U594 (N_594,N_447,N_204);
or U595 (N_595,N_232,N_121);
nor U596 (N_596,N_17,N_242);
or U597 (N_597,N_377,N_409);
or U598 (N_598,N_188,N_245);
or U599 (N_599,N_432,N_258);
nand U600 (N_600,N_90,N_402);
or U601 (N_601,N_490,N_351);
or U602 (N_602,N_317,N_71);
or U603 (N_603,N_69,N_396);
and U604 (N_604,N_403,N_481);
nor U605 (N_605,N_57,N_128);
or U606 (N_606,N_299,N_388);
or U607 (N_607,N_152,N_286);
or U608 (N_608,N_201,N_53);
and U609 (N_609,N_387,N_183);
and U610 (N_610,N_163,N_360);
nor U611 (N_611,N_70,N_407);
nand U612 (N_612,N_325,N_149);
or U613 (N_613,N_368,N_342);
nor U614 (N_614,N_233,N_375);
nand U615 (N_615,N_230,N_227);
or U616 (N_616,N_173,N_425);
and U617 (N_617,N_496,N_56);
nand U618 (N_618,N_493,N_63);
nor U619 (N_619,N_381,N_146);
or U620 (N_620,N_28,N_273);
and U621 (N_621,N_215,N_297);
nand U622 (N_622,N_34,N_16);
or U623 (N_623,N_25,N_174);
and U624 (N_624,N_102,N_213);
or U625 (N_625,N_167,N_446);
nor U626 (N_626,N_337,N_228);
nand U627 (N_627,N_40,N_400);
nand U628 (N_628,N_330,N_176);
nand U629 (N_629,N_164,N_359);
or U630 (N_630,N_390,N_220);
and U631 (N_631,N_216,N_338);
nor U632 (N_632,N_302,N_208);
and U633 (N_633,N_418,N_251);
or U634 (N_634,N_275,N_457);
and U635 (N_635,N_456,N_205);
nor U636 (N_636,N_279,N_156);
and U637 (N_637,N_487,N_129);
nor U638 (N_638,N_196,N_99);
or U639 (N_639,N_340,N_259);
or U640 (N_640,N_486,N_22);
nor U641 (N_641,N_73,N_440);
nand U642 (N_642,N_92,N_127);
nor U643 (N_643,N_175,N_119);
nor U644 (N_644,N_229,N_124);
nand U645 (N_645,N_159,N_366);
nor U646 (N_646,N_262,N_449);
nand U647 (N_647,N_29,N_50);
nand U648 (N_648,N_79,N_143);
or U649 (N_649,N_316,N_198);
and U650 (N_650,N_74,N_224);
and U651 (N_651,N_307,N_428);
nand U652 (N_652,N_373,N_268);
nand U653 (N_653,N_82,N_367);
and U654 (N_654,N_112,N_287);
nand U655 (N_655,N_492,N_355);
and U656 (N_656,N_357,N_277);
and U657 (N_657,N_350,N_218);
nand U658 (N_658,N_154,N_435);
or U659 (N_659,N_107,N_193);
or U660 (N_660,N_470,N_475);
and U661 (N_661,N_369,N_467);
nor U662 (N_662,N_59,N_284);
nor U663 (N_663,N_466,N_210);
nor U664 (N_664,N_35,N_382);
and U665 (N_665,N_160,N_474);
and U666 (N_666,N_248,N_452);
nor U667 (N_667,N_274,N_424);
or U668 (N_668,N_253,N_177);
or U669 (N_669,N_133,N_298);
nor U670 (N_670,N_371,N_364);
nand U671 (N_671,N_3,N_453);
and U672 (N_672,N_329,N_398);
nor U673 (N_673,N_155,N_443);
and U674 (N_674,N_293,N_24);
or U675 (N_675,N_185,N_328);
nor U676 (N_676,N_393,N_15);
and U677 (N_677,N_178,N_485);
nor U678 (N_678,N_153,N_122);
or U679 (N_679,N_6,N_254);
or U680 (N_680,N_202,N_76);
nor U681 (N_681,N_283,N_348);
nand U682 (N_682,N_151,N_313);
and U683 (N_683,N_263,N_101);
or U684 (N_684,N_345,N_58);
nor U685 (N_685,N_219,N_309);
nand U686 (N_686,N_468,N_327);
nand U687 (N_687,N_410,N_5);
nor U688 (N_688,N_148,N_78);
nor U689 (N_689,N_80,N_131);
or U690 (N_690,N_255,N_179);
and U691 (N_691,N_67,N_27);
nor U692 (N_692,N_295,N_52);
nand U693 (N_693,N_300,N_111);
nand U694 (N_694,N_461,N_83);
or U695 (N_695,N_123,N_319);
or U696 (N_696,N_448,N_182);
nor U697 (N_697,N_88,N_349);
and U698 (N_698,N_323,N_480);
and U699 (N_699,N_206,N_412);
and U700 (N_700,N_427,N_441);
and U701 (N_701,N_9,N_93);
nor U702 (N_702,N_181,N_118);
or U703 (N_703,N_311,N_473);
or U704 (N_704,N_54,N_397);
and U705 (N_705,N_479,N_444);
and U706 (N_706,N_222,N_499);
or U707 (N_707,N_241,N_12);
or U708 (N_708,N_321,N_43);
nor U709 (N_709,N_138,N_419);
nor U710 (N_710,N_68,N_41);
nand U711 (N_711,N_89,N_32);
and U712 (N_712,N_4,N_235);
nor U713 (N_713,N_426,N_137);
and U714 (N_714,N_356,N_134);
and U715 (N_715,N_18,N_212);
or U716 (N_716,N_391,N_46);
or U717 (N_717,N_189,N_61);
nand U718 (N_718,N_272,N_105);
and U719 (N_719,N_135,N_445);
nor U720 (N_720,N_401,N_231);
and U721 (N_721,N_19,N_117);
nand U722 (N_722,N_266,N_62);
and U723 (N_723,N_186,N_31);
nand U724 (N_724,N_33,N_380);
and U725 (N_725,N_372,N_433);
nand U726 (N_726,N_301,N_197);
and U727 (N_727,N_417,N_147);
or U728 (N_728,N_37,N_472);
nor U729 (N_729,N_303,N_278);
and U730 (N_730,N_463,N_384);
nand U731 (N_731,N_385,N_166);
nor U732 (N_732,N_454,N_158);
nor U733 (N_733,N_497,N_194);
nor U734 (N_734,N_26,N_437);
nand U735 (N_735,N_23,N_476);
and U736 (N_736,N_404,N_458);
and U737 (N_737,N_420,N_331);
and U738 (N_738,N_223,N_110);
nand U739 (N_739,N_290,N_234);
nand U740 (N_740,N_314,N_464);
nor U741 (N_741,N_374,N_65);
or U742 (N_742,N_450,N_64);
nor U743 (N_743,N_203,N_199);
nand U744 (N_744,N_113,N_250);
and U745 (N_745,N_484,N_494);
nand U746 (N_746,N_269,N_370);
nor U747 (N_747,N_320,N_13);
nor U748 (N_748,N_169,N_285);
or U749 (N_749,N_312,N_434);
and U750 (N_750,N_363,N_41);
or U751 (N_751,N_84,N_222);
and U752 (N_752,N_154,N_434);
nor U753 (N_753,N_233,N_219);
or U754 (N_754,N_499,N_275);
nor U755 (N_755,N_137,N_349);
or U756 (N_756,N_37,N_9);
xor U757 (N_757,N_394,N_391);
nor U758 (N_758,N_242,N_303);
nor U759 (N_759,N_115,N_436);
and U760 (N_760,N_177,N_143);
and U761 (N_761,N_160,N_0);
nor U762 (N_762,N_155,N_183);
nor U763 (N_763,N_321,N_413);
or U764 (N_764,N_457,N_421);
or U765 (N_765,N_124,N_117);
nor U766 (N_766,N_373,N_361);
xnor U767 (N_767,N_403,N_427);
nor U768 (N_768,N_493,N_132);
nand U769 (N_769,N_105,N_381);
nand U770 (N_770,N_324,N_31);
nand U771 (N_771,N_380,N_112);
nand U772 (N_772,N_181,N_95);
nor U773 (N_773,N_223,N_88);
or U774 (N_774,N_5,N_433);
nor U775 (N_775,N_262,N_428);
and U776 (N_776,N_334,N_414);
and U777 (N_777,N_472,N_336);
or U778 (N_778,N_467,N_280);
xor U779 (N_779,N_115,N_10);
or U780 (N_780,N_166,N_390);
or U781 (N_781,N_470,N_463);
and U782 (N_782,N_461,N_1);
nor U783 (N_783,N_210,N_294);
or U784 (N_784,N_201,N_420);
nand U785 (N_785,N_81,N_18);
xor U786 (N_786,N_226,N_353);
and U787 (N_787,N_135,N_179);
nand U788 (N_788,N_5,N_278);
or U789 (N_789,N_368,N_20);
and U790 (N_790,N_368,N_430);
nand U791 (N_791,N_122,N_256);
nand U792 (N_792,N_11,N_376);
nor U793 (N_793,N_386,N_93);
and U794 (N_794,N_151,N_391);
and U795 (N_795,N_379,N_190);
nand U796 (N_796,N_392,N_88);
nand U797 (N_797,N_331,N_427);
nand U798 (N_798,N_246,N_380);
nor U799 (N_799,N_157,N_146);
and U800 (N_800,N_39,N_144);
and U801 (N_801,N_48,N_257);
and U802 (N_802,N_76,N_126);
nor U803 (N_803,N_134,N_468);
or U804 (N_804,N_285,N_418);
and U805 (N_805,N_160,N_136);
or U806 (N_806,N_368,N_275);
or U807 (N_807,N_361,N_108);
nor U808 (N_808,N_180,N_193);
nand U809 (N_809,N_2,N_138);
or U810 (N_810,N_235,N_345);
nand U811 (N_811,N_51,N_233);
nand U812 (N_812,N_74,N_171);
and U813 (N_813,N_466,N_129);
nor U814 (N_814,N_244,N_492);
or U815 (N_815,N_49,N_63);
nor U816 (N_816,N_250,N_111);
and U817 (N_817,N_150,N_217);
and U818 (N_818,N_7,N_346);
nor U819 (N_819,N_88,N_103);
nor U820 (N_820,N_474,N_91);
nand U821 (N_821,N_463,N_16);
nor U822 (N_822,N_28,N_256);
nand U823 (N_823,N_413,N_231);
or U824 (N_824,N_195,N_208);
and U825 (N_825,N_386,N_473);
and U826 (N_826,N_412,N_363);
nand U827 (N_827,N_18,N_418);
nor U828 (N_828,N_100,N_134);
nand U829 (N_829,N_300,N_374);
nand U830 (N_830,N_459,N_10);
or U831 (N_831,N_113,N_218);
and U832 (N_832,N_218,N_76);
nand U833 (N_833,N_459,N_422);
nor U834 (N_834,N_343,N_107);
or U835 (N_835,N_151,N_284);
nand U836 (N_836,N_122,N_271);
nand U837 (N_837,N_346,N_404);
and U838 (N_838,N_78,N_418);
nand U839 (N_839,N_423,N_422);
and U840 (N_840,N_138,N_33);
nand U841 (N_841,N_64,N_394);
xor U842 (N_842,N_82,N_228);
nand U843 (N_843,N_336,N_113);
nor U844 (N_844,N_296,N_24);
nor U845 (N_845,N_135,N_53);
nand U846 (N_846,N_100,N_468);
nand U847 (N_847,N_198,N_6);
nor U848 (N_848,N_302,N_205);
or U849 (N_849,N_387,N_66);
or U850 (N_850,N_341,N_334);
or U851 (N_851,N_306,N_186);
or U852 (N_852,N_290,N_126);
and U853 (N_853,N_425,N_318);
or U854 (N_854,N_268,N_485);
nor U855 (N_855,N_253,N_291);
or U856 (N_856,N_141,N_118);
and U857 (N_857,N_13,N_336);
or U858 (N_858,N_156,N_346);
and U859 (N_859,N_326,N_342);
nand U860 (N_860,N_283,N_218);
or U861 (N_861,N_77,N_256);
or U862 (N_862,N_77,N_4);
nor U863 (N_863,N_150,N_359);
nor U864 (N_864,N_71,N_192);
and U865 (N_865,N_492,N_218);
nor U866 (N_866,N_156,N_416);
and U867 (N_867,N_335,N_128);
or U868 (N_868,N_366,N_107);
nor U869 (N_869,N_323,N_181);
nand U870 (N_870,N_272,N_206);
and U871 (N_871,N_49,N_19);
nor U872 (N_872,N_52,N_65);
and U873 (N_873,N_103,N_455);
or U874 (N_874,N_55,N_489);
and U875 (N_875,N_387,N_93);
nor U876 (N_876,N_225,N_317);
and U877 (N_877,N_99,N_484);
or U878 (N_878,N_47,N_237);
nand U879 (N_879,N_60,N_134);
or U880 (N_880,N_475,N_117);
and U881 (N_881,N_97,N_69);
and U882 (N_882,N_17,N_77);
or U883 (N_883,N_53,N_91);
nand U884 (N_884,N_112,N_327);
nor U885 (N_885,N_190,N_96);
nand U886 (N_886,N_289,N_36);
and U887 (N_887,N_10,N_217);
nor U888 (N_888,N_107,N_361);
nand U889 (N_889,N_195,N_146);
and U890 (N_890,N_298,N_424);
nand U891 (N_891,N_407,N_291);
nor U892 (N_892,N_124,N_114);
or U893 (N_893,N_59,N_16);
nand U894 (N_894,N_275,N_456);
nor U895 (N_895,N_65,N_325);
xnor U896 (N_896,N_369,N_170);
nor U897 (N_897,N_338,N_270);
nand U898 (N_898,N_54,N_475);
or U899 (N_899,N_372,N_388);
or U900 (N_900,N_92,N_268);
nand U901 (N_901,N_286,N_401);
or U902 (N_902,N_462,N_417);
nand U903 (N_903,N_224,N_471);
nor U904 (N_904,N_273,N_174);
or U905 (N_905,N_376,N_249);
nor U906 (N_906,N_499,N_462);
nand U907 (N_907,N_89,N_222);
or U908 (N_908,N_446,N_93);
nand U909 (N_909,N_24,N_359);
nand U910 (N_910,N_91,N_93);
or U911 (N_911,N_340,N_458);
nand U912 (N_912,N_391,N_415);
nand U913 (N_913,N_473,N_479);
nand U914 (N_914,N_25,N_161);
and U915 (N_915,N_173,N_414);
or U916 (N_916,N_15,N_244);
xor U917 (N_917,N_78,N_160);
nor U918 (N_918,N_209,N_250);
nand U919 (N_919,N_251,N_181);
xor U920 (N_920,N_169,N_81);
or U921 (N_921,N_424,N_262);
or U922 (N_922,N_345,N_189);
nand U923 (N_923,N_341,N_433);
or U924 (N_924,N_146,N_156);
or U925 (N_925,N_70,N_304);
nand U926 (N_926,N_225,N_82);
nand U927 (N_927,N_328,N_476);
or U928 (N_928,N_311,N_235);
and U929 (N_929,N_365,N_173);
nor U930 (N_930,N_368,N_239);
or U931 (N_931,N_241,N_332);
or U932 (N_932,N_250,N_162);
nor U933 (N_933,N_499,N_334);
nor U934 (N_934,N_247,N_439);
nand U935 (N_935,N_89,N_238);
nand U936 (N_936,N_99,N_59);
nor U937 (N_937,N_175,N_309);
nor U938 (N_938,N_58,N_488);
xnor U939 (N_939,N_212,N_281);
nand U940 (N_940,N_185,N_335);
and U941 (N_941,N_400,N_364);
nand U942 (N_942,N_242,N_58);
nand U943 (N_943,N_57,N_294);
nand U944 (N_944,N_469,N_196);
and U945 (N_945,N_196,N_120);
xnor U946 (N_946,N_395,N_272);
and U947 (N_947,N_300,N_201);
nor U948 (N_948,N_349,N_136);
nand U949 (N_949,N_97,N_186);
or U950 (N_950,N_475,N_353);
and U951 (N_951,N_257,N_130);
xor U952 (N_952,N_282,N_29);
and U953 (N_953,N_56,N_168);
nor U954 (N_954,N_164,N_478);
and U955 (N_955,N_208,N_213);
nand U956 (N_956,N_205,N_55);
or U957 (N_957,N_484,N_162);
nor U958 (N_958,N_254,N_398);
nand U959 (N_959,N_481,N_50);
nand U960 (N_960,N_236,N_300);
or U961 (N_961,N_149,N_4);
or U962 (N_962,N_47,N_64);
nor U963 (N_963,N_442,N_5);
nand U964 (N_964,N_311,N_350);
and U965 (N_965,N_386,N_409);
nor U966 (N_966,N_327,N_1);
and U967 (N_967,N_308,N_370);
nor U968 (N_968,N_131,N_7);
nand U969 (N_969,N_42,N_117);
or U970 (N_970,N_169,N_296);
or U971 (N_971,N_120,N_378);
or U972 (N_972,N_297,N_208);
or U973 (N_973,N_52,N_264);
and U974 (N_974,N_185,N_397);
nand U975 (N_975,N_308,N_66);
and U976 (N_976,N_269,N_454);
and U977 (N_977,N_208,N_393);
and U978 (N_978,N_375,N_440);
xnor U979 (N_979,N_93,N_225);
nor U980 (N_980,N_213,N_123);
nor U981 (N_981,N_219,N_49);
or U982 (N_982,N_256,N_338);
nand U983 (N_983,N_129,N_365);
nor U984 (N_984,N_264,N_84);
nor U985 (N_985,N_224,N_99);
and U986 (N_986,N_435,N_246);
nor U987 (N_987,N_253,N_228);
nor U988 (N_988,N_208,N_44);
or U989 (N_989,N_477,N_116);
nand U990 (N_990,N_482,N_384);
nor U991 (N_991,N_394,N_399);
nor U992 (N_992,N_364,N_27);
nand U993 (N_993,N_367,N_336);
nand U994 (N_994,N_369,N_345);
nor U995 (N_995,N_130,N_360);
and U996 (N_996,N_399,N_267);
and U997 (N_997,N_120,N_328);
nor U998 (N_998,N_485,N_279);
or U999 (N_999,N_94,N_419);
nand U1000 (N_1000,N_529,N_633);
or U1001 (N_1001,N_601,N_688);
xnor U1002 (N_1002,N_854,N_807);
and U1003 (N_1003,N_751,N_883);
or U1004 (N_1004,N_581,N_746);
nand U1005 (N_1005,N_742,N_717);
and U1006 (N_1006,N_936,N_701);
or U1007 (N_1007,N_938,N_882);
or U1008 (N_1008,N_800,N_921);
xor U1009 (N_1009,N_690,N_985);
or U1010 (N_1010,N_755,N_747);
nand U1011 (N_1011,N_712,N_886);
or U1012 (N_1012,N_665,N_649);
or U1013 (N_1013,N_924,N_514);
xnor U1014 (N_1014,N_906,N_692);
nor U1015 (N_1015,N_887,N_796);
or U1016 (N_1016,N_743,N_720);
and U1017 (N_1017,N_585,N_607);
or U1018 (N_1018,N_542,N_651);
and U1019 (N_1019,N_675,N_845);
nor U1020 (N_1020,N_672,N_741);
nand U1021 (N_1021,N_940,N_805);
and U1022 (N_1022,N_899,N_830);
nand U1023 (N_1023,N_918,N_713);
nor U1024 (N_1024,N_782,N_991);
or U1025 (N_1025,N_867,N_826);
or U1026 (N_1026,N_729,N_892);
nand U1027 (N_1027,N_863,N_605);
or U1028 (N_1028,N_731,N_547);
nand U1029 (N_1029,N_669,N_614);
nor U1030 (N_1030,N_656,N_652);
nand U1031 (N_1031,N_990,N_997);
and U1032 (N_1032,N_943,N_659);
nor U1033 (N_1033,N_785,N_726);
or U1034 (N_1034,N_803,N_880);
xor U1035 (N_1035,N_523,N_853);
or U1036 (N_1036,N_591,N_513);
or U1037 (N_1037,N_630,N_655);
nand U1038 (N_1038,N_543,N_679);
nand U1039 (N_1039,N_502,N_801);
nor U1040 (N_1040,N_986,N_587);
nor U1041 (N_1041,N_761,N_709);
and U1042 (N_1042,N_572,N_508);
nand U1043 (N_1043,N_610,N_766);
or U1044 (N_1044,N_848,N_916);
nand U1045 (N_1045,N_932,N_973);
nand U1046 (N_1046,N_745,N_628);
or U1047 (N_1047,N_645,N_597);
nor U1048 (N_1048,N_603,N_919);
nor U1049 (N_1049,N_788,N_862);
nand U1050 (N_1050,N_784,N_974);
or U1051 (N_1051,N_933,N_522);
nand U1052 (N_1052,N_507,N_964);
nor U1053 (N_1053,N_976,N_898);
nor U1054 (N_1054,N_811,N_617);
or U1055 (N_1055,N_846,N_517);
and U1056 (N_1056,N_632,N_576);
and U1057 (N_1057,N_714,N_871);
nor U1058 (N_1058,N_842,N_825);
and U1059 (N_1059,N_643,N_901);
and U1060 (N_1060,N_978,N_759);
and U1061 (N_1061,N_841,N_627);
and U1062 (N_1062,N_577,N_773);
or U1063 (N_1063,N_935,N_639);
nor U1064 (N_1064,N_828,N_872);
and U1065 (N_1065,N_571,N_954);
nand U1066 (N_1066,N_903,N_735);
nor U1067 (N_1067,N_822,N_718);
nor U1068 (N_1068,N_550,N_777);
nor U1069 (N_1069,N_516,N_667);
and U1070 (N_1070,N_972,N_604);
nand U1071 (N_1071,N_793,N_691);
nor U1072 (N_1072,N_531,N_538);
nor U1073 (N_1073,N_913,N_911);
nand U1074 (N_1074,N_948,N_677);
and U1075 (N_1075,N_570,N_536);
nor U1076 (N_1076,N_917,N_928);
nor U1077 (N_1077,N_860,N_855);
nor U1078 (N_1078,N_982,N_699);
xor U1079 (N_1079,N_551,N_975);
nand U1080 (N_1080,N_923,N_983);
and U1081 (N_1081,N_635,N_795);
xnor U1082 (N_1082,N_874,N_806);
nand U1083 (N_1083,N_897,N_590);
nor U1084 (N_1084,N_967,N_922);
nor U1085 (N_1085,N_599,N_647);
nor U1086 (N_1086,N_808,N_984);
nand U1087 (N_1087,N_900,N_721);
or U1088 (N_1088,N_566,N_840);
nand U1089 (N_1089,N_578,N_998);
and U1090 (N_1090,N_787,N_686);
and U1091 (N_1091,N_774,N_624);
or U1092 (N_1092,N_650,N_733);
nor U1093 (N_1093,N_579,N_783);
or U1094 (N_1094,N_682,N_750);
or U1095 (N_1095,N_512,N_560);
nand U1096 (N_1096,N_958,N_956);
nand U1097 (N_1097,N_953,N_879);
or U1098 (N_1098,N_518,N_562);
or U1099 (N_1099,N_676,N_891);
or U1100 (N_1100,N_563,N_920);
xnor U1101 (N_1101,N_817,N_980);
nor U1102 (N_1102,N_625,N_569);
nand U1103 (N_1103,N_809,N_963);
and U1104 (N_1104,N_820,N_937);
and U1105 (N_1105,N_565,N_559);
nand U1106 (N_1106,N_832,N_949);
nand U1107 (N_1107,N_705,N_707);
nor U1108 (N_1108,N_827,N_979);
and U1109 (N_1109,N_541,N_893);
or U1110 (N_1110,N_525,N_527);
and U1111 (N_1111,N_763,N_754);
nand U1112 (N_1112,N_545,N_671);
nor U1113 (N_1113,N_866,N_668);
nand U1114 (N_1114,N_528,N_544);
or U1115 (N_1115,N_503,N_837);
and U1116 (N_1116,N_524,N_584);
nand U1117 (N_1117,N_697,N_670);
or U1118 (N_1118,N_770,N_810);
and U1119 (N_1119,N_574,N_902);
and U1120 (N_1120,N_798,N_723);
or U1121 (N_1121,N_548,N_957);
or U1122 (N_1122,N_619,N_869);
xor U1123 (N_1123,N_553,N_646);
nand U1124 (N_1124,N_878,N_909);
and U1125 (N_1125,N_724,N_642);
nand U1126 (N_1126,N_678,N_595);
nand U1127 (N_1127,N_533,N_849);
or U1128 (N_1128,N_873,N_926);
or U1129 (N_1129,N_818,N_945);
or U1130 (N_1130,N_965,N_996);
and U1131 (N_1131,N_775,N_521);
or U1132 (N_1132,N_950,N_737);
nor U1133 (N_1133,N_764,N_987);
or U1134 (N_1134,N_526,N_685);
or U1135 (N_1135,N_895,N_698);
and U1136 (N_1136,N_684,N_988);
or U1137 (N_1137,N_567,N_561);
nor U1138 (N_1138,N_716,N_575);
nor U1139 (N_1139,N_749,N_725);
nor U1140 (N_1140,N_905,N_658);
nor U1141 (N_1141,N_977,N_680);
and U1142 (N_1142,N_884,N_532);
and U1143 (N_1143,N_520,N_865);
or U1144 (N_1144,N_621,N_703);
or U1145 (N_1145,N_776,N_802);
nor U1146 (N_1146,N_812,N_674);
nand U1147 (N_1147,N_952,N_598);
or U1148 (N_1148,N_637,N_934);
nor U1149 (N_1149,N_947,N_816);
nand U1150 (N_1150,N_641,N_704);
and U1151 (N_1151,N_765,N_758);
nand U1152 (N_1152,N_715,N_992);
or U1153 (N_1153,N_780,N_653);
or U1154 (N_1154,N_583,N_861);
nand U1155 (N_1155,N_748,N_804);
and U1156 (N_1156,N_836,N_552);
or U1157 (N_1157,N_711,N_589);
or U1158 (N_1158,N_555,N_819);
or U1159 (N_1159,N_896,N_593);
nor U1160 (N_1160,N_994,N_944);
or U1161 (N_1161,N_689,N_654);
nand U1162 (N_1162,N_968,N_662);
and U1163 (N_1163,N_626,N_960);
and U1164 (N_1164,N_888,N_885);
or U1165 (N_1165,N_814,N_852);
or U1166 (N_1166,N_657,N_702);
nor U1167 (N_1167,N_694,N_821);
and U1168 (N_1168,N_600,N_500);
and U1169 (N_1169,N_999,N_843);
or U1170 (N_1170,N_681,N_663);
nor U1171 (N_1171,N_790,N_823);
nand U1172 (N_1172,N_615,N_847);
and U1173 (N_1173,N_908,N_835);
nor U1174 (N_1174,N_606,N_586);
or U1175 (N_1175,N_534,N_970);
nand U1176 (N_1176,N_505,N_719);
nand U1177 (N_1177,N_875,N_666);
and U1178 (N_1178,N_969,N_622);
or U1179 (N_1179,N_580,N_734);
and U1180 (N_1180,N_789,N_915);
nor U1181 (N_1181,N_907,N_504);
nor U1182 (N_1182,N_501,N_596);
and U1183 (N_1183,N_673,N_594);
nor U1184 (N_1184,N_611,N_772);
nand U1185 (N_1185,N_582,N_870);
or U1186 (N_1186,N_740,N_588);
or U1187 (N_1187,N_881,N_834);
nor U1188 (N_1188,N_608,N_592);
or U1189 (N_1189,N_638,N_760);
nor U1190 (N_1190,N_797,N_894);
and U1191 (N_1191,N_959,N_941);
nor U1192 (N_1192,N_564,N_831);
and U1193 (N_1193,N_939,N_786);
and U1194 (N_1194,N_540,N_955);
nor U1195 (N_1195,N_912,N_813);
and U1196 (N_1196,N_993,N_864);
xnor U1197 (N_1197,N_558,N_781);
and U1198 (N_1198,N_696,N_877);
or U1199 (N_1199,N_556,N_769);
and U1200 (N_1200,N_573,N_931);
nor U1201 (N_1201,N_549,N_660);
and U1202 (N_1202,N_539,N_644);
nand U1203 (N_1203,N_868,N_929);
nand U1204 (N_1204,N_791,N_951);
nand U1205 (N_1205,N_620,N_616);
and U1206 (N_1206,N_962,N_857);
nor U1207 (N_1207,N_876,N_752);
nand U1208 (N_1208,N_613,N_925);
nor U1209 (N_1209,N_708,N_609);
nor U1210 (N_1210,N_732,N_930);
nor U1211 (N_1211,N_727,N_554);
and U1212 (N_1212,N_792,N_664);
and U1213 (N_1213,N_757,N_744);
nor U1214 (N_1214,N_768,N_966);
nor U1215 (N_1215,N_506,N_889);
and U1216 (N_1216,N_511,N_850);
nand U1217 (N_1217,N_636,N_629);
and U1218 (N_1218,N_634,N_833);
and U1219 (N_1219,N_736,N_537);
and U1220 (N_1220,N_693,N_722);
nand U1221 (N_1221,N_858,N_910);
and U1222 (N_1222,N_859,N_989);
nand U1223 (N_1223,N_683,N_710);
nand U1224 (N_1224,N_509,N_568);
or U1225 (N_1225,N_927,N_839);
or U1226 (N_1226,N_648,N_631);
and U1227 (N_1227,N_612,N_728);
nand U1228 (N_1228,N_794,N_838);
nand U1229 (N_1229,N_971,N_762);
nand U1230 (N_1230,N_890,N_535);
or U1231 (N_1231,N_530,N_946);
nor U1232 (N_1232,N_687,N_738);
nor U1233 (N_1233,N_623,N_942);
nand U1234 (N_1234,N_851,N_515);
nor U1235 (N_1235,N_557,N_904);
nor U1236 (N_1236,N_661,N_995);
and U1237 (N_1237,N_753,N_730);
or U1238 (N_1238,N_829,N_778);
nor U1239 (N_1239,N_700,N_981);
nor U1240 (N_1240,N_706,N_618);
nor U1241 (N_1241,N_640,N_767);
or U1242 (N_1242,N_961,N_771);
or U1243 (N_1243,N_856,N_546);
nand U1244 (N_1244,N_914,N_824);
nand U1245 (N_1245,N_510,N_799);
nand U1246 (N_1246,N_695,N_815);
and U1247 (N_1247,N_844,N_756);
nor U1248 (N_1248,N_779,N_602);
nand U1249 (N_1249,N_739,N_519);
nand U1250 (N_1250,N_693,N_910);
nand U1251 (N_1251,N_819,N_742);
nor U1252 (N_1252,N_651,N_725);
and U1253 (N_1253,N_799,N_743);
nor U1254 (N_1254,N_874,N_578);
or U1255 (N_1255,N_820,N_687);
nand U1256 (N_1256,N_564,N_715);
and U1257 (N_1257,N_957,N_608);
nand U1258 (N_1258,N_623,N_615);
or U1259 (N_1259,N_564,N_804);
nor U1260 (N_1260,N_927,N_983);
and U1261 (N_1261,N_816,N_608);
or U1262 (N_1262,N_855,N_606);
or U1263 (N_1263,N_681,N_814);
and U1264 (N_1264,N_948,N_551);
nand U1265 (N_1265,N_911,N_833);
nor U1266 (N_1266,N_819,N_545);
or U1267 (N_1267,N_977,N_708);
nor U1268 (N_1268,N_821,N_558);
nand U1269 (N_1269,N_927,N_988);
and U1270 (N_1270,N_794,N_984);
and U1271 (N_1271,N_651,N_669);
nand U1272 (N_1272,N_851,N_670);
nor U1273 (N_1273,N_622,N_787);
and U1274 (N_1274,N_908,N_916);
and U1275 (N_1275,N_651,N_627);
or U1276 (N_1276,N_945,N_843);
and U1277 (N_1277,N_901,N_978);
or U1278 (N_1278,N_780,N_887);
xor U1279 (N_1279,N_622,N_814);
and U1280 (N_1280,N_899,N_637);
nor U1281 (N_1281,N_647,N_871);
nor U1282 (N_1282,N_613,N_642);
nand U1283 (N_1283,N_915,N_783);
nand U1284 (N_1284,N_739,N_515);
nor U1285 (N_1285,N_785,N_566);
nand U1286 (N_1286,N_574,N_528);
nor U1287 (N_1287,N_636,N_891);
nand U1288 (N_1288,N_519,N_924);
nor U1289 (N_1289,N_636,N_526);
nand U1290 (N_1290,N_637,N_784);
or U1291 (N_1291,N_720,N_588);
nor U1292 (N_1292,N_795,N_902);
and U1293 (N_1293,N_830,N_987);
nand U1294 (N_1294,N_911,N_580);
or U1295 (N_1295,N_972,N_921);
and U1296 (N_1296,N_680,N_911);
nor U1297 (N_1297,N_713,N_806);
and U1298 (N_1298,N_715,N_557);
nor U1299 (N_1299,N_986,N_878);
or U1300 (N_1300,N_979,N_730);
nand U1301 (N_1301,N_513,N_757);
nand U1302 (N_1302,N_753,N_934);
nor U1303 (N_1303,N_864,N_906);
nand U1304 (N_1304,N_629,N_582);
xnor U1305 (N_1305,N_896,N_828);
nor U1306 (N_1306,N_760,N_923);
nor U1307 (N_1307,N_661,N_688);
or U1308 (N_1308,N_766,N_532);
nand U1309 (N_1309,N_649,N_691);
and U1310 (N_1310,N_569,N_610);
and U1311 (N_1311,N_978,N_910);
nor U1312 (N_1312,N_779,N_937);
or U1313 (N_1313,N_725,N_901);
nor U1314 (N_1314,N_660,N_747);
and U1315 (N_1315,N_870,N_561);
and U1316 (N_1316,N_966,N_619);
nand U1317 (N_1317,N_984,N_788);
nor U1318 (N_1318,N_787,N_743);
nor U1319 (N_1319,N_593,N_659);
nand U1320 (N_1320,N_714,N_611);
or U1321 (N_1321,N_572,N_900);
nor U1322 (N_1322,N_848,N_979);
or U1323 (N_1323,N_649,N_859);
and U1324 (N_1324,N_817,N_705);
and U1325 (N_1325,N_834,N_807);
and U1326 (N_1326,N_611,N_618);
nand U1327 (N_1327,N_718,N_834);
nand U1328 (N_1328,N_796,N_624);
nand U1329 (N_1329,N_917,N_963);
xor U1330 (N_1330,N_755,N_873);
and U1331 (N_1331,N_809,N_804);
nor U1332 (N_1332,N_648,N_668);
nand U1333 (N_1333,N_927,N_824);
or U1334 (N_1334,N_587,N_589);
nand U1335 (N_1335,N_921,N_629);
xor U1336 (N_1336,N_667,N_540);
nand U1337 (N_1337,N_943,N_547);
and U1338 (N_1338,N_785,N_586);
nor U1339 (N_1339,N_720,N_671);
or U1340 (N_1340,N_626,N_755);
or U1341 (N_1341,N_524,N_638);
nor U1342 (N_1342,N_978,N_998);
or U1343 (N_1343,N_870,N_801);
nor U1344 (N_1344,N_943,N_895);
and U1345 (N_1345,N_775,N_574);
or U1346 (N_1346,N_812,N_715);
nand U1347 (N_1347,N_849,N_704);
and U1348 (N_1348,N_544,N_693);
nor U1349 (N_1349,N_819,N_731);
or U1350 (N_1350,N_597,N_923);
or U1351 (N_1351,N_594,N_661);
nor U1352 (N_1352,N_853,N_929);
nand U1353 (N_1353,N_686,N_601);
or U1354 (N_1354,N_612,N_785);
nand U1355 (N_1355,N_841,N_849);
nor U1356 (N_1356,N_982,N_822);
nand U1357 (N_1357,N_588,N_654);
nand U1358 (N_1358,N_953,N_667);
and U1359 (N_1359,N_883,N_774);
or U1360 (N_1360,N_792,N_812);
and U1361 (N_1361,N_875,N_572);
nand U1362 (N_1362,N_987,N_541);
nand U1363 (N_1363,N_994,N_559);
and U1364 (N_1364,N_792,N_718);
or U1365 (N_1365,N_855,N_782);
or U1366 (N_1366,N_521,N_678);
nand U1367 (N_1367,N_562,N_686);
or U1368 (N_1368,N_992,N_733);
nand U1369 (N_1369,N_970,N_547);
and U1370 (N_1370,N_845,N_850);
or U1371 (N_1371,N_525,N_586);
and U1372 (N_1372,N_764,N_610);
nor U1373 (N_1373,N_890,N_772);
and U1374 (N_1374,N_546,N_542);
nor U1375 (N_1375,N_710,N_902);
or U1376 (N_1376,N_733,N_567);
or U1377 (N_1377,N_671,N_522);
and U1378 (N_1378,N_831,N_709);
nor U1379 (N_1379,N_509,N_519);
or U1380 (N_1380,N_705,N_715);
nor U1381 (N_1381,N_993,N_902);
or U1382 (N_1382,N_998,N_718);
and U1383 (N_1383,N_898,N_809);
nor U1384 (N_1384,N_857,N_680);
nand U1385 (N_1385,N_649,N_962);
or U1386 (N_1386,N_994,N_779);
and U1387 (N_1387,N_640,N_656);
nand U1388 (N_1388,N_533,N_728);
nand U1389 (N_1389,N_772,N_706);
nand U1390 (N_1390,N_867,N_833);
xnor U1391 (N_1391,N_727,N_544);
and U1392 (N_1392,N_902,N_858);
and U1393 (N_1393,N_817,N_617);
or U1394 (N_1394,N_570,N_706);
and U1395 (N_1395,N_514,N_974);
nor U1396 (N_1396,N_765,N_742);
nor U1397 (N_1397,N_689,N_569);
nor U1398 (N_1398,N_559,N_558);
and U1399 (N_1399,N_983,N_641);
nand U1400 (N_1400,N_627,N_660);
and U1401 (N_1401,N_964,N_838);
or U1402 (N_1402,N_639,N_885);
or U1403 (N_1403,N_867,N_642);
or U1404 (N_1404,N_532,N_833);
or U1405 (N_1405,N_826,N_672);
and U1406 (N_1406,N_666,N_784);
nor U1407 (N_1407,N_742,N_504);
nor U1408 (N_1408,N_843,N_867);
nand U1409 (N_1409,N_657,N_756);
or U1410 (N_1410,N_992,N_595);
or U1411 (N_1411,N_999,N_768);
xnor U1412 (N_1412,N_563,N_789);
or U1413 (N_1413,N_682,N_951);
nand U1414 (N_1414,N_718,N_780);
or U1415 (N_1415,N_675,N_564);
nand U1416 (N_1416,N_626,N_775);
nand U1417 (N_1417,N_824,N_761);
nand U1418 (N_1418,N_530,N_904);
nand U1419 (N_1419,N_995,N_683);
or U1420 (N_1420,N_705,N_902);
nand U1421 (N_1421,N_762,N_987);
or U1422 (N_1422,N_547,N_920);
or U1423 (N_1423,N_974,N_517);
or U1424 (N_1424,N_657,N_678);
nand U1425 (N_1425,N_883,N_547);
nor U1426 (N_1426,N_747,N_619);
nand U1427 (N_1427,N_866,N_618);
nand U1428 (N_1428,N_930,N_618);
nor U1429 (N_1429,N_941,N_568);
nand U1430 (N_1430,N_995,N_600);
nor U1431 (N_1431,N_823,N_894);
and U1432 (N_1432,N_507,N_631);
or U1433 (N_1433,N_681,N_662);
or U1434 (N_1434,N_713,N_628);
nor U1435 (N_1435,N_606,N_814);
or U1436 (N_1436,N_737,N_580);
and U1437 (N_1437,N_912,N_995);
and U1438 (N_1438,N_611,N_746);
nand U1439 (N_1439,N_531,N_626);
nand U1440 (N_1440,N_942,N_885);
and U1441 (N_1441,N_774,N_527);
or U1442 (N_1442,N_617,N_940);
nor U1443 (N_1443,N_586,N_562);
or U1444 (N_1444,N_598,N_660);
nor U1445 (N_1445,N_801,N_869);
nor U1446 (N_1446,N_965,N_627);
nor U1447 (N_1447,N_749,N_630);
or U1448 (N_1448,N_859,N_824);
nand U1449 (N_1449,N_931,N_671);
and U1450 (N_1450,N_945,N_937);
or U1451 (N_1451,N_873,N_602);
and U1452 (N_1452,N_791,N_907);
and U1453 (N_1453,N_837,N_794);
xnor U1454 (N_1454,N_646,N_636);
nor U1455 (N_1455,N_703,N_626);
and U1456 (N_1456,N_905,N_974);
and U1457 (N_1457,N_750,N_861);
and U1458 (N_1458,N_853,N_665);
or U1459 (N_1459,N_848,N_773);
or U1460 (N_1460,N_569,N_628);
nand U1461 (N_1461,N_612,N_804);
and U1462 (N_1462,N_892,N_678);
and U1463 (N_1463,N_928,N_670);
and U1464 (N_1464,N_995,N_622);
and U1465 (N_1465,N_791,N_671);
and U1466 (N_1466,N_655,N_853);
nand U1467 (N_1467,N_601,N_707);
and U1468 (N_1468,N_677,N_645);
nand U1469 (N_1469,N_986,N_953);
and U1470 (N_1470,N_791,N_868);
nor U1471 (N_1471,N_938,N_833);
and U1472 (N_1472,N_965,N_990);
nor U1473 (N_1473,N_882,N_833);
nor U1474 (N_1474,N_954,N_695);
nor U1475 (N_1475,N_883,N_677);
and U1476 (N_1476,N_629,N_502);
or U1477 (N_1477,N_930,N_720);
and U1478 (N_1478,N_887,N_655);
and U1479 (N_1479,N_825,N_519);
nand U1480 (N_1480,N_553,N_666);
and U1481 (N_1481,N_735,N_641);
nand U1482 (N_1482,N_836,N_897);
or U1483 (N_1483,N_535,N_641);
nor U1484 (N_1484,N_988,N_696);
or U1485 (N_1485,N_907,N_533);
nor U1486 (N_1486,N_998,N_993);
xor U1487 (N_1487,N_767,N_618);
nor U1488 (N_1488,N_610,N_563);
nor U1489 (N_1489,N_688,N_684);
nand U1490 (N_1490,N_719,N_962);
or U1491 (N_1491,N_857,N_691);
nand U1492 (N_1492,N_726,N_994);
and U1493 (N_1493,N_527,N_840);
or U1494 (N_1494,N_627,N_701);
nand U1495 (N_1495,N_649,N_674);
nor U1496 (N_1496,N_968,N_702);
and U1497 (N_1497,N_783,N_664);
xnor U1498 (N_1498,N_697,N_903);
or U1499 (N_1499,N_907,N_820);
nor U1500 (N_1500,N_1255,N_1159);
and U1501 (N_1501,N_1069,N_1136);
nor U1502 (N_1502,N_1470,N_1102);
nand U1503 (N_1503,N_1172,N_1037);
and U1504 (N_1504,N_1140,N_1410);
or U1505 (N_1505,N_1022,N_1385);
and U1506 (N_1506,N_1349,N_1454);
nor U1507 (N_1507,N_1263,N_1230);
nand U1508 (N_1508,N_1074,N_1226);
nand U1509 (N_1509,N_1082,N_1103);
and U1510 (N_1510,N_1482,N_1256);
or U1511 (N_1511,N_1208,N_1447);
or U1512 (N_1512,N_1291,N_1416);
nor U1513 (N_1513,N_1429,N_1465);
or U1514 (N_1514,N_1408,N_1290);
nor U1515 (N_1515,N_1424,N_1235);
or U1516 (N_1516,N_1307,N_1079);
and U1517 (N_1517,N_1154,N_1005);
or U1518 (N_1518,N_1171,N_1342);
and U1519 (N_1519,N_1064,N_1483);
nand U1520 (N_1520,N_1043,N_1497);
nand U1521 (N_1521,N_1271,N_1071);
nor U1522 (N_1522,N_1295,N_1180);
or U1523 (N_1523,N_1213,N_1117);
nand U1524 (N_1524,N_1135,N_1219);
nand U1525 (N_1525,N_1306,N_1457);
nor U1526 (N_1526,N_1467,N_1355);
or U1527 (N_1527,N_1280,N_1458);
nand U1528 (N_1528,N_1293,N_1088);
or U1529 (N_1529,N_1459,N_1194);
nand U1530 (N_1530,N_1354,N_1125);
or U1531 (N_1531,N_1370,N_1215);
nor U1532 (N_1532,N_1128,N_1020);
or U1533 (N_1533,N_1121,N_1151);
nand U1534 (N_1534,N_1145,N_1203);
nor U1535 (N_1535,N_1216,N_1392);
and U1536 (N_1536,N_1233,N_1024);
and U1537 (N_1537,N_1270,N_1273);
nand U1538 (N_1538,N_1132,N_1100);
xor U1539 (N_1539,N_1432,N_1415);
or U1540 (N_1540,N_1195,N_1218);
and U1541 (N_1541,N_1302,N_1089);
nor U1542 (N_1542,N_1225,N_1409);
and U1543 (N_1543,N_1127,N_1210);
or U1544 (N_1544,N_1214,N_1019);
and U1545 (N_1545,N_1221,N_1201);
or U1546 (N_1546,N_1453,N_1332);
xnor U1547 (N_1547,N_1228,N_1288);
nand U1548 (N_1548,N_1285,N_1443);
nor U1549 (N_1549,N_1407,N_1435);
or U1550 (N_1550,N_1445,N_1404);
and U1551 (N_1551,N_1016,N_1311);
nand U1552 (N_1552,N_1240,N_1181);
and U1553 (N_1553,N_1436,N_1442);
and U1554 (N_1554,N_1394,N_1420);
or U1555 (N_1555,N_1179,N_1199);
and U1556 (N_1556,N_1399,N_1462);
nand U1557 (N_1557,N_1169,N_1264);
or U1558 (N_1558,N_1391,N_1058);
nor U1559 (N_1559,N_1384,N_1249);
nand U1560 (N_1560,N_1490,N_1417);
nand U1561 (N_1561,N_1015,N_1113);
or U1562 (N_1562,N_1041,N_1346);
and U1563 (N_1563,N_1315,N_1124);
nor U1564 (N_1564,N_1418,N_1011);
or U1565 (N_1565,N_1395,N_1223);
or U1566 (N_1566,N_1039,N_1044);
nor U1567 (N_1567,N_1205,N_1473);
and U1568 (N_1568,N_1004,N_1092);
or U1569 (N_1569,N_1091,N_1431);
and U1570 (N_1570,N_1373,N_1345);
nand U1571 (N_1571,N_1419,N_1437);
nand U1572 (N_1572,N_1374,N_1107);
and U1573 (N_1573,N_1364,N_1206);
and U1574 (N_1574,N_1301,N_1237);
nor U1575 (N_1575,N_1254,N_1184);
and U1576 (N_1576,N_1002,N_1193);
nor U1577 (N_1577,N_1006,N_1081);
nand U1578 (N_1578,N_1493,N_1277);
nor U1579 (N_1579,N_1283,N_1001);
nand U1580 (N_1580,N_1086,N_1158);
nand U1581 (N_1581,N_1025,N_1328);
xor U1582 (N_1582,N_1248,N_1455);
nor U1583 (N_1583,N_1098,N_1338);
nand U1584 (N_1584,N_1460,N_1192);
and U1585 (N_1585,N_1087,N_1104);
and U1586 (N_1586,N_1250,N_1350);
or U1587 (N_1587,N_1278,N_1110);
nand U1588 (N_1588,N_1075,N_1475);
or U1589 (N_1589,N_1236,N_1010);
or U1590 (N_1590,N_1109,N_1023);
nand U1591 (N_1591,N_1234,N_1402);
nor U1592 (N_1592,N_1003,N_1094);
nor U1593 (N_1593,N_1351,N_1008);
and U1594 (N_1594,N_1366,N_1065);
nor U1595 (N_1595,N_1299,N_1449);
or U1596 (N_1596,N_1485,N_1347);
nand U1597 (N_1597,N_1292,N_1463);
and U1598 (N_1598,N_1057,N_1472);
nor U1599 (N_1599,N_1247,N_1428);
nor U1600 (N_1600,N_1045,N_1319);
nor U1601 (N_1601,N_1365,N_1260);
nand U1602 (N_1602,N_1155,N_1186);
nor U1603 (N_1603,N_1481,N_1498);
xor U1604 (N_1604,N_1360,N_1489);
nand U1605 (N_1605,N_1294,N_1324);
or U1606 (N_1606,N_1267,N_1153);
nor U1607 (N_1607,N_1251,N_1055);
nor U1608 (N_1608,N_1339,N_1000);
and U1609 (N_1609,N_1170,N_1072);
and U1610 (N_1610,N_1372,N_1448);
or U1611 (N_1611,N_1269,N_1231);
nor U1612 (N_1612,N_1190,N_1007);
or U1613 (N_1613,N_1161,N_1232);
and U1614 (N_1614,N_1330,N_1461);
nor U1615 (N_1615,N_1492,N_1341);
or U1616 (N_1616,N_1376,N_1406);
and U1617 (N_1617,N_1095,N_1242);
nor U1618 (N_1618,N_1176,N_1333);
nor U1619 (N_1619,N_1164,N_1122);
nor U1620 (N_1620,N_1083,N_1411);
or U1621 (N_1621,N_1427,N_1050);
or U1622 (N_1622,N_1438,N_1308);
nor U1623 (N_1623,N_1238,N_1147);
and U1624 (N_1624,N_1452,N_1141);
nand U1625 (N_1625,N_1134,N_1093);
nor U1626 (N_1626,N_1352,N_1137);
nor U1627 (N_1627,N_1476,N_1028);
or U1628 (N_1628,N_1211,N_1266);
and U1629 (N_1629,N_1451,N_1097);
nor U1630 (N_1630,N_1486,N_1099);
nand U1631 (N_1631,N_1059,N_1314);
or U1632 (N_1632,N_1325,N_1337);
nor U1633 (N_1633,N_1297,N_1488);
nor U1634 (N_1634,N_1390,N_1111);
nor U1635 (N_1635,N_1412,N_1054);
nand U1636 (N_1636,N_1101,N_1133);
nor U1637 (N_1637,N_1413,N_1329);
and U1638 (N_1638,N_1320,N_1165);
nand U1639 (N_1639,N_1080,N_1067);
or U1640 (N_1640,N_1336,N_1130);
nand U1641 (N_1641,N_1156,N_1157);
nor U1642 (N_1642,N_1227,N_1393);
nand U1643 (N_1643,N_1163,N_1116);
nand U1644 (N_1644,N_1243,N_1274);
nor U1645 (N_1645,N_1279,N_1353);
nor U1646 (N_1646,N_1479,N_1033);
or U1647 (N_1647,N_1426,N_1388);
and U1648 (N_1648,N_1178,N_1496);
and U1649 (N_1649,N_1123,N_1356);
and U1650 (N_1650,N_1188,N_1035);
or U1651 (N_1651,N_1026,N_1046);
or U1652 (N_1652,N_1009,N_1371);
and U1653 (N_1653,N_1403,N_1491);
xor U1654 (N_1654,N_1316,N_1368);
and U1655 (N_1655,N_1422,N_1143);
nor U1656 (N_1656,N_1217,N_1499);
and U1657 (N_1657,N_1400,N_1450);
or U1658 (N_1658,N_1129,N_1090);
and U1659 (N_1659,N_1272,N_1262);
nand U1660 (N_1660,N_1150,N_1173);
nand U1661 (N_1661,N_1120,N_1160);
nor U1662 (N_1662,N_1114,N_1348);
and U1663 (N_1663,N_1146,N_1335);
and U1664 (N_1664,N_1220,N_1017);
nor U1665 (N_1665,N_1300,N_1477);
nor U1666 (N_1666,N_1466,N_1187);
and U1667 (N_1667,N_1253,N_1284);
and U1668 (N_1668,N_1175,N_1468);
and U1669 (N_1669,N_1139,N_1375);
or U1670 (N_1670,N_1387,N_1068);
nor U1671 (N_1671,N_1398,N_1027);
nand U1672 (N_1672,N_1268,N_1040);
or U1673 (N_1673,N_1085,N_1259);
and U1674 (N_1674,N_1439,N_1484);
nand U1675 (N_1675,N_1474,N_1189);
or U1676 (N_1676,N_1062,N_1167);
nand U1677 (N_1677,N_1317,N_1357);
and U1678 (N_1678,N_1036,N_1197);
or U1679 (N_1679,N_1084,N_1245);
and U1680 (N_1680,N_1367,N_1389);
nand U1681 (N_1681,N_1191,N_1275);
and U1682 (N_1682,N_1287,N_1198);
nand U1683 (N_1683,N_1282,N_1401);
or U1684 (N_1684,N_1444,N_1405);
nor U1685 (N_1685,N_1304,N_1289);
nand U1686 (N_1686,N_1108,N_1321);
nor U1687 (N_1687,N_1362,N_1106);
nor U1688 (N_1688,N_1031,N_1464);
nor U1689 (N_1689,N_1185,N_1433);
nor U1690 (N_1690,N_1014,N_1322);
nand U1691 (N_1691,N_1257,N_1430);
nand U1692 (N_1692,N_1344,N_1309);
or U1693 (N_1693,N_1303,N_1142);
nor U1694 (N_1694,N_1241,N_1029);
or U1695 (N_1695,N_1144,N_1052);
or U1696 (N_1696,N_1048,N_1061);
nor U1697 (N_1697,N_1246,N_1343);
or U1698 (N_1698,N_1305,N_1310);
nor U1699 (N_1699,N_1131,N_1494);
nor U1700 (N_1700,N_1340,N_1182);
nor U1701 (N_1701,N_1363,N_1207);
xor U1702 (N_1702,N_1162,N_1258);
nand U1703 (N_1703,N_1077,N_1381);
nor U1704 (N_1704,N_1204,N_1047);
nor U1705 (N_1705,N_1331,N_1382);
or U1706 (N_1706,N_1032,N_1383);
or U1707 (N_1707,N_1379,N_1377);
or U1708 (N_1708,N_1441,N_1471);
and U1709 (N_1709,N_1149,N_1239);
and U1710 (N_1710,N_1049,N_1323);
and U1711 (N_1711,N_1060,N_1361);
nor U1712 (N_1712,N_1495,N_1177);
or U1713 (N_1713,N_1423,N_1286);
nand U1714 (N_1714,N_1183,N_1119);
nor U1715 (N_1715,N_1440,N_1212);
and U1716 (N_1716,N_1224,N_1229);
or U1717 (N_1717,N_1096,N_1038);
nor U1718 (N_1718,N_1148,N_1030);
or U1719 (N_1719,N_1380,N_1112);
and U1720 (N_1720,N_1327,N_1115);
nor U1721 (N_1721,N_1078,N_1202);
and U1722 (N_1722,N_1076,N_1386);
nor U1723 (N_1723,N_1456,N_1359);
nand U1724 (N_1724,N_1244,N_1478);
nor U1725 (N_1725,N_1053,N_1209);
and U1726 (N_1726,N_1222,N_1166);
or U1727 (N_1727,N_1051,N_1414);
nand U1728 (N_1728,N_1369,N_1265);
or U1729 (N_1729,N_1358,N_1298);
or U1730 (N_1730,N_1034,N_1200);
nor U1731 (N_1731,N_1174,N_1042);
or U1732 (N_1732,N_1446,N_1421);
nor U1733 (N_1733,N_1021,N_1276);
nor U1734 (N_1734,N_1138,N_1261);
nor U1735 (N_1735,N_1196,N_1281);
or U1736 (N_1736,N_1326,N_1012);
nand U1737 (N_1737,N_1118,N_1296);
and U1738 (N_1738,N_1126,N_1425);
and U1739 (N_1739,N_1318,N_1397);
and U1740 (N_1740,N_1070,N_1018);
xor U1741 (N_1741,N_1056,N_1334);
nand U1742 (N_1742,N_1105,N_1434);
nor U1743 (N_1743,N_1312,N_1073);
or U1744 (N_1744,N_1480,N_1313);
or U1745 (N_1745,N_1469,N_1168);
nor U1746 (N_1746,N_1378,N_1396);
or U1747 (N_1747,N_1252,N_1063);
nand U1748 (N_1748,N_1066,N_1013);
nor U1749 (N_1749,N_1152,N_1487);
nor U1750 (N_1750,N_1080,N_1283);
xnor U1751 (N_1751,N_1182,N_1004);
nand U1752 (N_1752,N_1211,N_1038);
or U1753 (N_1753,N_1157,N_1467);
or U1754 (N_1754,N_1000,N_1175);
or U1755 (N_1755,N_1300,N_1026);
nand U1756 (N_1756,N_1247,N_1016);
nand U1757 (N_1757,N_1421,N_1427);
nor U1758 (N_1758,N_1160,N_1423);
nor U1759 (N_1759,N_1451,N_1397);
nand U1760 (N_1760,N_1029,N_1274);
nor U1761 (N_1761,N_1304,N_1328);
or U1762 (N_1762,N_1415,N_1123);
nand U1763 (N_1763,N_1188,N_1144);
or U1764 (N_1764,N_1015,N_1362);
or U1765 (N_1765,N_1411,N_1098);
nand U1766 (N_1766,N_1019,N_1405);
nand U1767 (N_1767,N_1038,N_1360);
nor U1768 (N_1768,N_1005,N_1095);
nand U1769 (N_1769,N_1138,N_1377);
nor U1770 (N_1770,N_1308,N_1338);
and U1771 (N_1771,N_1147,N_1265);
nor U1772 (N_1772,N_1164,N_1317);
nand U1773 (N_1773,N_1016,N_1279);
nor U1774 (N_1774,N_1102,N_1246);
or U1775 (N_1775,N_1296,N_1430);
nand U1776 (N_1776,N_1355,N_1152);
nand U1777 (N_1777,N_1294,N_1269);
nand U1778 (N_1778,N_1334,N_1170);
nand U1779 (N_1779,N_1063,N_1024);
nand U1780 (N_1780,N_1490,N_1319);
and U1781 (N_1781,N_1093,N_1333);
and U1782 (N_1782,N_1100,N_1434);
nor U1783 (N_1783,N_1077,N_1113);
nor U1784 (N_1784,N_1445,N_1039);
or U1785 (N_1785,N_1097,N_1001);
or U1786 (N_1786,N_1426,N_1116);
nor U1787 (N_1787,N_1267,N_1361);
nor U1788 (N_1788,N_1000,N_1390);
nand U1789 (N_1789,N_1469,N_1263);
or U1790 (N_1790,N_1228,N_1180);
nor U1791 (N_1791,N_1069,N_1409);
nor U1792 (N_1792,N_1410,N_1068);
nand U1793 (N_1793,N_1262,N_1292);
and U1794 (N_1794,N_1186,N_1299);
nand U1795 (N_1795,N_1113,N_1484);
nor U1796 (N_1796,N_1158,N_1307);
and U1797 (N_1797,N_1389,N_1018);
nor U1798 (N_1798,N_1335,N_1322);
nand U1799 (N_1799,N_1261,N_1371);
nand U1800 (N_1800,N_1072,N_1236);
nor U1801 (N_1801,N_1239,N_1194);
nor U1802 (N_1802,N_1115,N_1100);
xor U1803 (N_1803,N_1072,N_1498);
and U1804 (N_1804,N_1337,N_1303);
nor U1805 (N_1805,N_1093,N_1280);
or U1806 (N_1806,N_1416,N_1287);
and U1807 (N_1807,N_1048,N_1087);
or U1808 (N_1808,N_1017,N_1475);
or U1809 (N_1809,N_1194,N_1245);
nor U1810 (N_1810,N_1201,N_1153);
and U1811 (N_1811,N_1425,N_1292);
nand U1812 (N_1812,N_1425,N_1212);
nor U1813 (N_1813,N_1198,N_1299);
xnor U1814 (N_1814,N_1309,N_1244);
nor U1815 (N_1815,N_1107,N_1021);
or U1816 (N_1816,N_1457,N_1116);
or U1817 (N_1817,N_1012,N_1297);
nor U1818 (N_1818,N_1117,N_1026);
nor U1819 (N_1819,N_1006,N_1380);
nand U1820 (N_1820,N_1185,N_1105);
and U1821 (N_1821,N_1062,N_1094);
and U1822 (N_1822,N_1284,N_1408);
or U1823 (N_1823,N_1285,N_1280);
or U1824 (N_1824,N_1209,N_1004);
or U1825 (N_1825,N_1419,N_1438);
and U1826 (N_1826,N_1002,N_1054);
or U1827 (N_1827,N_1191,N_1361);
nand U1828 (N_1828,N_1214,N_1304);
nor U1829 (N_1829,N_1246,N_1480);
nor U1830 (N_1830,N_1498,N_1251);
nor U1831 (N_1831,N_1109,N_1145);
or U1832 (N_1832,N_1058,N_1355);
or U1833 (N_1833,N_1098,N_1287);
nor U1834 (N_1834,N_1433,N_1176);
nor U1835 (N_1835,N_1464,N_1038);
and U1836 (N_1836,N_1441,N_1416);
or U1837 (N_1837,N_1067,N_1086);
nor U1838 (N_1838,N_1239,N_1294);
nand U1839 (N_1839,N_1137,N_1471);
or U1840 (N_1840,N_1361,N_1423);
or U1841 (N_1841,N_1104,N_1263);
and U1842 (N_1842,N_1335,N_1267);
nand U1843 (N_1843,N_1228,N_1187);
nand U1844 (N_1844,N_1464,N_1264);
and U1845 (N_1845,N_1306,N_1267);
and U1846 (N_1846,N_1285,N_1490);
and U1847 (N_1847,N_1068,N_1230);
nor U1848 (N_1848,N_1199,N_1432);
nor U1849 (N_1849,N_1494,N_1445);
xor U1850 (N_1850,N_1163,N_1382);
nand U1851 (N_1851,N_1415,N_1484);
nand U1852 (N_1852,N_1030,N_1175);
nand U1853 (N_1853,N_1353,N_1382);
or U1854 (N_1854,N_1017,N_1322);
and U1855 (N_1855,N_1110,N_1144);
nor U1856 (N_1856,N_1405,N_1478);
or U1857 (N_1857,N_1031,N_1363);
and U1858 (N_1858,N_1106,N_1248);
or U1859 (N_1859,N_1271,N_1448);
nor U1860 (N_1860,N_1267,N_1396);
nand U1861 (N_1861,N_1299,N_1438);
nor U1862 (N_1862,N_1495,N_1248);
nor U1863 (N_1863,N_1490,N_1034);
or U1864 (N_1864,N_1422,N_1106);
nor U1865 (N_1865,N_1389,N_1178);
and U1866 (N_1866,N_1336,N_1074);
and U1867 (N_1867,N_1094,N_1110);
xnor U1868 (N_1868,N_1388,N_1183);
nand U1869 (N_1869,N_1046,N_1365);
and U1870 (N_1870,N_1467,N_1269);
nand U1871 (N_1871,N_1148,N_1239);
nor U1872 (N_1872,N_1356,N_1054);
or U1873 (N_1873,N_1051,N_1006);
or U1874 (N_1874,N_1222,N_1154);
nor U1875 (N_1875,N_1221,N_1126);
and U1876 (N_1876,N_1125,N_1081);
and U1877 (N_1877,N_1444,N_1290);
or U1878 (N_1878,N_1143,N_1394);
or U1879 (N_1879,N_1227,N_1280);
nor U1880 (N_1880,N_1367,N_1104);
nand U1881 (N_1881,N_1490,N_1395);
or U1882 (N_1882,N_1152,N_1147);
and U1883 (N_1883,N_1423,N_1279);
or U1884 (N_1884,N_1255,N_1135);
nor U1885 (N_1885,N_1029,N_1493);
nor U1886 (N_1886,N_1195,N_1352);
or U1887 (N_1887,N_1448,N_1163);
or U1888 (N_1888,N_1444,N_1248);
nand U1889 (N_1889,N_1122,N_1036);
or U1890 (N_1890,N_1299,N_1056);
or U1891 (N_1891,N_1347,N_1498);
nor U1892 (N_1892,N_1327,N_1114);
and U1893 (N_1893,N_1480,N_1214);
or U1894 (N_1894,N_1422,N_1217);
nor U1895 (N_1895,N_1360,N_1349);
or U1896 (N_1896,N_1269,N_1135);
or U1897 (N_1897,N_1299,N_1276);
nor U1898 (N_1898,N_1149,N_1130);
or U1899 (N_1899,N_1032,N_1252);
xor U1900 (N_1900,N_1313,N_1071);
nand U1901 (N_1901,N_1228,N_1307);
nor U1902 (N_1902,N_1012,N_1082);
and U1903 (N_1903,N_1218,N_1281);
or U1904 (N_1904,N_1349,N_1391);
nand U1905 (N_1905,N_1364,N_1270);
nor U1906 (N_1906,N_1426,N_1325);
nand U1907 (N_1907,N_1369,N_1099);
or U1908 (N_1908,N_1133,N_1370);
and U1909 (N_1909,N_1262,N_1334);
or U1910 (N_1910,N_1158,N_1031);
nand U1911 (N_1911,N_1079,N_1343);
nand U1912 (N_1912,N_1432,N_1405);
nand U1913 (N_1913,N_1415,N_1106);
and U1914 (N_1914,N_1047,N_1091);
and U1915 (N_1915,N_1101,N_1007);
nand U1916 (N_1916,N_1417,N_1391);
and U1917 (N_1917,N_1151,N_1329);
or U1918 (N_1918,N_1274,N_1132);
nor U1919 (N_1919,N_1217,N_1417);
nor U1920 (N_1920,N_1311,N_1040);
nand U1921 (N_1921,N_1189,N_1192);
and U1922 (N_1922,N_1415,N_1453);
nand U1923 (N_1923,N_1237,N_1431);
or U1924 (N_1924,N_1086,N_1106);
nor U1925 (N_1925,N_1475,N_1271);
nor U1926 (N_1926,N_1027,N_1272);
and U1927 (N_1927,N_1104,N_1079);
nand U1928 (N_1928,N_1004,N_1180);
nor U1929 (N_1929,N_1217,N_1160);
nor U1930 (N_1930,N_1047,N_1431);
or U1931 (N_1931,N_1045,N_1345);
or U1932 (N_1932,N_1445,N_1258);
or U1933 (N_1933,N_1253,N_1010);
nand U1934 (N_1934,N_1172,N_1310);
and U1935 (N_1935,N_1194,N_1296);
nand U1936 (N_1936,N_1042,N_1184);
or U1937 (N_1937,N_1398,N_1438);
or U1938 (N_1938,N_1064,N_1126);
and U1939 (N_1939,N_1337,N_1427);
and U1940 (N_1940,N_1405,N_1145);
nor U1941 (N_1941,N_1413,N_1488);
nand U1942 (N_1942,N_1404,N_1319);
and U1943 (N_1943,N_1462,N_1220);
nor U1944 (N_1944,N_1330,N_1084);
nor U1945 (N_1945,N_1479,N_1365);
nand U1946 (N_1946,N_1335,N_1225);
xnor U1947 (N_1947,N_1418,N_1449);
or U1948 (N_1948,N_1159,N_1439);
nor U1949 (N_1949,N_1218,N_1367);
nand U1950 (N_1950,N_1071,N_1194);
and U1951 (N_1951,N_1136,N_1101);
nand U1952 (N_1952,N_1390,N_1442);
nor U1953 (N_1953,N_1191,N_1215);
and U1954 (N_1954,N_1349,N_1347);
xor U1955 (N_1955,N_1456,N_1085);
or U1956 (N_1956,N_1222,N_1470);
and U1957 (N_1957,N_1416,N_1498);
and U1958 (N_1958,N_1229,N_1090);
or U1959 (N_1959,N_1058,N_1260);
nor U1960 (N_1960,N_1391,N_1133);
nor U1961 (N_1961,N_1398,N_1431);
nand U1962 (N_1962,N_1320,N_1278);
and U1963 (N_1963,N_1378,N_1036);
nand U1964 (N_1964,N_1033,N_1138);
or U1965 (N_1965,N_1178,N_1407);
xnor U1966 (N_1966,N_1470,N_1392);
or U1967 (N_1967,N_1252,N_1107);
and U1968 (N_1968,N_1470,N_1406);
nand U1969 (N_1969,N_1243,N_1367);
or U1970 (N_1970,N_1441,N_1132);
nand U1971 (N_1971,N_1462,N_1078);
nor U1972 (N_1972,N_1167,N_1292);
and U1973 (N_1973,N_1006,N_1367);
nand U1974 (N_1974,N_1375,N_1104);
nor U1975 (N_1975,N_1474,N_1163);
or U1976 (N_1976,N_1278,N_1167);
and U1977 (N_1977,N_1018,N_1353);
nor U1978 (N_1978,N_1457,N_1369);
or U1979 (N_1979,N_1194,N_1301);
nor U1980 (N_1980,N_1233,N_1182);
or U1981 (N_1981,N_1131,N_1180);
nand U1982 (N_1982,N_1024,N_1238);
xnor U1983 (N_1983,N_1171,N_1213);
and U1984 (N_1984,N_1442,N_1295);
nor U1985 (N_1985,N_1497,N_1191);
nand U1986 (N_1986,N_1108,N_1239);
nor U1987 (N_1987,N_1330,N_1234);
nand U1988 (N_1988,N_1105,N_1166);
or U1989 (N_1989,N_1124,N_1094);
and U1990 (N_1990,N_1488,N_1025);
nand U1991 (N_1991,N_1294,N_1412);
or U1992 (N_1992,N_1139,N_1396);
nor U1993 (N_1993,N_1083,N_1323);
nor U1994 (N_1994,N_1148,N_1432);
nand U1995 (N_1995,N_1045,N_1336);
nor U1996 (N_1996,N_1322,N_1010);
nand U1997 (N_1997,N_1201,N_1139);
nand U1998 (N_1998,N_1123,N_1060);
nand U1999 (N_1999,N_1076,N_1229);
nor U2000 (N_2000,N_1597,N_1932);
nor U2001 (N_2001,N_1929,N_1869);
nand U2002 (N_2002,N_1758,N_1826);
xor U2003 (N_2003,N_1855,N_1730);
nor U2004 (N_2004,N_1754,N_1947);
or U2005 (N_2005,N_1797,N_1736);
nand U2006 (N_2006,N_1615,N_1681);
and U2007 (N_2007,N_1726,N_1931);
and U2008 (N_2008,N_1908,N_1960);
nor U2009 (N_2009,N_1545,N_1766);
nand U2010 (N_2010,N_1577,N_1630);
nor U2011 (N_2011,N_1704,N_1712);
nand U2012 (N_2012,N_1665,N_1919);
xor U2013 (N_2013,N_1941,N_1884);
or U2014 (N_2014,N_1689,N_1574);
and U2015 (N_2015,N_1868,N_1567);
nor U2016 (N_2016,N_1557,N_1666);
nand U2017 (N_2017,N_1696,N_1688);
xor U2018 (N_2018,N_1512,N_1638);
nand U2019 (N_2019,N_1786,N_1983);
nor U2020 (N_2020,N_1904,N_1602);
or U2021 (N_2021,N_1737,N_1825);
nor U2022 (N_2022,N_1782,N_1686);
nand U2023 (N_2023,N_1575,N_1639);
and U2024 (N_2024,N_1763,N_1768);
nor U2025 (N_2025,N_1981,N_1711);
and U2026 (N_2026,N_1986,N_1742);
nand U2027 (N_2027,N_1671,N_1971);
or U2028 (N_2028,N_1790,N_1824);
nor U2029 (N_2029,N_1569,N_1540);
nor U2030 (N_2030,N_1857,N_1674);
and U2031 (N_2031,N_1695,N_1753);
nand U2032 (N_2032,N_1834,N_1939);
nand U2033 (N_2033,N_1676,N_1700);
and U2034 (N_2034,N_1649,N_1603);
or U2035 (N_2035,N_1852,N_1579);
and U2036 (N_2036,N_1982,N_1586);
xnor U2037 (N_2037,N_1668,N_1903);
nand U2038 (N_2038,N_1890,N_1535);
nor U2039 (N_2039,N_1769,N_1648);
nor U2040 (N_2040,N_1589,N_1651);
nand U2041 (N_2041,N_1664,N_1654);
and U2042 (N_2042,N_1808,N_1799);
nand U2043 (N_2043,N_1588,N_1678);
nor U2044 (N_2044,N_1605,N_1815);
nor U2045 (N_2045,N_1895,N_1902);
or U2046 (N_2046,N_1999,N_1514);
or U2047 (N_2047,N_1593,N_1778);
nor U2048 (N_2048,N_1988,N_1634);
and U2049 (N_2049,N_1820,N_1523);
and U2050 (N_2050,N_1622,N_1755);
nor U2051 (N_2051,N_1706,N_1838);
and U2052 (N_2052,N_1800,N_1858);
or U2053 (N_2053,N_1905,N_1746);
nand U2054 (N_2054,N_1827,N_1504);
nor U2055 (N_2055,N_1814,N_1894);
or U2056 (N_2056,N_1608,N_1672);
xor U2057 (N_2057,N_1566,N_1546);
nand U2058 (N_2058,N_1954,N_1631);
and U2059 (N_2059,N_1796,N_1604);
nor U2060 (N_2060,N_1750,N_1946);
nor U2061 (N_2061,N_1531,N_1701);
nand U2062 (N_2062,N_1515,N_1990);
nand U2063 (N_2063,N_1585,N_1937);
nor U2064 (N_2064,N_1773,N_1793);
nor U2065 (N_2065,N_1658,N_1744);
and U2066 (N_2066,N_1979,N_1859);
and U2067 (N_2067,N_1560,N_1973);
and U2068 (N_2068,N_1707,N_1779);
nor U2069 (N_2069,N_1819,N_1770);
nand U2070 (N_2070,N_1916,N_1760);
or U2071 (N_2071,N_1961,N_1691);
xor U2072 (N_2072,N_1740,N_1774);
and U2073 (N_2073,N_1538,N_1853);
nand U2074 (N_2074,N_1980,N_1771);
nor U2075 (N_2075,N_1644,N_1974);
xnor U2076 (N_2076,N_1835,N_1731);
nor U2077 (N_2077,N_1636,N_1612);
and U2078 (N_2078,N_1611,N_1992);
and U2079 (N_2079,N_1616,N_1866);
nand U2080 (N_2080,N_1831,N_1762);
and U2081 (N_2081,N_1870,N_1518);
or U2082 (N_2082,N_1969,N_1710);
xnor U2083 (N_2083,N_1703,N_1867);
nand U2084 (N_2084,N_1993,N_1759);
nand U2085 (N_2085,N_1801,N_1875);
or U2086 (N_2086,N_1544,N_1617);
or U2087 (N_2087,N_1502,N_1930);
and U2088 (N_2088,N_1886,N_1956);
and U2089 (N_2089,N_1832,N_1907);
nor U2090 (N_2090,N_1529,N_1526);
nor U2091 (N_2091,N_1887,N_1692);
nor U2092 (N_2092,N_1508,N_1807);
and U2093 (N_2093,N_1896,N_1547);
or U2094 (N_2094,N_1909,N_1849);
and U2095 (N_2095,N_1965,N_1717);
nor U2096 (N_2096,N_1606,N_1977);
or U2097 (N_2097,N_1967,N_1976);
or U2098 (N_2098,N_1739,N_1923);
and U2099 (N_2099,N_1581,N_1830);
nand U2100 (N_2100,N_1794,N_1513);
and U2101 (N_2101,N_1662,N_1901);
nor U2102 (N_2102,N_1959,N_1541);
or U2103 (N_2103,N_1618,N_1747);
and U2104 (N_2104,N_1511,N_1848);
and U2105 (N_2105,N_1705,N_1724);
or U2106 (N_2106,N_1532,N_1863);
nor U2107 (N_2107,N_1576,N_1880);
and U2108 (N_2108,N_1558,N_1922);
nand U2109 (N_2109,N_1955,N_1765);
nor U2110 (N_2110,N_1891,N_1600);
or U2111 (N_2111,N_1893,N_1856);
and U2112 (N_2112,N_1554,N_1530);
nand U2113 (N_2113,N_1687,N_1876);
nand U2114 (N_2114,N_1964,N_1524);
and U2115 (N_2115,N_1989,N_1548);
and U2116 (N_2116,N_1879,N_1985);
xor U2117 (N_2117,N_1670,N_1645);
nand U2118 (N_2118,N_1877,N_1623);
nor U2119 (N_2119,N_1728,N_1564);
or U2120 (N_2120,N_1520,N_1667);
and U2121 (N_2121,N_1836,N_1915);
and U2122 (N_2122,N_1663,N_1503);
and U2123 (N_2123,N_1738,N_1940);
nor U2124 (N_2124,N_1713,N_1935);
and U2125 (N_2125,N_1972,N_1818);
nor U2126 (N_2126,N_1934,N_1551);
nand U2127 (N_2127,N_1571,N_1539);
nand U2128 (N_2128,N_1556,N_1632);
and U2129 (N_2129,N_1963,N_1673);
nand U2130 (N_2130,N_1805,N_1791);
or U2131 (N_2131,N_1889,N_1998);
nand U2132 (N_2132,N_1783,N_1719);
or U2133 (N_2133,N_1806,N_1629);
and U2134 (N_2134,N_1614,N_1698);
nor U2135 (N_2135,N_1563,N_1913);
and U2136 (N_2136,N_1748,N_1709);
nor U2137 (N_2137,N_1810,N_1823);
and U2138 (N_2138,N_1573,N_1910);
nand U2139 (N_2139,N_1509,N_1860);
and U2140 (N_2140,N_1635,N_1613);
nor U2141 (N_2141,N_1735,N_1792);
nand U2142 (N_2142,N_1975,N_1525);
and U2143 (N_2143,N_1817,N_1987);
nor U2144 (N_2144,N_1897,N_1950);
and U2145 (N_2145,N_1685,N_1920);
nor U2146 (N_2146,N_1995,N_1777);
and U2147 (N_2147,N_1693,N_1840);
nand U2148 (N_2148,N_1854,N_1669);
or U2149 (N_2149,N_1591,N_1592);
or U2150 (N_2150,N_1928,N_1552);
nor U2151 (N_2151,N_1590,N_1565);
and U2152 (N_2152,N_1751,N_1694);
nor U2153 (N_2153,N_1561,N_1568);
nor U2154 (N_2154,N_1752,N_1756);
and U2155 (N_2155,N_1528,N_1659);
nor U2156 (N_2156,N_1862,N_1757);
nand U2157 (N_2157,N_1533,N_1828);
or U2158 (N_2158,N_1723,N_1882);
or U2159 (N_2159,N_1843,N_1656);
or U2160 (N_2160,N_1516,N_1720);
and U2161 (N_2161,N_1802,N_1921);
nand U2162 (N_2162,N_1761,N_1690);
nor U2163 (N_2163,N_1583,N_1924);
or U2164 (N_2164,N_1521,N_1850);
nand U2165 (N_2165,N_1610,N_1708);
xor U2166 (N_2166,N_1637,N_1749);
or U2167 (N_2167,N_1718,N_1958);
nor U2168 (N_2168,N_1732,N_1549);
nor U2169 (N_2169,N_1625,N_1596);
and U2170 (N_2170,N_1957,N_1871);
and U2171 (N_2171,N_1599,N_1714);
nor U2172 (N_2172,N_1675,N_1865);
and U2173 (N_2173,N_1925,N_1609);
and U2174 (N_2174,N_1679,N_1944);
nor U2175 (N_2175,N_1519,N_1580);
and U2176 (N_2176,N_1507,N_1813);
nor U2177 (N_2177,N_1809,N_1842);
nor U2178 (N_2178,N_1517,N_1780);
or U2179 (N_2179,N_1727,N_1966);
and U2180 (N_2180,N_1968,N_1626);
nor U2181 (N_2181,N_1506,N_1847);
nor U2182 (N_2182,N_1646,N_1888);
nor U2183 (N_2183,N_1510,N_1945);
nor U2184 (N_2184,N_1785,N_1788);
and U2185 (N_2185,N_1845,N_1984);
nand U2186 (N_2186,N_1846,N_1822);
or U2187 (N_2187,N_1741,N_1733);
nor U2188 (N_2188,N_1627,N_1899);
nor U2189 (N_2189,N_1505,N_1816);
xnor U2190 (N_2190,N_1917,N_1864);
or U2191 (N_2191,N_1715,N_1628);
nand U2192 (N_2192,N_1951,N_1952);
or U2193 (N_2193,N_1620,N_1833);
nor U2194 (N_2194,N_1595,N_1578);
or U2195 (N_2195,N_1680,N_1559);
nor U2196 (N_2196,N_1655,N_1885);
or U2197 (N_2197,N_1949,N_1798);
and U2198 (N_2198,N_1878,N_1699);
xnor U2199 (N_2199,N_1997,N_1542);
nor U2200 (N_2200,N_1789,N_1572);
and U2201 (N_2201,N_1594,N_1772);
xor U2202 (N_2202,N_1953,N_1661);
and U2203 (N_2203,N_1943,N_1522);
nand U2204 (N_2204,N_1643,N_1642);
and U2205 (N_2205,N_1537,N_1653);
or U2206 (N_2206,N_1501,N_1500);
nor U2207 (N_2207,N_1861,N_1702);
and U2208 (N_2208,N_1640,N_1550);
or U2209 (N_2209,N_1652,N_1804);
or U2210 (N_2210,N_1641,N_1978);
and U2211 (N_2211,N_1660,N_1781);
nor U2212 (N_2212,N_1633,N_1918);
nand U2213 (N_2213,N_1725,N_1872);
or U2214 (N_2214,N_1795,N_1844);
nand U2215 (N_2215,N_1619,N_1722);
nor U2216 (N_2216,N_1811,N_1948);
or U2217 (N_2217,N_1892,N_1812);
or U2218 (N_2218,N_1926,N_1803);
nor U2219 (N_2219,N_1684,N_1898);
nand U2220 (N_2220,N_1874,N_1734);
nor U2221 (N_2221,N_1677,N_1621);
nor U2222 (N_2222,N_1587,N_1942);
and U2223 (N_2223,N_1562,N_1821);
or U2224 (N_2224,N_1570,N_1657);
nor U2225 (N_2225,N_1697,N_1962);
or U2226 (N_2226,N_1775,N_1914);
or U2227 (N_2227,N_1994,N_1873);
nor U2228 (N_2228,N_1936,N_1624);
and U2229 (N_2229,N_1927,N_1683);
and U2230 (N_2230,N_1991,N_1912);
nor U2231 (N_2231,N_1598,N_1534);
or U2232 (N_2232,N_1716,N_1787);
nand U2233 (N_2233,N_1601,N_1584);
nand U2234 (N_2234,N_1933,N_1527);
and U2235 (N_2235,N_1970,N_1829);
or U2236 (N_2236,N_1881,N_1841);
or U2237 (N_2237,N_1911,N_1839);
or U2238 (N_2238,N_1837,N_1883);
and U2239 (N_2239,N_1582,N_1743);
nor U2240 (N_2240,N_1721,N_1851);
or U2241 (N_2241,N_1650,N_1906);
and U2242 (N_2242,N_1767,N_1553);
nor U2243 (N_2243,N_1938,N_1543);
nor U2244 (N_2244,N_1647,N_1536);
nor U2245 (N_2245,N_1607,N_1776);
or U2246 (N_2246,N_1900,N_1682);
and U2247 (N_2247,N_1764,N_1996);
nand U2248 (N_2248,N_1745,N_1784);
nand U2249 (N_2249,N_1729,N_1555);
xor U2250 (N_2250,N_1534,N_1656);
or U2251 (N_2251,N_1704,N_1542);
nor U2252 (N_2252,N_1949,N_1822);
nand U2253 (N_2253,N_1790,N_1562);
or U2254 (N_2254,N_1708,N_1553);
nand U2255 (N_2255,N_1815,N_1834);
and U2256 (N_2256,N_1900,N_1666);
nor U2257 (N_2257,N_1725,N_1715);
or U2258 (N_2258,N_1520,N_1953);
and U2259 (N_2259,N_1671,N_1806);
nor U2260 (N_2260,N_1748,N_1508);
and U2261 (N_2261,N_1635,N_1781);
nand U2262 (N_2262,N_1955,N_1852);
nand U2263 (N_2263,N_1543,N_1949);
nor U2264 (N_2264,N_1807,N_1672);
nor U2265 (N_2265,N_1745,N_1503);
or U2266 (N_2266,N_1901,N_1668);
nand U2267 (N_2267,N_1507,N_1804);
nand U2268 (N_2268,N_1681,N_1612);
nand U2269 (N_2269,N_1718,N_1940);
nand U2270 (N_2270,N_1928,N_1757);
and U2271 (N_2271,N_1655,N_1794);
nand U2272 (N_2272,N_1842,N_1730);
and U2273 (N_2273,N_1500,N_1829);
or U2274 (N_2274,N_1988,N_1661);
or U2275 (N_2275,N_1841,N_1888);
nor U2276 (N_2276,N_1577,N_1805);
nand U2277 (N_2277,N_1976,N_1700);
or U2278 (N_2278,N_1724,N_1868);
nor U2279 (N_2279,N_1796,N_1999);
or U2280 (N_2280,N_1846,N_1718);
nor U2281 (N_2281,N_1910,N_1811);
or U2282 (N_2282,N_1595,N_1563);
or U2283 (N_2283,N_1870,N_1673);
nor U2284 (N_2284,N_1912,N_1551);
nand U2285 (N_2285,N_1505,N_1720);
nor U2286 (N_2286,N_1690,N_1998);
or U2287 (N_2287,N_1595,N_1728);
or U2288 (N_2288,N_1878,N_1695);
nand U2289 (N_2289,N_1898,N_1966);
nand U2290 (N_2290,N_1874,N_1772);
nand U2291 (N_2291,N_1759,N_1620);
nor U2292 (N_2292,N_1542,N_1863);
nor U2293 (N_2293,N_1921,N_1790);
nor U2294 (N_2294,N_1605,N_1670);
and U2295 (N_2295,N_1574,N_1663);
nand U2296 (N_2296,N_1515,N_1940);
and U2297 (N_2297,N_1722,N_1948);
nor U2298 (N_2298,N_1904,N_1937);
nor U2299 (N_2299,N_1958,N_1554);
nand U2300 (N_2300,N_1878,N_1652);
and U2301 (N_2301,N_1774,N_1504);
or U2302 (N_2302,N_1872,N_1813);
nand U2303 (N_2303,N_1617,N_1938);
and U2304 (N_2304,N_1749,N_1922);
nor U2305 (N_2305,N_1660,N_1776);
nand U2306 (N_2306,N_1614,N_1607);
and U2307 (N_2307,N_1550,N_1875);
nand U2308 (N_2308,N_1814,N_1509);
nand U2309 (N_2309,N_1835,N_1966);
or U2310 (N_2310,N_1652,N_1506);
and U2311 (N_2311,N_1911,N_1685);
and U2312 (N_2312,N_1531,N_1655);
or U2313 (N_2313,N_1502,N_1911);
and U2314 (N_2314,N_1801,N_1639);
nand U2315 (N_2315,N_1997,N_1988);
and U2316 (N_2316,N_1845,N_1803);
nor U2317 (N_2317,N_1557,N_1577);
and U2318 (N_2318,N_1634,N_1970);
and U2319 (N_2319,N_1957,N_1626);
nand U2320 (N_2320,N_1664,N_1826);
nor U2321 (N_2321,N_1911,N_1782);
nand U2322 (N_2322,N_1725,N_1796);
and U2323 (N_2323,N_1708,N_1876);
nor U2324 (N_2324,N_1617,N_1963);
nor U2325 (N_2325,N_1924,N_1715);
nor U2326 (N_2326,N_1952,N_1509);
and U2327 (N_2327,N_1749,N_1853);
or U2328 (N_2328,N_1680,N_1659);
or U2329 (N_2329,N_1840,N_1771);
or U2330 (N_2330,N_1764,N_1941);
nand U2331 (N_2331,N_1708,N_1850);
nand U2332 (N_2332,N_1698,N_1779);
and U2333 (N_2333,N_1565,N_1779);
and U2334 (N_2334,N_1807,N_1747);
and U2335 (N_2335,N_1507,N_1612);
and U2336 (N_2336,N_1745,N_1712);
nand U2337 (N_2337,N_1790,N_1685);
nand U2338 (N_2338,N_1921,N_1586);
xor U2339 (N_2339,N_1805,N_1853);
nor U2340 (N_2340,N_1825,N_1984);
nor U2341 (N_2341,N_1608,N_1600);
and U2342 (N_2342,N_1942,N_1965);
and U2343 (N_2343,N_1727,N_1701);
nand U2344 (N_2344,N_1580,N_1687);
or U2345 (N_2345,N_1583,N_1527);
and U2346 (N_2346,N_1918,N_1580);
nand U2347 (N_2347,N_1598,N_1639);
nand U2348 (N_2348,N_1799,N_1665);
xor U2349 (N_2349,N_1579,N_1778);
and U2350 (N_2350,N_1553,N_1648);
xnor U2351 (N_2351,N_1922,N_1748);
and U2352 (N_2352,N_1914,N_1511);
or U2353 (N_2353,N_1516,N_1733);
nand U2354 (N_2354,N_1741,N_1781);
nand U2355 (N_2355,N_1921,N_1581);
or U2356 (N_2356,N_1893,N_1761);
nand U2357 (N_2357,N_1996,N_1792);
nand U2358 (N_2358,N_1715,N_1606);
or U2359 (N_2359,N_1899,N_1648);
nand U2360 (N_2360,N_1810,N_1544);
nor U2361 (N_2361,N_1793,N_1917);
nand U2362 (N_2362,N_1932,N_1676);
and U2363 (N_2363,N_1726,N_1986);
and U2364 (N_2364,N_1580,N_1825);
and U2365 (N_2365,N_1712,N_1912);
and U2366 (N_2366,N_1866,N_1967);
and U2367 (N_2367,N_1644,N_1764);
and U2368 (N_2368,N_1842,N_1998);
nor U2369 (N_2369,N_1883,N_1946);
and U2370 (N_2370,N_1930,N_1877);
or U2371 (N_2371,N_1854,N_1760);
and U2372 (N_2372,N_1955,N_1827);
nor U2373 (N_2373,N_1600,N_1604);
nor U2374 (N_2374,N_1789,N_1529);
nand U2375 (N_2375,N_1649,N_1970);
nor U2376 (N_2376,N_1761,N_1606);
nor U2377 (N_2377,N_1626,N_1722);
or U2378 (N_2378,N_1686,N_1911);
nor U2379 (N_2379,N_1767,N_1667);
nor U2380 (N_2380,N_1884,N_1646);
nor U2381 (N_2381,N_1568,N_1634);
or U2382 (N_2382,N_1938,N_1571);
or U2383 (N_2383,N_1884,N_1591);
nor U2384 (N_2384,N_1575,N_1541);
xnor U2385 (N_2385,N_1809,N_1605);
and U2386 (N_2386,N_1912,N_1862);
nor U2387 (N_2387,N_1615,N_1610);
and U2388 (N_2388,N_1980,N_1751);
nor U2389 (N_2389,N_1926,N_1734);
and U2390 (N_2390,N_1807,N_1947);
or U2391 (N_2391,N_1864,N_1714);
nor U2392 (N_2392,N_1855,N_1770);
nand U2393 (N_2393,N_1797,N_1934);
nor U2394 (N_2394,N_1847,N_1746);
or U2395 (N_2395,N_1512,N_1696);
xor U2396 (N_2396,N_1942,N_1627);
nor U2397 (N_2397,N_1893,N_1503);
and U2398 (N_2398,N_1689,N_1985);
and U2399 (N_2399,N_1660,N_1609);
nor U2400 (N_2400,N_1784,N_1506);
nand U2401 (N_2401,N_1759,N_1778);
and U2402 (N_2402,N_1728,N_1898);
nand U2403 (N_2403,N_1660,N_1908);
or U2404 (N_2404,N_1523,N_1537);
nand U2405 (N_2405,N_1591,N_1506);
nor U2406 (N_2406,N_1527,N_1600);
nand U2407 (N_2407,N_1732,N_1936);
and U2408 (N_2408,N_1749,N_1949);
nand U2409 (N_2409,N_1842,N_1970);
nand U2410 (N_2410,N_1904,N_1623);
or U2411 (N_2411,N_1703,N_1926);
and U2412 (N_2412,N_1849,N_1781);
and U2413 (N_2413,N_1645,N_1543);
nand U2414 (N_2414,N_1885,N_1719);
nand U2415 (N_2415,N_1997,N_1527);
nand U2416 (N_2416,N_1670,N_1715);
and U2417 (N_2417,N_1772,N_1881);
nand U2418 (N_2418,N_1945,N_1587);
and U2419 (N_2419,N_1637,N_1784);
and U2420 (N_2420,N_1806,N_1996);
nand U2421 (N_2421,N_1773,N_1799);
xnor U2422 (N_2422,N_1765,N_1863);
or U2423 (N_2423,N_1831,N_1700);
and U2424 (N_2424,N_1795,N_1902);
nand U2425 (N_2425,N_1938,N_1940);
and U2426 (N_2426,N_1826,N_1835);
or U2427 (N_2427,N_1657,N_1722);
or U2428 (N_2428,N_1530,N_1622);
nor U2429 (N_2429,N_1907,N_1928);
or U2430 (N_2430,N_1698,N_1644);
nand U2431 (N_2431,N_1653,N_1783);
nor U2432 (N_2432,N_1998,N_1777);
nor U2433 (N_2433,N_1664,N_1920);
or U2434 (N_2434,N_1992,N_1563);
nand U2435 (N_2435,N_1994,N_1595);
nor U2436 (N_2436,N_1570,N_1697);
nand U2437 (N_2437,N_1667,N_1772);
nor U2438 (N_2438,N_1537,N_1700);
or U2439 (N_2439,N_1611,N_1561);
or U2440 (N_2440,N_1673,N_1868);
and U2441 (N_2441,N_1915,N_1657);
and U2442 (N_2442,N_1918,N_1514);
or U2443 (N_2443,N_1805,N_1894);
and U2444 (N_2444,N_1573,N_1793);
nor U2445 (N_2445,N_1996,N_1583);
and U2446 (N_2446,N_1867,N_1736);
nor U2447 (N_2447,N_1535,N_1725);
or U2448 (N_2448,N_1532,N_1669);
and U2449 (N_2449,N_1753,N_1507);
nand U2450 (N_2450,N_1949,N_1850);
or U2451 (N_2451,N_1976,N_1680);
and U2452 (N_2452,N_1708,N_1982);
nand U2453 (N_2453,N_1558,N_1573);
nand U2454 (N_2454,N_1680,N_1648);
xor U2455 (N_2455,N_1684,N_1875);
and U2456 (N_2456,N_1879,N_1680);
and U2457 (N_2457,N_1583,N_1726);
nand U2458 (N_2458,N_1713,N_1514);
nand U2459 (N_2459,N_1901,N_1836);
and U2460 (N_2460,N_1622,N_1823);
and U2461 (N_2461,N_1935,N_1865);
nand U2462 (N_2462,N_1945,N_1616);
or U2463 (N_2463,N_1600,N_1816);
and U2464 (N_2464,N_1698,N_1608);
nand U2465 (N_2465,N_1968,N_1969);
and U2466 (N_2466,N_1998,N_1775);
or U2467 (N_2467,N_1915,N_1858);
or U2468 (N_2468,N_1717,N_1667);
or U2469 (N_2469,N_1940,N_1994);
or U2470 (N_2470,N_1540,N_1584);
nand U2471 (N_2471,N_1900,N_1500);
or U2472 (N_2472,N_1856,N_1742);
nor U2473 (N_2473,N_1756,N_1909);
or U2474 (N_2474,N_1604,N_1512);
nor U2475 (N_2475,N_1560,N_1674);
and U2476 (N_2476,N_1702,N_1684);
or U2477 (N_2477,N_1764,N_1586);
nand U2478 (N_2478,N_1711,N_1611);
nor U2479 (N_2479,N_1503,N_1844);
or U2480 (N_2480,N_1868,N_1590);
or U2481 (N_2481,N_1788,N_1759);
and U2482 (N_2482,N_1644,N_1731);
or U2483 (N_2483,N_1776,N_1601);
or U2484 (N_2484,N_1623,N_1532);
and U2485 (N_2485,N_1807,N_1679);
nand U2486 (N_2486,N_1936,N_1673);
or U2487 (N_2487,N_1961,N_1638);
nor U2488 (N_2488,N_1832,N_1897);
and U2489 (N_2489,N_1970,N_1557);
nor U2490 (N_2490,N_1540,N_1734);
nand U2491 (N_2491,N_1929,N_1626);
or U2492 (N_2492,N_1586,N_1780);
and U2493 (N_2493,N_1566,N_1572);
or U2494 (N_2494,N_1568,N_1818);
nand U2495 (N_2495,N_1794,N_1816);
and U2496 (N_2496,N_1890,N_1665);
nor U2497 (N_2497,N_1503,N_1694);
and U2498 (N_2498,N_1675,N_1666);
nand U2499 (N_2499,N_1979,N_1875);
and U2500 (N_2500,N_2229,N_2387);
and U2501 (N_2501,N_2187,N_2327);
nand U2502 (N_2502,N_2468,N_2351);
nor U2503 (N_2503,N_2049,N_2272);
or U2504 (N_2504,N_2076,N_2415);
or U2505 (N_2505,N_2451,N_2246);
nand U2506 (N_2506,N_2131,N_2066);
nand U2507 (N_2507,N_2305,N_2354);
nor U2508 (N_2508,N_2494,N_2133);
and U2509 (N_2509,N_2158,N_2064);
and U2510 (N_2510,N_2046,N_2202);
or U2511 (N_2511,N_2132,N_2166);
nand U2512 (N_2512,N_2241,N_2162);
and U2513 (N_2513,N_2325,N_2143);
nand U2514 (N_2514,N_2389,N_2273);
nand U2515 (N_2515,N_2038,N_2425);
or U2516 (N_2516,N_2279,N_2465);
and U2517 (N_2517,N_2439,N_2269);
nand U2518 (N_2518,N_2460,N_2237);
nand U2519 (N_2519,N_2270,N_2088);
and U2520 (N_2520,N_2264,N_2379);
and U2521 (N_2521,N_2247,N_2287);
or U2522 (N_2522,N_2381,N_2400);
or U2523 (N_2523,N_2234,N_2386);
nand U2524 (N_2524,N_2320,N_2375);
and U2525 (N_2525,N_2142,N_2337);
and U2526 (N_2526,N_2371,N_2321);
or U2527 (N_2527,N_2115,N_2316);
or U2528 (N_2528,N_2488,N_2182);
nor U2529 (N_2529,N_2150,N_2051);
and U2530 (N_2530,N_2000,N_2409);
nand U2531 (N_2531,N_2188,N_2256);
nor U2532 (N_2532,N_2239,N_2003);
nor U2533 (N_2533,N_2446,N_2498);
or U2534 (N_2534,N_2392,N_2267);
or U2535 (N_2535,N_2346,N_2455);
nor U2536 (N_2536,N_2324,N_2159);
nor U2537 (N_2537,N_2342,N_2277);
and U2538 (N_2538,N_2199,N_2429);
nand U2539 (N_2539,N_2096,N_2084);
and U2540 (N_2540,N_2418,N_2459);
and U2541 (N_2541,N_2200,N_2313);
nand U2542 (N_2542,N_2222,N_2216);
and U2543 (N_2543,N_2397,N_2058);
or U2544 (N_2544,N_2147,N_2353);
or U2545 (N_2545,N_2413,N_2444);
nand U2546 (N_2546,N_2110,N_2406);
and U2547 (N_2547,N_2228,N_2181);
and U2548 (N_2548,N_2016,N_2426);
nand U2549 (N_2549,N_2334,N_2335);
nand U2550 (N_2550,N_2121,N_2274);
and U2551 (N_2551,N_2043,N_2201);
or U2552 (N_2552,N_2242,N_2052);
nor U2553 (N_2553,N_2364,N_2262);
and U2554 (N_2554,N_2411,N_2250);
or U2555 (N_2555,N_2018,N_2490);
or U2556 (N_2556,N_2174,N_2081);
nor U2557 (N_2557,N_2449,N_2124);
nor U2558 (N_2558,N_2231,N_2464);
or U2559 (N_2559,N_2252,N_2218);
xnor U2560 (N_2560,N_2317,N_2170);
or U2561 (N_2561,N_2045,N_2343);
and U2562 (N_2562,N_2394,N_2310);
nor U2563 (N_2563,N_2303,N_2336);
and U2564 (N_2564,N_2326,N_2189);
nand U2565 (N_2565,N_2034,N_2055);
nand U2566 (N_2566,N_2367,N_2276);
or U2567 (N_2567,N_2391,N_2028);
or U2568 (N_2568,N_2295,N_2235);
and U2569 (N_2569,N_2373,N_2308);
or U2570 (N_2570,N_2136,N_2118);
or U2571 (N_2571,N_2022,N_2160);
and U2572 (N_2572,N_2248,N_2315);
nand U2573 (N_2573,N_2238,N_2333);
and U2574 (N_2574,N_2259,N_2141);
nand U2575 (N_2575,N_2251,N_2230);
and U2576 (N_2576,N_2128,N_2447);
or U2577 (N_2577,N_2225,N_2024);
nand U2578 (N_2578,N_2461,N_2497);
and U2579 (N_2579,N_2107,N_2278);
nor U2580 (N_2580,N_2472,N_2332);
or U2581 (N_2581,N_2163,N_2300);
nor U2582 (N_2582,N_2109,N_2341);
or U2583 (N_2583,N_2347,N_2001);
nor U2584 (N_2584,N_2434,N_2035);
and U2585 (N_2585,N_2266,N_2388);
and U2586 (N_2586,N_2258,N_2116);
nand U2587 (N_2587,N_2179,N_2298);
and U2588 (N_2588,N_2029,N_2499);
nor U2589 (N_2589,N_2286,N_2176);
and U2590 (N_2590,N_2099,N_2477);
and U2591 (N_2591,N_2212,N_2495);
nand U2592 (N_2592,N_2196,N_2443);
nand U2593 (N_2593,N_2227,N_2138);
nor U2594 (N_2594,N_2487,N_2173);
or U2595 (N_2595,N_2309,N_2186);
nor U2596 (N_2596,N_2101,N_2011);
or U2597 (N_2597,N_2345,N_2193);
nor U2598 (N_2598,N_2007,N_2338);
nand U2599 (N_2599,N_2184,N_2412);
nor U2600 (N_2600,N_2294,N_2061);
nand U2601 (N_2601,N_2355,N_2289);
or U2602 (N_2602,N_2293,N_2349);
and U2603 (N_2603,N_2169,N_2482);
or U2604 (N_2604,N_2368,N_2220);
nor U2605 (N_2605,N_2493,N_2134);
and U2606 (N_2606,N_2363,N_2476);
or U2607 (N_2607,N_2486,N_2036);
or U2608 (N_2608,N_2438,N_2021);
nand U2609 (N_2609,N_2405,N_2361);
nor U2610 (N_2610,N_2190,N_2205);
nor U2611 (N_2611,N_2430,N_2261);
nand U2612 (N_2612,N_2360,N_2203);
nand U2613 (N_2613,N_2245,N_2090);
and U2614 (N_2614,N_2318,N_2440);
or U2615 (N_2615,N_2466,N_2086);
xnor U2616 (N_2616,N_2208,N_2408);
and U2617 (N_2617,N_2183,N_2232);
nor U2618 (N_2618,N_2399,N_2380);
and U2619 (N_2619,N_2478,N_2078);
and U2620 (N_2620,N_2417,N_2445);
or U2621 (N_2621,N_2129,N_2039);
nor U2622 (N_2622,N_2155,N_2070);
nor U2623 (N_2623,N_2281,N_2023);
nor U2624 (N_2624,N_2019,N_2144);
or U2625 (N_2625,N_2221,N_2005);
xor U2626 (N_2626,N_2057,N_2263);
nor U2627 (N_2627,N_2311,N_2467);
and U2628 (N_2628,N_2420,N_2020);
or U2629 (N_2629,N_2350,N_2180);
nor U2630 (N_2630,N_2114,N_2017);
or U2631 (N_2631,N_2257,N_2204);
nor U2632 (N_2632,N_2106,N_2401);
nor U2633 (N_2633,N_2092,N_2077);
nand U2634 (N_2634,N_2469,N_2140);
nand U2635 (N_2635,N_2376,N_2191);
and U2636 (N_2636,N_2097,N_2479);
nor U2637 (N_2637,N_2284,N_2108);
nand U2638 (N_2638,N_2357,N_2059);
or U2639 (N_2639,N_2348,N_2178);
and U2640 (N_2640,N_2080,N_2285);
xor U2641 (N_2641,N_2312,N_2433);
and U2642 (N_2642,N_2075,N_2253);
nand U2643 (N_2643,N_2123,N_2006);
xor U2644 (N_2644,N_2111,N_2025);
nor U2645 (N_2645,N_2254,N_2172);
or U2646 (N_2646,N_2053,N_2102);
and U2647 (N_2647,N_2307,N_2098);
and U2648 (N_2648,N_2157,N_2044);
and U2649 (N_2649,N_2063,N_2054);
nor U2650 (N_2650,N_2060,N_2339);
nand U2651 (N_2651,N_2456,N_2014);
nand U2652 (N_2652,N_2314,N_2302);
nor U2653 (N_2653,N_2328,N_2291);
nand U2654 (N_2654,N_2359,N_2422);
and U2655 (N_2655,N_2040,N_2026);
nor U2656 (N_2656,N_2441,N_2165);
and U2657 (N_2657,N_2079,N_2062);
and U2658 (N_2658,N_2319,N_2423);
or U2659 (N_2659,N_2370,N_2374);
and U2660 (N_2660,N_2296,N_2395);
or U2661 (N_2661,N_2344,N_2095);
nor U2662 (N_2662,N_2240,N_2330);
nor U2663 (N_2663,N_2483,N_2085);
or U2664 (N_2664,N_2306,N_2475);
and U2665 (N_2665,N_2301,N_2154);
or U2666 (N_2666,N_2236,N_2421);
nand U2667 (N_2667,N_2117,N_2323);
nor U2668 (N_2668,N_2125,N_2027);
nand U2669 (N_2669,N_2175,N_2414);
nor U2670 (N_2670,N_2463,N_2491);
and U2671 (N_2671,N_2292,N_2042);
or U2672 (N_2672,N_2265,N_2452);
and U2673 (N_2673,N_2378,N_2382);
nor U2674 (N_2674,N_2071,N_2083);
and U2675 (N_2675,N_2473,N_2282);
and U2676 (N_2676,N_2072,N_2470);
nor U2677 (N_2677,N_2424,N_2104);
xnor U2678 (N_2678,N_2074,N_2496);
nand U2679 (N_2679,N_2067,N_2219);
or U2680 (N_2680,N_2050,N_2480);
nor U2681 (N_2681,N_2008,N_2145);
nor U2682 (N_2682,N_2171,N_2384);
and U2683 (N_2683,N_2432,N_2177);
nand U2684 (N_2684,N_2304,N_2198);
nor U2685 (N_2685,N_2322,N_2002);
nand U2686 (N_2686,N_2402,N_2185);
nor U2687 (N_2687,N_2358,N_2137);
and U2688 (N_2688,N_2398,N_2105);
nand U2689 (N_2689,N_2094,N_2009);
and U2690 (N_2690,N_2366,N_2103);
and U2691 (N_2691,N_2197,N_2223);
or U2692 (N_2692,N_2037,N_2299);
nor U2693 (N_2693,N_2419,N_2404);
nand U2694 (N_2694,N_2122,N_2195);
nor U2695 (N_2695,N_2288,N_2331);
nor U2696 (N_2696,N_2207,N_2089);
or U2697 (N_2697,N_2087,N_2268);
and U2698 (N_2698,N_2485,N_2416);
or U2699 (N_2699,N_2093,N_2377);
and U2700 (N_2700,N_2120,N_2167);
nor U2701 (N_2701,N_2244,N_2233);
and U2702 (N_2702,N_2436,N_2004);
nand U2703 (N_2703,N_2448,N_2194);
and U2704 (N_2704,N_2091,N_2015);
or U2705 (N_2705,N_2471,N_2290);
or U2706 (N_2706,N_2056,N_2403);
nand U2707 (N_2707,N_2280,N_2489);
nand U2708 (N_2708,N_2492,N_2100);
nand U2709 (N_2709,N_2127,N_2442);
and U2710 (N_2710,N_2032,N_2130);
or U2711 (N_2711,N_2073,N_2151);
xnor U2712 (N_2712,N_2156,N_2393);
nand U2713 (N_2713,N_2012,N_2214);
and U2714 (N_2714,N_2030,N_2457);
nand U2715 (N_2715,N_2010,N_2474);
nand U2716 (N_2716,N_2224,N_2431);
nand U2717 (N_2717,N_2372,N_2340);
nand U2718 (N_2718,N_2329,N_2065);
nor U2719 (N_2719,N_2271,N_2390);
xnor U2720 (N_2720,N_2112,N_2126);
and U2721 (N_2721,N_2210,N_2152);
and U2722 (N_2722,N_2410,N_2135);
and U2723 (N_2723,N_2428,N_2450);
nor U2724 (N_2724,N_2215,N_2396);
or U2725 (N_2725,N_2068,N_2255);
nand U2726 (N_2726,N_2069,N_2148);
or U2727 (N_2727,N_2031,N_2462);
and U2728 (N_2728,N_2033,N_2297);
or U2729 (N_2729,N_2164,N_2048);
nand U2730 (N_2730,N_2484,N_2435);
nor U2731 (N_2731,N_2243,N_2213);
or U2732 (N_2732,N_2454,N_2082);
nor U2733 (N_2733,N_2047,N_2260);
and U2734 (N_2734,N_2211,N_2458);
and U2735 (N_2735,N_2161,N_2153);
nor U2736 (N_2736,N_2013,N_2249);
and U2737 (N_2737,N_2209,N_2206);
or U2738 (N_2738,N_2352,N_2365);
nand U2739 (N_2739,N_2407,N_2226);
and U2740 (N_2740,N_2437,N_2168);
nor U2741 (N_2741,N_2283,N_2146);
or U2742 (N_2742,N_2139,N_2217);
nand U2743 (N_2743,N_2481,N_2119);
nor U2744 (N_2744,N_2369,N_2427);
nand U2745 (N_2745,N_2362,N_2113);
nand U2746 (N_2746,N_2356,N_2192);
nand U2747 (N_2747,N_2149,N_2385);
or U2748 (N_2748,N_2275,N_2041);
nor U2749 (N_2749,N_2453,N_2383);
nor U2750 (N_2750,N_2218,N_2426);
and U2751 (N_2751,N_2458,N_2047);
and U2752 (N_2752,N_2171,N_2014);
nor U2753 (N_2753,N_2063,N_2183);
nor U2754 (N_2754,N_2298,N_2155);
and U2755 (N_2755,N_2475,N_2140);
xnor U2756 (N_2756,N_2433,N_2088);
and U2757 (N_2757,N_2317,N_2054);
nand U2758 (N_2758,N_2099,N_2328);
nand U2759 (N_2759,N_2356,N_2171);
nand U2760 (N_2760,N_2218,N_2339);
nand U2761 (N_2761,N_2463,N_2483);
and U2762 (N_2762,N_2283,N_2148);
nor U2763 (N_2763,N_2401,N_2160);
and U2764 (N_2764,N_2268,N_2303);
or U2765 (N_2765,N_2383,N_2328);
nand U2766 (N_2766,N_2211,N_2027);
nand U2767 (N_2767,N_2359,N_2180);
nor U2768 (N_2768,N_2004,N_2218);
nand U2769 (N_2769,N_2067,N_2472);
or U2770 (N_2770,N_2230,N_2312);
nand U2771 (N_2771,N_2213,N_2220);
nor U2772 (N_2772,N_2402,N_2413);
and U2773 (N_2773,N_2083,N_2085);
nor U2774 (N_2774,N_2186,N_2282);
nor U2775 (N_2775,N_2426,N_2065);
nand U2776 (N_2776,N_2044,N_2195);
nor U2777 (N_2777,N_2093,N_2345);
nor U2778 (N_2778,N_2302,N_2040);
nor U2779 (N_2779,N_2461,N_2296);
or U2780 (N_2780,N_2125,N_2349);
xnor U2781 (N_2781,N_2481,N_2040);
nand U2782 (N_2782,N_2317,N_2366);
xor U2783 (N_2783,N_2160,N_2340);
nor U2784 (N_2784,N_2382,N_2326);
nor U2785 (N_2785,N_2284,N_2303);
nor U2786 (N_2786,N_2116,N_2429);
and U2787 (N_2787,N_2093,N_2347);
nor U2788 (N_2788,N_2003,N_2038);
nor U2789 (N_2789,N_2300,N_2499);
and U2790 (N_2790,N_2036,N_2344);
nor U2791 (N_2791,N_2460,N_2274);
nand U2792 (N_2792,N_2058,N_2123);
or U2793 (N_2793,N_2183,N_2122);
nor U2794 (N_2794,N_2045,N_2376);
nor U2795 (N_2795,N_2473,N_2422);
nand U2796 (N_2796,N_2010,N_2446);
nand U2797 (N_2797,N_2488,N_2408);
and U2798 (N_2798,N_2217,N_2090);
and U2799 (N_2799,N_2367,N_2072);
nor U2800 (N_2800,N_2330,N_2165);
and U2801 (N_2801,N_2294,N_2131);
and U2802 (N_2802,N_2098,N_2040);
and U2803 (N_2803,N_2051,N_2476);
or U2804 (N_2804,N_2116,N_2430);
and U2805 (N_2805,N_2347,N_2449);
or U2806 (N_2806,N_2166,N_2356);
and U2807 (N_2807,N_2328,N_2373);
nand U2808 (N_2808,N_2207,N_2234);
or U2809 (N_2809,N_2406,N_2486);
nor U2810 (N_2810,N_2038,N_2079);
or U2811 (N_2811,N_2195,N_2031);
or U2812 (N_2812,N_2211,N_2427);
nand U2813 (N_2813,N_2047,N_2438);
nor U2814 (N_2814,N_2420,N_2101);
xnor U2815 (N_2815,N_2293,N_2129);
and U2816 (N_2816,N_2339,N_2123);
nor U2817 (N_2817,N_2458,N_2262);
and U2818 (N_2818,N_2410,N_2461);
nor U2819 (N_2819,N_2288,N_2261);
nand U2820 (N_2820,N_2069,N_2311);
nand U2821 (N_2821,N_2025,N_2245);
or U2822 (N_2822,N_2105,N_2189);
or U2823 (N_2823,N_2005,N_2245);
nand U2824 (N_2824,N_2414,N_2077);
nor U2825 (N_2825,N_2146,N_2415);
or U2826 (N_2826,N_2369,N_2091);
and U2827 (N_2827,N_2461,N_2245);
nand U2828 (N_2828,N_2028,N_2108);
and U2829 (N_2829,N_2227,N_2319);
nor U2830 (N_2830,N_2409,N_2312);
or U2831 (N_2831,N_2289,N_2391);
nand U2832 (N_2832,N_2062,N_2180);
or U2833 (N_2833,N_2320,N_2111);
or U2834 (N_2834,N_2470,N_2171);
or U2835 (N_2835,N_2384,N_2489);
nor U2836 (N_2836,N_2388,N_2461);
and U2837 (N_2837,N_2193,N_2395);
nand U2838 (N_2838,N_2380,N_2488);
nor U2839 (N_2839,N_2398,N_2383);
and U2840 (N_2840,N_2154,N_2429);
nand U2841 (N_2841,N_2395,N_2413);
or U2842 (N_2842,N_2069,N_2444);
and U2843 (N_2843,N_2026,N_2446);
nor U2844 (N_2844,N_2180,N_2463);
xnor U2845 (N_2845,N_2350,N_2055);
or U2846 (N_2846,N_2013,N_2163);
nand U2847 (N_2847,N_2104,N_2180);
nor U2848 (N_2848,N_2250,N_2394);
nor U2849 (N_2849,N_2316,N_2095);
and U2850 (N_2850,N_2332,N_2255);
or U2851 (N_2851,N_2095,N_2187);
nor U2852 (N_2852,N_2381,N_2448);
and U2853 (N_2853,N_2219,N_2364);
and U2854 (N_2854,N_2430,N_2130);
and U2855 (N_2855,N_2193,N_2180);
nand U2856 (N_2856,N_2139,N_2092);
or U2857 (N_2857,N_2222,N_2413);
nor U2858 (N_2858,N_2009,N_2271);
or U2859 (N_2859,N_2001,N_2325);
or U2860 (N_2860,N_2113,N_2314);
or U2861 (N_2861,N_2134,N_2474);
nand U2862 (N_2862,N_2202,N_2313);
and U2863 (N_2863,N_2344,N_2076);
nand U2864 (N_2864,N_2133,N_2337);
nor U2865 (N_2865,N_2225,N_2142);
nor U2866 (N_2866,N_2048,N_2114);
and U2867 (N_2867,N_2253,N_2170);
nand U2868 (N_2868,N_2385,N_2346);
nor U2869 (N_2869,N_2029,N_2046);
and U2870 (N_2870,N_2400,N_2289);
nand U2871 (N_2871,N_2460,N_2076);
and U2872 (N_2872,N_2066,N_2204);
nor U2873 (N_2873,N_2383,N_2332);
nor U2874 (N_2874,N_2397,N_2381);
and U2875 (N_2875,N_2164,N_2259);
or U2876 (N_2876,N_2322,N_2493);
or U2877 (N_2877,N_2161,N_2280);
and U2878 (N_2878,N_2297,N_2478);
or U2879 (N_2879,N_2438,N_2072);
or U2880 (N_2880,N_2400,N_2391);
xor U2881 (N_2881,N_2047,N_2171);
and U2882 (N_2882,N_2183,N_2221);
xor U2883 (N_2883,N_2004,N_2339);
nand U2884 (N_2884,N_2376,N_2066);
or U2885 (N_2885,N_2140,N_2219);
or U2886 (N_2886,N_2184,N_2053);
nor U2887 (N_2887,N_2132,N_2099);
nand U2888 (N_2888,N_2440,N_2036);
xnor U2889 (N_2889,N_2129,N_2178);
nand U2890 (N_2890,N_2126,N_2495);
and U2891 (N_2891,N_2106,N_2265);
and U2892 (N_2892,N_2269,N_2295);
xnor U2893 (N_2893,N_2172,N_2286);
or U2894 (N_2894,N_2171,N_2390);
nor U2895 (N_2895,N_2043,N_2121);
nand U2896 (N_2896,N_2179,N_2365);
nor U2897 (N_2897,N_2231,N_2412);
nor U2898 (N_2898,N_2376,N_2402);
xnor U2899 (N_2899,N_2030,N_2461);
nor U2900 (N_2900,N_2320,N_2472);
or U2901 (N_2901,N_2005,N_2259);
nand U2902 (N_2902,N_2010,N_2205);
xnor U2903 (N_2903,N_2141,N_2124);
or U2904 (N_2904,N_2496,N_2493);
nor U2905 (N_2905,N_2216,N_2296);
nand U2906 (N_2906,N_2431,N_2197);
or U2907 (N_2907,N_2494,N_2208);
nor U2908 (N_2908,N_2427,N_2160);
nor U2909 (N_2909,N_2277,N_2134);
nor U2910 (N_2910,N_2427,N_2002);
and U2911 (N_2911,N_2356,N_2160);
nor U2912 (N_2912,N_2042,N_2261);
xnor U2913 (N_2913,N_2232,N_2315);
nor U2914 (N_2914,N_2046,N_2243);
nand U2915 (N_2915,N_2171,N_2362);
nor U2916 (N_2916,N_2456,N_2116);
and U2917 (N_2917,N_2286,N_2053);
or U2918 (N_2918,N_2277,N_2382);
or U2919 (N_2919,N_2434,N_2349);
and U2920 (N_2920,N_2460,N_2481);
nand U2921 (N_2921,N_2479,N_2091);
or U2922 (N_2922,N_2187,N_2460);
nor U2923 (N_2923,N_2447,N_2153);
and U2924 (N_2924,N_2419,N_2272);
nor U2925 (N_2925,N_2051,N_2138);
nor U2926 (N_2926,N_2220,N_2018);
nand U2927 (N_2927,N_2152,N_2340);
and U2928 (N_2928,N_2498,N_2369);
or U2929 (N_2929,N_2272,N_2297);
nand U2930 (N_2930,N_2314,N_2187);
nand U2931 (N_2931,N_2346,N_2336);
nor U2932 (N_2932,N_2465,N_2113);
nor U2933 (N_2933,N_2151,N_2113);
nor U2934 (N_2934,N_2036,N_2370);
nand U2935 (N_2935,N_2143,N_2211);
or U2936 (N_2936,N_2495,N_2039);
nor U2937 (N_2937,N_2499,N_2488);
and U2938 (N_2938,N_2083,N_2328);
nand U2939 (N_2939,N_2493,N_2258);
and U2940 (N_2940,N_2109,N_2133);
nor U2941 (N_2941,N_2420,N_2204);
nor U2942 (N_2942,N_2113,N_2175);
xnor U2943 (N_2943,N_2355,N_2375);
or U2944 (N_2944,N_2186,N_2382);
or U2945 (N_2945,N_2161,N_2382);
nor U2946 (N_2946,N_2344,N_2418);
or U2947 (N_2947,N_2021,N_2493);
and U2948 (N_2948,N_2143,N_2370);
or U2949 (N_2949,N_2100,N_2134);
nor U2950 (N_2950,N_2166,N_2025);
nor U2951 (N_2951,N_2069,N_2426);
or U2952 (N_2952,N_2255,N_2078);
or U2953 (N_2953,N_2370,N_2043);
nand U2954 (N_2954,N_2019,N_2229);
nor U2955 (N_2955,N_2379,N_2332);
or U2956 (N_2956,N_2151,N_2313);
or U2957 (N_2957,N_2377,N_2068);
and U2958 (N_2958,N_2423,N_2052);
xnor U2959 (N_2959,N_2447,N_2386);
or U2960 (N_2960,N_2280,N_2323);
and U2961 (N_2961,N_2445,N_2027);
or U2962 (N_2962,N_2213,N_2358);
nor U2963 (N_2963,N_2137,N_2294);
nor U2964 (N_2964,N_2132,N_2425);
nand U2965 (N_2965,N_2436,N_2149);
nor U2966 (N_2966,N_2423,N_2223);
or U2967 (N_2967,N_2406,N_2269);
xor U2968 (N_2968,N_2164,N_2326);
or U2969 (N_2969,N_2300,N_2374);
nand U2970 (N_2970,N_2299,N_2007);
nand U2971 (N_2971,N_2355,N_2162);
or U2972 (N_2972,N_2125,N_2203);
xor U2973 (N_2973,N_2374,N_2413);
nor U2974 (N_2974,N_2470,N_2413);
and U2975 (N_2975,N_2335,N_2223);
and U2976 (N_2976,N_2347,N_2146);
nor U2977 (N_2977,N_2357,N_2092);
nor U2978 (N_2978,N_2033,N_2226);
or U2979 (N_2979,N_2362,N_2218);
and U2980 (N_2980,N_2221,N_2334);
and U2981 (N_2981,N_2182,N_2356);
or U2982 (N_2982,N_2135,N_2102);
and U2983 (N_2983,N_2421,N_2319);
and U2984 (N_2984,N_2229,N_2036);
nor U2985 (N_2985,N_2061,N_2193);
and U2986 (N_2986,N_2040,N_2394);
nor U2987 (N_2987,N_2280,N_2236);
nand U2988 (N_2988,N_2348,N_2000);
nor U2989 (N_2989,N_2152,N_2473);
nor U2990 (N_2990,N_2392,N_2252);
xor U2991 (N_2991,N_2006,N_2131);
nor U2992 (N_2992,N_2096,N_2131);
or U2993 (N_2993,N_2138,N_2197);
nor U2994 (N_2994,N_2348,N_2025);
and U2995 (N_2995,N_2003,N_2496);
nor U2996 (N_2996,N_2432,N_2238);
and U2997 (N_2997,N_2276,N_2180);
and U2998 (N_2998,N_2290,N_2059);
nor U2999 (N_2999,N_2277,N_2360);
nand U3000 (N_3000,N_2867,N_2929);
nor U3001 (N_3001,N_2646,N_2891);
and U3002 (N_3002,N_2824,N_2710);
nor U3003 (N_3003,N_2656,N_2980);
or U3004 (N_3004,N_2733,N_2946);
and U3005 (N_3005,N_2574,N_2928);
or U3006 (N_3006,N_2709,N_2786);
and U3007 (N_3007,N_2608,N_2758);
nand U3008 (N_3008,N_2887,N_2866);
nand U3009 (N_3009,N_2901,N_2588);
or U3010 (N_3010,N_2586,N_2926);
and U3011 (N_3011,N_2869,N_2550);
nand U3012 (N_3012,N_2868,N_2723);
nand U3013 (N_3013,N_2533,N_2585);
nand U3014 (N_3014,N_2833,N_2689);
and U3015 (N_3015,N_2968,N_2834);
nand U3016 (N_3016,N_2616,N_2697);
nand U3017 (N_3017,N_2982,N_2546);
or U3018 (N_3018,N_2937,N_2587);
or U3019 (N_3019,N_2910,N_2986);
and U3020 (N_3020,N_2857,N_2878);
nand U3021 (N_3021,N_2724,N_2798);
nand U3022 (N_3022,N_2850,N_2781);
or U3023 (N_3023,N_2805,N_2749);
or U3024 (N_3024,N_2516,N_2815);
nor U3025 (N_3025,N_2776,N_2800);
or U3026 (N_3026,N_2806,N_2747);
and U3027 (N_3027,N_2692,N_2995);
or U3028 (N_3028,N_2513,N_2948);
nor U3029 (N_3029,N_2707,N_2602);
nand U3030 (N_3030,N_2969,N_2530);
xnor U3031 (N_3031,N_2638,N_2903);
and U3032 (N_3032,N_2635,N_2790);
or U3033 (N_3033,N_2793,N_2764);
nor U3034 (N_3034,N_2832,N_2782);
nand U3035 (N_3035,N_2503,N_2770);
or U3036 (N_3036,N_2556,N_2994);
or U3037 (N_3037,N_2898,N_2897);
nor U3038 (N_3038,N_2951,N_2807);
nand U3039 (N_3039,N_2693,N_2779);
or U3040 (N_3040,N_2892,N_2900);
or U3041 (N_3041,N_2729,N_2979);
nor U3042 (N_3042,N_2597,N_2902);
or U3043 (N_3043,N_2886,N_2642);
or U3044 (N_3044,N_2988,N_2727);
xnor U3045 (N_3045,N_2541,N_2877);
and U3046 (N_3046,N_2792,N_2610);
nand U3047 (N_3047,N_2543,N_2852);
nor U3048 (N_3048,N_2680,N_2939);
and U3049 (N_3049,N_2531,N_2744);
nor U3050 (N_3050,N_2880,N_2768);
or U3051 (N_3051,N_2913,N_2978);
and U3052 (N_3052,N_2835,N_2737);
and U3053 (N_3053,N_2548,N_2873);
and U3054 (N_3054,N_2820,N_2535);
and U3055 (N_3055,N_2812,N_2767);
and U3056 (N_3056,N_2771,N_2645);
nor U3057 (N_3057,N_2829,N_2853);
nand U3058 (N_3058,N_2904,N_2593);
nand U3059 (N_3059,N_2931,N_2644);
or U3060 (N_3060,N_2917,N_2778);
or U3061 (N_3061,N_2840,N_2662);
and U3062 (N_3062,N_2571,N_2589);
and U3063 (N_3063,N_2705,N_2554);
nand U3064 (N_3064,N_2759,N_2676);
nand U3065 (N_3065,N_2669,N_2651);
or U3066 (N_3066,N_2665,N_2943);
and U3067 (N_3067,N_2906,N_2508);
or U3068 (N_3068,N_2804,N_2801);
or U3069 (N_3069,N_2679,N_2912);
nand U3070 (N_3070,N_2997,N_2769);
and U3071 (N_3071,N_2990,N_2510);
or U3072 (N_3072,N_2506,N_2861);
nor U3073 (N_3073,N_2884,N_2848);
nor U3074 (N_3074,N_2915,N_2675);
and U3075 (N_3075,N_2989,N_2713);
nor U3076 (N_3076,N_2971,N_2624);
and U3077 (N_3077,N_2843,N_2681);
nand U3078 (N_3078,N_2722,N_2636);
or U3079 (N_3079,N_2717,N_2564);
nand U3080 (N_3080,N_2984,N_2736);
or U3081 (N_3081,N_2844,N_2514);
xor U3082 (N_3082,N_2562,N_2935);
or U3083 (N_3083,N_2975,N_2592);
nor U3084 (N_3084,N_2615,N_2696);
and U3085 (N_3085,N_2598,N_2753);
and U3086 (N_3086,N_2816,N_2673);
or U3087 (N_3087,N_2613,N_2629);
and U3088 (N_3088,N_2558,N_2687);
nand U3089 (N_3089,N_2742,N_2750);
and U3090 (N_3090,N_2607,N_2938);
and U3091 (N_3091,N_2691,N_2936);
or U3092 (N_3092,N_2596,N_2667);
or U3093 (N_3093,N_2991,N_2703);
nand U3094 (N_3094,N_2871,N_2811);
or U3095 (N_3095,N_2559,N_2502);
nor U3096 (N_3096,N_2909,N_2817);
nor U3097 (N_3097,N_2796,N_2976);
nand U3098 (N_3098,N_2981,N_2858);
and U3099 (N_3099,N_2860,N_2738);
nor U3100 (N_3100,N_2582,N_2519);
nand U3101 (N_3101,N_2743,N_2841);
nor U3102 (N_3102,N_2973,N_2830);
and U3103 (N_3103,N_2787,N_2594);
xor U3104 (N_3104,N_2575,N_2785);
nand U3105 (N_3105,N_2634,N_2760);
and U3106 (N_3106,N_2958,N_2955);
nor U3107 (N_3107,N_2657,N_2987);
and U3108 (N_3108,N_2640,N_2777);
nor U3109 (N_3109,N_2735,N_2515);
and U3110 (N_3110,N_2956,N_2966);
nand U3111 (N_3111,N_2525,N_2549);
nand U3112 (N_3112,N_2950,N_2619);
nand U3113 (N_3113,N_2583,N_2763);
and U3114 (N_3114,N_2576,N_2916);
nor U3115 (N_3115,N_2992,N_2754);
or U3116 (N_3116,N_2745,N_2947);
and U3117 (N_3117,N_2625,N_2577);
nor U3118 (N_3118,N_2808,N_2797);
and U3119 (N_3119,N_2773,N_2639);
or U3120 (N_3120,N_2920,N_2802);
or U3121 (N_3121,N_2688,N_2846);
nor U3122 (N_3122,N_2751,N_2762);
nand U3123 (N_3123,N_2605,N_2627);
and U3124 (N_3124,N_2874,N_2967);
and U3125 (N_3125,N_2755,N_2544);
nand U3126 (N_3126,N_2828,N_2836);
or U3127 (N_3127,N_2591,N_2849);
nand U3128 (N_3128,N_2614,N_2819);
nor U3129 (N_3129,N_2560,N_2631);
and U3130 (N_3130,N_2512,N_2501);
nand U3131 (N_3131,N_2682,N_2963);
nor U3132 (N_3132,N_2505,N_2944);
nand U3133 (N_3133,N_2658,N_2630);
nor U3134 (N_3134,N_2766,N_2563);
nand U3135 (N_3135,N_2641,N_2686);
and U3136 (N_3136,N_2704,N_2998);
nor U3137 (N_3137,N_2953,N_2783);
xor U3138 (N_3138,N_2500,N_2606);
and U3139 (N_3139,N_2919,N_2789);
nor U3140 (N_3140,N_2842,N_2761);
nor U3141 (N_3141,N_2603,N_2579);
nand U3142 (N_3142,N_2522,N_2628);
and U3143 (N_3143,N_2914,N_2611);
nor U3144 (N_3144,N_2573,N_2540);
and U3145 (N_3145,N_2542,N_2694);
or U3146 (N_3146,N_2677,N_2799);
and U3147 (N_3147,N_2881,N_2637);
and U3148 (N_3148,N_2668,N_2730);
nor U3149 (N_3149,N_2654,N_2536);
nor U3150 (N_3150,N_2626,N_2566);
nand U3151 (N_3151,N_2617,N_2555);
nor U3152 (N_3152,N_2527,N_2601);
or U3153 (N_3153,N_2810,N_2712);
and U3154 (N_3154,N_2962,N_2826);
nor U3155 (N_3155,N_2894,N_2720);
and U3156 (N_3156,N_2794,N_2674);
or U3157 (N_3157,N_2604,N_2721);
nor U3158 (N_3158,N_2526,N_2814);
or U3159 (N_3159,N_2595,N_2839);
or U3160 (N_3160,N_2622,N_2701);
nand U3161 (N_3161,N_2934,N_2584);
nand U3162 (N_3162,N_2647,N_2923);
and U3163 (N_3163,N_2918,N_2740);
or U3164 (N_3164,N_2600,N_2854);
nor U3165 (N_3165,N_2977,N_2827);
and U3166 (N_3166,N_2803,N_2561);
nand U3167 (N_3167,N_2568,N_2983);
nor U3168 (N_3168,N_2883,N_2695);
and U3169 (N_3169,N_2921,N_2734);
or U3170 (N_3170,N_2539,N_2507);
and U3171 (N_3171,N_2972,N_2518);
and U3172 (N_3172,N_2572,N_2567);
nand U3173 (N_3173,N_2719,N_2664);
and U3174 (N_3174,N_2774,N_2581);
and U3175 (N_3175,N_2899,N_2859);
and U3176 (N_3176,N_2633,N_2509);
or U3177 (N_3177,N_2856,N_2537);
nor U3178 (N_3178,N_2700,N_2746);
and U3179 (N_3179,N_2952,N_2925);
or U3180 (N_3180,N_2557,N_2911);
or U3181 (N_3181,N_2570,N_2532);
nand U3182 (N_3182,N_2748,N_2908);
nand U3183 (N_3183,N_2716,N_2553);
or U3184 (N_3184,N_2845,N_2864);
nand U3185 (N_3185,N_2960,N_2663);
nor U3186 (N_3186,N_2565,N_2708);
or U3187 (N_3187,N_2772,N_2905);
and U3188 (N_3188,N_2732,N_2957);
and U3189 (N_3189,N_2959,N_2940);
and U3190 (N_3190,N_2726,N_2961);
nor U3191 (N_3191,N_2684,N_2964);
nand U3192 (N_3192,N_2780,N_2757);
nand U3193 (N_3193,N_2547,N_2599);
or U3194 (N_3194,N_2965,N_2823);
or U3195 (N_3195,N_2511,N_2851);
and U3196 (N_3196,N_2993,N_2578);
xor U3197 (N_3197,N_2711,N_2791);
nor U3198 (N_3198,N_2756,N_2552);
nor U3199 (N_3199,N_2813,N_2890);
nor U3200 (N_3200,N_2818,N_2702);
xor U3201 (N_3201,N_2788,N_2643);
and U3202 (N_3202,N_2821,N_2752);
nor U3203 (N_3203,N_2590,N_2670);
nand U3204 (N_3204,N_2837,N_2520);
or U3205 (N_3205,N_2660,N_2545);
nor U3206 (N_3206,N_2924,N_2862);
or U3207 (N_3207,N_2907,N_2949);
nand U3208 (N_3208,N_2623,N_2731);
nand U3209 (N_3209,N_2784,N_2620);
nor U3210 (N_3210,N_2504,N_2974);
and U3211 (N_3211,N_2896,N_2885);
nand U3212 (N_3212,N_2683,N_2932);
and U3213 (N_3213,N_2685,N_2739);
and U3214 (N_3214,N_2942,N_2876);
and U3215 (N_3215,N_2825,N_2882);
nor U3216 (N_3216,N_2699,N_2678);
and U3217 (N_3217,N_2945,N_2927);
nor U3218 (N_3218,N_2875,N_2985);
nor U3219 (N_3219,N_2698,N_2838);
nor U3220 (N_3220,N_2672,N_2690);
nor U3221 (N_3221,N_2999,N_2725);
and U3222 (N_3222,N_2865,N_2895);
nand U3223 (N_3223,N_2863,N_2728);
nor U3224 (N_3224,N_2618,N_2765);
nor U3225 (N_3225,N_2671,N_2879);
nor U3226 (N_3226,N_2652,N_2648);
nand U3227 (N_3227,N_2870,N_2715);
and U3228 (N_3228,N_2889,N_2933);
and U3229 (N_3229,N_2521,N_2650);
and U3230 (N_3230,N_2551,N_2569);
nand U3231 (N_3231,N_2831,N_2893);
nand U3232 (N_3232,N_2621,N_2741);
nand U3233 (N_3233,N_2822,N_2524);
or U3234 (N_3234,N_2632,N_2795);
or U3235 (N_3235,N_2922,N_2653);
nor U3236 (N_3236,N_2666,N_2872);
nor U3237 (N_3237,N_2649,N_2661);
and U3238 (N_3238,N_2855,N_2954);
and U3239 (N_3239,N_2529,N_2609);
or U3240 (N_3240,N_2706,N_2659);
nor U3241 (N_3241,N_2847,N_2538);
or U3242 (N_3242,N_2996,N_2534);
xor U3243 (N_3243,N_2809,N_2775);
nor U3244 (N_3244,N_2888,N_2612);
or U3245 (N_3245,N_2655,N_2718);
nor U3246 (N_3246,N_2580,N_2714);
nand U3247 (N_3247,N_2970,N_2941);
and U3248 (N_3248,N_2523,N_2528);
nand U3249 (N_3249,N_2517,N_2930);
nand U3250 (N_3250,N_2520,N_2672);
or U3251 (N_3251,N_2965,N_2926);
or U3252 (N_3252,N_2921,N_2672);
nand U3253 (N_3253,N_2634,N_2882);
nand U3254 (N_3254,N_2504,N_2522);
or U3255 (N_3255,N_2878,N_2782);
and U3256 (N_3256,N_2946,N_2734);
and U3257 (N_3257,N_2912,N_2919);
nor U3258 (N_3258,N_2971,N_2716);
nand U3259 (N_3259,N_2930,N_2512);
nand U3260 (N_3260,N_2681,N_2748);
and U3261 (N_3261,N_2971,N_2607);
nand U3262 (N_3262,N_2553,N_2712);
nor U3263 (N_3263,N_2801,N_2891);
nor U3264 (N_3264,N_2714,N_2948);
nor U3265 (N_3265,N_2701,N_2510);
nor U3266 (N_3266,N_2882,N_2717);
and U3267 (N_3267,N_2523,N_2816);
and U3268 (N_3268,N_2851,N_2634);
or U3269 (N_3269,N_2947,N_2660);
and U3270 (N_3270,N_2773,N_2838);
and U3271 (N_3271,N_2758,N_2933);
nor U3272 (N_3272,N_2945,N_2595);
and U3273 (N_3273,N_2830,N_2707);
nand U3274 (N_3274,N_2917,N_2896);
nand U3275 (N_3275,N_2885,N_2521);
nor U3276 (N_3276,N_2952,N_2767);
nor U3277 (N_3277,N_2954,N_2546);
nor U3278 (N_3278,N_2898,N_2795);
nor U3279 (N_3279,N_2888,N_2526);
and U3280 (N_3280,N_2531,N_2996);
or U3281 (N_3281,N_2596,N_2541);
or U3282 (N_3282,N_2509,N_2835);
or U3283 (N_3283,N_2854,N_2653);
nand U3284 (N_3284,N_2551,N_2663);
nor U3285 (N_3285,N_2530,N_2779);
nand U3286 (N_3286,N_2639,N_2953);
and U3287 (N_3287,N_2782,N_2661);
and U3288 (N_3288,N_2879,N_2512);
and U3289 (N_3289,N_2598,N_2813);
and U3290 (N_3290,N_2772,N_2588);
or U3291 (N_3291,N_2761,N_2784);
and U3292 (N_3292,N_2737,N_2855);
nand U3293 (N_3293,N_2720,N_2793);
nand U3294 (N_3294,N_2828,N_2965);
nand U3295 (N_3295,N_2744,N_2733);
nor U3296 (N_3296,N_2656,N_2790);
or U3297 (N_3297,N_2666,N_2553);
nor U3298 (N_3298,N_2819,N_2654);
nor U3299 (N_3299,N_2587,N_2725);
or U3300 (N_3300,N_2695,N_2567);
or U3301 (N_3301,N_2957,N_2935);
nand U3302 (N_3302,N_2915,N_2957);
nand U3303 (N_3303,N_2628,N_2721);
or U3304 (N_3304,N_2955,N_2524);
or U3305 (N_3305,N_2921,N_2951);
and U3306 (N_3306,N_2647,N_2541);
nor U3307 (N_3307,N_2848,N_2794);
nor U3308 (N_3308,N_2841,N_2948);
nor U3309 (N_3309,N_2994,N_2517);
or U3310 (N_3310,N_2604,N_2827);
xnor U3311 (N_3311,N_2616,N_2572);
nand U3312 (N_3312,N_2886,N_2623);
nor U3313 (N_3313,N_2558,N_2574);
and U3314 (N_3314,N_2584,N_2785);
nor U3315 (N_3315,N_2557,N_2754);
and U3316 (N_3316,N_2556,N_2817);
or U3317 (N_3317,N_2648,N_2782);
or U3318 (N_3318,N_2595,N_2648);
or U3319 (N_3319,N_2576,N_2861);
nand U3320 (N_3320,N_2973,N_2951);
nand U3321 (N_3321,N_2837,N_2853);
xor U3322 (N_3322,N_2988,N_2816);
or U3323 (N_3323,N_2994,N_2698);
nor U3324 (N_3324,N_2500,N_2922);
and U3325 (N_3325,N_2798,N_2932);
nor U3326 (N_3326,N_2705,N_2977);
or U3327 (N_3327,N_2707,N_2658);
nand U3328 (N_3328,N_2678,N_2816);
nor U3329 (N_3329,N_2901,N_2518);
or U3330 (N_3330,N_2670,N_2897);
and U3331 (N_3331,N_2917,N_2994);
nand U3332 (N_3332,N_2582,N_2984);
nand U3333 (N_3333,N_2708,N_2624);
nand U3334 (N_3334,N_2952,N_2582);
or U3335 (N_3335,N_2763,N_2639);
and U3336 (N_3336,N_2741,N_2721);
and U3337 (N_3337,N_2980,N_2621);
or U3338 (N_3338,N_2978,N_2699);
or U3339 (N_3339,N_2610,N_2868);
or U3340 (N_3340,N_2711,N_2586);
and U3341 (N_3341,N_2901,N_2779);
or U3342 (N_3342,N_2517,N_2601);
xor U3343 (N_3343,N_2683,N_2951);
nand U3344 (N_3344,N_2744,N_2936);
nand U3345 (N_3345,N_2751,N_2942);
and U3346 (N_3346,N_2738,N_2907);
or U3347 (N_3347,N_2625,N_2803);
nor U3348 (N_3348,N_2843,N_2555);
and U3349 (N_3349,N_2957,N_2595);
and U3350 (N_3350,N_2573,N_2511);
or U3351 (N_3351,N_2501,N_2588);
nand U3352 (N_3352,N_2869,N_2933);
nor U3353 (N_3353,N_2652,N_2635);
and U3354 (N_3354,N_2759,N_2913);
or U3355 (N_3355,N_2767,N_2768);
nor U3356 (N_3356,N_2614,N_2608);
and U3357 (N_3357,N_2686,N_2588);
nand U3358 (N_3358,N_2694,N_2570);
and U3359 (N_3359,N_2876,N_2667);
and U3360 (N_3360,N_2681,N_2853);
xnor U3361 (N_3361,N_2627,N_2696);
and U3362 (N_3362,N_2547,N_2658);
nor U3363 (N_3363,N_2566,N_2575);
and U3364 (N_3364,N_2676,N_2761);
nor U3365 (N_3365,N_2865,N_2679);
or U3366 (N_3366,N_2892,N_2543);
nand U3367 (N_3367,N_2606,N_2748);
and U3368 (N_3368,N_2810,N_2924);
or U3369 (N_3369,N_2575,N_2747);
and U3370 (N_3370,N_2818,N_2517);
nand U3371 (N_3371,N_2817,N_2583);
nor U3372 (N_3372,N_2655,N_2703);
nor U3373 (N_3373,N_2643,N_2507);
nand U3374 (N_3374,N_2812,N_2582);
nor U3375 (N_3375,N_2911,N_2718);
and U3376 (N_3376,N_2544,N_2937);
or U3377 (N_3377,N_2602,N_2700);
or U3378 (N_3378,N_2961,N_2851);
or U3379 (N_3379,N_2705,N_2682);
and U3380 (N_3380,N_2903,N_2631);
and U3381 (N_3381,N_2917,N_2651);
or U3382 (N_3382,N_2967,N_2902);
nand U3383 (N_3383,N_2541,N_2876);
or U3384 (N_3384,N_2954,N_2836);
and U3385 (N_3385,N_2593,N_2637);
nor U3386 (N_3386,N_2572,N_2610);
or U3387 (N_3387,N_2650,N_2902);
nor U3388 (N_3388,N_2948,N_2626);
nand U3389 (N_3389,N_2678,N_2547);
and U3390 (N_3390,N_2794,N_2578);
or U3391 (N_3391,N_2713,N_2932);
or U3392 (N_3392,N_2877,N_2756);
nor U3393 (N_3393,N_2765,N_2966);
or U3394 (N_3394,N_2692,N_2796);
or U3395 (N_3395,N_2548,N_2933);
or U3396 (N_3396,N_2635,N_2533);
or U3397 (N_3397,N_2999,N_2717);
or U3398 (N_3398,N_2640,N_2507);
nor U3399 (N_3399,N_2967,N_2932);
and U3400 (N_3400,N_2952,N_2694);
or U3401 (N_3401,N_2875,N_2822);
nand U3402 (N_3402,N_2566,N_2615);
or U3403 (N_3403,N_2714,N_2983);
and U3404 (N_3404,N_2837,N_2508);
nand U3405 (N_3405,N_2733,N_2838);
nand U3406 (N_3406,N_2534,N_2542);
nand U3407 (N_3407,N_2593,N_2943);
and U3408 (N_3408,N_2583,N_2637);
or U3409 (N_3409,N_2673,N_2827);
and U3410 (N_3410,N_2512,N_2614);
nand U3411 (N_3411,N_2740,N_2886);
or U3412 (N_3412,N_2914,N_2680);
or U3413 (N_3413,N_2549,N_2521);
or U3414 (N_3414,N_2711,N_2780);
and U3415 (N_3415,N_2884,N_2538);
and U3416 (N_3416,N_2518,N_2994);
nor U3417 (N_3417,N_2542,N_2934);
and U3418 (N_3418,N_2764,N_2539);
and U3419 (N_3419,N_2763,N_2784);
or U3420 (N_3420,N_2839,N_2812);
or U3421 (N_3421,N_2777,N_2825);
and U3422 (N_3422,N_2892,N_2926);
nand U3423 (N_3423,N_2967,N_2656);
nor U3424 (N_3424,N_2537,N_2773);
and U3425 (N_3425,N_2661,N_2982);
nor U3426 (N_3426,N_2709,N_2908);
nor U3427 (N_3427,N_2515,N_2847);
or U3428 (N_3428,N_2824,N_2680);
nor U3429 (N_3429,N_2579,N_2978);
nand U3430 (N_3430,N_2522,N_2781);
nor U3431 (N_3431,N_2829,N_2529);
and U3432 (N_3432,N_2668,N_2705);
nand U3433 (N_3433,N_2557,N_2778);
or U3434 (N_3434,N_2671,N_2951);
or U3435 (N_3435,N_2563,N_2874);
or U3436 (N_3436,N_2927,N_2502);
nand U3437 (N_3437,N_2561,N_2980);
nor U3438 (N_3438,N_2504,N_2970);
and U3439 (N_3439,N_2862,N_2855);
or U3440 (N_3440,N_2834,N_2601);
or U3441 (N_3441,N_2662,N_2535);
xor U3442 (N_3442,N_2880,N_2602);
nor U3443 (N_3443,N_2710,N_2938);
or U3444 (N_3444,N_2510,N_2695);
nand U3445 (N_3445,N_2649,N_2563);
or U3446 (N_3446,N_2609,N_2508);
nor U3447 (N_3447,N_2879,N_2574);
nand U3448 (N_3448,N_2820,N_2845);
nor U3449 (N_3449,N_2588,N_2798);
and U3450 (N_3450,N_2770,N_2960);
and U3451 (N_3451,N_2627,N_2821);
nand U3452 (N_3452,N_2874,N_2859);
nand U3453 (N_3453,N_2684,N_2611);
or U3454 (N_3454,N_2688,N_2538);
or U3455 (N_3455,N_2909,N_2615);
or U3456 (N_3456,N_2918,N_2855);
xor U3457 (N_3457,N_2579,N_2583);
and U3458 (N_3458,N_2530,N_2880);
and U3459 (N_3459,N_2825,N_2673);
nand U3460 (N_3460,N_2924,N_2910);
nand U3461 (N_3461,N_2775,N_2935);
nor U3462 (N_3462,N_2838,N_2795);
or U3463 (N_3463,N_2749,N_2898);
nand U3464 (N_3464,N_2588,N_2759);
nor U3465 (N_3465,N_2628,N_2624);
nor U3466 (N_3466,N_2945,N_2602);
nand U3467 (N_3467,N_2537,N_2859);
nand U3468 (N_3468,N_2896,N_2506);
nor U3469 (N_3469,N_2722,N_2937);
nand U3470 (N_3470,N_2738,N_2657);
nor U3471 (N_3471,N_2502,N_2826);
and U3472 (N_3472,N_2803,N_2565);
and U3473 (N_3473,N_2641,N_2783);
nor U3474 (N_3474,N_2816,N_2712);
nor U3475 (N_3475,N_2859,N_2614);
nor U3476 (N_3476,N_2794,N_2613);
nand U3477 (N_3477,N_2520,N_2696);
and U3478 (N_3478,N_2719,N_2695);
nor U3479 (N_3479,N_2667,N_2707);
nor U3480 (N_3480,N_2511,N_2568);
nand U3481 (N_3481,N_2677,N_2899);
nor U3482 (N_3482,N_2634,N_2759);
or U3483 (N_3483,N_2734,N_2612);
and U3484 (N_3484,N_2500,N_2643);
or U3485 (N_3485,N_2561,N_2697);
and U3486 (N_3486,N_2709,N_2876);
nand U3487 (N_3487,N_2685,N_2611);
or U3488 (N_3488,N_2868,N_2541);
or U3489 (N_3489,N_2990,N_2806);
and U3490 (N_3490,N_2579,N_2591);
nand U3491 (N_3491,N_2740,N_2614);
and U3492 (N_3492,N_2820,N_2544);
nand U3493 (N_3493,N_2887,N_2959);
and U3494 (N_3494,N_2594,N_2940);
nor U3495 (N_3495,N_2766,N_2545);
nor U3496 (N_3496,N_2808,N_2633);
nor U3497 (N_3497,N_2842,N_2937);
and U3498 (N_3498,N_2806,N_2861);
or U3499 (N_3499,N_2679,N_2880);
or U3500 (N_3500,N_3124,N_3451);
or U3501 (N_3501,N_3210,N_3417);
nand U3502 (N_3502,N_3020,N_3479);
and U3503 (N_3503,N_3302,N_3033);
and U3504 (N_3504,N_3461,N_3038);
nand U3505 (N_3505,N_3359,N_3392);
nor U3506 (N_3506,N_3364,N_3162);
nand U3507 (N_3507,N_3036,N_3045);
nand U3508 (N_3508,N_3431,N_3012);
nor U3509 (N_3509,N_3254,N_3197);
nor U3510 (N_3510,N_3488,N_3151);
nand U3511 (N_3511,N_3326,N_3433);
or U3512 (N_3512,N_3329,N_3126);
or U3513 (N_3513,N_3063,N_3094);
nand U3514 (N_3514,N_3410,N_3444);
nand U3515 (N_3515,N_3145,N_3498);
and U3516 (N_3516,N_3131,N_3374);
nand U3517 (N_3517,N_3196,N_3277);
and U3518 (N_3518,N_3005,N_3436);
nand U3519 (N_3519,N_3096,N_3270);
or U3520 (N_3520,N_3032,N_3158);
or U3521 (N_3521,N_3052,N_3076);
and U3522 (N_3522,N_3089,N_3297);
xnor U3523 (N_3523,N_3017,N_3071);
nor U3524 (N_3524,N_3135,N_3120);
or U3525 (N_3525,N_3305,N_3116);
nor U3526 (N_3526,N_3260,N_3328);
nand U3527 (N_3527,N_3007,N_3073);
nand U3528 (N_3528,N_3100,N_3293);
nand U3529 (N_3529,N_3405,N_3109);
and U3530 (N_3530,N_3320,N_3291);
nand U3531 (N_3531,N_3455,N_3236);
or U3532 (N_3532,N_3138,N_3221);
or U3533 (N_3533,N_3230,N_3044);
or U3534 (N_3534,N_3435,N_3106);
nor U3535 (N_3535,N_3478,N_3189);
nand U3536 (N_3536,N_3251,N_3027);
and U3537 (N_3537,N_3030,N_3396);
and U3538 (N_3538,N_3264,N_3213);
nand U3539 (N_3539,N_3003,N_3415);
or U3540 (N_3540,N_3467,N_3039);
nand U3541 (N_3541,N_3341,N_3241);
nor U3542 (N_3542,N_3295,N_3304);
and U3543 (N_3543,N_3091,N_3049);
nand U3544 (N_3544,N_3041,N_3307);
or U3545 (N_3545,N_3087,N_3011);
or U3546 (N_3546,N_3015,N_3407);
nand U3547 (N_3547,N_3119,N_3220);
and U3548 (N_3548,N_3406,N_3029);
nor U3549 (N_3549,N_3425,N_3292);
nor U3550 (N_3550,N_3460,N_3025);
and U3551 (N_3551,N_3393,N_3153);
and U3552 (N_3552,N_3483,N_3466);
and U3553 (N_3553,N_3043,N_3022);
or U3554 (N_3554,N_3303,N_3084);
nor U3555 (N_3555,N_3101,N_3112);
or U3556 (N_3556,N_3016,N_3265);
xnor U3557 (N_3557,N_3110,N_3399);
and U3558 (N_3558,N_3285,N_3249);
nand U3559 (N_3559,N_3137,N_3200);
or U3560 (N_3560,N_3459,N_3177);
xor U3561 (N_3561,N_3170,N_3141);
and U3562 (N_3562,N_3456,N_3227);
and U3563 (N_3563,N_3000,N_3372);
and U3564 (N_3564,N_3256,N_3178);
nor U3565 (N_3565,N_3412,N_3118);
nor U3566 (N_3566,N_3057,N_3385);
nand U3567 (N_3567,N_3055,N_3376);
and U3568 (N_3568,N_3259,N_3133);
or U3569 (N_3569,N_3381,N_3093);
or U3570 (N_3570,N_3186,N_3275);
nand U3571 (N_3571,N_3075,N_3490);
and U3572 (N_3572,N_3185,N_3179);
or U3573 (N_3573,N_3064,N_3199);
or U3574 (N_3574,N_3050,N_3365);
nand U3575 (N_3575,N_3095,N_3155);
nand U3576 (N_3576,N_3484,N_3319);
or U3577 (N_3577,N_3438,N_3062);
nand U3578 (N_3578,N_3281,N_3008);
or U3579 (N_3579,N_3114,N_3493);
nor U3580 (N_3580,N_3477,N_3378);
nor U3581 (N_3581,N_3345,N_3487);
nor U3582 (N_3582,N_3351,N_3327);
or U3583 (N_3583,N_3115,N_3318);
and U3584 (N_3584,N_3497,N_3492);
and U3585 (N_3585,N_3248,N_3072);
and U3586 (N_3586,N_3289,N_3111);
or U3587 (N_3587,N_3004,N_3382);
nand U3588 (N_3588,N_3325,N_3139);
nand U3589 (N_3589,N_3054,N_3391);
and U3590 (N_3590,N_3413,N_3229);
and U3591 (N_3591,N_3010,N_3343);
nand U3592 (N_3592,N_3102,N_3383);
or U3593 (N_3593,N_3489,N_3469);
or U3594 (N_3594,N_3334,N_3163);
or U3595 (N_3595,N_3006,N_3166);
nor U3596 (N_3596,N_3463,N_3122);
and U3597 (N_3597,N_3395,N_3360);
nor U3598 (N_3598,N_3280,N_3387);
or U3599 (N_3599,N_3182,N_3184);
nand U3600 (N_3600,N_3068,N_3198);
nor U3601 (N_3601,N_3272,N_3400);
nor U3602 (N_3602,N_3268,N_3140);
or U3603 (N_3603,N_3338,N_3299);
or U3604 (N_3604,N_3380,N_3428);
nor U3605 (N_3605,N_3384,N_3028);
and U3606 (N_3606,N_3283,N_3352);
nand U3607 (N_3607,N_3085,N_3188);
or U3608 (N_3608,N_3098,N_3271);
nand U3609 (N_3609,N_3389,N_3083);
nor U3610 (N_3610,N_3361,N_3247);
or U3611 (N_3611,N_3430,N_3202);
nor U3612 (N_3612,N_3205,N_3214);
nor U3613 (N_3613,N_3201,N_3279);
or U3614 (N_3614,N_3146,N_3239);
nor U3615 (N_3615,N_3237,N_3276);
and U3616 (N_3616,N_3437,N_3123);
nor U3617 (N_3617,N_3315,N_3287);
and U3618 (N_3618,N_3401,N_3058);
and U3619 (N_3619,N_3342,N_3423);
and U3620 (N_3620,N_3224,N_3377);
and U3621 (N_3621,N_3117,N_3161);
and U3622 (N_3622,N_3077,N_3426);
xor U3623 (N_3623,N_3298,N_3448);
and U3624 (N_3624,N_3215,N_3132);
nand U3625 (N_3625,N_3313,N_3231);
or U3626 (N_3626,N_3445,N_3160);
or U3627 (N_3627,N_3499,N_3009);
and U3628 (N_3628,N_3422,N_3240);
and U3629 (N_3629,N_3261,N_3193);
and U3630 (N_3630,N_3209,N_3099);
and U3631 (N_3631,N_3223,N_3147);
nand U3632 (N_3632,N_3403,N_3103);
or U3633 (N_3633,N_3250,N_3439);
and U3634 (N_3634,N_3286,N_3144);
and U3635 (N_3635,N_3127,N_3398);
and U3636 (N_3636,N_3217,N_3226);
and U3637 (N_3637,N_3150,N_3421);
or U3638 (N_3638,N_3294,N_3397);
nor U3639 (N_3639,N_3440,N_3424);
nor U3640 (N_3640,N_3154,N_3243);
nor U3641 (N_3641,N_3252,N_3157);
xor U3642 (N_3642,N_3346,N_3024);
or U3643 (N_3643,N_3092,N_3457);
nand U3644 (N_3644,N_3037,N_3404);
or U3645 (N_3645,N_3324,N_3206);
nand U3646 (N_3646,N_3233,N_3362);
and U3647 (N_3647,N_3255,N_3207);
xor U3648 (N_3648,N_3034,N_3330);
nor U3649 (N_3649,N_3339,N_3308);
xor U3650 (N_3650,N_3253,N_3462);
or U3651 (N_3651,N_3486,N_3290);
or U3652 (N_3652,N_3273,N_3317);
and U3653 (N_3653,N_3482,N_3323);
nand U3654 (N_3654,N_3332,N_3427);
xor U3655 (N_3655,N_3187,N_3344);
and U3656 (N_3656,N_3067,N_3473);
nand U3657 (N_3657,N_3368,N_3059);
or U3658 (N_3658,N_3322,N_3061);
and U3659 (N_3659,N_3419,N_3056);
nor U3660 (N_3660,N_3136,N_3105);
and U3661 (N_3661,N_3066,N_3171);
and U3662 (N_3662,N_3386,N_3356);
nor U3663 (N_3663,N_3078,N_3104);
and U3664 (N_3664,N_3375,N_3447);
or U3665 (N_3665,N_3080,N_3195);
or U3666 (N_3666,N_3065,N_3454);
or U3667 (N_3667,N_3296,N_3165);
and U3668 (N_3668,N_3367,N_3042);
or U3669 (N_3669,N_3358,N_3432);
or U3670 (N_3670,N_3107,N_3300);
and U3671 (N_3671,N_3495,N_3468);
nor U3672 (N_3672,N_3194,N_3046);
or U3673 (N_3673,N_3494,N_3449);
nor U3674 (N_3674,N_3347,N_3465);
nand U3675 (N_3675,N_3174,N_3013);
nor U3676 (N_3676,N_3169,N_3242);
or U3677 (N_3677,N_3191,N_3336);
or U3678 (N_3678,N_3369,N_3245);
and U3679 (N_3679,N_3018,N_3409);
nand U3680 (N_3680,N_3121,N_3232);
nor U3681 (N_3681,N_3216,N_3402);
or U3682 (N_3682,N_3314,N_3167);
nand U3683 (N_3683,N_3159,N_3014);
nand U3684 (N_3684,N_3208,N_3321);
or U3685 (N_3685,N_3443,N_3176);
nor U3686 (N_3686,N_3371,N_3051);
and U3687 (N_3687,N_3394,N_3446);
nand U3688 (N_3688,N_3458,N_3074);
nor U3689 (N_3689,N_3001,N_3235);
and U3690 (N_3690,N_3262,N_3354);
xor U3691 (N_3691,N_3258,N_3349);
and U3692 (N_3692,N_3306,N_3337);
nor U3693 (N_3693,N_3048,N_3238);
and U3694 (N_3694,N_3472,N_3274);
xor U3695 (N_3695,N_3244,N_3225);
nand U3696 (N_3696,N_3450,N_3370);
nand U3697 (N_3697,N_3464,N_3481);
or U3698 (N_3698,N_3353,N_3496);
nor U3699 (N_3699,N_3416,N_3379);
or U3700 (N_3700,N_3366,N_3434);
nor U3701 (N_3701,N_3388,N_3418);
nand U3702 (N_3702,N_3002,N_3088);
or U3703 (N_3703,N_3278,N_3181);
nor U3704 (N_3704,N_3129,N_3453);
nor U3705 (N_3705,N_3452,N_3282);
and U3706 (N_3706,N_3152,N_3125);
nor U3707 (N_3707,N_3190,N_3470);
and U3708 (N_3708,N_3333,N_3168);
and U3709 (N_3709,N_3491,N_3228);
nand U3710 (N_3710,N_3480,N_3309);
or U3711 (N_3711,N_3173,N_3090);
nor U3712 (N_3712,N_3355,N_3390);
nand U3713 (N_3713,N_3203,N_3476);
nand U3714 (N_3714,N_3211,N_3474);
nand U3715 (N_3715,N_3442,N_3429);
nor U3716 (N_3716,N_3301,N_3149);
nand U3717 (N_3717,N_3097,N_3053);
and U3718 (N_3718,N_3021,N_3234);
nor U3719 (N_3719,N_3081,N_3172);
nand U3720 (N_3720,N_3218,N_3411);
nand U3721 (N_3721,N_3180,N_3079);
and U3722 (N_3722,N_3257,N_3373);
or U3723 (N_3723,N_3284,N_3363);
and U3724 (N_3724,N_3212,N_3164);
nor U3725 (N_3725,N_3113,N_3023);
nor U3726 (N_3726,N_3263,N_3035);
and U3727 (N_3727,N_3143,N_3156);
and U3728 (N_3728,N_3267,N_3420);
nand U3729 (N_3729,N_3031,N_3148);
and U3730 (N_3730,N_3414,N_3288);
or U3731 (N_3731,N_3475,N_3269);
nand U3732 (N_3732,N_3219,N_3086);
nand U3733 (N_3733,N_3060,N_3175);
nand U3734 (N_3734,N_3082,N_3441);
nand U3735 (N_3735,N_3070,N_3204);
nand U3736 (N_3736,N_3142,N_3357);
or U3737 (N_3737,N_3340,N_3350);
or U3738 (N_3738,N_3108,N_3040);
or U3739 (N_3739,N_3130,N_3331);
and U3740 (N_3740,N_3348,N_3310);
and U3741 (N_3741,N_3266,N_3128);
nor U3742 (N_3742,N_3471,N_3019);
and U3743 (N_3743,N_3335,N_3183);
and U3744 (N_3744,N_3192,N_3222);
nand U3745 (N_3745,N_3408,N_3246);
nor U3746 (N_3746,N_3047,N_3069);
and U3747 (N_3747,N_3026,N_3134);
nand U3748 (N_3748,N_3312,N_3311);
or U3749 (N_3749,N_3485,N_3316);
nand U3750 (N_3750,N_3449,N_3329);
and U3751 (N_3751,N_3020,N_3098);
nand U3752 (N_3752,N_3326,N_3419);
and U3753 (N_3753,N_3291,N_3157);
or U3754 (N_3754,N_3255,N_3205);
nand U3755 (N_3755,N_3483,N_3351);
and U3756 (N_3756,N_3389,N_3111);
or U3757 (N_3757,N_3092,N_3375);
nand U3758 (N_3758,N_3204,N_3423);
or U3759 (N_3759,N_3245,N_3151);
or U3760 (N_3760,N_3428,N_3158);
nand U3761 (N_3761,N_3130,N_3023);
nand U3762 (N_3762,N_3037,N_3381);
nor U3763 (N_3763,N_3359,N_3253);
nand U3764 (N_3764,N_3002,N_3316);
and U3765 (N_3765,N_3162,N_3271);
or U3766 (N_3766,N_3240,N_3030);
nor U3767 (N_3767,N_3261,N_3424);
and U3768 (N_3768,N_3297,N_3094);
nand U3769 (N_3769,N_3251,N_3441);
nand U3770 (N_3770,N_3105,N_3435);
nand U3771 (N_3771,N_3483,N_3309);
and U3772 (N_3772,N_3367,N_3376);
nand U3773 (N_3773,N_3356,N_3057);
nand U3774 (N_3774,N_3096,N_3192);
or U3775 (N_3775,N_3472,N_3461);
or U3776 (N_3776,N_3182,N_3056);
or U3777 (N_3777,N_3089,N_3453);
nor U3778 (N_3778,N_3330,N_3362);
or U3779 (N_3779,N_3331,N_3283);
and U3780 (N_3780,N_3382,N_3300);
or U3781 (N_3781,N_3022,N_3347);
nor U3782 (N_3782,N_3258,N_3221);
or U3783 (N_3783,N_3001,N_3439);
xnor U3784 (N_3784,N_3078,N_3004);
nand U3785 (N_3785,N_3295,N_3108);
nor U3786 (N_3786,N_3369,N_3340);
or U3787 (N_3787,N_3202,N_3180);
nor U3788 (N_3788,N_3194,N_3031);
and U3789 (N_3789,N_3024,N_3009);
nor U3790 (N_3790,N_3304,N_3182);
nand U3791 (N_3791,N_3010,N_3050);
nor U3792 (N_3792,N_3240,N_3079);
and U3793 (N_3793,N_3307,N_3227);
or U3794 (N_3794,N_3387,N_3388);
nor U3795 (N_3795,N_3334,N_3069);
xor U3796 (N_3796,N_3173,N_3369);
nor U3797 (N_3797,N_3102,N_3158);
and U3798 (N_3798,N_3337,N_3288);
or U3799 (N_3799,N_3259,N_3369);
nand U3800 (N_3800,N_3059,N_3450);
or U3801 (N_3801,N_3091,N_3374);
and U3802 (N_3802,N_3451,N_3012);
or U3803 (N_3803,N_3446,N_3216);
nor U3804 (N_3804,N_3114,N_3187);
xnor U3805 (N_3805,N_3413,N_3498);
nand U3806 (N_3806,N_3007,N_3267);
and U3807 (N_3807,N_3318,N_3460);
nor U3808 (N_3808,N_3371,N_3181);
nor U3809 (N_3809,N_3335,N_3369);
or U3810 (N_3810,N_3123,N_3039);
nand U3811 (N_3811,N_3095,N_3385);
nand U3812 (N_3812,N_3269,N_3430);
or U3813 (N_3813,N_3439,N_3428);
nor U3814 (N_3814,N_3143,N_3356);
and U3815 (N_3815,N_3022,N_3305);
and U3816 (N_3816,N_3135,N_3459);
nor U3817 (N_3817,N_3423,N_3144);
and U3818 (N_3818,N_3275,N_3401);
nor U3819 (N_3819,N_3012,N_3140);
or U3820 (N_3820,N_3270,N_3183);
and U3821 (N_3821,N_3248,N_3270);
nor U3822 (N_3822,N_3156,N_3408);
or U3823 (N_3823,N_3295,N_3076);
and U3824 (N_3824,N_3485,N_3197);
and U3825 (N_3825,N_3136,N_3484);
nor U3826 (N_3826,N_3307,N_3234);
xor U3827 (N_3827,N_3084,N_3457);
and U3828 (N_3828,N_3067,N_3359);
xor U3829 (N_3829,N_3277,N_3273);
or U3830 (N_3830,N_3126,N_3063);
nor U3831 (N_3831,N_3393,N_3018);
nand U3832 (N_3832,N_3228,N_3340);
xor U3833 (N_3833,N_3481,N_3204);
nand U3834 (N_3834,N_3379,N_3267);
and U3835 (N_3835,N_3159,N_3128);
nor U3836 (N_3836,N_3472,N_3483);
nor U3837 (N_3837,N_3490,N_3188);
and U3838 (N_3838,N_3093,N_3231);
nand U3839 (N_3839,N_3182,N_3376);
nor U3840 (N_3840,N_3140,N_3497);
nor U3841 (N_3841,N_3145,N_3221);
nand U3842 (N_3842,N_3401,N_3168);
nand U3843 (N_3843,N_3022,N_3361);
and U3844 (N_3844,N_3402,N_3437);
or U3845 (N_3845,N_3004,N_3085);
and U3846 (N_3846,N_3029,N_3089);
nand U3847 (N_3847,N_3260,N_3399);
nand U3848 (N_3848,N_3335,N_3427);
and U3849 (N_3849,N_3405,N_3116);
nand U3850 (N_3850,N_3212,N_3403);
nand U3851 (N_3851,N_3022,N_3316);
nand U3852 (N_3852,N_3250,N_3173);
nand U3853 (N_3853,N_3380,N_3044);
nor U3854 (N_3854,N_3480,N_3125);
and U3855 (N_3855,N_3103,N_3180);
nor U3856 (N_3856,N_3019,N_3415);
or U3857 (N_3857,N_3128,N_3107);
and U3858 (N_3858,N_3269,N_3012);
and U3859 (N_3859,N_3225,N_3432);
nor U3860 (N_3860,N_3420,N_3339);
nor U3861 (N_3861,N_3294,N_3290);
and U3862 (N_3862,N_3232,N_3066);
xnor U3863 (N_3863,N_3011,N_3153);
nand U3864 (N_3864,N_3454,N_3277);
nand U3865 (N_3865,N_3443,N_3217);
nand U3866 (N_3866,N_3345,N_3119);
and U3867 (N_3867,N_3101,N_3354);
and U3868 (N_3868,N_3146,N_3176);
xor U3869 (N_3869,N_3468,N_3303);
and U3870 (N_3870,N_3351,N_3478);
and U3871 (N_3871,N_3070,N_3012);
or U3872 (N_3872,N_3077,N_3319);
and U3873 (N_3873,N_3440,N_3173);
nand U3874 (N_3874,N_3349,N_3441);
nand U3875 (N_3875,N_3243,N_3120);
and U3876 (N_3876,N_3360,N_3210);
or U3877 (N_3877,N_3216,N_3489);
nor U3878 (N_3878,N_3232,N_3378);
and U3879 (N_3879,N_3376,N_3343);
nand U3880 (N_3880,N_3348,N_3398);
or U3881 (N_3881,N_3400,N_3121);
nor U3882 (N_3882,N_3463,N_3451);
and U3883 (N_3883,N_3492,N_3216);
nor U3884 (N_3884,N_3194,N_3230);
or U3885 (N_3885,N_3139,N_3309);
nor U3886 (N_3886,N_3495,N_3381);
nand U3887 (N_3887,N_3051,N_3077);
or U3888 (N_3888,N_3165,N_3338);
nand U3889 (N_3889,N_3172,N_3484);
nand U3890 (N_3890,N_3146,N_3333);
nor U3891 (N_3891,N_3050,N_3487);
and U3892 (N_3892,N_3158,N_3008);
or U3893 (N_3893,N_3059,N_3108);
nor U3894 (N_3894,N_3197,N_3320);
xnor U3895 (N_3895,N_3361,N_3104);
nor U3896 (N_3896,N_3035,N_3201);
or U3897 (N_3897,N_3366,N_3128);
nor U3898 (N_3898,N_3336,N_3430);
nor U3899 (N_3899,N_3054,N_3215);
nand U3900 (N_3900,N_3296,N_3267);
or U3901 (N_3901,N_3348,N_3487);
nand U3902 (N_3902,N_3047,N_3410);
or U3903 (N_3903,N_3089,N_3000);
and U3904 (N_3904,N_3328,N_3417);
and U3905 (N_3905,N_3283,N_3139);
and U3906 (N_3906,N_3114,N_3421);
nand U3907 (N_3907,N_3400,N_3476);
nor U3908 (N_3908,N_3127,N_3096);
and U3909 (N_3909,N_3291,N_3295);
or U3910 (N_3910,N_3285,N_3476);
and U3911 (N_3911,N_3249,N_3212);
and U3912 (N_3912,N_3498,N_3177);
or U3913 (N_3913,N_3175,N_3136);
nor U3914 (N_3914,N_3166,N_3259);
nand U3915 (N_3915,N_3167,N_3454);
and U3916 (N_3916,N_3040,N_3113);
nand U3917 (N_3917,N_3267,N_3386);
nor U3918 (N_3918,N_3072,N_3168);
and U3919 (N_3919,N_3296,N_3303);
nand U3920 (N_3920,N_3028,N_3314);
nand U3921 (N_3921,N_3124,N_3375);
nor U3922 (N_3922,N_3414,N_3029);
or U3923 (N_3923,N_3000,N_3401);
nor U3924 (N_3924,N_3193,N_3446);
or U3925 (N_3925,N_3395,N_3246);
or U3926 (N_3926,N_3232,N_3014);
nand U3927 (N_3927,N_3286,N_3412);
or U3928 (N_3928,N_3327,N_3216);
and U3929 (N_3929,N_3130,N_3493);
nor U3930 (N_3930,N_3079,N_3066);
nor U3931 (N_3931,N_3013,N_3078);
or U3932 (N_3932,N_3028,N_3083);
or U3933 (N_3933,N_3326,N_3165);
and U3934 (N_3934,N_3302,N_3431);
and U3935 (N_3935,N_3065,N_3037);
and U3936 (N_3936,N_3475,N_3384);
nand U3937 (N_3937,N_3496,N_3166);
or U3938 (N_3938,N_3309,N_3454);
nor U3939 (N_3939,N_3323,N_3407);
nand U3940 (N_3940,N_3066,N_3252);
nor U3941 (N_3941,N_3085,N_3087);
nand U3942 (N_3942,N_3091,N_3485);
or U3943 (N_3943,N_3297,N_3217);
xnor U3944 (N_3944,N_3302,N_3425);
and U3945 (N_3945,N_3403,N_3236);
or U3946 (N_3946,N_3023,N_3391);
nand U3947 (N_3947,N_3123,N_3088);
and U3948 (N_3948,N_3097,N_3050);
nand U3949 (N_3949,N_3227,N_3064);
and U3950 (N_3950,N_3096,N_3011);
and U3951 (N_3951,N_3441,N_3257);
and U3952 (N_3952,N_3096,N_3117);
nor U3953 (N_3953,N_3122,N_3335);
nor U3954 (N_3954,N_3485,N_3257);
xnor U3955 (N_3955,N_3320,N_3110);
or U3956 (N_3956,N_3073,N_3221);
nand U3957 (N_3957,N_3271,N_3409);
nor U3958 (N_3958,N_3122,N_3124);
or U3959 (N_3959,N_3181,N_3275);
or U3960 (N_3960,N_3263,N_3445);
or U3961 (N_3961,N_3170,N_3191);
and U3962 (N_3962,N_3470,N_3493);
nand U3963 (N_3963,N_3127,N_3481);
nand U3964 (N_3964,N_3204,N_3306);
nor U3965 (N_3965,N_3338,N_3013);
or U3966 (N_3966,N_3362,N_3426);
or U3967 (N_3967,N_3381,N_3389);
nor U3968 (N_3968,N_3221,N_3191);
and U3969 (N_3969,N_3415,N_3420);
nor U3970 (N_3970,N_3143,N_3068);
nor U3971 (N_3971,N_3328,N_3381);
nand U3972 (N_3972,N_3425,N_3453);
nand U3973 (N_3973,N_3154,N_3117);
and U3974 (N_3974,N_3497,N_3368);
nor U3975 (N_3975,N_3302,N_3392);
nand U3976 (N_3976,N_3026,N_3109);
and U3977 (N_3977,N_3016,N_3310);
and U3978 (N_3978,N_3152,N_3451);
or U3979 (N_3979,N_3132,N_3147);
or U3980 (N_3980,N_3113,N_3151);
or U3981 (N_3981,N_3464,N_3472);
nor U3982 (N_3982,N_3467,N_3043);
and U3983 (N_3983,N_3088,N_3229);
or U3984 (N_3984,N_3107,N_3374);
and U3985 (N_3985,N_3418,N_3358);
nand U3986 (N_3986,N_3215,N_3447);
and U3987 (N_3987,N_3256,N_3265);
or U3988 (N_3988,N_3205,N_3244);
or U3989 (N_3989,N_3429,N_3042);
nor U3990 (N_3990,N_3196,N_3320);
nand U3991 (N_3991,N_3180,N_3102);
nand U3992 (N_3992,N_3037,N_3203);
xor U3993 (N_3993,N_3340,N_3124);
nand U3994 (N_3994,N_3432,N_3155);
or U3995 (N_3995,N_3173,N_3034);
xnor U3996 (N_3996,N_3452,N_3462);
and U3997 (N_3997,N_3424,N_3455);
nand U3998 (N_3998,N_3214,N_3493);
nand U3999 (N_3999,N_3454,N_3014);
or U4000 (N_4000,N_3669,N_3698);
or U4001 (N_4001,N_3999,N_3855);
nand U4002 (N_4002,N_3977,N_3997);
nor U4003 (N_4003,N_3646,N_3601);
or U4004 (N_4004,N_3735,N_3627);
or U4005 (N_4005,N_3919,N_3776);
or U4006 (N_4006,N_3801,N_3725);
nor U4007 (N_4007,N_3633,N_3750);
nor U4008 (N_4008,N_3791,N_3928);
or U4009 (N_4009,N_3962,N_3586);
nand U4010 (N_4010,N_3677,N_3513);
nor U4011 (N_4011,N_3571,N_3993);
nor U4012 (N_4012,N_3834,N_3604);
nor U4013 (N_4013,N_3672,N_3754);
nand U4014 (N_4014,N_3810,N_3667);
or U4015 (N_4015,N_3583,N_3897);
nand U4016 (N_4016,N_3679,N_3610);
nor U4017 (N_4017,N_3642,N_3840);
and U4018 (N_4018,N_3971,N_3572);
and U4019 (N_4019,N_3934,N_3920);
and U4020 (N_4020,N_3518,N_3552);
xor U4021 (N_4021,N_3546,N_3884);
and U4022 (N_4022,N_3852,N_3980);
and U4023 (N_4023,N_3998,N_3770);
nor U4024 (N_4024,N_3841,N_3961);
nand U4025 (N_4025,N_3848,N_3868);
or U4026 (N_4026,N_3696,N_3932);
nand U4027 (N_4027,N_3638,N_3674);
nor U4028 (N_4028,N_3773,N_3579);
or U4029 (N_4029,N_3907,N_3875);
and U4030 (N_4030,N_3626,N_3511);
and U4031 (N_4031,N_3746,N_3715);
nand U4032 (N_4032,N_3592,N_3559);
nand U4033 (N_4033,N_3635,N_3764);
nor U4034 (N_4034,N_3719,N_3905);
or U4035 (N_4035,N_3712,N_3573);
or U4036 (N_4036,N_3726,N_3662);
and U4037 (N_4037,N_3976,N_3734);
nand U4038 (N_4038,N_3869,N_3979);
nor U4039 (N_4039,N_3590,N_3947);
and U4040 (N_4040,N_3664,N_3645);
nand U4041 (N_4041,N_3942,N_3866);
nand U4042 (N_4042,N_3703,N_3960);
nand U4043 (N_4043,N_3783,N_3524);
and U4044 (N_4044,N_3623,N_3737);
nand U4045 (N_4045,N_3930,N_3545);
nand U4046 (N_4046,N_3851,N_3804);
nand U4047 (N_4047,N_3671,N_3847);
or U4048 (N_4048,N_3506,N_3500);
nor U4049 (N_4049,N_3954,N_3582);
nand U4050 (N_4050,N_3793,N_3882);
and U4051 (N_4051,N_3892,N_3955);
nand U4052 (N_4052,N_3517,N_3742);
or U4053 (N_4053,N_3901,N_3588);
nor U4054 (N_4054,N_3758,N_3609);
or U4055 (N_4055,N_3876,N_3686);
nand U4056 (N_4056,N_3649,N_3702);
and U4057 (N_4057,N_3654,N_3641);
nand U4058 (N_4058,N_3913,N_3585);
nor U4059 (N_4059,N_3606,N_3807);
nor U4060 (N_4060,N_3822,N_3800);
or U4061 (N_4061,N_3661,N_3561);
nor U4062 (N_4062,N_3877,N_3631);
xor U4063 (N_4063,N_3666,N_3676);
and U4064 (N_4064,N_3630,N_3888);
nor U4065 (N_4065,N_3535,N_3973);
nand U4066 (N_4066,N_3587,N_3713);
nor U4067 (N_4067,N_3827,N_3727);
nand U4068 (N_4068,N_3914,N_3906);
or U4069 (N_4069,N_3943,N_3835);
or U4070 (N_4070,N_3844,N_3574);
nor U4071 (N_4071,N_3689,N_3933);
and U4072 (N_4072,N_3927,N_3755);
nand U4073 (N_4073,N_3789,N_3534);
nand U4074 (N_4074,N_3615,N_3828);
or U4075 (N_4075,N_3527,N_3519);
and U4076 (N_4076,N_3864,N_3597);
nor U4077 (N_4077,N_3724,N_3799);
and U4078 (N_4078,N_3687,N_3628);
nand U4079 (N_4079,N_3613,N_3826);
and U4080 (N_4080,N_3902,N_3707);
nor U4081 (N_4081,N_3910,N_3802);
nor U4082 (N_4082,N_3915,N_3714);
and U4083 (N_4083,N_3784,N_3854);
nand U4084 (N_4084,N_3565,N_3538);
nand U4085 (N_4085,N_3681,N_3651);
nand U4086 (N_4086,N_3818,N_3871);
and U4087 (N_4087,N_3832,N_3539);
and U4088 (N_4088,N_3772,N_3656);
nand U4089 (N_4089,N_3551,N_3767);
or U4090 (N_4090,N_3536,N_3952);
nor U4091 (N_4091,N_3863,N_3540);
and U4092 (N_4092,N_3987,N_3521);
nor U4093 (N_4093,N_3811,N_3577);
and U4094 (N_4094,N_3831,N_3945);
nor U4095 (N_4095,N_3872,N_3537);
nor U4096 (N_4096,N_3929,N_3984);
nand U4097 (N_4097,N_3838,N_3515);
nor U4098 (N_4098,N_3562,N_3706);
or U4099 (N_4099,N_3680,N_3723);
nor U4100 (N_4100,N_3529,N_3821);
or U4101 (N_4101,N_3760,N_3693);
or U4102 (N_4102,N_3603,N_3946);
nand U4103 (N_4103,N_3716,N_3570);
nand U4104 (N_4104,N_3958,N_3584);
nor U4105 (N_4105,N_3950,N_3568);
or U4106 (N_4106,N_3805,N_3599);
nand U4107 (N_4107,N_3820,N_3815);
or U4108 (N_4108,N_3777,N_3786);
or U4109 (N_4109,N_3912,N_3739);
nor U4110 (N_4110,N_3505,N_3873);
or U4111 (N_4111,N_3862,N_3925);
nor U4112 (N_4112,N_3660,N_3576);
nor U4113 (N_4113,N_3708,N_3652);
nor U4114 (N_4114,N_3553,N_3636);
nand U4115 (N_4115,N_3580,N_3629);
and U4116 (N_4116,N_3894,N_3775);
and U4117 (N_4117,N_3963,N_3618);
or U4118 (N_4118,N_3885,N_3602);
nand U4119 (N_4119,N_3850,N_3625);
nor U4120 (N_4120,N_3718,N_3640);
nand U4121 (N_4121,N_3996,N_3981);
nor U4122 (N_4122,N_3616,N_3830);
or U4123 (N_4123,N_3814,N_3556);
and U4124 (N_4124,N_3849,N_3607);
or U4125 (N_4125,N_3544,N_3532);
nand U4126 (N_4126,N_3798,N_3525);
nand U4127 (N_4127,N_3936,N_3989);
or U4128 (N_4128,N_3663,N_3992);
nand U4129 (N_4129,N_3756,N_3508);
nand U4130 (N_4130,N_3722,N_3874);
nor U4131 (N_4131,N_3622,N_3694);
nor U4132 (N_4132,N_3825,N_3939);
or U4133 (N_4133,N_3655,N_3731);
or U4134 (N_4134,N_3721,N_3757);
nand U4135 (N_4135,N_3909,N_3659);
or U4136 (N_4136,N_3878,N_3697);
and U4137 (N_4137,N_3780,N_3918);
nor U4138 (N_4138,N_3741,N_3951);
and U4139 (N_4139,N_3833,N_3774);
nand U4140 (N_4140,N_3900,N_3803);
and U4141 (N_4141,N_3937,N_3503);
nand U4142 (N_4142,N_3608,N_3891);
nand U4143 (N_4143,N_3895,N_3765);
or U4144 (N_4144,N_3717,N_3509);
and U4145 (N_4145,N_3904,N_3566);
nor U4146 (N_4146,N_3510,N_3879);
and U4147 (N_4147,N_3637,N_3729);
nand U4148 (N_4148,N_3978,N_3931);
nand U4149 (N_4149,N_3809,N_3682);
and U4150 (N_4150,N_3889,N_3795);
nand U4151 (N_4151,N_3787,N_3528);
and U4152 (N_4152,N_3598,N_3526);
nand U4153 (N_4153,N_3812,N_3563);
and U4154 (N_4154,N_3688,N_3881);
and U4155 (N_4155,N_3670,N_3883);
nor U4156 (N_4156,N_3639,N_3824);
nor U4157 (N_4157,N_3685,N_3970);
nand U4158 (N_4158,N_3614,N_3744);
or U4159 (N_4159,N_3968,N_3533);
and U4160 (N_4160,N_3782,N_3853);
nand U4161 (N_4161,N_3549,N_3763);
nor U4162 (N_4162,N_3569,N_3748);
nor U4163 (N_4163,N_3762,N_3771);
and U4164 (N_4164,N_3695,N_3857);
xor U4165 (N_4165,N_3589,N_3747);
and U4166 (N_4166,N_3781,N_3709);
nand U4167 (N_4167,N_3541,N_3745);
nand U4168 (N_4168,N_3966,N_3917);
or U4169 (N_4169,N_3531,N_3957);
nor U4170 (N_4170,N_3797,N_3880);
or U4171 (N_4171,N_3959,N_3557);
and U4172 (N_4172,N_3736,N_3938);
nand U4173 (N_4173,N_3520,N_3893);
nor U4174 (N_4174,N_3740,N_3859);
or U4175 (N_4175,N_3752,N_3792);
or U4176 (N_4176,N_3507,N_3898);
nand U4177 (N_4177,N_3543,N_3701);
nand U4178 (N_4178,N_3778,N_3547);
nand U4179 (N_4179,N_3710,N_3967);
nor U4180 (N_4180,N_3911,N_3972);
nor U4181 (N_4181,N_3720,N_3548);
nand U4182 (N_4182,N_3982,N_3819);
and U4183 (N_4183,N_3870,N_3665);
or U4184 (N_4184,N_3829,N_3949);
nand U4185 (N_4185,N_3964,N_3941);
or U4186 (N_4186,N_3594,N_3705);
nand U4187 (N_4187,N_3899,N_3948);
nor U4188 (N_4188,N_3617,N_3690);
nand U4189 (N_4189,N_3504,N_3704);
nor U4190 (N_4190,N_3643,N_3836);
nand U4191 (N_4191,N_3502,N_3823);
or U4192 (N_4192,N_3896,N_3845);
nand U4193 (N_4193,N_3650,N_3522);
or U4194 (N_4194,N_3953,N_3605);
and U4195 (N_4195,N_3751,N_3794);
and U4196 (N_4196,N_3985,N_3691);
nor U4197 (N_4197,N_3788,N_3839);
nor U4198 (N_4198,N_3624,N_3550);
or U4199 (N_4199,N_3619,N_3514);
xnor U4200 (N_4200,N_3890,N_3621);
nand U4201 (N_4201,N_3575,N_3634);
nand U4202 (N_4202,N_3501,N_3842);
nand U4203 (N_4203,N_3806,N_3983);
and U4204 (N_4204,N_3860,N_3908);
or U4205 (N_4205,N_3995,N_3887);
or U4206 (N_4206,N_3816,N_3657);
or U4207 (N_4207,N_3769,N_3865);
nand U4208 (N_4208,N_3935,N_3578);
or U4209 (N_4209,N_3916,N_3658);
nand U4210 (N_4210,N_3986,N_3523);
nand U4211 (N_4211,N_3940,N_3903);
nand U4212 (N_4212,N_3974,N_3856);
or U4213 (N_4213,N_3647,N_3738);
xnor U4214 (N_4214,N_3922,N_3567);
and U4215 (N_4215,N_3564,N_3595);
nand U4216 (N_4216,N_3969,N_3733);
nand U4217 (N_4217,N_3768,N_3994);
and U4218 (N_4218,N_3813,N_3796);
nand U4219 (N_4219,N_3684,N_3558);
nand U4220 (N_4220,N_3620,N_3790);
nand U4221 (N_4221,N_3542,N_3648);
and U4222 (N_4222,N_3730,N_3673);
nor U4223 (N_4223,N_3678,N_3944);
xor U4224 (N_4224,N_3581,N_3596);
and U4225 (N_4225,N_3728,N_3711);
xnor U4226 (N_4226,N_3843,N_3512);
nand U4227 (N_4227,N_3611,N_3591);
nand U4228 (N_4228,N_3921,N_3808);
nor U4229 (N_4229,N_3990,N_3886);
nor U4230 (N_4230,N_3761,N_3766);
and U4231 (N_4231,N_3516,N_3612);
nor U4232 (N_4232,N_3632,N_3600);
or U4233 (N_4233,N_3530,N_3785);
and U4234 (N_4234,N_3554,N_3749);
and U4235 (N_4235,N_3560,N_3683);
or U4236 (N_4236,N_3653,N_3975);
and U4237 (N_4237,N_3965,N_3759);
and U4238 (N_4238,N_3924,N_3926);
or U4239 (N_4239,N_3988,N_3668);
and U4240 (N_4240,N_3675,N_3991);
nand U4241 (N_4241,N_3692,N_3956);
nand U4242 (N_4242,N_3837,N_3699);
or U4243 (N_4243,N_3867,N_3700);
or U4244 (N_4244,N_3779,N_3858);
or U4245 (N_4245,N_3644,N_3593);
nor U4246 (N_4246,N_3817,N_3923);
nor U4247 (N_4247,N_3743,N_3846);
nor U4248 (N_4248,N_3555,N_3753);
nand U4249 (N_4249,N_3732,N_3861);
nor U4250 (N_4250,N_3612,N_3828);
nand U4251 (N_4251,N_3676,N_3793);
or U4252 (N_4252,N_3883,N_3845);
nand U4253 (N_4253,N_3764,N_3599);
nand U4254 (N_4254,N_3782,N_3876);
or U4255 (N_4255,N_3728,N_3760);
nor U4256 (N_4256,N_3551,N_3618);
nand U4257 (N_4257,N_3886,N_3519);
nand U4258 (N_4258,N_3866,N_3757);
nor U4259 (N_4259,N_3778,N_3936);
or U4260 (N_4260,N_3768,N_3948);
or U4261 (N_4261,N_3937,N_3643);
and U4262 (N_4262,N_3884,N_3544);
xnor U4263 (N_4263,N_3754,N_3646);
nand U4264 (N_4264,N_3882,N_3746);
or U4265 (N_4265,N_3726,N_3518);
xnor U4266 (N_4266,N_3740,N_3821);
or U4267 (N_4267,N_3907,N_3519);
nor U4268 (N_4268,N_3616,N_3526);
nand U4269 (N_4269,N_3790,N_3721);
nand U4270 (N_4270,N_3612,N_3576);
or U4271 (N_4271,N_3814,N_3563);
nand U4272 (N_4272,N_3914,N_3772);
and U4273 (N_4273,N_3849,N_3538);
and U4274 (N_4274,N_3740,N_3753);
nor U4275 (N_4275,N_3917,N_3703);
or U4276 (N_4276,N_3685,N_3818);
and U4277 (N_4277,N_3637,N_3894);
nand U4278 (N_4278,N_3935,N_3604);
nand U4279 (N_4279,N_3763,N_3582);
or U4280 (N_4280,N_3705,N_3778);
or U4281 (N_4281,N_3820,N_3760);
nor U4282 (N_4282,N_3523,N_3879);
nor U4283 (N_4283,N_3961,N_3567);
nor U4284 (N_4284,N_3754,N_3558);
or U4285 (N_4285,N_3686,N_3909);
or U4286 (N_4286,N_3660,N_3604);
nor U4287 (N_4287,N_3566,N_3686);
nand U4288 (N_4288,N_3933,N_3697);
nor U4289 (N_4289,N_3755,N_3916);
and U4290 (N_4290,N_3507,N_3504);
nor U4291 (N_4291,N_3775,N_3650);
and U4292 (N_4292,N_3761,N_3987);
and U4293 (N_4293,N_3543,N_3751);
nor U4294 (N_4294,N_3613,N_3592);
and U4295 (N_4295,N_3864,N_3625);
nor U4296 (N_4296,N_3521,N_3633);
nand U4297 (N_4297,N_3766,N_3767);
nor U4298 (N_4298,N_3980,N_3516);
nor U4299 (N_4299,N_3586,N_3887);
xor U4300 (N_4300,N_3742,N_3743);
nor U4301 (N_4301,N_3751,N_3674);
and U4302 (N_4302,N_3797,N_3856);
and U4303 (N_4303,N_3960,N_3601);
or U4304 (N_4304,N_3695,N_3788);
nand U4305 (N_4305,N_3836,N_3765);
nand U4306 (N_4306,N_3638,N_3879);
xor U4307 (N_4307,N_3611,N_3688);
or U4308 (N_4308,N_3873,N_3559);
nand U4309 (N_4309,N_3945,N_3707);
nor U4310 (N_4310,N_3809,N_3761);
nor U4311 (N_4311,N_3871,N_3886);
and U4312 (N_4312,N_3657,N_3526);
and U4313 (N_4313,N_3897,N_3841);
nor U4314 (N_4314,N_3727,N_3568);
nor U4315 (N_4315,N_3800,N_3847);
or U4316 (N_4316,N_3872,N_3735);
or U4317 (N_4317,N_3880,N_3926);
or U4318 (N_4318,N_3941,N_3589);
and U4319 (N_4319,N_3637,N_3772);
nand U4320 (N_4320,N_3922,N_3752);
nor U4321 (N_4321,N_3695,N_3766);
and U4322 (N_4322,N_3822,N_3620);
nor U4323 (N_4323,N_3636,N_3952);
or U4324 (N_4324,N_3610,N_3645);
nand U4325 (N_4325,N_3878,N_3680);
nor U4326 (N_4326,N_3958,N_3726);
and U4327 (N_4327,N_3802,N_3932);
nand U4328 (N_4328,N_3842,N_3662);
or U4329 (N_4329,N_3948,N_3777);
nand U4330 (N_4330,N_3836,N_3849);
nor U4331 (N_4331,N_3883,N_3753);
or U4332 (N_4332,N_3696,N_3575);
or U4333 (N_4333,N_3708,N_3856);
nand U4334 (N_4334,N_3887,N_3574);
nand U4335 (N_4335,N_3818,N_3551);
or U4336 (N_4336,N_3774,N_3691);
nand U4337 (N_4337,N_3572,N_3744);
nand U4338 (N_4338,N_3754,N_3699);
and U4339 (N_4339,N_3526,N_3535);
xor U4340 (N_4340,N_3734,N_3918);
nand U4341 (N_4341,N_3622,N_3804);
or U4342 (N_4342,N_3923,N_3511);
nor U4343 (N_4343,N_3979,N_3721);
xor U4344 (N_4344,N_3913,N_3637);
and U4345 (N_4345,N_3979,N_3578);
nand U4346 (N_4346,N_3718,N_3789);
and U4347 (N_4347,N_3619,N_3871);
nor U4348 (N_4348,N_3807,N_3563);
nor U4349 (N_4349,N_3920,N_3649);
and U4350 (N_4350,N_3872,N_3811);
nor U4351 (N_4351,N_3529,N_3968);
and U4352 (N_4352,N_3867,N_3533);
xnor U4353 (N_4353,N_3579,N_3787);
nand U4354 (N_4354,N_3843,N_3969);
nand U4355 (N_4355,N_3627,N_3898);
and U4356 (N_4356,N_3523,N_3546);
nand U4357 (N_4357,N_3693,N_3808);
and U4358 (N_4358,N_3816,N_3520);
nor U4359 (N_4359,N_3547,N_3620);
or U4360 (N_4360,N_3839,N_3994);
nor U4361 (N_4361,N_3580,N_3679);
and U4362 (N_4362,N_3594,N_3848);
and U4363 (N_4363,N_3761,N_3903);
and U4364 (N_4364,N_3637,N_3611);
nor U4365 (N_4365,N_3561,N_3502);
and U4366 (N_4366,N_3573,N_3793);
and U4367 (N_4367,N_3968,N_3659);
and U4368 (N_4368,N_3702,N_3644);
or U4369 (N_4369,N_3602,N_3904);
and U4370 (N_4370,N_3896,N_3851);
nand U4371 (N_4371,N_3736,N_3630);
nand U4372 (N_4372,N_3537,N_3991);
nand U4373 (N_4373,N_3576,N_3898);
or U4374 (N_4374,N_3819,N_3985);
nand U4375 (N_4375,N_3862,N_3761);
and U4376 (N_4376,N_3566,N_3939);
nand U4377 (N_4377,N_3722,N_3725);
or U4378 (N_4378,N_3558,N_3553);
or U4379 (N_4379,N_3677,N_3536);
nand U4380 (N_4380,N_3937,N_3628);
and U4381 (N_4381,N_3894,N_3654);
nor U4382 (N_4382,N_3515,N_3616);
nand U4383 (N_4383,N_3631,N_3938);
nand U4384 (N_4384,N_3521,N_3836);
or U4385 (N_4385,N_3592,N_3914);
nand U4386 (N_4386,N_3943,N_3996);
or U4387 (N_4387,N_3874,N_3964);
or U4388 (N_4388,N_3865,N_3570);
or U4389 (N_4389,N_3753,N_3767);
nand U4390 (N_4390,N_3826,N_3622);
nand U4391 (N_4391,N_3569,N_3839);
nand U4392 (N_4392,N_3560,N_3784);
nor U4393 (N_4393,N_3670,N_3998);
and U4394 (N_4394,N_3600,N_3511);
nand U4395 (N_4395,N_3869,N_3611);
or U4396 (N_4396,N_3872,N_3591);
or U4397 (N_4397,N_3925,N_3989);
nor U4398 (N_4398,N_3691,N_3863);
xnor U4399 (N_4399,N_3742,N_3956);
or U4400 (N_4400,N_3979,N_3906);
or U4401 (N_4401,N_3919,N_3609);
nor U4402 (N_4402,N_3970,N_3551);
or U4403 (N_4403,N_3783,N_3731);
or U4404 (N_4404,N_3855,N_3926);
and U4405 (N_4405,N_3549,N_3774);
or U4406 (N_4406,N_3769,N_3713);
nand U4407 (N_4407,N_3848,N_3904);
nor U4408 (N_4408,N_3839,N_3673);
nand U4409 (N_4409,N_3763,N_3817);
nor U4410 (N_4410,N_3544,N_3935);
and U4411 (N_4411,N_3528,N_3608);
nand U4412 (N_4412,N_3699,N_3565);
xor U4413 (N_4413,N_3853,N_3915);
nand U4414 (N_4414,N_3726,N_3538);
nand U4415 (N_4415,N_3658,N_3742);
nor U4416 (N_4416,N_3818,N_3849);
or U4417 (N_4417,N_3839,N_3880);
xnor U4418 (N_4418,N_3616,N_3794);
nor U4419 (N_4419,N_3895,N_3712);
xnor U4420 (N_4420,N_3917,N_3522);
and U4421 (N_4421,N_3744,N_3571);
or U4422 (N_4422,N_3645,N_3580);
and U4423 (N_4423,N_3817,N_3703);
or U4424 (N_4424,N_3724,N_3977);
nand U4425 (N_4425,N_3738,N_3723);
or U4426 (N_4426,N_3705,N_3907);
nor U4427 (N_4427,N_3558,N_3721);
and U4428 (N_4428,N_3585,N_3692);
and U4429 (N_4429,N_3785,N_3971);
nand U4430 (N_4430,N_3770,N_3710);
and U4431 (N_4431,N_3579,N_3532);
and U4432 (N_4432,N_3986,N_3550);
and U4433 (N_4433,N_3552,N_3842);
nor U4434 (N_4434,N_3946,N_3691);
and U4435 (N_4435,N_3938,N_3567);
and U4436 (N_4436,N_3717,N_3558);
nand U4437 (N_4437,N_3959,N_3660);
and U4438 (N_4438,N_3791,N_3878);
or U4439 (N_4439,N_3774,N_3631);
or U4440 (N_4440,N_3595,N_3713);
nor U4441 (N_4441,N_3887,N_3676);
and U4442 (N_4442,N_3718,N_3909);
nand U4443 (N_4443,N_3768,N_3893);
and U4444 (N_4444,N_3671,N_3739);
nor U4445 (N_4445,N_3847,N_3810);
nor U4446 (N_4446,N_3558,N_3848);
nor U4447 (N_4447,N_3574,N_3842);
or U4448 (N_4448,N_3559,N_3851);
and U4449 (N_4449,N_3993,N_3969);
and U4450 (N_4450,N_3719,N_3770);
and U4451 (N_4451,N_3763,N_3561);
or U4452 (N_4452,N_3628,N_3861);
or U4453 (N_4453,N_3534,N_3694);
or U4454 (N_4454,N_3991,N_3658);
nand U4455 (N_4455,N_3829,N_3935);
nor U4456 (N_4456,N_3881,N_3558);
or U4457 (N_4457,N_3801,N_3993);
or U4458 (N_4458,N_3969,N_3826);
or U4459 (N_4459,N_3839,N_3713);
or U4460 (N_4460,N_3512,N_3694);
or U4461 (N_4461,N_3954,N_3931);
nor U4462 (N_4462,N_3703,N_3948);
or U4463 (N_4463,N_3980,N_3620);
or U4464 (N_4464,N_3876,N_3705);
nand U4465 (N_4465,N_3938,N_3932);
nand U4466 (N_4466,N_3831,N_3901);
nor U4467 (N_4467,N_3834,N_3992);
or U4468 (N_4468,N_3648,N_3631);
nand U4469 (N_4469,N_3805,N_3840);
or U4470 (N_4470,N_3585,N_3730);
nor U4471 (N_4471,N_3961,N_3772);
or U4472 (N_4472,N_3612,N_3676);
nand U4473 (N_4473,N_3920,N_3892);
xnor U4474 (N_4474,N_3630,N_3862);
nor U4475 (N_4475,N_3822,N_3538);
nor U4476 (N_4476,N_3551,N_3760);
nand U4477 (N_4477,N_3636,N_3563);
nand U4478 (N_4478,N_3723,N_3881);
or U4479 (N_4479,N_3756,N_3739);
and U4480 (N_4480,N_3839,N_3935);
nor U4481 (N_4481,N_3685,N_3583);
nand U4482 (N_4482,N_3810,N_3789);
nand U4483 (N_4483,N_3504,N_3703);
nand U4484 (N_4484,N_3740,N_3876);
nand U4485 (N_4485,N_3928,N_3871);
or U4486 (N_4486,N_3767,N_3794);
nand U4487 (N_4487,N_3883,N_3652);
nand U4488 (N_4488,N_3610,N_3974);
and U4489 (N_4489,N_3750,N_3643);
xnor U4490 (N_4490,N_3984,N_3777);
nand U4491 (N_4491,N_3715,N_3635);
nand U4492 (N_4492,N_3673,N_3578);
nand U4493 (N_4493,N_3820,N_3974);
and U4494 (N_4494,N_3611,N_3622);
and U4495 (N_4495,N_3777,N_3847);
or U4496 (N_4496,N_3929,N_3731);
nand U4497 (N_4497,N_3929,N_3581);
nand U4498 (N_4498,N_3743,N_3709);
nand U4499 (N_4499,N_3812,N_3943);
or U4500 (N_4500,N_4268,N_4042);
nor U4501 (N_4501,N_4453,N_4437);
nor U4502 (N_4502,N_4390,N_4252);
nor U4503 (N_4503,N_4298,N_4196);
nand U4504 (N_4504,N_4466,N_4074);
nor U4505 (N_4505,N_4379,N_4398);
nor U4506 (N_4506,N_4475,N_4280);
nand U4507 (N_4507,N_4295,N_4053);
xor U4508 (N_4508,N_4380,N_4355);
nand U4509 (N_4509,N_4394,N_4415);
nor U4510 (N_4510,N_4184,N_4465);
or U4511 (N_4511,N_4309,N_4271);
or U4512 (N_4512,N_4425,N_4121);
and U4513 (N_4513,N_4476,N_4222);
nand U4514 (N_4514,N_4468,N_4301);
nand U4515 (N_4515,N_4435,N_4323);
nand U4516 (N_4516,N_4395,N_4027);
and U4517 (N_4517,N_4081,N_4099);
or U4518 (N_4518,N_4140,N_4009);
or U4519 (N_4519,N_4063,N_4236);
nor U4520 (N_4520,N_4373,N_4489);
and U4521 (N_4521,N_4024,N_4003);
or U4522 (N_4522,N_4467,N_4039);
or U4523 (N_4523,N_4242,N_4080);
nor U4524 (N_4524,N_4017,N_4103);
nand U4525 (N_4525,N_4441,N_4360);
nand U4526 (N_4526,N_4311,N_4033);
nand U4527 (N_4527,N_4424,N_4075);
and U4528 (N_4528,N_4334,N_4105);
nand U4529 (N_4529,N_4123,N_4018);
nor U4530 (N_4530,N_4345,N_4212);
and U4531 (N_4531,N_4240,N_4115);
and U4532 (N_4532,N_4219,N_4186);
or U4533 (N_4533,N_4317,N_4166);
or U4534 (N_4534,N_4091,N_4176);
nor U4535 (N_4535,N_4384,N_4217);
and U4536 (N_4536,N_4291,N_4329);
and U4537 (N_4537,N_4431,N_4088);
or U4538 (N_4538,N_4193,N_4104);
nand U4539 (N_4539,N_4070,N_4092);
or U4540 (N_4540,N_4327,N_4410);
or U4541 (N_4541,N_4264,N_4332);
or U4542 (N_4542,N_4257,N_4248);
and U4543 (N_4543,N_4019,N_4457);
nand U4544 (N_4544,N_4383,N_4482);
nand U4545 (N_4545,N_4443,N_4245);
and U4546 (N_4546,N_4270,N_4470);
nor U4547 (N_4547,N_4031,N_4396);
nand U4548 (N_4548,N_4071,N_4138);
nor U4549 (N_4549,N_4374,N_4141);
or U4550 (N_4550,N_4029,N_4224);
and U4551 (N_4551,N_4045,N_4249);
nand U4552 (N_4552,N_4417,N_4126);
nand U4553 (N_4553,N_4096,N_4203);
and U4554 (N_4554,N_4343,N_4206);
nand U4555 (N_4555,N_4218,N_4116);
and U4556 (N_4556,N_4066,N_4168);
nand U4557 (N_4557,N_4162,N_4259);
nand U4558 (N_4558,N_4172,N_4055);
nor U4559 (N_4559,N_4117,N_4354);
xnor U4560 (N_4560,N_4461,N_4335);
or U4561 (N_4561,N_4296,N_4174);
nand U4562 (N_4562,N_4064,N_4118);
and U4563 (N_4563,N_4388,N_4269);
and U4564 (N_4564,N_4223,N_4399);
nand U4565 (N_4565,N_4178,N_4146);
nand U4566 (N_4566,N_4190,N_4130);
nor U4567 (N_4567,N_4488,N_4287);
nand U4568 (N_4568,N_4049,N_4378);
and U4569 (N_4569,N_4273,N_4450);
nand U4570 (N_4570,N_4459,N_4095);
and U4571 (N_4571,N_4256,N_4237);
nand U4572 (N_4572,N_4397,N_4032);
nand U4573 (N_4573,N_4142,N_4175);
nor U4574 (N_4574,N_4386,N_4285);
xnor U4575 (N_4575,N_4226,N_4061);
nand U4576 (N_4576,N_4479,N_4065);
and U4577 (N_4577,N_4491,N_4098);
or U4578 (N_4578,N_4127,N_4026);
nand U4579 (N_4579,N_4004,N_4315);
nand U4580 (N_4580,N_4407,N_4434);
and U4581 (N_4581,N_4093,N_4179);
nor U4582 (N_4582,N_4128,N_4154);
nand U4583 (N_4583,N_4367,N_4180);
and U4584 (N_4584,N_4144,N_4238);
nand U4585 (N_4585,N_4101,N_4318);
nor U4586 (N_4586,N_4233,N_4173);
nand U4587 (N_4587,N_4089,N_4356);
or U4588 (N_4588,N_4052,N_4243);
nand U4589 (N_4589,N_4119,N_4361);
nor U4590 (N_4590,N_4136,N_4008);
or U4591 (N_4591,N_4021,N_4062);
nand U4592 (N_4592,N_4312,N_4023);
and U4593 (N_4593,N_4428,N_4325);
nor U4594 (N_4594,N_4451,N_4215);
and U4595 (N_4595,N_4349,N_4283);
nor U4596 (N_4596,N_4346,N_4412);
or U4597 (N_4597,N_4342,N_4068);
nand U4598 (N_4598,N_4494,N_4151);
or U4599 (N_4599,N_4200,N_4035);
nor U4600 (N_4600,N_4170,N_4389);
nor U4601 (N_4601,N_4492,N_4133);
nor U4602 (N_4602,N_4198,N_4387);
or U4603 (N_4603,N_4446,N_4082);
nor U4604 (N_4604,N_4007,N_4185);
and U4605 (N_4605,N_4051,N_4368);
nor U4606 (N_4606,N_4111,N_4421);
and U4607 (N_4607,N_4213,N_4205);
or U4608 (N_4608,N_4013,N_4228);
nor U4609 (N_4609,N_4038,N_4278);
or U4610 (N_4610,N_4258,N_4404);
nand U4611 (N_4611,N_4324,N_4385);
nand U4612 (N_4612,N_4015,N_4057);
nand U4613 (N_4613,N_4294,N_4197);
xor U4614 (N_4614,N_4282,N_4471);
nand U4615 (N_4615,N_4498,N_4487);
and U4616 (N_4616,N_4267,N_4316);
nand U4617 (N_4617,N_4485,N_4211);
and U4618 (N_4618,N_4192,N_4375);
and U4619 (N_4619,N_4303,N_4432);
nor U4620 (N_4620,N_4352,N_4181);
nor U4621 (N_4621,N_4382,N_4430);
and U4622 (N_4622,N_4107,N_4194);
or U4623 (N_4623,N_4293,N_4177);
or U4624 (N_4624,N_4137,N_4094);
and U4625 (N_4625,N_4261,N_4069);
nor U4626 (N_4626,N_4182,N_4260);
nor U4627 (N_4627,N_4159,N_4490);
nor U4628 (N_4628,N_4108,N_4158);
or U4629 (N_4629,N_4125,N_4429);
and U4630 (N_4630,N_4363,N_4114);
and U4631 (N_4631,N_4497,N_4416);
nand U4632 (N_4632,N_4310,N_4148);
nand U4633 (N_4633,N_4155,N_4207);
nand U4634 (N_4634,N_4244,N_4201);
nand U4635 (N_4635,N_4037,N_4247);
nand U4636 (N_4636,N_4326,N_4290);
or U4637 (N_4637,N_4251,N_4420);
and U4638 (N_4638,N_4321,N_4406);
and U4639 (N_4639,N_4411,N_4231);
and U4640 (N_4640,N_4357,N_4254);
or U4641 (N_4641,N_4030,N_4036);
nand U4642 (N_4642,N_4433,N_4348);
nor U4643 (N_4643,N_4391,N_4145);
xnor U4644 (N_4644,N_4085,N_4135);
nand U4645 (N_4645,N_4110,N_4072);
and U4646 (N_4646,N_4376,N_4333);
and U4647 (N_4647,N_4050,N_4350);
and U4648 (N_4648,N_4447,N_4149);
and U4649 (N_4649,N_4143,N_4302);
and U4650 (N_4650,N_4187,N_4167);
nand U4651 (N_4651,N_4478,N_4477);
nand U4652 (N_4652,N_4448,N_4454);
or U4653 (N_4653,N_4084,N_4010);
nor U4654 (N_4654,N_4402,N_4371);
or U4655 (N_4655,N_4444,N_4191);
or U4656 (N_4656,N_4022,N_4163);
nor U4657 (N_4657,N_4460,N_4043);
or U4658 (N_4658,N_4210,N_4235);
or U4659 (N_4659,N_4372,N_4147);
nand U4660 (N_4660,N_4202,N_4308);
nand U4661 (N_4661,N_4073,N_4359);
and U4662 (N_4662,N_4328,N_4006);
or U4663 (N_4663,N_4486,N_4161);
or U4664 (N_4664,N_4239,N_4083);
or U4665 (N_4665,N_4409,N_4358);
nand U4666 (N_4666,N_4274,N_4067);
and U4667 (N_4667,N_4165,N_4455);
nand U4668 (N_4668,N_4279,N_4129);
or U4669 (N_4669,N_4299,N_4436);
nand U4670 (N_4670,N_4208,N_4336);
nand U4671 (N_4671,N_4134,N_4253);
nor U4672 (N_4672,N_4120,N_4225);
or U4673 (N_4673,N_4124,N_4289);
and U4674 (N_4674,N_4044,N_4422);
nor U4675 (N_4675,N_4364,N_4054);
nor U4676 (N_4676,N_4047,N_4304);
nand U4677 (N_4677,N_4427,N_4353);
nor U4678 (N_4678,N_4189,N_4370);
nand U4679 (N_4679,N_4106,N_4087);
nand U4680 (N_4680,N_4195,N_4493);
and U4681 (N_4681,N_4014,N_4331);
or U4682 (N_4682,N_4495,N_4306);
and U4683 (N_4683,N_4473,N_4276);
nand U4684 (N_4684,N_4481,N_4419);
nand U4685 (N_4685,N_4499,N_4322);
and U4686 (N_4686,N_4011,N_4000);
or U4687 (N_4687,N_4438,N_4262);
nor U4688 (N_4688,N_4418,N_4059);
nand U4689 (N_4689,N_4340,N_4246);
nor U4690 (N_4690,N_4401,N_4028);
or U4691 (N_4691,N_4220,N_4169);
and U4692 (N_4692,N_4277,N_4077);
or U4693 (N_4693,N_4463,N_4100);
nand U4694 (N_4694,N_4265,N_4232);
or U4695 (N_4695,N_4034,N_4392);
or U4696 (N_4696,N_4483,N_4016);
and U4697 (N_4697,N_4171,N_4097);
nor U4698 (N_4698,N_4164,N_4408);
nand U4699 (N_4699,N_4230,N_4403);
and U4700 (N_4700,N_4377,N_4480);
or U4701 (N_4701,N_4040,N_4400);
nor U4702 (N_4702,N_4250,N_4351);
nor U4703 (N_4703,N_4458,N_4362);
nor U4704 (N_4704,N_4079,N_4426);
nand U4705 (N_4705,N_4439,N_4314);
and U4706 (N_4706,N_4381,N_4307);
or U4707 (N_4707,N_4440,N_4413);
nand U4708 (N_4708,N_4229,N_4109);
nor U4709 (N_4709,N_4060,N_4442);
or U4710 (N_4710,N_4339,N_4313);
or U4711 (N_4711,N_4474,N_4405);
nand U4712 (N_4712,N_4157,N_4112);
nand U4713 (N_4713,N_4496,N_4320);
nor U4714 (N_4714,N_4150,N_4338);
or U4715 (N_4715,N_4020,N_4469);
nor U4716 (N_4716,N_4058,N_4209);
and U4717 (N_4717,N_4366,N_4160);
nand U4718 (N_4718,N_4005,N_4263);
and U4719 (N_4719,N_4241,N_4369);
or U4720 (N_4720,N_4456,N_4472);
nor U4721 (N_4721,N_4292,N_4305);
and U4722 (N_4722,N_4462,N_4156);
or U4723 (N_4723,N_4341,N_4041);
nand U4724 (N_4724,N_4423,N_4076);
nand U4725 (N_4725,N_4086,N_4090);
and U4726 (N_4726,N_4266,N_4214);
nor U4727 (N_4727,N_4227,N_4025);
or U4728 (N_4728,N_4464,N_4132);
and U4729 (N_4729,N_4046,N_4216);
and U4730 (N_4730,N_4297,N_4199);
xor U4731 (N_4731,N_4393,N_4330);
nor U4732 (N_4732,N_4286,N_4139);
nand U4733 (N_4733,N_4188,N_4153);
or U4734 (N_4734,N_4344,N_4001);
and U4735 (N_4735,N_4056,N_4445);
or U4736 (N_4736,N_4221,N_4449);
nand U4737 (N_4737,N_4078,N_4204);
or U4738 (N_4738,N_4272,N_4288);
nor U4739 (N_4739,N_4152,N_4281);
and U4740 (N_4740,N_4284,N_4183);
nor U4741 (N_4741,N_4347,N_4012);
or U4742 (N_4742,N_4102,N_4300);
and U4743 (N_4743,N_4122,N_4365);
nand U4744 (N_4744,N_4113,N_4131);
nor U4745 (N_4745,N_4414,N_4337);
nand U4746 (N_4746,N_4452,N_4275);
xnor U4747 (N_4747,N_4002,N_4484);
nor U4748 (N_4748,N_4319,N_4234);
or U4749 (N_4749,N_4048,N_4255);
and U4750 (N_4750,N_4144,N_4355);
or U4751 (N_4751,N_4496,N_4466);
or U4752 (N_4752,N_4026,N_4325);
nand U4753 (N_4753,N_4337,N_4341);
and U4754 (N_4754,N_4290,N_4293);
and U4755 (N_4755,N_4334,N_4076);
nor U4756 (N_4756,N_4188,N_4135);
and U4757 (N_4757,N_4131,N_4365);
or U4758 (N_4758,N_4220,N_4353);
nor U4759 (N_4759,N_4061,N_4493);
and U4760 (N_4760,N_4215,N_4344);
or U4761 (N_4761,N_4101,N_4201);
and U4762 (N_4762,N_4312,N_4053);
nor U4763 (N_4763,N_4347,N_4458);
and U4764 (N_4764,N_4144,N_4416);
nor U4765 (N_4765,N_4457,N_4371);
nor U4766 (N_4766,N_4223,N_4427);
or U4767 (N_4767,N_4259,N_4136);
nor U4768 (N_4768,N_4025,N_4147);
or U4769 (N_4769,N_4058,N_4276);
or U4770 (N_4770,N_4177,N_4121);
nand U4771 (N_4771,N_4042,N_4355);
xor U4772 (N_4772,N_4352,N_4407);
nor U4773 (N_4773,N_4489,N_4152);
and U4774 (N_4774,N_4267,N_4248);
nand U4775 (N_4775,N_4174,N_4097);
nand U4776 (N_4776,N_4101,N_4001);
nand U4777 (N_4777,N_4097,N_4090);
nor U4778 (N_4778,N_4119,N_4086);
nand U4779 (N_4779,N_4339,N_4391);
or U4780 (N_4780,N_4255,N_4154);
and U4781 (N_4781,N_4046,N_4016);
nand U4782 (N_4782,N_4207,N_4012);
nand U4783 (N_4783,N_4494,N_4032);
and U4784 (N_4784,N_4053,N_4417);
nand U4785 (N_4785,N_4047,N_4040);
nor U4786 (N_4786,N_4156,N_4185);
nand U4787 (N_4787,N_4139,N_4221);
xnor U4788 (N_4788,N_4486,N_4156);
nand U4789 (N_4789,N_4018,N_4450);
xor U4790 (N_4790,N_4192,N_4018);
and U4791 (N_4791,N_4360,N_4472);
xnor U4792 (N_4792,N_4248,N_4402);
nor U4793 (N_4793,N_4489,N_4092);
or U4794 (N_4794,N_4191,N_4430);
nand U4795 (N_4795,N_4128,N_4095);
and U4796 (N_4796,N_4209,N_4358);
or U4797 (N_4797,N_4468,N_4111);
xnor U4798 (N_4798,N_4236,N_4180);
and U4799 (N_4799,N_4176,N_4476);
or U4800 (N_4800,N_4326,N_4452);
and U4801 (N_4801,N_4118,N_4054);
nor U4802 (N_4802,N_4403,N_4212);
or U4803 (N_4803,N_4329,N_4454);
nand U4804 (N_4804,N_4158,N_4331);
or U4805 (N_4805,N_4069,N_4141);
nand U4806 (N_4806,N_4046,N_4262);
and U4807 (N_4807,N_4098,N_4112);
nor U4808 (N_4808,N_4185,N_4166);
nand U4809 (N_4809,N_4038,N_4216);
and U4810 (N_4810,N_4012,N_4452);
or U4811 (N_4811,N_4323,N_4072);
nand U4812 (N_4812,N_4306,N_4206);
and U4813 (N_4813,N_4248,N_4349);
nor U4814 (N_4814,N_4046,N_4105);
nor U4815 (N_4815,N_4412,N_4260);
nand U4816 (N_4816,N_4245,N_4129);
nand U4817 (N_4817,N_4267,N_4214);
nor U4818 (N_4818,N_4279,N_4201);
nand U4819 (N_4819,N_4282,N_4387);
nor U4820 (N_4820,N_4203,N_4198);
nand U4821 (N_4821,N_4348,N_4246);
or U4822 (N_4822,N_4411,N_4429);
or U4823 (N_4823,N_4197,N_4018);
nand U4824 (N_4824,N_4025,N_4368);
nor U4825 (N_4825,N_4213,N_4234);
and U4826 (N_4826,N_4069,N_4125);
or U4827 (N_4827,N_4455,N_4288);
nand U4828 (N_4828,N_4252,N_4413);
nand U4829 (N_4829,N_4272,N_4258);
and U4830 (N_4830,N_4320,N_4272);
nand U4831 (N_4831,N_4036,N_4241);
or U4832 (N_4832,N_4017,N_4007);
nor U4833 (N_4833,N_4379,N_4200);
nor U4834 (N_4834,N_4492,N_4392);
or U4835 (N_4835,N_4445,N_4267);
or U4836 (N_4836,N_4185,N_4378);
nor U4837 (N_4837,N_4309,N_4376);
nor U4838 (N_4838,N_4354,N_4127);
nand U4839 (N_4839,N_4353,N_4304);
or U4840 (N_4840,N_4488,N_4448);
or U4841 (N_4841,N_4420,N_4319);
xor U4842 (N_4842,N_4028,N_4352);
and U4843 (N_4843,N_4274,N_4123);
nand U4844 (N_4844,N_4223,N_4221);
and U4845 (N_4845,N_4078,N_4360);
nor U4846 (N_4846,N_4268,N_4338);
or U4847 (N_4847,N_4184,N_4201);
nand U4848 (N_4848,N_4329,N_4204);
nand U4849 (N_4849,N_4336,N_4403);
nand U4850 (N_4850,N_4095,N_4169);
xnor U4851 (N_4851,N_4115,N_4022);
and U4852 (N_4852,N_4421,N_4159);
and U4853 (N_4853,N_4095,N_4312);
xnor U4854 (N_4854,N_4304,N_4118);
or U4855 (N_4855,N_4166,N_4394);
or U4856 (N_4856,N_4469,N_4485);
nand U4857 (N_4857,N_4307,N_4186);
nand U4858 (N_4858,N_4011,N_4086);
nand U4859 (N_4859,N_4051,N_4420);
and U4860 (N_4860,N_4492,N_4126);
or U4861 (N_4861,N_4348,N_4316);
or U4862 (N_4862,N_4255,N_4301);
or U4863 (N_4863,N_4347,N_4497);
or U4864 (N_4864,N_4067,N_4053);
nor U4865 (N_4865,N_4392,N_4221);
and U4866 (N_4866,N_4262,N_4268);
nand U4867 (N_4867,N_4126,N_4250);
nor U4868 (N_4868,N_4209,N_4333);
and U4869 (N_4869,N_4045,N_4447);
and U4870 (N_4870,N_4433,N_4009);
and U4871 (N_4871,N_4073,N_4206);
or U4872 (N_4872,N_4326,N_4460);
and U4873 (N_4873,N_4117,N_4414);
or U4874 (N_4874,N_4020,N_4054);
xnor U4875 (N_4875,N_4351,N_4046);
and U4876 (N_4876,N_4264,N_4402);
or U4877 (N_4877,N_4287,N_4414);
nand U4878 (N_4878,N_4413,N_4114);
nor U4879 (N_4879,N_4375,N_4186);
nand U4880 (N_4880,N_4258,N_4289);
nand U4881 (N_4881,N_4135,N_4286);
nand U4882 (N_4882,N_4254,N_4076);
nor U4883 (N_4883,N_4030,N_4119);
nor U4884 (N_4884,N_4373,N_4435);
nor U4885 (N_4885,N_4257,N_4474);
nand U4886 (N_4886,N_4252,N_4376);
nor U4887 (N_4887,N_4218,N_4453);
nor U4888 (N_4888,N_4126,N_4437);
xnor U4889 (N_4889,N_4072,N_4388);
or U4890 (N_4890,N_4372,N_4310);
nand U4891 (N_4891,N_4417,N_4036);
and U4892 (N_4892,N_4446,N_4016);
and U4893 (N_4893,N_4109,N_4440);
nand U4894 (N_4894,N_4226,N_4272);
or U4895 (N_4895,N_4255,N_4020);
nand U4896 (N_4896,N_4241,N_4495);
nand U4897 (N_4897,N_4077,N_4386);
nand U4898 (N_4898,N_4261,N_4297);
nand U4899 (N_4899,N_4245,N_4304);
nand U4900 (N_4900,N_4293,N_4204);
nor U4901 (N_4901,N_4003,N_4082);
and U4902 (N_4902,N_4128,N_4351);
nand U4903 (N_4903,N_4013,N_4432);
nor U4904 (N_4904,N_4456,N_4032);
nor U4905 (N_4905,N_4241,N_4005);
xnor U4906 (N_4906,N_4333,N_4277);
nand U4907 (N_4907,N_4232,N_4249);
nand U4908 (N_4908,N_4323,N_4070);
and U4909 (N_4909,N_4310,N_4045);
or U4910 (N_4910,N_4361,N_4132);
or U4911 (N_4911,N_4238,N_4088);
nand U4912 (N_4912,N_4427,N_4000);
nor U4913 (N_4913,N_4244,N_4242);
nor U4914 (N_4914,N_4139,N_4463);
nand U4915 (N_4915,N_4286,N_4053);
xnor U4916 (N_4916,N_4149,N_4044);
nor U4917 (N_4917,N_4333,N_4346);
or U4918 (N_4918,N_4379,N_4444);
and U4919 (N_4919,N_4376,N_4115);
or U4920 (N_4920,N_4221,N_4074);
nor U4921 (N_4921,N_4273,N_4267);
nor U4922 (N_4922,N_4340,N_4373);
nor U4923 (N_4923,N_4068,N_4425);
or U4924 (N_4924,N_4496,N_4058);
and U4925 (N_4925,N_4480,N_4137);
xor U4926 (N_4926,N_4173,N_4346);
nand U4927 (N_4927,N_4414,N_4111);
or U4928 (N_4928,N_4054,N_4179);
nand U4929 (N_4929,N_4331,N_4313);
nand U4930 (N_4930,N_4085,N_4459);
nor U4931 (N_4931,N_4125,N_4247);
nand U4932 (N_4932,N_4334,N_4019);
nand U4933 (N_4933,N_4393,N_4486);
and U4934 (N_4934,N_4167,N_4242);
nand U4935 (N_4935,N_4229,N_4492);
nor U4936 (N_4936,N_4405,N_4361);
or U4937 (N_4937,N_4315,N_4216);
or U4938 (N_4938,N_4171,N_4467);
or U4939 (N_4939,N_4461,N_4322);
and U4940 (N_4940,N_4089,N_4458);
nor U4941 (N_4941,N_4282,N_4081);
nand U4942 (N_4942,N_4468,N_4164);
nand U4943 (N_4943,N_4240,N_4279);
nor U4944 (N_4944,N_4455,N_4294);
nand U4945 (N_4945,N_4064,N_4121);
and U4946 (N_4946,N_4452,N_4046);
xnor U4947 (N_4947,N_4064,N_4025);
or U4948 (N_4948,N_4256,N_4172);
nand U4949 (N_4949,N_4405,N_4045);
xnor U4950 (N_4950,N_4081,N_4139);
or U4951 (N_4951,N_4487,N_4348);
nor U4952 (N_4952,N_4445,N_4455);
nor U4953 (N_4953,N_4472,N_4220);
nor U4954 (N_4954,N_4235,N_4331);
or U4955 (N_4955,N_4309,N_4148);
and U4956 (N_4956,N_4455,N_4157);
nand U4957 (N_4957,N_4158,N_4168);
and U4958 (N_4958,N_4443,N_4268);
nand U4959 (N_4959,N_4016,N_4173);
or U4960 (N_4960,N_4254,N_4082);
nand U4961 (N_4961,N_4299,N_4410);
or U4962 (N_4962,N_4368,N_4224);
and U4963 (N_4963,N_4321,N_4315);
and U4964 (N_4964,N_4291,N_4111);
nor U4965 (N_4965,N_4192,N_4428);
nor U4966 (N_4966,N_4361,N_4400);
nor U4967 (N_4967,N_4262,N_4083);
and U4968 (N_4968,N_4333,N_4210);
and U4969 (N_4969,N_4304,N_4475);
and U4970 (N_4970,N_4112,N_4392);
nand U4971 (N_4971,N_4279,N_4471);
and U4972 (N_4972,N_4124,N_4065);
nor U4973 (N_4973,N_4325,N_4117);
nand U4974 (N_4974,N_4334,N_4435);
and U4975 (N_4975,N_4194,N_4205);
or U4976 (N_4976,N_4208,N_4098);
and U4977 (N_4977,N_4421,N_4003);
nor U4978 (N_4978,N_4481,N_4138);
nand U4979 (N_4979,N_4047,N_4338);
nand U4980 (N_4980,N_4166,N_4251);
and U4981 (N_4981,N_4294,N_4056);
or U4982 (N_4982,N_4014,N_4287);
nand U4983 (N_4983,N_4035,N_4433);
nor U4984 (N_4984,N_4108,N_4295);
nand U4985 (N_4985,N_4018,N_4496);
or U4986 (N_4986,N_4318,N_4089);
nor U4987 (N_4987,N_4186,N_4260);
nand U4988 (N_4988,N_4459,N_4190);
nor U4989 (N_4989,N_4445,N_4486);
or U4990 (N_4990,N_4306,N_4310);
and U4991 (N_4991,N_4446,N_4277);
or U4992 (N_4992,N_4263,N_4420);
and U4993 (N_4993,N_4074,N_4215);
or U4994 (N_4994,N_4145,N_4442);
nand U4995 (N_4995,N_4267,N_4231);
and U4996 (N_4996,N_4495,N_4104);
nand U4997 (N_4997,N_4081,N_4120);
nor U4998 (N_4998,N_4390,N_4263);
xnor U4999 (N_4999,N_4166,N_4064);
nor UO_0 (O_0,N_4720,N_4930);
xnor UO_1 (O_1,N_4602,N_4641);
nand UO_2 (O_2,N_4960,N_4903);
or UO_3 (O_3,N_4500,N_4701);
nor UO_4 (O_4,N_4689,N_4978);
nor UO_5 (O_5,N_4841,N_4652);
nand UO_6 (O_6,N_4775,N_4900);
nand UO_7 (O_7,N_4654,N_4699);
nand UO_8 (O_8,N_4547,N_4536);
or UO_9 (O_9,N_4564,N_4620);
nand UO_10 (O_10,N_4845,N_4924);
nand UO_11 (O_11,N_4661,N_4669);
or UO_12 (O_12,N_4736,N_4678);
nor UO_13 (O_13,N_4799,N_4835);
nand UO_14 (O_14,N_4862,N_4713);
or UO_15 (O_15,N_4864,N_4861);
nor UO_16 (O_16,N_4842,N_4828);
or UO_17 (O_17,N_4839,N_4541);
and UO_18 (O_18,N_4853,N_4762);
nor UO_19 (O_19,N_4994,N_4626);
and UO_20 (O_20,N_4525,N_4923);
or UO_21 (O_21,N_4926,N_4642);
nand UO_22 (O_22,N_4907,N_4848);
nor UO_23 (O_23,N_4532,N_4975);
and UO_24 (O_24,N_4553,N_4570);
nand UO_25 (O_25,N_4790,N_4821);
nor UO_26 (O_26,N_4581,N_4798);
and UO_27 (O_27,N_4727,N_4992);
or UO_28 (O_28,N_4885,N_4528);
nand UO_29 (O_29,N_4721,N_4941);
nor UO_30 (O_30,N_4719,N_4988);
and UO_31 (O_31,N_4991,N_4748);
or UO_32 (O_32,N_4769,N_4554);
nand UO_33 (O_33,N_4890,N_4706);
or UO_34 (O_34,N_4916,N_4674);
and UO_35 (O_35,N_4901,N_4793);
nand UO_36 (O_36,N_4921,N_4869);
and UO_37 (O_37,N_4632,N_4952);
nor UO_38 (O_38,N_4953,N_4568);
nor UO_39 (O_39,N_4716,N_4755);
or UO_40 (O_40,N_4605,N_4857);
nand UO_41 (O_41,N_4973,N_4780);
and UO_42 (O_42,N_4740,N_4644);
and UO_43 (O_43,N_4956,N_4730);
nand UO_44 (O_44,N_4792,N_4750);
nand UO_45 (O_45,N_4659,N_4741);
nor UO_46 (O_46,N_4932,N_4823);
nand UO_47 (O_47,N_4601,N_4722);
and UO_48 (O_48,N_4985,N_4922);
nand UO_49 (O_49,N_4779,N_4647);
nor UO_50 (O_50,N_4807,N_4888);
or UO_51 (O_51,N_4756,N_4809);
and UO_52 (O_52,N_4757,N_4688);
or UO_53 (O_53,N_4550,N_4855);
nand UO_54 (O_54,N_4598,N_4827);
or UO_55 (O_55,N_4627,N_4667);
and UO_56 (O_56,N_4612,N_4505);
nand UO_57 (O_57,N_4503,N_4993);
nand UO_58 (O_58,N_4970,N_4502);
nor UO_59 (O_59,N_4840,N_4518);
and UO_60 (O_60,N_4585,N_4977);
or UO_61 (O_61,N_4774,N_4843);
nor UO_62 (O_62,N_4596,N_4889);
nand UO_63 (O_63,N_4566,N_4844);
or UO_64 (O_64,N_4815,N_4574);
or UO_65 (O_65,N_4946,N_4898);
nor UO_66 (O_66,N_4990,N_4535);
nor UO_67 (O_67,N_4651,N_4653);
nand UO_68 (O_68,N_4909,N_4682);
or UO_69 (O_69,N_4506,N_4634);
or UO_70 (O_70,N_4707,N_4710);
and UO_71 (O_71,N_4943,N_4819);
nor UO_72 (O_72,N_4781,N_4666);
nand UO_73 (O_73,N_4982,N_4751);
or UO_74 (O_74,N_4562,N_4934);
and UO_75 (O_75,N_4747,N_4812);
xnor UO_76 (O_76,N_4618,N_4715);
nor UO_77 (O_77,N_4868,N_4530);
nand UO_78 (O_78,N_4734,N_4754);
and UO_79 (O_79,N_4725,N_4964);
nand UO_80 (O_80,N_4529,N_4696);
and UO_81 (O_81,N_4548,N_4965);
and UO_82 (O_82,N_4969,N_4694);
nand UO_83 (O_83,N_4692,N_4732);
xnor UO_84 (O_84,N_4789,N_4829);
or UO_85 (O_85,N_4933,N_4928);
nand UO_86 (O_86,N_4507,N_4940);
or UO_87 (O_87,N_4739,N_4860);
nand UO_88 (O_88,N_4545,N_4884);
or UO_89 (O_89,N_4847,N_4588);
and UO_90 (O_90,N_4501,N_4577);
or UO_91 (O_91,N_4981,N_4705);
nor UO_92 (O_92,N_4737,N_4818);
and UO_93 (O_93,N_4939,N_4886);
and UO_94 (O_94,N_4670,N_4595);
and UO_95 (O_95,N_4766,N_4521);
nand UO_96 (O_96,N_4572,N_4519);
nand UO_97 (O_97,N_4899,N_4947);
nand UO_98 (O_98,N_4656,N_4663);
and UO_99 (O_99,N_4534,N_4945);
or UO_100 (O_100,N_4557,N_4931);
and UO_101 (O_101,N_4524,N_4555);
and UO_102 (O_102,N_4785,N_4565);
and UO_103 (O_103,N_4830,N_4571);
and UO_104 (O_104,N_4797,N_4679);
or UO_105 (O_105,N_4735,N_4558);
nand UO_106 (O_106,N_4784,N_4971);
nor UO_107 (O_107,N_4879,N_4814);
nor UO_108 (O_108,N_4896,N_4984);
nor UO_109 (O_109,N_4673,N_4643);
nor UO_110 (O_110,N_4599,N_4915);
and UO_111 (O_111,N_4838,N_4594);
or UO_112 (O_112,N_4623,N_4802);
nand UO_113 (O_113,N_4708,N_4700);
or UO_114 (O_114,N_4579,N_4996);
or UO_115 (O_115,N_4801,N_4833);
nand UO_116 (O_116,N_4582,N_4718);
or UO_117 (O_117,N_4622,N_4972);
or UO_118 (O_118,N_4777,N_4877);
and UO_119 (O_119,N_4874,N_4948);
and UO_120 (O_120,N_4597,N_4794);
or UO_121 (O_121,N_4959,N_4825);
nand UO_122 (O_122,N_4675,N_4600);
nor UO_123 (O_123,N_4616,N_4995);
and UO_124 (O_124,N_4693,N_4662);
or UO_125 (O_125,N_4968,N_4808);
nor UO_126 (O_126,N_4504,N_4824);
or UO_127 (O_127,N_4559,N_4871);
nor UO_128 (O_128,N_4569,N_4983);
nor UO_129 (O_129,N_4687,N_4587);
nor UO_130 (O_130,N_4726,N_4752);
or UO_131 (O_131,N_4937,N_4786);
nor UO_132 (O_132,N_4731,N_4583);
or UO_133 (O_133,N_4925,N_4635);
nand UO_134 (O_134,N_4542,N_4552);
or UO_135 (O_135,N_4619,N_4677);
nor UO_136 (O_136,N_4614,N_4810);
nor UO_137 (O_137,N_4997,N_4998);
nand UO_138 (O_138,N_4893,N_4650);
or UO_139 (O_139,N_4544,N_4850);
xnor UO_140 (O_140,N_4849,N_4509);
xor UO_141 (O_141,N_4986,N_4686);
or UO_142 (O_142,N_4966,N_4580);
and UO_143 (O_143,N_4791,N_4753);
nor UO_144 (O_144,N_4962,N_4944);
nand UO_145 (O_145,N_4646,N_4717);
or UO_146 (O_146,N_4854,N_4846);
nor UO_147 (O_147,N_4743,N_4697);
nand UO_148 (O_148,N_4892,N_4665);
and UO_149 (O_149,N_4887,N_4578);
and UO_150 (O_150,N_4902,N_4856);
nor UO_151 (O_151,N_4549,N_4576);
nor UO_152 (O_152,N_4613,N_4684);
or UO_153 (O_153,N_4540,N_4629);
nand UO_154 (O_154,N_4607,N_4728);
and UO_155 (O_155,N_4526,N_4672);
and UO_156 (O_156,N_4639,N_4560);
nor UO_157 (O_157,N_4733,N_4767);
nand UO_158 (O_158,N_4522,N_4782);
nor UO_159 (O_159,N_4974,N_4563);
nand UO_160 (O_160,N_4624,N_4891);
nor UO_161 (O_161,N_4515,N_4875);
nor UO_162 (O_162,N_4745,N_4538);
and UO_163 (O_163,N_4852,N_4655);
and UO_164 (O_164,N_4537,N_4770);
and UO_165 (O_165,N_4744,N_4912);
and UO_166 (O_166,N_4698,N_4905);
nor UO_167 (O_167,N_4604,N_4691);
nor UO_168 (O_168,N_4917,N_4832);
nor UO_169 (O_169,N_4778,N_4546);
nor UO_170 (O_170,N_4609,N_4584);
or UO_171 (O_171,N_4951,N_4816);
nand UO_172 (O_172,N_4593,N_4904);
and UO_173 (O_173,N_4768,N_4954);
or UO_174 (O_174,N_4863,N_4615);
nor UO_175 (O_175,N_4938,N_4795);
and UO_176 (O_176,N_4764,N_4817);
or UO_177 (O_177,N_4551,N_4514);
or UO_178 (O_178,N_4870,N_4831);
or UO_179 (O_179,N_4950,N_4936);
nor UO_180 (O_180,N_4834,N_4883);
nand UO_181 (O_181,N_4906,N_4668);
or UO_182 (O_182,N_4603,N_4820);
nor UO_183 (O_183,N_4591,N_4702);
or UO_184 (O_184,N_4695,N_4703);
nand UO_185 (O_185,N_4586,N_4649);
or UO_186 (O_186,N_4573,N_4836);
nand UO_187 (O_187,N_4657,N_4908);
nand UO_188 (O_188,N_4685,N_4633);
nand UO_189 (O_189,N_4872,N_4920);
and UO_190 (O_190,N_4617,N_4935);
nand UO_191 (O_191,N_4837,N_4895);
nor UO_192 (O_192,N_4523,N_4771);
nand UO_193 (O_193,N_4592,N_4880);
or UO_194 (O_194,N_4631,N_4664);
nor UO_195 (O_195,N_4918,N_4967);
nor UO_196 (O_196,N_4712,N_4760);
or UO_197 (O_197,N_4957,N_4796);
and UO_198 (O_198,N_4758,N_4826);
nand UO_199 (O_199,N_4910,N_4671);
or UO_200 (O_200,N_4876,N_4513);
and UO_201 (O_201,N_4681,N_4683);
or UO_202 (O_202,N_4645,N_4999);
nor UO_203 (O_203,N_4919,N_4867);
nand UO_204 (O_204,N_4531,N_4927);
and UO_205 (O_205,N_4527,N_4800);
nand UO_206 (O_206,N_4512,N_4787);
nand UO_207 (O_207,N_4813,N_4711);
nand UO_208 (O_208,N_4961,N_4776);
nand UO_209 (O_209,N_4773,N_4676);
and UO_210 (O_210,N_4567,N_4783);
and UO_211 (O_211,N_4508,N_4628);
or UO_212 (O_212,N_4963,N_4987);
or UO_213 (O_213,N_4881,N_4606);
or UO_214 (O_214,N_4746,N_4714);
or UO_215 (O_215,N_4851,N_4866);
and UO_216 (O_216,N_4772,N_4822);
or UO_217 (O_217,N_4690,N_4805);
nand UO_218 (O_218,N_4803,N_4859);
nor UO_219 (O_219,N_4761,N_4949);
and UO_220 (O_220,N_4759,N_4873);
nand UO_221 (O_221,N_4704,N_4858);
nor UO_222 (O_222,N_4894,N_4729);
and UO_223 (O_223,N_4621,N_4897);
nand UO_224 (O_224,N_4680,N_4630);
nor UO_225 (O_225,N_4811,N_4958);
or UO_226 (O_226,N_4723,N_4638);
and UO_227 (O_227,N_4511,N_4543);
nor UO_228 (O_228,N_4648,N_4911);
or UO_229 (O_229,N_4516,N_4640);
or UO_230 (O_230,N_4742,N_4878);
nor UO_231 (O_231,N_4636,N_4590);
nand UO_232 (O_232,N_4589,N_4980);
nor UO_233 (O_233,N_4979,N_4608);
and UO_234 (O_234,N_4637,N_4520);
nor UO_235 (O_235,N_4914,N_4882);
nand UO_236 (O_236,N_4533,N_4942);
or UO_237 (O_237,N_4804,N_4976);
nand UO_238 (O_238,N_4611,N_4749);
nor UO_239 (O_239,N_4955,N_4625);
or UO_240 (O_240,N_4913,N_4806);
or UO_241 (O_241,N_4724,N_4575);
or UO_242 (O_242,N_4738,N_4763);
nor UO_243 (O_243,N_4788,N_4929);
and UO_244 (O_244,N_4765,N_4561);
and UO_245 (O_245,N_4539,N_4660);
nor UO_246 (O_246,N_4556,N_4510);
and UO_247 (O_247,N_4709,N_4658);
and UO_248 (O_248,N_4517,N_4865);
or UO_249 (O_249,N_4610,N_4989);
and UO_250 (O_250,N_4886,N_4770);
or UO_251 (O_251,N_4723,N_4747);
and UO_252 (O_252,N_4592,N_4941);
nor UO_253 (O_253,N_4640,N_4730);
and UO_254 (O_254,N_4642,N_4938);
xor UO_255 (O_255,N_4969,N_4524);
nand UO_256 (O_256,N_4596,N_4755);
nand UO_257 (O_257,N_4738,N_4942);
or UO_258 (O_258,N_4770,N_4782);
nor UO_259 (O_259,N_4887,N_4556);
nor UO_260 (O_260,N_4709,N_4916);
and UO_261 (O_261,N_4595,N_4510);
nand UO_262 (O_262,N_4658,N_4852);
nand UO_263 (O_263,N_4787,N_4726);
and UO_264 (O_264,N_4546,N_4755);
nor UO_265 (O_265,N_4937,N_4981);
and UO_266 (O_266,N_4754,N_4523);
or UO_267 (O_267,N_4656,N_4713);
and UO_268 (O_268,N_4535,N_4552);
nand UO_269 (O_269,N_4855,N_4718);
or UO_270 (O_270,N_4793,N_4652);
xnor UO_271 (O_271,N_4719,N_4853);
or UO_272 (O_272,N_4616,N_4877);
nor UO_273 (O_273,N_4553,N_4823);
nor UO_274 (O_274,N_4563,N_4522);
xnor UO_275 (O_275,N_4545,N_4666);
or UO_276 (O_276,N_4613,N_4648);
xnor UO_277 (O_277,N_4778,N_4911);
and UO_278 (O_278,N_4717,N_4732);
nand UO_279 (O_279,N_4686,N_4618);
xor UO_280 (O_280,N_4901,N_4683);
and UO_281 (O_281,N_4937,N_4611);
nand UO_282 (O_282,N_4544,N_4507);
nand UO_283 (O_283,N_4565,N_4672);
nor UO_284 (O_284,N_4713,N_4673);
and UO_285 (O_285,N_4719,N_4810);
nand UO_286 (O_286,N_4757,N_4656);
xnor UO_287 (O_287,N_4927,N_4674);
nor UO_288 (O_288,N_4538,N_4874);
nor UO_289 (O_289,N_4689,N_4619);
nor UO_290 (O_290,N_4983,N_4746);
or UO_291 (O_291,N_4855,N_4653);
nand UO_292 (O_292,N_4749,N_4593);
or UO_293 (O_293,N_4716,N_4670);
nand UO_294 (O_294,N_4743,N_4588);
nand UO_295 (O_295,N_4524,N_4716);
nor UO_296 (O_296,N_4910,N_4807);
or UO_297 (O_297,N_4932,N_4586);
or UO_298 (O_298,N_4684,N_4888);
xor UO_299 (O_299,N_4859,N_4770);
nand UO_300 (O_300,N_4510,N_4704);
nor UO_301 (O_301,N_4669,N_4505);
or UO_302 (O_302,N_4796,N_4612);
or UO_303 (O_303,N_4872,N_4559);
nand UO_304 (O_304,N_4666,N_4566);
or UO_305 (O_305,N_4690,N_4762);
nor UO_306 (O_306,N_4815,N_4662);
nor UO_307 (O_307,N_4643,N_4881);
nand UO_308 (O_308,N_4655,N_4691);
nor UO_309 (O_309,N_4527,N_4703);
nand UO_310 (O_310,N_4597,N_4676);
nand UO_311 (O_311,N_4715,N_4948);
and UO_312 (O_312,N_4791,N_4557);
nor UO_313 (O_313,N_4634,N_4986);
and UO_314 (O_314,N_4746,N_4889);
nor UO_315 (O_315,N_4583,N_4559);
and UO_316 (O_316,N_4609,N_4823);
nor UO_317 (O_317,N_4680,N_4946);
nand UO_318 (O_318,N_4769,N_4618);
nor UO_319 (O_319,N_4515,N_4930);
nand UO_320 (O_320,N_4530,N_4881);
and UO_321 (O_321,N_4996,N_4864);
nand UO_322 (O_322,N_4971,N_4604);
nand UO_323 (O_323,N_4621,N_4874);
nor UO_324 (O_324,N_4645,N_4983);
or UO_325 (O_325,N_4696,N_4820);
nand UO_326 (O_326,N_4628,N_4592);
or UO_327 (O_327,N_4564,N_4932);
or UO_328 (O_328,N_4588,N_4563);
nand UO_329 (O_329,N_4677,N_4920);
and UO_330 (O_330,N_4761,N_4843);
nor UO_331 (O_331,N_4689,N_4866);
or UO_332 (O_332,N_4643,N_4796);
nand UO_333 (O_333,N_4817,N_4587);
nor UO_334 (O_334,N_4849,N_4710);
and UO_335 (O_335,N_4523,N_4669);
nand UO_336 (O_336,N_4961,N_4712);
and UO_337 (O_337,N_4821,N_4920);
nand UO_338 (O_338,N_4828,N_4625);
nor UO_339 (O_339,N_4576,N_4581);
and UO_340 (O_340,N_4601,N_4554);
nor UO_341 (O_341,N_4966,N_4804);
or UO_342 (O_342,N_4670,N_4926);
nor UO_343 (O_343,N_4668,N_4681);
nand UO_344 (O_344,N_4709,N_4590);
or UO_345 (O_345,N_4992,N_4574);
nand UO_346 (O_346,N_4839,N_4922);
or UO_347 (O_347,N_4713,N_4680);
and UO_348 (O_348,N_4638,N_4669);
nor UO_349 (O_349,N_4867,N_4863);
and UO_350 (O_350,N_4892,N_4883);
nor UO_351 (O_351,N_4549,N_4746);
and UO_352 (O_352,N_4957,N_4845);
or UO_353 (O_353,N_4872,N_4688);
nand UO_354 (O_354,N_4723,N_4940);
nor UO_355 (O_355,N_4753,N_4861);
nor UO_356 (O_356,N_4655,N_4617);
nor UO_357 (O_357,N_4523,N_4968);
and UO_358 (O_358,N_4573,N_4707);
or UO_359 (O_359,N_4881,N_4505);
nand UO_360 (O_360,N_4585,N_4571);
nor UO_361 (O_361,N_4895,N_4947);
or UO_362 (O_362,N_4613,N_4985);
nor UO_363 (O_363,N_4587,N_4977);
and UO_364 (O_364,N_4819,N_4833);
and UO_365 (O_365,N_4602,N_4687);
nand UO_366 (O_366,N_4999,N_4930);
and UO_367 (O_367,N_4835,N_4842);
nand UO_368 (O_368,N_4875,N_4892);
nand UO_369 (O_369,N_4760,N_4908);
nand UO_370 (O_370,N_4812,N_4962);
and UO_371 (O_371,N_4651,N_4900);
or UO_372 (O_372,N_4955,N_4720);
or UO_373 (O_373,N_4748,N_4649);
or UO_374 (O_374,N_4875,N_4945);
or UO_375 (O_375,N_4727,N_4937);
xnor UO_376 (O_376,N_4588,N_4710);
and UO_377 (O_377,N_4979,N_4928);
and UO_378 (O_378,N_4751,N_4900);
nand UO_379 (O_379,N_4955,N_4521);
or UO_380 (O_380,N_4993,N_4942);
and UO_381 (O_381,N_4710,N_4955);
xor UO_382 (O_382,N_4757,N_4934);
and UO_383 (O_383,N_4663,N_4828);
nor UO_384 (O_384,N_4601,N_4887);
and UO_385 (O_385,N_4647,N_4753);
nand UO_386 (O_386,N_4779,N_4580);
nand UO_387 (O_387,N_4812,N_4720);
nand UO_388 (O_388,N_4629,N_4590);
nand UO_389 (O_389,N_4814,N_4894);
nor UO_390 (O_390,N_4755,N_4812);
nand UO_391 (O_391,N_4953,N_4764);
and UO_392 (O_392,N_4667,N_4692);
nor UO_393 (O_393,N_4783,N_4865);
nor UO_394 (O_394,N_4627,N_4949);
and UO_395 (O_395,N_4582,N_4550);
or UO_396 (O_396,N_4565,N_4644);
and UO_397 (O_397,N_4537,N_4952);
nand UO_398 (O_398,N_4827,N_4828);
nor UO_399 (O_399,N_4751,N_4774);
nand UO_400 (O_400,N_4748,N_4866);
nand UO_401 (O_401,N_4547,N_4987);
and UO_402 (O_402,N_4747,N_4785);
nor UO_403 (O_403,N_4520,N_4956);
nor UO_404 (O_404,N_4556,N_4644);
nor UO_405 (O_405,N_4926,N_4707);
nand UO_406 (O_406,N_4770,N_4703);
nor UO_407 (O_407,N_4929,N_4533);
nand UO_408 (O_408,N_4720,N_4610);
and UO_409 (O_409,N_4521,N_4925);
or UO_410 (O_410,N_4827,N_4610);
or UO_411 (O_411,N_4590,N_4769);
or UO_412 (O_412,N_4759,N_4953);
or UO_413 (O_413,N_4976,N_4667);
and UO_414 (O_414,N_4841,N_4582);
and UO_415 (O_415,N_4675,N_4875);
nand UO_416 (O_416,N_4976,N_4977);
or UO_417 (O_417,N_4960,N_4984);
nor UO_418 (O_418,N_4951,N_4803);
nand UO_419 (O_419,N_4552,N_4617);
nand UO_420 (O_420,N_4706,N_4873);
nand UO_421 (O_421,N_4549,N_4560);
and UO_422 (O_422,N_4565,N_4534);
or UO_423 (O_423,N_4924,N_4836);
nor UO_424 (O_424,N_4739,N_4994);
nor UO_425 (O_425,N_4986,N_4637);
nand UO_426 (O_426,N_4732,N_4761);
nand UO_427 (O_427,N_4920,N_4577);
nor UO_428 (O_428,N_4809,N_4690);
nor UO_429 (O_429,N_4881,N_4681);
and UO_430 (O_430,N_4703,N_4728);
nor UO_431 (O_431,N_4523,N_4624);
nand UO_432 (O_432,N_4573,N_4535);
nand UO_433 (O_433,N_4658,N_4689);
and UO_434 (O_434,N_4522,N_4701);
xnor UO_435 (O_435,N_4733,N_4584);
and UO_436 (O_436,N_4953,N_4896);
nor UO_437 (O_437,N_4566,N_4930);
xor UO_438 (O_438,N_4901,N_4970);
or UO_439 (O_439,N_4714,N_4958);
or UO_440 (O_440,N_4714,N_4509);
nand UO_441 (O_441,N_4589,N_4631);
and UO_442 (O_442,N_4957,N_4510);
nand UO_443 (O_443,N_4607,N_4965);
nand UO_444 (O_444,N_4778,N_4585);
nand UO_445 (O_445,N_4931,N_4556);
nand UO_446 (O_446,N_4637,N_4744);
or UO_447 (O_447,N_4640,N_4884);
or UO_448 (O_448,N_4598,N_4846);
nand UO_449 (O_449,N_4670,N_4540);
and UO_450 (O_450,N_4995,N_4901);
and UO_451 (O_451,N_4575,N_4883);
or UO_452 (O_452,N_4858,N_4998);
nand UO_453 (O_453,N_4813,N_4632);
nand UO_454 (O_454,N_4572,N_4889);
or UO_455 (O_455,N_4876,N_4534);
nand UO_456 (O_456,N_4718,N_4815);
nor UO_457 (O_457,N_4819,N_4879);
nand UO_458 (O_458,N_4953,N_4521);
and UO_459 (O_459,N_4868,N_4609);
or UO_460 (O_460,N_4502,N_4576);
nor UO_461 (O_461,N_4860,N_4567);
or UO_462 (O_462,N_4771,N_4762);
and UO_463 (O_463,N_4815,N_4887);
and UO_464 (O_464,N_4747,N_4761);
nand UO_465 (O_465,N_4802,N_4793);
and UO_466 (O_466,N_4535,N_4780);
nand UO_467 (O_467,N_4509,N_4725);
nor UO_468 (O_468,N_4787,N_4500);
xnor UO_469 (O_469,N_4945,N_4839);
and UO_470 (O_470,N_4722,N_4655);
or UO_471 (O_471,N_4853,N_4709);
and UO_472 (O_472,N_4863,N_4541);
nand UO_473 (O_473,N_4621,N_4958);
or UO_474 (O_474,N_4733,N_4554);
nand UO_475 (O_475,N_4605,N_4887);
or UO_476 (O_476,N_4769,N_4832);
nor UO_477 (O_477,N_4982,N_4822);
nand UO_478 (O_478,N_4565,N_4800);
nand UO_479 (O_479,N_4857,N_4871);
nor UO_480 (O_480,N_4755,N_4920);
or UO_481 (O_481,N_4685,N_4634);
xnor UO_482 (O_482,N_4830,N_4943);
nand UO_483 (O_483,N_4815,N_4732);
nand UO_484 (O_484,N_4735,N_4649);
or UO_485 (O_485,N_4974,N_4899);
nor UO_486 (O_486,N_4915,N_4971);
or UO_487 (O_487,N_4664,N_4803);
nor UO_488 (O_488,N_4747,N_4880);
nor UO_489 (O_489,N_4580,N_4950);
or UO_490 (O_490,N_4500,N_4958);
or UO_491 (O_491,N_4866,N_4667);
or UO_492 (O_492,N_4667,N_4674);
or UO_493 (O_493,N_4962,N_4570);
or UO_494 (O_494,N_4613,N_4847);
or UO_495 (O_495,N_4766,N_4809);
and UO_496 (O_496,N_4579,N_4599);
nor UO_497 (O_497,N_4685,N_4889);
nor UO_498 (O_498,N_4985,N_4648);
nand UO_499 (O_499,N_4836,N_4630);
nand UO_500 (O_500,N_4871,N_4686);
nand UO_501 (O_501,N_4979,N_4879);
nand UO_502 (O_502,N_4936,N_4637);
nor UO_503 (O_503,N_4986,N_4708);
xor UO_504 (O_504,N_4677,N_4764);
nor UO_505 (O_505,N_4524,N_4767);
nand UO_506 (O_506,N_4987,N_4602);
or UO_507 (O_507,N_4957,N_4718);
or UO_508 (O_508,N_4638,N_4962);
nor UO_509 (O_509,N_4776,N_4739);
or UO_510 (O_510,N_4904,N_4736);
nor UO_511 (O_511,N_4861,N_4526);
and UO_512 (O_512,N_4849,N_4637);
and UO_513 (O_513,N_4672,N_4568);
nand UO_514 (O_514,N_4558,N_4569);
xor UO_515 (O_515,N_4592,N_4664);
xor UO_516 (O_516,N_4930,N_4523);
and UO_517 (O_517,N_4826,N_4573);
nor UO_518 (O_518,N_4655,N_4566);
and UO_519 (O_519,N_4997,N_4828);
or UO_520 (O_520,N_4639,N_4618);
and UO_521 (O_521,N_4615,N_4649);
or UO_522 (O_522,N_4912,N_4575);
or UO_523 (O_523,N_4575,N_4917);
and UO_524 (O_524,N_4877,N_4985);
and UO_525 (O_525,N_4954,N_4671);
nand UO_526 (O_526,N_4844,N_4690);
nand UO_527 (O_527,N_4526,N_4953);
and UO_528 (O_528,N_4691,N_4784);
nor UO_529 (O_529,N_4566,N_4896);
nand UO_530 (O_530,N_4637,N_4538);
and UO_531 (O_531,N_4763,N_4848);
nor UO_532 (O_532,N_4733,N_4969);
nor UO_533 (O_533,N_4546,N_4863);
nor UO_534 (O_534,N_4695,N_4928);
and UO_535 (O_535,N_4742,N_4515);
nor UO_536 (O_536,N_4689,N_4994);
and UO_537 (O_537,N_4709,N_4652);
and UO_538 (O_538,N_4987,N_4614);
or UO_539 (O_539,N_4738,N_4543);
or UO_540 (O_540,N_4718,N_4570);
nand UO_541 (O_541,N_4607,N_4519);
nor UO_542 (O_542,N_4513,N_4700);
nor UO_543 (O_543,N_4707,N_4845);
nand UO_544 (O_544,N_4793,N_4940);
nand UO_545 (O_545,N_4906,N_4840);
nor UO_546 (O_546,N_4762,N_4814);
nand UO_547 (O_547,N_4726,N_4754);
nor UO_548 (O_548,N_4686,N_4567);
and UO_549 (O_549,N_4791,N_4553);
and UO_550 (O_550,N_4554,N_4740);
or UO_551 (O_551,N_4554,N_4822);
or UO_552 (O_552,N_4562,N_4920);
and UO_553 (O_553,N_4898,N_4956);
and UO_554 (O_554,N_4501,N_4759);
nand UO_555 (O_555,N_4605,N_4565);
nand UO_556 (O_556,N_4585,N_4507);
nor UO_557 (O_557,N_4988,N_4687);
xnor UO_558 (O_558,N_4615,N_4573);
nand UO_559 (O_559,N_4536,N_4541);
nand UO_560 (O_560,N_4619,N_4838);
or UO_561 (O_561,N_4678,N_4991);
or UO_562 (O_562,N_4528,N_4894);
nor UO_563 (O_563,N_4773,N_4607);
nand UO_564 (O_564,N_4942,N_4616);
nand UO_565 (O_565,N_4641,N_4786);
and UO_566 (O_566,N_4959,N_4729);
or UO_567 (O_567,N_4683,N_4986);
nand UO_568 (O_568,N_4848,N_4820);
xnor UO_569 (O_569,N_4952,N_4894);
nor UO_570 (O_570,N_4526,N_4613);
xnor UO_571 (O_571,N_4770,N_4980);
and UO_572 (O_572,N_4782,N_4876);
nor UO_573 (O_573,N_4916,N_4834);
nand UO_574 (O_574,N_4592,N_4655);
and UO_575 (O_575,N_4952,N_4508);
and UO_576 (O_576,N_4600,N_4579);
and UO_577 (O_577,N_4611,N_4980);
and UO_578 (O_578,N_4757,N_4815);
nand UO_579 (O_579,N_4574,N_4810);
or UO_580 (O_580,N_4507,N_4575);
or UO_581 (O_581,N_4524,N_4778);
and UO_582 (O_582,N_4599,N_4690);
and UO_583 (O_583,N_4937,N_4561);
nor UO_584 (O_584,N_4738,N_4620);
or UO_585 (O_585,N_4928,N_4967);
or UO_586 (O_586,N_4948,N_4860);
or UO_587 (O_587,N_4943,N_4803);
nand UO_588 (O_588,N_4678,N_4683);
nor UO_589 (O_589,N_4920,N_4544);
nand UO_590 (O_590,N_4892,N_4972);
nor UO_591 (O_591,N_4948,N_4556);
nand UO_592 (O_592,N_4712,N_4883);
or UO_593 (O_593,N_4873,N_4807);
and UO_594 (O_594,N_4594,N_4737);
or UO_595 (O_595,N_4788,N_4623);
or UO_596 (O_596,N_4699,N_4516);
nor UO_597 (O_597,N_4918,N_4599);
nor UO_598 (O_598,N_4746,N_4664);
nor UO_599 (O_599,N_4856,N_4792);
or UO_600 (O_600,N_4831,N_4891);
and UO_601 (O_601,N_4857,N_4577);
nor UO_602 (O_602,N_4834,N_4866);
nor UO_603 (O_603,N_4554,N_4687);
and UO_604 (O_604,N_4804,N_4800);
nor UO_605 (O_605,N_4524,N_4637);
nor UO_606 (O_606,N_4895,N_4552);
nor UO_607 (O_607,N_4803,N_4814);
nor UO_608 (O_608,N_4514,N_4651);
or UO_609 (O_609,N_4820,N_4845);
or UO_610 (O_610,N_4596,N_4798);
nand UO_611 (O_611,N_4725,N_4644);
and UO_612 (O_612,N_4948,N_4869);
or UO_613 (O_613,N_4761,N_4905);
nand UO_614 (O_614,N_4654,N_4671);
or UO_615 (O_615,N_4848,N_4797);
or UO_616 (O_616,N_4614,N_4705);
nand UO_617 (O_617,N_4804,N_4740);
and UO_618 (O_618,N_4713,N_4640);
or UO_619 (O_619,N_4522,N_4986);
or UO_620 (O_620,N_4669,N_4703);
or UO_621 (O_621,N_4575,N_4547);
nor UO_622 (O_622,N_4875,N_4855);
nor UO_623 (O_623,N_4553,N_4761);
and UO_624 (O_624,N_4663,N_4877);
nor UO_625 (O_625,N_4905,N_4879);
nand UO_626 (O_626,N_4705,N_4717);
and UO_627 (O_627,N_4513,N_4833);
nor UO_628 (O_628,N_4714,N_4877);
or UO_629 (O_629,N_4622,N_4700);
or UO_630 (O_630,N_4676,N_4780);
and UO_631 (O_631,N_4535,N_4723);
or UO_632 (O_632,N_4791,N_4537);
nand UO_633 (O_633,N_4992,N_4912);
nor UO_634 (O_634,N_4594,N_4765);
nand UO_635 (O_635,N_4622,N_4653);
xor UO_636 (O_636,N_4752,N_4510);
and UO_637 (O_637,N_4693,N_4748);
or UO_638 (O_638,N_4575,N_4633);
nor UO_639 (O_639,N_4961,N_4931);
nand UO_640 (O_640,N_4802,N_4838);
nor UO_641 (O_641,N_4648,N_4585);
and UO_642 (O_642,N_4782,N_4998);
nand UO_643 (O_643,N_4785,N_4594);
nor UO_644 (O_644,N_4621,N_4639);
nand UO_645 (O_645,N_4766,N_4606);
and UO_646 (O_646,N_4565,N_4686);
nand UO_647 (O_647,N_4687,N_4847);
or UO_648 (O_648,N_4776,N_4977);
and UO_649 (O_649,N_4967,N_4632);
nand UO_650 (O_650,N_4563,N_4850);
xnor UO_651 (O_651,N_4654,N_4947);
nand UO_652 (O_652,N_4599,N_4590);
and UO_653 (O_653,N_4676,N_4614);
nor UO_654 (O_654,N_4990,N_4845);
nor UO_655 (O_655,N_4651,N_4683);
and UO_656 (O_656,N_4582,N_4781);
nand UO_657 (O_657,N_4744,N_4677);
and UO_658 (O_658,N_4523,N_4715);
nand UO_659 (O_659,N_4780,N_4957);
nand UO_660 (O_660,N_4900,N_4818);
or UO_661 (O_661,N_4582,N_4640);
nand UO_662 (O_662,N_4999,N_4663);
and UO_663 (O_663,N_4971,N_4631);
and UO_664 (O_664,N_4737,N_4967);
and UO_665 (O_665,N_4692,N_4907);
nand UO_666 (O_666,N_4605,N_4774);
or UO_667 (O_667,N_4846,N_4851);
nor UO_668 (O_668,N_4691,N_4563);
and UO_669 (O_669,N_4904,N_4549);
and UO_670 (O_670,N_4642,N_4727);
and UO_671 (O_671,N_4832,N_4706);
or UO_672 (O_672,N_4868,N_4948);
and UO_673 (O_673,N_4890,N_4865);
xnor UO_674 (O_674,N_4549,N_4995);
nor UO_675 (O_675,N_4598,N_4547);
or UO_676 (O_676,N_4766,N_4624);
nor UO_677 (O_677,N_4868,N_4564);
nand UO_678 (O_678,N_4804,N_4701);
or UO_679 (O_679,N_4982,N_4578);
or UO_680 (O_680,N_4820,N_4673);
or UO_681 (O_681,N_4706,N_4967);
and UO_682 (O_682,N_4935,N_4836);
or UO_683 (O_683,N_4907,N_4651);
or UO_684 (O_684,N_4964,N_4514);
and UO_685 (O_685,N_4962,N_4717);
and UO_686 (O_686,N_4811,N_4772);
or UO_687 (O_687,N_4556,N_4534);
nand UO_688 (O_688,N_4852,N_4756);
nand UO_689 (O_689,N_4731,N_4816);
or UO_690 (O_690,N_4975,N_4630);
nor UO_691 (O_691,N_4900,N_4873);
or UO_692 (O_692,N_4540,N_4886);
xnor UO_693 (O_693,N_4557,N_4880);
nand UO_694 (O_694,N_4928,N_4849);
xor UO_695 (O_695,N_4615,N_4852);
and UO_696 (O_696,N_4665,N_4560);
and UO_697 (O_697,N_4756,N_4816);
or UO_698 (O_698,N_4531,N_4642);
and UO_699 (O_699,N_4911,N_4522);
nor UO_700 (O_700,N_4836,N_4851);
or UO_701 (O_701,N_4652,N_4704);
nand UO_702 (O_702,N_4794,N_4966);
and UO_703 (O_703,N_4916,N_4737);
and UO_704 (O_704,N_4585,N_4686);
or UO_705 (O_705,N_4996,N_4553);
nand UO_706 (O_706,N_4742,N_4828);
and UO_707 (O_707,N_4760,N_4546);
or UO_708 (O_708,N_4800,N_4957);
and UO_709 (O_709,N_4841,N_4974);
and UO_710 (O_710,N_4800,N_4994);
and UO_711 (O_711,N_4881,N_4628);
and UO_712 (O_712,N_4605,N_4886);
nand UO_713 (O_713,N_4832,N_4652);
or UO_714 (O_714,N_4529,N_4653);
or UO_715 (O_715,N_4684,N_4577);
nand UO_716 (O_716,N_4653,N_4504);
or UO_717 (O_717,N_4747,N_4923);
nand UO_718 (O_718,N_4584,N_4503);
or UO_719 (O_719,N_4873,N_4912);
nand UO_720 (O_720,N_4899,N_4932);
and UO_721 (O_721,N_4967,N_4535);
or UO_722 (O_722,N_4954,N_4965);
and UO_723 (O_723,N_4798,N_4629);
and UO_724 (O_724,N_4643,N_4888);
nand UO_725 (O_725,N_4837,N_4635);
nor UO_726 (O_726,N_4830,N_4516);
xnor UO_727 (O_727,N_4852,N_4752);
and UO_728 (O_728,N_4780,N_4802);
nor UO_729 (O_729,N_4783,N_4921);
nand UO_730 (O_730,N_4543,N_4990);
nand UO_731 (O_731,N_4981,N_4686);
nor UO_732 (O_732,N_4707,N_4625);
nor UO_733 (O_733,N_4897,N_4762);
or UO_734 (O_734,N_4796,N_4726);
nand UO_735 (O_735,N_4644,N_4831);
and UO_736 (O_736,N_4817,N_4979);
and UO_737 (O_737,N_4774,N_4763);
nor UO_738 (O_738,N_4539,N_4662);
or UO_739 (O_739,N_4903,N_4706);
nand UO_740 (O_740,N_4574,N_4736);
and UO_741 (O_741,N_4922,N_4633);
nand UO_742 (O_742,N_4914,N_4722);
and UO_743 (O_743,N_4793,N_4993);
and UO_744 (O_744,N_4646,N_4669);
nor UO_745 (O_745,N_4764,N_4816);
and UO_746 (O_746,N_4653,N_4602);
nor UO_747 (O_747,N_4530,N_4922);
nand UO_748 (O_748,N_4655,N_4881);
or UO_749 (O_749,N_4680,N_4766);
nor UO_750 (O_750,N_4558,N_4859);
nand UO_751 (O_751,N_4703,N_4567);
or UO_752 (O_752,N_4617,N_4567);
nor UO_753 (O_753,N_4618,N_4795);
nor UO_754 (O_754,N_4781,N_4748);
or UO_755 (O_755,N_4503,N_4733);
and UO_756 (O_756,N_4988,N_4798);
nand UO_757 (O_757,N_4941,N_4949);
and UO_758 (O_758,N_4660,N_4500);
xor UO_759 (O_759,N_4572,N_4608);
and UO_760 (O_760,N_4768,N_4877);
and UO_761 (O_761,N_4761,N_4584);
nand UO_762 (O_762,N_4774,N_4790);
nand UO_763 (O_763,N_4617,N_4536);
and UO_764 (O_764,N_4861,N_4589);
or UO_765 (O_765,N_4525,N_4548);
and UO_766 (O_766,N_4823,N_4730);
nand UO_767 (O_767,N_4669,N_4641);
or UO_768 (O_768,N_4627,N_4868);
nor UO_769 (O_769,N_4996,N_4801);
nand UO_770 (O_770,N_4575,N_4960);
or UO_771 (O_771,N_4822,N_4718);
nand UO_772 (O_772,N_4554,N_4896);
nand UO_773 (O_773,N_4614,N_4808);
or UO_774 (O_774,N_4754,N_4937);
and UO_775 (O_775,N_4594,N_4813);
nand UO_776 (O_776,N_4543,N_4663);
nor UO_777 (O_777,N_4637,N_4845);
and UO_778 (O_778,N_4618,N_4601);
or UO_779 (O_779,N_4925,N_4623);
nand UO_780 (O_780,N_4966,N_4741);
nand UO_781 (O_781,N_4812,N_4944);
nand UO_782 (O_782,N_4687,N_4541);
nor UO_783 (O_783,N_4717,N_4609);
nor UO_784 (O_784,N_4637,N_4664);
or UO_785 (O_785,N_4927,N_4914);
nor UO_786 (O_786,N_4553,N_4503);
nand UO_787 (O_787,N_4964,N_4606);
and UO_788 (O_788,N_4515,N_4788);
nand UO_789 (O_789,N_4563,N_4581);
or UO_790 (O_790,N_4825,N_4785);
and UO_791 (O_791,N_4704,N_4611);
nand UO_792 (O_792,N_4566,N_4889);
and UO_793 (O_793,N_4997,N_4747);
and UO_794 (O_794,N_4945,N_4812);
nor UO_795 (O_795,N_4556,N_4574);
or UO_796 (O_796,N_4788,N_4508);
nand UO_797 (O_797,N_4542,N_4501);
nor UO_798 (O_798,N_4810,N_4818);
nor UO_799 (O_799,N_4610,N_4857);
or UO_800 (O_800,N_4639,N_4548);
or UO_801 (O_801,N_4702,N_4513);
nand UO_802 (O_802,N_4879,N_4947);
or UO_803 (O_803,N_4738,N_4966);
or UO_804 (O_804,N_4592,N_4864);
or UO_805 (O_805,N_4767,N_4618);
nand UO_806 (O_806,N_4748,N_4876);
nor UO_807 (O_807,N_4607,N_4977);
and UO_808 (O_808,N_4660,N_4861);
and UO_809 (O_809,N_4714,N_4643);
and UO_810 (O_810,N_4949,N_4683);
and UO_811 (O_811,N_4941,N_4974);
or UO_812 (O_812,N_4873,N_4688);
nor UO_813 (O_813,N_4515,N_4675);
or UO_814 (O_814,N_4887,N_4947);
nand UO_815 (O_815,N_4844,N_4923);
nor UO_816 (O_816,N_4631,N_4504);
nor UO_817 (O_817,N_4635,N_4715);
and UO_818 (O_818,N_4897,N_4955);
nor UO_819 (O_819,N_4776,N_4968);
nor UO_820 (O_820,N_4883,N_4811);
and UO_821 (O_821,N_4691,N_4845);
or UO_822 (O_822,N_4785,N_4523);
and UO_823 (O_823,N_4657,N_4577);
nand UO_824 (O_824,N_4583,N_4501);
or UO_825 (O_825,N_4956,N_4631);
xor UO_826 (O_826,N_4536,N_4690);
nor UO_827 (O_827,N_4570,N_4636);
or UO_828 (O_828,N_4710,N_4799);
nor UO_829 (O_829,N_4923,N_4976);
or UO_830 (O_830,N_4880,N_4670);
xnor UO_831 (O_831,N_4585,N_4514);
or UO_832 (O_832,N_4552,N_4978);
or UO_833 (O_833,N_4938,N_4917);
or UO_834 (O_834,N_4711,N_4725);
or UO_835 (O_835,N_4893,N_4516);
or UO_836 (O_836,N_4792,N_4668);
and UO_837 (O_837,N_4887,N_4629);
or UO_838 (O_838,N_4589,N_4516);
nand UO_839 (O_839,N_4795,N_4764);
nor UO_840 (O_840,N_4668,N_4708);
and UO_841 (O_841,N_4599,N_4946);
and UO_842 (O_842,N_4537,N_4605);
nor UO_843 (O_843,N_4997,N_4614);
or UO_844 (O_844,N_4551,N_4591);
and UO_845 (O_845,N_4688,N_4539);
nor UO_846 (O_846,N_4628,N_4997);
and UO_847 (O_847,N_4787,N_4622);
and UO_848 (O_848,N_4769,N_4873);
nor UO_849 (O_849,N_4527,N_4859);
xor UO_850 (O_850,N_4544,N_4883);
and UO_851 (O_851,N_4943,N_4773);
nand UO_852 (O_852,N_4827,N_4746);
nor UO_853 (O_853,N_4927,N_4620);
or UO_854 (O_854,N_4501,N_4889);
and UO_855 (O_855,N_4890,N_4658);
nand UO_856 (O_856,N_4810,N_4950);
or UO_857 (O_857,N_4772,N_4756);
nor UO_858 (O_858,N_4694,N_4828);
and UO_859 (O_859,N_4896,N_4647);
or UO_860 (O_860,N_4865,N_4842);
nor UO_861 (O_861,N_4532,N_4520);
nor UO_862 (O_862,N_4918,N_4669);
and UO_863 (O_863,N_4932,N_4650);
and UO_864 (O_864,N_4838,N_4777);
and UO_865 (O_865,N_4942,N_4587);
and UO_866 (O_866,N_4500,N_4687);
and UO_867 (O_867,N_4608,N_4813);
nor UO_868 (O_868,N_4929,N_4566);
nor UO_869 (O_869,N_4574,N_4588);
or UO_870 (O_870,N_4945,N_4516);
and UO_871 (O_871,N_4871,N_4670);
and UO_872 (O_872,N_4770,N_4811);
nor UO_873 (O_873,N_4719,N_4830);
and UO_874 (O_874,N_4977,N_4595);
nand UO_875 (O_875,N_4641,N_4579);
or UO_876 (O_876,N_4566,N_4921);
nand UO_877 (O_877,N_4685,N_4696);
or UO_878 (O_878,N_4639,N_4605);
or UO_879 (O_879,N_4513,N_4589);
nor UO_880 (O_880,N_4546,N_4735);
xor UO_881 (O_881,N_4838,N_4966);
or UO_882 (O_882,N_4554,N_4578);
or UO_883 (O_883,N_4659,N_4693);
or UO_884 (O_884,N_4575,N_4671);
nor UO_885 (O_885,N_4680,N_4919);
and UO_886 (O_886,N_4772,N_4885);
nand UO_887 (O_887,N_4932,N_4519);
nor UO_888 (O_888,N_4674,N_4561);
nor UO_889 (O_889,N_4945,N_4757);
or UO_890 (O_890,N_4868,N_4922);
or UO_891 (O_891,N_4804,N_4860);
or UO_892 (O_892,N_4631,N_4797);
nand UO_893 (O_893,N_4839,N_4792);
nand UO_894 (O_894,N_4842,N_4900);
nor UO_895 (O_895,N_4623,N_4755);
and UO_896 (O_896,N_4746,N_4742);
and UO_897 (O_897,N_4702,N_4668);
and UO_898 (O_898,N_4556,N_4789);
nand UO_899 (O_899,N_4827,N_4930);
nor UO_900 (O_900,N_4765,N_4773);
nor UO_901 (O_901,N_4649,N_4655);
nor UO_902 (O_902,N_4590,N_4808);
and UO_903 (O_903,N_4743,N_4910);
and UO_904 (O_904,N_4960,N_4962);
or UO_905 (O_905,N_4613,N_4592);
nor UO_906 (O_906,N_4721,N_4691);
or UO_907 (O_907,N_4682,N_4966);
nor UO_908 (O_908,N_4529,N_4807);
or UO_909 (O_909,N_4674,N_4926);
or UO_910 (O_910,N_4737,N_4859);
and UO_911 (O_911,N_4941,N_4664);
or UO_912 (O_912,N_4744,N_4985);
nand UO_913 (O_913,N_4772,N_4564);
or UO_914 (O_914,N_4615,N_4563);
nand UO_915 (O_915,N_4977,N_4602);
or UO_916 (O_916,N_4614,N_4795);
nand UO_917 (O_917,N_4758,N_4882);
or UO_918 (O_918,N_4660,N_4544);
nor UO_919 (O_919,N_4643,N_4758);
nand UO_920 (O_920,N_4702,N_4567);
nand UO_921 (O_921,N_4951,N_4994);
nand UO_922 (O_922,N_4941,N_4882);
and UO_923 (O_923,N_4922,N_4577);
nor UO_924 (O_924,N_4745,N_4880);
and UO_925 (O_925,N_4741,N_4958);
xnor UO_926 (O_926,N_4942,N_4918);
and UO_927 (O_927,N_4791,N_4884);
nor UO_928 (O_928,N_4665,N_4737);
and UO_929 (O_929,N_4885,N_4705);
nand UO_930 (O_930,N_4852,N_4522);
nand UO_931 (O_931,N_4806,N_4914);
and UO_932 (O_932,N_4883,N_4793);
and UO_933 (O_933,N_4627,N_4571);
nor UO_934 (O_934,N_4912,N_4776);
nor UO_935 (O_935,N_4707,N_4635);
or UO_936 (O_936,N_4844,N_4756);
or UO_937 (O_937,N_4789,N_4788);
nand UO_938 (O_938,N_4530,N_4722);
nor UO_939 (O_939,N_4564,N_4682);
nor UO_940 (O_940,N_4809,N_4914);
and UO_941 (O_941,N_4516,N_4865);
nor UO_942 (O_942,N_4853,N_4570);
nand UO_943 (O_943,N_4657,N_4950);
or UO_944 (O_944,N_4872,N_4750);
and UO_945 (O_945,N_4979,N_4941);
nor UO_946 (O_946,N_4774,N_4729);
or UO_947 (O_947,N_4958,N_4559);
nand UO_948 (O_948,N_4758,N_4611);
xnor UO_949 (O_949,N_4953,N_4716);
nor UO_950 (O_950,N_4854,N_4554);
or UO_951 (O_951,N_4709,N_4806);
nand UO_952 (O_952,N_4642,N_4820);
xor UO_953 (O_953,N_4803,N_4643);
nand UO_954 (O_954,N_4967,N_4717);
nor UO_955 (O_955,N_4866,N_4539);
nand UO_956 (O_956,N_4966,N_4510);
xnor UO_957 (O_957,N_4736,N_4585);
or UO_958 (O_958,N_4832,N_4744);
nand UO_959 (O_959,N_4714,N_4614);
nor UO_960 (O_960,N_4937,N_4911);
nor UO_961 (O_961,N_4704,N_4990);
and UO_962 (O_962,N_4713,N_4931);
and UO_963 (O_963,N_4529,N_4901);
or UO_964 (O_964,N_4847,N_4716);
or UO_965 (O_965,N_4645,N_4535);
or UO_966 (O_966,N_4785,N_4693);
nand UO_967 (O_967,N_4718,N_4539);
nor UO_968 (O_968,N_4748,N_4762);
nor UO_969 (O_969,N_4911,N_4945);
or UO_970 (O_970,N_4719,N_4775);
nor UO_971 (O_971,N_4607,N_4676);
and UO_972 (O_972,N_4569,N_4764);
and UO_973 (O_973,N_4588,N_4841);
nand UO_974 (O_974,N_4802,N_4955);
nand UO_975 (O_975,N_4662,N_4907);
nand UO_976 (O_976,N_4601,N_4692);
nor UO_977 (O_977,N_4672,N_4900);
and UO_978 (O_978,N_4877,N_4621);
nor UO_979 (O_979,N_4641,N_4730);
and UO_980 (O_980,N_4558,N_4737);
and UO_981 (O_981,N_4574,N_4508);
xnor UO_982 (O_982,N_4715,N_4535);
and UO_983 (O_983,N_4700,N_4910);
or UO_984 (O_984,N_4743,N_4735);
nor UO_985 (O_985,N_4831,N_4833);
or UO_986 (O_986,N_4777,N_4533);
or UO_987 (O_987,N_4978,N_4752);
nor UO_988 (O_988,N_4626,N_4846);
and UO_989 (O_989,N_4999,N_4925);
or UO_990 (O_990,N_4912,N_4895);
nor UO_991 (O_991,N_4634,N_4637);
or UO_992 (O_992,N_4914,N_4814);
and UO_993 (O_993,N_4718,N_4968);
nor UO_994 (O_994,N_4507,N_4782);
or UO_995 (O_995,N_4883,N_4741);
or UO_996 (O_996,N_4946,N_4973);
and UO_997 (O_997,N_4889,N_4595);
and UO_998 (O_998,N_4958,N_4571);
and UO_999 (O_999,N_4679,N_4773);
endmodule