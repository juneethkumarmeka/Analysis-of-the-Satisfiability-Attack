module basic_1000_10000_1500_20_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_755,In_101);
or U1 (N_1,In_27,In_576);
nand U2 (N_2,In_707,In_886);
nand U3 (N_3,In_650,In_443);
and U4 (N_4,In_590,In_750);
nor U5 (N_5,In_458,In_697);
nand U6 (N_6,In_641,In_669);
nand U7 (N_7,In_52,In_398);
or U8 (N_8,In_730,In_778);
nor U9 (N_9,In_912,In_162);
and U10 (N_10,In_579,In_46);
nand U11 (N_11,In_689,In_43);
nand U12 (N_12,In_905,In_935);
nand U13 (N_13,In_508,In_713);
or U14 (N_14,In_553,In_524);
nand U15 (N_15,In_676,In_878);
nand U16 (N_16,In_543,In_488);
nand U17 (N_17,In_188,In_725);
nor U18 (N_18,In_341,In_628);
nand U19 (N_19,In_933,In_966);
and U20 (N_20,In_603,In_996);
nor U21 (N_21,In_578,In_89);
nor U22 (N_22,In_678,In_313);
or U23 (N_23,In_120,In_840);
nand U24 (N_24,In_112,In_836);
and U25 (N_25,In_583,In_181);
and U26 (N_26,In_479,In_829);
or U27 (N_27,In_53,In_177);
nand U28 (N_28,In_139,In_586);
or U29 (N_29,In_946,In_584);
nand U30 (N_30,In_604,In_668);
and U31 (N_31,In_514,In_70);
or U32 (N_32,In_384,In_827);
xnor U33 (N_33,In_351,In_273);
nand U34 (N_34,In_263,In_42);
nand U35 (N_35,In_688,In_223);
nor U36 (N_36,In_38,In_11);
nand U37 (N_37,In_560,In_324);
or U38 (N_38,In_761,In_904);
xnor U39 (N_39,In_902,In_800);
or U40 (N_40,In_483,In_787);
nor U41 (N_41,In_719,In_471);
nand U42 (N_42,In_348,In_410);
and U43 (N_43,In_539,In_346);
nand U44 (N_44,In_985,In_216);
xnor U45 (N_45,In_503,In_360);
xor U46 (N_46,In_283,In_942);
nor U47 (N_47,In_805,In_964);
and U48 (N_48,In_1,In_659);
nor U49 (N_49,In_212,In_694);
nand U50 (N_50,In_848,In_489);
and U51 (N_51,In_357,In_298);
nor U52 (N_52,In_501,In_498);
xor U53 (N_53,In_986,In_815);
nand U54 (N_54,In_698,In_230);
nand U55 (N_55,In_484,In_679);
nand U56 (N_56,In_781,In_500);
or U57 (N_57,In_366,In_209);
nor U58 (N_58,In_531,In_981);
nor U59 (N_59,In_41,In_189);
and U60 (N_60,In_404,In_83);
nand U61 (N_61,In_782,In_548);
and U62 (N_62,In_322,In_444);
nand U63 (N_63,In_552,In_16);
or U64 (N_64,In_577,In_587);
or U65 (N_65,In_739,In_540);
or U66 (N_66,In_467,In_36);
nor U67 (N_67,In_460,In_627);
xnor U68 (N_68,In_474,In_285);
nor U69 (N_69,In_370,In_340);
or U70 (N_70,In_461,In_85);
or U71 (N_71,In_646,In_673);
or U72 (N_72,In_248,In_751);
and U73 (N_73,In_464,In_895);
nor U74 (N_74,In_839,In_279);
or U75 (N_75,In_930,In_447);
and U76 (N_76,In_561,In_862);
or U77 (N_77,In_870,In_541);
or U78 (N_78,In_394,In_103);
and U79 (N_79,In_670,In_795);
xnor U80 (N_80,In_21,In_924);
nand U81 (N_81,In_20,In_476);
and U82 (N_82,In_451,In_665);
nor U83 (N_83,In_907,In_264);
and U84 (N_84,In_12,In_417);
and U85 (N_85,In_256,In_148);
nand U86 (N_86,In_431,In_871);
and U87 (N_87,In_411,In_432);
or U88 (N_88,In_90,In_95);
nand U89 (N_89,In_801,In_413);
nand U90 (N_90,In_399,In_92);
nor U91 (N_91,In_824,In_622);
nor U92 (N_92,In_10,In_429);
or U93 (N_93,In_626,In_130);
nand U94 (N_94,In_408,In_314);
nand U95 (N_95,In_94,In_851);
or U96 (N_96,In_378,In_359);
nor U97 (N_97,In_412,In_822);
or U98 (N_98,In_271,In_395);
and U99 (N_99,In_18,In_149);
nor U100 (N_100,In_915,In_232);
nand U101 (N_101,In_845,In_506);
and U102 (N_102,In_485,In_956);
or U103 (N_103,In_73,In_200);
or U104 (N_104,In_396,In_535);
nand U105 (N_105,In_407,In_282);
nand U106 (N_106,In_423,In_393);
nor U107 (N_107,In_262,In_362);
or U108 (N_108,In_61,In_455);
and U109 (N_109,In_704,In_463);
xnor U110 (N_110,In_126,In_969);
nand U111 (N_111,In_178,In_846);
nand U112 (N_112,In_601,In_316);
or U113 (N_113,In_909,In_140);
nor U114 (N_114,In_147,In_733);
or U115 (N_115,In_754,In_23);
nor U116 (N_116,In_437,In_660);
and U117 (N_117,In_142,In_50);
and U118 (N_118,In_480,In_244);
or U119 (N_119,In_299,In_206);
nand U120 (N_120,In_328,In_816);
or U121 (N_121,In_616,In_826);
or U122 (N_122,In_242,In_452);
nand U123 (N_123,In_786,In_374);
xnor U124 (N_124,In_714,In_179);
nand U125 (N_125,In_596,In_325);
nor U126 (N_126,In_847,In_170);
or U127 (N_127,In_40,In_903);
and U128 (N_128,In_236,In_887);
and U129 (N_129,In_486,In_893);
nor U130 (N_130,In_172,In_640);
xor U131 (N_131,In_819,In_572);
nand U132 (N_132,In_368,In_699);
nand U133 (N_133,In_208,In_286);
nor U134 (N_134,In_65,In_278);
nand U135 (N_135,In_758,In_997);
nand U136 (N_136,In_387,In_834);
or U137 (N_137,In_849,In_833);
xor U138 (N_138,In_537,In_250);
or U139 (N_139,In_775,In_898);
nor U140 (N_140,In_84,In_723);
and U141 (N_141,In_96,In_550);
nor U142 (N_142,In_375,In_692);
or U143 (N_143,In_854,In_643);
nand U144 (N_144,In_502,In_218);
or U145 (N_145,In_219,In_88);
or U146 (N_146,In_133,In_803);
nor U147 (N_147,In_740,In_320);
and U148 (N_148,In_722,In_495);
or U149 (N_149,In_617,In_418);
nor U150 (N_150,In_174,In_873);
nand U151 (N_151,In_857,In_465);
or U152 (N_152,In_490,In_303);
nor U153 (N_153,In_134,In_598);
nand U154 (N_154,In_970,In_309);
and U155 (N_155,In_861,In_306);
or U156 (N_156,In_770,In_589);
nor U157 (N_157,In_630,In_13);
nor U158 (N_158,In_118,In_321);
nand U159 (N_159,In_386,In_760);
nand U160 (N_160,In_406,In_482);
nand U161 (N_161,In_735,In_439);
nand U162 (N_162,In_908,In_239);
nand U163 (N_163,In_204,In_233);
and U164 (N_164,In_512,In_762);
nand U165 (N_165,In_339,In_76);
nor U166 (N_166,In_457,In_390);
nor U167 (N_167,In_425,In_235);
xnor U168 (N_168,In_156,In_509);
nor U169 (N_169,In_599,In_806);
or U170 (N_170,In_5,In_664);
or U171 (N_171,In_241,In_881);
nor U172 (N_172,In_654,In_110);
and U173 (N_173,In_213,In_292);
or U174 (N_174,In_98,In_333);
or U175 (N_175,In_113,In_810);
or U176 (N_176,In_927,In_54);
nand U177 (N_177,In_753,In_135);
or U178 (N_178,In_459,In_247);
nor U179 (N_179,In_534,In_513);
xor U180 (N_180,In_825,In_337);
and U181 (N_181,In_568,In_349);
xnor U182 (N_182,In_789,In_549);
and U183 (N_183,In_675,In_127);
nor U184 (N_184,In_72,In_75);
nor U185 (N_185,In_45,In_334);
and U186 (N_186,In_493,In_949);
xor U187 (N_187,In_690,In_746);
nand U188 (N_188,In_645,In_655);
or U189 (N_189,In_661,In_709);
or U190 (N_190,In_69,In_528);
or U191 (N_191,In_975,In_693);
or U192 (N_192,In_987,In_807);
nor U193 (N_193,In_582,In_131);
nand U194 (N_194,In_545,In_859);
nor U195 (N_195,In_352,In_995);
nor U196 (N_196,In_154,In_542);
nand U197 (N_197,In_581,In_117);
nand U198 (N_198,In_97,In_729);
xor U199 (N_199,In_663,In_365);
xor U200 (N_200,In_82,In_648);
nor U201 (N_201,In_635,In_294);
and U202 (N_202,In_115,In_892);
or U203 (N_203,In_748,In_427);
nor U204 (N_204,In_379,In_757);
nor U205 (N_205,In_420,In_295);
nand U206 (N_206,In_56,In_965);
or U207 (N_207,In_104,In_402);
xnor U208 (N_208,In_510,In_342);
xor U209 (N_209,In_944,In_202);
nor U210 (N_210,In_214,In_547);
nand U211 (N_211,In_973,In_642);
nand U212 (N_212,In_151,In_380);
or U213 (N_213,In_22,In_565);
nor U214 (N_214,In_477,In_153);
or U215 (N_215,In_100,In_980);
nand U216 (N_216,In_732,In_637);
or U217 (N_217,In_122,In_877);
nand U218 (N_218,In_446,In_132);
and U219 (N_219,In_564,In_916);
or U220 (N_220,In_287,In_33);
and U221 (N_221,In_945,In_428);
or U222 (N_222,In_367,In_950);
nor U223 (N_223,In_632,In_240);
or U224 (N_224,In_989,In_60);
and U225 (N_225,In_338,In_718);
nand U226 (N_226,In_918,In_369);
nor U227 (N_227,In_731,In_491);
nor U228 (N_228,In_392,In_487);
nor U229 (N_229,In_926,In_720);
and U230 (N_230,In_64,In_880);
nor U231 (N_231,In_830,In_813);
or U232 (N_232,In_738,In_624);
nand U233 (N_233,In_363,In_835);
or U234 (N_234,In_968,In_958);
nand U235 (N_235,In_614,In_726);
nand U236 (N_236,In_456,In_959);
xor U237 (N_237,In_260,In_809);
nand U238 (N_238,In_941,In_921);
nand U239 (N_239,In_184,In_728);
and U240 (N_240,In_14,In_137);
or U241 (N_241,In_672,In_288);
or U242 (N_242,In_961,In_529);
or U243 (N_243,In_421,In_507);
nand U244 (N_244,In_37,In_121);
or U245 (N_245,In_66,In_194);
and U246 (N_246,In_74,In_414);
and U247 (N_247,In_435,In_925);
or U248 (N_248,In_466,In_255);
or U249 (N_249,In_867,In_215);
or U250 (N_250,In_114,In_585);
nor U251 (N_251,In_814,In_607);
nor U252 (N_252,In_159,In_792);
and U253 (N_253,In_703,In_163);
or U254 (N_254,In_505,In_119);
or U255 (N_255,In_526,In_424);
and U256 (N_256,In_323,In_784);
nor U257 (N_257,In_221,In_998);
xor U258 (N_258,In_554,In_332);
nand U259 (N_259,In_19,In_677);
and U260 (N_260,In_150,In_558);
nand U261 (N_261,In_680,In_785);
or U262 (N_262,In_138,In_928);
nand U263 (N_263,In_319,In_169);
or U264 (N_264,In_35,In_290);
nand U265 (N_265,In_963,In_780);
nor U266 (N_266,In_329,In_793);
xor U267 (N_267,In_207,In_710);
nor U268 (N_268,In_331,In_875);
or U269 (N_269,In_812,In_796);
nand U270 (N_270,In_666,In_518);
or U271 (N_271,In_727,In_81);
nor U272 (N_272,In_195,In_494);
nor U273 (N_273,In_844,In_804);
and U274 (N_274,In_939,In_571);
and U275 (N_275,In_934,In_951);
or U276 (N_276,In_237,In_953);
nand U277 (N_277,In_797,In_312);
and U278 (N_278,In_521,In_936);
nand U279 (N_279,In_940,In_6);
and U280 (N_280,In_350,In_91);
nand U281 (N_281,In_261,In_695);
nor U282 (N_282,In_982,In_275);
nand U283 (N_283,In_289,In_343);
nand U284 (N_284,In_656,In_606);
nand U285 (N_285,In_382,In_201);
or U286 (N_286,In_176,In_192);
nor U287 (N_287,In_225,In_744);
nor U288 (N_288,In_838,In_304);
or U289 (N_289,In_28,In_745);
nor U290 (N_290,In_8,In_284);
and U291 (N_291,In_625,In_633);
and U292 (N_292,In_802,In_621);
nor U293 (N_293,In_575,In_522);
nor U294 (N_294,In_954,In_619);
nor U295 (N_295,In_696,In_922);
xor U296 (N_296,In_224,In_318);
nor U297 (N_297,In_449,In_496);
or U298 (N_298,In_899,In_798);
nor U299 (N_299,In_371,In_865);
nand U300 (N_300,In_869,In_492);
nand U301 (N_301,In_884,In_258);
or U302 (N_302,In_765,In_741);
nor U303 (N_303,In_409,In_674);
nand U304 (N_304,In_266,In_611);
or U305 (N_305,In_345,In_106);
nor U306 (N_306,In_856,In_469);
and U307 (N_307,In_281,In_769);
and U308 (N_308,In_734,In_715);
nand U309 (N_309,In_419,In_3);
and U310 (N_310,In_377,In_948);
nor U311 (N_311,In_914,In_817);
and U312 (N_312,In_952,In_251);
or U313 (N_313,In_853,In_164);
or U314 (N_314,In_876,In_634);
nand U315 (N_315,In_280,In_57);
xor U316 (N_316,In_516,In_882);
or U317 (N_317,In_708,In_55);
and U318 (N_318,In_852,In_855);
or U319 (N_319,In_58,In_124);
nand U320 (N_320,In_533,In_270);
nor U321 (N_321,In_187,In_183);
nor U322 (N_322,In_570,In_504);
and U323 (N_323,In_992,In_311);
or U324 (N_324,In_62,In_711);
nor U325 (N_325,In_600,In_647);
nand U326 (N_326,In_450,In_358);
nand U327 (N_327,In_984,In_268);
nand U328 (N_328,In_706,In_977);
or U329 (N_329,In_551,In_681);
nand U330 (N_330,In_34,In_821);
and U331 (N_331,In_228,In_841);
and U332 (N_332,In_71,In_910);
and U333 (N_333,In_145,In_434);
nor U334 (N_334,In_957,In_649);
or U335 (N_335,In_771,In_631);
nor U336 (N_336,In_974,In_897);
and U337 (N_337,In_297,In_597);
or U338 (N_338,In_900,In_252);
nor U339 (N_339,In_426,In_511);
or U340 (N_340,In_983,In_197);
and U341 (N_341,In_629,In_129);
or U342 (N_342,In_705,In_49);
nand U343 (N_343,In_198,In_779);
or U344 (N_344,In_685,In_296);
nand U345 (N_345,In_161,In_227);
nand U346 (N_346,In_267,In_837);
and U347 (N_347,In_310,In_315);
or U348 (N_348,In_519,In_691);
and U349 (N_349,In_759,In_17);
or U350 (N_350,In_4,In_749);
nand U351 (N_351,In_453,In_454);
nand U352 (N_352,In_919,In_277);
or U353 (N_353,In_932,In_874);
xor U354 (N_354,In_355,In_473);
nand U355 (N_355,In_863,In_243);
nor U356 (N_356,In_994,In_422);
nor U357 (N_357,In_917,In_116);
and U358 (N_358,In_108,In_879);
or U359 (N_359,In_971,In_595);
and U360 (N_360,In_51,In_667);
nor U361 (N_361,In_580,In_109);
or U362 (N_362,In_712,In_858);
nor U363 (N_363,In_107,In_864);
nor U364 (N_364,In_405,In_823);
and U365 (N_365,In_307,In_608);
nor U366 (N_366,In_440,In_210);
nor U367 (N_367,In_86,In_373);
or U368 (N_368,In_217,In_790);
nand U369 (N_369,In_48,In_756);
nor U370 (N_370,In_136,In_885);
nor U371 (N_371,In_143,In_185);
and U372 (N_372,In_684,In_77);
or U373 (N_373,In_818,In_475);
nor U374 (N_374,In_525,In_574);
or U375 (N_375,In_566,In_229);
or U376 (N_376,In_913,In_636);
nor U377 (N_377,In_653,In_671);
or U378 (N_378,In_389,In_63);
and U379 (N_379,In_774,In_31);
or U380 (N_380,In_620,In_354);
and U381 (N_381,In_220,In_436);
nor U382 (N_382,In_272,In_901);
and U383 (N_383,In_385,In_9);
nor U384 (N_384,In_923,In_850);
nor U385 (N_385,In_190,In_445);
or U386 (N_386,In_573,In_752);
nand U387 (N_387,In_929,In_972);
nor U388 (N_388,In_364,In_356);
nand U389 (N_389,In_544,In_976);
nand U390 (N_390,In_191,In_766);
nor U391 (N_391,In_173,In_246);
or U392 (N_392,In_125,In_743);
and U393 (N_393,In_828,In_93);
nand U394 (N_394,In_683,In_610);
xor U395 (N_395,In_569,In_555);
and U396 (N_396,In_532,In_152);
and U397 (N_397,In_920,In_438);
and U398 (N_398,In_894,In_591);
and U399 (N_399,In_559,In_39);
xor U400 (N_400,In_615,In_468);
nand U401 (N_401,In_196,In_888);
nand U402 (N_402,In_254,In_317);
nand U403 (N_403,In_556,In_716);
nor U404 (N_404,In_794,In_890);
and U405 (N_405,In_943,In_274);
nand U406 (N_406,In_80,In_168);
or U407 (N_407,In_144,In_978);
or U408 (N_408,In_563,In_433);
and U409 (N_409,In_896,In_257);
xnor U410 (N_410,In_300,In_991);
or U411 (N_411,In_687,In_7);
nand U412 (N_412,In_265,In_231);
nand U413 (N_413,In_777,In_376);
nand U414 (N_414,In_737,In_523);
and U415 (N_415,In_400,In_175);
nand U416 (N_416,In_166,In_520);
nor U417 (N_417,In_146,In_517);
nand U418 (N_418,In_401,In_160);
nor U419 (N_419,In_165,In_658);
nor U420 (N_420,In_605,In_763);
nand U421 (N_421,In_906,In_831);
or U422 (N_422,In_682,In_245);
or U423 (N_423,In_768,In_613);
nand U424 (N_424,In_128,In_736);
nor U425 (N_425,In_609,In_481);
nor U426 (N_426,In_889,In_742);
or U427 (N_427,In_592,In_843);
or U428 (N_428,In_527,In_403);
or U429 (N_429,In_955,In_193);
nand U430 (N_430,In_87,In_335);
nor U431 (N_431,In_623,In_155);
or U432 (N_432,In_868,In_947);
and U433 (N_433,In_811,In_747);
or U434 (N_434,In_962,In_68);
nand U435 (N_435,In_259,In_472);
nor U436 (N_436,In_788,In_562);
nand U437 (N_437,In_866,In_883);
nand U438 (N_438,In_416,In_353);
nor U439 (N_439,In_302,In_442);
nand U440 (N_440,In_639,In_515);
or U441 (N_441,In_700,In_499);
or U442 (N_442,In_291,In_47);
nor U443 (N_443,In_26,In_618);
nor U444 (N_444,In_462,In_347);
nor U445 (N_445,In_249,In_808);
or U446 (N_446,In_293,In_24);
and U447 (N_447,In_203,In_967);
nand U448 (N_448,In_2,In_330);
nor U449 (N_449,In_791,In_651);
nand U450 (N_450,In_538,In_171);
nor U451 (N_451,In_724,In_105);
nor U452 (N_452,In_764,In_326);
and U453 (N_453,In_701,In_721);
and U454 (N_454,In_594,In_783);
or U455 (N_455,In_842,In_772);
nand U456 (N_456,In_536,In_657);
and U457 (N_457,In_123,In_29);
nor U458 (N_458,In_99,In_344);
or U459 (N_459,In_397,In_182);
nand U460 (N_460,In_717,In_226);
and U461 (N_461,In_820,In_391);
or U462 (N_462,In_911,In_59);
nand U463 (N_463,In_530,In_832);
nor U464 (N_464,In_993,In_860);
nand U465 (N_465,In_301,In_336);
or U466 (N_466,In_15,In_662);
or U467 (N_467,In_931,In_470);
or U468 (N_468,In_30,In_567);
and U469 (N_469,In_478,In_872);
nand U470 (N_470,In_638,In_238);
nor U471 (N_471,In_111,In_686);
nand U472 (N_472,In_78,In_0);
nand U473 (N_473,In_186,In_305);
nor U474 (N_474,In_546,In_102);
or U475 (N_475,In_588,In_497);
xor U476 (N_476,In_157,In_67);
nand U477 (N_477,In_767,In_799);
nor U478 (N_478,In_211,In_199);
nor U479 (N_479,In_938,In_388);
and U480 (N_480,In_644,In_891);
and U481 (N_481,In_773,In_276);
nor U482 (N_482,In_593,In_372);
nor U483 (N_483,In_234,In_141);
nand U484 (N_484,In_960,In_180);
nand U485 (N_485,In_430,In_222);
nor U486 (N_486,In_441,In_557);
nand U487 (N_487,In_937,In_988);
and U488 (N_488,In_327,In_44);
or U489 (N_489,In_205,In_448);
nand U490 (N_490,In_361,In_253);
and U491 (N_491,In_308,In_979);
or U492 (N_492,In_702,In_25);
nand U493 (N_493,In_269,In_79);
xnor U494 (N_494,In_167,In_383);
nand U495 (N_495,In_612,In_415);
nor U496 (N_496,In_381,In_158);
and U497 (N_497,In_652,In_602);
nor U498 (N_498,In_32,In_776);
nor U499 (N_499,In_990,In_999);
and U500 (N_500,N_295,N_423);
nor U501 (N_501,N_86,N_268);
or U502 (N_502,N_139,N_461);
or U503 (N_503,N_89,N_110);
or U504 (N_504,N_364,N_55);
nor U505 (N_505,N_355,N_68);
nand U506 (N_506,N_272,N_386);
nand U507 (N_507,N_486,N_450);
or U508 (N_508,N_121,N_326);
or U509 (N_509,N_494,N_77);
or U510 (N_510,N_356,N_490);
and U511 (N_511,N_84,N_399);
nor U512 (N_512,N_368,N_344);
or U513 (N_513,N_307,N_444);
and U514 (N_514,N_184,N_473);
nor U515 (N_515,N_384,N_303);
or U516 (N_516,N_449,N_391);
or U517 (N_517,N_103,N_111);
and U518 (N_518,N_32,N_238);
nor U519 (N_519,N_403,N_443);
nor U520 (N_520,N_151,N_148);
xor U521 (N_521,N_446,N_117);
and U522 (N_522,N_210,N_59);
and U523 (N_523,N_310,N_434);
nand U524 (N_524,N_369,N_7);
and U525 (N_525,N_455,N_476);
and U526 (N_526,N_388,N_253);
nor U527 (N_527,N_281,N_235);
and U528 (N_528,N_414,N_173);
and U529 (N_529,N_123,N_390);
nand U530 (N_530,N_379,N_229);
or U531 (N_531,N_36,N_27);
or U532 (N_532,N_319,N_382);
or U533 (N_533,N_69,N_149);
nand U534 (N_534,N_201,N_362);
or U535 (N_535,N_257,N_31);
and U536 (N_536,N_381,N_130);
nand U537 (N_537,N_311,N_453);
or U538 (N_538,N_339,N_158);
nand U539 (N_539,N_366,N_26);
nand U540 (N_540,N_65,N_10);
nor U541 (N_541,N_8,N_135);
or U542 (N_542,N_291,N_419);
nor U543 (N_543,N_394,N_39);
nand U544 (N_544,N_258,N_371);
or U545 (N_545,N_109,N_165);
nor U546 (N_546,N_346,N_197);
nand U547 (N_547,N_312,N_246);
or U548 (N_548,N_13,N_144);
nand U549 (N_549,N_38,N_383);
and U550 (N_550,N_285,N_408);
and U551 (N_551,N_485,N_199);
and U552 (N_552,N_497,N_207);
or U553 (N_553,N_420,N_79);
and U554 (N_554,N_83,N_251);
nand U555 (N_555,N_466,N_236);
nor U556 (N_556,N_283,N_270);
or U557 (N_557,N_498,N_249);
and U558 (N_558,N_416,N_47);
nor U559 (N_559,N_88,N_266);
nor U560 (N_560,N_70,N_133);
and U561 (N_561,N_67,N_357);
and U562 (N_562,N_113,N_341);
nor U563 (N_563,N_3,N_24);
or U564 (N_564,N_457,N_180);
nor U565 (N_565,N_194,N_465);
nand U566 (N_566,N_361,N_392);
nand U567 (N_567,N_256,N_489);
and U568 (N_568,N_264,N_273);
nand U569 (N_569,N_178,N_183);
or U570 (N_570,N_101,N_499);
xor U571 (N_571,N_128,N_20);
nand U572 (N_572,N_374,N_153);
or U573 (N_573,N_452,N_134);
and U574 (N_574,N_395,N_492);
and U575 (N_575,N_202,N_234);
or U576 (N_576,N_6,N_138);
or U577 (N_577,N_49,N_370);
or U578 (N_578,N_198,N_46);
nand U579 (N_579,N_299,N_54);
nand U580 (N_580,N_318,N_222);
nand U581 (N_581,N_402,N_66);
or U582 (N_582,N_116,N_432);
xnor U583 (N_583,N_214,N_34);
nor U584 (N_584,N_274,N_112);
and U585 (N_585,N_367,N_422);
nor U586 (N_586,N_174,N_204);
or U587 (N_587,N_12,N_407);
nand U588 (N_588,N_484,N_331);
nor U589 (N_589,N_206,N_470);
xor U590 (N_590,N_475,N_263);
xnor U591 (N_591,N_171,N_433);
and U592 (N_592,N_411,N_172);
or U593 (N_593,N_271,N_43);
nor U594 (N_594,N_195,N_82);
and U595 (N_595,N_301,N_211);
and U596 (N_596,N_168,N_333);
and U597 (N_597,N_146,N_150);
or U598 (N_598,N_231,N_205);
and U599 (N_599,N_438,N_290);
nand U600 (N_600,N_320,N_136);
or U601 (N_601,N_64,N_413);
or U602 (N_602,N_445,N_440);
nor U603 (N_603,N_353,N_17);
nand U604 (N_604,N_358,N_293);
nand U605 (N_605,N_375,N_21);
nand U606 (N_606,N_418,N_480);
and U607 (N_607,N_230,N_488);
nand U608 (N_608,N_309,N_430);
and U609 (N_609,N_305,N_481);
or U610 (N_610,N_247,N_218);
or U611 (N_611,N_426,N_226);
nand U612 (N_612,N_286,N_163);
nand U613 (N_613,N_460,N_314);
nor U614 (N_614,N_23,N_275);
nand U615 (N_615,N_188,N_196);
nor U616 (N_616,N_471,N_294);
nand U617 (N_617,N_169,N_306);
nand U618 (N_618,N_406,N_53);
nand U619 (N_619,N_260,N_477);
nand U620 (N_620,N_254,N_217);
xor U621 (N_621,N_487,N_332);
nor U622 (N_622,N_267,N_131);
and U623 (N_623,N_107,N_115);
nor U624 (N_624,N_51,N_252);
nor U625 (N_625,N_335,N_127);
or U626 (N_626,N_142,N_462);
nor U627 (N_627,N_209,N_304);
or U628 (N_628,N_122,N_345);
nor U629 (N_629,N_323,N_324);
nand U630 (N_630,N_192,N_448);
and U631 (N_631,N_57,N_15);
and U632 (N_632,N_317,N_170);
nand U633 (N_633,N_493,N_190);
nand U634 (N_634,N_189,N_308);
nor U635 (N_635,N_467,N_316);
nor U636 (N_636,N_92,N_396);
or U637 (N_637,N_97,N_321);
or U638 (N_638,N_336,N_94);
or U639 (N_639,N_200,N_297);
nand U640 (N_640,N_11,N_187);
nand U641 (N_641,N_50,N_237);
nor U642 (N_642,N_398,N_126);
and U643 (N_643,N_108,N_152);
and U644 (N_644,N_141,N_428);
and U645 (N_645,N_223,N_387);
nor U646 (N_646,N_262,N_389);
and U647 (N_647,N_104,N_224);
and U648 (N_648,N_292,N_227);
nor U649 (N_649,N_417,N_330);
nor U650 (N_650,N_327,N_186);
and U651 (N_651,N_373,N_63);
or U652 (N_652,N_380,N_41);
nor U653 (N_653,N_240,N_482);
nor U654 (N_654,N_185,N_228);
and U655 (N_655,N_491,N_87);
xnor U656 (N_656,N_298,N_114);
nand U657 (N_657,N_410,N_447);
xnor U658 (N_658,N_162,N_56);
nand U659 (N_659,N_5,N_159);
nand U660 (N_660,N_284,N_348);
and U661 (N_661,N_359,N_242);
nor U662 (N_662,N_378,N_459);
or U663 (N_663,N_145,N_175);
or U664 (N_664,N_393,N_289);
or U665 (N_665,N_14,N_424);
nand U666 (N_666,N_81,N_322);
nor U667 (N_667,N_102,N_95);
or U668 (N_668,N_80,N_161);
nand U669 (N_669,N_90,N_456);
and U670 (N_670,N_243,N_255);
nor U671 (N_671,N_349,N_400);
nand U672 (N_672,N_415,N_313);
nor U673 (N_673,N_239,N_33);
nand U674 (N_674,N_377,N_119);
nand U675 (N_675,N_125,N_61);
nand U676 (N_676,N_1,N_451);
xnor U677 (N_677,N_100,N_360);
or U678 (N_678,N_248,N_421);
or U679 (N_679,N_435,N_96);
and U680 (N_680,N_454,N_468);
nor U681 (N_681,N_176,N_37);
nor U682 (N_682,N_212,N_129);
or U683 (N_683,N_179,N_425);
xnor U684 (N_684,N_437,N_372);
and U685 (N_685,N_350,N_220);
and U686 (N_686,N_85,N_340);
and U687 (N_687,N_215,N_405);
nor U688 (N_688,N_203,N_265);
or U689 (N_689,N_436,N_397);
or U690 (N_690,N_155,N_35);
or U691 (N_691,N_282,N_181);
nor U692 (N_692,N_431,N_60);
and U693 (N_693,N_329,N_164);
nor U694 (N_694,N_48,N_52);
nand U695 (N_695,N_132,N_269);
or U696 (N_696,N_412,N_479);
nand U697 (N_697,N_337,N_363);
nand U698 (N_698,N_105,N_458);
or U699 (N_699,N_118,N_58);
nor U700 (N_700,N_72,N_296);
nor U701 (N_701,N_124,N_75);
or U702 (N_702,N_338,N_343);
and U703 (N_703,N_4,N_9);
nor U704 (N_704,N_167,N_137);
and U705 (N_705,N_280,N_351);
nand U706 (N_706,N_29,N_427);
and U707 (N_707,N_28,N_385);
nor U708 (N_708,N_19,N_22);
and U709 (N_709,N_365,N_44);
or U710 (N_710,N_140,N_245);
nand U711 (N_711,N_442,N_474);
nand U712 (N_712,N_232,N_472);
nand U713 (N_713,N_496,N_334);
and U714 (N_714,N_160,N_276);
nand U715 (N_715,N_120,N_78);
nand U716 (N_716,N_241,N_495);
nand U717 (N_717,N_193,N_91);
and U718 (N_718,N_62,N_2);
and U719 (N_719,N_287,N_225);
nor U720 (N_720,N_71,N_213);
xnor U721 (N_721,N_464,N_208);
and U722 (N_722,N_0,N_478);
or U723 (N_723,N_328,N_376);
nand U724 (N_724,N_99,N_279);
nand U725 (N_725,N_45,N_221);
and U726 (N_726,N_463,N_352);
and U727 (N_727,N_233,N_325);
nor U728 (N_728,N_300,N_250);
and U729 (N_729,N_439,N_469);
or U730 (N_730,N_404,N_288);
and U731 (N_731,N_441,N_354);
nor U732 (N_732,N_42,N_106);
xor U733 (N_733,N_18,N_261);
xnor U734 (N_734,N_166,N_347);
nand U735 (N_735,N_278,N_74);
nand U736 (N_736,N_259,N_315);
nand U737 (N_737,N_409,N_483);
nor U738 (N_738,N_277,N_429);
or U739 (N_739,N_157,N_143);
and U740 (N_740,N_40,N_191);
nand U741 (N_741,N_177,N_73);
and U742 (N_742,N_16,N_76);
nor U743 (N_743,N_182,N_302);
and U744 (N_744,N_147,N_219);
and U745 (N_745,N_30,N_401);
or U746 (N_746,N_154,N_244);
nand U747 (N_747,N_98,N_93);
nor U748 (N_748,N_216,N_25);
or U749 (N_749,N_156,N_342);
or U750 (N_750,N_272,N_469);
and U751 (N_751,N_122,N_433);
nor U752 (N_752,N_335,N_315);
nor U753 (N_753,N_437,N_147);
nor U754 (N_754,N_407,N_426);
or U755 (N_755,N_242,N_494);
or U756 (N_756,N_70,N_370);
nor U757 (N_757,N_63,N_235);
or U758 (N_758,N_81,N_279);
xnor U759 (N_759,N_229,N_315);
nor U760 (N_760,N_390,N_224);
nor U761 (N_761,N_306,N_10);
nor U762 (N_762,N_145,N_205);
and U763 (N_763,N_323,N_490);
and U764 (N_764,N_221,N_436);
and U765 (N_765,N_344,N_157);
nor U766 (N_766,N_473,N_202);
nand U767 (N_767,N_379,N_264);
xor U768 (N_768,N_131,N_482);
nor U769 (N_769,N_40,N_287);
and U770 (N_770,N_268,N_394);
or U771 (N_771,N_263,N_390);
nand U772 (N_772,N_387,N_40);
nand U773 (N_773,N_353,N_365);
and U774 (N_774,N_495,N_380);
nand U775 (N_775,N_24,N_341);
nor U776 (N_776,N_274,N_187);
nor U777 (N_777,N_175,N_352);
nand U778 (N_778,N_15,N_324);
or U779 (N_779,N_43,N_171);
or U780 (N_780,N_154,N_49);
nand U781 (N_781,N_142,N_274);
and U782 (N_782,N_0,N_416);
and U783 (N_783,N_454,N_234);
nor U784 (N_784,N_201,N_302);
or U785 (N_785,N_139,N_326);
or U786 (N_786,N_327,N_100);
nand U787 (N_787,N_218,N_477);
nor U788 (N_788,N_213,N_427);
and U789 (N_789,N_82,N_174);
nand U790 (N_790,N_279,N_459);
or U791 (N_791,N_468,N_392);
or U792 (N_792,N_267,N_284);
nor U793 (N_793,N_163,N_452);
nor U794 (N_794,N_422,N_218);
nor U795 (N_795,N_130,N_96);
nor U796 (N_796,N_430,N_155);
nand U797 (N_797,N_185,N_491);
nand U798 (N_798,N_438,N_337);
or U799 (N_799,N_363,N_57);
nor U800 (N_800,N_473,N_249);
or U801 (N_801,N_489,N_396);
nand U802 (N_802,N_54,N_13);
nand U803 (N_803,N_310,N_363);
and U804 (N_804,N_444,N_327);
and U805 (N_805,N_33,N_217);
or U806 (N_806,N_167,N_480);
and U807 (N_807,N_62,N_144);
nor U808 (N_808,N_420,N_231);
and U809 (N_809,N_238,N_438);
or U810 (N_810,N_472,N_260);
nand U811 (N_811,N_36,N_113);
and U812 (N_812,N_445,N_361);
or U813 (N_813,N_91,N_147);
xnor U814 (N_814,N_321,N_181);
or U815 (N_815,N_386,N_377);
nand U816 (N_816,N_452,N_301);
nor U817 (N_817,N_388,N_356);
or U818 (N_818,N_117,N_453);
and U819 (N_819,N_15,N_224);
nand U820 (N_820,N_14,N_378);
nor U821 (N_821,N_247,N_75);
nand U822 (N_822,N_58,N_311);
nand U823 (N_823,N_70,N_333);
and U824 (N_824,N_65,N_211);
and U825 (N_825,N_231,N_272);
or U826 (N_826,N_472,N_418);
nand U827 (N_827,N_413,N_244);
nor U828 (N_828,N_386,N_21);
xnor U829 (N_829,N_124,N_187);
or U830 (N_830,N_382,N_91);
or U831 (N_831,N_382,N_31);
nor U832 (N_832,N_82,N_483);
xor U833 (N_833,N_446,N_184);
nand U834 (N_834,N_457,N_199);
nand U835 (N_835,N_69,N_330);
nand U836 (N_836,N_24,N_302);
nor U837 (N_837,N_297,N_481);
or U838 (N_838,N_218,N_487);
nor U839 (N_839,N_390,N_136);
and U840 (N_840,N_350,N_258);
nor U841 (N_841,N_315,N_23);
nor U842 (N_842,N_249,N_280);
or U843 (N_843,N_423,N_15);
and U844 (N_844,N_290,N_196);
or U845 (N_845,N_274,N_94);
nand U846 (N_846,N_91,N_357);
or U847 (N_847,N_255,N_346);
and U848 (N_848,N_465,N_169);
nand U849 (N_849,N_4,N_123);
nor U850 (N_850,N_419,N_263);
and U851 (N_851,N_36,N_344);
and U852 (N_852,N_41,N_401);
and U853 (N_853,N_299,N_439);
xnor U854 (N_854,N_317,N_164);
nand U855 (N_855,N_228,N_377);
or U856 (N_856,N_89,N_167);
or U857 (N_857,N_236,N_20);
or U858 (N_858,N_200,N_111);
or U859 (N_859,N_18,N_330);
and U860 (N_860,N_292,N_115);
nor U861 (N_861,N_478,N_114);
nand U862 (N_862,N_458,N_366);
and U863 (N_863,N_27,N_31);
and U864 (N_864,N_82,N_323);
and U865 (N_865,N_474,N_361);
xnor U866 (N_866,N_411,N_357);
nand U867 (N_867,N_495,N_153);
nand U868 (N_868,N_206,N_297);
nand U869 (N_869,N_85,N_345);
nor U870 (N_870,N_452,N_68);
or U871 (N_871,N_87,N_477);
and U872 (N_872,N_351,N_230);
and U873 (N_873,N_273,N_269);
or U874 (N_874,N_291,N_86);
nand U875 (N_875,N_155,N_237);
and U876 (N_876,N_480,N_387);
or U877 (N_877,N_479,N_12);
nor U878 (N_878,N_246,N_98);
and U879 (N_879,N_209,N_257);
nand U880 (N_880,N_181,N_215);
nor U881 (N_881,N_247,N_367);
nor U882 (N_882,N_78,N_9);
or U883 (N_883,N_409,N_372);
and U884 (N_884,N_115,N_72);
and U885 (N_885,N_314,N_161);
nand U886 (N_886,N_423,N_355);
xnor U887 (N_887,N_449,N_443);
nand U888 (N_888,N_149,N_461);
or U889 (N_889,N_365,N_496);
nor U890 (N_890,N_197,N_279);
nand U891 (N_891,N_323,N_236);
nand U892 (N_892,N_287,N_369);
nand U893 (N_893,N_228,N_485);
nand U894 (N_894,N_115,N_157);
nor U895 (N_895,N_421,N_240);
and U896 (N_896,N_181,N_79);
or U897 (N_897,N_419,N_83);
xor U898 (N_898,N_44,N_189);
nand U899 (N_899,N_221,N_442);
nand U900 (N_900,N_67,N_361);
and U901 (N_901,N_398,N_352);
nand U902 (N_902,N_366,N_39);
or U903 (N_903,N_15,N_321);
and U904 (N_904,N_442,N_393);
xnor U905 (N_905,N_482,N_285);
and U906 (N_906,N_277,N_400);
and U907 (N_907,N_405,N_341);
and U908 (N_908,N_461,N_321);
nand U909 (N_909,N_241,N_106);
and U910 (N_910,N_34,N_204);
nor U911 (N_911,N_419,N_17);
nand U912 (N_912,N_141,N_160);
nand U913 (N_913,N_298,N_331);
nand U914 (N_914,N_337,N_46);
nand U915 (N_915,N_316,N_171);
nor U916 (N_916,N_49,N_372);
and U917 (N_917,N_453,N_184);
and U918 (N_918,N_318,N_406);
and U919 (N_919,N_411,N_247);
nand U920 (N_920,N_89,N_173);
and U921 (N_921,N_28,N_60);
nand U922 (N_922,N_475,N_117);
nor U923 (N_923,N_471,N_87);
or U924 (N_924,N_142,N_101);
and U925 (N_925,N_453,N_91);
nand U926 (N_926,N_405,N_22);
or U927 (N_927,N_79,N_393);
and U928 (N_928,N_474,N_366);
and U929 (N_929,N_138,N_390);
or U930 (N_930,N_73,N_412);
and U931 (N_931,N_400,N_135);
nand U932 (N_932,N_278,N_212);
nor U933 (N_933,N_274,N_361);
and U934 (N_934,N_113,N_383);
and U935 (N_935,N_315,N_384);
nor U936 (N_936,N_18,N_352);
or U937 (N_937,N_459,N_453);
nand U938 (N_938,N_56,N_366);
nor U939 (N_939,N_229,N_278);
and U940 (N_940,N_213,N_280);
or U941 (N_941,N_295,N_59);
and U942 (N_942,N_499,N_116);
or U943 (N_943,N_310,N_260);
nor U944 (N_944,N_450,N_449);
or U945 (N_945,N_267,N_58);
and U946 (N_946,N_185,N_258);
and U947 (N_947,N_488,N_135);
nand U948 (N_948,N_201,N_117);
or U949 (N_949,N_301,N_114);
nand U950 (N_950,N_306,N_167);
nor U951 (N_951,N_243,N_323);
or U952 (N_952,N_23,N_48);
and U953 (N_953,N_15,N_402);
and U954 (N_954,N_382,N_89);
nor U955 (N_955,N_84,N_417);
and U956 (N_956,N_386,N_468);
or U957 (N_957,N_116,N_341);
and U958 (N_958,N_211,N_250);
and U959 (N_959,N_240,N_492);
and U960 (N_960,N_272,N_38);
and U961 (N_961,N_200,N_413);
or U962 (N_962,N_162,N_264);
and U963 (N_963,N_291,N_173);
nor U964 (N_964,N_318,N_288);
nand U965 (N_965,N_358,N_110);
and U966 (N_966,N_467,N_470);
nand U967 (N_967,N_353,N_462);
or U968 (N_968,N_148,N_327);
xor U969 (N_969,N_374,N_269);
nand U970 (N_970,N_133,N_125);
and U971 (N_971,N_84,N_192);
and U972 (N_972,N_107,N_196);
and U973 (N_973,N_471,N_377);
nand U974 (N_974,N_495,N_75);
nor U975 (N_975,N_137,N_465);
and U976 (N_976,N_491,N_305);
nand U977 (N_977,N_499,N_397);
and U978 (N_978,N_167,N_492);
and U979 (N_979,N_162,N_201);
and U980 (N_980,N_272,N_114);
or U981 (N_981,N_491,N_307);
or U982 (N_982,N_326,N_193);
nand U983 (N_983,N_5,N_19);
nand U984 (N_984,N_462,N_145);
and U985 (N_985,N_491,N_12);
nand U986 (N_986,N_454,N_422);
nor U987 (N_987,N_219,N_95);
and U988 (N_988,N_450,N_320);
nand U989 (N_989,N_343,N_496);
nor U990 (N_990,N_3,N_197);
and U991 (N_991,N_112,N_25);
or U992 (N_992,N_263,N_10);
and U993 (N_993,N_171,N_400);
nand U994 (N_994,N_170,N_207);
and U995 (N_995,N_204,N_243);
nor U996 (N_996,N_41,N_400);
and U997 (N_997,N_101,N_222);
and U998 (N_998,N_147,N_494);
nor U999 (N_999,N_176,N_50);
nand U1000 (N_1000,N_849,N_967);
nand U1001 (N_1001,N_891,N_912);
nand U1002 (N_1002,N_673,N_884);
or U1003 (N_1003,N_504,N_826);
nor U1004 (N_1004,N_992,N_877);
or U1005 (N_1005,N_615,N_719);
or U1006 (N_1006,N_677,N_747);
nand U1007 (N_1007,N_553,N_732);
and U1008 (N_1008,N_627,N_995);
and U1009 (N_1009,N_901,N_856);
and U1010 (N_1010,N_923,N_612);
and U1011 (N_1011,N_694,N_675);
nand U1012 (N_1012,N_520,N_532);
nand U1013 (N_1013,N_969,N_723);
or U1014 (N_1014,N_803,N_822);
nand U1015 (N_1015,N_588,N_623);
nand U1016 (N_1016,N_528,N_687);
nor U1017 (N_1017,N_538,N_853);
and U1018 (N_1018,N_578,N_866);
or U1019 (N_1019,N_907,N_679);
nor U1020 (N_1020,N_643,N_961);
or U1021 (N_1021,N_745,N_775);
and U1022 (N_1022,N_962,N_781);
nand U1023 (N_1023,N_734,N_990);
and U1024 (N_1024,N_517,N_640);
or U1025 (N_1025,N_832,N_742);
nor U1026 (N_1026,N_562,N_552);
nand U1027 (N_1027,N_988,N_945);
nor U1028 (N_1028,N_737,N_851);
or U1029 (N_1029,N_610,N_598);
and U1030 (N_1030,N_916,N_974);
and U1031 (N_1031,N_569,N_502);
and U1032 (N_1032,N_978,N_593);
nor U1033 (N_1033,N_872,N_509);
nand U1034 (N_1034,N_536,N_940);
nand U1035 (N_1035,N_513,N_540);
nand U1036 (N_1036,N_772,N_902);
and U1037 (N_1037,N_507,N_931);
and U1038 (N_1038,N_883,N_823);
and U1039 (N_1039,N_767,N_702);
nor U1040 (N_1040,N_638,N_946);
or U1041 (N_1041,N_965,N_881);
nand U1042 (N_1042,N_928,N_736);
nor U1043 (N_1043,N_631,N_587);
and U1044 (N_1044,N_676,N_942);
nor U1045 (N_1045,N_893,N_604);
nor U1046 (N_1046,N_860,N_875);
nor U1047 (N_1047,N_722,N_700);
nand U1048 (N_1048,N_503,N_739);
and U1049 (N_1049,N_956,N_871);
or U1050 (N_1050,N_903,N_614);
or U1051 (N_1051,N_657,N_889);
nand U1052 (N_1052,N_580,N_595);
and U1053 (N_1053,N_611,N_999);
and U1054 (N_1054,N_649,N_852);
and U1055 (N_1055,N_648,N_798);
and U1056 (N_1056,N_548,N_760);
and U1057 (N_1057,N_591,N_617);
nand U1058 (N_1058,N_865,N_996);
and U1059 (N_1059,N_980,N_518);
nand U1060 (N_1060,N_994,N_779);
or U1061 (N_1061,N_761,N_787);
nand U1062 (N_1062,N_692,N_879);
nand U1063 (N_1063,N_824,N_844);
nand U1064 (N_1064,N_574,N_653);
nand U1065 (N_1065,N_905,N_756);
or U1066 (N_1066,N_589,N_966);
and U1067 (N_1067,N_914,N_937);
and U1068 (N_1068,N_973,N_867);
or U1069 (N_1069,N_519,N_650);
nor U1070 (N_1070,N_782,N_510);
and U1071 (N_1071,N_656,N_701);
nor U1072 (N_1072,N_618,N_819);
nand U1073 (N_1073,N_897,N_957);
and U1074 (N_1074,N_987,N_663);
nand U1075 (N_1075,N_689,N_601);
nand U1076 (N_1076,N_876,N_955);
nand U1077 (N_1077,N_514,N_697);
and U1078 (N_1078,N_930,N_830);
nor U1079 (N_1079,N_555,N_726);
nor U1080 (N_1080,N_911,N_765);
or U1081 (N_1081,N_546,N_972);
or U1082 (N_1082,N_695,N_783);
nand U1083 (N_1083,N_516,N_915);
nand U1084 (N_1084,N_743,N_843);
nand U1085 (N_1085,N_597,N_926);
and U1086 (N_1086,N_838,N_810);
and U1087 (N_1087,N_836,N_599);
or U1088 (N_1088,N_848,N_573);
or U1089 (N_1089,N_568,N_837);
or U1090 (N_1090,N_885,N_887);
and U1091 (N_1091,N_585,N_768);
and U1092 (N_1092,N_949,N_952);
nand U1093 (N_1093,N_935,N_845);
nor U1094 (N_1094,N_661,N_964);
and U1095 (N_1095,N_556,N_682);
and U1096 (N_1096,N_985,N_954);
and U1097 (N_1097,N_533,N_602);
nand U1098 (N_1098,N_850,N_629);
and U1099 (N_1099,N_936,N_549);
nand U1100 (N_1100,N_842,N_963);
nand U1101 (N_1101,N_806,N_545);
or U1102 (N_1102,N_725,N_672);
nand U1103 (N_1103,N_791,N_804);
or U1104 (N_1104,N_763,N_869);
or U1105 (N_1105,N_635,N_951);
nand U1106 (N_1106,N_691,N_724);
nor U1107 (N_1107,N_859,N_619);
nor U1108 (N_1108,N_641,N_799);
nand U1109 (N_1109,N_829,N_809);
or U1110 (N_1110,N_727,N_854);
and U1111 (N_1111,N_714,N_862);
and U1112 (N_1112,N_645,N_764);
or U1113 (N_1113,N_939,N_835);
xor U1114 (N_1114,N_758,N_913);
nand U1115 (N_1115,N_655,N_784);
nand U1116 (N_1116,N_906,N_831);
or U1117 (N_1117,N_728,N_792);
xor U1118 (N_1118,N_515,N_566);
and U1119 (N_1119,N_886,N_741);
nor U1120 (N_1120,N_626,N_530);
or U1121 (N_1121,N_584,N_525);
nor U1122 (N_1122,N_733,N_633);
or U1123 (N_1123,N_878,N_710);
and U1124 (N_1124,N_704,N_534);
xor U1125 (N_1125,N_646,N_561);
nand U1126 (N_1126,N_984,N_802);
nor U1127 (N_1127,N_526,N_828);
or U1128 (N_1128,N_609,N_505);
and U1129 (N_1129,N_894,N_947);
or U1130 (N_1130,N_993,N_753);
or U1131 (N_1131,N_581,N_715);
or U1132 (N_1132,N_681,N_698);
and U1133 (N_1133,N_735,N_958);
xnor U1134 (N_1134,N_696,N_861);
nand U1135 (N_1135,N_751,N_523);
or U1136 (N_1136,N_795,N_582);
and U1137 (N_1137,N_636,N_716);
nor U1138 (N_1138,N_757,N_818);
and U1139 (N_1139,N_680,N_814);
nand U1140 (N_1140,N_943,N_571);
nand U1141 (N_1141,N_748,N_991);
or U1142 (N_1142,N_986,N_846);
or U1143 (N_1143,N_801,N_896);
or U1144 (N_1144,N_977,N_731);
and U1145 (N_1145,N_855,N_586);
nor U1146 (N_1146,N_554,N_535);
and U1147 (N_1147,N_909,N_821);
nor U1148 (N_1148,N_620,N_521);
nor U1149 (N_1149,N_808,N_729);
nand U1150 (N_1150,N_605,N_770);
or U1151 (N_1151,N_576,N_669);
nand U1152 (N_1152,N_600,N_684);
nor U1153 (N_1153,N_630,N_531);
nor U1154 (N_1154,N_975,N_671);
and U1155 (N_1155,N_637,N_550);
nand U1156 (N_1156,N_709,N_793);
and U1157 (N_1157,N_558,N_982);
or U1158 (N_1158,N_929,N_820);
or U1159 (N_1159,N_752,N_922);
xor U1160 (N_1160,N_537,N_740);
or U1161 (N_1161,N_738,N_932);
nor U1162 (N_1162,N_847,N_693);
nor U1163 (N_1163,N_890,N_707);
and U1164 (N_1164,N_579,N_577);
nand U1165 (N_1165,N_812,N_685);
nand U1166 (N_1166,N_639,N_864);
or U1167 (N_1167,N_543,N_624);
nand U1168 (N_1168,N_665,N_927);
and U1169 (N_1169,N_933,N_938);
nor U1170 (N_1170,N_570,N_750);
nor U1171 (N_1171,N_690,N_882);
nor U1172 (N_1172,N_572,N_892);
nor U1173 (N_1173,N_688,N_796);
xor U1174 (N_1174,N_904,N_529);
and U1175 (N_1175,N_919,N_563);
or U1176 (N_1176,N_934,N_950);
nand U1177 (N_1177,N_621,N_730);
nor U1178 (N_1178,N_632,N_785);
nand U1179 (N_1179,N_642,N_777);
nor U1180 (N_1180,N_979,N_788);
nor U1181 (N_1181,N_834,N_717);
and U1182 (N_1182,N_652,N_590);
nand U1183 (N_1183,N_551,N_983);
nand U1184 (N_1184,N_908,N_759);
or U1185 (N_1185,N_564,N_773);
xnor U1186 (N_1186,N_989,N_501);
nor U1187 (N_1187,N_721,N_868);
nand U1188 (N_1188,N_805,N_705);
nand U1189 (N_1189,N_976,N_910);
and U1190 (N_1190,N_666,N_664);
nand U1191 (N_1191,N_713,N_613);
nand U1192 (N_1192,N_662,N_522);
nand U1193 (N_1193,N_895,N_997);
and U1194 (N_1194,N_557,N_873);
nor U1195 (N_1195,N_888,N_660);
nand U1196 (N_1196,N_651,N_658);
nand U1197 (N_1197,N_678,N_944);
and U1198 (N_1198,N_527,N_815);
nor U1199 (N_1199,N_790,N_771);
xor U1200 (N_1200,N_718,N_863);
nand U1201 (N_1201,N_924,N_744);
or U1202 (N_1202,N_817,N_769);
nand U1203 (N_1203,N_712,N_647);
or U1204 (N_1204,N_825,N_711);
and U1205 (N_1205,N_827,N_789);
xor U1206 (N_1206,N_925,N_880);
nor U1207 (N_1207,N_606,N_559);
nand U1208 (N_1208,N_634,N_720);
or U1209 (N_1209,N_800,N_583);
nor U1210 (N_1210,N_592,N_616);
nor U1211 (N_1211,N_544,N_508);
nand U1212 (N_1212,N_674,N_998);
and U1213 (N_1213,N_512,N_628);
or U1214 (N_1214,N_500,N_607);
nand U1215 (N_1215,N_667,N_668);
nand U1216 (N_1216,N_541,N_654);
and U1217 (N_1217,N_766,N_778);
nor U1218 (N_1218,N_959,N_813);
nor U1219 (N_1219,N_703,N_560);
nand U1220 (N_1220,N_857,N_776);
nand U1221 (N_1221,N_603,N_575);
and U1222 (N_1222,N_708,N_797);
nand U1223 (N_1223,N_960,N_941);
nand U1224 (N_1224,N_858,N_625);
or U1225 (N_1225,N_594,N_547);
nand U1226 (N_1226,N_567,N_921);
and U1227 (N_1227,N_870,N_981);
and U1228 (N_1228,N_746,N_699);
nand U1229 (N_1229,N_899,N_706);
nand U1230 (N_1230,N_898,N_511);
nand U1231 (N_1231,N_542,N_659);
xor U1232 (N_1232,N_953,N_971);
nand U1233 (N_1233,N_608,N_644);
nor U1234 (N_1234,N_755,N_524);
and U1235 (N_1235,N_683,N_774);
nor U1236 (N_1236,N_686,N_565);
nor U1237 (N_1237,N_816,N_948);
and U1238 (N_1238,N_670,N_811);
nor U1239 (N_1239,N_762,N_506);
xnor U1240 (N_1240,N_807,N_841);
or U1241 (N_1241,N_968,N_794);
nand U1242 (N_1242,N_917,N_970);
and U1243 (N_1243,N_918,N_596);
and U1244 (N_1244,N_840,N_874);
nor U1245 (N_1245,N_539,N_786);
or U1246 (N_1246,N_839,N_780);
or U1247 (N_1247,N_622,N_900);
nor U1248 (N_1248,N_833,N_920);
and U1249 (N_1249,N_749,N_754);
or U1250 (N_1250,N_723,N_682);
nand U1251 (N_1251,N_766,N_536);
nand U1252 (N_1252,N_583,N_762);
or U1253 (N_1253,N_569,N_973);
or U1254 (N_1254,N_752,N_725);
and U1255 (N_1255,N_787,N_875);
nand U1256 (N_1256,N_740,N_969);
or U1257 (N_1257,N_808,N_919);
nand U1258 (N_1258,N_520,N_512);
or U1259 (N_1259,N_591,N_527);
nand U1260 (N_1260,N_752,N_562);
or U1261 (N_1261,N_551,N_783);
nor U1262 (N_1262,N_708,N_813);
and U1263 (N_1263,N_949,N_983);
or U1264 (N_1264,N_904,N_727);
or U1265 (N_1265,N_896,N_616);
or U1266 (N_1266,N_811,N_926);
nor U1267 (N_1267,N_888,N_934);
or U1268 (N_1268,N_720,N_970);
xnor U1269 (N_1269,N_680,N_641);
nand U1270 (N_1270,N_975,N_839);
or U1271 (N_1271,N_713,N_892);
xnor U1272 (N_1272,N_935,N_503);
nor U1273 (N_1273,N_921,N_726);
and U1274 (N_1274,N_614,N_734);
or U1275 (N_1275,N_545,N_669);
nand U1276 (N_1276,N_740,N_887);
xnor U1277 (N_1277,N_616,N_859);
nor U1278 (N_1278,N_934,N_608);
and U1279 (N_1279,N_888,N_576);
nand U1280 (N_1280,N_623,N_634);
nor U1281 (N_1281,N_562,N_988);
nand U1282 (N_1282,N_923,N_561);
nor U1283 (N_1283,N_721,N_548);
nand U1284 (N_1284,N_774,N_891);
and U1285 (N_1285,N_997,N_950);
nand U1286 (N_1286,N_891,N_926);
xnor U1287 (N_1287,N_561,N_913);
and U1288 (N_1288,N_544,N_659);
and U1289 (N_1289,N_664,N_682);
nand U1290 (N_1290,N_628,N_665);
nor U1291 (N_1291,N_603,N_553);
nand U1292 (N_1292,N_990,N_980);
nand U1293 (N_1293,N_823,N_538);
and U1294 (N_1294,N_945,N_934);
nor U1295 (N_1295,N_753,N_800);
and U1296 (N_1296,N_839,N_996);
nand U1297 (N_1297,N_968,N_797);
and U1298 (N_1298,N_753,N_734);
nor U1299 (N_1299,N_988,N_918);
nor U1300 (N_1300,N_882,N_587);
or U1301 (N_1301,N_632,N_856);
nand U1302 (N_1302,N_704,N_724);
and U1303 (N_1303,N_629,N_977);
and U1304 (N_1304,N_808,N_598);
nand U1305 (N_1305,N_690,N_957);
or U1306 (N_1306,N_788,N_676);
and U1307 (N_1307,N_803,N_799);
xor U1308 (N_1308,N_860,N_539);
nand U1309 (N_1309,N_863,N_942);
and U1310 (N_1310,N_765,N_632);
or U1311 (N_1311,N_804,N_874);
nor U1312 (N_1312,N_727,N_715);
nand U1313 (N_1313,N_896,N_515);
or U1314 (N_1314,N_606,N_940);
nor U1315 (N_1315,N_656,N_714);
and U1316 (N_1316,N_555,N_528);
and U1317 (N_1317,N_715,N_962);
or U1318 (N_1318,N_836,N_759);
nand U1319 (N_1319,N_602,N_974);
nand U1320 (N_1320,N_977,N_514);
and U1321 (N_1321,N_576,N_909);
nor U1322 (N_1322,N_930,N_711);
nand U1323 (N_1323,N_530,N_882);
or U1324 (N_1324,N_844,N_998);
and U1325 (N_1325,N_758,N_571);
nor U1326 (N_1326,N_938,N_661);
or U1327 (N_1327,N_895,N_970);
nand U1328 (N_1328,N_949,N_750);
nor U1329 (N_1329,N_839,N_695);
or U1330 (N_1330,N_992,N_888);
or U1331 (N_1331,N_723,N_566);
nand U1332 (N_1332,N_765,N_501);
or U1333 (N_1333,N_518,N_834);
or U1334 (N_1334,N_935,N_724);
nor U1335 (N_1335,N_669,N_717);
nand U1336 (N_1336,N_856,N_935);
or U1337 (N_1337,N_672,N_665);
nand U1338 (N_1338,N_576,N_611);
nor U1339 (N_1339,N_998,N_626);
or U1340 (N_1340,N_666,N_786);
nand U1341 (N_1341,N_835,N_975);
and U1342 (N_1342,N_547,N_728);
xnor U1343 (N_1343,N_780,N_571);
or U1344 (N_1344,N_524,N_986);
nand U1345 (N_1345,N_540,N_671);
nor U1346 (N_1346,N_630,N_922);
nand U1347 (N_1347,N_920,N_952);
nor U1348 (N_1348,N_831,N_738);
and U1349 (N_1349,N_525,N_590);
nor U1350 (N_1350,N_967,N_638);
and U1351 (N_1351,N_844,N_554);
nor U1352 (N_1352,N_930,N_506);
nor U1353 (N_1353,N_783,N_756);
nand U1354 (N_1354,N_533,N_592);
and U1355 (N_1355,N_960,N_991);
nor U1356 (N_1356,N_677,N_922);
nand U1357 (N_1357,N_814,N_601);
nand U1358 (N_1358,N_756,N_596);
nor U1359 (N_1359,N_777,N_725);
nor U1360 (N_1360,N_885,N_673);
nand U1361 (N_1361,N_765,N_693);
and U1362 (N_1362,N_546,N_657);
nand U1363 (N_1363,N_567,N_551);
nor U1364 (N_1364,N_618,N_670);
and U1365 (N_1365,N_730,N_890);
or U1366 (N_1366,N_621,N_884);
and U1367 (N_1367,N_966,N_761);
or U1368 (N_1368,N_796,N_604);
nand U1369 (N_1369,N_784,N_727);
or U1370 (N_1370,N_618,N_757);
or U1371 (N_1371,N_642,N_855);
nand U1372 (N_1372,N_706,N_503);
and U1373 (N_1373,N_796,N_939);
nand U1374 (N_1374,N_806,N_840);
and U1375 (N_1375,N_650,N_891);
and U1376 (N_1376,N_738,N_844);
and U1377 (N_1377,N_549,N_800);
nor U1378 (N_1378,N_732,N_736);
nand U1379 (N_1379,N_928,N_659);
nor U1380 (N_1380,N_960,N_775);
and U1381 (N_1381,N_882,N_971);
nand U1382 (N_1382,N_679,N_982);
or U1383 (N_1383,N_862,N_513);
nand U1384 (N_1384,N_840,N_633);
or U1385 (N_1385,N_824,N_806);
nand U1386 (N_1386,N_588,N_620);
nand U1387 (N_1387,N_976,N_543);
or U1388 (N_1388,N_740,N_856);
nand U1389 (N_1389,N_729,N_509);
nand U1390 (N_1390,N_934,N_600);
or U1391 (N_1391,N_580,N_952);
nor U1392 (N_1392,N_700,N_883);
or U1393 (N_1393,N_537,N_706);
xor U1394 (N_1394,N_744,N_959);
nor U1395 (N_1395,N_854,N_932);
nor U1396 (N_1396,N_837,N_554);
nor U1397 (N_1397,N_971,N_931);
nand U1398 (N_1398,N_698,N_506);
nand U1399 (N_1399,N_952,N_953);
or U1400 (N_1400,N_764,N_805);
nand U1401 (N_1401,N_916,N_767);
and U1402 (N_1402,N_796,N_852);
nand U1403 (N_1403,N_790,N_641);
or U1404 (N_1404,N_519,N_793);
or U1405 (N_1405,N_799,N_544);
and U1406 (N_1406,N_922,N_708);
and U1407 (N_1407,N_765,N_609);
and U1408 (N_1408,N_573,N_718);
or U1409 (N_1409,N_718,N_794);
nor U1410 (N_1410,N_671,N_939);
and U1411 (N_1411,N_502,N_520);
or U1412 (N_1412,N_500,N_524);
nand U1413 (N_1413,N_610,N_956);
and U1414 (N_1414,N_958,N_558);
nor U1415 (N_1415,N_896,N_645);
nand U1416 (N_1416,N_751,N_872);
nand U1417 (N_1417,N_995,N_928);
or U1418 (N_1418,N_675,N_945);
nor U1419 (N_1419,N_635,N_886);
nor U1420 (N_1420,N_634,N_925);
and U1421 (N_1421,N_957,N_558);
or U1422 (N_1422,N_577,N_606);
nor U1423 (N_1423,N_985,N_967);
and U1424 (N_1424,N_992,N_670);
nand U1425 (N_1425,N_705,N_614);
or U1426 (N_1426,N_598,N_717);
and U1427 (N_1427,N_642,N_709);
or U1428 (N_1428,N_687,N_526);
or U1429 (N_1429,N_790,N_909);
and U1430 (N_1430,N_977,N_522);
or U1431 (N_1431,N_525,N_683);
nand U1432 (N_1432,N_757,N_603);
nor U1433 (N_1433,N_586,N_947);
or U1434 (N_1434,N_821,N_813);
and U1435 (N_1435,N_914,N_589);
nand U1436 (N_1436,N_717,N_589);
nand U1437 (N_1437,N_713,N_757);
nor U1438 (N_1438,N_847,N_550);
nor U1439 (N_1439,N_624,N_581);
nand U1440 (N_1440,N_608,N_513);
nand U1441 (N_1441,N_603,N_584);
nand U1442 (N_1442,N_675,N_960);
and U1443 (N_1443,N_865,N_935);
or U1444 (N_1444,N_762,N_897);
and U1445 (N_1445,N_931,N_562);
nand U1446 (N_1446,N_697,N_635);
nor U1447 (N_1447,N_767,N_909);
nand U1448 (N_1448,N_531,N_609);
nor U1449 (N_1449,N_969,N_530);
and U1450 (N_1450,N_638,N_741);
or U1451 (N_1451,N_707,N_979);
or U1452 (N_1452,N_646,N_921);
nand U1453 (N_1453,N_997,N_887);
and U1454 (N_1454,N_716,N_912);
or U1455 (N_1455,N_835,N_825);
nand U1456 (N_1456,N_667,N_736);
or U1457 (N_1457,N_947,N_787);
and U1458 (N_1458,N_881,N_943);
and U1459 (N_1459,N_783,N_776);
and U1460 (N_1460,N_544,N_916);
or U1461 (N_1461,N_829,N_954);
and U1462 (N_1462,N_810,N_653);
nor U1463 (N_1463,N_911,N_743);
nand U1464 (N_1464,N_925,N_730);
or U1465 (N_1465,N_843,N_600);
nor U1466 (N_1466,N_778,N_756);
nor U1467 (N_1467,N_713,N_994);
or U1468 (N_1468,N_600,N_962);
and U1469 (N_1469,N_534,N_583);
nand U1470 (N_1470,N_887,N_761);
or U1471 (N_1471,N_626,N_872);
and U1472 (N_1472,N_773,N_779);
nor U1473 (N_1473,N_657,N_744);
and U1474 (N_1474,N_845,N_744);
nor U1475 (N_1475,N_619,N_765);
or U1476 (N_1476,N_584,N_595);
and U1477 (N_1477,N_582,N_881);
nand U1478 (N_1478,N_555,N_527);
and U1479 (N_1479,N_594,N_597);
and U1480 (N_1480,N_885,N_897);
nor U1481 (N_1481,N_789,N_842);
or U1482 (N_1482,N_987,N_697);
or U1483 (N_1483,N_830,N_988);
nor U1484 (N_1484,N_581,N_951);
and U1485 (N_1485,N_576,N_799);
or U1486 (N_1486,N_937,N_930);
nand U1487 (N_1487,N_631,N_694);
nand U1488 (N_1488,N_980,N_970);
or U1489 (N_1489,N_939,N_624);
nor U1490 (N_1490,N_871,N_786);
and U1491 (N_1491,N_952,N_564);
and U1492 (N_1492,N_802,N_769);
and U1493 (N_1493,N_693,N_745);
and U1494 (N_1494,N_724,N_869);
or U1495 (N_1495,N_564,N_552);
nor U1496 (N_1496,N_779,N_807);
and U1497 (N_1497,N_772,N_507);
and U1498 (N_1498,N_778,N_564);
nor U1499 (N_1499,N_779,N_502);
or U1500 (N_1500,N_1368,N_1154);
and U1501 (N_1501,N_1150,N_1067);
or U1502 (N_1502,N_1495,N_1032);
or U1503 (N_1503,N_1078,N_1369);
nand U1504 (N_1504,N_1351,N_1395);
nand U1505 (N_1505,N_1217,N_1004);
nor U1506 (N_1506,N_1125,N_1255);
and U1507 (N_1507,N_1337,N_1149);
nor U1508 (N_1508,N_1047,N_1325);
nand U1509 (N_1509,N_1073,N_1466);
or U1510 (N_1510,N_1106,N_1181);
or U1511 (N_1511,N_1431,N_1418);
nand U1512 (N_1512,N_1044,N_1222);
nor U1513 (N_1513,N_1002,N_1173);
or U1514 (N_1514,N_1463,N_1184);
nand U1515 (N_1515,N_1072,N_1135);
and U1516 (N_1516,N_1287,N_1063);
or U1517 (N_1517,N_1052,N_1464);
nand U1518 (N_1518,N_1429,N_1486);
and U1519 (N_1519,N_1472,N_1126);
xor U1520 (N_1520,N_1039,N_1269);
or U1521 (N_1521,N_1299,N_1153);
or U1522 (N_1522,N_1417,N_1275);
nand U1523 (N_1523,N_1372,N_1103);
and U1524 (N_1524,N_1005,N_1192);
and U1525 (N_1525,N_1271,N_1068);
and U1526 (N_1526,N_1300,N_1127);
nor U1527 (N_1527,N_1454,N_1168);
or U1528 (N_1528,N_1460,N_1379);
and U1529 (N_1529,N_1499,N_1478);
and U1530 (N_1530,N_1470,N_1292);
nand U1531 (N_1531,N_1183,N_1388);
and U1532 (N_1532,N_1290,N_1357);
and U1533 (N_1533,N_1145,N_1137);
nor U1534 (N_1534,N_1489,N_1331);
nor U1535 (N_1535,N_1237,N_1266);
and U1536 (N_1536,N_1311,N_1169);
nand U1537 (N_1537,N_1254,N_1383);
or U1538 (N_1538,N_1128,N_1438);
nor U1539 (N_1539,N_1256,N_1323);
nand U1540 (N_1540,N_1029,N_1170);
nor U1541 (N_1541,N_1278,N_1406);
nand U1542 (N_1542,N_1229,N_1028);
or U1543 (N_1543,N_1310,N_1131);
or U1544 (N_1544,N_1442,N_1057);
and U1545 (N_1545,N_1398,N_1353);
and U1546 (N_1546,N_1015,N_1240);
nand U1547 (N_1547,N_1257,N_1187);
nand U1548 (N_1548,N_1307,N_1496);
and U1549 (N_1549,N_1286,N_1411);
nand U1550 (N_1550,N_1247,N_1262);
or U1551 (N_1551,N_1041,N_1136);
and U1552 (N_1552,N_1021,N_1394);
nor U1553 (N_1553,N_1043,N_1324);
and U1554 (N_1554,N_1318,N_1061);
nor U1555 (N_1555,N_1077,N_1194);
or U1556 (N_1556,N_1322,N_1373);
nor U1557 (N_1557,N_1098,N_1200);
or U1558 (N_1558,N_1280,N_1296);
or U1559 (N_1559,N_1444,N_1282);
nand U1560 (N_1560,N_1109,N_1025);
nand U1561 (N_1561,N_1377,N_1189);
xnor U1562 (N_1562,N_1349,N_1000);
and U1563 (N_1563,N_1160,N_1402);
and U1564 (N_1564,N_1422,N_1102);
or U1565 (N_1565,N_1301,N_1390);
nor U1566 (N_1566,N_1405,N_1093);
or U1567 (N_1567,N_1066,N_1343);
nor U1568 (N_1568,N_1295,N_1273);
or U1569 (N_1569,N_1451,N_1453);
nand U1570 (N_1570,N_1082,N_1233);
or U1571 (N_1571,N_1224,N_1013);
nand U1572 (N_1572,N_1235,N_1308);
or U1573 (N_1573,N_1027,N_1081);
or U1574 (N_1574,N_1441,N_1058);
nor U1575 (N_1575,N_1230,N_1070);
and U1576 (N_1576,N_1448,N_1342);
or U1577 (N_1577,N_1420,N_1205);
or U1578 (N_1578,N_1366,N_1344);
nor U1579 (N_1579,N_1085,N_1414);
and U1580 (N_1580,N_1320,N_1216);
nor U1581 (N_1581,N_1111,N_1167);
nand U1582 (N_1582,N_1370,N_1449);
or U1583 (N_1583,N_1242,N_1246);
xor U1584 (N_1584,N_1363,N_1151);
or U1585 (N_1585,N_1272,N_1143);
nor U1586 (N_1586,N_1392,N_1202);
and U1587 (N_1587,N_1226,N_1010);
nand U1588 (N_1588,N_1421,N_1424);
or U1589 (N_1589,N_1380,N_1386);
or U1590 (N_1590,N_1313,N_1371);
nor U1591 (N_1591,N_1447,N_1129);
and U1592 (N_1592,N_1274,N_1465);
nor U1593 (N_1593,N_1139,N_1018);
nand U1594 (N_1594,N_1014,N_1118);
and U1595 (N_1595,N_1212,N_1482);
nor U1596 (N_1596,N_1034,N_1211);
xnor U1597 (N_1597,N_1091,N_1361);
nor U1598 (N_1598,N_1455,N_1413);
and U1599 (N_1599,N_1459,N_1297);
nor U1600 (N_1600,N_1471,N_1396);
nand U1601 (N_1601,N_1206,N_1060);
nor U1602 (N_1602,N_1488,N_1201);
nor U1603 (N_1603,N_1355,N_1326);
nand U1604 (N_1604,N_1031,N_1279);
and U1605 (N_1605,N_1214,N_1384);
nor U1606 (N_1606,N_1439,N_1327);
or U1607 (N_1607,N_1283,N_1458);
and U1608 (N_1608,N_1003,N_1095);
nand U1609 (N_1609,N_1116,N_1191);
and U1610 (N_1610,N_1046,N_1195);
nand U1611 (N_1611,N_1354,N_1223);
nor U1612 (N_1612,N_1490,N_1140);
or U1613 (N_1613,N_1409,N_1336);
and U1614 (N_1614,N_1219,N_1258);
nand U1615 (N_1615,N_1239,N_1190);
or U1616 (N_1616,N_1281,N_1412);
or U1617 (N_1617,N_1374,N_1023);
nor U1618 (N_1618,N_1410,N_1026);
or U1619 (N_1619,N_1265,N_1450);
nor U1620 (N_1620,N_1248,N_1427);
nand U1621 (N_1621,N_1251,N_1376);
and U1622 (N_1622,N_1339,N_1425);
nand U1623 (N_1623,N_1113,N_1285);
and U1624 (N_1624,N_1393,N_1443);
nor U1625 (N_1625,N_1075,N_1227);
nor U1626 (N_1626,N_1110,N_1074);
or U1627 (N_1627,N_1294,N_1302);
or U1628 (N_1628,N_1094,N_1011);
nand U1629 (N_1629,N_1435,N_1172);
and U1630 (N_1630,N_1048,N_1391);
or U1631 (N_1631,N_1008,N_1457);
nor U1632 (N_1632,N_1468,N_1155);
nand U1633 (N_1633,N_1232,N_1213);
and U1634 (N_1634,N_1261,N_1434);
and U1635 (N_1635,N_1341,N_1007);
and U1636 (N_1636,N_1188,N_1130);
nand U1637 (N_1637,N_1346,N_1364);
and U1638 (N_1638,N_1108,N_1433);
and U1639 (N_1639,N_1186,N_1267);
nand U1640 (N_1640,N_1303,N_1001);
nand U1641 (N_1641,N_1174,N_1132);
and U1642 (N_1642,N_1315,N_1062);
or U1643 (N_1643,N_1166,N_1289);
or U1644 (N_1644,N_1356,N_1087);
nor U1645 (N_1645,N_1185,N_1494);
nor U1646 (N_1646,N_1220,N_1157);
and U1647 (N_1647,N_1399,N_1179);
nand U1648 (N_1648,N_1334,N_1092);
nand U1649 (N_1649,N_1430,N_1104);
and U1650 (N_1650,N_1119,N_1141);
nand U1651 (N_1651,N_1484,N_1309);
and U1652 (N_1652,N_1176,N_1350);
nand U1653 (N_1653,N_1375,N_1475);
and U1654 (N_1654,N_1483,N_1117);
or U1655 (N_1655,N_1319,N_1249);
and U1656 (N_1656,N_1403,N_1099);
or U1657 (N_1657,N_1020,N_1012);
and U1658 (N_1658,N_1493,N_1264);
and U1659 (N_1659,N_1407,N_1291);
nand U1660 (N_1660,N_1316,N_1175);
nor U1661 (N_1661,N_1298,N_1097);
and U1662 (N_1662,N_1071,N_1133);
or U1663 (N_1663,N_1122,N_1218);
and U1664 (N_1664,N_1045,N_1147);
or U1665 (N_1665,N_1462,N_1144);
and U1666 (N_1666,N_1263,N_1481);
or U1667 (N_1667,N_1452,N_1332);
nor U1668 (N_1668,N_1204,N_1193);
nor U1669 (N_1669,N_1474,N_1378);
and U1670 (N_1670,N_1114,N_1345);
nand U1671 (N_1671,N_1006,N_1069);
or U1672 (N_1672,N_1284,N_1050);
or U1673 (N_1673,N_1096,N_1142);
or U1674 (N_1674,N_1423,N_1146);
nand U1675 (N_1675,N_1059,N_1196);
nor U1676 (N_1676,N_1024,N_1162);
and U1677 (N_1677,N_1033,N_1253);
nor U1678 (N_1678,N_1415,N_1365);
or U1679 (N_1679,N_1340,N_1105);
nand U1680 (N_1680,N_1042,N_1035);
nand U1681 (N_1681,N_1270,N_1260);
nor U1682 (N_1682,N_1030,N_1446);
and U1683 (N_1683,N_1065,N_1054);
nor U1684 (N_1684,N_1440,N_1485);
or U1685 (N_1685,N_1487,N_1243);
and U1686 (N_1686,N_1416,N_1362);
and U1687 (N_1687,N_1497,N_1208);
nand U1688 (N_1688,N_1215,N_1330);
or U1689 (N_1689,N_1277,N_1123);
nor U1690 (N_1690,N_1231,N_1498);
nand U1691 (N_1691,N_1360,N_1088);
and U1692 (N_1692,N_1080,N_1009);
nor U1693 (N_1693,N_1469,N_1178);
or U1694 (N_1694,N_1120,N_1049);
and U1695 (N_1695,N_1428,N_1252);
and U1696 (N_1696,N_1401,N_1225);
nor U1697 (N_1697,N_1038,N_1473);
nand U1698 (N_1698,N_1036,N_1382);
and U1699 (N_1699,N_1304,N_1437);
and U1700 (N_1700,N_1419,N_1461);
nor U1701 (N_1701,N_1124,N_1335);
nand U1702 (N_1702,N_1305,N_1138);
nor U1703 (N_1703,N_1228,N_1051);
nand U1704 (N_1704,N_1134,N_1017);
nor U1705 (N_1705,N_1101,N_1019);
nand U1706 (N_1706,N_1210,N_1359);
or U1707 (N_1707,N_1100,N_1209);
and U1708 (N_1708,N_1480,N_1159);
and U1709 (N_1709,N_1387,N_1241);
nor U1710 (N_1710,N_1329,N_1436);
nand U1711 (N_1711,N_1321,N_1040);
or U1712 (N_1712,N_1400,N_1306);
nand U1713 (N_1713,N_1314,N_1389);
or U1714 (N_1714,N_1083,N_1076);
nand U1715 (N_1715,N_1221,N_1056);
nand U1716 (N_1716,N_1317,N_1203);
or U1717 (N_1717,N_1158,N_1426);
nor U1718 (N_1718,N_1171,N_1333);
nor U1719 (N_1719,N_1408,N_1352);
xnor U1720 (N_1720,N_1328,N_1112);
nor U1721 (N_1721,N_1385,N_1207);
and U1722 (N_1722,N_1347,N_1338);
nor U1723 (N_1723,N_1084,N_1404);
or U1724 (N_1724,N_1152,N_1492);
or U1725 (N_1725,N_1182,N_1053);
nand U1726 (N_1726,N_1381,N_1467);
nor U1727 (N_1727,N_1238,N_1445);
nand U1728 (N_1728,N_1016,N_1163);
nor U1729 (N_1729,N_1358,N_1037);
nand U1730 (N_1730,N_1165,N_1090);
nand U1731 (N_1731,N_1161,N_1397);
nand U1732 (N_1732,N_1177,N_1432);
nand U1733 (N_1733,N_1479,N_1055);
nor U1734 (N_1734,N_1086,N_1234);
or U1735 (N_1735,N_1236,N_1276);
or U1736 (N_1736,N_1198,N_1022);
nand U1737 (N_1737,N_1268,N_1079);
nand U1738 (N_1738,N_1064,N_1491);
nor U1739 (N_1739,N_1259,N_1156);
or U1740 (N_1740,N_1456,N_1367);
and U1741 (N_1741,N_1288,N_1476);
and U1742 (N_1742,N_1164,N_1244);
or U1743 (N_1743,N_1245,N_1115);
or U1744 (N_1744,N_1089,N_1148);
nor U1745 (N_1745,N_1199,N_1312);
or U1746 (N_1746,N_1121,N_1293);
and U1747 (N_1747,N_1348,N_1107);
nand U1748 (N_1748,N_1180,N_1197);
and U1749 (N_1749,N_1250,N_1477);
nand U1750 (N_1750,N_1315,N_1130);
nand U1751 (N_1751,N_1318,N_1091);
nand U1752 (N_1752,N_1315,N_1414);
nand U1753 (N_1753,N_1081,N_1348);
nand U1754 (N_1754,N_1087,N_1256);
nor U1755 (N_1755,N_1257,N_1045);
nor U1756 (N_1756,N_1140,N_1333);
or U1757 (N_1757,N_1038,N_1045);
nor U1758 (N_1758,N_1385,N_1418);
or U1759 (N_1759,N_1129,N_1367);
nor U1760 (N_1760,N_1388,N_1150);
or U1761 (N_1761,N_1109,N_1231);
nor U1762 (N_1762,N_1088,N_1493);
and U1763 (N_1763,N_1033,N_1367);
and U1764 (N_1764,N_1218,N_1222);
nor U1765 (N_1765,N_1371,N_1413);
nand U1766 (N_1766,N_1363,N_1041);
and U1767 (N_1767,N_1442,N_1022);
and U1768 (N_1768,N_1444,N_1189);
nor U1769 (N_1769,N_1083,N_1233);
nand U1770 (N_1770,N_1279,N_1420);
and U1771 (N_1771,N_1060,N_1353);
and U1772 (N_1772,N_1341,N_1406);
and U1773 (N_1773,N_1393,N_1354);
nor U1774 (N_1774,N_1365,N_1058);
and U1775 (N_1775,N_1303,N_1283);
nor U1776 (N_1776,N_1095,N_1348);
nand U1777 (N_1777,N_1389,N_1395);
nand U1778 (N_1778,N_1457,N_1204);
nor U1779 (N_1779,N_1157,N_1335);
nand U1780 (N_1780,N_1267,N_1428);
nor U1781 (N_1781,N_1479,N_1334);
or U1782 (N_1782,N_1489,N_1079);
nor U1783 (N_1783,N_1292,N_1257);
nor U1784 (N_1784,N_1477,N_1174);
or U1785 (N_1785,N_1023,N_1141);
xnor U1786 (N_1786,N_1448,N_1238);
or U1787 (N_1787,N_1083,N_1471);
or U1788 (N_1788,N_1194,N_1232);
and U1789 (N_1789,N_1093,N_1389);
nor U1790 (N_1790,N_1432,N_1233);
nor U1791 (N_1791,N_1183,N_1456);
nand U1792 (N_1792,N_1434,N_1367);
and U1793 (N_1793,N_1284,N_1238);
nand U1794 (N_1794,N_1309,N_1267);
and U1795 (N_1795,N_1356,N_1233);
and U1796 (N_1796,N_1304,N_1411);
or U1797 (N_1797,N_1070,N_1025);
nor U1798 (N_1798,N_1363,N_1167);
nand U1799 (N_1799,N_1046,N_1479);
nand U1800 (N_1800,N_1219,N_1230);
nor U1801 (N_1801,N_1161,N_1300);
and U1802 (N_1802,N_1300,N_1098);
and U1803 (N_1803,N_1270,N_1258);
and U1804 (N_1804,N_1124,N_1411);
nand U1805 (N_1805,N_1140,N_1101);
nand U1806 (N_1806,N_1106,N_1146);
xor U1807 (N_1807,N_1231,N_1381);
or U1808 (N_1808,N_1388,N_1105);
nand U1809 (N_1809,N_1386,N_1279);
or U1810 (N_1810,N_1446,N_1217);
xnor U1811 (N_1811,N_1062,N_1329);
nor U1812 (N_1812,N_1330,N_1074);
nor U1813 (N_1813,N_1019,N_1104);
xor U1814 (N_1814,N_1150,N_1422);
nand U1815 (N_1815,N_1032,N_1320);
nor U1816 (N_1816,N_1031,N_1181);
nand U1817 (N_1817,N_1433,N_1381);
and U1818 (N_1818,N_1346,N_1117);
nand U1819 (N_1819,N_1292,N_1494);
or U1820 (N_1820,N_1161,N_1108);
and U1821 (N_1821,N_1207,N_1306);
nor U1822 (N_1822,N_1456,N_1483);
nor U1823 (N_1823,N_1455,N_1140);
nor U1824 (N_1824,N_1405,N_1189);
and U1825 (N_1825,N_1062,N_1015);
nor U1826 (N_1826,N_1182,N_1499);
nor U1827 (N_1827,N_1206,N_1496);
and U1828 (N_1828,N_1008,N_1403);
nand U1829 (N_1829,N_1057,N_1349);
or U1830 (N_1830,N_1309,N_1411);
or U1831 (N_1831,N_1361,N_1063);
or U1832 (N_1832,N_1432,N_1016);
nor U1833 (N_1833,N_1149,N_1226);
nand U1834 (N_1834,N_1356,N_1393);
nor U1835 (N_1835,N_1057,N_1195);
or U1836 (N_1836,N_1273,N_1225);
nand U1837 (N_1837,N_1444,N_1279);
nand U1838 (N_1838,N_1317,N_1038);
nor U1839 (N_1839,N_1041,N_1468);
and U1840 (N_1840,N_1066,N_1150);
nand U1841 (N_1841,N_1228,N_1251);
nor U1842 (N_1842,N_1105,N_1223);
xnor U1843 (N_1843,N_1386,N_1321);
nand U1844 (N_1844,N_1192,N_1076);
or U1845 (N_1845,N_1034,N_1225);
nand U1846 (N_1846,N_1131,N_1082);
nor U1847 (N_1847,N_1236,N_1080);
and U1848 (N_1848,N_1043,N_1337);
nand U1849 (N_1849,N_1386,N_1195);
or U1850 (N_1850,N_1416,N_1056);
nor U1851 (N_1851,N_1130,N_1452);
and U1852 (N_1852,N_1095,N_1159);
and U1853 (N_1853,N_1423,N_1282);
and U1854 (N_1854,N_1170,N_1101);
and U1855 (N_1855,N_1153,N_1089);
or U1856 (N_1856,N_1021,N_1029);
or U1857 (N_1857,N_1370,N_1479);
and U1858 (N_1858,N_1416,N_1321);
nor U1859 (N_1859,N_1296,N_1082);
nor U1860 (N_1860,N_1016,N_1469);
or U1861 (N_1861,N_1281,N_1221);
or U1862 (N_1862,N_1078,N_1391);
nand U1863 (N_1863,N_1038,N_1393);
nor U1864 (N_1864,N_1186,N_1026);
or U1865 (N_1865,N_1465,N_1368);
or U1866 (N_1866,N_1477,N_1086);
nor U1867 (N_1867,N_1337,N_1455);
and U1868 (N_1868,N_1209,N_1311);
or U1869 (N_1869,N_1352,N_1253);
nor U1870 (N_1870,N_1277,N_1355);
nor U1871 (N_1871,N_1274,N_1241);
nand U1872 (N_1872,N_1172,N_1048);
nand U1873 (N_1873,N_1451,N_1122);
nor U1874 (N_1874,N_1149,N_1044);
nor U1875 (N_1875,N_1061,N_1053);
and U1876 (N_1876,N_1405,N_1403);
and U1877 (N_1877,N_1234,N_1300);
nand U1878 (N_1878,N_1384,N_1389);
nor U1879 (N_1879,N_1496,N_1181);
nand U1880 (N_1880,N_1065,N_1031);
xnor U1881 (N_1881,N_1246,N_1311);
and U1882 (N_1882,N_1299,N_1119);
nand U1883 (N_1883,N_1055,N_1119);
and U1884 (N_1884,N_1341,N_1204);
and U1885 (N_1885,N_1355,N_1258);
nor U1886 (N_1886,N_1326,N_1171);
nand U1887 (N_1887,N_1304,N_1112);
or U1888 (N_1888,N_1124,N_1104);
or U1889 (N_1889,N_1258,N_1180);
nand U1890 (N_1890,N_1273,N_1236);
nor U1891 (N_1891,N_1241,N_1263);
or U1892 (N_1892,N_1422,N_1499);
nor U1893 (N_1893,N_1308,N_1062);
nor U1894 (N_1894,N_1441,N_1251);
nor U1895 (N_1895,N_1091,N_1461);
and U1896 (N_1896,N_1161,N_1145);
or U1897 (N_1897,N_1491,N_1327);
nand U1898 (N_1898,N_1215,N_1133);
nor U1899 (N_1899,N_1288,N_1281);
nand U1900 (N_1900,N_1311,N_1166);
nand U1901 (N_1901,N_1335,N_1491);
or U1902 (N_1902,N_1435,N_1441);
or U1903 (N_1903,N_1379,N_1167);
nand U1904 (N_1904,N_1121,N_1291);
and U1905 (N_1905,N_1064,N_1231);
nor U1906 (N_1906,N_1065,N_1306);
or U1907 (N_1907,N_1048,N_1209);
nor U1908 (N_1908,N_1381,N_1141);
or U1909 (N_1909,N_1303,N_1068);
or U1910 (N_1910,N_1008,N_1090);
nor U1911 (N_1911,N_1042,N_1441);
or U1912 (N_1912,N_1019,N_1178);
nand U1913 (N_1913,N_1444,N_1072);
nand U1914 (N_1914,N_1483,N_1376);
xnor U1915 (N_1915,N_1386,N_1033);
and U1916 (N_1916,N_1374,N_1445);
and U1917 (N_1917,N_1404,N_1178);
and U1918 (N_1918,N_1113,N_1004);
and U1919 (N_1919,N_1132,N_1184);
nand U1920 (N_1920,N_1034,N_1494);
nand U1921 (N_1921,N_1142,N_1129);
nand U1922 (N_1922,N_1249,N_1358);
and U1923 (N_1923,N_1003,N_1400);
nor U1924 (N_1924,N_1177,N_1363);
nor U1925 (N_1925,N_1135,N_1000);
nor U1926 (N_1926,N_1200,N_1289);
and U1927 (N_1927,N_1439,N_1052);
or U1928 (N_1928,N_1098,N_1192);
xor U1929 (N_1929,N_1083,N_1152);
nand U1930 (N_1930,N_1326,N_1042);
and U1931 (N_1931,N_1152,N_1273);
nand U1932 (N_1932,N_1032,N_1202);
or U1933 (N_1933,N_1325,N_1416);
and U1934 (N_1934,N_1237,N_1242);
xor U1935 (N_1935,N_1407,N_1364);
or U1936 (N_1936,N_1047,N_1145);
and U1937 (N_1937,N_1198,N_1419);
nand U1938 (N_1938,N_1259,N_1102);
nor U1939 (N_1939,N_1056,N_1000);
nor U1940 (N_1940,N_1491,N_1354);
and U1941 (N_1941,N_1257,N_1124);
or U1942 (N_1942,N_1446,N_1462);
nor U1943 (N_1943,N_1414,N_1069);
nand U1944 (N_1944,N_1105,N_1429);
nor U1945 (N_1945,N_1278,N_1247);
nand U1946 (N_1946,N_1246,N_1410);
nor U1947 (N_1947,N_1031,N_1385);
nor U1948 (N_1948,N_1119,N_1147);
nand U1949 (N_1949,N_1346,N_1272);
nor U1950 (N_1950,N_1026,N_1431);
nand U1951 (N_1951,N_1145,N_1458);
xnor U1952 (N_1952,N_1374,N_1414);
nand U1953 (N_1953,N_1152,N_1338);
or U1954 (N_1954,N_1287,N_1141);
nor U1955 (N_1955,N_1414,N_1495);
nor U1956 (N_1956,N_1233,N_1490);
nand U1957 (N_1957,N_1369,N_1041);
nor U1958 (N_1958,N_1294,N_1326);
nand U1959 (N_1959,N_1330,N_1264);
nor U1960 (N_1960,N_1297,N_1137);
nor U1961 (N_1961,N_1261,N_1436);
nand U1962 (N_1962,N_1132,N_1488);
nor U1963 (N_1963,N_1182,N_1421);
nor U1964 (N_1964,N_1177,N_1345);
and U1965 (N_1965,N_1173,N_1089);
nor U1966 (N_1966,N_1316,N_1215);
or U1967 (N_1967,N_1151,N_1024);
and U1968 (N_1968,N_1084,N_1425);
nand U1969 (N_1969,N_1344,N_1432);
or U1970 (N_1970,N_1498,N_1167);
and U1971 (N_1971,N_1485,N_1305);
and U1972 (N_1972,N_1102,N_1437);
and U1973 (N_1973,N_1458,N_1176);
and U1974 (N_1974,N_1265,N_1457);
and U1975 (N_1975,N_1189,N_1076);
nor U1976 (N_1976,N_1424,N_1110);
nand U1977 (N_1977,N_1328,N_1431);
or U1978 (N_1978,N_1212,N_1139);
nor U1979 (N_1979,N_1085,N_1499);
or U1980 (N_1980,N_1410,N_1483);
nand U1981 (N_1981,N_1420,N_1312);
nand U1982 (N_1982,N_1335,N_1113);
nor U1983 (N_1983,N_1476,N_1206);
nand U1984 (N_1984,N_1033,N_1348);
nor U1985 (N_1985,N_1368,N_1447);
nor U1986 (N_1986,N_1449,N_1239);
nand U1987 (N_1987,N_1273,N_1174);
or U1988 (N_1988,N_1161,N_1353);
or U1989 (N_1989,N_1250,N_1119);
nor U1990 (N_1990,N_1256,N_1108);
or U1991 (N_1991,N_1058,N_1060);
nand U1992 (N_1992,N_1002,N_1349);
or U1993 (N_1993,N_1204,N_1038);
or U1994 (N_1994,N_1134,N_1430);
nor U1995 (N_1995,N_1378,N_1396);
nor U1996 (N_1996,N_1344,N_1119);
and U1997 (N_1997,N_1196,N_1213);
nand U1998 (N_1998,N_1042,N_1023);
nand U1999 (N_1999,N_1085,N_1422);
or U2000 (N_2000,N_1947,N_1965);
and U2001 (N_2001,N_1725,N_1964);
nand U2002 (N_2002,N_1738,N_1872);
nand U2003 (N_2003,N_1758,N_1993);
or U2004 (N_2004,N_1855,N_1522);
nor U2005 (N_2005,N_1541,N_1691);
nand U2006 (N_2006,N_1946,N_1882);
or U2007 (N_2007,N_1710,N_1692);
and U2008 (N_2008,N_1870,N_1874);
and U2009 (N_2009,N_1624,N_1625);
and U2010 (N_2010,N_1816,N_1718);
nor U2011 (N_2011,N_1622,N_1626);
and U2012 (N_2012,N_1927,N_1811);
or U2013 (N_2013,N_1999,N_1919);
and U2014 (N_2014,N_1835,N_1801);
nor U2015 (N_2015,N_1650,N_1614);
nor U2016 (N_2016,N_1575,N_1770);
or U2017 (N_2017,N_1950,N_1745);
nand U2018 (N_2018,N_1716,N_1617);
and U2019 (N_2019,N_1581,N_1956);
nand U2020 (N_2020,N_1648,N_1900);
nor U2021 (N_2021,N_1905,N_1852);
nor U2022 (N_2022,N_1539,N_1551);
and U2023 (N_2023,N_1748,N_1849);
or U2024 (N_2024,N_1721,N_1932);
or U2025 (N_2025,N_1991,N_1589);
nand U2026 (N_2026,N_1880,N_1657);
and U2027 (N_2027,N_1961,N_1808);
or U2028 (N_2028,N_1830,N_1684);
and U2029 (N_2029,N_1877,N_1963);
nand U2030 (N_2030,N_1634,N_1600);
or U2031 (N_2031,N_1926,N_1596);
or U2032 (N_2032,N_1747,N_1876);
nor U2033 (N_2033,N_1798,N_1968);
nand U2034 (N_2034,N_1777,N_1543);
nand U2035 (N_2035,N_1845,N_1854);
nor U2036 (N_2036,N_1733,N_1537);
nor U2037 (N_2037,N_1992,N_1916);
nand U2038 (N_2038,N_1520,N_1941);
or U2039 (N_2039,N_1586,N_1613);
nor U2040 (N_2040,N_1558,N_1731);
nand U2041 (N_2041,N_1741,N_1661);
or U2042 (N_2042,N_1720,N_1682);
or U2043 (N_2043,N_1860,N_1742);
and U2044 (N_2044,N_1579,N_1591);
nor U2045 (N_2045,N_1636,N_1750);
nand U2046 (N_2046,N_1853,N_1549);
nor U2047 (N_2047,N_1890,N_1995);
or U2048 (N_2048,N_1913,N_1670);
nand U2049 (N_2049,N_1989,N_1701);
nor U2050 (N_2050,N_1704,N_1669);
nor U2051 (N_2051,N_1793,N_1935);
and U2052 (N_2052,N_1667,N_1513);
nand U2053 (N_2053,N_1527,N_1676);
and U2054 (N_2054,N_1556,N_1826);
nor U2055 (N_2055,N_1775,N_1663);
nand U2056 (N_2056,N_1912,N_1978);
and U2057 (N_2057,N_1732,N_1842);
nand U2058 (N_2058,N_1555,N_1562);
nand U2059 (N_2059,N_1898,N_1807);
nand U2060 (N_2060,N_1547,N_1630);
or U2061 (N_2061,N_1871,N_1752);
nor U2062 (N_2062,N_1700,N_1837);
and U2063 (N_2063,N_1795,N_1531);
and U2064 (N_2064,N_1706,N_1683);
nand U2065 (N_2065,N_1550,N_1571);
and U2066 (N_2066,N_1792,N_1789);
nor U2067 (N_2067,N_1815,N_1885);
xnor U2068 (N_2068,N_1627,N_1938);
or U2069 (N_2069,N_1820,N_1615);
nor U2070 (N_2070,N_1583,N_1666);
nor U2071 (N_2071,N_1904,N_1560);
nand U2072 (N_2072,N_1573,N_1962);
and U2073 (N_2073,N_1759,N_1986);
and U2074 (N_2074,N_1894,N_1825);
nand U2075 (N_2075,N_1577,N_1569);
and U2076 (N_2076,N_1535,N_1867);
nand U2077 (N_2077,N_1698,N_1804);
and U2078 (N_2078,N_1847,N_1763);
nor U2079 (N_2079,N_1769,N_1843);
or U2080 (N_2080,N_1603,N_1781);
and U2081 (N_2081,N_1561,N_1973);
or U2082 (N_2082,N_1511,N_1509);
nand U2083 (N_2083,N_1857,N_1884);
or U2084 (N_2084,N_1695,N_1907);
nor U2085 (N_2085,N_1533,N_1996);
nand U2086 (N_2086,N_1639,N_1841);
nor U2087 (N_2087,N_1929,N_1552);
nand U2088 (N_2088,N_1590,N_1730);
nor U2089 (N_2089,N_1805,N_1505);
nand U2090 (N_2090,N_1608,N_1736);
or U2091 (N_2091,N_1887,N_1728);
nor U2092 (N_2092,N_1618,N_1844);
or U2093 (N_2093,N_1526,N_1909);
or U2094 (N_2094,N_1637,N_1969);
nor U2095 (N_2095,N_1580,N_1819);
nand U2096 (N_2096,N_1640,N_1754);
nor U2097 (N_2097,N_1799,N_1655);
xnor U2098 (N_2098,N_1516,N_1779);
xor U2099 (N_2099,N_1765,N_1506);
and U2100 (N_2100,N_1863,N_1631);
or U2101 (N_2101,N_1739,N_1914);
nand U2102 (N_2102,N_1931,N_1756);
or U2103 (N_2103,N_1515,N_1766);
and U2104 (N_2104,N_1800,N_1883);
or U2105 (N_2105,N_1861,N_1508);
nor U2106 (N_2106,N_1782,N_1990);
or U2107 (N_2107,N_1697,N_1559);
xor U2108 (N_2108,N_1671,N_1582);
and U2109 (N_2109,N_1501,N_1790);
nor U2110 (N_2110,N_1873,N_1729);
nor U2111 (N_2111,N_1967,N_1647);
or U2112 (N_2112,N_1868,N_1621);
or U2113 (N_2113,N_1974,N_1783);
and U2114 (N_2114,N_1619,N_1774);
nand U2115 (N_2115,N_1895,N_1784);
nand U2116 (N_2116,N_1584,N_1512);
xnor U2117 (N_2117,N_1760,N_1664);
nor U2118 (N_2118,N_1665,N_1719);
nand U2119 (N_2119,N_1681,N_1605);
and U2120 (N_2120,N_1532,N_1864);
nand U2121 (N_2121,N_1651,N_1534);
nand U2122 (N_2122,N_1940,N_1524);
and U2123 (N_2123,N_1859,N_1960);
nand U2124 (N_2124,N_1910,N_1565);
nand U2125 (N_2125,N_1821,N_1972);
nor U2126 (N_2126,N_1711,N_1881);
or U2127 (N_2127,N_1628,N_1834);
or U2128 (N_2128,N_1921,N_1553);
or U2129 (N_2129,N_1544,N_1983);
nor U2130 (N_2130,N_1592,N_1839);
and U2131 (N_2131,N_1578,N_1817);
nand U2132 (N_2132,N_1942,N_1959);
nor U2133 (N_2133,N_1893,N_1680);
or U2134 (N_2134,N_1542,N_1674);
nor U2135 (N_2135,N_1629,N_1502);
nand U2136 (N_2136,N_1948,N_1813);
or U2137 (N_2137,N_1705,N_1862);
nor U2138 (N_2138,N_1500,N_1507);
and U2139 (N_2139,N_1944,N_1724);
and U2140 (N_2140,N_1751,N_1797);
nand U2141 (N_2141,N_1928,N_1521);
nor U2142 (N_2142,N_1635,N_1897);
nand U2143 (N_2143,N_1593,N_1656);
nand U2144 (N_2144,N_1977,N_1930);
nor U2145 (N_2145,N_1755,N_1994);
nand U2146 (N_2146,N_1952,N_1924);
nor U2147 (N_2147,N_1778,N_1903);
and U2148 (N_2148,N_1675,N_1594);
nor U2149 (N_2149,N_1823,N_1540);
nand U2150 (N_2150,N_1828,N_1984);
nand U2151 (N_2151,N_1557,N_1574);
and U2152 (N_2152,N_1970,N_1660);
and U2153 (N_2153,N_1850,N_1564);
nor U2154 (N_2154,N_1519,N_1686);
nor U2155 (N_2155,N_1523,N_1632);
and U2156 (N_2156,N_1891,N_1567);
nand U2157 (N_2157,N_1827,N_1764);
nor U2158 (N_2158,N_1875,N_1818);
nand U2159 (N_2159,N_1988,N_1685);
nand U2160 (N_2160,N_1749,N_1982);
nor U2161 (N_2161,N_1514,N_1727);
and U2162 (N_2162,N_1794,N_1997);
or U2163 (N_2163,N_1901,N_1953);
nor U2164 (N_2164,N_1677,N_1786);
nand U2165 (N_2165,N_1712,N_1643);
nor U2166 (N_2166,N_1937,N_1714);
nor U2167 (N_2167,N_1906,N_1803);
and U2168 (N_2168,N_1696,N_1642);
xnor U2169 (N_2169,N_1856,N_1971);
nor U2170 (N_2170,N_1693,N_1546);
or U2171 (N_2171,N_1673,N_1788);
nor U2172 (N_2172,N_1588,N_1679);
nor U2173 (N_2173,N_1776,N_1886);
and U2174 (N_2174,N_1858,N_1644);
nor U2175 (N_2175,N_1746,N_1672);
nor U2176 (N_2176,N_1908,N_1915);
and U2177 (N_2177,N_1899,N_1998);
and U2178 (N_2178,N_1652,N_1572);
nor U2179 (N_2179,N_1662,N_1517);
and U2180 (N_2180,N_1668,N_1772);
and U2181 (N_2181,N_1824,N_1678);
nor U2182 (N_2182,N_1773,N_1762);
or U2183 (N_2183,N_1703,N_1954);
and U2184 (N_2184,N_1722,N_1570);
nor U2185 (N_2185,N_1585,N_1641);
or U2186 (N_2186,N_1687,N_1529);
nor U2187 (N_2187,N_1735,N_1918);
nand U2188 (N_2188,N_1838,N_1743);
nand U2189 (N_2189,N_1945,N_1598);
or U2190 (N_2190,N_1923,N_1925);
nand U2191 (N_2191,N_1538,N_1865);
nand U2192 (N_2192,N_1768,N_1576);
nor U2193 (N_2193,N_1814,N_1638);
or U2194 (N_2194,N_1757,N_1958);
nand U2195 (N_2195,N_1688,N_1610);
nor U2196 (N_2196,N_1896,N_1597);
and U2197 (N_2197,N_1806,N_1831);
and U2198 (N_2198,N_1510,N_1771);
or U2199 (N_2199,N_1653,N_1791);
or U2200 (N_2200,N_1933,N_1889);
nand U2201 (N_2201,N_1654,N_1699);
nor U2202 (N_2202,N_1980,N_1737);
and U2203 (N_2203,N_1911,N_1554);
or U2204 (N_2204,N_1602,N_1796);
xnor U2205 (N_2205,N_1633,N_1702);
nor U2206 (N_2206,N_1659,N_1694);
nor U2207 (N_2207,N_1545,N_1604);
nand U2208 (N_2208,N_1595,N_1740);
and U2209 (N_2209,N_1611,N_1620);
or U2210 (N_2210,N_1785,N_1949);
or U2211 (N_2211,N_1902,N_1734);
nor U2212 (N_2212,N_1787,N_1943);
and U2213 (N_2213,N_1708,N_1832);
nand U2214 (N_2214,N_1726,N_1690);
nor U2215 (N_2215,N_1566,N_1528);
nand U2216 (N_2216,N_1623,N_1936);
or U2217 (N_2217,N_1536,N_1985);
or U2218 (N_2218,N_1518,N_1599);
and U2219 (N_2219,N_1869,N_1836);
nor U2220 (N_2220,N_1723,N_1548);
nor U2221 (N_2221,N_1616,N_1846);
nor U2222 (N_2222,N_1976,N_1645);
and U2223 (N_2223,N_1892,N_1504);
nor U2224 (N_2224,N_1525,N_1987);
nor U2225 (N_2225,N_1713,N_1957);
and U2226 (N_2226,N_1809,N_1646);
or U2227 (N_2227,N_1833,N_1607);
nor U2228 (N_2228,N_1802,N_1568);
nor U2229 (N_2229,N_1866,N_1606);
nor U2230 (N_2230,N_1879,N_1812);
nand U2231 (N_2231,N_1709,N_1851);
or U2232 (N_2232,N_1587,N_1767);
and U2233 (N_2233,N_1753,N_1689);
and U2234 (N_2234,N_1979,N_1966);
or U2235 (N_2235,N_1780,N_1878);
nand U2236 (N_2236,N_1658,N_1955);
nor U2237 (N_2237,N_1934,N_1939);
nor U2238 (N_2238,N_1810,N_1888);
or U2239 (N_2239,N_1922,N_1920);
and U2240 (N_2240,N_1829,N_1612);
nor U2241 (N_2241,N_1822,N_1649);
nor U2242 (N_2242,N_1609,N_1917);
or U2243 (N_2243,N_1563,N_1530);
or U2244 (N_2244,N_1761,N_1744);
nand U2245 (N_2245,N_1951,N_1601);
nor U2246 (N_2246,N_1715,N_1981);
or U2247 (N_2247,N_1840,N_1848);
or U2248 (N_2248,N_1717,N_1975);
nand U2249 (N_2249,N_1707,N_1503);
nor U2250 (N_2250,N_1916,N_1612);
nand U2251 (N_2251,N_1683,N_1619);
nor U2252 (N_2252,N_1738,N_1559);
nor U2253 (N_2253,N_1558,N_1936);
nor U2254 (N_2254,N_1954,N_1957);
nand U2255 (N_2255,N_1885,N_1705);
or U2256 (N_2256,N_1872,N_1644);
and U2257 (N_2257,N_1909,N_1574);
and U2258 (N_2258,N_1521,N_1923);
or U2259 (N_2259,N_1963,N_1620);
and U2260 (N_2260,N_1740,N_1957);
nor U2261 (N_2261,N_1531,N_1985);
or U2262 (N_2262,N_1809,N_1702);
or U2263 (N_2263,N_1594,N_1617);
nor U2264 (N_2264,N_1742,N_1624);
nor U2265 (N_2265,N_1820,N_1895);
and U2266 (N_2266,N_1601,N_1547);
nand U2267 (N_2267,N_1678,N_1967);
nor U2268 (N_2268,N_1576,N_1835);
nor U2269 (N_2269,N_1770,N_1574);
nand U2270 (N_2270,N_1940,N_1700);
or U2271 (N_2271,N_1841,N_1548);
or U2272 (N_2272,N_1993,N_1665);
nand U2273 (N_2273,N_1784,N_1946);
nor U2274 (N_2274,N_1923,N_1912);
or U2275 (N_2275,N_1707,N_1681);
and U2276 (N_2276,N_1848,N_1568);
or U2277 (N_2277,N_1803,N_1935);
nor U2278 (N_2278,N_1604,N_1661);
or U2279 (N_2279,N_1660,N_1679);
or U2280 (N_2280,N_1630,N_1991);
nand U2281 (N_2281,N_1839,N_1533);
nor U2282 (N_2282,N_1870,N_1817);
and U2283 (N_2283,N_1709,N_1926);
nand U2284 (N_2284,N_1773,N_1578);
and U2285 (N_2285,N_1765,N_1705);
xor U2286 (N_2286,N_1538,N_1629);
and U2287 (N_2287,N_1844,N_1677);
and U2288 (N_2288,N_1925,N_1808);
and U2289 (N_2289,N_1760,N_1811);
or U2290 (N_2290,N_1970,N_1746);
nor U2291 (N_2291,N_1820,N_1732);
or U2292 (N_2292,N_1567,N_1594);
nor U2293 (N_2293,N_1986,N_1720);
nand U2294 (N_2294,N_1878,N_1621);
nor U2295 (N_2295,N_1610,N_1975);
or U2296 (N_2296,N_1883,N_1768);
nor U2297 (N_2297,N_1682,N_1730);
or U2298 (N_2298,N_1549,N_1679);
and U2299 (N_2299,N_1667,N_1985);
and U2300 (N_2300,N_1519,N_1658);
and U2301 (N_2301,N_1998,N_1577);
nand U2302 (N_2302,N_1764,N_1786);
or U2303 (N_2303,N_1965,N_1708);
xor U2304 (N_2304,N_1835,N_1505);
nand U2305 (N_2305,N_1578,N_1506);
nand U2306 (N_2306,N_1892,N_1526);
nand U2307 (N_2307,N_1601,N_1636);
or U2308 (N_2308,N_1894,N_1889);
nor U2309 (N_2309,N_1650,N_1566);
or U2310 (N_2310,N_1663,N_1544);
nor U2311 (N_2311,N_1837,N_1754);
nand U2312 (N_2312,N_1723,N_1916);
or U2313 (N_2313,N_1862,N_1913);
and U2314 (N_2314,N_1535,N_1847);
nor U2315 (N_2315,N_1686,N_1760);
or U2316 (N_2316,N_1824,N_1804);
nand U2317 (N_2317,N_1934,N_1543);
or U2318 (N_2318,N_1656,N_1755);
or U2319 (N_2319,N_1579,N_1622);
nor U2320 (N_2320,N_1846,N_1640);
xor U2321 (N_2321,N_1669,N_1803);
and U2322 (N_2322,N_1722,N_1642);
or U2323 (N_2323,N_1510,N_1610);
nor U2324 (N_2324,N_1535,N_1646);
or U2325 (N_2325,N_1974,N_1816);
or U2326 (N_2326,N_1948,N_1566);
nand U2327 (N_2327,N_1533,N_1584);
or U2328 (N_2328,N_1617,N_1549);
nand U2329 (N_2329,N_1513,N_1771);
xnor U2330 (N_2330,N_1722,N_1923);
and U2331 (N_2331,N_1656,N_1757);
xor U2332 (N_2332,N_1662,N_1778);
or U2333 (N_2333,N_1905,N_1733);
nor U2334 (N_2334,N_1725,N_1970);
or U2335 (N_2335,N_1670,N_1986);
and U2336 (N_2336,N_1650,N_1887);
or U2337 (N_2337,N_1634,N_1824);
nand U2338 (N_2338,N_1541,N_1654);
nand U2339 (N_2339,N_1798,N_1766);
nand U2340 (N_2340,N_1514,N_1782);
nand U2341 (N_2341,N_1938,N_1591);
nand U2342 (N_2342,N_1857,N_1859);
nand U2343 (N_2343,N_1539,N_1929);
nand U2344 (N_2344,N_1561,N_1971);
or U2345 (N_2345,N_1966,N_1719);
or U2346 (N_2346,N_1597,N_1997);
or U2347 (N_2347,N_1656,N_1840);
nor U2348 (N_2348,N_1916,N_1555);
xor U2349 (N_2349,N_1723,N_1810);
and U2350 (N_2350,N_1720,N_1750);
nor U2351 (N_2351,N_1903,N_1593);
and U2352 (N_2352,N_1593,N_1500);
or U2353 (N_2353,N_1788,N_1789);
or U2354 (N_2354,N_1969,N_1874);
and U2355 (N_2355,N_1906,N_1891);
nor U2356 (N_2356,N_1912,N_1595);
nor U2357 (N_2357,N_1943,N_1965);
and U2358 (N_2358,N_1691,N_1864);
nand U2359 (N_2359,N_1647,N_1758);
and U2360 (N_2360,N_1733,N_1713);
or U2361 (N_2361,N_1886,N_1771);
nand U2362 (N_2362,N_1991,N_1869);
nand U2363 (N_2363,N_1854,N_1707);
nor U2364 (N_2364,N_1841,N_1816);
nand U2365 (N_2365,N_1731,N_1692);
nand U2366 (N_2366,N_1746,N_1674);
nor U2367 (N_2367,N_1565,N_1557);
and U2368 (N_2368,N_1876,N_1650);
or U2369 (N_2369,N_1511,N_1732);
nand U2370 (N_2370,N_1603,N_1794);
and U2371 (N_2371,N_1691,N_1913);
nor U2372 (N_2372,N_1701,N_1985);
and U2373 (N_2373,N_1623,N_1569);
and U2374 (N_2374,N_1629,N_1733);
or U2375 (N_2375,N_1522,N_1969);
nand U2376 (N_2376,N_1556,N_1917);
and U2377 (N_2377,N_1843,N_1589);
and U2378 (N_2378,N_1984,N_1633);
xnor U2379 (N_2379,N_1693,N_1518);
or U2380 (N_2380,N_1922,N_1588);
and U2381 (N_2381,N_1811,N_1708);
and U2382 (N_2382,N_1600,N_1728);
nor U2383 (N_2383,N_1943,N_1791);
nand U2384 (N_2384,N_1978,N_1940);
nor U2385 (N_2385,N_1714,N_1628);
and U2386 (N_2386,N_1967,N_1663);
or U2387 (N_2387,N_1665,N_1734);
or U2388 (N_2388,N_1764,N_1970);
nor U2389 (N_2389,N_1869,N_1934);
nand U2390 (N_2390,N_1850,N_1639);
xor U2391 (N_2391,N_1856,N_1830);
or U2392 (N_2392,N_1908,N_1519);
or U2393 (N_2393,N_1647,N_1888);
and U2394 (N_2394,N_1770,N_1819);
nor U2395 (N_2395,N_1634,N_1656);
or U2396 (N_2396,N_1672,N_1737);
nor U2397 (N_2397,N_1937,N_1622);
nor U2398 (N_2398,N_1930,N_1925);
nor U2399 (N_2399,N_1539,N_1691);
and U2400 (N_2400,N_1798,N_1838);
xnor U2401 (N_2401,N_1660,N_1984);
or U2402 (N_2402,N_1796,N_1527);
and U2403 (N_2403,N_1600,N_1897);
nor U2404 (N_2404,N_1927,N_1574);
or U2405 (N_2405,N_1905,N_1917);
or U2406 (N_2406,N_1535,N_1738);
and U2407 (N_2407,N_1804,N_1520);
and U2408 (N_2408,N_1614,N_1640);
or U2409 (N_2409,N_1559,N_1557);
nor U2410 (N_2410,N_1823,N_1853);
or U2411 (N_2411,N_1513,N_1744);
nor U2412 (N_2412,N_1712,N_1862);
and U2413 (N_2413,N_1707,N_1775);
and U2414 (N_2414,N_1736,N_1546);
nor U2415 (N_2415,N_1906,N_1876);
nand U2416 (N_2416,N_1783,N_1954);
or U2417 (N_2417,N_1564,N_1589);
or U2418 (N_2418,N_1863,N_1710);
nand U2419 (N_2419,N_1746,N_1857);
nor U2420 (N_2420,N_1968,N_1938);
or U2421 (N_2421,N_1754,N_1890);
or U2422 (N_2422,N_1934,N_1680);
nor U2423 (N_2423,N_1813,N_1859);
nor U2424 (N_2424,N_1620,N_1762);
nand U2425 (N_2425,N_1795,N_1624);
and U2426 (N_2426,N_1922,N_1873);
nor U2427 (N_2427,N_1918,N_1634);
or U2428 (N_2428,N_1989,N_1694);
or U2429 (N_2429,N_1928,N_1594);
nor U2430 (N_2430,N_1754,N_1574);
nor U2431 (N_2431,N_1640,N_1998);
or U2432 (N_2432,N_1738,N_1815);
or U2433 (N_2433,N_1986,N_1929);
and U2434 (N_2434,N_1942,N_1591);
nand U2435 (N_2435,N_1935,N_1701);
or U2436 (N_2436,N_1943,N_1702);
and U2437 (N_2437,N_1810,N_1649);
nand U2438 (N_2438,N_1828,N_1551);
or U2439 (N_2439,N_1715,N_1797);
nand U2440 (N_2440,N_1887,N_1882);
nor U2441 (N_2441,N_1854,N_1777);
and U2442 (N_2442,N_1508,N_1551);
or U2443 (N_2443,N_1894,N_1988);
or U2444 (N_2444,N_1756,N_1564);
or U2445 (N_2445,N_1657,N_1717);
nand U2446 (N_2446,N_1518,N_1728);
and U2447 (N_2447,N_1873,N_1994);
or U2448 (N_2448,N_1583,N_1831);
nand U2449 (N_2449,N_1535,N_1852);
nand U2450 (N_2450,N_1868,N_1928);
or U2451 (N_2451,N_1606,N_1731);
nor U2452 (N_2452,N_1781,N_1902);
and U2453 (N_2453,N_1886,N_1778);
and U2454 (N_2454,N_1739,N_1549);
nor U2455 (N_2455,N_1541,N_1987);
and U2456 (N_2456,N_1884,N_1747);
or U2457 (N_2457,N_1963,N_1817);
nand U2458 (N_2458,N_1854,N_1681);
nor U2459 (N_2459,N_1587,N_1826);
nand U2460 (N_2460,N_1701,N_1895);
nand U2461 (N_2461,N_1532,N_1796);
and U2462 (N_2462,N_1779,N_1886);
or U2463 (N_2463,N_1916,N_1941);
or U2464 (N_2464,N_1574,N_1609);
or U2465 (N_2465,N_1763,N_1989);
or U2466 (N_2466,N_1884,N_1892);
and U2467 (N_2467,N_1983,N_1515);
nor U2468 (N_2468,N_1852,N_1503);
or U2469 (N_2469,N_1536,N_1838);
or U2470 (N_2470,N_1956,N_1896);
nand U2471 (N_2471,N_1782,N_1932);
and U2472 (N_2472,N_1996,N_1797);
and U2473 (N_2473,N_1579,N_1643);
nand U2474 (N_2474,N_1525,N_1865);
xor U2475 (N_2475,N_1975,N_1571);
and U2476 (N_2476,N_1762,N_1610);
nand U2477 (N_2477,N_1802,N_1629);
or U2478 (N_2478,N_1697,N_1658);
nor U2479 (N_2479,N_1863,N_1683);
or U2480 (N_2480,N_1545,N_1655);
nand U2481 (N_2481,N_1709,N_1591);
nand U2482 (N_2482,N_1798,N_1666);
or U2483 (N_2483,N_1900,N_1552);
nand U2484 (N_2484,N_1726,N_1982);
and U2485 (N_2485,N_1876,N_1947);
and U2486 (N_2486,N_1939,N_1536);
nand U2487 (N_2487,N_1969,N_1892);
nand U2488 (N_2488,N_1895,N_1530);
nor U2489 (N_2489,N_1708,N_1918);
or U2490 (N_2490,N_1993,N_1945);
or U2491 (N_2491,N_1820,N_1643);
nor U2492 (N_2492,N_1966,N_1754);
nand U2493 (N_2493,N_1562,N_1678);
or U2494 (N_2494,N_1520,N_1887);
or U2495 (N_2495,N_1818,N_1660);
nand U2496 (N_2496,N_1966,N_1671);
and U2497 (N_2497,N_1751,N_1955);
and U2498 (N_2498,N_1546,N_1723);
nor U2499 (N_2499,N_1910,N_1822);
and U2500 (N_2500,N_2350,N_2005);
and U2501 (N_2501,N_2296,N_2078);
nor U2502 (N_2502,N_2135,N_2320);
nand U2503 (N_2503,N_2165,N_2129);
nor U2504 (N_2504,N_2010,N_2204);
or U2505 (N_2505,N_2409,N_2353);
nand U2506 (N_2506,N_2289,N_2406);
xor U2507 (N_2507,N_2214,N_2004);
nor U2508 (N_2508,N_2140,N_2325);
nor U2509 (N_2509,N_2461,N_2341);
or U2510 (N_2510,N_2076,N_2260);
and U2511 (N_2511,N_2039,N_2047);
or U2512 (N_2512,N_2456,N_2372);
and U2513 (N_2513,N_2333,N_2332);
or U2514 (N_2514,N_2153,N_2079);
nand U2515 (N_2515,N_2111,N_2142);
and U2516 (N_2516,N_2432,N_2403);
or U2517 (N_2517,N_2478,N_2218);
xor U2518 (N_2518,N_2200,N_2131);
nor U2519 (N_2519,N_2173,N_2246);
or U2520 (N_2520,N_2171,N_2124);
nor U2521 (N_2521,N_2477,N_2217);
or U2522 (N_2522,N_2343,N_2418);
or U2523 (N_2523,N_2286,N_2197);
xor U2524 (N_2524,N_2185,N_2376);
or U2525 (N_2525,N_2150,N_2455);
and U2526 (N_2526,N_2147,N_2479);
or U2527 (N_2527,N_2169,N_2349);
and U2528 (N_2528,N_2265,N_2025);
and U2529 (N_2529,N_2112,N_2064);
nor U2530 (N_2530,N_2364,N_2166);
and U2531 (N_2531,N_2449,N_2283);
nor U2532 (N_2532,N_2100,N_2253);
and U2533 (N_2533,N_2020,N_2107);
nor U2534 (N_2534,N_2399,N_2168);
nand U2535 (N_2535,N_2413,N_2003);
and U2536 (N_2536,N_2336,N_2271);
or U2537 (N_2537,N_2037,N_2300);
nor U2538 (N_2538,N_2021,N_2034);
nand U2539 (N_2539,N_2338,N_2137);
or U2540 (N_2540,N_2266,N_2091);
nand U2541 (N_2541,N_2408,N_2414);
and U2542 (N_2542,N_2314,N_2030);
nor U2543 (N_2543,N_2081,N_2292);
nand U2544 (N_2544,N_2105,N_2396);
nor U2545 (N_2545,N_2213,N_2211);
nand U2546 (N_2546,N_2497,N_2101);
and U2547 (N_2547,N_2278,N_2201);
or U2548 (N_2548,N_2486,N_2196);
nor U2549 (N_2549,N_2002,N_2464);
or U2550 (N_2550,N_2476,N_2309);
nand U2551 (N_2551,N_2389,N_2382);
and U2552 (N_2552,N_2006,N_2458);
or U2553 (N_2553,N_2095,N_2352);
xnor U2554 (N_2554,N_2245,N_2425);
or U2555 (N_2555,N_2381,N_2075);
and U2556 (N_2556,N_2182,N_2344);
nor U2557 (N_2557,N_2008,N_2264);
nand U2558 (N_2558,N_2489,N_2239);
or U2559 (N_2559,N_2454,N_2295);
and U2560 (N_2560,N_2402,N_2102);
nand U2561 (N_2561,N_2334,N_2090);
and U2562 (N_2562,N_2015,N_2386);
nor U2563 (N_2563,N_2206,N_2322);
and U2564 (N_2564,N_2234,N_2238);
or U2565 (N_2565,N_2035,N_2189);
xnor U2566 (N_2566,N_2326,N_2146);
nand U2567 (N_2567,N_2345,N_2491);
nand U2568 (N_2568,N_2466,N_2248);
nor U2569 (N_2569,N_2080,N_2063);
xnor U2570 (N_2570,N_2235,N_2417);
nand U2571 (N_2571,N_2280,N_2226);
nor U2572 (N_2572,N_2054,N_2138);
and U2573 (N_2573,N_2068,N_2220);
nand U2574 (N_2574,N_2244,N_2184);
nor U2575 (N_2575,N_2016,N_2032);
and U2576 (N_2576,N_2052,N_2222);
nand U2577 (N_2577,N_2228,N_2074);
or U2578 (N_2578,N_2041,N_2242);
or U2579 (N_2579,N_2042,N_2324);
and U2580 (N_2580,N_2293,N_2066);
nor U2581 (N_2581,N_2070,N_2116);
nand U2582 (N_2582,N_2391,N_2415);
xor U2583 (N_2583,N_2272,N_2233);
or U2584 (N_2584,N_2269,N_2367);
and U2585 (N_2585,N_2323,N_2291);
nor U2586 (N_2586,N_2436,N_2018);
or U2587 (N_2587,N_2001,N_2475);
xnor U2588 (N_2588,N_2487,N_2051);
xor U2589 (N_2589,N_2420,N_2268);
and U2590 (N_2590,N_2401,N_2071);
and U2591 (N_2591,N_2232,N_2328);
nand U2592 (N_2592,N_2430,N_2306);
nand U2593 (N_2593,N_2469,N_2368);
nor U2594 (N_2594,N_2434,N_2060);
and U2595 (N_2595,N_2160,N_2251);
or U2596 (N_2596,N_2023,N_2067);
nor U2597 (N_2597,N_2031,N_2227);
nor U2598 (N_2598,N_2050,N_2249);
and U2599 (N_2599,N_2261,N_2256);
and U2600 (N_2600,N_2044,N_2488);
nor U2601 (N_2601,N_2317,N_2483);
or U2602 (N_2602,N_2086,N_2012);
or U2603 (N_2603,N_2433,N_2384);
nor U2604 (N_2604,N_2207,N_2127);
nand U2605 (N_2605,N_2045,N_2318);
nor U2606 (N_2606,N_2453,N_2115);
nand U2607 (N_2607,N_2462,N_2022);
or U2608 (N_2608,N_2029,N_2307);
or U2609 (N_2609,N_2040,N_2496);
nand U2610 (N_2610,N_2194,N_2495);
nor U2611 (N_2611,N_2250,N_2036);
nand U2612 (N_2612,N_2437,N_2121);
and U2613 (N_2613,N_2210,N_2172);
xnor U2614 (N_2614,N_2387,N_2471);
or U2615 (N_2615,N_2277,N_2321);
nor U2616 (N_2616,N_2069,N_2099);
xor U2617 (N_2617,N_2059,N_2442);
nor U2618 (N_2618,N_2118,N_2061);
or U2619 (N_2619,N_2065,N_2311);
or U2620 (N_2620,N_2457,N_2017);
or U2621 (N_2621,N_2445,N_2164);
nor U2622 (N_2622,N_2428,N_2084);
nor U2623 (N_2623,N_2013,N_2410);
or U2624 (N_2624,N_2092,N_2177);
nand U2625 (N_2625,N_2103,N_2247);
nand U2626 (N_2626,N_2011,N_2043);
nand U2627 (N_2627,N_2120,N_2148);
nor U2628 (N_2628,N_2082,N_2134);
xnor U2629 (N_2629,N_2459,N_2114);
or U2630 (N_2630,N_2240,N_2481);
and U2631 (N_2631,N_2024,N_2360);
nor U2632 (N_2632,N_2363,N_2374);
and U2633 (N_2633,N_2499,N_2305);
and U2634 (N_2634,N_2405,N_2474);
or U2635 (N_2635,N_2198,N_2274);
and U2636 (N_2636,N_2282,N_2243);
and U2637 (N_2637,N_2450,N_2303);
xor U2638 (N_2638,N_2181,N_2404);
nor U2639 (N_2639,N_2028,N_2056);
or U2640 (N_2640,N_2255,N_2361);
nor U2641 (N_2641,N_2046,N_2193);
and U2642 (N_2642,N_2183,N_2117);
nand U2643 (N_2643,N_2014,N_2154);
and U2644 (N_2644,N_2109,N_2275);
nor U2645 (N_2645,N_2494,N_2347);
or U2646 (N_2646,N_2151,N_2163);
and U2647 (N_2647,N_2421,N_2237);
or U2648 (N_2648,N_2208,N_2085);
and U2649 (N_2649,N_2298,N_2152);
nand U2650 (N_2650,N_2429,N_2190);
nor U2651 (N_2651,N_2254,N_2388);
nand U2652 (N_2652,N_2221,N_2273);
and U2653 (N_2653,N_2288,N_2423);
or U2654 (N_2654,N_2355,N_2175);
nand U2655 (N_2655,N_2383,N_2392);
nor U2656 (N_2656,N_2072,N_2301);
or U2657 (N_2657,N_2230,N_2132);
nor U2658 (N_2658,N_2302,N_2395);
nor U2659 (N_2659,N_2088,N_2136);
nor U2660 (N_2660,N_2191,N_2335);
and U2661 (N_2661,N_2212,N_2098);
or U2662 (N_2662,N_2180,N_2231);
nor U2663 (N_2663,N_2267,N_2186);
nor U2664 (N_2664,N_2270,N_2480);
or U2665 (N_2665,N_2393,N_2465);
nand U2666 (N_2666,N_2252,N_2241);
and U2667 (N_2667,N_2315,N_2113);
nand U2668 (N_2668,N_2412,N_2472);
and U2669 (N_2669,N_2262,N_2149);
nand U2670 (N_2670,N_2195,N_2158);
nor U2671 (N_2671,N_2219,N_2482);
and U2672 (N_2672,N_2205,N_2145);
or U2673 (N_2673,N_2490,N_2276);
nor U2674 (N_2674,N_2312,N_2225);
nand U2675 (N_2675,N_2139,N_2342);
or U2676 (N_2676,N_2192,N_2365);
nand U2677 (N_2677,N_2359,N_2258);
nor U2678 (N_2678,N_2125,N_2346);
nor U2679 (N_2679,N_2294,N_2416);
nand U2680 (N_2680,N_2093,N_2259);
nand U2681 (N_2681,N_2348,N_2161);
or U2682 (N_2682,N_2463,N_2257);
or U2683 (N_2683,N_2444,N_2019);
nor U2684 (N_2684,N_2285,N_2223);
nor U2685 (N_2685,N_2162,N_2287);
nor U2686 (N_2686,N_2083,N_2354);
and U2687 (N_2687,N_2284,N_2058);
nand U2688 (N_2688,N_2187,N_2202);
and U2689 (N_2689,N_2000,N_2224);
or U2690 (N_2690,N_2236,N_2130);
and U2691 (N_2691,N_2026,N_2178);
nand U2692 (N_2692,N_2123,N_2087);
nand U2693 (N_2693,N_2426,N_2073);
nand U2694 (N_2694,N_2371,N_2209);
and U2695 (N_2695,N_2319,N_2297);
nand U2696 (N_2696,N_2133,N_2062);
nand U2697 (N_2697,N_2339,N_2229);
nor U2698 (N_2698,N_2407,N_2337);
nand U2699 (N_2699,N_2380,N_2167);
or U2700 (N_2700,N_2316,N_2077);
or U2701 (N_2701,N_2452,N_2263);
or U2702 (N_2702,N_2170,N_2157);
and U2703 (N_2703,N_2055,N_2009);
nand U2704 (N_2704,N_2493,N_2089);
nand U2705 (N_2705,N_2340,N_2438);
and U2706 (N_2706,N_2443,N_2373);
and U2707 (N_2707,N_2447,N_2203);
nand U2708 (N_2708,N_2144,N_2143);
nor U2709 (N_2709,N_2308,N_2199);
nor U2710 (N_2710,N_2104,N_2128);
nor U2711 (N_2711,N_2435,N_2394);
or U2712 (N_2712,N_2216,N_2156);
nor U2713 (N_2713,N_2448,N_2097);
or U2714 (N_2714,N_2439,N_2027);
nand U2715 (N_2715,N_2159,N_2281);
nand U2716 (N_2716,N_2358,N_2485);
and U2717 (N_2717,N_2048,N_2290);
nand U2718 (N_2718,N_2362,N_2106);
nor U2719 (N_2719,N_2357,N_2351);
nor U2720 (N_2720,N_2378,N_2188);
nor U2721 (N_2721,N_2431,N_2310);
and U2722 (N_2722,N_2155,N_2424);
and U2723 (N_2723,N_2094,N_2313);
nor U2724 (N_2724,N_2377,N_2108);
or U2725 (N_2725,N_2356,N_2007);
nand U2726 (N_2726,N_2126,N_2398);
and U2727 (N_2727,N_2122,N_2390);
nand U2728 (N_2728,N_2441,N_2304);
nand U2729 (N_2729,N_2460,N_2470);
nand U2730 (N_2730,N_2411,N_2375);
nand U2731 (N_2731,N_2427,N_2053);
or U2732 (N_2732,N_2038,N_2049);
nand U2733 (N_2733,N_2330,N_2057);
nor U2734 (N_2734,N_2484,N_2331);
and U2735 (N_2735,N_2370,N_2419);
and U2736 (N_2736,N_2119,N_2446);
and U2737 (N_2737,N_2110,N_2385);
or U2738 (N_2738,N_2327,N_2440);
nor U2739 (N_2739,N_2369,N_2467);
and U2740 (N_2740,N_2473,N_2141);
nor U2741 (N_2741,N_2215,N_2366);
nand U2742 (N_2742,N_2397,N_2174);
nand U2743 (N_2743,N_2179,N_2096);
nor U2744 (N_2744,N_2299,N_2422);
or U2745 (N_2745,N_2279,N_2451);
nand U2746 (N_2746,N_2033,N_2400);
nand U2747 (N_2747,N_2468,N_2498);
or U2748 (N_2748,N_2492,N_2176);
and U2749 (N_2749,N_2329,N_2379);
nand U2750 (N_2750,N_2060,N_2305);
or U2751 (N_2751,N_2303,N_2061);
or U2752 (N_2752,N_2298,N_2248);
and U2753 (N_2753,N_2041,N_2182);
and U2754 (N_2754,N_2236,N_2021);
xor U2755 (N_2755,N_2128,N_2099);
nor U2756 (N_2756,N_2350,N_2495);
or U2757 (N_2757,N_2169,N_2056);
nand U2758 (N_2758,N_2496,N_2039);
nor U2759 (N_2759,N_2262,N_2157);
nor U2760 (N_2760,N_2192,N_2487);
and U2761 (N_2761,N_2463,N_2184);
nor U2762 (N_2762,N_2212,N_2221);
and U2763 (N_2763,N_2301,N_2052);
and U2764 (N_2764,N_2080,N_2174);
nor U2765 (N_2765,N_2222,N_2056);
nand U2766 (N_2766,N_2061,N_2070);
nor U2767 (N_2767,N_2354,N_2183);
or U2768 (N_2768,N_2085,N_2334);
nor U2769 (N_2769,N_2111,N_2037);
nand U2770 (N_2770,N_2375,N_2356);
nand U2771 (N_2771,N_2202,N_2497);
and U2772 (N_2772,N_2240,N_2151);
nor U2773 (N_2773,N_2172,N_2123);
or U2774 (N_2774,N_2029,N_2051);
nand U2775 (N_2775,N_2211,N_2330);
nor U2776 (N_2776,N_2499,N_2097);
nor U2777 (N_2777,N_2492,N_2140);
or U2778 (N_2778,N_2206,N_2455);
nand U2779 (N_2779,N_2199,N_2158);
and U2780 (N_2780,N_2359,N_2270);
nand U2781 (N_2781,N_2301,N_2212);
nor U2782 (N_2782,N_2276,N_2229);
nor U2783 (N_2783,N_2056,N_2355);
and U2784 (N_2784,N_2186,N_2361);
nor U2785 (N_2785,N_2252,N_2300);
nand U2786 (N_2786,N_2129,N_2211);
and U2787 (N_2787,N_2337,N_2464);
or U2788 (N_2788,N_2175,N_2104);
or U2789 (N_2789,N_2078,N_2154);
or U2790 (N_2790,N_2215,N_2290);
and U2791 (N_2791,N_2124,N_2259);
or U2792 (N_2792,N_2374,N_2482);
nand U2793 (N_2793,N_2218,N_2095);
or U2794 (N_2794,N_2152,N_2025);
or U2795 (N_2795,N_2026,N_2034);
and U2796 (N_2796,N_2049,N_2417);
or U2797 (N_2797,N_2488,N_2412);
nand U2798 (N_2798,N_2397,N_2186);
nor U2799 (N_2799,N_2033,N_2433);
or U2800 (N_2800,N_2324,N_2225);
or U2801 (N_2801,N_2311,N_2280);
and U2802 (N_2802,N_2300,N_2199);
nand U2803 (N_2803,N_2304,N_2011);
nor U2804 (N_2804,N_2078,N_2124);
or U2805 (N_2805,N_2229,N_2343);
nor U2806 (N_2806,N_2303,N_2309);
nand U2807 (N_2807,N_2380,N_2106);
xnor U2808 (N_2808,N_2018,N_2205);
nor U2809 (N_2809,N_2256,N_2015);
nand U2810 (N_2810,N_2354,N_2391);
nand U2811 (N_2811,N_2295,N_2373);
or U2812 (N_2812,N_2487,N_2017);
and U2813 (N_2813,N_2482,N_2081);
and U2814 (N_2814,N_2023,N_2077);
nor U2815 (N_2815,N_2461,N_2065);
or U2816 (N_2816,N_2272,N_2478);
and U2817 (N_2817,N_2039,N_2260);
nor U2818 (N_2818,N_2036,N_2317);
nor U2819 (N_2819,N_2028,N_2329);
or U2820 (N_2820,N_2135,N_2099);
and U2821 (N_2821,N_2439,N_2056);
or U2822 (N_2822,N_2080,N_2401);
nor U2823 (N_2823,N_2075,N_2446);
or U2824 (N_2824,N_2121,N_2175);
nor U2825 (N_2825,N_2296,N_2120);
or U2826 (N_2826,N_2278,N_2049);
nor U2827 (N_2827,N_2265,N_2485);
nor U2828 (N_2828,N_2100,N_2318);
and U2829 (N_2829,N_2232,N_2156);
or U2830 (N_2830,N_2059,N_2497);
nand U2831 (N_2831,N_2360,N_2078);
nand U2832 (N_2832,N_2187,N_2244);
nand U2833 (N_2833,N_2236,N_2304);
or U2834 (N_2834,N_2208,N_2167);
nor U2835 (N_2835,N_2373,N_2422);
and U2836 (N_2836,N_2136,N_2035);
nand U2837 (N_2837,N_2278,N_2286);
nor U2838 (N_2838,N_2425,N_2442);
nor U2839 (N_2839,N_2413,N_2068);
or U2840 (N_2840,N_2424,N_2416);
nor U2841 (N_2841,N_2403,N_2365);
nand U2842 (N_2842,N_2169,N_2298);
nor U2843 (N_2843,N_2280,N_2467);
nand U2844 (N_2844,N_2028,N_2352);
nand U2845 (N_2845,N_2206,N_2332);
nor U2846 (N_2846,N_2346,N_2399);
and U2847 (N_2847,N_2348,N_2458);
nand U2848 (N_2848,N_2053,N_2166);
and U2849 (N_2849,N_2306,N_2237);
nand U2850 (N_2850,N_2300,N_2482);
nand U2851 (N_2851,N_2204,N_2057);
nor U2852 (N_2852,N_2297,N_2443);
or U2853 (N_2853,N_2201,N_2061);
nand U2854 (N_2854,N_2068,N_2009);
nand U2855 (N_2855,N_2154,N_2275);
or U2856 (N_2856,N_2006,N_2290);
nand U2857 (N_2857,N_2469,N_2189);
nand U2858 (N_2858,N_2010,N_2106);
nor U2859 (N_2859,N_2441,N_2178);
nand U2860 (N_2860,N_2450,N_2017);
nor U2861 (N_2861,N_2362,N_2363);
and U2862 (N_2862,N_2271,N_2153);
nor U2863 (N_2863,N_2269,N_2176);
and U2864 (N_2864,N_2340,N_2482);
nand U2865 (N_2865,N_2451,N_2215);
nor U2866 (N_2866,N_2122,N_2029);
and U2867 (N_2867,N_2051,N_2140);
or U2868 (N_2868,N_2196,N_2050);
and U2869 (N_2869,N_2039,N_2073);
nand U2870 (N_2870,N_2492,N_2370);
nand U2871 (N_2871,N_2210,N_2443);
or U2872 (N_2872,N_2401,N_2285);
nand U2873 (N_2873,N_2013,N_2373);
nand U2874 (N_2874,N_2161,N_2261);
and U2875 (N_2875,N_2451,N_2124);
nand U2876 (N_2876,N_2439,N_2018);
or U2877 (N_2877,N_2352,N_2372);
or U2878 (N_2878,N_2405,N_2138);
nor U2879 (N_2879,N_2270,N_2353);
and U2880 (N_2880,N_2043,N_2214);
nand U2881 (N_2881,N_2152,N_2392);
nand U2882 (N_2882,N_2288,N_2165);
and U2883 (N_2883,N_2429,N_2408);
or U2884 (N_2884,N_2413,N_2133);
and U2885 (N_2885,N_2185,N_2138);
nand U2886 (N_2886,N_2129,N_2017);
nor U2887 (N_2887,N_2207,N_2239);
nor U2888 (N_2888,N_2356,N_2222);
and U2889 (N_2889,N_2345,N_2206);
or U2890 (N_2890,N_2285,N_2179);
or U2891 (N_2891,N_2249,N_2476);
and U2892 (N_2892,N_2445,N_2455);
or U2893 (N_2893,N_2395,N_2287);
nand U2894 (N_2894,N_2374,N_2331);
nor U2895 (N_2895,N_2462,N_2281);
nand U2896 (N_2896,N_2264,N_2084);
nand U2897 (N_2897,N_2316,N_2355);
and U2898 (N_2898,N_2216,N_2320);
nor U2899 (N_2899,N_2394,N_2127);
or U2900 (N_2900,N_2175,N_2243);
or U2901 (N_2901,N_2234,N_2201);
or U2902 (N_2902,N_2382,N_2142);
or U2903 (N_2903,N_2409,N_2364);
nand U2904 (N_2904,N_2379,N_2333);
or U2905 (N_2905,N_2419,N_2174);
or U2906 (N_2906,N_2386,N_2243);
or U2907 (N_2907,N_2448,N_2397);
nand U2908 (N_2908,N_2382,N_2238);
nor U2909 (N_2909,N_2473,N_2016);
nor U2910 (N_2910,N_2374,N_2439);
nand U2911 (N_2911,N_2233,N_2248);
and U2912 (N_2912,N_2195,N_2363);
and U2913 (N_2913,N_2041,N_2123);
nand U2914 (N_2914,N_2434,N_2256);
or U2915 (N_2915,N_2375,N_2431);
or U2916 (N_2916,N_2314,N_2464);
nor U2917 (N_2917,N_2483,N_2463);
nor U2918 (N_2918,N_2102,N_2106);
and U2919 (N_2919,N_2321,N_2411);
nor U2920 (N_2920,N_2176,N_2488);
nor U2921 (N_2921,N_2221,N_2301);
nor U2922 (N_2922,N_2392,N_2220);
nand U2923 (N_2923,N_2130,N_2061);
nand U2924 (N_2924,N_2012,N_2340);
or U2925 (N_2925,N_2409,N_2293);
and U2926 (N_2926,N_2452,N_2398);
or U2927 (N_2927,N_2143,N_2389);
or U2928 (N_2928,N_2374,N_2345);
and U2929 (N_2929,N_2137,N_2263);
nor U2930 (N_2930,N_2296,N_2013);
and U2931 (N_2931,N_2195,N_2367);
or U2932 (N_2932,N_2376,N_2192);
and U2933 (N_2933,N_2353,N_2446);
nor U2934 (N_2934,N_2400,N_2389);
nand U2935 (N_2935,N_2105,N_2170);
nand U2936 (N_2936,N_2085,N_2445);
nand U2937 (N_2937,N_2121,N_2393);
nand U2938 (N_2938,N_2358,N_2235);
nand U2939 (N_2939,N_2090,N_2478);
or U2940 (N_2940,N_2000,N_2087);
or U2941 (N_2941,N_2417,N_2234);
nor U2942 (N_2942,N_2127,N_2099);
nor U2943 (N_2943,N_2308,N_2317);
nor U2944 (N_2944,N_2032,N_2010);
or U2945 (N_2945,N_2052,N_2109);
and U2946 (N_2946,N_2364,N_2352);
or U2947 (N_2947,N_2462,N_2447);
xnor U2948 (N_2948,N_2141,N_2153);
nand U2949 (N_2949,N_2157,N_2315);
or U2950 (N_2950,N_2139,N_2152);
or U2951 (N_2951,N_2088,N_2216);
or U2952 (N_2952,N_2488,N_2172);
and U2953 (N_2953,N_2402,N_2390);
and U2954 (N_2954,N_2102,N_2340);
nand U2955 (N_2955,N_2454,N_2140);
or U2956 (N_2956,N_2297,N_2379);
and U2957 (N_2957,N_2099,N_2195);
or U2958 (N_2958,N_2279,N_2447);
nand U2959 (N_2959,N_2184,N_2170);
nand U2960 (N_2960,N_2295,N_2288);
and U2961 (N_2961,N_2381,N_2404);
or U2962 (N_2962,N_2155,N_2034);
nor U2963 (N_2963,N_2384,N_2274);
and U2964 (N_2964,N_2420,N_2466);
nand U2965 (N_2965,N_2481,N_2354);
and U2966 (N_2966,N_2444,N_2377);
nand U2967 (N_2967,N_2468,N_2110);
nor U2968 (N_2968,N_2008,N_2382);
nor U2969 (N_2969,N_2400,N_2017);
and U2970 (N_2970,N_2377,N_2389);
xnor U2971 (N_2971,N_2022,N_2442);
nand U2972 (N_2972,N_2443,N_2290);
and U2973 (N_2973,N_2277,N_2314);
and U2974 (N_2974,N_2451,N_2449);
or U2975 (N_2975,N_2460,N_2329);
nor U2976 (N_2976,N_2010,N_2407);
or U2977 (N_2977,N_2333,N_2401);
nor U2978 (N_2978,N_2274,N_2044);
nand U2979 (N_2979,N_2448,N_2055);
and U2980 (N_2980,N_2379,N_2041);
nand U2981 (N_2981,N_2231,N_2401);
nor U2982 (N_2982,N_2344,N_2293);
nor U2983 (N_2983,N_2181,N_2207);
or U2984 (N_2984,N_2211,N_2424);
or U2985 (N_2985,N_2481,N_2476);
or U2986 (N_2986,N_2179,N_2350);
nor U2987 (N_2987,N_2030,N_2115);
nand U2988 (N_2988,N_2315,N_2419);
or U2989 (N_2989,N_2024,N_2130);
or U2990 (N_2990,N_2370,N_2438);
nand U2991 (N_2991,N_2160,N_2104);
nor U2992 (N_2992,N_2376,N_2411);
or U2993 (N_2993,N_2401,N_2102);
or U2994 (N_2994,N_2293,N_2458);
or U2995 (N_2995,N_2484,N_2294);
or U2996 (N_2996,N_2021,N_2149);
nand U2997 (N_2997,N_2374,N_2209);
or U2998 (N_2998,N_2441,N_2255);
nor U2999 (N_2999,N_2088,N_2424);
or U3000 (N_3000,N_2904,N_2530);
or U3001 (N_3001,N_2880,N_2714);
and U3002 (N_3002,N_2973,N_2785);
and U3003 (N_3003,N_2589,N_2801);
or U3004 (N_3004,N_2662,N_2734);
and U3005 (N_3005,N_2501,N_2542);
and U3006 (N_3006,N_2572,N_2675);
nor U3007 (N_3007,N_2590,N_2868);
nand U3008 (N_3008,N_2964,N_2978);
or U3009 (N_3009,N_2751,N_2667);
nor U3010 (N_3010,N_2933,N_2583);
nor U3011 (N_3011,N_2552,N_2676);
nor U3012 (N_3012,N_2762,N_2640);
xor U3013 (N_3013,N_2943,N_2780);
nor U3014 (N_3014,N_2889,N_2900);
nand U3015 (N_3015,N_2961,N_2723);
or U3016 (N_3016,N_2617,N_2733);
nor U3017 (N_3017,N_2525,N_2775);
nand U3018 (N_3018,N_2674,N_2659);
nand U3019 (N_3019,N_2963,N_2596);
or U3020 (N_3020,N_2953,N_2895);
nand U3021 (N_3021,N_2571,N_2870);
nand U3022 (N_3022,N_2894,N_2577);
or U3023 (N_3023,N_2586,N_2557);
nand U3024 (N_3024,N_2917,N_2546);
or U3025 (N_3025,N_2587,N_2950);
nand U3026 (N_3026,N_2830,N_2720);
nor U3027 (N_3027,N_2710,N_2845);
and U3028 (N_3028,N_2837,N_2938);
and U3029 (N_3029,N_2912,N_2665);
nand U3030 (N_3030,N_2823,N_2891);
or U3031 (N_3031,N_2739,N_2520);
or U3032 (N_3032,N_2568,N_2502);
nand U3033 (N_3033,N_2813,N_2570);
nor U3034 (N_3034,N_2805,N_2609);
nor U3035 (N_3035,N_2545,N_2729);
and U3036 (N_3036,N_2914,N_2614);
nor U3037 (N_3037,N_2716,N_2819);
nand U3038 (N_3038,N_2913,N_2608);
nand U3039 (N_3039,N_2585,N_2555);
or U3040 (N_3040,N_2976,N_2712);
nand U3041 (N_3041,N_2782,N_2772);
nand U3042 (N_3042,N_2576,N_2503);
and U3043 (N_3043,N_2646,N_2928);
nand U3044 (N_3044,N_2983,N_2745);
or U3045 (N_3045,N_2599,N_2853);
and U3046 (N_3046,N_2936,N_2701);
or U3047 (N_3047,N_2875,N_2907);
or U3048 (N_3048,N_2550,N_2651);
nor U3049 (N_3049,N_2768,N_2954);
xor U3050 (N_3050,N_2524,N_2728);
or U3051 (N_3051,N_2696,N_2629);
or U3052 (N_3052,N_2737,N_2746);
nand U3053 (N_3053,N_2564,N_2942);
nand U3054 (N_3054,N_2937,N_2831);
or U3055 (N_3055,N_2932,N_2673);
and U3056 (N_3056,N_2538,N_2803);
nand U3057 (N_3057,N_2818,N_2686);
nand U3058 (N_3058,N_2621,N_2529);
nand U3059 (N_3059,N_2774,N_2725);
xor U3060 (N_3060,N_2666,N_2984);
and U3061 (N_3061,N_2994,N_2533);
nor U3062 (N_3062,N_2579,N_2602);
and U3063 (N_3063,N_2692,N_2977);
or U3064 (N_3064,N_2652,N_2876);
xor U3065 (N_3065,N_2862,N_2829);
nand U3066 (N_3066,N_2613,N_2776);
and U3067 (N_3067,N_2540,N_2559);
and U3068 (N_3068,N_2655,N_2697);
nand U3069 (N_3069,N_2885,N_2832);
nand U3070 (N_3070,N_2606,N_2625);
nor U3071 (N_3071,N_2680,N_2612);
and U3072 (N_3072,N_2563,N_2883);
nand U3073 (N_3073,N_2882,N_2653);
nand U3074 (N_3074,N_2523,N_2987);
nor U3075 (N_3075,N_2826,N_2506);
and U3076 (N_3076,N_2906,N_2787);
and U3077 (N_3077,N_2873,N_2635);
or U3078 (N_3078,N_2974,N_2702);
nor U3079 (N_3079,N_2514,N_2750);
xor U3080 (N_3080,N_2593,N_2962);
nand U3081 (N_3081,N_2634,N_2945);
nand U3082 (N_3082,N_2763,N_2929);
or U3083 (N_3083,N_2627,N_2537);
nand U3084 (N_3084,N_2700,N_2838);
and U3085 (N_3085,N_2584,N_2531);
and U3086 (N_3086,N_2628,N_2784);
nor U3087 (N_3087,N_2508,N_2753);
and U3088 (N_3088,N_2821,N_2660);
or U3089 (N_3089,N_2671,N_2939);
nand U3090 (N_3090,N_2802,N_2810);
or U3091 (N_3091,N_2910,N_2594);
and U3092 (N_3092,N_2742,N_2850);
nor U3093 (N_3093,N_2988,N_2598);
or U3094 (N_3094,N_2835,N_2521);
or U3095 (N_3095,N_2715,N_2681);
and U3096 (N_3096,N_2844,N_2636);
and U3097 (N_3097,N_2897,N_2949);
xnor U3098 (N_3098,N_2709,N_2558);
nand U3099 (N_3099,N_2777,N_2547);
nor U3100 (N_3100,N_2565,N_2694);
and U3101 (N_3101,N_2597,N_2812);
and U3102 (N_3102,N_2619,N_2638);
or U3103 (N_3103,N_2717,N_2690);
nand U3104 (N_3104,N_2708,N_2946);
nand U3105 (N_3105,N_2624,N_2543);
or U3106 (N_3106,N_2935,N_2644);
and U3107 (N_3107,N_2718,N_2797);
or U3108 (N_3108,N_2998,N_2944);
nand U3109 (N_3109,N_2903,N_2981);
nand U3110 (N_3110,N_2730,N_2857);
nand U3111 (N_3111,N_2893,N_2990);
or U3112 (N_3112,N_2767,N_2670);
nor U3113 (N_3113,N_2901,N_2811);
nor U3114 (N_3114,N_2504,N_2643);
nor U3115 (N_3115,N_2847,N_2573);
and U3116 (N_3116,N_2689,N_2687);
and U3117 (N_3117,N_2663,N_2796);
and U3118 (N_3118,N_2748,N_2856);
nor U3119 (N_3119,N_2808,N_2877);
nor U3120 (N_3120,N_2795,N_2664);
nor U3121 (N_3121,N_2757,N_2927);
or U3122 (N_3122,N_2726,N_2707);
nor U3123 (N_3123,N_2685,N_2760);
nor U3124 (N_3124,N_2711,N_2781);
nor U3125 (N_3125,N_2560,N_2959);
nor U3126 (N_3126,N_2920,N_2649);
nand U3127 (N_3127,N_2874,N_2836);
or U3128 (N_3128,N_2869,N_2863);
nand U3129 (N_3129,N_2713,N_2861);
or U3130 (N_3130,N_2582,N_2526);
and U3131 (N_3131,N_2616,N_2769);
nand U3132 (N_3132,N_2919,N_2648);
nand U3133 (N_3133,N_2980,N_2601);
or U3134 (N_3134,N_2672,N_2815);
nand U3135 (N_3135,N_2500,N_2905);
nor U3136 (N_3136,N_2682,N_2872);
nor U3137 (N_3137,N_2691,N_2807);
or U3138 (N_3138,N_2605,N_2522);
nor U3139 (N_3139,N_2908,N_2548);
nor U3140 (N_3140,N_2747,N_2758);
and U3141 (N_3141,N_2592,N_2699);
nand U3142 (N_3142,N_2567,N_2968);
or U3143 (N_3143,N_2724,N_2637);
nand U3144 (N_3144,N_2820,N_2541);
nand U3145 (N_3145,N_2886,N_2771);
or U3146 (N_3146,N_2551,N_2595);
nand U3147 (N_3147,N_2852,N_2575);
nand U3148 (N_3148,N_2822,N_2827);
nor U3149 (N_3149,N_2654,N_2607);
nand U3150 (N_3150,N_2957,N_2925);
nor U3151 (N_3151,N_2562,N_2817);
nand U3152 (N_3152,N_2930,N_2722);
or U3153 (N_3153,N_2956,N_2966);
nor U3154 (N_3154,N_2790,N_2678);
and U3155 (N_3155,N_2727,N_2825);
or U3156 (N_3156,N_2794,N_2849);
or U3157 (N_3157,N_2955,N_2512);
or U3158 (N_3158,N_2855,N_2622);
or U3159 (N_3159,N_2986,N_2510);
nand U3160 (N_3160,N_2765,N_2693);
nor U3161 (N_3161,N_2911,N_2798);
and U3162 (N_3162,N_2834,N_2631);
or U3163 (N_3163,N_2866,N_2871);
xor U3164 (N_3164,N_2752,N_2705);
and U3165 (N_3165,N_2890,N_2887);
or U3166 (N_3166,N_2704,N_2915);
nor U3167 (N_3167,N_2735,N_2985);
nor U3168 (N_3168,N_2941,N_2668);
nand U3169 (N_3169,N_2528,N_2878);
nor U3170 (N_3170,N_2683,N_2719);
nand U3171 (N_3171,N_2618,N_2744);
nor U3172 (N_3172,N_2574,N_2809);
or U3173 (N_3173,N_2641,N_2569);
xor U3174 (N_3174,N_2766,N_2773);
nand U3175 (N_3175,N_2741,N_2695);
nand U3176 (N_3176,N_2864,N_2884);
nor U3177 (N_3177,N_2656,N_2738);
or U3178 (N_3178,N_2623,N_2833);
nand U3179 (N_3179,N_2519,N_2934);
or U3180 (N_3180,N_2677,N_2881);
or U3181 (N_3181,N_2867,N_2517);
or U3182 (N_3182,N_2839,N_2556);
or U3183 (N_3183,N_2604,N_2539);
nand U3184 (N_3184,N_2860,N_2969);
or U3185 (N_3185,N_2951,N_2661);
and U3186 (N_3186,N_2967,N_2918);
and U3187 (N_3187,N_2923,N_2620);
or U3188 (N_3188,N_2650,N_2764);
and U3189 (N_3189,N_2979,N_2865);
and U3190 (N_3190,N_2997,N_2515);
and U3191 (N_3191,N_2926,N_2846);
nand U3192 (N_3192,N_2633,N_2898);
and U3193 (N_3193,N_2561,N_2982);
nand U3194 (N_3194,N_2960,N_2679);
and U3195 (N_3195,N_2858,N_2828);
or U3196 (N_3196,N_2658,N_2721);
or U3197 (N_3197,N_2580,N_2732);
or U3198 (N_3198,N_2511,N_2786);
or U3199 (N_3199,N_2761,N_2824);
or U3200 (N_3200,N_2793,N_2749);
and U3201 (N_3201,N_2971,N_2581);
nor U3202 (N_3202,N_2975,N_2842);
nand U3203 (N_3203,N_2804,N_2645);
or U3204 (N_3204,N_2783,N_2922);
nand U3205 (N_3205,N_2989,N_2947);
and U3206 (N_3206,N_2684,N_2999);
or U3207 (N_3207,N_2603,N_2909);
xor U3208 (N_3208,N_2516,N_2892);
or U3209 (N_3209,N_2518,N_2657);
nand U3210 (N_3210,N_2996,N_2791);
xor U3211 (N_3211,N_2535,N_2743);
and U3212 (N_3212,N_2896,N_2806);
nand U3213 (N_3213,N_2532,N_2779);
nor U3214 (N_3214,N_2840,N_2505);
nand U3215 (N_3215,N_2706,N_2848);
nor U3216 (N_3216,N_2755,N_2799);
and U3217 (N_3217,N_2843,N_2993);
and U3218 (N_3218,N_2940,N_2626);
and U3219 (N_3219,N_2600,N_2698);
and U3220 (N_3220,N_2591,N_2688);
and U3221 (N_3221,N_2736,N_2800);
nand U3222 (N_3222,N_2754,N_2924);
nand U3223 (N_3223,N_2647,N_2854);
and U3224 (N_3224,N_2995,N_2992);
nor U3225 (N_3225,N_2788,N_2615);
or U3226 (N_3226,N_2888,N_2527);
nand U3227 (N_3227,N_2916,N_2879);
and U3228 (N_3228,N_2958,N_2566);
or U3229 (N_3229,N_2544,N_2534);
nand U3230 (N_3230,N_2740,N_2816);
nand U3231 (N_3231,N_2814,N_2789);
nor U3232 (N_3232,N_2899,N_2902);
nand U3233 (N_3233,N_2952,N_2770);
or U3234 (N_3234,N_2970,N_2509);
nor U3235 (N_3235,N_2507,N_2610);
nor U3236 (N_3236,N_2921,N_2972);
nor U3237 (N_3237,N_2553,N_2731);
nor U3238 (N_3238,N_2588,N_2536);
nor U3239 (N_3239,N_2554,N_2931);
and U3240 (N_3240,N_2792,N_2549);
nor U3241 (N_3241,N_2578,N_2639);
or U3242 (N_3242,N_2756,N_2642);
and U3243 (N_3243,N_2841,N_2630);
or U3244 (N_3244,N_2669,N_2991);
or U3245 (N_3245,N_2859,N_2703);
nand U3246 (N_3246,N_2851,N_2778);
and U3247 (N_3247,N_2965,N_2632);
and U3248 (N_3248,N_2948,N_2611);
nand U3249 (N_3249,N_2513,N_2759);
and U3250 (N_3250,N_2979,N_2975);
and U3251 (N_3251,N_2897,N_2676);
or U3252 (N_3252,N_2524,N_2689);
or U3253 (N_3253,N_2568,N_2604);
or U3254 (N_3254,N_2780,N_2545);
nor U3255 (N_3255,N_2776,N_2553);
nand U3256 (N_3256,N_2560,N_2955);
or U3257 (N_3257,N_2940,N_2523);
nand U3258 (N_3258,N_2879,N_2919);
nor U3259 (N_3259,N_2528,N_2607);
nor U3260 (N_3260,N_2526,N_2928);
nand U3261 (N_3261,N_2658,N_2605);
or U3262 (N_3262,N_2884,N_2557);
or U3263 (N_3263,N_2837,N_2816);
nand U3264 (N_3264,N_2734,N_2998);
nor U3265 (N_3265,N_2524,N_2870);
and U3266 (N_3266,N_2555,N_2997);
and U3267 (N_3267,N_2596,N_2663);
or U3268 (N_3268,N_2872,N_2800);
nand U3269 (N_3269,N_2828,N_2582);
and U3270 (N_3270,N_2534,N_2555);
nand U3271 (N_3271,N_2930,N_2846);
or U3272 (N_3272,N_2830,N_2939);
nor U3273 (N_3273,N_2675,N_2938);
and U3274 (N_3274,N_2860,N_2880);
nand U3275 (N_3275,N_2671,N_2623);
and U3276 (N_3276,N_2746,N_2515);
and U3277 (N_3277,N_2814,N_2684);
or U3278 (N_3278,N_2721,N_2538);
nand U3279 (N_3279,N_2660,N_2699);
nand U3280 (N_3280,N_2982,N_2979);
and U3281 (N_3281,N_2599,N_2716);
and U3282 (N_3282,N_2513,N_2935);
nor U3283 (N_3283,N_2575,N_2817);
and U3284 (N_3284,N_2640,N_2596);
and U3285 (N_3285,N_2681,N_2892);
and U3286 (N_3286,N_2971,N_2765);
or U3287 (N_3287,N_2592,N_2600);
nor U3288 (N_3288,N_2794,N_2619);
nor U3289 (N_3289,N_2533,N_2741);
nand U3290 (N_3290,N_2637,N_2869);
nand U3291 (N_3291,N_2993,N_2938);
and U3292 (N_3292,N_2930,N_2781);
or U3293 (N_3293,N_2764,N_2748);
and U3294 (N_3294,N_2798,N_2542);
or U3295 (N_3295,N_2957,N_2840);
nand U3296 (N_3296,N_2653,N_2870);
and U3297 (N_3297,N_2833,N_2606);
or U3298 (N_3298,N_2944,N_2788);
nand U3299 (N_3299,N_2552,N_2791);
nor U3300 (N_3300,N_2872,N_2975);
and U3301 (N_3301,N_2845,N_2794);
and U3302 (N_3302,N_2600,N_2718);
or U3303 (N_3303,N_2502,N_2836);
or U3304 (N_3304,N_2699,N_2770);
nor U3305 (N_3305,N_2727,N_2737);
nor U3306 (N_3306,N_2740,N_2990);
or U3307 (N_3307,N_2915,N_2555);
nand U3308 (N_3308,N_2513,N_2604);
nand U3309 (N_3309,N_2672,N_2505);
and U3310 (N_3310,N_2588,N_2655);
nand U3311 (N_3311,N_2903,N_2840);
nand U3312 (N_3312,N_2807,N_2846);
nor U3313 (N_3313,N_2801,N_2510);
and U3314 (N_3314,N_2919,N_2813);
nand U3315 (N_3315,N_2775,N_2663);
or U3316 (N_3316,N_2758,N_2880);
or U3317 (N_3317,N_2994,N_2848);
or U3318 (N_3318,N_2520,N_2991);
or U3319 (N_3319,N_2730,N_2874);
nand U3320 (N_3320,N_2666,N_2829);
or U3321 (N_3321,N_2736,N_2940);
nand U3322 (N_3322,N_2832,N_2557);
nor U3323 (N_3323,N_2679,N_2589);
and U3324 (N_3324,N_2657,N_2606);
nand U3325 (N_3325,N_2711,N_2570);
and U3326 (N_3326,N_2937,N_2617);
and U3327 (N_3327,N_2648,N_2991);
and U3328 (N_3328,N_2554,N_2504);
nor U3329 (N_3329,N_2535,N_2745);
or U3330 (N_3330,N_2636,N_2627);
nor U3331 (N_3331,N_2897,N_2940);
or U3332 (N_3332,N_2720,N_2834);
nand U3333 (N_3333,N_2525,N_2723);
xnor U3334 (N_3334,N_2715,N_2669);
or U3335 (N_3335,N_2730,N_2893);
and U3336 (N_3336,N_2599,N_2997);
nand U3337 (N_3337,N_2825,N_2552);
nand U3338 (N_3338,N_2979,N_2873);
and U3339 (N_3339,N_2660,N_2854);
nand U3340 (N_3340,N_2724,N_2879);
nand U3341 (N_3341,N_2860,N_2907);
nand U3342 (N_3342,N_2893,N_2957);
or U3343 (N_3343,N_2961,N_2665);
and U3344 (N_3344,N_2580,N_2628);
or U3345 (N_3345,N_2794,N_2966);
and U3346 (N_3346,N_2564,N_2631);
nand U3347 (N_3347,N_2695,N_2609);
nor U3348 (N_3348,N_2945,N_2978);
and U3349 (N_3349,N_2578,N_2697);
and U3350 (N_3350,N_2691,N_2616);
nor U3351 (N_3351,N_2774,N_2539);
or U3352 (N_3352,N_2838,N_2706);
nand U3353 (N_3353,N_2600,N_2758);
nor U3354 (N_3354,N_2931,N_2539);
nand U3355 (N_3355,N_2960,N_2541);
nor U3356 (N_3356,N_2644,N_2584);
and U3357 (N_3357,N_2684,N_2652);
nand U3358 (N_3358,N_2616,N_2554);
or U3359 (N_3359,N_2691,N_2893);
nor U3360 (N_3360,N_2558,N_2618);
and U3361 (N_3361,N_2658,N_2977);
nor U3362 (N_3362,N_2816,N_2726);
or U3363 (N_3363,N_2503,N_2668);
nor U3364 (N_3364,N_2929,N_2765);
nor U3365 (N_3365,N_2747,N_2845);
or U3366 (N_3366,N_2964,N_2624);
or U3367 (N_3367,N_2805,N_2813);
and U3368 (N_3368,N_2647,N_2974);
nand U3369 (N_3369,N_2789,N_2934);
or U3370 (N_3370,N_2780,N_2591);
nor U3371 (N_3371,N_2603,N_2689);
and U3372 (N_3372,N_2786,N_2785);
and U3373 (N_3373,N_2835,N_2851);
or U3374 (N_3374,N_2663,N_2749);
or U3375 (N_3375,N_2920,N_2509);
nand U3376 (N_3376,N_2521,N_2755);
nand U3377 (N_3377,N_2930,N_2963);
nor U3378 (N_3378,N_2761,N_2748);
nand U3379 (N_3379,N_2838,N_2655);
xnor U3380 (N_3380,N_2601,N_2710);
and U3381 (N_3381,N_2622,N_2632);
nand U3382 (N_3382,N_2725,N_2699);
nor U3383 (N_3383,N_2738,N_2716);
and U3384 (N_3384,N_2618,N_2626);
nand U3385 (N_3385,N_2622,N_2767);
nor U3386 (N_3386,N_2830,N_2649);
nor U3387 (N_3387,N_2721,N_2708);
or U3388 (N_3388,N_2829,N_2585);
and U3389 (N_3389,N_2538,N_2865);
and U3390 (N_3390,N_2969,N_2688);
and U3391 (N_3391,N_2713,N_2707);
and U3392 (N_3392,N_2508,N_2655);
nand U3393 (N_3393,N_2845,N_2851);
nor U3394 (N_3394,N_2865,N_2646);
and U3395 (N_3395,N_2512,N_2501);
nand U3396 (N_3396,N_2685,N_2887);
nor U3397 (N_3397,N_2747,N_2636);
and U3398 (N_3398,N_2589,N_2987);
and U3399 (N_3399,N_2873,N_2720);
and U3400 (N_3400,N_2712,N_2619);
or U3401 (N_3401,N_2798,N_2941);
nand U3402 (N_3402,N_2753,N_2770);
and U3403 (N_3403,N_2676,N_2982);
and U3404 (N_3404,N_2639,N_2767);
nand U3405 (N_3405,N_2854,N_2767);
nand U3406 (N_3406,N_2969,N_2727);
and U3407 (N_3407,N_2804,N_2848);
or U3408 (N_3408,N_2536,N_2781);
xnor U3409 (N_3409,N_2753,N_2754);
nor U3410 (N_3410,N_2590,N_2759);
and U3411 (N_3411,N_2975,N_2905);
nor U3412 (N_3412,N_2679,N_2824);
and U3413 (N_3413,N_2839,N_2626);
or U3414 (N_3414,N_2553,N_2788);
nand U3415 (N_3415,N_2741,N_2870);
nand U3416 (N_3416,N_2704,N_2552);
nor U3417 (N_3417,N_2943,N_2950);
and U3418 (N_3418,N_2694,N_2680);
or U3419 (N_3419,N_2887,N_2782);
nor U3420 (N_3420,N_2551,N_2699);
nand U3421 (N_3421,N_2649,N_2577);
nor U3422 (N_3422,N_2540,N_2877);
nor U3423 (N_3423,N_2687,N_2656);
xnor U3424 (N_3424,N_2589,N_2800);
nor U3425 (N_3425,N_2578,N_2569);
nand U3426 (N_3426,N_2944,N_2818);
nand U3427 (N_3427,N_2786,N_2702);
nand U3428 (N_3428,N_2767,N_2770);
or U3429 (N_3429,N_2957,N_2788);
xor U3430 (N_3430,N_2768,N_2751);
xnor U3431 (N_3431,N_2884,N_2522);
nor U3432 (N_3432,N_2816,N_2685);
and U3433 (N_3433,N_2571,N_2903);
nor U3434 (N_3434,N_2818,N_2559);
or U3435 (N_3435,N_2783,N_2679);
and U3436 (N_3436,N_2694,N_2719);
nor U3437 (N_3437,N_2884,N_2526);
or U3438 (N_3438,N_2994,N_2842);
nor U3439 (N_3439,N_2853,N_2510);
and U3440 (N_3440,N_2788,N_2927);
nand U3441 (N_3441,N_2562,N_2978);
nand U3442 (N_3442,N_2539,N_2737);
or U3443 (N_3443,N_2996,N_2839);
nor U3444 (N_3444,N_2804,N_2577);
nand U3445 (N_3445,N_2625,N_2683);
nor U3446 (N_3446,N_2745,N_2677);
or U3447 (N_3447,N_2586,N_2556);
and U3448 (N_3448,N_2858,N_2718);
nor U3449 (N_3449,N_2643,N_2896);
nand U3450 (N_3450,N_2607,N_2897);
nand U3451 (N_3451,N_2547,N_2900);
nor U3452 (N_3452,N_2923,N_2627);
nand U3453 (N_3453,N_2905,N_2625);
nand U3454 (N_3454,N_2952,N_2766);
nor U3455 (N_3455,N_2825,N_2855);
and U3456 (N_3456,N_2540,N_2547);
nand U3457 (N_3457,N_2683,N_2903);
xor U3458 (N_3458,N_2955,N_2994);
and U3459 (N_3459,N_2881,N_2713);
and U3460 (N_3460,N_2561,N_2792);
nand U3461 (N_3461,N_2794,N_2751);
nand U3462 (N_3462,N_2685,N_2763);
xor U3463 (N_3463,N_2690,N_2698);
nor U3464 (N_3464,N_2565,N_2742);
nor U3465 (N_3465,N_2919,N_2646);
nand U3466 (N_3466,N_2669,N_2898);
nand U3467 (N_3467,N_2643,N_2962);
nor U3468 (N_3468,N_2854,N_2736);
and U3469 (N_3469,N_2988,N_2618);
and U3470 (N_3470,N_2748,N_2901);
and U3471 (N_3471,N_2898,N_2818);
nor U3472 (N_3472,N_2736,N_2898);
and U3473 (N_3473,N_2979,N_2840);
or U3474 (N_3474,N_2557,N_2597);
or U3475 (N_3475,N_2560,N_2973);
or U3476 (N_3476,N_2685,N_2860);
nand U3477 (N_3477,N_2526,N_2868);
and U3478 (N_3478,N_2828,N_2697);
nand U3479 (N_3479,N_2574,N_2971);
nand U3480 (N_3480,N_2867,N_2615);
nor U3481 (N_3481,N_2830,N_2936);
nor U3482 (N_3482,N_2521,N_2712);
nand U3483 (N_3483,N_2871,N_2551);
nand U3484 (N_3484,N_2686,N_2534);
or U3485 (N_3485,N_2526,N_2946);
or U3486 (N_3486,N_2589,N_2736);
or U3487 (N_3487,N_2573,N_2529);
nor U3488 (N_3488,N_2790,N_2985);
and U3489 (N_3489,N_2516,N_2988);
or U3490 (N_3490,N_2715,N_2825);
nor U3491 (N_3491,N_2553,N_2743);
nor U3492 (N_3492,N_2899,N_2805);
and U3493 (N_3493,N_2532,N_2536);
nand U3494 (N_3494,N_2667,N_2723);
nand U3495 (N_3495,N_2829,N_2714);
or U3496 (N_3496,N_2733,N_2803);
nor U3497 (N_3497,N_2645,N_2547);
nand U3498 (N_3498,N_2855,N_2797);
and U3499 (N_3499,N_2846,N_2673);
nor U3500 (N_3500,N_3223,N_3464);
nand U3501 (N_3501,N_3422,N_3045);
nor U3502 (N_3502,N_3100,N_3062);
nand U3503 (N_3503,N_3297,N_3111);
nand U3504 (N_3504,N_3063,N_3316);
nand U3505 (N_3505,N_3109,N_3147);
nor U3506 (N_3506,N_3435,N_3009);
nand U3507 (N_3507,N_3451,N_3126);
or U3508 (N_3508,N_3014,N_3463);
or U3509 (N_3509,N_3124,N_3005);
nor U3510 (N_3510,N_3467,N_3097);
xor U3511 (N_3511,N_3168,N_3036);
and U3512 (N_3512,N_3074,N_3145);
nor U3513 (N_3513,N_3098,N_3397);
and U3514 (N_3514,N_3362,N_3341);
and U3515 (N_3515,N_3001,N_3418);
nor U3516 (N_3516,N_3123,N_3255);
nand U3517 (N_3517,N_3188,N_3204);
nand U3518 (N_3518,N_3459,N_3018);
or U3519 (N_3519,N_3020,N_3049);
nor U3520 (N_3520,N_3402,N_3056);
or U3521 (N_3521,N_3305,N_3284);
nand U3522 (N_3522,N_3162,N_3154);
nand U3523 (N_3523,N_3432,N_3006);
or U3524 (N_3524,N_3291,N_3114);
nand U3525 (N_3525,N_3071,N_3338);
and U3526 (N_3526,N_3233,N_3192);
nor U3527 (N_3527,N_3383,N_3398);
nand U3528 (N_3528,N_3299,N_3053);
or U3529 (N_3529,N_3148,N_3248);
nor U3530 (N_3530,N_3271,N_3019);
and U3531 (N_3531,N_3160,N_3215);
nor U3532 (N_3532,N_3129,N_3121);
or U3533 (N_3533,N_3391,N_3473);
or U3534 (N_3534,N_3158,N_3348);
nor U3535 (N_3535,N_3242,N_3417);
nand U3536 (N_3536,N_3280,N_3149);
or U3537 (N_3537,N_3293,N_3039);
and U3538 (N_3538,N_3198,N_3441);
or U3539 (N_3539,N_3450,N_3170);
nor U3540 (N_3540,N_3414,N_3484);
or U3541 (N_3541,N_3183,N_3349);
nand U3542 (N_3542,N_3191,N_3252);
nor U3543 (N_3543,N_3285,N_3048);
or U3544 (N_3544,N_3073,N_3259);
or U3545 (N_3545,N_3120,N_3491);
xor U3546 (N_3546,N_3337,N_3013);
nand U3547 (N_3547,N_3246,N_3393);
nand U3548 (N_3548,N_3262,N_3258);
or U3549 (N_3549,N_3064,N_3031);
nand U3550 (N_3550,N_3260,N_3446);
or U3551 (N_3551,N_3241,N_3361);
nand U3552 (N_3552,N_3288,N_3156);
and U3553 (N_3553,N_3218,N_3408);
nand U3554 (N_3554,N_3167,N_3263);
nor U3555 (N_3555,N_3323,N_3221);
and U3556 (N_3556,N_3294,N_3070);
nor U3557 (N_3557,N_3139,N_3388);
or U3558 (N_3558,N_3261,N_3104);
nand U3559 (N_3559,N_3022,N_3000);
or U3560 (N_3560,N_3365,N_3180);
nor U3561 (N_3561,N_3310,N_3272);
and U3562 (N_3562,N_3201,N_3407);
or U3563 (N_3563,N_3225,N_3436);
and U3564 (N_3564,N_3151,N_3222);
and U3565 (N_3565,N_3496,N_3395);
or U3566 (N_3566,N_3283,N_3102);
or U3567 (N_3567,N_3229,N_3003);
or U3568 (N_3568,N_3159,N_3041);
nor U3569 (N_3569,N_3057,N_3356);
nand U3570 (N_3570,N_3421,N_3430);
nor U3571 (N_3571,N_3286,N_3081);
and U3572 (N_3572,N_3174,N_3083);
and U3573 (N_3573,N_3250,N_3352);
or U3574 (N_3574,N_3406,N_3029);
or U3575 (N_3575,N_3219,N_3091);
and U3576 (N_3576,N_3217,N_3420);
nand U3577 (N_3577,N_3405,N_3131);
or U3578 (N_3578,N_3208,N_3290);
nand U3579 (N_3579,N_3309,N_3419);
and U3580 (N_3580,N_3375,N_3134);
nor U3581 (N_3581,N_3460,N_3412);
and U3582 (N_3582,N_3313,N_3302);
nor U3583 (N_3583,N_3269,N_3021);
nand U3584 (N_3584,N_3240,N_3401);
nand U3585 (N_3585,N_3171,N_3426);
nor U3586 (N_3586,N_3343,N_3153);
nand U3587 (N_3587,N_3178,N_3227);
or U3588 (N_3588,N_3187,N_3437);
nor U3589 (N_3589,N_3157,N_3060);
nand U3590 (N_3590,N_3366,N_3199);
nor U3591 (N_3591,N_3237,N_3433);
nor U3592 (N_3592,N_3332,N_3253);
or U3593 (N_3593,N_3330,N_3085);
xor U3594 (N_3594,N_3303,N_3068);
nand U3595 (N_3595,N_3108,N_3236);
or U3596 (N_3596,N_3069,N_3054);
or U3597 (N_3597,N_3354,N_3127);
nor U3598 (N_3598,N_3251,N_3386);
and U3599 (N_3599,N_3358,N_3184);
nand U3600 (N_3600,N_3080,N_3175);
nand U3601 (N_3601,N_3257,N_3472);
and U3602 (N_3602,N_3470,N_3359);
nand U3603 (N_3603,N_3346,N_3497);
nand U3604 (N_3604,N_3044,N_3442);
nand U3605 (N_3605,N_3007,N_3445);
or U3606 (N_3606,N_3276,N_3385);
and U3607 (N_3607,N_3231,N_3119);
and U3608 (N_3608,N_3243,N_3090);
and U3609 (N_3609,N_3480,N_3440);
or U3610 (N_3610,N_3249,N_3471);
nor U3611 (N_3611,N_3220,N_3452);
xnor U3612 (N_3612,N_3469,N_3169);
nor U3613 (N_3613,N_3125,N_3392);
nor U3614 (N_3614,N_3270,N_3319);
and U3615 (N_3615,N_3334,N_3403);
and U3616 (N_3616,N_3015,N_3328);
xnor U3617 (N_3617,N_3034,N_3457);
and U3618 (N_3618,N_3027,N_3304);
nand U3619 (N_3619,N_3117,N_3380);
or U3620 (N_3620,N_3038,N_3382);
and U3621 (N_3621,N_3494,N_3481);
and U3622 (N_3622,N_3458,N_3110);
xor U3623 (N_3623,N_3128,N_3295);
or U3624 (N_3624,N_3166,N_3389);
nand U3625 (N_3625,N_3072,N_3493);
nand U3626 (N_3626,N_3321,N_3378);
and U3627 (N_3627,N_3092,N_3028);
nand U3628 (N_3628,N_3101,N_3492);
nand U3629 (N_3629,N_3112,N_3331);
nor U3630 (N_3630,N_3194,N_3279);
nor U3631 (N_3631,N_3143,N_3483);
nand U3632 (N_3632,N_3344,N_3468);
nor U3633 (N_3633,N_3339,N_3146);
nor U3634 (N_3634,N_3353,N_3179);
xnor U3635 (N_3635,N_3043,N_3274);
nand U3636 (N_3636,N_3399,N_3444);
nor U3637 (N_3637,N_3089,N_3379);
nand U3638 (N_3638,N_3144,N_3454);
nand U3639 (N_3639,N_3202,N_3059);
and U3640 (N_3640,N_3413,N_3161);
nand U3641 (N_3641,N_3372,N_3448);
nor U3642 (N_3642,N_3315,N_3118);
nor U3643 (N_3643,N_3106,N_3396);
and U3644 (N_3644,N_3335,N_3008);
and U3645 (N_3645,N_3498,N_3115);
and U3646 (N_3646,N_3163,N_3487);
and U3647 (N_3647,N_3244,N_3010);
nand U3648 (N_3648,N_3189,N_3004);
nor U3649 (N_3649,N_3046,N_3278);
and U3650 (N_3650,N_3411,N_3226);
nand U3651 (N_3651,N_3181,N_3096);
nand U3652 (N_3652,N_3076,N_3176);
or U3653 (N_3653,N_3475,N_3256);
nor U3654 (N_3654,N_3340,N_3336);
and U3655 (N_3655,N_3416,N_3326);
nor U3656 (N_3656,N_3314,N_3488);
nor U3657 (N_3657,N_3002,N_3431);
nor U3658 (N_3658,N_3023,N_3351);
nand U3659 (N_3659,N_3363,N_3322);
nor U3660 (N_3660,N_3479,N_3387);
nand U3661 (N_3661,N_3087,N_3084);
or U3662 (N_3662,N_3301,N_3245);
and U3663 (N_3663,N_3312,N_3094);
nand U3664 (N_3664,N_3055,N_3474);
nor U3665 (N_3665,N_3093,N_3429);
nor U3666 (N_3666,N_3200,N_3230);
or U3667 (N_3667,N_3224,N_3462);
or U3668 (N_3668,N_3499,N_3186);
nand U3669 (N_3669,N_3424,N_3207);
and U3670 (N_3670,N_3369,N_3275);
or U3671 (N_3671,N_3376,N_3026);
and U3672 (N_3672,N_3485,N_3364);
or U3673 (N_3673,N_3374,N_3177);
nand U3674 (N_3674,N_3132,N_3265);
nand U3675 (N_3675,N_3113,N_3235);
nand U3676 (N_3676,N_3105,N_3409);
nor U3677 (N_3677,N_3486,N_3152);
nor U3678 (N_3678,N_3035,N_3453);
nand U3679 (N_3679,N_3052,N_3185);
xor U3680 (N_3680,N_3012,N_3423);
and U3681 (N_3681,N_3317,N_3078);
or U3682 (N_3682,N_3357,N_3032);
nor U3683 (N_3683,N_3306,N_3228);
nand U3684 (N_3684,N_3033,N_3211);
or U3685 (N_3685,N_3050,N_3307);
nand U3686 (N_3686,N_3190,N_3209);
and U3687 (N_3687,N_3086,N_3368);
or U3688 (N_3688,N_3427,N_3047);
and U3689 (N_3689,N_3287,N_3327);
nor U3690 (N_3690,N_3193,N_3282);
and U3691 (N_3691,N_3206,N_3267);
or U3692 (N_3692,N_3449,N_3333);
and U3693 (N_3693,N_3040,N_3042);
nor U3694 (N_3694,N_3088,N_3140);
nand U3695 (N_3695,N_3425,N_3077);
nand U3696 (N_3696,N_3212,N_3030);
and U3697 (N_3697,N_3173,N_3277);
nand U3698 (N_3698,N_3067,N_3325);
and U3699 (N_3699,N_3273,N_3011);
nand U3700 (N_3700,N_3490,N_3311);
nor U3701 (N_3701,N_3238,N_3371);
and U3702 (N_3702,N_3350,N_3400);
nor U3703 (N_3703,N_3136,N_3107);
nand U3704 (N_3704,N_3196,N_3443);
nand U3705 (N_3705,N_3320,N_3075);
or U3706 (N_3706,N_3234,N_3016);
nor U3707 (N_3707,N_3347,N_3342);
or U3708 (N_3708,N_3197,N_3203);
xor U3709 (N_3709,N_3345,N_3438);
nand U3710 (N_3710,N_3439,N_3103);
nand U3711 (N_3711,N_3355,N_3037);
nand U3712 (N_3712,N_3182,N_3130);
nor U3713 (N_3713,N_3298,N_3165);
nor U3714 (N_3714,N_3377,N_3456);
nor U3715 (N_3715,N_3482,N_3466);
nand U3716 (N_3716,N_3410,N_3150);
and U3717 (N_3717,N_3254,N_3434);
nor U3718 (N_3718,N_3142,N_3061);
nor U3719 (N_3719,N_3082,N_3195);
and U3720 (N_3720,N_3058,N_3205);
and U3721 (N_3721,N_3210,N_3318);
nand U3722 (N_3722,N_3264,N_3268);
and U3723 (N_3723,N_3477,N_3370);
xnor U3724 (N_3724,N_3360,N_3164);
or U3725 (N_3725,N_3384,N_3465);
nand U3726 (N_3726,N_3135,N_3478);
or U3727 (N_3727,N_3172,N_3247);
nor U3728 (N_3728,N_3415,N_3116);
or U3729 (N_3729,N_3495,N_3079);
and U3730 (N_3730,N_3099,N_3373);
and U3731 (N_3731,N_3394,N_3367);
or U3732 (N_3732,N_3025,N_3017);
or U3733 (N_3733,N_3447,N_3051);
nor U3734 (N_3734,N_3213,N_3289);
or U3735 (N_3735,N_3232,N_3381);
and U3736 (N_3736,N_3095,N_3214);
nand U3737 (N_3737,N_3404,N_3300);
or U3738 (N_3738,N_3296,N_3266);
or U3739 (N_3739,N_3141,N_3137);
and U3740 (N_3740,N_3138,N_3329);
nand U3741 (N_3741,N_3390,N_3239);
and U3742 (N_3742,N_3324,N_3281);
and U3743 (N_3743,N_3216,N_3489);
or U3744 (N_3744,N_3461,N_3066);
and U3745 (N_3745,N_3065,N_3476);
and U3746 (N_3746,N_3133,N_3122);
nor U3747 (N_3747,N_3292,N_3428);
and U3748 (N_3748,N_3024,N_3455);
or U3749 (N_3749,N_3155,N_3308);
and U3750 (N_3750,N_3104,N_3041);
or U3751 (N_3751,N_3088,N_3029);
nor U3752 (N_3752,N_3264,N_3223);
and U3753 (N_3753,N_3374,N_3419);
and U3754 (N_3754,N_3089,N_3032);
nand U3755 (N_3755,N_3165,N_3439);
nor U3756 (N_3756,N_3229,N_3343);
and U3757 (N_3757,N_3101,N_3244);
or U3758 (N_3758,N_3385,N_3236);
and U3759 (N_3759,N_3478,N_3091);
or U3760 (N_3760,N_3468,N_3021);
or U3761 (N_3761,N_3410,N_3022);
nand U3762 (N_3762,N_3000,N_3266);
or U3763 (N_3763,N_3058,N_3005);
nor U3764 (N_3764,N_3148,N_3044);
and U3765 (N_3765,N_3225,N_3459);
or U3766 (N_3766,N_3184,N_3108);
and U3767 (N_3767,N_3333,N_3061);
and U3768 (N_3768,N_3330,N_3087);
or U3769 (N_3769,N_3323,N_3244);
or U3770 (N_3770,N_3462,N_3104);
nor U3771 (N_3771,N_3421,N_3291);
or U3772 (N_3772,N_3457,N_3071);
nor U3773 (N_3773,N_3381,N_3143);
or U3774 (N_3774,N_3483,N_3048);
nand U3775 (N_3775,N_3183,N_3180);
nand U3776 (N_3776,N_3288,N_3153);
or U3777 (N_3777,N_3476,N_3034);
or U3778 (N_3778,N_3476,N_3164);
or U3779 (N_3779,N_3298,N_3199);
nor U3780 (N_3780,N_3144,N_3222);
nand U3781 (N_3781,N_3129,N_3109);
or U3782 (N_3782,N_3445,N_3364);
nand U3783 (N_3783,N_3365,N_3461);
nand U3784 (N_3784,N_3490,N_3072);
or U3785 (N_3785,N_3404,N_3442);
nor U3786 (N_3786,N_3246,N_3437);
or U3787 (N_3787,N_3445,N_3170);
and U3788 (N_3788,N_3159,N_3277);
nand U3789 (N_3789,N_3044,N_3134);
nor U3790 (N_3790,N_3135,N_3231);
and U3791 (N_3791,N_3048,N_3320);
and U3792 (N_3792,N_3161,N_3336);
or U3793 (N_3793,N_3012,N_3326);
nor U3794 (N_3794,N_3332,N_3105);
nor U3795 (N_3795,N_3376,N_3319);
nor U3796 (N_3796,N_3450,N_3421);
and U3797 (N_3797,N_3145,N_3107);
nand U3798 (N_3798,N_3034,N_3018);
and U3799 (N_3799,N_3142,N_3372);
nor U3800 (N_3800,N_3091,N_3377);
nand U3801 (N_3801,N_3250,N_3022);
and U3802 (N_3802,N_3423,N_3300);
nand U3803 (N_3803,N_3126,N_3406);
nor U3804 (N_3804,N_3088,N_3136);
nor U3805 (N_3805,N_3032,N_3028);
and U3806 (N_3806,N_3428,N_3205);
or U3807 (N_3807,N_3263,N_3050);
nor U3808 (N_3808,N_3366,N_3309);
or U3809 (N_3809,N_3429,N_3137);
nor U3810 (N_3810,N_3295,N_3031);
nand U3811 (N_3811,N_3295,N_3451);
and U3812 (N_3812,N_3194,N_3269);
or U3813 (N_3813,N_3347,N_3300);
or U3814 (N_3814,N_3390,N_3167);
or U3815 (N_3815,N_3478,N_3000);
nand U3816 (N_3816,N_3369,N_3160);
or U3817 (N_3817,N_3111,N_3315);
nand U3818 (N_3818,N_3338,N_3239);
or U3819 (N_3819,N_3438,N_3350);
nor U3820 (N_3820,N_3395,N_3347);
nor U3821 (N_3821,N_3211,N_3021);
xor U3822 (N_3822,N_3287,N_3315);
or U3823 (N_3823,N_3004,N_3249);
nand U3824 (N_3824,N_3278,N_3024);
nor U3825 (N_3825,N_3104,N_3406);
nor U3826 (N_3826,N_3088,N_3284);
nor U3827 (N_3827,N_3275,N_3399);
and U3828 (N_3828,N_3027,N_3026);
or U3829 (N_3829,N_3027,N_3386);
nand U3830 (N_3830,N_3241,N_3036);
nand U3831 (N_3831,N_3108,N_3175);
nor U3832 (N_3832,N_3228,N_3142);
nor U3833 (N_3833,N_3128,N_3131);
or U3834 (N_3834,N_3161,N_3120);
nand U3835 (N_3835,N_3094,N_3332);
and U3836 (N_3836,N_3191,N_3140);
and U3837 (N_3837,N_3156,N_3420);
nand U3838 (N_3838,N_3186,N_3394);
or U3839 (N_3839,N_3259,N_3093);
and U3840 (N_3840,N_3489,N_3466);
and U3841 (N_3841,N_3404,N_3343);
and U3842 (N_3842,N_3225,N_3019);
and U3843 (N_3843,N_3261,N_3102);
and U3844 (N_3844,N_3295,N_3472);
nor U3845 (N_3845,N_3052,N_3200);
nor U3846 (N_3846,N_3428,N_3235);
and U3847 (N_3847,N_3203,N_3082);
and U3848 (N_3848,N_3389,N_3059);
xor U3849 (N_3849,N_3369,N_3276);
nand U3850 (N_3850,N_3168,N_3084);
nor U3851 (N_3851,N_3188,N_3489);
nor U3852 (N_3852,N_3367,N_3028);
nor U3853 (N_3853,N_3042,N_3405);
or U3854 (N_3854,N_3392,N_3478);
nand U3855 (N_3855,N_3437,N_3165);
nor U3856 (N_3856,N_3433,N_3221);
and U3857 (N_3857,N_3307,N_3433);
and U3858 (N_3858,N_3372,N_3453);
and U3859 (N_3859,N_3139,N_3157);
and U3860 (N_3860,N_3380,N_3319);
nand U3861 (N_3861,N_3278,N_3362);
nand U3862 (N_3862,N_3265,N_3220);
and U3863 (N_3863,N_3275,N_3414);
nor U3864 (N_3864,N_3038,N_3081);
nor U3865 (N_3865,N_3381,N_3061);
nor U3866 (N_3866,N_3351,N_3172);
xnor U3867 (N_3867,N_3112,N_3442);
nor U3868 (N_3868,N_3162,N_3398);
and U3869 (N_3869,N_3188,N_3423);
or U3870 (N_3870,N_3101,N_3145);
nor U3871 (N_3871,N_3379,N_3219);
nor U3872 (N_3872,N_3108,N_3411);
and U3873 (N_3873,N_3128,N_3321);
and U3874 (N_3874,N_3410,N_3067);
or U3875 (N_3875,N_3104,N_3216);
nor U3876 (N_3876,N_3451,N_3382);
nor U3877 (N_3877,N_3074,N_3352);
and U3878 (N_3878,N_3030,N_3386);
and U3879 (N_3879,N_3002,N_3106);
and U3880 (N_3880,N_3170,N_3473);
nand U3881 (N_3881,N_3357,N_3053);
and U3882 (N_3882,N_3295,N_3453);
nor U3883 (N_3883,N_3338,N_3352);
or U3884 (N_3884,N_3387,N_3020);
nand U3885 (N_3885,N_3186,N_3079);
and U3886 (N_3886,N_3425,N_3278);
nand U3887 (N_3887,N_3106,N_3205);
and U3888 (N_3888,N_3428,N_3490);
and U3889 (N_3889,N_3368,N_3472);
and U3890 (N_3890,N_3169,N_3196);
nand U3891 (N_3891,N_3394,N_3441);
nor U3892 (N_3892,N_3032,N_3429);
and U3893 (N_3893,N_3262,N_3158);
nor U3894 (N_3894,N_3315,N_3430);
or U3895 (N_3895,N_3430,N_3132);
or U3896 (N_3896,N_3348,N_3498);
nor U3897 (N_3897,N_3484,N_3451);
nor U3898 (N_3898,N_3337,N_3155);
and U3899 (N_3899,N_3029,N_3004);
nand U3900 (N_3900,N_3303,N_3074);
nand U3901 (N_3901,N_3256,N_3170);
and U3902 (N_3902,N_3203,N_3317);
or U3903 (N_3903,N_3181,N_3447);
nor U3904 (N_3904,N_3269,N_3100);
xor U3905 (N_3905,N_3193,N_3023);
nor U3906 (N_3906,N_3217,N_3442);
and U3907 (N_3907,N_3047,N_3025);
and U3908 (N_3908,N_3239,N_3172);
and U3909 (N_3909,N_3294,N_3174);
and U3910 (N_3910,N_3158,N_3320);
or U3911 (N_3911,N_3393,N_3103);
or U3912 (N_3912,N_3483,N_3387);
xor U3913 (N_3913,N_3284,N_3082);
nor U3914 (N_3914,N_3127,N_3005);
xnor U3915 (N_3915,N_3429,N_3158);
nor U3916 (N_3916,N_3488,N_3254);
nand U3917 (N_3917,N_3180,N_3499);
and U3918 (N_3918,N_3133,N_3498);
and U3919 (N_3919,N_3484,N_3327);
or U3920 (N_3920,N_3361,N_3427);
nor U3921 (N_3921,N_3436,N_3339);
nand U3922 (N_3922,N_3348,N_3491);
nor U3923 (N_3923,N_3155,N_3362);
or U3924 (N_3924,N_3284,N_3017);
nor U3925 (N_3925,N_3400,N_3478);
and U3926 (N_3926,N_3347,N_3492);
or U3927 (N_3927,N_3446,N_3144);
nor U3928 (N_3928,N_3087,N_3299);
and U3929 (N_3929,N_3409,N_3270);
or U3930 (N_3930,N_3210,N_3392);
and U3931 (N_3931,N_3399,N_3159);
nor U3932 (N_3932,N_3410,N_3018);
nand U3933 (N_3933,N_3390,N_3488);
nor U3934 (N_3934,N_3089,N_3497);
nand U3935 (N_3935,N_3167,N_3395);
nand U3936 (N_3936,N_3336,N_3164);
nor U3937 (N_3937,N_3076,N_3287);
nand U3938 (N_3938,N_3192,N_3377);
nand U3939 (N_3939,N_3167,N_3360);
xor U3940 (N_3940,N_3483,N_3372);
or U3941 (N_3941,N_3117,N_3047);
nor U3942 (N_3942,N_3022,N_3498);
nand U3943 (N_3943,N_3022,N_3261);
nor U3944 (N_3944,N_3017,N_3107);
and U3945 (N_3945,N_3212,N_3173);
nand U3946 (N_3946,N_3227,N_3406);
nand U3947 (N_3947,N_3394,N_3134);
or U3948 (N_3948,N_3178,N_3335);
nor U3949 (N_3949,N_3040,N_3313);
and U3950 (N_3950,N_3164,N_3017);
or U3951 (N_3951,N_3436,N_3437);
and U3952 (N_3952,N_3014,N_3371);
or U3953 (N_3953,N_3427,N_3059);
nor U3954 (N_3954,N_3163,N_3084);
nor U3955 (N_3955,N_3372,N_3460);
and U3956 (N_3956,N_3490,N_3226);
nand U3957 (N_3957,N_3022,N_3017);
or U3958 (N_3958,N_3473,N_3359);
xnor U3959 (N_3959,N_3392,N_3183);
or U3960 (N_3960,N_3245,N_3193);
and U3961 (N_3961,N_3074,N_3080);
and U3962 (N_3962,N_3217,N_3318);
xor U3963 (N_3963,N_3394,N_3387);
or U3964 (N_3964,N_3005,N_3192);
xor U3965 (N_3965,N_3111,N_3337);
nor U3966 (N_3966,N_3262,N_3093);
or U3967 (N_3967,N_3166,N_3377);
and U3968 (N_3968,N_3313,N_3358);
and U3969 (N_3969,N_3282,N_3293);
or U3970 (N_3970,N_3391,N_3076);
nand U3971 (N_3971,N_3004,N_3401);
or U3972 (N_3972,N_3316,N_3183);
nand U3973 (N_3973,N_3454,N_3237);
and U3974 (N_3974,N_3472,N_3088);
nor U3975 (N_3975,N_3131,N_3145);
or U3976 (N_3976,N_3004,N_3130);
nand U3977 (N_3977,N_3150,N_3202);
nor U3978 (N_3978,N_3244,N_3357);
nand U3979 (N_3979,N_3489,N_3112);
nor U3980 (N_3980,N_3378,N_3115);
and U3981 (N_3981,N_3186,N_3002);
or U3982 (N_3982,N_3148,N_3147);
or U3983 (N_3983,N_3135,N_3243);
xor U3984 (N_3984,N_3483,N_3095);
and U3985 (N_3985,N_3118,N_3037);
and U3986 (N_3986,N_3426,N_3090);
or U3987 (N_3987,N_3412,N_3226);
or U3988 (N_3988,N_3006,N_3105);
nand U3989 (N_3989,N_3072,N_3316);
or U3990 (N_3990,N_3073,N_3277);
nor U3991 (N_3991,N_3055,N_3477);
and U3992 (N_3992,N_3121,N_3003);
nor U3993 (N_3993,N_3480,N_3335);
nor U3994 (N_3994,N_3166,N_3231);
nor U3995 (N_3995,N_3452,N_3338);
xor U3996 (N_3996,N_3463,N_3446);
or U3997 (N_3997,N_3448,N_3115);
and U3998 (N_3998,N_3299,N_3409);
nand U3999 (N_3999,N_3226,N_3125);
and U4000 (N_4000,N_3635,N_3629);
and U4001 (N_4001,N_3519,N_3749);
or U4002 (N_4002,N_3618,N_3526);
and U4003 (N_4003,N_3632,N_3910);
or U4004 (N_4004,N_3995,N_3872);
and U4005 (N_4005,N_3556,N_3883);
and U4006 (N_4006,N_3863,N_3642);
and U4007 (N_4007,N_3805,N_3668);
and U4008 (N_4008,N_3921,N_3891);
or U4009 (N_4009,N_3583,N_3820);
and U4010 (N_4010,N_3747,N_3829);
or U4011 (N_4011,N_3649,N_3616);
and U4012 (N_4012,N_3544,N_3599);
nor U4013 (N_4013,N_3865,N_3907);
or U4014 (N_4014,N_3550,N_3906);
or U4015 (N_4015,N_3680,N_3740);
and U4016 (N_4016,N_3662,N_3617);
xnor U4017 (N_4017,N_3693,N_3752);
nand U4018 (N_4018,N_3535,N_3842);
and U4019 (N_4019,N_3890,N_3646);
and U4020 (N_4020,N_3847,N_3584);
or U4021 (N_4021,N_3553,N_3620);
nand U4022 (N_4022,N_3887,N_3835);
or U4023 (N_4023,N_3857,N_3575);
nor U4024 (N_4024,N_3688,N_3705);
nor U4025 (N_4025,N_3561,N_3798);
and U4026 (N_4026,N_3716,N_3679);
nor U4027 (N_4027,N_3904,N_3937);
xnor U4028 (N_4028,N_3993,N_3969);
nand U4029 (N_4029,N_3508,N_3780);
or U4030 (N_4030,N_3729,N_3502);
nand U4031 (N_4031,N_3673,N_3771);
and U4032 (N_4032,N_3999,N_3717);
nor U4033 (N_4033,N_3855,N_3725);
or U4034 (N_4034,N_3784,N_3726);
nor U4035 (N_4035,N_3742,N_3597);
or U4036 (N_4036,N_3785,N_3852);
or U4037 (N_4037,N_3922,N_3657);
nand U4038 (N_4038,N_3702,N_3875);
nor U4039 (N_4039,N_3861,N_3941);
or U4040 (N_4040,N_3723,N_3984);
nor U4041 (N_4041,N_3958,N_3968);
or U4042 (N_4042,N_3713,N_3607);
nor U4043 (N_4043,N_3671,N_3568);
nand U4044 (N_4044,N_3640,N_3631);
nand U4045 (N_4045,N_3858,N_3976);
nand U4046 (N_4046,N_3707,N_3722);
or U4047 (N_4047,N_3848,N_3677);
nor U4048 (N_4048,N_3555,N_3945);
and U4049 (N_4049,N_3776,N_3572);
nor U4050 (N_4050,N_3912,N_3648);
or U4051 (N_4051,N_3990,N_3503);
nor U4052 (N_4052,N_3903,N_3719);
and U4053 (N_4053,N_3956,N_3889);
nand U4054 (N_4054,N_3734,N_3926);
nor U4055 (N_4055,N_3661,N_3695);
or U4056 (N_4056,N_3739,N_3938);
nand U4057 (N_4057,N_3586,N_3853);
or U4058 (N_4058,N_3982,N_3510);
and U4059 (N_4059,N_3626,N_3806);
or U4060 (N_4060,N_3892,N_3779);
and U4061 (N_4061,N_3778,N_3754);
nand U4062 (N_4062,N_3675,N_3953);
nor U4063 (N_4063,N_3957,N_3621);
and U4064 (N_4064,N_3975,N_3745);
nand U4065 (N_4065,N_3582,N_3951);
and U4066 (N_4066,N_3913,N_3727);
nor U4067 (N_4067,N_3610,N_3560);
nor U4068 (N_4068,N_3652,N_3691);
and U4069 (N_4069,N_3793,N_3974);
nand U4070 (N_4070,N_3682,N_3638);
or U4071 (N_4071,N_3894,N_3714);
nand U4072 (N_4072,N_3542,N_3522);
nor U4073 (N_4073,N_3833,N_3843);
and U4074 (N_4074,N_3708,N_3971);
or U4075 (N_4075,N_3602,N_3543);
nand U4076 (N_4076,N_3942,N_3998);
nor U4077 (N_4077,N_3670,N_3573);
or U4078 (N_4078,N_3834,N_3751);
xnor U4079 (N_4079,N_3647,N_3686);
nor U4080 (N_4080,N_3789,N_3905);
nand U4081 (N_4081,N_3733,N_3523);
nor U4082 (N_4082,N_3548,N_3792);
xor U4083 (N_4083,N_3783,N_3914);
xor U4084 (N_4084,N_3917,N_3770);
nand U4085 (N_4085,N_3655,N_3940);
or U4086 (N_4086,N_3732,N_3637);
and U4087 (N_4087,N_3870,N_3797);
or U4088 (N_4088,N_3966,N_3815);
nand U4089 (N_4089,N_3939,N_3593);
nand U4090 (N_4090,N_3932,N_3881);
nand U4091 (N_4091,N_3669,N_3823);
xnor U4092 (N_4092,N_3816,N_3501);
or U4093 (N_4093,N_3918,N_3933);
and U4094 (N_4094,N_3860,N_3769);
nor U4095 (N_4095,N_3827,N_3554);
or U4096 (N_4096,N_3868,N_3692);
nor U4097 (N_4097,N_3962,N_3694);
nand U4098 (N_4098,N_3529,N_3651);
and U4099 (N_4099,N_3928,N_3831);
or U4100 (N_4100,N_3633,N_3521);
and U4101 (N_4101,N_3867,N_3660);
nand U4102 (N_4102,N_3977,N_3799);
or U4103 (N_4103,N_3600,N_3753);
or U4104 (N_4104,N_3514,N_3934);
nand U4105 (N_4105,N_3886,N_3871);
xnor U4106 (N_4106,N_3624,N_3796);
nor U4107 (N_4107,N_3809,N_3609);
or U4108 (N_4108,N_3737,N_3768);
and U4109 (N_4109,N_3813,N_3577);
and U4110 (N_4110,N_3674,N_3988);
and U4111 (N_4111,N_3516,N_3760);
nor U4112 (N_4112,N_3690,N_3930);
or U4113 (N_4113,N_3985,N_3558);
and U4114 (N_4114,N_3672,N_3505);
nand U4115 (N_4115,N_3534,N_3955);
or U4116 (N_4116,N_3807,N_3791);
and U4117 (N_4117,N_3808,N_3866);
and U4118 (N_4118,N_3664,N_3736);
nor U4119 (N_4119,N_3997,N_3927);
nor U4120 (N_4120,N_3830,N_3764);
nand U4121 (N_4121,N_3720,N_3828);
nand U4122 (N_4122,N_3517,N_3588);
nand U4123 (N_4123,N_3884,N_3836);
or U4124 (N_4124,N_3810,N_3619);
nor U4125 (N_4125,N_3876,N_3520);
nand U4126 (N_4126,N_3538,N_3518);
nor U4127 (N_4127,N_3731,N_3859);
nor U4128 (N_4128,N_3525,N_3874);
and U4129 (N_4129,N_3724,N_3949);
and U4130 (N_4130,N_3856,N_3512);
nor U4131 (N_4131,N_3781,N_3775);
and U4132 (N_4132,N_3978,N_3511);
nand U4133 (N_4133,N_3580,N_3551);
or U4134 (N_4134,N_3946,N_3825);
nor U4135 (N_4135,N_3678,N_3862);
nor U4136 (N_4136,N_3822,N_3546);
nand U4137 (N_4137,N_3909,N_3804);
nor U4138 (N_4138,N_3954,N_3541);
or U4139 (N_4139,N_3948,N_3832);
xor U4140 (N_4140,N_3959,N_3826);
and U4141 (N_4141,N_3574,N_3645);
or U4142 (N_4142,N_3824,N_3794);
nor U4143 (N_4143,N_3559,N_3986);
or U4144 (N_4144,N_3960,N_3801);
or U4145 (N_4145,N_3812,N_3636);
nor U4146 (N_4146,N_3601,N_3895);
xnor U4147 (N_4147,N_3701,N_3681);
and U4148 (N_4148,N_3613,N_3911);
nor U4149 (N_4149,N_3898,N_3961);
xnor U4150 (N_4150,N_3689,N_3899);
nor U4151 (N_4151,N_3598,N_3735);
and U4152 (N_4152,N_3973,N_3612);
and U4153 (N_4153,N_3579,N_3924);
nand U4154 (N_4154,N_3515,N_3786);
xnor U4155 (N_4155,N_3614,N_3592);
nand U4156 (N_4156,N_3897,N_3545);
nand U4157 (N_4157,N_3700,N_3650);
nand U4158 (N_4158,N_3623,N_3654);
nand U4159 (N_4159,N_3659,N_3566);
and U4160 (N_4160,N_3838,N_3991);
or U4161 (N_4161,N_3811,N_3715);
or U4162 (N_4162,N_3880,N_3916);
or U4163 (N_4163,N_3711,N_3685);
and U4164 (N_4164,N_3531,N_3981);
nand U4165 (N_4165,N_3504,N_3676);
nand U4166 (N_4166,N_3996,N_3802);
and U4167 (N_4167,N_3712,N_3721);
nor U4168 (N_4168,N_3819,N_3761);
and U4169 (N_4169,N_3885,N_3596);
or U4170 (N_4170,N_3625,N_3639);
nand U4171 (N_4171,N_3604,N_3622);
and U4172 (N_4172,N_3697,N_3589);
nor U4173 (N_4173,N_3536,N_3901);
and U4174 (N_4174,N_3746,N_3594);
or U4175 (N_4175,N_3506,N_3571);
nand U4176 (N_4176,N_3743,N_3509);
or U4177 (N_4177,N_3931,N_3972);
xor U4178 (N_4178,N_3718,N_3943);
and U4179 (N_4179,N_3947,N_3790);
or U4180 (N_4180,N_3864,N_3795);
nand U4181 (N_4181,N_3565,N_3663);
nand U4182 (N_4182,N_3524,N_3845);
and U4183 (N_4183,N_3570,N_3630);
nor U4184 (N_4184,N_3709,N_3634);
nand U4185 (N_4185,N_3595,N_3666);
or U4186 (N_4186,N_3537,N_3562);
and U4187 (N_4187,N_3569,N_3952);
nor U4188 (N_4188,N_3567,N_3557);
or U4189 (N_4189,N_3530,N_3564);
nand U4190 (N_4190,N_3900,N_3627);
or U4191 (N_4191,N_3696,N_3765);
nor U4192 (N_4192,N_3849,N_3644);
nand U4193 (N_4193,N_3896,N_3590);
nand U4194 (N_4194,N_3994,N_3919);
nand U4195 (N_4195,N_3513,N_3665);
nand U4196 (N_4196,N_3656,N_3915);
and U4197 (N_4197,N_3605,N_3767);
and U4198 (N_4198,N_3839,N_3882);
and U4199 (N_4199,N_3762,N_3628);
nand U4200 (N_4200,N_3850,N_3980);
and U4201 (N_4201,N_3840,N_3888);
nand U4202 (N_4202,N_3773,N_3774);
nor U4203 (N_4203,N_3787,N_3758);
and U4204 (N_4204,N_3851,N_3532);
nor U4205 (N_4205,N_3533,N_3741);
and U4206 (N_4206,N_3684,N_3563);
and U4207 (N_4207,N_3967,N_3615);
and U4208 (N_4208,N_3788,N_3963);
or U4209 (N_4209,N_3983,N_3706);
and U4210 (N_4210,N_3821,N_3759);
nor U4211 (N_4211,N_3935,N_3877);
or U4212 (N_4212,N_3641,N_3687);
or U4213 (N_4213,N_3818,N_3920);
nand U4214 (N_4214,N_3539,N_3925);
or U4215 (N_4215,N_3527,N_3965);
nor U4216 (N_4216,N_3964,N_3869);
nand U4217 (N_4217,N_3606,N_3611);
nand U4218 (N_4218,N_3528,N_3970);
and U4219 (N_4219,N_3710,N_3944);
and U4220 (N_4220,N_3699,N_3581);
and U4221 (N_4221,N_3844,N_3540);
and U4222 (N_4222,N_3507,N_3750);
nand U4223 (N_4223,N_3578,N_3814);
or U4224 (N_4224,N_3591,N_3757);
nand U4225 (N_4225,N_3653,N_3667);
or U4226 (N_4226,N_3936,N_3817);
or U4227 (N_4227,N_3908,N_3552);
and U4228 (N_4228,N_3730,N_3603);
or U4229 (N_4229,N_3846,N_3587);
and U4230 (N_4230,N_3992,N_3800);
or U4231 (N_4231,N_3728,N_3837);
xnor U4232 (N_4232,N_3748,N_3879);
or U4233 (N_4233,N_3683,N_3500);
nand U4234 (N_4234,N_3763,N_3772);
nand U4235 (N_4235,N_3756,N_3744);
xnor U4236 (N_4236,N_3658,N_3854);
nand U4237 (N_4237,N_3777,N_3987);
nor U4238 (N_4238,N_3878,N_3893);
or U4239 (N_4239,N_3547,N_3549);
and U4240 (N_4240,N_3782,N_3738);
or U4241 (N_4241,N_3704,N_3698);
and U4242 (N_4242,N_3755,N_3585);
nand U4243 (N_4243,N_3576,N_3841);
or U4244 (N_4244,N_3608,N_3643);
xor U4245 (N_4245,N_3803,N_3979);
nor U4246 (N_4246,N_3989,N_3703);
xor U4247 (N_4247,N_3929,N_3766);
nor U4248 (N_4248,N_3873,N_3923);
and U4249 (N_4249,N_3950,N_3902);
and U4250 (N_4250,N_3726,N_3960);
nor U4251 (N_4251,N_3976,N_3950);
and U4252 (N_4252,N_3656,N_3512);
nand U4253 (N_4253,N_3846,N_3731);
and U4254 (N_4254,N_3885,N_3789);
nand U4255 (N_4255,N_3723,N_3671);
or U4256 (N_4256,N_3535,N_3999);
nor U4257 (N_4257,N_3692,N_3762);
or U4258 (N_4258,N_3992,N_3887);
or U4259 (N_4259,N_3957,N_3906);
or U4260 (N_4260,N_3629,N_3980);
and U4261 (N_4261,N_3918,N_3827);
nor U4262 (N_4262,N_3624,N_3587);
or U4263 (N_4263,N_3914,N_3689);
nand U4264 (N_4264,N_3552,N_3935);
nor U4265 (N_4265,N_3958,N_3636);
and U4266 (N_4266,N_3931,N_3616);
and U4267 (N_4267,N_3803,N_3624);
nor U4268 (N_4268,N_3986,N_3631);
or U4269 (N_4269,N_3576,N_3510);
and U4270 (N_4270,N_3881,N_3988);
nor U4271 (N_4271,N_3704,N_3910);
nor U4272 (N_4272,N_3929,N_3893);
nand U4273 (N_4273,N_3644,N_3901);
nor U4274 (N_4274,N_3884,N_3549);
nor U4275 (N_4275,N_3900,N_3841);
nand U4276 (N_4276,N_3985,N_3716);
xnor U4277 (N_4277,N_3582,N_3627);
nor U4278 (N_4278,N_3956,N_3557);
nor U4279 (N_4279,N_3794,N_3575);
nand U4280 (N_4280,N_3987,N_3533);
or U4281 (N_4281,N_3526,N_3993);
nand U4282 (N_4282,N_3653,N_3984);
nor U4283 (N_4283,N_3912,N_3903);
nand U4284 (N_4284,N_3668,N_3784);
nand U4285 (N_4285,N_3537,N_3775);
and U4286 (N_4286,N_3874,N_3721);
nand U4287 (N_4287,N_3615,N_3561);
xnor U4288 (N_4288,N_3660,N_3805);
and U4289 (N_4289,N_3553,N_3942);
nand U4290 (N_4290,N_3608,N_3854);
and U4291 (N_4291,N_3640,N_3981);
or U4292 (N_4292,N_3586,N_3836);
nand U4293 (N_4293,N_3653,N_3970);
nor U4294 (N_4294,N_3602,N_3978);
or U4295 (N_4295,N_3603,N_3946);
nand U4296 (N_4296,N_3664,N_3801);
and U4297 (N_4297,N_3893,N_3649);
nor U4298 (N_4298,N_3554,N_3671);
nand U4299 (N_4299,N_3674,N_3886);
or U4300 (N_4300,N_3516,N_3945);
and U4301 (N_4301,N_3679,N_3708);
or U4302 (N_4302,N_3842,N_3869);
nor U4303 (N_4303,N_3536,N_3719);
or U4304 (N_4304,N_3712,N_3951);
or U4305 (N_4305,N_3965,N_3973);
nand U4306 (N_4306,N_3669,N_3919);
and U4307 (N_4307,N_3577,N_3888);
nand U4308 (N_4308,N_3745,N_3768);
or U4309 (N_4309,N_3810,N_3512);
nand U4310 (N_4310,N_3709,N_3788);
and U4311 (N_4311,N_3820,N_3642);
nand U4312 (N_4312,N_3884,N_3671);
and U4313 (N_4313,N_3734,N_3814);
nand U4314 (N_4314,N_3699,N_3577);
nand U4315 (N_4315,N_3936,N_3860);
or U4316 (N_4316,N_3924,N_3887);
nand U4317 (N_4317,N_3678,N_3524);
or U4318 (N_4318,N_3747,N_3568);
and U4319 (N_4319,N_3767,N_3576);
and U4320 (N_4320,N_3722,N_3547);
and U4321 (N_4321,N_3512,N_3598);
nor U4322 (N_4322,N_3710,N_3595);
nand U4323 (N_4323,N_3962,N_3603);
nand U4324 (N_4324,N_3513,N_3621);
nand U4325 (N_4325,N_3951,N_3608);
or U4326 (N_4326,N_3646,N_3979);
nor U4327 (N_4327,N_3848,N_3563);
nor U4328 (N_4328,N_3686,N_3893);
nor U4329 (N_4329,N_3665,N_3515);
nor U4330 (N_4330,N_3953,N_3588);
or U4331 (N_4331,N_3681,N_3634);
or U4332 (N_4332,N_3809,N_3769);
nand U4333 (N_4333,N_3559,N_3519);
nor U4334 (N_4334,N_3956,N_3671);
nor U4335 (N_4335,N_3571,N_3863);
nand U4336 (N_4336,N_3949,N_3791);
and U4337 (N_4337,N_3603,N_3594);
or U4338 (N_4338,N_3652,N_3740);
or U4339 (N_4339,N_3789,N_3673);
and U4340 (N_4340,N_3701,N_3821);
or U4341 (N_4341,N_3829,N_3606);
or U4342 (N_4342,N_3954,N_3526);
or U4343 (N_4343,N_3685,N_3902);
or U4344 (N_4344,N_3676,N_3593);
xor U4345 (N_4345,N_3883,N_3990);
nand U4346 (N_4346,N_3874,N_3573);
or U4347 (N_4347,N_3899,N_3941);
or U4348 (N_4348,N_3929,N_3964);
and U4349 (N_4349,N_3935,N_3825);
and U4350 (N_4350,N_3878,N_3547);
or U4351 (N_4351,N_3748,N_3714);
or U4352 (N_4352,N_3817,N_3958);
nand U4353 (N_4353,N_3904,N_3528);
nor U4354 (N_4354,N_3690,N_3520);
nor U4355 (N_4355,N_3974,N_3845);
or U4356 (N_4356,N_3818,N_3636);
nand U4357 (N_4357,N_3667,N_3723);
nand U4358 (N_4358,N_3705,N_3528);
or U4359 (N_4359,N_3686,N_3835);
or U4360 (N_4360,N_3888,N_3596);
nand U4361 (N_4361,N_3668,N_3667);
or U4362 (N_4362,N_3694,N_3670);
and U4363 (N_4363,N_3665,N_3993);
and U4364 (N_4364,N_3521,N_3980);
nand U4365 (N_4365,N_3713,N_3724);
and U4366 (N_4366,N_3623,N_3747);
nor U4367 (N_4367,N_3996,N_3725);
nand U4368 (N_4368,N_3791,N_3814);
nand U4369 (N_4369,N_3634,N_3955);
and U4370 (N_4370,N_3503,N_3560);
or U4371 (N_4371,N_3986,N_3827);
or U4372 (N_4372,N_3784,N_3686);
nand U4373 (N_4373,N_3878,N_3717);
nand U4374 (N_4374,N_3935,N_3504);
nand U4375 (N_4375,N_3993,N_3799);
nand U4376 (N_4376,N_3593,N_3844);
nor U4377 (N_4377,N_3896,N_3899);
or U4378 (N_4378,N_3534,N_3948);
nor U4379 (N_4379,N_3894,N_3850);
and U4380 (N_4380,N_3590,N_3981);
or U4381 (N_4381,N_3711,N_3837);
nor U4382 (N_4382,N_3593,N_3739);
and U4383 (N_4383,N_3813,N_3950);
or U4384 (N_4384,N_3952,N_3841);
nor U4385 (N_4385,N_3738,N_3843);
or U4386 (N_4386,N_3976,N_3754);
nor U4387 (N_4387,N_3762,N_3944);
or U4388 (N_4388,N_3974,N_3528);
and U4389 (N_4389,N_3535,N_3700);
or U4390 (N_4390,N_3545,N_3584);
nor U4391 (N_4391,N_3528,N_3666);
or U4392 (N_4392,N_3533,N_3584);
or U4393 (N_4393,N_3626,N_3579);
and U4394 (N_4394,N_3603,N_3503);
and U4395 (N_4395,N_3804,N_3715);
or U4396 (N_4396,N_3641,N_3710);
nand U4397 (N_4397,N_3510,N_3796);
nand U4398 (N_4398,N_3902,N_3791);
or U4399 (N_4399,N_3687,N_3556);
and U4400 (N_4400,N_3876,N_3919);
or U4401 (N_4401,N_3552,N_3755);
nand U4402 (N_4402,N_3981,N_3831);
nor U4403 (N_4403,N_3673,N_3532);
nor U4404 (N_4404,N_3567,N_3767);
and U4405 (N_4405,N_3579,N_3568);
nand U4406 (N_4406,N_3785,N_3848);
nand U4407 (N_4407,N_3796,N_3900);
or U4408 (N_4408,N_3884,N_3567);
nand U4409 (N_4409,N_3745,N_3680);
nor U4410 (N_4410,N_3737,N_3586);
or U4411 (N_4411,N_3837,N_3619);
nor U4412 (N_4412,N_3940,N_3957);
and U4413 (N_4413,N_3611,N_3752);
xnor U4414 (N_4414,N_3537,N_3554);
and U4415 (N_4415,N_3937,N_3968);
or U4416 (N_4416,N_3974,N_3722);
xnor U4417 (N_4417,N_3939,N_3628);
xnor U4418 (N_4418,N_3987,N_3775);
nor U4419 (N_4419,N_3520,N_3861);
nand U4420 (N_4420,N_3983,N_3931);
nor U4421 (N_4421,N_3658,N_3938);
or U4422 (N_4422,N_3719,N_3951);
nand U4423 (N_4423,N_3501,N_3878);
nor U4424 (N_4424,N_3939,N_3946);
or U4425 (N_4425,N_3888,N_3654);
or U4426 (N_4426,N_3945,N_3908);
nand U4427 (N_4427,N_3580,N_3754);
nor U4428 (N_4428,N_3531,N_3780);
and U4429 (N_4429,N_3605,N_3685);
nor U4430 (N_4430,N_3536,N_3895);
or U4431 (N_4431,N_3632,N_3670);
and U4432 (N_4432,N_3924,N_3589);
and U4433 (N_4433,N_3636,N_3867);
nor U4434 (N_4434,N_3708,N_3524);
nor U4435 (N_4435,N_3869,N_3691);
or U4436 (N_4436,N_3993,N_3724);
nand U4437 (N_4437,N_3546,N_3890);
nand U4438 (N_4438,N_3506,N_3833);
nor U4439 (N_4439,N_3509,N_3562);
and U4440 (N_4440,N_3797,N_3698);
nor U4441 (N_4441,N_3546,N_3555);
nor U4442 (N_4442,N_3619,N_3647);
nor U4443 (N_4443,N_3585,N_3996);
or U4444 (N_4444,N_3939,N_3589);
or U4445 (N_4445,N_3508,N_3997);
and U4446 (N_4446,N_3611,N_3992);
and U4447 (N_4447,N_3887,N_3742);
nand U4448 (N_4448,N_3621,N_3655);
or U4449 (N_4449,N_3788,N_3762);
nand U4450 (N_4450,N_3782,N_3741);
or U4451 (N_4451,N_3673,N_3581);
nand U4452 (N_4452,N_3821,N_3844);
or U4453 (N_4453,N_3556,N_3969);
and U4454 (N_4454,N_3620,N_3883);
and U4455 (N_4455,N_3814,N_3781);
and U4456 (N_4456,N_3500,N_3753);
nor U4457 (N_4457,N_3684,N_3912);
nand U4458 (N_4458,N_3873,N_3595);
or U4459 (N_4459,N_3717,N_3574);
nor U4460 (N_4460,N_3849,N_3770);
or U4461 (N_4461,N_3532,N_3951);
nor U4462 (N_4462,N_3971,N_3806);
and U4463 (N_4463,N_3760,N_3580);
and U4464 (N_4464,N_3575,N_3622);
nand U4465 (N_4465,N_3986,N_3989);
nand U4466 (N_4466,N_3620,N_3678);
nor U4467 (N_4467,N_3950,N_3892);
nor U4468 (N_4468,N_3951,N_3955);
or U4469 (N_4469,N_3922,N_3702);
and U4470 (N_4470,N_3568,N_3502);
nand U4471 (N_4471,N_3720,N_3803);
and U4472 (N_4472,N_3546,N_3855);
nand U4473 (N_4473,N_3783,N_3761);
and U4474 (N_4474,N_3868,N_3857);
nand U4475 (N_4475,N_3969,N_3544);
or U4476 (N_4476,N_3521,N_3765);
xnor U4477 (N_4477,N_3566,N_3875);
nor U4478 (N_4478,N_3904,N_3894);
nor U4479 (N_4479,N_3825,N_3674);
and U4480 (N_4480,N_3873,N_3619);
nor U4481 (N_4481,N_3977,N_3625);
and U4482 (N_4482,N_3542,N_3831);
or U4483 (N_4483,N_3789,N_3541);
or U4484 (N_4484,N_3630,N_3861);
nor U4485 (N_4485,N_3935,N_3526);
nand U4486 (N_4486,N_3652,N_3568);
nand U4487 (N_4487,N_3973,N_3643);
nor U4488 (N_4488,N_3708,N_3768);
or U4489 (N_4489,N_3572,N_3855);
or U4490 (N_4490,N_3882,N_3823);
and U4491 (N_4491,N_3815,N_3591);
nor U4492 (N_4492,N_3519,N_3522);
nor U4493 (N_4493,N_3983,N_3525);
and U4494 (N_4494,N_3934,N_3615);
or U4495 (N_4495,N_3765,N_3527);
and U4496 (N_4496,N_3753,N_3742);
or U4497 (N_4497,N_3568,N_3800);
or U4498 (N_4498,N_3759,N_3568);
and U4499 (N_4499,N_3523,N_3509);
or U4500 (N_4500,N_4489,N_4391);
and U4501 (N_4501,N_4321,N_4298);
or U4502 (N_4502,N_4337,N_4451);
and U4503 (N_4503,N_4468,N_4294);
nand U4504 (N_4504,N_4223,N_4062);
nor U4505 (N_4505,N_4148,N_4410);
or U4506 (N_4506,N_4487,N_4003);
nand U4507 (N_4507,N_4393,N_4403);
nand U4508 (N_4508,N_4118,N_4089);
nor U4509 (N_4509,N_4137,N_4115);
or U4510 (N_4510,N_4280,N_4203);
nand U4511 (N_4511,N_4212,N_4225);
or U4512 (N_4512,N_4154,N_4078);
nand U4513 (N_4513,N_4344,N_4052);
nor U4514 (N_4514,N_4352,N_4098);
nand U4515 (N_4515,N_4422,N_4481);
and U4516 (N_4516,N_4301,N_4087);
and U4517 (N_4517,N_4017,N_4398);
and U4518 (N_4518,N_4260,N_4303);
or U4519 (N_4519,N_4354,N_4143);
and U4520 (N_4520,N_4176,N_4359);
and U4521 (N_4521,N_4379,N_4282);
nor U4522 (N_4522,N_4328,N_4082);
and U4523 (N_4523,N_4307,N_4112);
and U4524 (N_4524,N_4155,N_4267);
nor U4525 (N_4525,N_4306,N_4350);
nand U4526 (N_4526,N_4269,N_4404);
or U4527 (N_4527,N_4424,N_4497);
or U4528 (N_4528,N_4432,N_4185);
and U4529 (N_4529,N_4274,N_4139);
nor U4530 (N_4530,N_4334,N_4475);
and U4531 (N_4531,N_4129,N_4229);
nor U4532 (N_4532,N_4116,N_4132);
and U4533 (N_4533,N_4244,N_4057);
nor U4534 (N_4534,N_4317,N_4300);
or U4535 (N_4535,N_4006,N_4259);
nand U4536 (N_4536,N_4415,N_4073);
or U4537 (N_4537,N_4405,N_4462);
and U4538 (N_4538,N_4285,N_4210);
nor U4539 (N_4539,N_4341,N_4314);
nand U4540 (N_4540,N_4069,N_4195);
nand U4541 (N_4541,N_4053,N_4182);
or U4542 (N_4542,N_4316,N_4295);
or U4543 (N_4543,N_4136,N_4370);
and U4544 (N_4544,N_4079,N_4378);
nand U4545 (N_4545,N_4222,N_4390);
or U4546 (N_4546,N_4367,N_4252);
xor U4547 (N_4547,N_4320,N_4059);
nand U4548 (N_4548,N_4105,N_4077);
nand U4549 (N_4549,N_4254,N_4058);
or U4550 (N_4550,N_4327,N_4171);
nor U4551 (N_4551,N_4029,N_4331);
or U4552 (N_4552,N_4042,N_4189);
and U4553 (N_4553,N_4251,N_4455);
nand U4554 (N_4554,N_4375,N_4392);
and U4555 (N_4555,N_4117,N_4168);
xnor U4556 (N_4556,N_4031,N_4040);
nor U4557 (N_4557,N_4343,N_4308);
or U4558 (N_4558,N_4471,N_4369);
or U4559 (N_4559,N_4099,N_4499);
nand U4560 (N_4560,N_4091,N_4101);
nor U4561 (N_4561,N_4217,N_4479);
nand U4562 (N_4562,N_4239,N_4216);
or U4563 (N_4563,N_4094,N_4163);
nor U4564 (N_4564,N_4026,N_4281);
and U4565 (N_4565,N_4081,N_4243);
or U4566 (N_4566,N_4181,N_4414);
or U4567 (N_4567,N_4012,N_4202);
nor U4568 (N_4568,N_4355,N_4147);
nor U4569 (N_4569,N_4371,N_4402);
nor U4570 (N_4570,N_4289,N_4443);
or U4571 (N_4571,N_4149,N_4093);
nand U4572 (N_4572,N_4237,N_4450);
nor U4573 (N_4573,N_4262,N_4135);
nor U4574 (N_4574,N_4326,N_4278);
or U4575 (N_4575,N_4102,N_4111);
nand U4576 (N_4576,N_4299,N_4036);
xnor U4577 (N_4577,N_4448,N_4348);
nor U4578 (N_4578,N_4035,N_4399);
and U4579 (N_4579,N_4201,N_4151);
and U4580 (N_4580,N_4075,N_4454);
nor U4581 (N_4581,N_4275,N_4472);
nand U4582 (N_4582,N_4085,N_4109);
nor U4583 (N_4583,N_4213,N_4068);
nand U4584 (N_4584,N_4114,N_4047);
and U4585 (N_4585,N_4412,N_4240);
and U4586 (N_4586,N_4383,N_4256);
xor U4587 (N_4587,N_4146,N_4070);
and U4588 (N_4588,N_4054,N_4119);
and U4589 (N_4589,N_4442,N_4207);
nor U4590 (N_4590,N_4128,N_4048);
or U4591 (N_4591,N_4358,N_4276);
and U4592 (N_4592,N_4457,N_4257);
and U4593 (N_4593,N_4033,N_4236);
or U4594 (N_4594,N_4198,N_4486);
nand U4595 (N_4595,N_4142,N_4192);
or U4596 (N_4596,N_4156,N_4366);
or U4597 (N_4597,N_4473,N_4446);
xnor U4598 (N_4598,N_4064,N_4368);
nor U4599 (N_4599,N_4384,N_4041);
xor U4600 (N_4600,N_4365,N_4453);
nor U4601 (N_4601,N_4050,N_4034);
or U4602 (N_4602,N_4494,N_4286);
nand U4603 (N_4603,N_4437,N_4086);
and U4604 (N_4604,N_4123,N_4108);
or U4605 (N_4605,N_4401,N_4227);
or U4606 (N_4606,N_4090,N_4461);
and U4607 (N_4607,N_4152,N_4218);
nand U4608 (N_4608,N_4263,N_4178);
and U4609 (N_4609,N_4421,N_4339);
nor U4610 (N_4610,N_4413,N_4092);
and U4611 (N_4611,N_4196,N_4209);
nor U4612 (N_4612,N_4361,N_4433);
nand U4613 (N_4613,N_4083,N_4005);
nand U4614 (N_4614,N_4459,N_4490);
nand U4615 (N_4615,N_4253,N_4107);
and U4616 (N_4616,N_4397,N_4120);
nand U4617 (N_4617,N_4485,N_4046);
and U4618 (N_4618,N_4039,N_4418);
or U4619 (N_4619,N_4190,N_4138);
nor U4620 (N_4620,N_4018,N_4387);
or U4621 (N_4621,N_4394,N_4206);
or U4622 (N_4622,N_4283,N_4150);
nor U4623 (N_4623,N_4045,N_4325);
nor U4624 (N_4624,N_4215,N_4408);
nand U4625 (N_4625,N_4400,N_4221);
nand U4626 (N_4626,N_4103,N_4242);
nand U4627 (N_4627,N_4141,N_4228);
nand U4628 (N_4628,N_4312,N_4277);
and U4629 (N_4629,N_4356,N_4435);
and U4630 (N_4630,N_4084,N_4349);
or U4631 (N_4631,N_4467,N_4049);
or U4632 (N_4632,N_4066,N_4271);
and U4633 (N_4633,N_4194,N_4248);
or U4634 (N_4634,N_4330,N_4015);
or U4635 (N_4635,N_4346,N_4126);
and U4636 (N_4636,N_4157,N_4169);
nor U4637 (N_4637,N_4110,N_4296);
or U4638 (N_4638,N_4007,N_4191);
and U4639 (N_4639,N_4231,N_4342);
or U4640 (N_4640,N_4235,N_4420);
nor U4641 (N_4641,N_4363,N_4060);
nor U4642 (N_4642,N_4428,N_4024);
nor U4643 (N_4643,N_4357,N_4372);
nand U4644 (N_4644,N_4179,N_4373);
and U4645 (N_4645,N_4491,N_4161);
xor U4646 (N_4646,N_4456,N_4272);
and U4647 (N_4647,N_4279,N_4417);
nor U4648 (N_4648,N_4360,N_4332);
nand U4649 (N_4649,N_4051,N_4160);
or U4650 (N_4650,N_4106,N_4319);
nor U4651 (N_4651,N_4416,N_4291);
or U4652 (N_4652,N_4477,N_4095);
nand U4653 (N_4653,N_4449,N_4027);
or U4654 (N_4654,N_4465,N_4121);
nand U4655 (N_4655,N_4174,N_4480);
or U4656 (N_4656,N_4389,N_4322);
or U4657 (N_4657,N_4310,N_4019);
and U4658 (N_4658,N_4302,N_4021);
nor U4659 (N_4659,N_4199,N_4130);
or U4660 (N_4660,N_4407,N_4258);
or U4661 (N_4661,N_4311,N_4113);
nor U4662 (N_4662,N_4495,N_4436);
and U4663 (N_4663,N_4318,N_4340);
xnor U4664 (N_4664,N_4315,N_4385);
or U4665 (N_4665,N_4463,N_4043);
and U4666 (N_4666,N_4096,N_4388);
nor U4667 (N_4667,N_4376,N_4431);
xnor U4668 (N_4668,N_4484,N_4032);
nor U4669 (N_4669,N_4430,N_4288);
nor U4670 (N_4670,N_4447,N_4374);
nor U4671 (N_4671,N_4180,N_4028);
and U4672 (N_4672,N_4010,N_4232);
and U4673 (N_4673,N_4268,N_4020);
and U4674 (N_4674,N_4261,N_4464);
and U4675 (N_4675,N_4411,N_4297);
or U4676 (N_4676,N_4097,N_4014);
or U4677 (N_4677,N_4197,N_4234);
nand U4678 (N_4678,N_4406,N_4329);
or U4679 (N_4679,N_4226,N_4211);
nand U4680 (N_4680,N_4444,N_4336);
or U4681 (N_4681,N_4183,N_4466);
nor U4682 (N_4682,N_4438,N_4074);
nand U4683 (N_4683,N_4351,N_4347);
and U4684 (N_4684,N_4165,N_4122);
or U4685 (N_4685,N_4270,N_4381);
nor U4686 (N_4686,N_4233,N_4304);
or U4687 (N_4687,N_4309,N_4184);
and U4688 (N_4688,N_4247,N_4458);
nand U4689 (N_4689,N_4002,N_4063);
or U4690 (N_4690,N_4246,N_4044);
or U4691 (N_4691,N_4164,N_4364);
nor U4692 (N_4692,N_4476,N_4004);
and U4693 (N_4693,N_4153,N_4055);
nor U4694 (N_4694,N_4425,N_4145);
nand U4695 (N_4695,N_4395,N_4377);
or U4696 (N_4696,N_4439,N_4001);
nand U4697 (N_4697,N_4025,N_4441);
and U4698 (N_4698,N_4323,N_4345);
nand U4699 (N_4699,N_4460,N_4427);
or U4700 (N_4700,N_4162,N_4292);
nand U4701 (N_4701,N_4013,N_4186);
or U4702 (N_4702,N_4167,N_4219);
and U4703 (N_4703,N_4159,N_4238);
xor U4704 (N_4704,N_4305,N_4076);
or U4705 (N_4705,N_4488,N_4496);
xor U4706 (N_4706,N_4173,N_4200);
or U4707 (N_4707,N_4080,N_4293);
nor U4708 (N_4708,N_4474,N_4170);
nor U4709 (N_4709,N_4264,N_4250);
nor U4710 (N_4710,N_4030,N_4140);
nand U4711 (N_4711,N_4335,N_4224);
nand U4712 (N_4712,N_4088,N_4241);
nand U4713 (N_4713,N_4265,N_4125);
nor U4714 (N_4714,N_4067,N_4193);
nor U4715 (N_4715,N_4452,N_4172);
or U4716 (N_4716,N_4419,N_4426);
nand U4717 (N_4717,N_4000,N_4124);
nor U4718 (N_4718,N_4134,N_4144);
or U4719 (N_4719,N_4038,N_4287);
xnor U4720 (N_4720,N_4273,N_4208);
or U4721 (N_4721,N_4290,N_4470);
nor U4722 (N_4722,N_4266,N_4333);
and U4723 (N_4723,N_4061,N_4008);
nor U4724 (N_4724,N_4440,N_4423);
and U4725 (N_4725,N_4127,N_4284);
nand U4726 (N_4726,N_4492,N_4056);
or U4727 (N_4727,N_4022,N_4023);
nor U4728 (N_4728,N_4133,N_4409);
nor U4729 (N_4729,N_4382,N_4434);
nor U4730 (N_4730,N_4429,N_4204);
or U4731 (N_4731,N_4037,N_4187);
or U4732 (N_4732,N_4249,N_4478);
nor U4733 (N_4733,N_4483,N_4188);
and U4734 (N_4734,N_4482,N_4071);
nand U4735 (N_4735,N_4362,N_4396);
and U4736 (N_4736,N_4245,N_4177);
nand U4737 (N_4737,N_4016,N_4255);
nand U4738 (N_4738,N_4100,N_4445);
nor U4739 (N_4739,N_4324,N_4230);
nor U4740 (N_4740,N_4065,N_4009);
nor U4741 (N_4741,N_4158,N_4214);
nand U4742 (N_4742,N_4386,N_4011);
nor U4743 (N_4743,N_4338,N_4205);
nand U4744 (N_4744,N_4220,N_4380);
or U4745 (N_4745,N_4469,N_4353);
or U4746 (N_4746,N_4175,N_4072);
or U4747 (N_4747,N_4498,N_4166);
nand U4748 (N_4748,N_4493,N_4131);
or U4749 (N_4749,N_4104,N_4313);
nor U4750 (N_4750,N_4244,N_4432);
or U4751 (N_4751,N_4004,N_4315);
or U4752 (N_4752,N_4099,N_4078);
nand U4753 (N_4753,N_4384,N_4292);
nor U4754 (N_4754,N_4376,N_4211);
nand U4755 (N_4755,N_4114,N_4339);
and U4756 (N_4756,N_4315,N_4189);
or U4757 (N_4757,N_4061,N_4206);
nor U4758 (N_4758,N_4269,N_4202);
nor U4759 (N_4759,N_4224,N_4372);
or U4760 (N_4760,N_4199,N_4054);
nor U4761 (N_4761,N_4010,N_4157);
nand U4762 (N_4762,N_4074,N_4422);
or U4763 (N_4763,N_4144,N_4274);
nand U4764 (N_4764,N_4313,N_4059);
nor U4765 (N_4765,N_4029,N_4321);
or U4766 (N_4766,N_4026,N_4235);
and U4767 (N_4767,N_4422,N_4381);
and U4768 (N_4768,N_4102,N_4495);
and U4769 (N_4769,N_4413,N_4000);
nor U4770 (N_4770,N_4453,N_4004);
xnor U4771 (N_4771,N_4442,N_4157);
or U4772 (N_4772,N_4089,N_4204);
nand U4773 (N_4773,N_4312,N_4470);
nand U4774 (N_4774,N_4412,N_4417);
and U4775 (N_4775,N_4047,N_4406);
nor U4776 (N_4776,N_4155,N_4426);
nand U4777 (N_4777,N_4407,N_4499);
or U4778 (N_4778,N_4352,N_4466);
nand U4779 (N_4779,N_4013,N_4343);
and U4780 (N_4780,N_4336,N_4330);
and U4781 (N_4781,N_4181,N_4437);
or U4782 (N_4782,N_4117,N_4006);
or U4783 (N_4783,N_4081,N_4248);
nand U4784 (N_4784,N_4228,N_4464);
and U4785 (N_4785,N_4380,N_4458);
or U4786 (N_4786,N_4066,N_4362);
and U4787 (N_4787,N_4130,N_4164);
nand U4788 (N_4788,N_4046,N_4118);
and U4789 (N_4789,N_4350,N_4421);
nand U4790 (N_4790,N_4226,N_4360);
or U4791 (N_4791,N_4017,N_4291);
nand U4792 (N_4792,N_4266,N_4429);
and U4793 (N_4793,N_4442,N_4391);
or U4794 (N_4794,N_4244,N_4106);
and U4795 (N_4795,N_4337,N_4447);
and U4796 (N_4796,N_4164,N_4491);
xnor U4797 (N_4797,N_4449,N_4026);
and U4798 (N_4798,N_4333,N_4216);
or U4799 (N_4799,N_4046,N_4116);
nor U4800 (N_4800,N_4037,N_4460);
or U4801 (N_4801,N_4254,N_4188);
nand U4802 (N_4802,N_4364,N_4380);
and U4803 (N_4803,N_4295,N_4458);
and U4804 (N_4804,N_4444,N_4055);
or U4805 (N_4805,N_4250,N_4342);
or U4806 (N_4806,N_4117,N_4299);
and U4807 (N_4807,N_4007,N_4181);
nand U4808 (N_4808,N_4238,N_4279);
or U4809 (N_4809,N_4204,N_4154);
nand U4810 (N_4810,N_4181,N_4271);
nor U4811 (N_4811,N_4449,N_4231);
nor U4812 (N_4812,N_4369,N_4040);
nor U4813 (N_4813,N_4084,N_4009);
or U4814 (N_4814,N_4152,N_4111);
or U4815 (N_4815,N_4336,N_4109);
and U4816 (N_4816,N_4487,N_4142);
and U4817 (N_4817,N_4386,N_4188);
nor U4818 (N_4818,N_4331,N_4417);
nand U4819 (N_4819,N_4402,N_4304);
or U4820 (N_4820,N_4305,N_4057);
and U4821 (N_4821,N_4352,N_4203);
or U4822 (N_4822,N_4379,N_4291);
or U4823 (N_4823,N_4436,N_4345);
and U4824 (N_4824,N_4231,N_4093);
nor U4825 (N_4825,N_4297,N_4462);
nand U4826 (N_4826,N_4451,N_4496);
nand U4827 (N_4827,N_4279,N_4452);
or U4828 (N_4828,N_4236,N_4431);
or U4829 (N_4829,N_4243,N_4383);
nor U4830 (N_4830,N_4147,N_4281);
or U4831 (N_4831,N_4361,N_4338);
or U4832 (N_4832,N_4155,N_4079);
nor U4833 (N_4833,N_4443,N_4002);
xor U4834 (N_4834,N_4212,N_4415);
nand U4835 (N_4835,N_4062,N_4479);
nand U4836 (N_4836,N_4382,N_4116);
nand U4837 (N_4837,N_4228,N_4445);
and U4838 (N_4838,N_4104,N_4466);
or U4839 (N_4839,N_4343,N_4074);
and U4840 (N_4840,N_4113,N_4457);
or U4841 (N_4841,N_4193,N_4217);
and U4842 (N_4842,N_4195,N_4178);
nor U4843 (N_4843,N_4327,N_4249);
nand U4844 (N_4844,N_4075,N_4401);
nor U4845 (N_4845,N_4412,N_4155);
xor U4846 (N_4846,N_4120,N_4468);
nor U4847 (N_4847,N_4465,N_4020);
nand U4848 (N_4848,N_4489,N_4086);
nor U4849 (N_4849,N_4071,N_4247);
and U4850 (N_4850,N_4083,N_4202);
nand U4851 (N_4851,N_4123,N_4346);
and U4852 (N_4852,N_4390,N_4395);
nand U4853 (N_4853,N_4285,N_4010);
and U4854 (N_4854,N_4399,N_4338);
or U4855 (N_4855,N_4272,N_4127);
nand U4856 (N_4856,N_4415,N_4026);
nand U4857 (N_4857,N_4452,N_4164);
or U4858 (N_4858,N_4499,N_4210);
nand U4859 (N_4859,N_4077,N_4326);
nand U4860 (N_4860,N_4006,N_4284);
nor U4861 (N_4861,N_4093,N_4345);
nand U4862 (N_4862,N_4477,N_4300);
nor U4863 (N_4863,N_4458,N_4028);
nand U4864 (N_4864,N_4476,N_4207);
nor U4865 (N_4865,N_4417,N_4117);
and U4866 (N_4866,N_4391,N_4387);
nor U4867 (N_4867,N_4364,N_4245);
or U4868 (N_4868,N_4254,N_4416);
and U4869 (N_4869,N_4153,N_4010);
or U4870 (N_4870,N_4010,N_4175);
nor U4871 (N_4871,N_4489,N_4290);
nor U4872 (N_4872,N_4419,N_4445);
and U4873 (N_4873,N_4261,N_4282);
nand U4874 (N_4874,N_4187,N_4168);
nor U4875 (N_4875,N_4193,N_4454);
and U4876 (N_4876,N_4033,N_4085);
or U4877 (N_4877,N_4234,N_4185);
or U4878 (N_4878,N_4022,N_4391);
and U4879 (N_4879,N_4262,N_4250);
nor U4880 (N_4880,N_4158,N_4482);
and U4881 (N_4881,N_4047,N_4011);
or U4882 (N_4882,N_4335,N_4443);
and U4883 (N_4883,N_4181,N_4048);
nand U4884 (N_4884,N_4176,N_4389);
nand U4885 (N_4885,N_4458,N_4066);
and U4886 (N_4886,N_4240,N_4127);
or U4887 (N_4887,N_4333,N_4374);
or U4888 (N_4888,N_4408,N_4081);
or U4889 (N_4889,N_4191,N_4097);
nor U4890 (N_4890,N_4290,N_4219);
and U4891 (N_4891,N_4147,N_4403);
nor U4892 (N_4892,N_4086,N_4045);
nand U4893 (N_4893,N_4124,N_4227);
and U4894 (N_4894,N_4426,N_4485);
nor U4895 (N_4895,N_4076,N_4339);
and U4896 (N_4896,N_4370,N_4358);
or U4897 (N_4897,N_4352,N_4057);
and U4898 (N_4898,N_4116,N_4492);
or U4899 (N_4899,N_4491,N_4482);
or U4900 (N_4900,N_4039,N_4014);
and U4901 (N_4901,N_4026,N_4400);
nor U4902 (N_4902,N_4160,N_4423);
or U4903 (N_4903,N_4246,N_4355);
nor U4904 (N_4904,N_4449,N_4294);
and U4905 (N_4905,N_4274,N_4183);
xor U4906 (N_4906,N_4234,N_4473);
and U4907 (N_4907,N_4181,N_4183);
or U4908 (N_4908,N_4461,N_4302);
xor U4909 (N_4909,N_4074,N_4044);
or U4910 (N_4910,N_4292,N_4114);
and U4911 (N_4911,N_4030,N_4412);
nor U4912 (N_4912,N_4458,N_4016);
and U4913 (N_4913,N_4160,N_4480);
nand U4914 (N_4914,N_4028,N_4438);
xor U4915 (N_4915,N_4266,N_4477);
nand U4916 (N_4916,N_4070,N_4264);
nor U4917 (N_4917,N_4001,N_4316);
nand U4918 (N_4918,N_4387,N_4228);
nor U4919 (N_4919,N_4276,N_4280);
and U4920 (N_4920,N_4456,N_4411);
nor U4921 (N_4921,N_4441,N_4328);
or U4922 (N_4922,N_4012,N_4477);
or U4923 (N_4923,N_4252,N_4156);
or U4924 (N_4924,N_4349,N_4273);
and U4925 (N_4925,N_4344,N_4250);
and U4926 (N_4926,N_4409,N_4250);
and U4927 (N_4927,N_4155,N_4052);
or U4928 (N_4928,N_4241,N_4397);
nor U4929 (N_4929,N_4411,N_4038);
and U4930 (N_4930,N_4440,N_4353);
and U4931 (N_4931,N_4396,N_4077);
nor U4932 (N_4932,N_4216,N_4214);
or U4933 (N_4933,N_4135,N_4326);
or U4934 (N_4934,N_4006,N_4001);
nand U4935 (N_4935,N_4231,N_4401);
nand U4936 (N_4936,N_4415,N_4065);
nand U4937 (N_4937,N_4152,N_4184);
nand U4938 (N_4938,N_4017,N_4317);
nor U4939 (N_4939,N_4097,N_4021);
nand U4940 (N_4940,N_4117,N_4318);
nand U4941 (N_4941,N_4464,N_4104);
xnor U4942 (N_4942,N_4281,N_4003);
or U4943 (N_4943,N_4316,N_4273);
and U4944 (N_4944,N_4381,N_4340);
or U4945 (N_4945,N_4362,N_4097);
and U4946 (N_4946,N_4052,N_4137);
nor U4947 (N_4947,N_4297,N_4325);
nand U4948 (N_4948,N_4188,N_4271);
nand U4949 (N_4949,N_4119,N_4452);
nand U4950 (N_4950,N_4402,N_4399);
nand U4951 (N_4951,N_4438,N_4337);
or U4952 (N_4952,N_4221,N_4466);
or U4953 (N_4953,N_4280,N_4251);
or U4954 (N_4954,N_4263,N_4340);
and U4955 (N_4955,N_4364,N_4318);
xor U4956 (N_4956,N_4070,N_4293);
or U4957 (N_4957,N_4244,N_4478);
nand U4958 (N_4958,N_4078,N_4251);
or U4959 (N_4959,N_4387,N_4311);
nand U4960 (N_4960,N_4456,N_4437);
nand U4961 (N_4961,N_4097,N_4410);
or U4962 (N_4962,N_4459,N_4103);
nand U4963 (N_4963,N_4053,N_4317);
or U4964 (N_4964,N_4214,N_4367);
or U4965 (N_4965,N_4179,N_4438);
and U4966 (N_4966,N_4444,N_4032);
or U4967 (N_4967,N_4092,N_4184);
nor U4968 (N_4968,N_4002,N_4022);
and U4969 (N_4969,N_4439,N_4327);
and U4970 (N_4970,N_4233,N_4235);
nor U4971 (N_4971,N_4214,N_4172);
nand U4972 (N_4972,N_4184,N_4082);
and U4973 (N_4973,N_4110,N_4479);
or U4974 (N_4974,N_4317,N_4411);
or U4975 (N_4975,N_4348,N_4231);
xnor U4976 (N_4976,N_4370,N_4070);
or U4977 (N_4977,N_4390,N_4210);
and U4978 (N_4978,N_4040,N_4362);
or U4979 (N_4979,N_4492,N_4007);
nand U4980 (N_4980,N_4354,N_4133);
nand U4981 (N_4981,N_4249,N_4264);
nor U4982 (N_4982,N_4156,N_4055);
or U4983 (N_4983,N_4231,N_4121);
and U4984 (N_4984,N_4143,N_4023);
or U4985 (N_4985,N_4228,N_4099);
nand U4986 (N_4986,N_4294,N_4254);
nand U4987 (N_4987,N_4065,N_4159);
and U4988 (N_4988,N_4218,N_4497);
and U4989 (N_4989,N_4309,N_4315);
nand U4990 (N_4990,N_4499,N_4317);
nor U4991 (N_4991,N_4118,N_4318);
and U4992 (N_4992,N_4274,N_4020);
nor U4993 (N_4993,N_4489,N_4446);
nand U4994 (N_4994,N_4058,N_4172);
nand U4995 (N_4995,N_4428,N_4069);
and U4996 (N_4996,N_4133,N_4079);
and U4997 (N_4997,N_4275,N_4098);
nand U4998 (N_4998,N_4497,N_4434);
and U4999 (N_4999,N_4101,N_4046);
nand U5000 (N_5000,N_4931,N_4619);
and U5001 (N_5001,N_4653,N_4906);
nor U5002 (N_5002,N_4613,N_4783);
or U5003 (N_5003,N_4511,N_4868);
nor U5004 (N_5004,N_4776,N_4763);
xnor U5005 (N_5005,N_4567,N_4647);
xnor U5006 (N_5006,N_4862,N_4750);
nand U5007 (N_5007,N_4688,N_4893);
nand U5008 (N_5008,N_4724,N_4822);
nand U5009 (N_5009,N_4861,N_4630);
and U5010 (N_5010,N_4690,N_4627);
or U5011 (N_5011,N_4741,N_4850);
nor U5012 (N_5012,N_4744,N_4795);
nor U5013 (N_5013,N_4569,N_4594);
nand U5014 (N_5014,N_4814,N_4896);
nand U5015 (N_5015,N_4932,N_4779);
nor U5016 (N_5016,N_4887,N_4946);
and U5017 (N_5017,N_4778,N_4948);
or U5018 (N_5018,N_4919,N_4823);
and U5019 (N_5019,N_4908,N_4642);
or U5020 (N_5020,N_4599,N_4758);
nand U5021 (N_5021,N_4677,N_4928);
nand U5022 (N_5022,N_4969,N_4798);
nor U5023 (N_5023,N_4657,N_4675);
nand U5024 (N_5024,N_4501,N_4623);
and U5025 (N_5025,N_4863,N_4894);
and U5026 (N_5026,N_4915,N_4835);
or U5027 (N_5027,N_4713,N_4684);
and U5028 (N_5028,N_4914,N_4582);
and U5029 (N_5029,N_4535,N_4517);
or U5030 (N_5030,N_4890,N_4526);
or U5031 (N_5031,N_4571,N_4748);
nor U5032 (N_5032,N_4612,N_4691);
nand U5033 (N_5033,N_4658,N_4864);
or U5034 (N_5034,N_4572,N_4838);
or U5035 (N_5035,N_4837,N_4704);
nor U5036 (N_5036,N_4707,N_4885);
nor U5037 (N_5037,N_4920,N_4829);
and U5038 (N_5038,N_4955,N_4602);
or U5039 (N_5039,N_4686,N_4762);
nand U5040 (N_5040,N_4929,N_4570);
nor U5041 (N_5041,N_4905,N_4548);
or U5042 (N_5042,N_4631,N_4502);
nand U5043 (N_5043,N_4553,N_4626);
and U5044 (N_5044,N_4967,N_4769);
nor U5045 (N_5045,N_4510,N_4655);
and U5046 (N_5046,N_4891,N_4976);
and U5047 (N_5047,N_4869,N_4678);
xnor U5048 (N_5048,N_4696,N_4557);
nand U5049 (N_5049,N_4938,N_4767);
or U5050 (N_5050,N_4895,N_4555);
nor U5051 (N_5051,N_4656,N_4811);
and U5052 (N_5052,N_4785,N_4537);
nand U5053 (N_5053,N_4968,N_4760);
and U5054 (N_5054,N_4827,N_4951);
nand U5055 (N_5055,N_4560,N_4710);
nand U5056 (N_5056,N_4958,N_4939);
or U5057 (N_5057,N_4576,N_4563);
xor U5058 (N_5058,N_4705,N_4680);
nand U5059 (N_5059,N_4789,N_4826);
and U5060 (N_5060,N_4971,N_4923);
nand U5061 (N_5061,N_4585,N_4756);
nand U5062 (N_5062,N_4803,N_4670);
nor U5063 (N_5063,N_4574,N_4935);
and U5064 (N_5064,N_4679,N_4947);
or U5065 (N_5065,N_4669,N_4733);
nor U5066 (N_5066,N_4745,N_4717);
xnor U5067 (N_5067,N_4739,N_4834);
nor U5068 (N_5068,N_4614,N_4721);
nor U5069 (N_5069,N_4638,N_4839);
or U5070 (N_5070,N_4963,N_4892);
or U5071 (N_5071,N_4729,N_4852);
nand U5072 (N_5072,N_4853,N_4978);
or U5073 (N_5073,N_4727,N_4715);
nand U5074 (N_5074,N_4792,N_4924);
and U5075 (N_5075,N_4970,N_4743);
and U5076 (N_5076,N_4507,N_4749);
or U5077 (N_5077,N_4546,N_4771);
and U5078 (N_5078,N_4747,N_4842);
nand U5079 (N_5079,N_4708,N_4793);
nor U5080 (N_5080,N_4554,N_4505);
nand U5081 (N_5081,N_4768,N_4556);
or U5082 (N_5082,N_4661,N_4595);
or U5083 (N_5083,N_4525,N_4573);
or U5084 (N_5084,N_4818,N_4590);
nor U5085 (N_5085,N_4592,N_4995);
nor U5086 (N_5086,N_4873,N_4695);
nand U5087 (N_5087,N_4722,N_4580);
or U5088 (N_5088,N_4797,N_4866);
nand U5089 (N_5089,N_4752,N_4941);
nand U5090 (N_5090,N_4990,N_4728);
and U5091 (N_5091,N_4565,N_4987);
and U5092 (N_5092,N_4693,N_4854);
or U5093 (N_5093,N_4828,N_4980);
nand U5094 (N_5094,N_4731,N_4791);
nand U5095 (N_5095,N_4593,N_4874);
or U5096 (N_5096,N_4662,N_4520);
and U5097 (N_5097,N_4966,N_4732);
and U5098 (N_5098,N_4819,N_4506);
or U5099 (N_5099,N_4983,N_4687);
nor U5100 (N_5100,N_4660,N_4579);
nand U5101 (N_5101,N_4876,N_4530);
nor U5102 (N_5102,N_4843,N_4904);
nor U5103 (N_5103,N_4694,N_4622);
xor U5104 (N_5104,N_4782,N_4856);
or U5105 (N_5105,N_4558,N_4667);
nand U5106 (N_5106,N_4886,N_4637);
or U5107 (N_5107,N_4700,N_4897);
nor U5108 (N_5108,N_4940,N_4956);
or U5109 (N_5109,N_4954,N_4755);
nand U5110 (N_5110,N_4531,N_4529);
and U5111 (N_5111,N_4641,N_4651);
nor U5112 (N_5112,N_4588,N_4907);
nor U5113 (N_5113,N_4740,N_4830);
and U5114 (N_5114,N_4999,N_4877);
nand U5115 (N_5115,N_4964,N_4512);
and U5116 (N_5116,N_4672,N_4735);
or U5117 (N_5117,N_4784,N_4539);
nor U5118 (N_5118,N_4836,N_4504);
and U5119 (N_5119,N_4532,N_4857);
nor U5120 (N_5120,N_4977,N_4833);
and U5121 (N_5121,N_4881,N_4764);
nor U5122 (N_5122,N_4581,N_4550);
nor U5123 (N_5123,N_4766,N_4591);
nand U5124 (N_5124,N_4577,N_4847);
and U5125 (N_5125,N_4518,N_4902);
nor U5126 (N_5126,N_4816,N_4682);
or U5127 (N_5127,N_4543,N_4773);
and U5128 (N_5128,N_4761,N_4736);
nor U5129 (N_5129,N_4878,N_4536);
or U5130 (N_5130,N_4988,N_4889);
and U5131 (N_5131,N_4775,N_4746);
nand U5132 (N_5132,N_4986,N_4701);
nand U5133 (N_5133,N_4945,N_4930);
nor U5134 (N_5134,N_4800,N_4806);
or U5135 (N_5135,N_4934,N_4676);
and U5136 (N_5136,N_4975,N_4730);
nor U5137 (N_5137,N_4711,N_4703);
nand U5138 (N_5138,N_4809,N_4960);
nand U5139 (N_5139,N_4604,N_4824);
nand U5140 (N_5140,N_4673,N_4805);
and U5141 (N_5141,N_4596,N_4645);
and U5142 (N_5142,N_4551,N_4522);
nand U5143 (N_5143,N_4719,N_4858);
nor U5144 (N_5144,N_4888,N_4855);
nand U5145 (N_5145,N_4926,N_4772);
nor U5146 (N_5146,N_4668,N_4547);
or U5147 (N_5147,N_4807,N_4982);
nor U5148 (N_5148,N_4916,N_4706);
nor U5149 (N_5149,N_4568,N_4561);
nor U5150 (N_5150,N_4949,N_4562);
and U5151 (N_5151,N_4911,N_4950);
and U5152 (N_5152,N_4759,N_4903);
and U5153 (N_5153,N_4608,N_4742);
nor U5154 (N_5154,N_4624,N_4559);
nor U5155 (N_5155,N_4870,N_4996);
nor U5156 (N_5156,N_4720,N_4544);
nor U5157 (N_5157,N_4654,N_4566);
and U5158 (N_5158,N_4846,N_4712);
nor U5159 (N_5159,N_4610,N_4664);
nand U5160 (N_5160,N_4629,N_4639);
and U5161 (N_5161,N_4821,N_4528);
and U5162 (N_5162,N_4882,N_4871);
or U5163 (N_5163,N_4867,N_4880);
nand U5164 (N_5164,N_4605,N_4578);
nor U5165 (N_5165,N_4523,N_4817);
or U5166 (N_5166,N_4663,N_4674);
nor U5167 (N_5167,N_4698,N_4985);
nand U5168 (N_5168,N_4848,N_4671);
or U5169 (N_5169,N_4564,N_4992);
and U5170 (N_5170,N_4552,N_4757);
nor U5171 (N_5171,N_4685,N_4597);
nand U5172 (N_5172,N_4944,N_4974);
nor U5173 (N_5173,N_4937,N_4633);
and U5174 (N_5174,N_4734,N_4840);
nand U5175 (N_5175,N_4628,N_4503);
xnor U5176 (N_5176,N_4514,N_4508);
or U5177 (N_5177,N_4575,N_4636);
and U5178 (N_5178,N_4860,N_4617);
or U5179 (N_5179,N_4865,N_4709);
or U5180 (N_5180,N_4692,N_4898);
nor U5181 (N_5181,N_4632,N_4618);
nor U5182 (N_5182,N_4603,N_4899);
or U5183 (N_5183,N_4957,N_4917);
nand U5184 (N_5184,N_4689,N_4943);
nor U5185 (N_5185,N_4927,N_4790);
nand U5186 (N_5186,N_4513,N_4786);
nand U5187 (N_5187,N_4774,N_4936);
or U5188 (N_5188,N_4723,N_4925);
nor U5189 (N_5189,N_4545,N_4804);
or U5190 (N_5190,N_4900,N_4584);
nand U5191 (N_5191,N_4962,N_4516);
nor U5192 (N_5192,N_4549,N_4859);
nand U5193 (N_5193,N_4991,N_4737);
nor U5194 (N_5194,N_4781,N_4831);
nand U5195 (N_5195,N_4601,N_4646);
nor U5196 (N_5196,N_4598,N_4820);
and U5197 (N_5197,N_4600,N_4611);
and U5198 (N_5198,N_4787,N_4972);
and U5199 (N_5199,N_4910,N_4918);
nor U5200 (N_5200,N_4524,N_4810);
and U5201 (N_5201,N_4659,N_4616);
and U5202 (N_5202,N_4912,N_4796);
or U5203 (N_5203,N_4714,N_4515);
and U5204 (N_5204,N_4812,N_4961);
nor U5205 (N_5205,N_4500,N_4725);
and U5206 (N_5206,N_4875,N_4583);
and U5207 (N_5207,N_4542,N_4994);
and U5208 (N_5208,N_4794,N_4521);
or U5209 (N_5209,N_4665,N_4620);
nand U5210 (N_5210,N_4716,N_4952);
nand U5211 (N_5211,N_4979,N_4799);
or U5212 (N_5212,N_4883,N_4699);
nor U5213 (N_5213,N_4738,N_4589);
or U5214 (N_5214,N_4998,N_4801);
nor U5215 (N_5215,N_4993,N_4649);
and U5216 (N_5216,N_4634,N_4644);
nand U5217 (N_5217,N_4997,N_4640);
and U5218 (N_5218,N_4533,N_4884);
or U5219 (N_5219,N_4849,N_4879);
and U5220 (N_5220,N_4702,N_4625);
and U5221 (N_5221,N_4765,N_4650);
nand U5222 (N_5222,N_4540,N_4984);
nor U5223 (N_5223,N_4942,N_4753);
xor U5224 (N_5224,N_4538,N_4770);
or U5225 (N_5225,N_4519,N_4606);
and U5226 (N_5226,N_4901,N_4802);
nor U5227 (N_5227,N_4652,N_4953);
nand U5228 (N_5228,N_4586,N_4643);
nor U5229 (N_5229,N_4754,N_4973);
nand U5230 (N_5230,N_4909,N_4621);
nand U5231 (N_5231,N_4913,N_4815);
and U5232 (N_5232,N_4527,N_4751);
nor U5233 (N_5233,N_4989,N_4780);
nor U5234 (N_5234,N_4825,N_4541);
nor U5235 (N_5235,N_4922,N_4718);
nand U5236 (N_5236,N_4832,N_4609);
nand U5237 (N_5237,N_4509,N_4648);
nor U5238 (N_5238,N_4788,N_4808);
nor U5239 (N_5239,N_4681,N_4933);
xnor U5240 (N_5240,N_4965,N_4697);
or U5241 (N_5241,N_4666,N_4813);
nand U5242 (N_5242,N_4587,N_4534);
and U5243 (N_5243,N_4726,N_4607);
or U5244 (N_5244,N_4981,N_4683);
nor U5245 (N_5245,N_4777,N_4921);
xor U5246 (N_5246,N_4841,N_4844);
or U5247 (N_5247,N_4851,N_4845);
nand U5248 (N_5248,N_4959,N_4615);
or U5249 (N_5249,N_4872,N_4635);
or U5250 (N_5250,N_4783,N_4902);
nand U5251 (N_5251,N_4801,N_4946);
and U5252 (N_5252,N_4857,N_4998);
nor U5253 (N_5253,N_4872,N_4860);
nor U5254 (N_5254,N_4820,N_4624);
nor U5255 (N_5255,N_4573,N_4628);
and U5256 (N_5256,N_4620,N_4608);
nor U5257 (N_5257,N_4516,N_4528);
nor U5258 (N_5258,N_4501,N_4759);
or U5259 (N_5259,N_4709,N_4647);
nand U5260 (N_5260,N_4575,N_4517);
nor U5261 (N_5261,N_4793,N_4565);
nand U5262 (N_5262,N_4754,N_4779);
nor U5263 (N_5263,N_4894,N_4746);
and U5264 (N_5264,N_4589,N_4754);
and U5265 (N_5265,N_4820,N_4945);
and U5266 (N_5266,N_4740,N_4848);
and U5267 (N_5267,N_4816,N_4832);
and U5268 (N_5268,N_4751,N_4941);
xor U5269 (N_5269,N_4889,N_4829);
or U5270 (N_5270,N_4864,N_4500);
and U5271 (N_5271,N_4612,N_4693);
nor U5272 (N_5272,N_4588,N_4901);
and U5273 (N_5273,N_4836,N_4823);
nor U5274 (N_5274,N_4975,N_4608);
or U5275 (N_5275,N_4765,N_4802);
nor U5276 (N_5276,N_4789,N_4948);
or U5277 (N_5277,N_4661,N_4930);
or U5278 (N_5278,N_4812,N_4789);
nand U5279 (N_5279,N_4699,N_4832);
or U5280 (N_5280,N_4589,N_4783);
nor U5281 (N_5281,N_4697,N_4583);
nand U5282 (N_5282,N_4935,N_4997);
nor U5283 (N_5283,N_4692,N_4767);
nor U5284 (N_5284,N_4804,N_4922);
nand U5285 (N_5285,N_4639,N_4807);
and U5286 (N_5286,N_4530,N_4717);
or U5287 (N_5287,N_4709,N_4785);
or U5288 (N_5288,N_4634,N_4872);
nand U5289 (N_5289,N_4549,N_4997);
nor U5290 (N_5290,N_4556,N_4875);
nor U5291 (N_5291,N_4831,N_4837);
or U5292 (N_5292,N_4985,N_4785);
and U5293 (N_5293,N_4994,N_4792);
and U5294 (N_5294,N_4514,N_4589);
nor U5295 (N_5295,N_4658,N_4714);
nor U5296 (N_5296,N_4716,N_4628);
and U5297 (N_5297,N_4992,N_4756);
xor U5298 (N_5298,N_4936,N_4573);
nor U5299 (N_5299,N_4863,N_4677);
nand U5300 (N_5300,N_4948,N_4655);
or U5301 (N_5301,N_4780,N_4810);
or U5302 (N_5302,N_4890,N_4912);
nand U5303 (N_5303,N_4799,N_4817);
and U5304 (N_5304,N_4529,N_4606);
or U5305 (N_5305,N_4679,N_4579);
xor U5306 (N_5306,N_4678,N_4709);
and U5307 (N_5307,N_4712,N_4601);
nor U5308 (N_5308,N_4630,N_4517);
and U5309 (N_5309,N_4937,N_4592);
or U5310 (N_5310,N_4765,N_4652);
nor U5311 (N_5311,N_4762,N_4966);
nand U5312 (N_5312,N_4802,N_4650);
nand U5313 (N_5313,N_4948,N_4943);
xnor U5314 (N_5314,N_4772,N_4510);
xor U5315 (N_5315,N_4706,N_4694);
nor U5316 (N_5316,N_4743,N_4851);
nor U5317 (N_5317,N_4975,N_4668);
and U5318 (N_5318,N_4792,N_4732);
or U5319 (N_5319,N_4662,N_4929);
nand U5320 (N_5320,N_4920,N_4506);
and U5321 (N_5321,N_4794,N_4849);
or U5322 (N_5322,N_4884,N_4583);
nand U5323 (N_5323,N_4788,N_4816);
nor U5324 (N_5324,N_4928,N_4909);
nand U5325 (N_5325,N_4518,N_4997);
xor U5326 (N_5326,N_4723,N_4828);
and U5327 (N_5327,N_4651,N_4753);
nor U5328 (N_5328,N_4545,N_4590);
or U5329 (N_5329,N_4506,N_4935);
and U5330 (N_5330,N_4844,N_4683);
nor U5331 (N_5331,N_4642,N_4851);
nand U5332 (N_5332,N_4989,N_4760);
nor U5333 (N_5333,N_4977,N_4597);
nor U5334 (N_5334,N_4855,N_4550);
nand U5335 (N_5335,N_4529,N_4660);
and U5336 (N_5336,N_4920,N_4683);
and U5337 (N_5337,N_4931,N_4692);
nand U5338 (N_5338,N_4887,N_4860);
or U5339 (N_5339,N_4614,N_4529);
and U5340 (N_5340,N_4885,N_4584);
nand U5341 (N_5341,N_4563,N_4812);
or U5342 (N_5342,N_4565,N_4685);
and U5343 (N_5343,N_4936,N_4505);
nor U5344 (N_5344,N_4797,N_4736);
nor U5345 (N_5345,N_4687,N_4513);
and U5346 (N_5346,N_4928,N_4791);
and U5347 (N_5347,N_4987,N_4657);
or U5348 (N_5348,N_4652,N_4846);
and U5349 (N_5349,N_4975,N_4708);
nand U5350 (N_5350,N_4690,N_4825);
nor U5351 (N_5351,N_4814,N_4783);
and U5352 (N_5352,N_4577,N_4571);
nor U5353 (N_5353,N_4607,N_4839);
and U5354 (N_5354,N_4920,N_4958);
or U5355 (N_5355,N_4914,N_4769);
nor U5356 (N_5356,N_4946,N_4587);
nand U5357 (N_5357,N_4606,N_4823);
and U5358 (N_5358,N_4968,N_4849);
nor U5359 (N_5359,N_4963,N_4940);
or U5360 (N_5360,N_4666,N_4539);
nand U5361 (N_5361,N_4777,N_4644);
nor U5362 (N_5362,N_4881,N_4836);
or U5363 (N_5363,N_4666,N_4534);
nor U5364 (N_5364,N_4649,N_4686);
nand U5365 (N_5365,N_4796,N_4682);
nor U5366 (N_5366,N_4587,N_4558);
and U5367 (N_5367,N_4872,N_4859);
or U5368 (N_5368,N_4764,N_4763);
or U5369 (N_5369,N_4870,N_4744);
and U5370 (N_5370,N_4636,N_4523);
xor U5371 (N_5371,N_4996,N_4644);
nor U5372 (N_5372,N_4693,N_4792);
and U5373 (N_5373,N_4778,N_4755);
nor U5374 (N_5374,N_4818,N_4705);
nor U5375 (N_5375,N_4951,N_4545);
nor U5376 (N_5376,N_4583,N_4795);
nand U5377 (N_5377,N_4701,N_4614);
and U5378 (N_5378,N_4966,N_4580);
xor U5379 (N_5379,N_4544,N_4502);
nand U5380 (N_5380,N_4582,N_4706);
nand U5381 (N_5381,N_4693,N_4779);
and U5382 (N_5382,N_4505,N_4516);
or U5383 (N_5383,N_4949,N_4670);
or U5384 (N_5384,N_4905,N_4572);
nand U5385 (N_5385,N_4628,N_4576);
or U5386 (N_5386,N_4708,N_4758);
or U5387 (N_5387,N_4839,N_4548);
nor U5388 (N_5388,N_4705,N_4703);
nand U5389 (N_5389,N_4682,N_4717);
nor U5390 (N_5390,N_4890,N_4511);
nor U5391 (N_5391,N_4806,N_4825);
or U5392 (N_5392,N_4596,N_4658);
and U5393 (N_5393,N_4535,N_4677);
nand U5394 (N_5394,N_4690,N_4937);
nand U5395 (N_5395,N_4949,N_4666);
or U5396 (N_5396,N_4880,N_4641);
nand U5397 (N_5397,N_4618,N_4615);
or U5398 (N_5398,N_4519,N_4676);
and U5399 (N_5399,N_4699,N_4518);
nand U5400 (N_5400,N_4811,N_4969);
nor U5401 (N_5401,N_4882,N_4518);
nor U5402 (N_5402,N_4589,N_4896);
nand U5403 (N_5403,N_4602,N_4624);
and U5404 (N_5404,N_4563,N_4772);
nand U5405 (N_5405,N_4943,N_4774);
nand U5406 (N_5406,N_4876,N_4842);
nand U5407 (N_5407,N_4948,N_4765);
nand U5408 (N_5408,N_4934,N_4850);
and U5409 (N_5409,N_4699,N_4608);
or U5410 (N_5410,N_4790,N_4559);
or U5411 (N_5411,N_4551,N_4915);
and U5412 (N_5412,N_4805,N_4608);
or U5413 (N_5413,N_4524,N_4855);
or U5414 (N_5414,N_4569,N_4871);
and U5415 (N_5415,N_4831,N_4783);
or U5416 (N_5416,N_4951,N_4945);
nor U5417 (N_5417,N_4523,N_4746);
nand U5418 (N_5418,N_4509,N_4865);
nor U5419 (N_5419,N_4793,N_4539);
or U5420 (N_5420,N_4779,N_4601);
and U5421 (N_5421,N_4782,N_4546);
and U5422 (N_5422,N_4658,N_4599);
or U5423 (N_5423,N_4894,N_4658);
and U5424 (N_5424,N_4678,N_4606);
nand U5425 (N_5425,N_4672,N_4632);
or U5426 (N_5426,N_4976,N_4591);
nand U5427 (N_5427,N_4958,N_4721);
nor U5428 (N_5428,N_4541,N_4863);
nand U5429 (N_5429,N_4852,N_4907);
or U5430 (N_5430,N_4717,N_4964);
or U5431 (N_5431,N_4900,N_4547);
and U5432 (N_5432,N_4790,N_4871);
nor U5433 (N_5433,N_4548,N_4778);
or U5434 (N_5434,N_4821,N_4653);
nor U5435 (N_5435,N_4836,N_4751);
xor U5436 (N_5436,N_4641,N_4712);
or U5437 (N_5437,N_4684,N_4991);
nand U5438 (N_5438,N_4545,N_4636);
nand U5439 (N_5439,N_4846,N_4545);
nor U5440 (N_5440,N_4556,N_4918);
nor U5441 (N_5441,N_4993,N_4946);
nand U5442 (N_5442,N_4998,N_4752);
nor U5443 (N_5443,N_4759,N_4684);
or U5444 (N_5444,N_4613,N_4831);
nor U5445 (N_5445,N_4998,N_4635);
nor U5446 (N_5446,N_4690,N_4951);
or U5447 (N_5447,N_4557,N_4854);
or U5448 (N_5448,N_4860,N_4854);
or U5449 (N_5449,N_4860,N_4729);
or U5450 (N_5450,N_4772,N_4916);
nor U5451 (N_5451,N_4680,N_4559);
or U5452 (N_5452,N_4597,N_4945);
nor U5453 (N_5453,N_4692,N_4834);
or U5454 (N_5454,N_4724,N_4960);
nand U5455 (N_5455,N_4517,N_4860);
and U5456 (N_5456,N_4609,N_4647);
nand U5457 (N_5457,N_4887,N_4523);
nand U5458 (N_5458,N_4953,N_4544);
and U5459 (N_5459,N_4896,N_4635);
nor U5460 (N_5460,N_4972,N_4903);
nor U5461 (N_5461,N_4902,N_4502);
nor U5462 (N_5462,N_4975,N_4571);
or U5463 (N_5463,N_4979,N_4634);
nand U5464 (N_5464,N_4678,N_4846);
and U5465 (N_5465,N_4718,N_4938);
nand U5466 (N_5466,N_4539,N_4810);
or U5467 (N_5467,N_4866,N_4975);
nand U5468 (N_5468,N_4700,N_4681);
nor U5469 (N_5469,N_4594,N_4640);
or U5470 (N_5470,N_4927,N_4872);
and U5471 (N_5471,N_4813,N_4851);
nor U5472 (N_5472,N_4664,N_4745);
nand U5473 (N_5473,N_4732,N_4538);
xor U5474 (N_5474,N_4510,N_4732);
nor U5475 (N_5475,N_4785,N_4512);
and U5476 (N_5476,N_4516,N_4689);
and U5477 (N_5477,N_4850,N_4988);
nor U5478 (N_5478,N_4798,N_4558);
and U5479 (N_5479,N_4701,N_4599);
nand U5480 (N_5480,N_4771,N_4936);
nor U5481 (N_5481,N_4979,N_4584);
and U5482 (N_5482,N_4726,N_4664);
nand U5483 (N_5483,N_4854,N_4515);
nor U5484 (N_5484,N_4727,N_4774);
nor U5485 (N_5485,N_4856,N_4770);
and U5486 (N_5486,N_4617,N_4772);
xnor U5487 (N_5487,N_4808,N_4840);
and U5488 (N_5488,N_4673,N_4622);
nor U5489 (N_5489,N_4934,N_4922);
or U5490 (N_5490,N_4970,N_4698);
and U5491 (N_5491,N_4944,N_4787);
nor U5492 (N_5492,N_4963,N_4522);
nand U5493 (N_5493,N_4874,N_4849);
nor U5494 (N_5494,N_4877,N_4667);
nor U5495 (N_5495,N_4827,N_4533);
nor U5496 (N_5496,N_4849,N_4841);
and U5497 (N_5497,N_4911,N_4744);
nor U5498 (N_5498,N_4887,N_4518);
and U5499 (N_5499,N_4692,N_4826);
nor U5500 (N_5500,N_5354,N_5239);
nor U5501 (N_5501,N_5424,N_5158);
or U5502 (N_5502,N_5088,N_5056);
nor U5503 (N_5503,N_5033,N_5059);
nand U5504 (N_5504,N_5460,N_5497);
or U5505 (N_5505,N_5325,N_5423);
nand U5506 (N_5506,N_5180,N_5147);
nand U5507 (N_5507,N_5435,N_5352);
and U5508 (N_5508,N_5048,N_5055);
and U5509 (N_5509,N_5288,N_5084);
and U5510 (N_5510,N_5282,N_5037);
xor U5511 (N_5511,N_5372,N_5350);
nand U5512 (N_5512,N_5198,N_5149);
nand U5513 (N_5513,N_5269,N_5258);
and U5514 (N_5514,N_5476,N_5225);
and U5515 (N_5515,N_5047,N_5197);
xor U5516 (N_5516,N_5151,N_5474);
or U5517 (N_5517,N_5000,N_5026);
and U5518 (N_5518,N_5215,N_5315);
and U5519 (N_5519,N_5445,N_5126);
and U5520 (N_5520,N_5112,N_5292);
nor U5521 (N_5521,N_5241,N_5275);
or U5522 (N_5522,N_5238,N_5066);
or U5523 (N_5523,N_5490,N_5220);
or U5524 (N_5524,N_5484,N_5155);
or U5525 (N_5525,N_5378,N_5256);
or U5526 (N_5526,N_5371,N_5345);
and U5527 (N_5527,N_5310,N_5464);
or U5528 (N_5528,N_5223,N_5322);
nand U5529 (N_5529,N_5312,N_5331);
and U5530 (N_5530,N_5163,N_5235);
nand U5531 (N_5531,N_5254,N_5039);
nand U5532 (N_5532,N_5391,N_5458);
nor U5533 (N_5533,N_5382,N_5038);
or U5534 (N_5534,N_5005,N_5092);
nor U5535 (N_5535,N_5478,N_5116);
nand U5536 (N_5536,N_5176,N_5347);
or U5537 (N_5537,N_5487,N_5205);
or U5538 (N_5538,N_5319,N_5025);
nor U5539 (N_5539,N_5366,N_5019);
nor U5540 (N_5540,N_5251,N_5363);
nand U5541 (N_5541,N_5496,N_5316);
nand U5542 (N_5542,N_5291,N_5014);
nand U5543 (N_5543,N_5070,N_5052);
and U5544 (N_5544,N_5448,N_5498);
nor U5545 (N_5545,N_5489,N_5379);
or U5546 (N_5546,N_5074,N_5044);
nor U5547 (N_5547,N_5168,N_5376);
or U5548 (N_5548,N_5323,N_5054);
or U5549 (N_5549,N_5188,N_5051);
nor U5550 (N_5550,N_5397,N_5427);
or U5551 (N_5551,N_5106,N_5479);
or U5552 (N_5552,N_5230,N_5078);
nand U5553 (N_5553,N_5399,N_5380);
nor U5554 (N_5554,N_5173,N_5404);
nand U5555 (N_5555,N_5160,N_5206);
and U5556 (N_5556,N_5193,N_5299);
and U5557 (N_5557,N_5185,N_5260);
nand U5558 (N_5558,N_5253,N_5200);
xor U5559 (N_5559,N_5061,N_5336);
and U5560 (N_5560,N_5456,N_5293);
nor U5561 (N_5561,N_5332,N_5166);
nand U5562 (N_5562,N_5271,N_5388);
and U5563 (N_5563,N_5086,N_5202);
and U5564 (N_5564,N_5094,N_5141);
nand U5565 (N_5565,N_5343,N_5221);
xnor U5566 (N_5566,N_5021,N_5276);
nand U5567 (N_5567,N_5060,N_5156);
or U5568 (N_5568,N_5255,N_5320);
nand U5569 (N_5569,N_5192,N_5344);
nand U5570 (N_5570,N_5194,N_5085);
or U5571 (N_5571,N_5053,N_5091);
and U5572 (N_5572,N_5407,N_5265);
nand U5573 (N_5573,N_5028,N_5381);
or U5574 (N_5574,N_5146,N_5229);
nor U5575 (N_5575,N_5280,N_5471);
or U5576 (N_5576,N_5032,N_5421);
and U5577 (N_5577,N_5453,N_5483);
or U5578 (N_5578,N_5353,N_5102);
nor U5579 (N_5579,N_5015,N_5017);
or U5580 (N_5580,N_5425,N_5357);
nor U5581 (N_5581,N_5400,N_5369);
or U5582 (N_5582,N_5289,N_5023);
or U5583 (N_5583,N_5481,N_5182);
nand U5584 (N_5584,N_5330,N_5297);
and U5585 (N_5585,N_5327,N_5281);
or U5586 (N_5586,N_5217,N_5428);
nand U5587 (N_5587,N_5351,N_5326);
xor U5588 (N_5588,N_5472,N_5268);
or U5589 (N_5589,N_5262,N_5298);
and U5590 (N_5590,N_5101,N_5461);
nor U5591 (N_5591,N_5204,N_5311);
and U5592 (N_5592,N_5348,N_5465);
or U5593 (N_5593,N_5042,N_5377);
nor U5594 (N_5594,N_5236,N_5375);
nand U5595 (N_5595,N_5247,N_5485);
or U5596 (N_5596,N_5090,N_5355);
and U5597 (N_5597,N_5099,N_5093);
nor U5598 (N_5598,N_5389,N_5294);
or U5599 (N_5599,N_5416,N_5267);
or U5600 (N_5600,N_5250,N_5113);
or U5601 (N_5601,N_5179,N_5475);
xnor U5602 (N_5602,N_5131,N_5008);
and U5603 (N_5603,N_5287,N_5171);
and U5604 (N_5604,N_5029,N_5145);
xnor U5605 (N_5605,N_5307,N_5115);
nor U5606 (N_5606,N_5277,N_5300);
and U5607 (N_5607,N_5279,N_5270);
or U5608 (N_5608,N_5161,N_5449);
nand U5609 (N_5609,N_5433,N_5429);
and U5610 (N_5610,N_5309,N_5257);
nand U5611 (N_5611,N_5076,N_5308);
and U5612 (N_5612,N_5001,N_5152);
and U5613 (N_5613,N_5367,N_5272);
or U5614 (N_5614,N_5227,N_5124);
xor U5615 (N_5615,N_5286,N_5383);
nor U5616 (N_5616,N_5360,N_5334);
nor U5617 (N_5617,N_5142,N_5219);
nor U5618 (N_5618,N_5395,N_5196);
or U5619 (N_5619,N_5234,N_5210);
nand U5620 (N_5620,N_5341,N_5089);
and U5621 (N_5621,N_5246,N_5153);
xor U5622 (N_5622,N_5263,N_5136);
or U5623 (N_5623,N_5412,N_5036);
or U5624 (N_5624,N_5467,N_5067);
or U5625 (N_5625,N_5027,N_5138);
and U5626 (N_5626,N_5415,N_5164);
or U5627 (N_5627,N_5438,N_5237);
and U5628 (N_5628,N_5466,N_5339);
nor U5629 (N_5629,N_5216,N_5314);
and U5630 (N_5630,N_5333,N_5318);
or U5631 (N_5631,N_5165,N_5420);
nor U5632 (N_5632,N_5049,N_5495);
nand U5633 (N_5633,N_5181,N_5401);
and U5634 (N_5634,N_5422,N_5480);
and U5635 (N_5635,N_5385,N_5259);
and U5636 (N_5636,N_5317,N_5045);
and U5637 (N_5637,N_5071,N_5139);
or U5638 (N_5638,N_5414,N_5432);
or U5639 (N_5639,N_5003,N_5177);
or U5640 (N_5640,N_5328,N_5486);
or U5641 (N_5641,N_5043,N_5356);
or U5642 (N_5642,N_5373,N_5174);
nor U5643 (N_5643,N_5172,N_5444);
or U5644 (N_5644,N_5468,N_5107);
nor U5645 (N_5645,N_5082,N_5451);
nand U5646 (N_5646,N_5103,N_5121);
and U5647 (N_5647,N_5413,N_5063);
or U5648 (N_5648,N_5175,N_5096);
or U5649 (N_5649,N_5162,N_5114);
and U5650 (N_5650,N_5390,N_5306);
nor U5651 (N_5651,N_5417,N_5492);
nor U5652 (N_5652,N_5018,N_5214);
or U5653 (N_5653,N_5240,N_5081);
and U5654 (N_5654,N_5128,N_5050);
and U5655 (N_5655,N_5183,N_5118);
nand U5656 (N_5656,N_5305,N_5170);
and U5657 (N_5657,N_5340,N_5443);
and U5658 (N_5658,N_5452,N_5100);
and U5659 (N_5659,N_5266,N_5104);
or U5660 (N_5660,N_5338,N_5013);
and U5661 (N_5661,N_5295,N_5184);
nand U5662 (N_5662,N_5321,N_5022);
nor U5663 (N_5663,N_5494,N_5064);
or U5664 (N_5664,N_5150,N_5057);
nand U5665 (N_5665,N_5396,N_5189);
nand U5666 (N_5666,N_5386,N_5313);
nor U5667 (N_5667,N_5191,N_5134);
or U5668 (N_5668,N_5491,N_5303);
or U5669 (N_5669,N_5359,N_5418);
nor U5670 (N_5670,N_5007,N_5224);
nand U5671 (N_5671,N_5358,N_5010);
or U5672 (N_5672,N_5199,N_5095);
nand U5673 (N_5673,N_5482,N_5446);
and U5674 (N_5674,N_5470,N_5137);
or U5675 (N_5675,N_5208,N_5387);
nor U5676 (N_5676,N_5245,N_5108);
nand U5677 (N_5677,N_5079,N_5035);
or U5678 (N_5678,N_5083,N_5329);
nand U5679 (N_5679,N_5127,N_5009);
xor U5680 (N_5680,N_5222,N_5169);
nor U5681 (N_5681,N_5419,N_5434);
and U5682 (N_5682,N_5098,N_5040);
and U5683 (N_5683,N_5290,N_5402);
nor U5684 (N_5684,N_5403,N_5368);
and U5685 (N_5685,N_5087,N_5190);
or U5686 (N_5686,N_5301,N_5337);
or U5687 (N_5687,N_5228,N_5248);
or U5688 (N_5688,N_5159,N_5075);
nand U5689 (N_5689,N_5477,N_5342);
or U5690 (N_5690,N_5186,N_5213);
nand U5691 (N_5691,N_5457,N_5374);
and U5692 (N_5692,N_5426,N_5109);
or U5693 (N_5693,N_5077,N_5157);
nor U5694 (N_5694,N_5006,N_5211);
or U5695 (N_5695,N_5441,N_5195);
and U5696 (N_5696,N_5144,N_5439);
nand U5697 (N_5697,N_5117,N_5178);
nor U5698 (N_5698,N_5030,N_5459);
nand U5699 (N_5699,N_5450,N_5285);
nor U5700 (N_5700,N_5011,N_5447);
nor U5701 (N_5701,N_5231,N_5002);
nor U5702 (N_5702,N_5135,N_5349);
nand U5703 (N_5703,N_5125,N_5454);
or U5704 (N_5704,N_5207,N_5004);
nand U5705 (N_5705,N_5278,N_5473);
nand U5706 (N_5706,N_5394,N_5252);
nand U5707 (N_5707,N_5273,N_5097);
or U5708 (N_5708,N_5405,N_5411);
nor U5709 (N_5709,N_5020,N_5324);
or U5710 (N_5710,N_5140,N_5201);
or U5711 (N_5711,N_5110,N_5072);
xnor U5712 (N_5712,N_5046,N_5080);
and U5713 (N_5713,N_5283,N_5410);
or U5714 (N_5714,N_5493,N_5132);
or U5715 (N_5715,N_5062,N_5365);
or U5716 (N_5716,N_5346,N_5302);
nand U5717 (N_5717,N_5362,N_5073);
nand U5718 (N_5718,N_5212,N_5148);
nor U5719 (N_5719,N_5261,N_5249);
or U5720 (N_5720,N_5154,N_5384);
xnor U5721 (N_5721,N_5119,N_5068);
and U5722 (N_5722,N_5304,N_5065);
nor U5723 (N_5723,N_5024,N_5130);
nor U5724 (N_5724,N_5209,N_5440);
or U5725 (N_5725,N_5244,N_5203);
or U5726 (N_5726,N_5123,N_5437);
and U5727 (N_5727,N_5406,N_5284);
or U5728 (N_5728,N_5233,N_5133);
nand U5729 (N_5729,N_5105,N_5436);
and U5730 (N_5730,N_5409,N_5226);
and U5731 (N_5731,N_5408,N_5499);
nor U5732 (N_5732,N_5120,N_5187);
and U5733 (N_5733,N_5431,N_5031);
or U5734 (N_5734,N_5167,N_5218);
and U5735 (N_5735,N_5012,N_5463);
or U5736 (N_5736,N_5430,N_5069);
or U5737 (N_5737,N_5243,N_5111);
and U5738 (N_5738,N_5016,N_5143);
or U5739 (N_5739,N_5122,N_5469);
nand U5740 (N_5740,N_5041,N_5364);
or U5741 (N_5741,N_5370,N_5335);
and U5742 (N_5742,N_5455,N_5393);
or U5743 (N_5743,N_5242,N_5034);
or U5744 (N_5744,N_5232,N_5361);
nand U5745 (N_5745,N_5129,N_5274);
and U5746 (N_5746,N_5058,N_5398);
nand U5747 (N_5747,N_5392,N_5488);
nor U5748 (N_5748,N_5442,N_5462);
nand U5749 (N_5749,N_5296,N_5264);
or U5750 (N_5750,N_5499,N_5369);
nand U5751 (N_5751,N_5172,N_5343);
or U5752 (N_5752,N_5242,N_5138);
nand U5753 (N_5753,N_5418,N_5402);
nor U5754 (N_5754,N_5160,N_5371);
nand U5755 (N_5755,N_5395,N_5326);
or U5756 (N_5756,N_5057,N_5083);
nor U5757 (N_5757,N_5422,N_5216);
nor U5758 (N_5758,N_5311,N_5289);
nand U5759 (N_5759,N_5125,N_5452);
or U5760 (N_5760,N_5095,N_5479);
nor U5761 (N_5761,N_5196,N_5160);
and U5762 (N_5762,N_5209,N_5144);
nand U5763 (N_5763,N_5428,N_5019);
nand U5764 (N_5764,N_5499,N_5221);
or U5765 (N_5765,N_5297,N_5431);
or U5766 (N_5766,N_5199,N_5082);
or U5767 (N_5767,N_5049,N_5066);
and U5768 (N_5768,N_5095,N_5189);
nand U5769 (N_5769,N_5140,N_5438);
or U5770 (N_5770,N_5446,N_5440);
or U5771 (N_5771,N_5352,N_5280);
or U5772 (N_5772,N_5198,N_5478);
and U5773 (N_5773,N_5369,N_5149);
or U5774 (N_5774,N_5305,N_5472);
nor U5775 (N_5775,N_5209,N_5488);
nand U5776 (N_5776,N_5180,N_5456);
nand U5777 (N_5777,N_5334,N_5213);
or U5778 (N_5778,N_5047,N_5393);
and U5779 (N_5779,N_5307,N_5205);
nor U5780 (N_5780,N_5007,N_5214);
or U5781 (N_5781,N_5359,N_5170);
nand U5782 (N_5782,N_5164,N_5169);
and U5783 (N_5783,N_5121,N_5228);
and U5784 (N_5784,N_5240,N_5469);
or U5785 (N_5785,N_5446,N_5068);
and U5786 (N_5786,N_5408,N_5281);
nor U5787 (N_5787,N_5390,N_5314);
and U5788 (N_5788,N_5139,N_5264);
and U5789 (N_5789,N_5225,N_5386);
nand U5790 (N_5790,N_5070,N_5464);
nand U5791 (N_5791,N_5319,N_5415);
nand U5792 (N_5792,N_5014,N_5183);
nand U5793 (N_5793,N_5034,N_5182);
or U5794 (N_5794,N_5129,N_5267);
or U5795 (N_5795,N_5132,N_5070);
nor U5796 (N_5796,N_5293,N_5358);
nor U5797 (N_5797,N_5099,N_5062);
and U5798 (N_5798,N_5174,N_5319);
or U5799 (N_5799,N_5263,N_5201);
or U5800 (N_5800,N_5072,N_5157);
and U5801 (N_5801,N_5346,N_5001);
nand U5802 (N_5802,N_5224,N_5098);
or U5803 (N_5803,N_5006,N_5096);
or U5804 (N_5804,N_5366,N_5173);
nand U5805 (N_5805,N_5198,N_5263);
xor U5806 (N_5806,N_5465,N_5195);
or U5807 (N_5807,N_5383,N_5146);
nor U5808 (N_5808,N_5243,N_5369);
and U5809 (N_5809,N_5377,N_5359);
and U5810 (N_5810,N_5221,N_5433);
nor U5811 (N_5811,N_5083,N_5493);
or U5812 (N_5812,N_5136,N_5490);
xor U5813 (N_5813,N_5305,N_5405);
nor U5814 (N_5814,N_5138,N_5375);
nor U5815 (N_5815,N_5196,N_5249);
and U5816 (N_5816,N_5491,N_5200);
and U5817 (N_5817,N_5097,N_5066);
nor U5818 (N_5818,N_5149,N_5033);
and U5819 (N_5819,N_5341,N_5469);
nand U5820 (N_5820,N_5148,N_5471);
and U5821 (N_5821,N_5151,N_5137);
nand U5822 (N_5822,N_5490,N_5357);
nor U5823 (N_5823,N_5082,N_5231);
nor U5824 (N_5824,N_5082,N_5213);
nor U5825 (N_5825,N_5292,N_5153);
or U5826 (N_5826,N_5268,N_5048);
nor U5827 (N_5827,N_5151,N_5357);
and U5828 (N_5828,N_5212,N_5008);
nand U5829 (N_5829,N_5098,N_5309);
or U5830 (N_5830,N_5158,N_5005);
nor U5831 (N_5831,N_5488,N_5217);
and U5832 (N_5832,N_5065,N_5318);
nand U5833 (N_5833,N_5349,N_5266);
and U5834 (N_5834,N_5061,N_5077);
nand U5835 (N_5835,N_5496,N_5310);
and U5836 (N_5836,N_5290,N_5020);
or U5837 (N_5837,N_5315,N_5014);
or U5838 (N_5838,N_5285,N_5113);
nor U5839 (N_5839,N_5244,N_5096);
nand U5840 (N_5840,N_5081,N_5324);
nand U5841 (N_5841,N_5148,N_5165);
xor U5842 (N_5842,N_5459,N_5271);
nor U5843 (N_5843,N_5439,N_5124);
nor U5844 (N_5844,N_5428,N_5110);
nor U5845 (N_5845,N_5027,N_5403);
or U5846 (N_5846,N_5193,N_5378);
xor U5847 (N_5847,N_5384,N_5179);
nor U5848 (N_5848,N_5240,N_5444);
or U5849 (N_5849,N_5078,N_5012);
or U5850 (N_5850,N_5381,N_5457);
and U5851 (N_5851,N_5367,N_5305);
nor U5852 (N_5852,N_5158,N_5001);
xnor U5853 (N_5853,N_5308,N_5253);
nor U5854 (N_5854,N_5035,N_5255);
or U5855 (N_5855,N_5024,N_5036);
and U5856 (N_5856,N_5472,N_5382);
or U5857 (N_5857,N_5378,N_5178);
nor U5858 (N_5858,N_5065,N_5017);
nand U5859 (N_5859,N_5222,N_5418);
or U5860 (N_5860,N_5465,N_5334);
nor U5861 (N_5861,N_5429,N_5063);
nand U5862 (N_5862,N_5423,N_5061);
nor U5863 (N_5863,N_5293,N_5183);
nor U5864 (N_5864,N_5127,N_5046);
nor U5865 (N_5865,N_5368,N_5150);
nand U5866 (N_5866,N_5400,N_5123);
nand U5867 (N_5867,N_5251,N_5100);
and U5868 (N_5868,N_5115,N_5458);
and U5869 (N_5869,N_5300,N_5218);
or U5870 (N_5870,N_5107,N_5285);
and U5871 (N_5871,N_5393,N_5138);
nor U5872 (N_5872,N_5258,N_5190);
nand U5873 (N_5873,N_5113,N_5251);
nor U5874 (N_5874,N_5020,N_5071);
nand U5875 (N_5875,N_5451,N_5437);
nand U5876 (N_5876,N_5385,N_5411);
xnor U5877 (N_5877,N_5144,N_5270);
or U5878 (N_5878,N_5355,N_5446);
nand U5879 (N_5879,N_5354,N_5257);
nor U5880 (N_5880,N_5296,N_5407);
nor U5881 (N_5881,N_5495,N_5329);
nor U5882 (N_5882,N_5396,N_5025);
and U5883 (N_5883,N_5448,N_5386);
nand U5884 (N_5884,N_5421,N_5180);
nand U5885 (N_5885,N_5100,N_5029);
nand U5886 (N_5886,N_5357,N_5294);
or U5887 (N_5887,N_5165,N_5292);
and U5888 (N_5888,N_5423,N_5332);
nor U5889 (N_5889,N_5394,N_5092);
or U5890 (N_5890,N_5067,N_5383);
or U5891 (N_5891,N_5107,N_5431);
and U5892 (N_5892,N_5330,N_5340);
and U5893 (N_5893,N_5127,N_5028);
nor U5894 (N_5894,N_5471,N_5215);
or U5895 (N_5895,N_5164,N_5094);
nor U5896 (N_5896,N_5007,N_5399);
nand U5897 (N_5897,N_5383,N_5120);
nor U5898 (N_5898,N_5060,N_5220);
or U5899 (N_5899,N_5179,N_5019);
nor U5900 (N_5900,N_5243,N_5236);
or U5901 (N_5901,N_5403,N_5351);
nand U5902 (N_5902,N_5370,N_5299);
nor U5903 (N_5903,N_5285,N_5263);
nand U5904 (N_5904,N_5052,N_5492);
or U5905 (N_5905,N_5452,N_5401);
nand U5906 (N_5906,N_5420,N_5330);
nor U5907 (N_5907,N_5012,N_5046);
and U5908 (N_5908,N_5052,N_5140);
or U5909 (N_5909,N_5318,N_5292);
and U5910 (N_5910,N_5485,N_5438);
or U5911 (N_5911,N_5256,N_5133);
nor U5912 (N_5912,N_5481,N_5012);
and U5913 (N_5913,N_5435,N_5240);
and U5914 (N_5914,N_5102,N_5219);
and U5915 (N_5915,N_5112,N_5312);
and U5916 (N_5916,N_5397,N_5244);
xnor U5917 (N_5917,N_5352,N_5205);
nor U5918 (N_5918,N_5411,N_5320);
nand U5919 (N_5919,N_5200,N_5314);
and U5920 (N_5920,N_5420,N_5217);
nand U5921 (N_5921,N_5346,N_5107);
or U5922 (N_5922,N_5100,N_5101);
nand U5923 (N_5923,N_5023,N_5072);
or U5924 (N_5924,N_5480,N_5042);
or U5925 (N_5925,N_5015,N_5411);
or U5926 (N_5926,N_5102,N_5445);
and U5927 (N_5927,N_5377,N_5062);
nand U5928 (N_5928,N_5336,N_5005);
nand U5929 (N_5929,N_5342,N_5190);
nand U5930 (N_5930,N_5499,N_5224);
or U5931 (N_5931,N_5288,N_5359);
nand U5932 (N_5932,N_5339,N_5478);
nand U5933 (N_5933,N_5361,N_5074);
or U5934 (N_5934,N_5061,N_5429);
nand U5935 (N_5935,N_5442,N_5356);
and U5936 (N_5936,N_5075,N_5324);
or U5937 (N_5937,N_5479,N_5126);
and U5938 (N_5938,N_5030,N_5290);
and U5939 (N_5939,N_5337,N_5066);
nand U5940 (N_5940,N_5375,N_5177);
nor U5941 (N_5941,N_5209,N_5328);
nand U5942 (N_5942,N_5382,N_5336);
nand U5943 (N_5943,N_5007,N_5229);
or U5944 (N_5944,N_5381,N_5341);
nor U5945 (N_5945,N_5299,N_5316);
nor U5946 (N_5946,N_5027,N_5421);
nor U5947 (N_5947,N_5370,N_5053);
nand U5948 (N_5948,N_5404,N_5022);
nor U5949 (N_5949,N_5272,N_5151);
and U5950 (N_5950,N_5203,N_5479);
or U5951 (N_5951,N_5303,N_5093);
and U5952 (N_5952,N_5497,N_5139);
or U5953 (N_5953,N_5103,N_5479);
or U5954 (N_5954,N_5258,N_5330);
nand U5955 (N_5955,N_5143,N_5216);
and U5956 (N_5956,N_5358,N_5257);
or U5957 (N_5957,N_5039,N_5312);
nor U5958 (N_5958,N_5268,N_5062);
or U5959 (N_5959,N_5009,N_5212);
nor U5960 (N_5960,N_5051,N_5469);
or U5961 (N_5961,N_5113,N_5052);
nand U5962 (N_5962,N_5295,N_5227);
nor U5963 (N_5963,N_5330,N_5426);
and U5964 (N_5964,N_5055,N_5171);
and U5965 (N_5965,N_5178,N_5043);
xnor U5966 (N_5966,N_5370,N_5282);
nor U5967 (N_5967,N_5365,N_5057);
and U5968 (N_5968,N_5005,N_5380);
or U5969 (N_5969,N_5133,N_5096);
xnor U5970 (N_5970,N_5231,N_5293);
nor U5971 (N_5971,N_5061,N_5130);
or U5972 (N_5972,N_5431,N_5162);
and U5973 (N_5973,N_5209,N_5354);
nand U5974 (N_5974,N_5032,N_5013);
xnor U5975 (N_5975,N_5136,N_5401);
and U5976 (N_5976,N_5321,N_5192);
nor U5977 (N_5977,N_5480,N_5138);
nor U5978 (N_5978,N_5447,N_5363);
nand U5979 (N_5979,N_5110,N_5389);
and U5980 (N_5980,N_5353,N_5235);
or U5981 (N_5981,N_5089,N_5334);
xnor U5982 (N_5982,N_5132,N_5246);
nand U5983 (N_5983,N_5214,N_5431);
or U5984 (N_5984,N_5484,N_5423);
or U5985 (N_5985,N_5008,N_5358);
nor U5986 (N_5986,N_5315,N_5435);
and U5987 (N_5987,N_5049,N_5297);
nand U5988 (N_5988,N_5347,N_5198);
nand U5989 (N_5989,N_5060,N_5490);
or U5990 (N_5990,N_5296,N_5203);
or U5991 (N_5991,N_5001,N_5488);
nand U5992 (N_5992,N_5097,N_5490);
or U5993 (N_5993,N_5229,N_5189);
nor U5994 (N_5994,N_5093,N_5254);
nor U5995 (N_5995,N_5016,N_5306);
and U5996 (N_5996,N_5241,N_5002);
nor U5997 (N_5997,N_5332,N_5346);
or U5998 (N_5998,N_5403,N_5422);
and U5999 (N_5999,N_5172,N_5213);
nor U6000 (N_6000,N_5932,N_5824);
nor U6001 (N_6001,N_5672,N_5797);
and U6002 (N_6002,N_5790,N_5584);
or U6003 (N_6003,N_5724,N_5854);
and U6004 (N_6004,N_5810,N_5506);
and U6005 (N_6005,N_5916,N_5757);
nor U6006 (N_6006,N_5684,N_5785);
or U6007 (N_6007,N_5691,N_5967);
or U6008 (N_6008,N_5938,N_5598);
and U6009 (N_6009,N_5934,N_5696);
or U6010 (N_6010,N_5791,N_5693);
nor U6011 (N_6011,N_5728,N_5620);
and U6012 (N_6012,N_5835,N_5540);
and U6013 (N_6013,N_5544,N_5906);
and U6014 (N_6014,N_5589,N_5813);
nand U6015 (N_6015,N_5914,N_5726);
and U6016 (N_6016,N_5919,N_5971);
and U6017 (N_6017,N_5963,N_5775);
and U6018 (N_6018,N_5863,N_5812);
nor U6019 (N_6019,N_5591,N_5892);
and U6020 (N_6020,N_5804,N_5543);
nand U6021 (N_6021,N_5516,N_5970);
nor U6022 (N_6022,N_5652,N_5510);
or U6023 (N_6023,N_5703,N_5943);
and U6024 (N_6024,N_5753,N_5607);
or U6025 (N_6025,N_5799,N_5641);
nor U6026 (N_6026,N_5993,N_5923);
nand U6027 (N_6027,N_5920,N_5975);
nor U6028 (N_6028,N_5711,N_5925);
nand U6029 (N_6029,N_5674,N_5682);
and U6030 (N_6030,N_5735,N_5864);
nand U6031 (N_6031,N_5670,N_5909);
or U6032 (N_6032,N_5865,N_5978);
xor U6033 (N_6033,N_5782,N_5819);
or U6034 (N_6034,N_5855,N_5657);
or U6035 (N_6035,N_5985,N_5936);
nor U6036 (N_6036,N_5847,N_5958);
nand U6037 (N_6037,N_5562,N_5722);
and U6038 (N_6038,N_5907,N_5692);
nand U6039 (N_6039,N_5681,N_5505);
nand U6040 (N_6040,N_5755,N_5667);
or U6041 (N_6041,N_5573,N_5877);
nor U6042 (N_6042,N_5525,N_5754);
or U6043 (N_6043,N_5802,N_5942);
or U6044 (N_6044,N_5974,N_5781);
xor U6045 (N_6045,N_5629,N_5746);
nand U6046 (N_6046,N_5986,N_5960);
xnor U6047 (N_6047,N_5683,N_5660);
and U6048 (N_6048,N_5921,N_5990);
or U6049 (N_6049,N_5537,N_5730);
nor U6050 (N_6050,N_5617,N_5772);
and U6051 (N_6051,N_5881,N_5519);
and U6052 (N_6052,N_5602,N_5874);
or U6053 (N_6053,N_5704,N_5846);
and U6054 (N_6054,N_5729,N_5902);
nor U6055 (N_6055,N_5756,N_5608);
or U6056 (N_6056,N_5664,N_5953);
xnor U6057 (N_6057,N_5642,N_5597);
or U6058 (N_6058,N_5995,N_5701);
and U6059 (N_6059,N_5595,N_5590);
and U6060 (N_6060,N_5644,N_5679);
nor U6061 (N_6061,N_5687,N_5520);
or U6062 (N_6062,N_5827,N_5758);
nand U6063 (N_6063,N_5945,N_5928);
nor U6064 (N_6064,N_5935,N_5710);
nor U6065 (N_6065,N_5913,N_5760);
or U6066 (N_6066,N_5850,N_5588);
nand U6067 (N_6067,N_5927,N_5955);
nand U6068 (N_6068,N_5898,N_5513);
nand U6069 (N_6069,N_5581,N_5952);
nand U6070 (N_6070,N_5699,N_5522);
nor U6071 (N_6071,N_5896,N_5976);
nand U6072 (N_6072,N_5825,N_5833);
nand U6073 (N_6073,N_5633,N_5600);
nand U6074 (N_6074,N_5700,N_5763);
nand U6075 (N_6075,N_5599,N_5817);
or U6076 (N_6076,N_5852,N_5697);
nor U6077 (N_6077,N_5648,N_5669);
nor U6078 (N_6078,N_5694,N_5605);
xor U6079 (N_6079,N_5840,N_5721);
nand U6080 (N_6080,N_5830,N_5832);
nor U6081 (N_6081,N_5899,N_5732);
nor U6082 (N_6082,N_5715,N_5764);
or U6083 (N_6083,N_5859,N_5621);
nand U6084 (N_6084,N_5552,N_5631);
nand U6085 (N_6085,N_5717,N_5716);
nor U6086 (N_6086,N_5841,N_5618);
nand U6087 (N_6087,N_5926,N_5713);
or U6088 (N_6088,N_5640,N_5845);
and U6089 (N_6089,N_5838,N_5839);
nand U6090 (N_6090,N_5622,N_5645);
nand U6091 (N_6091,N_5806,N_5737);
and U6092 (N_6092,N_5706,N_5509);
or U6093 (N_6093,N_5912,N_5593);
xnor U6094 (N_6094,N_5871,N_5964);
and U6095 (N_6095,N_5794,N_5529);
nand U6096 (N_6096,N_5594,N_5596);
and U6097 (N_6097,N_5649,N_5861);
or U6098 (N_6098,N_5826,N_5885);
nand U6099 (N_6099,N_5636,N_5507);
nor U6100 (N_6100,N_5527,N_5626);
nand U6101 (N_6101,N_5808,N_5747);
and U6102 (N_6102,N_5820,N_5702);
nand U6103 (N_6103,N_5731,N_5951);
nor U6104 (N_6104,N_5712,N_5613);
or U6105 (N_6105,N_5911,N_5879);
nor U6106 (N_6106,N_5766,N_5709);
and U6107 (N_6107,N_5744,N_5695);
nor U6108 (N_6108,N_5867,N_5603);
and U6109 (N_6109,N_5515,N_5957);
or U6110 (N_6110,N_5815,N_5654);
or U6111 (N_6111,N_5889,N_5745);
nand U6112 (N_6112,N_5587,N_5676);
nand U6113 (N_6113,N_5834,N_5612);
and U6114 (N_6114,N_5627,N_5569);
or U6115 (N_6115,N_5727,N_5580);
and U6116 (N_6116,N_5937,N_5559);
and U6117 (N_6117,N_5615,N_5872);
and U6118 (N_6118,N_5637,N_5518);
or U6119 (N_6119,N_5623,N_5528);
nand U6120 (N_6120,N_5910,N_5961);
or U6121 (N_6121,N_5857,N_5823);
or U6122 (N_6122,N_5579,N_5944);
and U6123 (N_6123,N_5886,N_5814);
nand U6124 (N_6124,N_5673,N_5770);
and U6125 (N_6125,N_5940,N_5947);
nor U6126 (N_6126,N_5742,N_5554);
and U6127 (N_6127,N_5816,N_5980);
or U6128 (N_6128,N_5571,N_5577);
and U6129 (N_6129,N_5965,N_5739);
and U6130 (N_6130,N_5897,N_5551);
and U6131 (N_6131,N_5643,N_5979);
nor U6132 (N_6132,N_5738,N_5860);
and U6133 (N_6133,N_5866,N_5807);
and U6134 (N_6134,N_5984,N_5604);
or U6135 (N_6135,N_5851,N_5788);
nand U6136 (N_6136,N_5610,N_5663);
nand U6137 (N_6137,N_5946,N_5888);
nand U6138 (N_6138,N_5586,N_5939);
nand U6139 (N_6139,N_5930,N_5992);
or U6140 (N_6140,N_5982,N_5658);
nand U6141 (N_6141,N_5989,N_5988);
or U6142 (N_6142,N_5968,N_5558);
nor U6143 (N_6143,N_5675,N_5550);
and U6144 (N_6144,N_5853,N_5685);
and U6145 (N_6145,N_5752,N_5625);
and U6146 (N_6146,N_5624,N_5875);
nor U6147 (N_6147,N_5572,N_5883);
or U6148 (N_6148,N_5796,N_5929);
or U6149 (N_6149,N_5891,N_5690);
and U6150 (N_6150,N_5628,N_5546);
or U6151 (N_6151,N_5856,N_5904);
nor U6152 (N_6152,N_5708,N_5678);
or U6153 (N_6153,N_5659,N_5526);
nand U6154 (N_6154,N_5779,N_5609);
or U6155 (N_6155,N_5821,N_5977);
or U6156 (N_6156,N_5530,N_5714);
nor U6157 (N_6157,N_5668,N_5688);
and U6158 (N_6158,N_5959,N_5619);
nor U6159 (N_6159,N_5759,N_5566);
or U6160 (N_6160,N_5948,N_5614);
or U6161 (N_6161,N_5553,N_5800);
and U6162 (N_6162,N_5858,N_5773);
nand U6163 (N_6163,N_5547,N_5719);
nand U6164 (N_6164,N_5565,N_5725);
and U6165 (N_6165,N_5698,N_5998);
or U6166 (N_6166,N_5511,N_5606);
and U6167 (N_6167,N_5822,N_5793);
nor U6168 (N_6168,N_5662,N_5592);
or U6169 (N_6169,N_5514,N_5705);
xnor U6170 (N_6170,N_5876,N_5776);
and U6171 (N_6171,N_5805,N_5941);
nand U6172 (N_6172,N_5931,N_5575);
or U6173 (N_6173,N_5720,N_5778);
nand U6174 (N_6174,N_5508,N_5862);
or U6175 (N_6175,N_5568,N_5532);
or U6176 (N_6176,N_5539,N_5647);
nor U6177 (N_6177,N_5521,N_5836);
and U6178 (N_6178,N_5769,N_5809);
or U6179 (N_6179,N_5656,N_5534);
or U6180 (N_6180,N_5570,N_5981);
nor U6181 (N_6181,N_5893,N_5924);
nand U6182 (N_6182,N_5922,N_5890);
nand U6183 (N_6183,N_5585,N_5878);
or U6184 (N_6184,N_5500,N_5634);
and U6185 (N_6185,N_5873,N_5818);
and U6186 (N_6186,N_5903,N_5677);
and U6187 (N_6187,N_5887,N_5650);
and U6188 (N_6188,N_5956,N_5842);
and U6189 (N_6189,N_5743,N_5646);
nor U6190 (N_6190,N_5749,N_5771);
nor U6191 (N_6191,N_5523,N_5868);
nand U6192 (N_6192,N_5582,N_5999);
or U6193 (N_6193,N_5991,N_5973);
or U6194 (N_6194,N_5996,N_5601);
and U6195 (N_6195,N_5762,N_5661);
nand U6196 (N_6196,N_5750,N_5578);
nand U6197 (N_6197,N_5616,N_5829);
nand U6198 (N_6198,N_5535,N_5734);
nor U6199 (N_6199,N_5895,N_5723);
nand U6200 (N_6200,N_5784,N_5789);
nor U6201 (N_6201,N_5635,N_5557);
and U6202 (N_6202,N_5741,N_5632);
or U6203 (N_6203,N_5767,N_5574);
or U6204 (N_6204,N_5843,N_5686);
and U6205 (N_6205,N_5560,N_5983);
nor U6206 (N_6206,N_5901,N_5718);
nand U6207 (N_6207,N_5564,N_5639);
xor U6208 (N_6208,N_5531,N_5777);
and U6209 (N_6209,N_5541,N_5900);
xor U6210 (N_6210,N_5576,N_5915);
and U6211 (N_6211,N_5761,N_5880);
xnor U6212 (N_6212,N_5556,N_5549);
or U6213 (N_6213,N_5567,N_5538);
nand U6214 (N_6214,N_5583,N_5548);
and U6215 (N_6215,N_5917,N_5536);
or U6216 (N_6216,N_5630,N_5504);
nor U6217 (N_6217,N_5918,N_5655);
nor U6218 (N_6218,N_5828,N_5811);
or U6219 (N_6219,N_5803,N_5680);
nand U6220 (N_6220,N_5954,N_5666);
and U6221 (N_6221,N_5795,N_5894);
and U6222 (N_6222,N_5949,N_5503);
and U6223 (N_6223,N_5882,N_5780);
or U6224 (N_6224,N_5848,N_5768);
and U6225 (N_6225,N_5517,N_5792);
nand U6226 (N_6226,N_5653,N_5997);
or U6227 (N_6227,N_5765,N_5783);
or U6228 (N_6228,N_5933,N_5966);
nor U6229 (N_6229,N_5707,N_5740);
nand U6230 (N_6230,N_5733,N_5972);
and U6231 (N_6231,N_5512,N_5524);
nand U6232 (N_6232,N_5563,N_5651);
nor U6233 (N_6233,N_5849,N_5844);
or U6234 (N_6234,N_5638,N_5748);
or U6235 (N_6235,N_5908,N_5665);
nand U6236 (N_6236,N_5798,N_5545);
or U6237 (N_6237,N_5869,N_5671);
nand U6238 (N_6238,N_5502,N_5736);
or U6239 (N_6239,N_5884,N_5870);
xnor U6240 (N_6240,N_5969,N_5611);
or U6241 (N_6241,N_5801,N_5555);
nor U6242 (N_6242,N_5994,N_5786);
nor U6243 (N_6243,N_5561,N_5787);
nand U6244 (N_6244,N_5751,N_5905);
nor U6245 (N_6245,N_5962,N_5987);
nor U6246 (N_6246,N_5831,N_5501);
or U6247 (N_6247,N_5533,N_5542);
or U6248 (N_6248,N_5837,N_5950);
nand U6249 (N_6249,N_5689,N_5774);
and U6250 (N_6250,N_5671,N_5682);
or U6251 (N_6251,N_5692,N_5989);
or U6252 (N_6252,N_5683,N_5591);
and U6253 (N_6253,N_5518,N_5511);
and U6254 (N_6254,N_5961,N_5578);
nand U6255 (N_6255,N_5675,N_5897);
nor U6256 (N_6256,N_5572,N_5579);
or U6257 (N_6257,N_5513,N_5532);
or U6258 (N_6258,N_5626,N_5872);
nand U6259 (N_6259,N_5574,N_5550);
or U6260 (N_6260,N_5778,N_5698);
nor U6261 (N_6261,N_5731,N_5546);
and U6262 (N_6262,N_5969,N_5678);
or U6263 (N_6263,N_5952,N_5668);
nand U6264 (N_6264,N_5607,N_5556);
or U6265 (N_6265,N_5893,N_5539);
nand U6266 (N_6266,N_5935,N_5717);
nor U6267 (N_6267,N_5898,N_5679);
and U6268 (N_6268,N_5812,N_5626);
and U6269 (N_6269,N_5835,N_5513);
nor U6270 (N_6270,N_5985,N_5716);
nand U6271 (N_6271,N_5895,N_5859);
nor U6272 (N_6272,N_5617,N_5755);
and U6273 (N_6273,N_5891,N_5878);
and U6274 (N_6274,N_5549,N_5818);
or U6275 (N_6275,N_5940,N_5548);
nor U6276 (N_6276,N_5779,N_5936);
nand U6277 (N_6277,N_5949,N_5827);
nor U6278 (N_6278,N_5608,N_5520);
and U6279 (N_6279,N_5962,N_5591);
xor U6280 (N_6280,N_5501,N_5551);
and U6281 (N_6281,N_5743,N_5560);
nand U6282 (N_6282,N_5554,N_5762);
and U6283 (N_6283,N_5587,N_5731);
or U6284 (N_6284,N_5857,N_5508);
nor U6285 (N_6285,N_5871,N_5542);
nand U6286 (N_6286,N_5593,N_5586);
and U6287 (N_6287,N_5572,N_5860);
nand U6288 (N_6288,N_5800,N_5960);
and U6289 (N_6289,N_5533,N_5662);
or U6290 (N_6290,N_5861,N_5844);
and U6291 (N_6291,N_5674,N_5590);
nor U6292 (N_6292,N_5501,N_5789);
and U6293 (N_6293,N_5903,N_5848);
nor U6294 (N_6294,N_5606,N_5696);
or U6295 (N_6295,N_5519,N_5746);
or U6296 (N_6296,N_5612,N_5842);
or U6297 (N_6297,N_5883,N_5688);
nor U6298 (N_6298,N_5813,N_5993);
nand U6299 (N_6299,N_5809,N_5674);
or U6300 (N_6300,N_5689,N_5564);
nand U6301 (N_6301,N_5806,N_5799);
nand U6302 (N_6302,N_5938,N_5987);
nor U6303 (N_6303,N_5906,N_5763);
nor U6304 (N_6304,N_5689,N_5749);
and U6305 (N_6305,N_5588,N_5558);
or U6306 (N_6306,N_5747,N_5757);
nor U6307 (N_6307,N_5646,N_5819);
or U6308 (N_6308,N_5871,N_5838);
and U6309 (N_6309,N_5942,N_5746);
nor U6310 (N_6310,N_5673,N_5690);
or U6311 (N_6311,N_5740,N_5774);
nand U6312 (N_6312,N_5774,N_5556);
nor U6313 (N_6313,N_5726,N_5817);
and U6314 (N_6314,N_5976,N_5646);
and U6315 (N_6315,N_5781,N_5518);
or U6316 (N_6316,N_5854,N_5579);
nor U6317 (N_6317,N_5956,N_5988);
nand U6318 (N_6318,N_5750,N_5612);
nor U6319 (N_6319,N_5766,N_5684);
nor U6320 (N_6320,N_5822,N_5785);
or U6321 (N_6321,N_5922,N_5935);
or U6322 (N_6322,N_5960,N_5771);
nor U6323 (N_6323,N_5691,N_5914);
or U6324 (N_6324,N_5960,N_5737);
or U6325 (N_6325,N_5619,N_5814);
or U6326 (N_6326,N_5576,N_5582);
or U6327 (N_6327,N_5532,N_5608);
nand U6328 (N_6328,N_5648,N_5560);
nor U6329 (N_6329,N_5757,N_5894);
nor U6330 (N_6330,N_5757,N_5808);
nand U6331 (N_6331,N_5610,N_5692);
or U6332 (N_6332,N_5610,N_5950);
xnor U6333 (N_6333,N_5724,N_5862);
xor U6334 (N_6334,N_5511,N_5910);
or U6335 (N_6335,N_5891,N_5736);
and U6336 (N_6336,N_5670,N_5779);
and U6337 (N_6337,N_5760,N_5676);
and U6338 (N_6338,N_5850,N_5506);
or U6339 (N_6339,N_5940,N_5919);
or U6340 (N_6340,N_5637,N_5619);
nor U6341 (N_6341,N_5945,N_5577);
or U6342 (N_6342,N_5730,N_5707);
nand U6343 (N_6343,N_5777,N_5995);
nand U6344 (N_6344,N_5622,N_5819);
and U6345 (N_6345,N_5760,N_5604);
nor U6346 (N_6346,N_5693,N_5939);
nor U6347 (N_6347,N_5891,N_5620);
xor U6348 (N_6348,N_5827,N_5527);
nor U6349 (N_6349,N_5859,N_5933);
nand U6350 (N_6350,N_5771,N_5897);
nor U6351 (N_6351,N_5899,N_5902);
nor U6352 (N_6352,N_5810,N_5758);
nor U6353 (N_6353,N_5595,N_5559);
or U6354 (N_6354,N_5819,N_5633);
or U6355 (N_6355,N_5564,N_5928);
nor U6356 (N_6356,N_5603,N_5709);
and U6357 (N_6357,N_5656,N_5543);
or U6358 (N_6358,N_5790,N_5644);
or U6359 (N_6359,N_5774,N_5580);
or U6360 (N_6360,N_5821,N_5583);
nand U6361 (N_6361,N_5587,N_5613);
nand U6362 (N_6362,N_5738,N_5649);
nand U6363 (N_6363,N_5860,N_5791);
nor U6364 (N_6364,N_5933,N_5731);
nand U6365 (N_6365,N_5906,N_5940);
nand U6366 (N_6366,N_5833,N_5647);
or U6367 (N_6367,N_5848,N_5582);
nand U6368 (N_6368,N_5600,N_5542);
and U6369 (N_6369,N_5687,N_5862);
nor U6370 (N_6370,N_5766,N_5930);
nor U6371 (N_6371,N_5612,N_5559);
nor U6372 (N_6372,N_5773,N_5920);
nor U6373 (N_6373,N_5969,N_5860);
or U6374 (N_6374,N_5582,N_5858);
and U6375 (N_6375,N_5892,N_5804);
nand U6376 (N_6376,N_5909,N_5665);
nor U6377 (N_6377,N_5890,N_5801);
or U6378 (N_6378,N_5995,N_5718);
nor U6379 (N_6379,N_5960,N_5580);
nand U6380 (N_6380,N_5918,N_5668);
nor U6381 (N_6381,N_5876,N_5556);
nor U6382 (N_6382,N_5800,N_5715);
nor U6383 (N_6383,N_5512,N_5798);
or U6384 (N_6384,N_5627,N_5800);
nand U6385 (N_6385,N_5866,N_5767);
and U6386 (N_6386,N_5820,N_5988);
and U6387 (N_6387,N_5800,N_5988);
nand U6388 (N_6388,N_5549,N_5547);
xnor U6389 (N_6389,N_5601,N_5807);
nor U6390 (N_6390,N_5530,N_5555);
xnor U6391 (N_6391,N_5866,N_5878);
nand U6392 (N_6392,N_5634,N_5993);
nor U6393 (N_6393,N_5541,N_5833);
and U6394 (N_6394,N_5588,N_5923);
nand U6395 (N_6395,N_5733,N_5598);
xnor U6396 (N_6396,N_5747,N_5627);
or U6397 (N_6397,N_5763,N_5997);
nor U6398 (N_6398,N_5570,N_5927);
and U6399 (N_6399,N_5851,N_5645);
nor U6400 (N_6400,N_5596,N_5731);
xor U6401 (N_6401,N_5821,N_5872);
or U6402 (N_6402,N_5612,N_5511);
nor U6403 (N_6403,N_5975,N_5804);
nand U6404 (N_6404,N_5880,N_5765);
nor U6405 (N_6405,N_5673,N_5551);
and U6406 (N_6406,N_5840,N_5573);
nor U6407 (N_6407,N_5623,N_5879);
and U6408 (N_6408,N_5848,N_5943);
nand U6409 (N_6409,N_5737,N_5657);
or U6410 (N_6410,N_5999,N_5609);
and U6411 (N_6411,N_5974,N_5721);
or U6412 (N_6412,N_5867,N_5644);
nand U6413 (N_6413,N_5786,N_5683);
or U6414 (N_6414,N_5802,N_5731);
or U6415 (N_6415,N_5812,N_5642);
xor U6416 (N_6416,N_5901,N_5809);
nor U6417 (N_6417,N_5958,N_5710);
and U6418 (N_6418,N_5658,N_5842);
nor U6419 (N_6419,N_5798,N_5974);
nor U6420 (N_6420,N_5703,N_5546);
or U6421 (N_6421,N_5632,N_5857);
nand U6422 (N_6422,N_5887,N_5989);
or U6423 (N_6423,N_5908,N_5631);
and U6424 (N_6424,N_5770,N_5713);
nand U6425 (N_6425,N_5730,N_5594);
or U6426 (N_6426,N_5860,N_5536);
nand U6427 (N_6427,N_5747,N_5522);
nor U6428 (N_6428,N_5836,N_5712);
nand U6429 (N_6429,N_5634,N_5959);
or U6430 (N_6430,N_5740,N_5629);
and U6431 (N_6431,N_5646,N_5857);
and U6432 (N_6432,N_5758,N_5946);
nand U6433 (N_6433,N_5588,N_5671);
and U6434 (N_6434,N_5893,N_5660);
and U6435 (N_6435,N_5775,N_5625);
and U6436 (N_6436,N_5669,N_5909);
nor U6437 (N_6437,N_5507,N_5706);
and U6438 (N_6438,N_5793,N_5645);
nor U6439 (N_6439,N_5907,N_5861);
or U6440 (N_6440,N_5773,N_5562);
or U6441 (N_6441,N_5961,N_5847);
or U6442 (N_6442,N_5786,N_5712);
and U6443 (N_6443,N_5758,N_5714);
nand U6444 (N_6444,N_5828,N_5836);
or U6445 (N_6445,N_5884,N_5509);
and U6446 (N_6446,N_5711,N_5701);
or U6447 (N_6447,N_5581,N_5708);
or U6448 (N_6448,N_5978,N_5909);
nand U6449 (N_6449,N_5651,N_5798);
and U6450 (N_6450,N_5697,N_5792);
nand U6451 (N_6451,N_5934,N_5850);
or U6452 (N_6452,N_5553,N_5608);
and U6453 (N_6453,N_5557,N_5953);
and U6454 (N_6454,N_5632,N_5952);
and U6455 (N_6455,N_5626,N_5904);
or U6456 (N_6456,N_5766,N_5948);
nor U6457 (N_6457,N_5937,N_5618);
nor U6458 (N_6458,N_5681,N_5643);
or U6459 (N_6459,N_5976,N_5526);
nand U6460 (N_6460,N_5750,N_5611);
nand U6461 (N_6461,N_5586,N_5639);
nand U6462 (N_6462,N_5637,N_5823);
nand U6463 (N_6463,N_5942,N_5592);
or U6464 (N_6464,N_5787,N_5916);
nand U6465 (N_6465,N_5606,N_5514);
nor U6466 (N_6466,N_5914,N_5849);
nor U6467 (N_6467,N_5729,N_5633);
and U6468 (N_6468,N_5656,N_5940);
nor U6469 (N_6469,N_5975,N_5974);
nor U6470 (N_6470,N_5582,N_5840);
nor U6471 (N_6471,N_5617,N_5542);
and U6472 (N_6472,N_5937,N_5795);
and U6473 (N_6473,N_5931,N_5680);
nand U6474 (N_6474,N_5708,N_5587);
xnor U6475 (N_6475,N_5830,N_5710);
or U6476 (N_6476,N_5998,N_5755);
xnor U6477 (N_6477,N_5626,N_5989);
and U6478 (N_6478,N_5723,N_5580);
and U6479 (N_6479,N_5699,N_5795);
or U6480 (N_6480,N_5721,N_5929);
and U6481 (N_6481,N_5618,N_5936);
nor U6482 (N_6482,N_5604,N_5781);
nor U6483 (N_6483,N_5695,N_5776);
nand U6484 (N_6484,N_5584,N_5549);
nand U6485 (N_6485,N_5578,N_5684);
or U6486 (N_6486,N_5873,N_5959);
nor U6487 (N_6487,N_5500,N_5669);
nand U6488 (N_6488,N_5599,N_5785);
nor U6489 (N_6489,N_5757,N_5769);
or U6490 (N_6490,N_5779,N_5868);
nor U6491 (N_6491,N_5821,N_5723);
nor U6492 (N_6492,N_5911,N_5547);
nand U6493 (N_6493,N_5731,N_5738);
or U6494 (N_6494,N_5644,N_5624);
and U6495 (N_6495,N_5518,N_5967);
nor U6496 (N_6496,N_5609,N_5789);
and U6497 (N_6497,N_5670,N_5680);
or U6498 (N_6498,N_5792,N_5838);
nand U6499 (N_6499,N_5614,N_5585);
and U6500 (N_6500,N_6441,N_6392);
nor U6501 (N_6501,N_6299,N_6166);
nand U6502 (N_6502,N_6195,N_6277);
nand U6503 (N_6503,N_6004,N_6152);
and U6504 (N_6504,N_6053,N_6282);
and U6505 (N_6505,N_6123,N_6258);
nor U6506 (N_6506,N_6481,N_6488);
or U6507 (N_6507,N_6240,N_6112);
nand U6508 (N_6508,N_6388,N_6080);
or U6509 (N_6509,N_6332,N_6070);
nand U6510 (N_6510,N_6171,N_6305);
or U6511 (N_6511,N_6413,N_6233);
nor U6512 (N_6512,N_6400,N_6414);
and U6513 (N_6513,N_6295,N_6106);
and U6514 (N_6514,N_6389,N_6269);
nand U6515 (N_6515,N_6293,N_6154);
or U6516 (N_6516,N_6463,N_6081);
nor U6517 (N_6517,N_6218,N_6022);
nand U6518 (N_6518,N_6329,N_6032);
or U6519 (N_6519,N_6102,N_6136);
nand U6520 (N_6520,N_6340,N_6460);
or U6521 (N_6521,N_6467,N_6067);
and U6522 (N_6522,N_6320,N_6003);
nor U6523 (N_6523,N_6058,N_6082);
or U6524 (N_6524,N_6242,N_6221);
xor U6525 (N_6525,N_6241,N_6380);
nor U6526 (N_6526,N_6177,N_6351);
or U6527 (N_6527,N_6087,N_6200);
nor U6528 (N_6528,N_6316,N_6279);
and U6529 (N_6529,N_6412,N_6182);
nand U6530 (N_6530,N_6122,N_6302);
or U6531 (N_6531,N_6077,N_6472);
and U6532 (N_6532,N_6193,N_6447);
nor U6533 (N_6533,N_6064,N_6104);
and U6534 (N_6534,N_6427,N_6033);
nor U6535 (N_6535,N_6446,N_6292);
nor U6536 (N_6536,N_6253,N_6317);
and U6537 (N_6537,N_6455,N_6274);
or U6538 (N_6538,N_6311,N_6084);
nand U6539 (N_6539,N_6284,N_6013);
nor U6540 (N_6540,N_6015,N_6006);
nand U6541 (N_6541,N_6155,N_6354);
nor U6542 (N_6542,N_6315,N_6150);
and U6543 (N_6543,N_6169,N_6301);
and U6544 (N_6544,N_6259,N_6217);
or U6545 (N_6545,N_6094,N_6156);
or U6546 (N_6546,N_6263,N_6191);
nor U6547 (N_6547,N_6403,N_6181);
nor U6548 (N_6548,N_6117,N_6345);
nand U6549 (N_6549,N_6050,N_6360);
xnor U6550 (N_6550,N_6344,N_6225);
or U6551 (N_6551,N_6348,N_6183);
nor U6552 (N_6552,N_6132,N_6237);
or U6553 (N_6553,N_6116,N_6339);
nor U6554 (N_6554,N_6027,N_6203);
and U6555 (N_6555,N_6436,N_6330);
nand U6556 (N_6556,N_6031,N_6044);
nand U6557 (N_6557,N_6484,N_6387);
nor U6558 (N_6558,N_6244,N_6465);
or U6559 (N_6559,N_6055,N_6100);
or U6560 (N_6560,N_6206,N_6493);
nor U6561 (N_6561,N_6395,N_6267);
or U6562 (N_6562,N_6452,N_6303);
nor U6563 (N_6563,N_6473,N_6135);
and U6564 (N_6564,N_6313,N_6223);
xnor U6565 (N_6565,N_6060,N_6337);
and U6566 (N_6566,N_6411,N_6280);
nor U6567 (N_6567,N_6246,N_6275);
or U6568 (N_6568,N_6017,N_6281);
nor U6569 (N_6569,N_6146,N_6023);
or U6570 (N_6570,N_6101,N_6083);
and U6571 (N_6571,N_6342,N_6066);
nor U6572 (N_6572,N_6393,N_6099);
nand U6573 (N_6573,N_6290,N_6390);
or U6574 (N_6574,N_6416,N_6434);
nor U6575 (N_6575,N_6459,N_6211);
or U6576 (N_6576,N_6334,N_6245);
nor U6577 (N_6577,N_6312,N_6347);
nand U6578 (N_6578,N_6196,N_6331);
or U6579 (N_6579,N_6034,N_6417);
or U6580 (N_6580,N_6318,N_6306);
or U6581 (N_6581,N_6139,N_6186);
or U6582 (N_6582,N_6212,N_6047);
and U6583 (N_6583,N_6103,N_6426);
nor U6584 (N_6584,N_6262,N_6376);
and U6585 (N_6585,N_6264,N_6418);
and U6586 (N_6586,N_6179,N_6046);
nand U6587 (N_6587,N_6238,N_6404);
nor U6588 (N_6588,N_6428,N_6073);
nand U6589 (N_6589,N_6197,N_6019);
nand U6590 (N_6590,N_6440,N_6439);
nand U6591 (N_6591,N_6420,N_6361);
nand U6592 (N_6592,N_6366,N_6375);
and U6593 (N_6593,N_6190,N_6283);
nor U6594 (N_6594,N_6325,N_6367);
nand U6595 (N_6595,N_6369,N_6466);
and U6596 (N_6596,N_6220,N_6498);
and U6597 (N_6597,N_6204,N_6054);
and U6598 (N_6598,N_6119,N_6343);
nand U6599 (N_6599,N_6297,N_6074);
nand U6600 (N_6600,N_6160,N_6296);
or U6601 (N_6601,N_6052,N_6443);
or U6602 (N_6602,N_6079,N_6114);
and U6603 (N_6603,N_6405,N_6268);
or U6604 (N_6604,N_6261,N_6391);
or U6605 (N_6605,N_6085,N_6232);
xor U6606 (N_6606,N_6321,N_6324);
nor U6607 (N_6607,N_6352,N_6071);
or U6608 (N_6608,N_6326,N_6185);
or U6609 (N_6609,N_6038,N_6062);
nor U6610 (N_6610,N_6250,N_6491);
or U6611 (N_6611,N_6453,N_6142);
or U6612 (N_6612,N_6454,N_6482);
nand U6613 (N_6613,N_6364,N_6000);
nand U6614 (N_6614,N_6368,N_6495);
nor U6615 (N_6615,N_6120,N_6239);
nand U6616 (N_6616,N_6162,N_6381);
and U6617 (N_6617,N_6021,N_6338);
and U6618 (N_6618,N_6188,N_6236);
and U6619 (N_6619,N_6307,N_6091);
nand U6620 (N_6620,N_6249,N_6230);
nor U6621 (N_6621,N_6202,N_6129);
nand U6622 (N_6622,N_6294,N_6149);
nor U6623 (N_6623,N_6068,N_6349);
or U6624 (N_6624,N_6143,N_6494);
and U6625 (N_6625,N_6430,N_6093);
nand U6626 (N_6626,N_6167,N_6134);
or U6627 (N_6627,N_6214,N_6172);
nor U6628 (N_6628,N_6399,N_6170);
or U6629 (N_6629,N_6398,N_6092);
nand U6630 (N_6630,N_6029,N_6096);
xnor U6631 (N_6631,N_6335,N_6045);
and U6632 (N_6632,N_6043,N_6438);
or U6633 (N_6633,N_6359,N_6018);
or U6634 (N_6634,N_6468,N_6433);
nand U6635 (N_6635,N_6041,N_6378);
and U6636 (N_6636,N_6346,N_6397);
nand U6637 (N_6637,N_6396,N_6379);
and U6638 (N_6638,N_6144,N_6291);
or U6639 (N_6639,N_6175,N_6161);
nand U6640 (N_6640,N_6108,N_6201);
nand U6641 (N_6641,N_6487,N_6141);
and U6642 (N_6642,N_6374,N_6247);
and U6643 (N_6643,N_6492,N_6355);
or U6644 (N_6644,N_6137,N_6222);
or U6645 (N_6645,N_6286,N_6304);
nand U6646 (N_6646,N_6298,N_6126);
xnor U6647 (N_6647,N_6048,N_6138);
and U6648 (N_6648,N_6386,N_6384);
nand U6649 (N_6649,N_6063,N_6159);
nand U6650 (N_6650,N_6252,N_6184);
or U6651 (N_6651,N_6121,N_6470);
or U6652 (N_6652,N_6219,N_6198);
or U6653 (N_6653,N_6051,N_6009);
and U6654 (N_6654,N_6229,N_6001);
nand U6655 (N_6655,N_6479,N_6231);
and U6656 (N_6656,N_6350,N_6435);
nor U6657 (N_6657,N_6042,N_6409);
nand U6658 (N_6658,N_6140,N_6464);
nor U6659 (N_6659,N_6109,N_6370);
nor U6660 (N_6660,N_6213,N_6012);
nor U6661 (N_6661,N_6444,N_6251);
or U6662 (N_6662,N_6028,N_6451);
nor U6663 (N_6663,N_6475,N_6278);
or U6664 (N_6664,N_6205,N_6078);
nor U6665 (N_6665,N_6097,N_6327);
or U6666 (N_6666,N_6007,N_6272);
and U6667 (N_6667,N_6497,N_6040);
or U6668 (N_6668,N_6477,N_6382);
nor U6669 (N_6669,N_6385,N_6025);
and U6670 (N_6670,N_6474,N_6228);
xnor U6671 (N_6671,N_6107,N_6158);
nor U6672 (N_6672,N_6131,N_6476);
or U6673 (N_6673,N_6133,N_6008);
nor U6674 (N_6674,N_6308,N_6128);
and U6675 (N_6675,N_6176,N_6059);
nor U6676 (N_6676,N_6310,N_6429);
nand U6677 (N_6677,N_6030,N_6088);
nor U6678 (N_6678,N_6147,N_6187);
nor U6679 (N_6679,N_6163,N_6377);
and U6680 (N_6680,N_6490,N_6069);
nand U6681 (N_6681,N_6151,N_6260);
or U6682 (N_6682,N_6394,N_6016);
and U6683 (N_6683,N_6153,N_6336);
and U6684 (N_6684,N_6289,N_6328);
and U6685 (N_6685,N_6148,N_6090);
and U6686 (N_6686,N_6363,N_6256);
nor U6687 (N_6687,N_6036,N_6026);
nand U6688 (N_6688,N_6424,N_6168);
or U6689 (N_6689,N_6180,N_6456);
and U6690 (N_6690,N_6450,N_6356);
and U6691 (N_6691,N_6020,N_6485);
nand U6692 (N_6692,N_6457,N_6118);
and U6693 (N_6693,N_6227,N_6471);
and U6694 (N_6694,N_6216,N_6049);
nand U6695 (N_6695,N_6265,N_6314);
nand U6696 (N_6696,N_6410,N_6437);
and U6697 (N_6697,N_6072,N_6127);
or U6698 (N_6698,N_6011,N_6111);
or U6699 (N_6699,N_6057,N_6319);
nor U6700 (N_6700,N_6266,N_6037);
and U6701 (N_6701,N_6421,N_6371);
and U6702 (N_6702,N_6415,N_6215);
nand U6703 (N_6703,N_6273,N_6365);
nor U6704 (N_6704,N_6483,N_6089);
nand U6705 (N_6705,N_6165,N_6445);
nand U6706 (N_6706,N_6014,N_6056);
and U6707 (N_6707,N_6234,N_6255);
nand U6708 (N_6708,N_6189,N_6362);
nand U6709 (N_6709,N_6486,N_6357);
or U6710 (N_6710,N_6407,N_6300);
and U6711 (N_6711,N_6401,N_6065);
nor U6712 (N_6712,N_6341,N_6105);
nor U6713 (N_6713,N_6192,N_6270);
xor U6714 (N_6714,N_6422,N_6210);
nand U6715 (N_6715,N_6431,N_6442);
nor U6716 (N_6716,N_6164,N_6499);
and U6717 (N_6717,N_6076,N_6035);
nor U6718 (N_6718,N_6496,N_6145);
nor U6719 (N_6719,N_6174,N_6208);
and U6720 (N_6720,N_6095,N_6207);
xor U6721 (N_6721,N_6408,N_6288);
nand U6722 (N_6722,N_6353,N_6173);
nand U6723 (N_6723,N_6402,N_6373);
or U6724 (N_6724,N_6098,N_6254);
nor U6725 (N_6725,N_6458,N_6480);
nand U6726 (N_6726,N_6243,N_6178);
nand U6727 (N_6727,N_6406,N_6248);
nand U6728 (N_6728,N_6271,N_6194);
or U6729 (N_6729,N_6489,N_6449);
nor U6730 (N_6730,N_6461,N_6423);
nor U6731 (N_6731,N_6209,N_6383);
or U6732 (N_6732,N_6322,N_6157);
or U6733 (N_6733,N_6419,N_6002);
and U6734 (N_6734,N_6024,N_6226);
and U6735 (N_6735,N_6113,N_6224);
or U6736 (N_6736,N_6309,N_6130);
nand U6737 (N_6737,N_6010,N_6358);
nand U6738 (N_6738,N_6061,N_6110);
nand U6739 (N_6739,N_6086,N_6235);
nand U6740 (N_6740,N_6075,N_6124);
nor U6741 (N_6741,N_6448,N_6199);
nand U6742 (N_6742,N_6005,N_6469);
nor U6743 (N_6743,N_6115,N_6432);
and U6744 (N_6744,N_6257,N_6276);
and U6745 (N_6745,N_6125,N_6323);
nand U6746 (N_6746,N_6039,N_6333);
nand U6747 (N_6747,N_6287,N_6372);
nand U6748 (N_6748,N_6285,N_6425);
and U6749 (N_6749,N_6462,N_6478);
nor U6750 (N_6750,N_6394,N_6300);
nand U6751 (N_6751,N_6066,N_6390);
nand U6752 (N_6752,N_6239,N_6312);
or U6753 (N_6753,N_6230,N_6226);
or U6754 (N_6754,N_6144,N_6294);
or U6755 (N_6755,N_6006,N_6430);
nand U6756 (N_6756,N_6040,N_6301);
or U6757 (N_6757,N_6332,N_6009);
or U6758 (N_6758,N_6380,N_6411);
nor U6759 (N_6759,N_6005,N_6445);
or U6760 (N_6760,N_6332,N_6048);
nor U6761 (N_6761,N_6316,N_6108);
nand U6762 (N_6762,N_6263,N_6330);
and U6763 (N_6763,N_6397,N_6110);
or U6764 (N_6764,N_6424,N_6033);
nand U6765 (N_6765,N_6273,N_6032);
and U6766 (N_6766,N_6374,N_6273);
or U6767 (N_6767,N_6311,N_6270);
and U6768 (N_6768,N_6169,N_6263);
or U6769 (N_6769,N_6049,N_6053);
nand U6770 (N_6770,N_6201,N_6037);
or U6771 (N_6771,N_6154,N_6413);
nand U6772 (N_6772,N_6019,N_6396);
or U6773 (N_6773,N_6133,N_6024);
nand U6774 (N_6774,N_6212,N_6263);
or U6775 (N_6775,N_6337,N_6054);
or U6776 (N_6776,N_6210,N_6330);
nor U6777 (N_6777,N_6204,N_6237);
nor U6778 (N_6778,N_6448,N_6237);
or U6779 (N_6779,N_6074,N_6457);
xor U6780 (N_6780,N_6106,N_6485);
and U6781 (N_6781,N_6098,N_6115);
or U6782 (N_6782,N_6495,N_6411);
and U6783 (N_6783,N_6283,N_6218);
nand U6784 (N_6784,N_6451,N_6274);
nand U6785 (N_6785,N_6425,N_6381);
and U6786 (N_6786,N_6392,N_6230);
nand U6787 (N_6787,N_6480,N_6206);
nor U6788 (N_6788,N_6342,N_6258);
nor U6789 (N_6789,N_6119,N_6431);
xnor U6790 (N_6790,N_6044,N_6405);
or U6791 (N_6791,N_6356,N_6485);
and U6792 (N_6792,N_6221,N_6188);
nand U6793 (N_6793,N_6440,N_6119);
and U6794 (N_6794,N_6036,N_6207);
nand U6795 (N_6795,N_6123,N_6465);
or U6796 (N_6796,N_6424,N_6294);
or U6797 (N_6797,N_6476,N_6185);
or U6798 (N_6798,N_6161,N_6225);
nand U6799 (N_6799,N_6039,N_6187);
nor U6800 (N_6800,N_6130,N_6157);
nor U6801 (N_6801,N_6005,N_6296);
nand U6802 (N_6802,N_6302,N_6362);
nand U6803 (N_6803,N_6414,N_6168);
nand U6804 (N_6804,N_6156,N_6289);
nor U6805 (N_6805,N_6115,N_6002);
and U6806 (N_6806,N_6052,N_6051);
nand U6807 (N_6807,N_6368,N_6162);
or U6808 (N_6808,N_6310,N_6450);
nand U6809 (N_6809,N_6143,N_6258);
nor U6810 (N_6810,N_6289,N_6479);
nand U6811 (N_6811,N_6163,N_6257);
nand U6812 (N_6812,N_6325,N_6337);
nor U6813 (N_6813,N_6282,N_6219);
nor U6814 (N_6814,N_6235,N_6400);
or U6815 (N_6815,N_6210,N_6154);
nand U6816 (N_6816,N_6336,N_6111);
nor U6817 (N_6817,N_6388,N_6281);
nor U6818 (N_6818,N_6244,N_6318);
and U6819 (N_6819,N_6210,N_6270);
and U6820 (N_6820,N_6207,N_6351);
nand U6821 (N_6821,N_6244,N_6388);
and U6822 (N_6822,N_6007,N_6296);
or U6823 (N_6823,N_6064,N_6487);
nor U6824 (N_6824,N_6069,N_6281);
nand U6825 (N_6825,N_6308,N_6072);
nor U6826 (N_6826,N_6245,N_6054);
nand U6827 (N_6827,N_6013,N_6447);
or U6828 (N_6828,N_6277,N_6094);
or U6829 (N_6829,N_6049,N_6351);
nor U6830 (N_6830,N_6078,N_6164);
and U6831 (N_6831,N_6191,N_6229);
or U6832 (N_6832,N_6357,N_6223);
nand U6833 (N_6833,N_6339,N_6111);
and U6834 (N_6834,N_6205,N_6319);
and U6835 (N_6835,N_6438,N_6229);
nor U6836 (N_6836,N_6009,N_6307);
nand U6837 (N_6837,N_6161,N_6212);
and U6838 (N_6838,N_6213,N_6164);
nand U6839 (N_6839,N_6169,N_6025);
or U6840 (N_6840,N_6409,N_6023);
or U6841 (N_6841,N_6218,N_6397);
or U6842 (N_6842,N_6336,N_6442);
and U6843 (N_6843,N_6252,N_6265);
or U6844 (N_6844,N_6347,N_6033);
xor U6845 (N_6845,N_6296,N_6234);
nor U6846 (N_6846,N_6018,N_6403);
and U6847 (N_6847,N_6116,N_6356);
or U6848 (N_6848,N_6302,N_6248);
and U6849 (N_6849,N_6157,N_6135);
xnor U6850 (N_6850,N_6267,N_6114);
and U6851 (N_6851,N_6113,N_6199);
nand U6852 (N_6852,N_6130,N_6310);
or U6853 (N_6853,N_6039,N_6061);
nand U6854 (N_6854,N_6033,N_6380);
or U6855 (N_6855,N_6154,N_6400);
and U6856 (N_6856,N_6166,N_6439);
nand U6857 (N_6857,N_6454,N_6171);
nor U6858 (N_6858,N_6022,N_6101);
nand U6859 (N_6859,N_6023,N_6301);
and U6860 (N_6860,N_6047,N_6327);
nor U6861 (N_6861,N_6169,N_6391);
nand U6862 (N_6862,N_6231,N_6259);
nand U6863 (N_6863,N_6145,N_6011);
or U6864 (N_6864,N_6145,N_6364);
nand U6865 (N_6865,N_6398,N_6421);
nand U6866 (N_6866,N_6477,N_6260);
and U6867 (N_6867,N_6465,N_6228);
nor U6868 (N_6868,N_6311,N_6044);
and U6869 (N_6869,N_6309,N_6253);
xor U6870 (N_6870,N_6224,N_6179);
or U6871 (N_6871,N_6016,N_6365);
nand U6872 (N_6872,N_6487,N_6479);
nor U6873 (N_6873,N_6296,N_6151);
and U6874 (N_6874,N_6434,N_6290);
and U6875 (N_6875,N_6152,N_6256);
nand U6876 (N_6876,N_6200,N_6431);
nand U6877 (N_6877,N_6312,N_6317);
and U6878 (N_6878,N_6449,N_6382);
or U6879 (N_6879,N_6042,N_6131);
and U6880 (N_6880,N_6179,N_6141);
and U6881 (N_6881,N_6473,N_6396);
and U6882 (N_6882,N_6410,N_6411);
or U6883 (N_6883,N_6038,N_6213);
nor U6884 (N_6884,N_6128,N_6023);
nand U6885 (N_6885,N_6276,N_6275);
and U6886 (N_6886,N_6125,N_6267);
nand U6887 (N_6887,N_6497,N_6418);
xor U6888 (N_6888,N_6389,N_6156);
or U6889 (N_6889,N_6400,N_6110);
or U6890 (N_6890,N_6429,N_6475);
or U6891 (N_6891,N_6099,N_6395);
nand U6892 (N_6892,N_6038,N_6045);
nand U6893 (N_6893,N_6196,N_6205);
nand U6894 (N_6894,N_6395,N_6323);
or U6895 (N_6895,N_6172,N_6127);
nand U6896 (N_6896,N_6253,N_6497);
nor U6897 (N_6897,N_6309,N_6212);
nor U6898 (N_6898,N_6075,N_6269);
and U6899 (N_6899,N_6481,N_6070);
or U6900 (N_6900,N_6015,N_6318);
and U6901 (N_6901,N_6095,N_6399);
and U6902 (N_6902,N_6069,N_6034);
or U6903 (N_6903,N_6249,N_6311);
and U6904 (N_6904,N_6417,N_6476);
nand U6905 (N_6905,N_6439,N_6455);
nand U6906 (N_6906,N_6052,N_6344);
nor U6907 (N_6907,N_6343,N_6338);
or U6908 (N_6908,N_6000,N_6426);
nor U6909 (N_6909,N_6366,N_6268);
nand U6910 (N_6910,N_6144,N_6224);
and U6911 (N_6911,N_6460,N_6061);
nor U6912 (N_6912,N_6014,N_6236);
nor U6913 (N_6913,N_6062,N_6022);
or U6914 (N_6914,N_6299,N_6399);
nand U6915 (N_6915,N_6376,N_6360);
nand U6916 (N_6916,N_6114,N_6199);
and U6917 (N_6917,N_6434,N_6333);
nor U6918 (N_6918,N_6339,N_6144);
xor U6919 (N_6919,N_6062,N_6116);
and U6920 (N_6920,N_6317,N_6238);
nand U6921 (N_6921,N_6324,N_6188);
nor U6922 (N_6922,N_6276,N_6304);
nand U6923 (N_6923,N_6143,N_6495);
and U6924 (N_6924,N_6455,N_6034);
nor U6925 (N_6925,N_6373,N_6260);
nand U6926 (N_6926,N_6004,N_6320);
and U6927 (N_6927,N_6021,N_6496);
nand U6928 (N_6928,N_6444,N_6094);
or U6929 (N_6929,N_6440,N_6487);
nor U6930 (N_6930,N_6254,N_6145);
nand U6931 (N_6931,N_6056,N_6316);
or U6932 (N_6932,N_6072,N_6191);
and U6933 (N_6933,N_6241,N_6153);
nor U6934 (N_6934,N_6169,N_6274);
or U6935 (N_6935,N_6350,N_6399);
or U6936 (N_6936,N_6023,N_6126);
nor U6937 (N_6937,N_6401,N_6349);
or U6938 (N_6938,N_6138,N_6006);
and U6939 (N_6939,N_6470,N_6203);
xor U6940 (N_6940,N_6349,N_6372);
and U6941 (N_6941,N_6102,N_6179);
or U6942 (N_6942,N_6477,N_6106);
or U6943 (N_6943,N_6005,N_6436);
nor U6944 (N_6944,N_6196,N_6197);
nand U6945 (N_6945,N_6011,N_6013);
nor U6946 (N_6946,N_6087,N_6431);
or U6947 (N_6947,N_6464,N_6310);
or U6948 (N_6948,N_6042,N_6290);
nor U6949 (N_6949,N_6401,N_6003);
nor U6950 (N_6950,N_6053,N_6201);
xor U6951 (N_6951,N_6385,N_6394);
or U6952 (N_6952,N_6441,N_6008);
and U6953 (N_6953,N_6012,N_6177);
nor U6954 (N_6954,N_6443,N_6149);
nor U6955 (N_6955,N_6059,N_6007);
nand U6956 (N_6956,N_6044,N_6003);
nor U6957 (N_6957,N_6113,N_6101);
nor U6958 (N_6958,N_6167,N_6411);
nand U6959 (N_6959,N_6266,N_6316);
nor U6960 (N_6960,N_6043,N_6413);
nor U6961 (N_6961,N_6288,N_6197);
and U6962 (N_6962,N_6239,N_6223);
and U6963 (N_6963,N_6209,N_6144);
nand U6964 (N_6964,N_6411,N_6192);
and U6965 (N_6965,N_6387,N_6202);
and U6966 (N_6966,N_6002,N_6095);
nor U6967 (N_6967,N_6223,N_6144);
nand U6968 (N_6968,N_6130,N_6223);
nand U6969 (N_6969,N_6247,N_6440);
or U6970 (N_6970,N_6193,N_6310);
and U6971 (N_6971,N_6228,N_6469);
nand U6972 (N_6972,N_6493,N_6413);
nand U6973 (N_6973,N_6156,N_6398);
and U6974 (N_6974,N_6106,N_6490);
nand U6975 (N_6975,N_6016,N_6018);
nand U6976 (N_6976,N_6320,N_6411);
or U6977 (N_6977,N_6193,N_6142);
or U6978 (N_6978,N_6259,N_6495);
and U6979 (N_6979,N_6235,N_6059);
nor U6980 (N_6980,N_6426,N_6178);
nor U6981 (N_6981,N_6244,N_6261);
nand U6982 (N_6982,N_6084,N_6030);
nor U6983 (N_6983,N_6005,N_6123);
nand U6984 (N_6984,N_6277,N_6034);
nand U6985 (N_6985,N_6445,N_6054);
xor U6986 (N_6986,N_6228,N_6481);
nand U6987 (N_6987,N_6310,N_6406);
or U6988 (N_6988,N_6167,N_6358);
nand U6989 (N_6989,N_6264,N_6078);
nand U6990 (N_6990,N_6371,N_6202);
and U6991 (N_6991,N_6313,N_6135);
and U6992 (N_6992,N_6340,N_6155);
nor U6993 (N_6993,N_6063,N_6413);
nor U6994 (N_6994,N_6248,N_6413);
and U6995 (N_6995,N_6493,N_6453);
nand U6996 (N_6996,N_6323,N_6278);
and U6997 (N_6997,N_6126,N_6300);
and U6998 (N_6998,N_6475,N_6101);
and U6999 (N_6999,N_6307,N_6086);
nor U7000 (N_7000,N_6813,N_6719);
nor U7001 (N_7001,N_6761,N_6980);
and U7002 (N_7002,N_6793,N_6577);
and U7003 (N_7003,N_6571,N_6915);
nor U7004 (N_7004,N_6704,N_6610);
and U7005 (N_7005,N_6946,N_6832);
nor U7006 (N_7006,N_6716,N_6994);
nor U7007 (N_7007,N_6865,N_6566);
or U7008 (N_7008,N_6609,N_6933);
nor U7009 (N_7009,N_6842,N_6876);
or U7010 (N_7010,N_6552,N_6673);
nor U7011 (N_7011,N_6968,N_6806);
or U7012 (N_7012,N_6991,N_6615);
or U7013 (N_7013,N_6530,N_6854);
nor U7014 (N_7014,N_6705,N_6618);
nand U7015 (N_7015,N_6712,N_6962);
and U7016 (N_7016,N_6599,N_6520);
nor U7017 (N_7017,N_6619,N_6906);
nand U7018 (N_7018,N_6836,N_6549);
nand U7019 (N_7019,N_6923,N_6846);
nor U7020 (N_7020,N_6623,N_6974);
nand U7021 (N_7021,N_6990,N_6844);
and U7022 (N_7022,N_6536,N_6722);
nand U7023 (N_7023,N_6714,N_6899);
or U7024 (N_7024,N_6872,N_6645);
and U7025 (N_7025,N_6878,N_6992);
or U7026 (N_7026,N_6829,N_6812);
nor U7027 (N_7027,N_6650,N_6871);
or U7028 (N_7028,N_6696,N_6734);
or U7029 (N_7029,N_6745,N_6819);
nor U7030 (N_7030,N_6922,N_6604);
or U7031 (N_7031,N_6797,N_6795);
and U7032 (N_7032,N_6694,N_6861);
or U7033 (N_7033,N_6746,N_6545);
and U7034 (N_7034,N_6572,N_6686);
and U7035 (N_7035,N_6807,N_6573);
nor U7036 (N_7036,N_6726,N_6943);
nand U7037 (N_7037,N_6900,N_6683);
and U7038 (N_7038,N_6788,N_6993);
and U7039 (N_7039,N_6699,N_6518);
and U7040 (N_7040,N_6730,N_6775);
or U7041 (N_7041,N_6748,N_6883);
xor U7042 (N_7042,N_6873,N_6798);
nand U7043 (N_7043,N_6939,N_6910);
or U7044 (N_7044,N_6856,N_6720);
nand U7045 (N_7045,N_6898,N_6998);
xor U7046 (N_7046,N_6759,N_6579);
and U7047 (N_7047,N_6786,N_6895);
nand U7048 (N_7048,N_6863,N_6710);
or U7049 (N_7049,N_6584,N_6676);
nand U7050 (N_7050,N_6517,N_6964);
nand U7051 (N_7051,N_6888,N_6987);
and U7052 (N_7052,N_6858,N_6791);
and U7053 (N_7053,N_6742,N_6560);
or U7054 (N_7054,N_6905,N_6516);
nor U7055 (N_7055,N_6612,N_6664);
or U7056 (N_7056,N_6736,N_6588);
and U7057 (N_7057,N_6866,N_6982);
xnor U7058 (N_7058,N_6592,N_6953);
nor U7059 (N_7059,N_6901,N_6521);
nor U7060 (N_7060,N_6654,N_6620);
nand U7061 (N_7061,N_6752,N_6638);
and U7062 (N_7062,N_6847,N_6697);
and U7063 (N_7063,N_6581,N_6624);
nand U7064 (N_7064,N_6892,N_6973);
or U7065 (N_7065,N_6862,N_6531);
nand U7066 (N_7066,N_6904,N_6631);
nor U7067 (N_7067,N_6784,N_6689);
and U7068 (N_7068,N_6978,N_6514);
nor U7069 (N_7069,N_6565,N_6838);
and U7070 (N_7070,N_6559,N_6702);
and U7071 (N_7071,N_6543,N_6525);
or U7072 (N_7072,N_6652,N_6695);
nand U7073 (N_7073,N_6938,N_6556);
nor U7074 (N_7074,N_6762,N_6988);
nor U7075 (N_7075,N_6680,N_6569);
or U7076 (N_7076,N_6504,N_6674);
nand U7077 (N_7077,N_6659,N_6582);
nand U7078 (N_7078,N_6586,N_6713);
and U7079 (N_7079,N_6541,N_6930);
nand U7080 (N_7080,N_6961,N_6502);
nor U7081 (N_7081,N_6526,N_6947);
and U7082 (N_7082,N_6542,N_6948);
and U7083 (N_7083,N_6550,N_6834);
nand U7084 (N_7084,N_6903,N_6537);
nor U7085 (N_7085,N_6692,N_6756);
or U7086 (N_7086,N_6755,N_6799);
nand U7087 (N_7087,N_6544,N_6907);
and U7088 (N_7088,N_6956,N_6877);
nor U7089 (N_7089,N_6849,N_6583);
xor U7090 (N_7090,N_6596,N_6882);
and U7091 (N_7091,N_6985,N_6796);
nor U7092 (N_7092,N_6663,N_6790);
and U7093 (N_7093,N_6954,N_6625);
nand U7094 (N_7094,N_6909,N_6794);
nand U7095 (N_7095,N_6926,N_6738);
nor U7096 (N_7096,N_6575,N_6669);
and U7097 (N_7097,N_6553,N_6647);
nor U7098 (N_7098,N_6920,N_6508);
and U7099 (N_7099,N_6833,N_6886);
and U7100 (N_7100,N_6934,N_6735);
or U7101 (N_7101,N_6787,N_6971);
and U7102 (N_7102,N_6658,N_6641);
nand U7103 (N_7103,N_6651,N_6608);
nor U7104 (N_7104,N_6598,N_6580);
or U7105 (N_7105,N_6678,N_6975);
and U7106 (N_7106,N_6955,N_6763);
nor U7107 (N_7107,N_6989,N_6808);
nor U7108 (N_7108,N_6519,N_6533);
nor U7109 (N_7109,N_6848,N_6845);
nor U7110 (N_7110,N_6958,N_6621);
or U7111 (N_7111,N_6839,N_6976);
xnor U7112 (N_7112,N_6887,N_6999);
or U7113 (N_7113,N_6523,N_6841);
nand U7114 (N_7114,N_6637,N_6614);
nand U7115 (N_7115,N_6595,N_6562);
nand U7116 (N_7116,N_6868,N_6657);
or U7117 (N_7117,N_6785,N_6966);
or U7118 (N_7118,N_6940,N_6707);
and U7119 (N_7119,N_6629,N_6715);
and U7120 (N_7120,N_6703,N_6660);
or U7121 (N_7121,N_6515,N_6779);
nand U7122 (N_7122,N_6731,N_6850);
and U7123 (N_7123,N_6532,N_6972);
and U7124 (N_7124,N_6805,N_6802);
and U7125 (N_7125,N_6607,N_6774);
or U7126 (N_7126,N_6733,N_6600);
nor U7127 (N_7127,N_6950,N_6995);
nor U7128 (N_7128,N_6820,N_6548);
or U7129 (N_7129,N_6666,N_6897);
and U7130 (N_7130,N_6709,N_6636);
nand U7131 (N_7131,N_6894,N_6935);
and U7132 (N_7132,N_6911,N_6821);
nor U7133 (N_7133,N_6632,N_6587);
and U7134 (N_7134,N_6981,N_6741);
or U7135 (N_7135,N_6538,N_6814);
xnor U7136 (N_7136,N_6853,N_6546);
nor U7137 (N_7137,N_6593,N_6815);
nor U7138 (N_7138,N_6648,N_6606);
and U7139 (N_7139,N_6800,N_6949);
and U7140 (N_7140,N_6524,N_6749);
or U7141 (N_7141,N_6723,N_6857);
and U7142 (N_7142,N_6792,N_6732);
or U7143 (N_7143,N_6568,N_6500);
nand U7144 (N_7144,N_6701,N_6855);
or U7145 (N_7145,N_6729,N_6564);
nand U7146 (N_7146,N_6661,N_6529);
and U7147 (N_7147,N_6522,N_6574);
and U7148 (N_7148,N_6916,N_6567);
xor U7149 (N_7149,N_6758,N_6768);
and U7150 (N_7150,N_6662,N_6879);
or U7151 (N_7151,N_6851,N_6936);
and U7152 (N_7152,N_6890,N_6534);
and U7153 (N_7153,N_6773,N_6557);
or U7154 (N_7154,N_6668,N_6893);
nand U7155 (N_7155,N_6983,N_6835);
and U7156 (N_7156,N_6816,N_6700);
xnor U7157 (N_7157,N_6764,N_6728);
nand U7158 (N_7158,N_6881,N_6919);
nor U7159 (N_7159,N_6507,N_6843);
and U7160 (N_7160,N_6670,N_6765);
nor U7161 (N_7161,N_6769,N_6766);
nand U7162 (N_7162,N_6688,N_6511);
and U7163 (N_7163,N_6914,N_6644);
and U7164 (N_7164,N_6590,N_6594);
and U7165 (N_7165,N_6864,N_6576);
or U7166 (N_7166,N_6750,N_6928);
xnor U7167 (N_7167,N_6611,N_6945);
and U7168 (N_7168,N_6602,N_6852);
and U7169 (N_7169,N_6503,N_6740);
and U7170 (N_7170,N_6667,N_6739);
and U7171 (N_7171,N_6628,N_6921);
and U7172 (N_7172,N_6528,N_6831);
nor U7173 (N_7173,N_6630,N_6721);
or U7174 (N_7174,N_6937,N_6957);
nor U7175 (N_7175,N_6917,N_6908);
and U7176 (N_7176,N_6711,N_6770);
nand U7177 (N_7177,N_6967,N_6760);
or U7178 (N_7178,N_6969,N_6626);
xor U7179 (N_7179,N_6984,N_6941);
and U7180 (N_7180,N_6540,N_6656);
or U7181 (N_7181,N_6642,N_6912);
or U7182 (N_7182,N_6591,N_6783);
nor U7183 (N_7183,N_6874,N_6627);
xnor U7184 (N_7184,N_6724,N_6727);
or U7185 (N_7185,N_6605,N_6810);
or U7186 (N_7186,N_6558,N_6860);
nand U7187 (N_7187,N_6776,N_6634);
nand U7188 (N_7188,N_6506,N_6554);
and U7189 (N_7189,N_6555,N_6589);
and U7190 (N_7190,N_6837,N_6649);
xor U7191 (N_7191,N_6687,N_6951);
nand U7192 (N_7192,N_6809,N_6782);
nor U7193 (N_7193,N_6828,N_6677);
or U7194 (N_7194,N_6944,N_6826);
or U7195 (N_7195,N_6977,N_6959);
nor U7196 (N_7196,N_6927,N_6902);
and U7197 (N_7197,N_6781,N_6771);
nor U7198 (N_7198,N_6918,N_6698);
nand U7199 (N_7199,N_6747,N_6965);
and U7200 (N_7200,N_6640,N_6880);
and U7201 (N_7201,N_6924,N_6639);
nand U7202 (N_7202,N_6743,N_6867);
and U7203 (N_7203,N_6803,N_6585);
nand U7204 (N_7204,N_6603,N_6859);
nor U7205 (N_7205,N_6622,N_6811);
or U7206 (N_7206,N_6718,N_6960);
nor U7207 (N_7207,N_6690,N_6633);
or U7208 (N_7208,N_6996,N_6597);
or U7209 (N_7209,N_6870,N_6840);
or U7210 (N_7210,N_6801,N_6535);
and U7211 (N_7211,N_6684,N_6942);
nand U7212 (N_7212,N_6643,N_6737);
or U7213 (N_7213,N_6997,N_6913);
nor U7214 (N_7214,N_6635,N_6963);
nor U7215 (N_7215,N_6753,N_6932);
and U7216 (N_7216,N_6706,N_6789);
nand U7217 (N_7217,N_6757,N_6925);
nand U7218 (N_7218,N_6527,N_6617);
or U7219 (N_7219,N_6754,N_6681);
nor U7220 (N_7220,N_6772,N_6601);
and U7221 (N_7221,N_6561,N_6505);
or U7222 (N_7222,N_6679,N_6780);
or U7223 (N_7223,N_6693,N_6818);
nor U7224 (N_7224,N_6875,N_6891);
and U7225 (N_7225,N_6929,N_6725);
nor U7226 (N_7226,N_6970,N_6884);
and U7227 (N_7227,N_6889,N_6767);
and U7228 (N_7228,N_6513,N_6896);
nor U7229 (N_7229,N_6744,N_6616);
and U7230 (N_7230,N_6563,N_6827);
or U7231 (N_7231,N_6671,N_6825);
nor U7232 (N_7232,N_6539,N_6979);
or U7233 (N_7233,N_6685,N_6869);
nor U7234 (N_7234,N_6665,N_6952);
and U7235 (N_7235,N_6509,N_6682);
nor U7236 (N_7236,N_6501,N_6675);
or U7237 (N_7237,N_6512,N_6822);
nor U7238 (N_7238,N_6547,N_6570);
nand U7239 (N_7239,N_6510,N_6817);
and U7240 (N_7240,N_6885,N_6578);
and U7241 (N_7241,N_6986,N_6778);
or U7242 (N_7242,N_6717,N_6751);
and U7243 (N_7243,N_6823,N_6708);
nand U7244 (N_7244,N_6804,N_6646);
or U7245 (N_7245,N_6830,N_6824);
nor U7246 (N_7246,N_6691,N_6655);
nand U7247 (N_7247,N_6672,N_6653);
or U7248 (N_7248,N_6777,N_6613);
or U7249 (N_7249,N_6551,N_6931);
or U7250 (N_7250,N_6618,N_6967);
nand U7251 (N_7251,N_6924,N_6719);
nor U7252 (N_7252,N_6686,N_6767);
nor U7253 (N_7253,N_6745,N_6541);
nand U7254 (N_7254,N_6573,N_6727);
and U7255 (N_7255,N_6964,N_6506);
and U7256 (N_7256,N_6510,N_6747);
and U7257 (N_7257,N_6761,N_6548);
or U7258 (N_7258,N_6616,N_6838);
nor U7259 (N_7259,N_6653,N_6933);
nor U7260 (N_7260,N_6977,N_6580);
and U7261 (N_7261,N_6724,N_6592);
and U7262 (N_7262,N_6636,N_6574);
and U7263 (N_7263,N_6994,N_6652);
nand U7264 (N_7264,N_6748,N_6784);
nor U7265 (N_7265,N_6894,N_6632);
or U7266 (N_7266,N_6724,N_6874);
nand U7267 (N_7267,N_6778,N_6968);
nor U7268 (N_7268,N_6997,N_6559);
nand U7269 (N_7269,N_6592,N_6923);
nor U7270 (N_7270,N_6981,N_6894);
nand U7271 (N_7271,N_6807,N_6515);
nor U7272 (N_7272,N_6822,N_6741);
nand U7273 (N_7273,N_6793,N_6760);
nor U7274 (N_7274,N_6664,N_6657);
nand U7275 (N_7275,N_6868,N_6731);
or U7276 (N_7276,N_6970,N_6655);
nor U7277 (N_7277,N_6561,N_6508);
nand U7278 (N_7278,N_6841,N_6825);
or U7279 (N_7279,N_6865,N_6963);
and U7280 (N_7280,N_6834,N_6956);
nand U7281 (N_7281,N_6974,N_6888);
and U7282 (N_7282,N_6689,N_6715);
nand U7283 (N_7283,N_6995,N_6646);
nand U7284 (N_7284,N_6884,N_6895);
nand U7285 (N_7285,N_6708,N_6505);
nor U7286 (N_7286,N_6681,N_6832);
and U7287 (N_7287,N_6889,N_6682);
or U7288 (N_7288,N_6797,N_6671);
nor U7289 (N_7289,N_6849,N_6611);
and U7290 (N_7290,N_6683,N_6898);
nor U7291 (N_7291,N_6993,N_6822);
nand U7292 (N_7292,N_6863,N_6518);
and U7293 (N_7293,N_6833,N_6726);
and U7294 (N_7294,N_6939,N_6941);
and U7295 (N_7295,N_6956,N_6711);
or U7296 (N_7296,N_6993,N_6507);
nor U7297 (N_7297,N_6764,N_6720);
nand U7298 (N_7298,N_6599,N_6561);
and U7299 (N_7299,N_6774,N_6938);
nor U7300 (N_7300,N_6769,N_6573);
nand U7301 (N_7301,N_6628,N_6622);
or U7302 (N_7302,N_6514,N_6537);
or U7303 (N_7303,N_6995,N_6873);
or U7304 (N_7304,N_6768,N_6707);
nor U7305 (N_7305,N_6546,N_6778);
and U7306 (N_7306,N_6784,N_6567);
nand U7307 (N_7307,N_6668,N_6758);
nor U7308 (N_7308,N_6620,N_6542);
or U7309 (N_7309,N_6603,N_6620);
xnor U7310 (N_7310,N_6772,N_6907);
nor U7311 (N_7311,N_6510,N_6622);
or U7312 (N_7312,N_6525,N_6732);
or U7313 (N_7313,N_6812,N_6642);
nor U7314 (N_7314,N_6962,N_6742);
nand U7315 (N_7315,N_6768,N_6622);
nand U7316 (N_7316,N_6699,N_6656);
or U7317 (N_7317,N_6769,N_6702);
nor U7318 (N_7318,N_6788,N_6791);
or U7319 (N_7319,N_6918,N_6753);
or U7320 (N_7320,N_6953,N_6879);
nor U7321 (N_7321,N_6947,N_6653);
and U7322 (N_7322,N_6643,N_6552);
nor U7323 (N_7323,N_6742,N_6717);
or U7324 (N_7324,N_6731,N_6650);
xor U7325 (N_7325,N_6769,N_6849);
or U7326 (N_7326,N_6709,N_6528);
or U7327 (N_7327,N_6509,N_6879);
nor U7328 (N_7328,N_6912,N_6842);
and U7329 (N_7329,N_6873,N_6692);
and U7330 (N_7330,N_6621,N_6911);
nor U7331 (N_7331,N_6583,N_6940);
nand U7332 (N_7332,N_6525,N_6662);
nor U7333 (N_7333,N_6513,N_6956);
and U7334 (N_7334,N_6590,N_6839);
nand U7335 (N_7335,N_6677,N_6736);
or U7336 (N_7336,N_6709,N_6816);
nor U7337 (N_7337,N_6742,N_6811);
or U7338 (N_7338,N_6596,N_6840);
or U7339 (N_7339,N_6668,N_6652);
or U7340 (N_7340,N_6717,N_6655);
nand U7341 (N_7341,N_6658,N_6908);
nor U7342 (N_7342,N_6672,N_6951);
or U7343 (N_7343,N_6744,N_6866);
nand U7344 (N_7344,N_6819,N_6553);
nand U7345 (N_7345,N_6602,N_6897);
nor U7346 (N_7346,N_6711,N_6805);
nor U7347 (N_7347,N_6890,N_6696);
or U7348 (N_7348,N_6810,N_6841);
and U7349 (N_7349,N_6766,N_6899);
nor U7350 (N_7350,N_6720,N_6620);
nand U7351 (N_7351,N_6984,N_6680);
xnor U7352 (N_7352,N_6672,N_6925);
or U7353 (N_7353,N_6553,N_6601);
nor U7354 (N_7354,N_6962,N_6790);
nand U7355 (N_7355,N_6764,N_6836);
nor U7356 (N_7356,N_6933,N_6849);
nor U7357 (N_7357,N_6649,N_6818);
or U7358 (N_7358,N_6544,N_6969);
nor U7359 (N_7359,N_6900,N_6762);
or U7360 (N_7360,N_6662,N_6633);
xnor U7361 (N_7361,N_6871,N_6969);
and U7362 (N_7362,N_6681,N_6652);
and U7363 (N_7363,N_6837,N_6813);
and U7364 (N_7364,N_6948,N_6820);
nand U7365 (N_7365,N_6541,N_6758);
and U7366 (N_7366,N_6749,N_6618);
or U7367 (N_7367,N_6693,N_6735);
or U7368 (N_7368,N_6813,N_6824);
and U7369 (N_7369,N_6878,N_6658);
and U7370 (N_7370,N_6983,N_6912);
or U7371 (N_7371,N_6585,N_6812);
nand U7372 (N_7372,N_6946,N_6595);
nor U7373 (N_7373,N_6980,N_6896);
nor U7374 (N_7374,N_6682,N_6818);
and U7375 (N_7375,N_6794,N_6821);
nand U7376 (N_7376,N_6814,N_6862);
nor U7377 (N_7377,N_6544,N_6758);
nand U7378 (N_7378,N_6778,N_6594);
xor U7379 (N_7379,N_6549,N_6847);
nand U7380 (N_7380,N_6869,N_6550);
nand U7381 (N_7381,N_6772,N_6513);
nor U7382 (N_7382,N_6938,N_6585);
nor U7383 (N_7383,N_6749,N_6984);
xor U7384 (N_7384,N_6822,N_6614);
or U7385 (N_7385,N_6921,N_6984);
nand U7386 (N_7386,N_6532,N_6982);
or U7387 (N_7387,N_6725,N_6928);
nand U7388 (N_7388,N_6689,N_6808);
and U7389 (N_7389,N_6832,N_6933);
or U7390 (N_7390,N_6582,N_6906);
nand U7391 (N_7391,N_6592,N_6713);
nand U7392 (N_7392,N_6871,N_6770);
nand U7393 (N_7393,N_6893,N_6876);
or U7394 (N_7394,N_6817,N_6798);
or U7395 (N_7395,N_6500,N_6881);
xor U7396 (N_7396,N_6913,N_6988);
nand U7397 (N_7397,N_6742,N_6934);
nand U7398 (N_7398,N_6853,N_6634);
nand U7399 (N_7399,N_6545,N_6736);
xor U7400 (N_7400,N_6557,N_6645);
and U7401 (N_7401,N_6865,N_6994);
nand U7402 (N_7402,N_6610,N_6594);
nand U7403 (N_7403,N_6557,N_6949);
nor U7404 (N_7404,N_6960,N_6908);
nand U7405 (N_7405,N_6952,N_6857);
nor U7406 (N_7406,N_6813,N_6782);
or U7407 (N_7407,N_6520,N_6650);
nor U7408 (N_7408,N_6516,N_6725);
nand U7409 (N_7409,N_6727,N_6795);
and U7410 (N_7410,N_6955,N_6984);
nand U7411 (N_7411,N_6866,N_6832);
nand U7412 (N_7412,N_6901,N_6519);
or U7413 (N_7413,N_6563,N_6925);
and U7414 (N_7414,N_6748,N_6977);
nor U7415 (N_7415,N_6640,N_6701);
or U7416 (N_7416,N_6813,N_6909);
and U7417 (N_7417,N_6808,N_6901);
nor U7418 (N_7418,N_6983,N_6618);
or U7419 (N_7419,N_6962,N_6771);
nand U7420 (N_7420,N_6944,N_6722);
nor U7421 (N_7421,N_6564,N_6773);
or U7422 (N_7422,N_6947,N_6641);
or U7423 (N_7423,N_6626,N_6593);
or U7424 (N_7424,N_6712,N_6821);
and U7425 (N_7425,N_6895,N_6879);
and U7426 (N_7426,N_6530,N_6532);
and U7427 (N_7427,N_6773,N_6994);
nand U7428 (N_7428,N_6767,N_6976);
and U7429 (N_7429,N_6525,N_6673);
nand U7430 (N_7430,N_6711,N_6522);
nor U7431 (N_7431,N_6787,N_6948);
and U7432 (N_7432,N_6699,N_6675);
or U7433 (N_7433,N_6913,N_6724);
or U7434 (N_7434,N_6579,N_6919);
nand U7435 (N_7435,N_6789,N_6834);
or U7436 (N_7436,N_6642,N_6846);
or U7437 (N_7437,N_6699,N_6743);
nor U7438 (N_7438,N_6898,N_6618);
or U7439 (N_7439,N_6969,N_6753);
or U7440 (N_7440,N_6960,N_6662);
and U7441 (N_7441,N_6878,N_6704);
nand U7442 (N_7442,N_6915,N_6846);
and U7443 (N_7443,N_6576,N_6643);
or U7444 (N_7444,N_6549,N_6949);
or U7445 (N_7445,N_6938,N_6674);
and U7446 (N_7446,N_6781,N_6796);
and U7447 (N_7447,N_6948,N_6607);
nand U7448 (N_7448,N_6791,N_6984);
or U7449 (N_7449,N_6906,N_6715);
and U7450 (N_7450,N_6562,N_6634);
nor U7451 (N_7451,N_6602,N_6606);
and U7452 (N_7452,N_6555,N_6547);
nand U7453 (N_7453,N_6938,N_6950);
xnor U7454 (N_7454,N_6971,N_6910);
and U7455 (N_7455,N_6759,N_6705);
and U7456 (N_7456,N_6899,N_6809);
and U7457 (N_7457,N_6796,N_6905);
and U7458 (N_7458,N_6781,N_6903);
or U7459 (N_7459,N_6549,N_6956);
nand U7460 (N_7460,N_6987,N_6659);
and U7461 (N_7461,N_6865,N_6679);
nand U7462 (N_7462,N_6797,N_6843);
and U7463 (N_7463,N_6574,N_6748);
nand U7464 (N_7464,N_6753,N_6931);
or U7465 (N_7465,N_6826,N_6709);
or U7466 (N_7466,N_6663,N_6718);
or U7467 (N_7467,N_6928,N_6679);
and U7468 (N_7468,N_6551,N_6823);
nor U7469 (N_7469,N_6898,N_6835);
nand U7470 (N_7470,N_6548,N_6568);
and U7471 (N_7471,N_6587,N_6854);
or U7472 (N_7472,N_6663,N_6909);
or U7473 (N_7473,N_6729,N_6745);
nor U7474 (N_7474,N_6829,N_6697);
and U7475 (N_7475,N_6664,N_6695);
or U7476 (N_7476,N_6743,N_6783);
or U7477 (N_7477,N_6803,N_6896);
nand U7478 (N_7478,N_6581,N_6779);
or U7479 (N_7479,N_6511,N_6767);
nand U7480 (N_7480,N_6771,N_6949);
or U7481 (N_7481,N_6566,N_6887);
nor U7482 (N_7482,N_6891,N_6657);
nor U7483 (N_7483,N_6819,N_6780);
nor U7484 (N_7484,N_6732,N_6712);
nor U7485 (N_7485,N_6676,N_6572);
or U7486 (N_7486,N_6588,N_6796);
nand U7487 (N_7487,N_6755,N_6653);
or U7488 (N_7488,N_6532,N_6825);
or U7489 (N_7489,N_6624,N_6904);
and U7490 (N_7490,N_6987,N_6648);
nand U7491 (N_7491,N_6709,N_6611);
or U7492 (N_7492,N_6516,N_6931);
nand U7493 (N_7493,N_6933,N_6548);
or U7494 (N_7494,N_6797,N_6677);
and U7495 (N_7495,N_6613,N_6547);
or U7496 (N_7496,N_6779,N_6887);
or U7497 (N_7497,N_6577,N_6919);
nand U7498 (N_7498,N_6684,N_6598);
and U7499 (N_7499,N_6763,N_6531);
nor U7500 (N_7500,N_7429,N_7208);
and U7501 (N_7501,N_7310,N_7067);
nand U7502 (N_7502,N_7283,N_7356);
and U7503 (N_7503,N_7244,N_7224);
or U7504 (N_7504,N_7021,N_7226);
nand U7505 (N_7505,N_7345,N_7033);
or U7506 (N_7506,N_7420,N_7426);
xor U7507 (N_7507,N_7452,N_7129);
nor U7508 (N_7508,N_7247,N_7222);
and U7509 (N_7509,N_7455,N_7489);
xor U7510 (N_7510,N_7256,N_7187);
or U7511 (N_7511,N_7272,N_7087);
nor U7512 (N_7512,N_7194,N_7182);
nor U7513 (N_7513,N_7269,N_7109);
and U7514 (N_7514,N_7495,N_7232);
and U7515 (N_7515,N_7442,N_7395);
nor U7516 (N_7516,N_7110,N_7064);
nor U7517 (N_7517,N_7173,N_7276);
nor U7518 (N_7518,N_7104,N_7063);
and U7519 (N_7519,N_7186,N_7282);
nand U7520 (N_7520,N_7262,N_7013);
or U7521 (N_7521,N_7046,N_7254);
and U7522 (N_7522,N_7462,N_7150);
or U7523 (N_7523,N_7170,N_7080);
or U7524 (N_7524,N_7294,N_7156);
nand U7525 (N_7525,N_7135,N_7003);
nand U7526 (N_7526,N_7327,N_7465);
nor U7527 (N_7527,N_7311,N_7346);
nand U7528 (N_7528,N_7120,N_7373);
xor U7529 (N_7529,N_7088,N_7390);
nand U7530 (N_7530,N_7062,N_7086);
nand U7531 (N_7531,N_7306,N_7301);
nor U7532 (N_7532,N_7317,N_7212);
xor U7533 (N_7533,N_7202,N_7409);
nand U7534 (N_7534,N_7281,N_7121);
xor U7535 (N_7535,N_7023,N_7319);
and U7536 (N_7536,N_7443,N_7148);
and U7537 (N_7537,N_7467,N_7011);
and U7538 (N_7538,N_7338,N_7027);
nand U7539 (N_7539,N_7153,N_7466);
or U7540 (N_7540,N_7459,N_7043);
nand U7541 (N_7541,N_7270,N_7217);
nor U7542 (N_7542,N_7246,N_7180);
and U7543 (N_7543,N_7491,N_7298);
nor U7544 (N_7544,N_7201,N_7478);
and U7545 (N_7545,N_7130,N_7024);
nand U7546 (N_7546,N_7206,N_7075);
nand U7547 (N_7547,N_7322,N_7077);
or U7548 (N_7548,N_7030,N_7248);
or U7549 (N_7549,N_7353,N_7473);
nor U7550 (N_7550,N_7387,N_7348);
and U7551 (N_7551,N_7111,N_7190);
and U7552 (N_7552,N_7259,N_7488);
or U7553 (N_7553,N_7384,N_7060);
or U7554 (N_7554,N_7159,N_7393);
or U7555 (N_7555,N_7421,N_7157);
nand U7556 (N_7556,N_7496,N_7287);
and U7557 (N_7557,N_7108,N_7475);
nor U7558 (N_7558,N_7418,N_7441);
nand U7559 (N_7559,N_7470,N_7131);
and U7560 (N_7560,N_7040,N_7017);
or U7561 (N_7561,N_7499,N_7242);
or U7562 (N_7562,N_7330,N_7307);
nor U7563 (N_7563,N_7410,N_7260);
nor U7564 (N_7564,N_7385,N_7227);
and U7565 (N_7565,N_7169,N_7084);
or U7566 (N_7566,N_7302,N_7101);
or U7567 (N_7567,N_7050,N_7422);
nor U7568 (N_7568,N_7451,N_7048);
or U7569 (N_7569,N_7095,N_7207);
nor U7570 (N_7570,N_7320,N_7263);
nor U7571 (N_7571,N_7349,N_7402);
or U7572 (N_7572,N_7364,N_7141);
and U7573 (N_7573,N_7144,N_7461);
or U7574 (N_7574,N_7371,N_7396);
nand U7575 (N_7575,N_7274,N_7031);
and U7576 (N_7576,N_7012,N_7070);
or U7577 (N_7577,N_7085,N_7204);
nand U7578 (N_7578,N_7160,N_7367);
xnor U7579 (N_7579,N_7229,N_7125);
nor U7580 (N_7580,N_7477,N_7342);
or U7581 (N_7581,N_7337,N_7325);
nor U7582 (N_7582,N_7164,N_7264);
nand U7583 (N_7583,N_7236,N_7333);
and U7584 (N_7584,N_7097,N_7008);
and U7585 (N_7585,N_7380,N_7009);
and U7586 (N_7586,N_7341,N_7365);
and U7587 (N_7587,N_7428,N_7216);
nand U7588 (N_7588,N_7436,N_7412);
and U7589 (N_7589,N_7126,N_7430);
and U7590 (N_7590,N_7056,N_7010);
or U7591 (N_7591,N_7432,N_7329);
or U7592 (N_7592,N_7123,N_7273);
and U7593 (N_7593,N_7146,N_7291);
nor U7594 (N_7594,N_7362,N_7416);
nand U7595 (N_7595,N_7018,N_7474);
nor U7596 (N_7596,N_7168,N_7147);
nor U7597 (N_7597,N_7230,N_7458);
or U7598 (N_7598,N_7163,N_7026);
xor U7599 (N_7599,N_7357,N_7136);
nand U7600 (N_7600,N_7460,N_7400);
nand U7601 (N_7601,N_7339,N_7425);
nand U7602 (N_7602,N_7280,N_7332);
or U7603 (N_7603,N_7198,N_7482);
nand U7604 (N_7604,N_7038,N_7007);
and U7605 (N_7605,N_7486,N_7480);
or U7606 (N_7606,N_7231,N_7044);
and U7607 (N_7607,N_7293,N_7028);
nor U7608 (N_7608,N_7149,N_7092);
nand U7609 (N_7609,N_7255,N_7392);
nor U7610 (N_7610,N_7289,N_7314);
or U7611 (N_7611,N_7331,N_7116);
and U7612 (N_7612,N_7360,N_7200);
nor U7613 (N_7613,N_7389,N_7343);
or U7614 (N_7614,N_7447,N_7174);
xor U7615 (N_7615,N_7464,N_7142);
and U7616 (N_7616,N_7408,N_7446);
nor U7617 (N_7617,N_7424,N_7350);
or U7618 (N_7618,N_7078,N_7098);
xor U7619 (N_7619,N_7093,N_7191);
and U7620 (N_7620,N_7020,N_7074);
and U7621 (N_7621,N_7165,N_7195);
nand U7622 (N_7622,N_7450,N_7181);
nand U7623 (N_7623,N_7241,N_7223);
nand U7624 (N_7624,N_7277,N_7225);
or U7625 (N_7625,N_7411,N_7415);
nor U7626 (N_7626,N_7266,N_7154);
or U7627 (N_7627,N_7440,N_7398);
nor U7628 (N_7628,N_7381,N_7113);
nor U7629 (N_7629,N_7404,N_7234);
nor U7630 (N_7630,N_7041,N_7453);
nand U7631 (N_7631,N_7284,N_7279);
nand U7632 (N_7632,N_7036,N_7361);
and U7633 (N_7633,N_7472,N_7072);
xor U7634 (N_7634,N_7312,N_7414);
and U7635 (N_7635,N_7107,N_7133);
nor U7636 (N_7636,N_7315,N_7448);
or U7637 (N_7637,N_7444,N_7347);
nand U7638 (N_7638,N_7145,N_7445);
and U7639 (N_7639,N_7378,N_7296);
nand U7640 (N_7640,N_7090,N_7297);
nor U7641 (N_7641,N_7213,N_7316);
or U7642 (N_7642,N_7323,N_7089);
nand U7643 (N_7643,N_7039,N_7369);
nor U7644 (N_7644,N_7340,N_7304);
or U7645 (N_7645,N_7119,N_7189);
nand U7646 (N_7646,N_7127,N_7383);
or U7647 (N_7647,N_7235,N_7102);
nand U7648 (N_7648,N_7372,N_7096);
or U7649 (N_7649,N_7377,N_7209);
and U7650 (N_7650,N_7016,N_7278);
and U7651 (N_7651,N_7490,N_7468);
nand U7652 (N_7652,N_7032,N_7292);
nor U7653 (N_7653,N_7494,N_7245);
or U7654 (N_7654,N_7433,N_7185);
or U7655 (N_7655,N_7406,N_7220);
xnor U7656 (N_7656,N_7029,N_7295);
and U7657 (N_7657,N_7099,N_7423);
nor U7658 (N_7658,N_7267,N_7359);
and U7659 (N_7659,N_7318,N_7268);
nand U7660 (N_7660,N_7037,N_7042);
xnor U7661 (N_7661,N_7275,N_7463);
nor U7662 (N_7662,N_7034,N_7352);
nand U7663 (N_7663,N_7243,N_7379);
and U7664 (N_7664,N_7167,N_7118);
nand U7665 (N_7665,N_7471,N_7166);
or U7666 (N_7666,N_7375,N_7370);
nor U7667 (N_7667,N_7328,N_7434);
nor U7668 (N_7668,N_7290,N_7069);
nand U7669 (N_7669,N_7485,N_7054);
nor U7670 (N_7670,N_7487,N_7497);
nor U7671 (N_7671,N_7271,N_7363);
and U7672 (N_7672,N_7103,N_7035);
or U7673 (N_7673,N_7238,N_7184);
nor U7674 (N_7674,N_7057,N_7205);
nor U7675 (N_7675,N_7193,N_7313);
and U7676 (N_7676,N_7161,N_7019);
and U7677 (N_7677,N_7479,N_7417);
nand U7678 (N_7678,N_7394,N_7483);
and U7679 (N_7679,N_7128,N_7240);
nor U7680 (N_7680,N_7334,N_7015);
and U7681 (N_7681,N_7162,N_7214);
nand U7682 (N_7682,N_7391,N_7336);
or U7683 (N_7683,N_7076,N_7253);
nand U7684 (N_7684,N_7025,N_7484);
and U7685 (N_7685,N_7258,N_7215);
or U7686 (N_7686,N_7065,N_7233);
or U7687 (N_7687,N_7250,N_7456);
or U7688 (N_7688,N_7082,N_7158);
nand U7689 (N_7689,N_7138,N_7324);
or U7690 (N_7690,N_7115,N_7376);
nand U7691 (N_7691,N_7493,N_7344);
nand U7692 (N_7692,N_7219,N_7326);
nor U7693 (N_7693,N_7100,N_7171);
and U7694 (N_7694,N_7091,N_7386);
or U7695 (N_7695,N_7051,N_7449);
nor U7696 (N_7696,N_7399,N_7265);
and U7697 (N_7697,N_7178,N_7094);
and U7698 (N_7698,N_7059,N_7438);
or U7699 (N_7699,N_7188,N_7176);
xor U7700 (N_7700,N_7221,N_7368);
nand U7701 (N_7701,N_7001,N_7405);
or U7702 (N_7702,N_7058,N_7172);
and U7703 (N_7703,N_7137,N_7068);
or U7704 (N_7704,N_7203,N_7492);
or U7705 (N_7705,N_7114,N_7006);
nand U7706 (N_7706,N_7066,N_7358);
or U7707 (N_7707,N_7305,N_7498);
or U7708 (N_7708,N_7239,N_7183);
nor U7709 (N_7709,N_7155,N_7403);
and U7710 (N_7710,N_7351,N_7457);
or U7711 (N_7711,N_7014,N_7132);
or U7712 (N_7712,N_7286,N_7237);
nand U7713 (N_7713,N_7261,N_7382);
or U7714 (N_7714,N_7431,N_7374);
and U7715 (N_7715,N_7397,N_7308);
or U7716 (N_7716,N_7083,N_7177);
nand U7717 (N_7717,N_7005,N_7112);
and U7718 (N_7718,N_7228,N_7335);
and U7719 (N_7719,N_7175,N_7303);
nand U7720 (N_7720,N_7288,N_7055);
nor U7721 (N_7721,N_7047,N_7053);
nand U7722 (N_7722,N_7419,N_7211);
nand U7723 (N_7723,N_7300,N_7199);
xnor U7724 (N_7724,N_7476,N_7257);
nand U7725 (N_7725,N_7321,N_7022);
or U7726 (N_7726,N_7192,N_7196);
or U7727 (N_7727,N_7004,N_7134);
and U7728 (N_7728,N_7117,N_7105);
and U7729 (N_7729,N_7401,N_7122);
and U7730 (N_7730,N_7073,N_7249);
or U7731 (N_7731,N_7309,N_7355);
or U7732 (N_7732,N_7049,N_7000);
nor U7733 (N_7733,N_7124,N_7469);
nand U7734 (N_7734,N_7139,N_7439);
nand U7735 (N_7735,N_7179,N_7252);
nand U7736 (N_7736,N_7427,N_7151);
nand U7737 (N_7737,N_7354,N_7143);
or U7738 (N_7738,N_7079,N_7435);
nand U7739 (N_7739,N_7081,N_7106);
or U7740 (N_7740,N_7140,N_7388);
or U7741 (N_7741,N_7061,N_7481);
and U7742 (N_7742,N_7045,N_7071);
or U7743 (N_7743,N_7285,N_7218);
or U7744 (N_7744,N_7299,N_7152);
or U7745 (N_7745,N_7366,N_7052);
or U7746 (N_7746,N_7454,N_7407);
or U7747 (N_7747,N_7002,N_7251);
or U7748 (N_7748,N_7413,N_7197);
nand U7749 (N_7749,N_7210,N_7437);
nand U7750 (N_7750,N_7061,N_7220);
or U7751 (N_7751,N_7377,N_7491);
nor U7752 (N_7752,N_7368,N_7321);
and U7753 (N_7753,N_7385,N_7251);
and U7754 (N_7754,N_7316,N_7041);
nand U7755 (N_7755,N_7391,N_7247);
nor U7756 (N_7756,N_7406,N_7437);
nor U7757 (N_7757,N_7491,N_7461);
nor U7758 (N_7758,N_7112,N_7453);
nor U7759 (N_7759,N_7466,N_7298);
or U7760 (N_7760,N_7386,N_7432);
and U7761 (N_7761,N_7007,N_7327);
or U7762 (N_7762,N_7162,N_7172);
or U7763 (N_7763,N_7216,N_7347);
and U7764 (N_7764,N_7162,N_7313);
or U7765 (N_7765,N_7219,N_7091);
and U7766 (N_7766,N_7325,N_7164);
nor U7767 (N_7767,N_7150,N_7427);
and U7768 (N_7768,N_7384,N_7217);
or U7769 (N_7769,N_7382,N_7110);
nand U7770 (N_7770,N_7410,N_7291);
or U7771 (N_7771,N_7236,N_7005);
nor U7772 (N_7772,N_7327,N_7260);
nor U7773 (N_7773,N_7221,N_7330);
or U7774 (N_7774,N_7138,N_7080);
xor U7775 (N_7775,N_7056,N_7151);
and U7776 (N_7776,N_7232,N_7180);
nor U7777 (N_7777,N_7022,N_7054);
nor U7778 (N_7778,N_7327,N_7084);
or U7779 (N_7779,N_7274,N_7021);
nor U7780 (N_7780,N_7267,N_7490);
nor U7781 (N_7781,N_7224,N_7234);
nor U7782 (N_7782,N_7040,N_7139);
and U7783 (N_7783,N_7073,N_7454);
or U7784 (N_7784,N_7229,N_7315);
or U7785 (N_7785,N_7323,N_7087);
or U7786 (N_7786,N_7440,N_7477);
nand U7787 (N_7787,N_7119,N_7008);
nor U7788 (N_7788,N_7019,N_7222);
nand U7789 (N_7789,N_7013,N_7497);
and U7790 (N_7790,N_7477,N_7280);
and U7791 (N_7791,N_7433,N_7097);
nor U7792 (N_7792,N_7019,N_7441);
and U7793 (N_7793,N_7067,N_7405);
and U7794 (N_7794,N_7082,N_7180);
nor U7795 (N_7795,N_7135,N_7447);
and U7796 (N_7796,N_7195,N_7177);
and U7797 (N_7797,N_7278,N_7010);
xnor U7798 (N_7798,N_7252,N_7324);
and U7799 (N_7799,N_7450,N_7106);
nand U7800 (N_7800,N_7219,N_7211);
nand U7801 (N_7801,N_7120,N_7151);
or U7802 (N_7802,N_7296,N_7110);
or U7803 (N_7803,N_7463,N_7299);
nand U7804 (N_7804,N_7344,N_7158);
nand U7805 (N_7805,N_7156,N_7226);
or U7806 (N_7806,N_7488,N_7317);
nor U7807 (N_7807,N_7106,N_7188);
or U7808 (N_7808,N_7259,N_7319);
or U7809 (N_7809,N_7026,N_7047);
nor U7810 (N_7810,N_7363,N_7329);
nor U7811 (N_7811,N_7049,N_7251);
or U7812 (N_7812,N_7170,N_7184);
or U7813 (N_7813,N_7399,N_7197);
nor U7814 (N_7814,N_7325,N_7375);
nand U7815 (N_7815,N_7022,N_7368);
or U7816 (N_7816,N_7062,N_7047);
and U7817 (N_7817,N_7350,N_7471);
or U7818 (N_7818,N_7120,N_7047);
nor U7819 (N_7819,N_7289,N_7000);
or U7820 (N_7820,N_7293,N_7459);
and U7821 (N_7821,N_7458,N_7294);
xnor U7822 (N_7822,N_7159,N_7268);
nand U7823 (N_7823,N_7065,N_7104);
or U7824 (N_7824,N_7014,N_7188);
nand U7825 (N_7825,N_7147,N_7122);
and U7826 (N_7826,N_7433,N_7395);
xor U7827 (N_7827,N_7293,N_7174);
and U7828 (N_7828,N_7486,N_7222);
nor U7829 (N_7829,N_7234,N_7283);
nor U7830 (N_7830,N_7413,N_7354);
nand U7831 (N_7831,N_7346,N_7003);
nand U7832 (N_7832,N_7483,N_7200);
and U7833 (N_7833,N_7492,N_7056);
nand U7834 (N_7834,N_7112,N_7018);
or U7835 (N_7835,N_7486,N_7479);
or U7836 (N_7836,N_7230,N_7142);
or U7837 (N_7837,N_7400,N_7130);
nand U7838 (N_7838,N_7152,N_7212);
nand U7839 (N_7839,N_7040,N_7162);
nor U7840 (N_7840,N_7405,N_7386);
or U7841 (N_7841,N_7449,N_7473);
and U7842 (N_7842,N_7106,N_7343);
nand U7843 (N_7843,N_7065,N_7082);
nand U7844 (N_7844,N_7294,N_7386);
nand U7845 (N_7845,N_7095,N_7048);
or U7846 (N_7846,N_7127,N_7067);
or U7847 (N_7847,N_7189,N_7336);
nand U7848 (N_7848,N_7109,N_7266);
nor U7849 (N_7849,N_7071,N_7185);
and U7850 (N_7850,N_7293,N_7317);
nand U7851 (N_7851,N_7134,N_7042);
and U7852 (N_7852,N_7419,N_7227);
or U7853 (N_7853,N_7038,N_7478);
or U7854 (N_7854,N_7312,N_7320);
nand U7855 (N_7855,N_7115,N_7295);
nand U7856 (N_7856,N_7146,N_7058);
nand U7857 (N_7857,N_7360,N_7279);
nor U7858 (N_7858,N_7021,N_7065);
or U7859 (N_7859,N_7385,N_7110);
xnor U7860 (N_7860,N_7479,N_7017);
nand U7861 (N_7861,N_7138,N_7356);
nand U7862 (N_7862,N_7105,N_7290);
nor U7863 (N_7863,N_7390,N_7262);
nor U7864 (N_7864,N_7292,N_7359);
nand U7865 (N_7865,N_7193,N_7259);
and U7866 (N_7866,N_7448,N_7146);
nor U7867 (N_7867,N_7241,N_7091);
and U7868 (N_7868,N_7293,N_7246);
nor U7869 (N_7869,N_7186,N_7373);
and U7870 (N_7870,N_7048,N_7194);
or U7871 (N_7871,N_7453,N_7190);
or U7872 (N_7872,N_7116,N_7390);
nand U7873 (N_7873,N_7362,N_7287);
nand U7874 (N_7874,N_7320,N_7324);
nand U7875 (N_7875,N_7085,N_7015);
or U7876 (N_7876,N_7437,N_7045);
and U7877 (N_7877,N_7211,N_7465);
nand U7878 (N_7878,N_7223,N_7390);
nand U7879 (N_7879,N_7119,N_7491);
nor U7880 (N_7880,N_7398,N_7038);
nand U7881 (N_7881,N_7319,N_7209);
nor U7882 (N_7882,N_7429,N_7130);
nand U7883 (N_7883,N_7364,N_7453);
nor U7884 (N_7884,N_7468,N_7157);
nor U7885 (N_7885,N_7288,N_7394);
and U7886 (N_7886,N_7239,N_7103);
and U7887 (N_7887,N_7039,N_7180);
or U7888 (N_7888,N_7063,N_7072);
and U7889 (N_7889,N_7025,N_7153);
nand U7890 (N_7890,N_7317,N_7328);
or U7891 (N_7891,N_7072,N_7029);
nor U7892 (N_7892,N_7109,N_7070);
nand U7893 (N_7893,N_7429,N_7084);
nor U7894 (N_7894,N_7377,N_7087);
nor U7895 (N_7895,N_7405,N_7176);
or U7896 (N_7896,N_7206,N_7491);
nor U7897 (N_7897,N_7089,N_7263);
or U7898 (N_7898,N_7122,N_7470);
or U7899 (N_7899,N_7132,N_7228);
and U7900 (N_7900,N_7190,N_7373);
and U7901 (N_7901,N_7234,N_7295);
nand U7902 (N_7902,N_7169,N_7260);
nor U7903 (N_7903,N_7446,N_7064);
and U7904 (N_7904,N_7403,N_7216);
or U7905 (N_7905,N_7191,N_7031);
or U7906 (N_7906,N_7266,N_7308);
nand U7907 (N_7907,N_7246,N_7060);
and U7908 (N_7908,N_7430,N_7459);
nor U7909 (N_7909,N_7068,N_7346);
nand U7910 (N_7910,N_7360,N_7180);
and U7911 (N_7911,N_7408,N_7303);
nand U7912 (N_7912,N_7065,N_7152);
and U7913 (N_7913,N_7168,N_7071);
nand U7914 (N_7914,N_7014,N_7106);
and U7915 (N_7915,N_7489,N_7240);
nand U7916 (N_7916,N_7171,N_7369);
nor U7917 (N_7917,N_7205,N_7447);
nor U7918 (N_7918,N_7463,N_7101);
nor U7919 (N_7919,N_7376,N_7083);
nor U7920 (N_7920,N_7360,N_7417);
nor U7921 (N_7921,N_7129,N_7048);
and U7922 (N_7922,N_7335,N_7244);
and U7923 (N_7923,N_7345,N_7045);
nand U7924 (N_7924,N_7224,N_7040);
nand U7925 (N_7925,N_7233,N_7391);
and U7926 (N_7926,N_7132,N_7118);
nor U7927 (N_7927,N_7092,N_7088);
and U7928 (N_7928,N_7440,N_7456);
or U7929 (N_7929,N_7387,N_7177);
xor U7930 (N_7930,N_7084,N_7302);
nand U7931 (N_7931,N_7282,N_7384);
or U7932 (N_7932,N_7197,N_7480);
nand U7933 (N_7933,N_7385,N_7250);
nand U7934 (N_7934,N_7088,N_7037);
or U7935 (N_7935,N_7248,N_7158);
nor U7936 (N_7936,N_7222,N_7471);
nor U7937 (N_7937,N_7364,N_7490);
nand U7938 (N_7938,N_7039,N_7218);
and U7939 (N_7939,N_7189,N_7283);
or U7940 (N_7940,N_7424,N_7169);
or U7941 (N_7941,N_7389,N_7368);
or U7942 (N_7942,N_7310,N_7100);
and U7943 (N_7943,N_7239,N_7410);
nand U7944 (N_7944,N_7312,N_7232);
nor U7945 (N_7945,N_7243,N_7327);
nand U7946 (N_7946,N_7299,N_7062);
nand U7947 (N_7947,N_7378,N_7445);
and U7948 (N_7948,N_7218,N_7238);
nor U7949 (N_7949,N_7018,N_7431);
nor U7950 (N_7950,N_7365,N_7179);
and U7951 (N_7951,N_7132,N_7144);
nor U7952 (N_7952,N_7197,N_7086);
and U7953 (N_7953,N_7310,N_7269);
nand U7954 (N_7954,N_7151,N_7267);
nor U7955 (N_7955,N_7382,N_7468);
nor U7956 (N_7956,N_7046,N_7464);
nand U7957 (N_7957,N_7004,N_7371);
nor U7958 (N_7958,N_7425,N_7363);
or U7959 (N_7959,N_7012,N_7049);
nor U7960 (N_7960,N_7204,N_7279);
nor U7961 (N_7961,N_7394,N_7016);
nand U7962 (N_7962,N_7171,N_7104);
and U7963 (N_7963,N_7463,N_7288);
or U7964 (N_7964,N_7007,N_7347);
nand U7965 (N_7965,N_7082,N_7236);
nor U7966 (N_7966,N_7373,N_7316);
nand U7967 (N_7967,N_7438,N_7401);
or U7968 (N_7968,N_7384,N_7488);
nor U7969 (N_7969,N_7347,N_7070);
xor U7970 (N_7970,N_7329,N_7326);
nand U7971 (N_7971,N_7330,N_7431);
and U7972 (N_7972,N_7347,N_7030);
and U7973 (N_7973,N_7270,N_7243);
nand U7974 (N_7974,N_7342,N_7329);
or U7975 (N_7975,N_7358,N_7265);
nand U7976 (N_7976,N_7048,N_7207);
or U7977 (N_7977,N_7047,N_7098);
nand U7978 (N_7978,N_7127,N_7487);
nor U7979 (N_7979,N_7244,N_7410);
nand U7980 (N_7980,N_7474,N_7032);
nand U7981 (N_7981,N_7365,N_7382);
or U7982 (N_7982,N_7081,N_7102);
and U7983 (N_7983,N_7047,N_7317);
or U7984 (N_7984,N_7237,N_7085);
nand U7985 (N_7985,N_7391,N_7401);
nand U7986 (N_7986,N_7324,N_7474);
nand U7987 (N_7987,N_7195,N_7337);
and U7988 (N_7988,N_7357,N_7205);
and U7989 (N_7989,N_7247,N_7083);
and U7990 (N_7990,N_7022,N_7166);
or U7991 (N_7991,N_7357,N_7151);
nor U7992 (N_7992,N_7187,N_7467);
and U7993 (N_7993,N_7450,N_7387);
nor U7994 (N_7994,N_7456,N_7345);
or U7995 (N_7995,N_7002,N_7145);
and U7996 (N_7996,N_7038,N_7191);
and U7997 (N_7997,N_7293,N_7332);
nor U7998 (N_7998,N_7246,N_7344);
nor U7999 (N_7999,N_7101,N_7471);
nor U8000 (N_8000,N_7594,N_7537);
nor U8001 (N_8001,N_7986,N_7991);
nor U8002 (N_8002,N_7860,N_7612);
nor U8003 (N_8003,N_7942,N_7791);
nand U8004 (N_8004,N_7602,N_7982);
or U8005 (N_8005,N_7784,N_7956);
and U8006 (N_8006,N_7894,N_7897);
xnor U8007 (N_8007,N_7905,N_7579);
and U8008 (N_8008,N_7933,N_7752);
nor U8009 (N_8009,N_7911,N_7560);
nor U8010 (N_8010,N_7528,N_7676);
and U8011 (N_8011,N_7989,N_7827);
and U8012 (N_8012,N_7955,N_7657);
or U8013 (N_8013,N_7624,N_7976);
nand U8014 (N_8014,N_7793,N_7704);
and U8015 (N_8015,N_7570,N_7867);
or U8016 (N_8016,N_7936,N_7984);
nand U8017 (N_8017,N_7925,N_7899);
nor U8018 (N_8018,N_7798,N_7943);
nand U8019 (N_8019,N_7950,N_7682);
or U8020 (N_8020,N_7954,N_7902);
nor U8021 (N_8021,N_7981,N_7951);
nand U8022 (N_8022,N_7694,N_7907);
or U8023 (N_8023,N_7618,N_7926);
nor U8024 (N_8024,N_7736,N_7609);
nor U8025 (N_8025,N_7585,N_7776);
and U8026 (N_8026,N_7615,N_7815);
or U8027 (N_8027,N_7686,N_7965);
and U8028 (N_8028,N_7562,N_7828);
nand U8029 (N_8029,N_7917,N_7935);
or U8030 (N_8030,N_7941,N_7649);
nand U8031 (N_8031,N_7653,N_7509);
nand U8032 (N_8032,N_7814,N_7802);
or U8033 (N_8033,N_7808,N_7913);
and U8034 (N_8034,N_7763,N_7619);
and U8035 (N_8035,N_7788,N_7568);
nor U8036 (N_8036,N_7931,N_7874);
and U8037 (N_8037,N_7861,N_7616);
nor U8038 (N_8038,N_7540,N_7718);
nand U8039 (N_8039,N_7549,N_7645);
nand U8040 (N_8040,N_7683,N_7884);
nand U8041 (N_8041,N_7522,N_7635);
and U8042 (N_8042,N_7758,N_7781);
nor U8043 (N_8043,N_7970,N_7766);
or U8044 (N_8044,N_7893,N_7608);
and U8045 (N_8045,N_7888,N_7969);
and U8046 (N_8046,N_7906,N_7852);
or U8047 (N_8047,N_7957,N_7895);
nand U8048 (N_8048,N_7980,N_7789);
or U8049 (N_8049,N_7504,N_7526);
and U8050 (N_8050,N_7679,N_7782);
nor U8051 (N_8051,N_7963,N_7865);
nor U8052 (N_8052,N_7524,N_7885);
nand U8053 (N_8053,N_7673,N_7859);
and U8054 (N_8054,N_7632,N_7819);
or U8055 (N_8055,N_7846,N_7997);
and U8056 (N_8056,N_7580,N_7934);
and U8057 (N_8057,N_7614,N_7995);
or U8058 (N_8058,N_7896,N_7968);
nor U8059 (N_8059,N_7557,N_7832);
and U8060 (N_8060,N_7741,N_7703);
and U8061 (N_8061,N_7765,N_7503);
nor U8062 (N_8062,N_7574,N_7840);
nand U8063 (N_8063,N_7523,N_7998);
nand U8064 (N_8064,N_7947,N_7625);
and U8065 (N_8065,N_7967,N_7555);
and U8066 (N_8066,N_7719,N_7601);
nor U8067 (N_8067,N_7660,N_7650);
or U8068 (N_8068,N_7924,N_7889);
nor U8069 (N_8069,N_7949,N_7887);
nand U8070 (N_8070,N_7746,N_7790);
nand U8071 (N_8071,N_7975,N_7909);
nor U8072 (N_8072,N_7738,N_7774);
or U8073 (N_8073,N_7783,N_7643);
nor U8074 (N_8074,N_7856,N_7755);
nand U8075 (N_8075,N_7709,N_7651);
nor U8076 (N_8076,N_7550,N_7851);
or U8077 (N_8077,N_7868,N_7515);
nand U8078 (N_8078,N_7713,N_7903);
nor U8079 (N_8079,N_7593,N_7561);
or U8080 (N_8080,N_7661,N_7743);
nor U8081 (N_8081,N_7990,N_7834);
or U8082 (N_8082,N_7667,N_7506);
nor U8083 (N_8083,N_7655,N_7729);
or U8084 (N_8084,N_7646,N_7690);
and U8085 (N_8085,N_7833,N_7575);
and U8086 (N_8086,N_7564,N_7987);
nand U8087 (N_8087,N_7724,N_7711);
and U8088 (N_8088,N_7835,N_7881);
and U8089 (N_8089,N_7551,N_7598);
nor U8090 (N_8090,N_7730,N_7876);
or U8091 (N_8091,N_7707,N_7569);
nand U8092 (N_8092,N_7797,N_7767);
nand U8093 (N_8093,N_7688,N_7800);
and U8094 (N_8094,N_7578,N_7677);
or U8095 (N_8095,N_7761,N_7929);
and U8096 (N_8096,N_7536,N_7531);
nor U8097 (N_8097,N_7807,N_7611);
nand U8098 (N_8098,N_7825,N_7753);
nand U8099 (N_8099,N_7666,N_7697);
xnor U8100 (N_8100,N_7691,N_7778);
nand U8101 (N_8101,N_7589,N_7922);
xor U8102 (N_8102,N_7573,N_7723);
nor U8103 (N_8103,N_7698,N_7584);
nand U8104 (N_8104,N_7775,N_7757);
nand U8105 (N_8105,N_7717,N_7546);
nor U8106 (N_8106,N_7824,N_7544);
or U8107 (N_8107,N_7638,N_7809);
or U8108 (N_8108,N_7539,N_7764);
or U8109 (N_8109,N_7672,N_7883);
and U8110 (N_8110,N_7599,N_7974);
xor U8111 (N_8111,N_7621,N_7731);
and U8112 (N_8112,N_7822,N_7988);
or U8113 (N_8113,N_7559,N_7525);
and U8114 (N_8114,N_7699,N_7680);
and U8115 (N_8115,N_7558,N_7854);
or U8116 (N_8116,N_7886,N_7668);
nor U8117 (N_8117,N_7908,N_7554);
nor U8118 (N_8118,N_7748,N_7543);
nor U8119 (N_8119,N_7786,N_7813);
nor U8120 (N_8120,N_7507,N_7912);
and U8121 (N_8121,N_7607,N_7582);
and U8122 (N_8122,N_7879,N_7952);
or U8123 (N_8123,N_7932,N_7572);
nor U8124 (N_8124,N_7756,N_7750);
or U8125 (N_8125,N_7514,N_7818);
nor U8126 (N_8126,N_7739,N_7633);
or U8127 (N_8127,N_7725,N_7862);
nor U8128 (N_8128,N_7629,N_7500);
xor U8129 (N_8129,N_7830,N_7831);
nor U8130 (N_8130,N_7512,N_7805);
or U8131 (N_8131,N_7556,N_7610);
nor U8132 (N_8132,N_7678,N_7596);
nand U8133 (N_8133,N_7983,N_7882);
and U8134 (N_8134,N_7613,N_7692);
nor U8135 (N_8135,N_7921,N_7946);
nand U8136 (N_8136,N_7644,N_7606);
and U8137 (N_8137,N_7794,N_7826);
or U8138 (N_8138,N_7547,N_7674);
and U8139 (N_8139,N_7873,N_7772);
nor U8140 (N_8140,N_7938,N_7771);
nand U8141 (N_8141,N_7744,N_7518);
nor U8142 (N_8142,N_7617,N_7627);
nand U8143 (N_8143,N_7904,N_7631);
and U8144 (N_8144,N_7880,N_7519);
nor U8145 (N_8145,N_7622,N_7538);
nand U8146 (N_8146,N_7640,N_7960);
or U8147 (N_8147,N_7816,N_7745);
nor U8148 (N_8148,N_7542,N_7773);
nor U8149 (N_8149,N_7641,N_7945);
or U8150 (N_8150,N_7985,N_7715);
nand U8151 (N_8151,N_7636,N_7695);
or U8152 (N_8152,N_7710,N_7978);
nand U8153 (N_8153,N_7787,N_7654);
nand U8154 (N_8154,N_7693,N_7634);
nor U8155 (N_8155,N_7669,N_7749);
nand U8156 (N_8156,N_7735,N_7812);
nand U8157 (N_8157,N_7508,N_7623);
or U8158 (N_8158,N_7684,N_7892);
nand U8159 (N_8159,N_7505,N_7754);
nor U8160 (N_8160,N_7552,N_7855);
nor U8161 (N_8161,N_7737,N_7529);
nand U8162 (N_8162,N_7670,N_7548);
nor U8163 (N_8163,N_7993,N_7804);
nand U8164 (N_8164,N_7626,N_7864);
or U8165 (N_8165,N_7877,N_7541);
or U8166 (N_8166,N_7687,N_7647);
and U8167 (N_8167,N_7663,N_7747);
and U8168 (N_8168,N_7857,N_7517);
xnor U8169 (N_8169,N_7733,N_7762);
nor U8170 (N_8170,N_7849,N_7656);
and U8171 (N_8171,N_7915,N_7702);
nand U8172 (N_8172,N_7532,N_7930);
nor U8173 (N_8173,N_7844,N_7590);
nand U8174 (N_8174,N_7586,N_7811);
or U8175 (N_8175,N_7628,N_7891);
nand U8176 (N_8176,N_7603,N_7553);
nand U8177 (N_8177,N_7652,N_7977);
and U8178 (N_8178,N_7959,N_7581);
and U8179 (N_8179,N_7900,N_7510);
nor U8180 (N_8180,N_7658,N_7962);
or U8181 (N_8181,N_7576,N_7705);
and U8182 (N_8182,N_7914,N_7973);
nor U8183 (N_8183,N_7801,N_7721);
nand U8184 (N_8184,N_7759,N_7696);
and U8185 (N_8185,N_7591,N_7820);
nand U8186 (N_8186,N_7732,N_7910);
nor U8187 (N_8187,N_7871,N_7769);
nand U8188 (N_8188,N_7742,N_7853);
or U8189 (N_8189,N_7777,N_7639);
and U8190 (N_8190,N_7642,N_7839);
and U8191 (N_8191,N_7996,N_7516);
nor U8192 (N_8192,N_7878,N_7999);
nand U8193 (N_8193,N_7821,N_7563);
or U8194 (N_8194,N_7533,N_7520);
nor U8195 (N_8195,N_7961,N_7706);
and U8196 (N_8196,N_7577,N_7940);
nand U8197 (N_8197,N_7600,N_7841);
nand U8198 (N_8198,N_7664,N_7845);
nor U8199 (N_8199,N_7944,N_7928);
nor U8200 (N_8200,N_7770,N_7720);
and U8201 (N_8201,N_7513,N_7535);
nor U8202 (N_8202,N_7620,N_7566);
and U8203 (N_8203,N_7890,N_7714);
nor U8204 (N_8204,N_7502,N_7901);
or U8205 (N_8205,N_7823,N_7665);
and U8206 (N_8206,N_7817,N_7842);
nor U8207 (N_8207,N_7521,N_7779);
and U8208 (N_8208,N_7918,N_7681);
nor U8209 (N_8209,N_7796,N_7799);
or U8210 (N_8210,N_7994,N_7964);
nand U8211 (N_8211,N_7592,N_7870);
and U8212 (N_8212,N_7875,N_7948);
nand U8213 (N_8213,N_7728,N_7604);
nand U8214 (N_8214,N_7630,N_7760);
nand U8215 (N_8215,N_7869,N_7836);
and U8216 (N_8216,N_7527,N_7768);
and U8217 (N_8217,N_7722,N_7939);
and U8218 (N_8218,N_7712,N_7829);
or U8219 (N_8219,N_7701,N_7838);
nor U8220 (N_8220,N_7685,N_7992);
nand U8221 (N_8221,N_7937,N_7872);
nor U8222 (N_8222,N_7511,N_7803);
and U8223 (N_8223,N_7806,N_7726);
and U8224 (N_8224,N_7605,N_7565);
nand U8225 (N_8225,N_7916,N_7659);
nor U8226 (N_8226,N_7567,N_7780);
nand U8227 (N_8227,N_7966,N_7953);
or U8228 (N_8228,N_7671,N_7587);
nor U8229 (N_8229,N_7595,N_7530);
nor U8230 (N_8230,N_7927,N_7648);
or U8231 (N_8231,N_7662,N_7923);
or U8232 (N_8232,N_7708,N_7534);
nand U8233 (N_8233,N_7843,N_7979);
or U8234 (N_8234,N_7785,N_7848);
nand U8235 (N_8235,N_7597,N_7740);
and U8236 (N_8236,N_7751,N_7689);
or U8237 (N_8237,N_7583,N_7971);
or U8238 (N_8238,N_7863,N_7716);
and U8239 (N_8239,N_7501,N_7920);
nor U8240 (N_8240,N_7588,N_7858);
and U8241 (N_8241,N_7898,N_7727);
or U8242 (N_8242,N_7571,N_7810);
nor U8243 (N_8243,N_7972,N_7675);
or U8244 (N_8244,N_7792,N_7795);
nand U8245 (N_8245,N_7637,N_7847);
nand U8246 (N_8246,N_7545,N_7866);
nor U8247 (N_8247,N_7837,N_7958);
nand U8248 (N_8248,N_7734,N_7850);
nor U8249 (N_8249,N_7919,N_7700);
nor U8250 (N_8250,N_7987,N_7787);
nor U8251 (N_8251,N_7782,N_7821);
or U8252 (N_8252,N_7636,N_7820);
and U8253 (N_8253,N_7587,N_7908);
nand U8254 (N_8254,N_7627,N_7821);
xnor U8255 (N_8255,N_7936,N_7694);
and U8256 (N_8256,N_7679,N_7952);
and U8257 (N_8257,N_7983,N_7538);
nor U8258 (N_8258,N_7909,N_7856);
nor U8259 (N_8259,N_7926,N_7838);
and U8260 (N_8260,N_7969,N_7915);
and U8261 (N_8261,N_7941,N_7854);
nand U8262 (N_8262,N_7636,N_7999);
nand U8263 (N_8263,N_7573,N_7707);
xor U8264 (N_8264,N_7548,N_7584);
and U8265 (N_8265,N_7849,N_7811);
or U8266 (N_8266,N_7991,N_7931);
nand U8267 (N_8267,N_7512,N_7657);
or U8268 (N_8268,N_7541,N_7578);
nand U8269 (N_8269,N_7872,N_7702);
nor U8270 (N_8270,N_7801,N_7832);
nand U8271 (N_8271,N_7758,N_7545);
or U8272 (N_8272,N_7551,N_7933);
and U8273 (N_8273,N_7733,N_7847);
or U8274 (N_8274,N_7717,N_7803);
nor U8275 (N_8275,N_7657,N_7533);
nand U8276 (N_8276,N_7740,N_7807);
or U8277 (N_8277,N_7576,N_7800);
nor U8278 (N_8278,N_7933,N_7808);
nand U8279 (N_8279,N_7501,N_7993);
nand U8280 (N_8280,N_7693,N_7832);
nand U8281 (N_8281,N_7668,N_7866);
or U8282 (N_8282,N_7674,N_7819);
or U8283 (N_8283,N_7959,N_7998);
and U8284 (N_8284,N_7637,N_7813);
nand U8285 (N_8285,N_7528,N_7745);
nand U8286 (N_8286,N_7866,N_7585);
nor U8287 (N_8287,N_7893,N_7706);
nor U8288 (N_8288,N_7541,N_7545);
nor U8289 (N_8289,N_7541,N_7904);
nor U8290 (N_8290,N_7724,N_7996);
and U8291 (N_8291,N_7564,N_7572);
or U8292 (N_8292,N_7952,N_7829);
or U8293 (N_8293,N_7674,N_7972);
nand U8294 (N_8294,N_7971,N_7951);
nand U8295 (N_8295,N_7782,N_7520);
and U8296 (N_8296,N_7934,N_7571);
and U8297 (N_8297,N_7891,N_7842);
nand U8298 (N_8298,N_7883,N_7573);
nand U8299 (N_8299,N_7717,N_7831);
and U8300 (N_8300,N_7989,N_7538);
nand U8301 (N_8301,N_7572,N_7997);
and U8302 (N_8302,N_7678,N_7829);
nand U8303 (N_8303,N_7516,N_7985);
and U8304 (N_8304,N_7831,N_7918);
nor U8305 (N_8305,N_7924,N_7545);
nand U8306 (N_8306,N_7790,N_7941);
or U8307 (N_8307,N_7797,N_7761);
and U8308 (N_8308,N_7847,N_7584);
nor U8309 (N_8309,N_7938,N_7595);
or U8310 (N_8310,N_7963,N_7851);
nand U8311 (N_8311,N_7764,N_7594);
or U8312 (N_8312,N_7980,N_7563);
and U8313 (N_8313,N_7955,N_7872);
and U8314 (N_8314,N_7794,N_7815);
or U8315 (N_8315,N_7957,N_7503);
nand U8316 (N_8316,N_7909,N_7543);
or U8317 (N_8317,N_7674,N_7977);
nor U8318 (N_8318,N_7916,N_7580);
or U8319 (N_8319,N_7726,N_7708);
nor U8320 (N_8320,N_7574,N_7650);
nand U8321 (N_8321,N_7626,N_7799);
nor U8322 (N_8322,N_7863,N_7704);
nor U8323 (N_8323,N_7967,N_7757);
nor U8324 (N_8324,N_7958,N_7799);
and U8325 (N_8325,N_7501,N_7505);
and U8326 (N_8326,N_7985,N_7867);
nand U8327 (N_8327,N_7924,N_7900);
nor U8328 (N_8328,N_7847,N_7857);
or U8329 (N_8329,N_7946,N_7986);
nand U8330 (N_8330,N_7720,N_7547);
or U8331 (N_8331,N_7613,N_7917);
or U8332 (N_8332,N_7702,N_7729);
or U8333 (N_8333,N_7560,N_7978);
nor U8334 (N_8334,N_7902,N_7573);
nor U8335 (N_8335,N_7742,N_7527);
nor U8336 (N_8336,N_7904,N_7528);
nand U8337 (N_8337,N_7512,N_7872);
nor U8338 (N_8338,N_7586,N_7536);
and U8339 (N_8339,N_7879,N_7741);
nor U8340 (N_8340,N_7774,N_7755);
and U8341 (N_8341,N_7920,N_7889);
nor U8342 (N_8342,N_7870,N_7576);
or U8343 (N_8343,N_7902,N_7557);
or U8344 (N_8344,N_7659,N_7979);
xor U8345 (N_8345,N_7607,N_7619);
or U8346 (N_8346,N_7518,N_7680);
and U8347 (N_8347,N_7725,N_7826);
and U8348 (N_8348,N_7805,N_7849);
or U8349 (N_8349,N_7722,N_7772);
or U8350 (N_8350,N_7714,N_7949);
nor U8351 (N_8351,N_7969,N_7642);
and U8352 (N_8352,N_7653,N_7799);
or U8353 (N_8353,N_7613,N_7652);
nand U8354 (N_8354,N_7613,N_7732);
nor U8355 (N_8355,N_7586,N_7527);
and U8356 (N_8356,N_7605,N_7667);
nand U8357 (N_8357,N_7600,N_7911);
or U8358 (N_8358,N_7921,N_7780);
nor U8359 (N_8359,N_7856,N_7940);
nor U8360 (N_8360,N_7540,N_7822);
or U8361 (N_8361,N_7943,N_7975);
or U8362 (N_8362,N_7563,N_7978);
nor U8363 (N_8363,N_7527,N_7650);
nand U8364 (N_8364,N_7729,N_7653);
and U8365 (N_8365,N_7560,N_7631);
nand U8366 (N_8366,N_7625,N_7846);
or U8367 (N_8367,N_7970,N_7648);
or U8368 (N_8368,N_7569,N_7819);
and U8369 (N_8369,N_7640,N_7681);
or U8370 (N_8370,N_7812,N_7628);
nor U8371 (N_8371,N_7713,N_7804);
nor U8372 (N_8372,N_7871,N_7642);
nand U8373 (N_8373,N_7974,N_7638);
or U8374 (N_8374,N_7600,N_7843);
nand U8375 (N_8375,N_7998,N_7688);
and U8376 (N_8376,N_7942,N_7978);
nand U8377 (N_8377,N_7559,N_7596);
nand U8378 (N_8378,N_7630,N_7889);
and U8379 (N_8379,N_7906,N_7602);
or U8380 (N_8380,N_7764,N_7736);
or U8381 (N_8381,N_7595,N_7591);
nor U8382 (N_8382,N_7891,N_7638);
nor U8383 (N_8383,N_7923,N_7600);
or U8384 (N_8384,N_7657,N_7778);
and U8385 (N_8385,N_7813,N_7743);
nor U8386 (N_8386,N_7689,N_7548);
and U8387 (N_8387,N_7919,N_7830);
nor U8388 (N_8388,N_7711,N_7844);
and U8389 (N_8389,N_7639,N_7515);
nand U8390 (N_8390,N_7648,N_7930);
nor U8391 (N_8391,N_7611,N_7625);
nor U8392 (N_8392,N_7901,N_7951);
and U8393 (N_8393,N_7812,N_7571);
nand U8394 (N_8394,N_7667,N_7651);
nand U8395 (N_8395,N_7693,N_7921);
nor U8396 (N_8396,N_7707,N_7697);
xor U8397 (N_8397,N_7670,N_7697);
xnor U8398 (N_8398,N_7755,N_7588);
nand U8399 (N_8399,N_7563,N_7718);
nand U8400 (N_8400,N_7617,N_7986);
nand U8401 (N_8401,N_7621,N_7975);
nand U8402 (N_8402,N_7643,N_7745);
nand U8403 (N_8403,N_7607,N_7777);
nor U8404 (N_8404,N_7892,N_7659);
nor U8405 (N_8405,N_7574,N_7636);
nor U8406 (N_8406,N_7931,N_7610);
nand U8407 (N_8407,N_7948,N_7720);
nor U8408 (N_8408,N_7801,N_7885);
nand U8409 (N_8409,N_7988,N_7638);
or U8410 (N_8410,N_7553,N_7881);
nand U8411 (N_8411,N_7746,N_7926);
nand U8412 (N_8412,N_7754,N_7920);
or U8413 (N_8413,N_7726,N_7609);
and U8414 (N_8414,N_7821,N_7800);
nor U8415 (N_8415,N_7513,N_7545);
or U8416 (N_8416,N_7954,N_7509);
and U8417 (N_8417,N_7984,N_7983);
and U8418 (N_8418,N_7973,N_7995);
nand U8419 (N_8419,N_7700,N_7927);
or U8420 (N_8420,N_7856,N_7853);
nand U8421 (N_8421,N_7572,N_7603);
and U8422 (N_8422,N_7634,N_7864);
xor U8423 (N_8423,N_7826,N_7610);
and U8424 (N_8424,N_7672,N_7634);
and U8425 (N_8425,N_7867,N_7808);
and U8426 (N_8426,N_7568,N_7986);
or U8427 (N_8427,N_7883,N_7732);
nand U8428 (N_8428,N_7627,N_7584);
and U8429 (N_8429,N_7609,N_7747);
and U8430 (N_8430,N_7679,N_7937);
nand U8431 (N_8431,N_7698,N_7856);
or U8432 (N_8432,N_7511,N_7937);
and U8433 (N_8433,N_7912,N_7883);
or U8434 (N_8434,N_7890,N_7863);
nand U8435 (N_8435,N_7635,N_7924);
xnor U8436 (N_8436,N_7707,N_7931);
and U8437 (N_8437,N_7526,N_7688);
nand U8438 (N_8438,N_7542,N_7604);
or U8439 (N_8439,N_7904,N_7572);
and U8440 (N_8440,N_7613,N_7796);
or U8441 (N_8441,N_7659,N_7913);
nand U8442 (N_8442,N_7659,N_7599);
nand U8443 (N_8443,N_7717,N_7820);
nor U8444 (N_8444,N_7722,N_7633);
nand U8445 (N_8445,N_7954,N_7815);
nand U8446 (N_8446,N_7814,N_7720);
or U8447 (N_8447,N_7543,N_7873);
nand U8448 (N_8448,N_7664,N_7518);
nand U8449 (N_8449,N_7674,N_7550);
and U8450 (N_8450,N_7745,N_7859);
and U8451 (N_8451,N_7719,N_7553);
or U8452 (N_8452,N_7831,N_7863);
nor U8453 (N_8453,N_7808,N_7886);
or U8454 (N_8454,N_7728,N_7944);
nand U8455 (N_8455,N_7949,N_7807);
nand U8456 (N_8456,N_7632,N_7830);
nor U8457 (N_8457,N_7627,N_7985);
nand U8458 (N_8458,N_7878,N_7742);
or U8459 (N_8459,N_7772,N_7611);
and U8460 (N_8460,N_7760,N_7632);
or U8461 (N_8461,N_7575,N_7899);
nor U8462 (N_8462,N_7749,N_7808);
nand U8463 (N_8463,N_7623,N_7634);
xnor U8464 (N_8464,N_7536,N_7780);
nand U8465 (N_8465,N_7502,N_7894);
and U8466 (N_8466,N_7805,N_7872);
and U8467 (N_8467,N_7915,N_7764);
nor U8468 (N_8468,N_7932,N_7648);
and U8469 (N_8469,N_7553,N_7676);
or U8470 (N_8470,N_7753,N_7834);
and U8471 (N_8471,N_7555,N_7806);
nand U8472 (N_8472,N_7900,N_7766);
nor U8473 (N_8473,N_7693,N_7829);
nand U8474 (N_8474,N_7818,N_7978);
or U8475 (N_8475,N_7884,N_7689);
nand U8476 (N_8476,N_7742,N_7557);
nand U8477 (N_8477,N_7854,N_7664);
or U8478 (N_8478,N_7870,N_7581);
nand U8479 (N_8479,N_7944,N_7830);
or U8480 (N_8480,N_7778,N_7663);
nand U8481 (N_8481,N_7987,N_7620);
nor U8482 (N_8482,N_7854,N_7580);
xor U8483 (N_8483,N_7763,N_7899);
nand U8484 (N_8484,N_7863,N_7687);
nor U8485 (N_8485,N_7681,N_7532);
nand U8486 (N_8486,N_7582,N_7748);
and U8487 (N_8487,N_7544,N_7771);
nand U8488 (N_8488,N_7959,N_7797);
and U8489 (N_8489,N_7862,N_7745);
or U8490 (N_8490,N_7531,N_7882);
and U8491 (N_8491,N_7724,N_7566);
nor U8492 (N_8492,N_7661,N_7631);
and U8493 (N_8493,N_7522,N_7747);
and U8494 (N_8494,N_7692,N_7625);
and U8495 (N_8495,N_7515,N_7793);
xnor U8496 (N_8496,N_7870,N_7674);
nor U8497 (N_8497,N_7714,N_7602);
nand U8498 (N_8498,N_7638,N_7901);
nand U8499 (N_8499,N_7714,N_7686);
and U8500 (N_8500,N_8058,N_8288);
nor U8501 (N_8501,N_8458,N_8066);
or U8502 (N_8502,N_8110,N_8206);
nand U8503 (N_8503,N_8452,N_8235);
nand U8504 (N_8504,N_8075,N_8013);
or U8505 (N_8505,N_8213,N_8364);
and U8506 (N_8506,N_8086,N_8064);
nor U8507 (N_8507,N_8355,N_8105);
or U8508 (N_8508,N_8014,N_8442);
and U8509 (N_8509,N_8264,N_8087);
and U8510 (N_8510,N_8112,N_8296);
or U8511 (N_8511,N_8084,N_8470);
or U8512 (N_8512,N_8226,N_8377);
or U8513 (N_8513,N_8358,N_8212);
or U8514 (N_8514,N_8186,N_8218);
and U8515 (N_8515,N_8029,N_8284);
or U8516 (N_8516,N_8426,N_8291);
or U8517 (N_8517,N_8404,N_8137);
xnor U8518 (N_8518,N_8131,N_8003);
xor U8519 (N_8519,N_8390,N_8190);
nor U8520 (N_8520,N_8198,N_8265);
or U8521 (N_8521,N_8300,N_8170);
or U8522 (N_8522,N_8059,N_8255);
xnor U8523 (N_8523,N_8046,N_8368);
nand U8524 (N_8524,N_8103,N_8178);
nor U8525 (N_8525,N_8323,N_8278);
and U8526 (N_8526,N_8373,N_8040);
nand U8527 (N_8527,N_8388,N_8182);
and U8528 (N_8528,N_8465,N_8466);
xor U8529 (N_8529,N_8293,N_8257);
nand U8530 (N_8530,N_8381,N_8322);
xnor U8531 (N_8531,N_8357,N_8267);
nor U8532 (N_8532,N_8242,N_8495);
and U8533 (N_8533,N_8340,N_8229);
nand U8534 (N_8534,N_8021,N_8150);
nor U8535 (N_8535,N_8455,N_8376);
nand U8536 (N_8536,N_8023,N_8155);
nor U8537 (N_8537,N_8425,N_8015);
and U8538 (N_8538,N_8001,N_8124);
nand U8539 (N_8539,N_8398,N_8175);
nand U8540 (N_8540,N_8069,N_8313);
nor U8541 (N_8541,N_8488,N_8083);
and U8542 (N_8542,N_8473,N_8494);
and U8543 (N_8543,N_8185,N_8018);
or U8544 (N_8544,N_8151,N_8268);
xnor U8545 (N_8545,N_8076,N_8335);
or U8546 (N_8546,N_8414,N_8026);
and U8547 (N_8547,N_8400,N_8041);
or U8548 (N_8548,N_8408,N_8431);
nand U8549 (N_8549,N_8342,N_8403);
nor U8550 (N_8550,N_8104,N_8312);
nor U8551 (N_8551,N_8308,N_8231);
nand U8552 (N_8552,N_8480,N_8096);
nor U8553 (N_8553,N_8223,N_8391);
and U8554 (N_8554,N_8347,N_8101);
and U8555 (N_8555,N_8251,N_8315);
nor U8556 (N_8556,N_8162,N_8147);
nor U8557 (N_8557,N_8445,N_8311);
nand U8558 (N_8558,N_8149,N_8166);
and U8559 (N_8559,N_8139,N_8049);
nand U8560 (N_8560,N_8309,N_8177);
nor U8561 (N_8561,N_8443,N_8446);
and U8562 (N_8562,N_8286,N_8220);
nor U8563 (N_8563,N_8197,N_8191);
and U8564 (N_8564,N_8294,N_8369);
or U8565 (N_8565,N_8419,N_8019);
or U8566 (N_8566,N_8352,N_8448);
or U8567 (N_8567,N_8454,N_8290);
nor U8568 (N_8568,N_8052,N_8384);
nand U8569 (N_8569,N_8138,N_8184);
or U8570 (N_8570,N_8215,N_8359);
nand U8571 (N_8571,N_8094,N_8028);
nand U8572 (N_8572,N_8476,N_8095);
nand U8573 (N_8573,N_8393,N_8421);
or U8574 (N_8574,N_8120,N_8459);
and U8575 (N_8575,N_8478,N_8319);
and U8576 (N_8576,N_8496,N_8475);
or U8577 (N_8577,N_8148,N_8256);
xor U8578 (N_8578,N_8092,N_8158);
nor U8579 (N_8579,N_8196,N_8063);
or U8580 (N_8580,N_8118,N_8362);
nor U8581 (N_8581,N_8238,N_8349);
or U8582 (N_8582,N_8067,N_8244);
nor U8583 (N_8583,N_8330,N_8202);
nor U8584 (N_8584,N_8438,N_8392);
nand U8585 (N_8585,N_8317,N_8119);
nand U8586 (N_8586,N_8114,N_8132);
and U8587 (N_8587,N_8042,N_8217);
and U8588 (N_8588,N_8201,N_8463);
and U8589 (N_8589,N_8062,N_8004);
nand U8590 (N_8590,N_8462,N_8387);
and U8591 (N_8591,N_8022,N_8273);
nand U8592 (N_8592,N_8295,N_8474);
nor U8593 (N_8593,N_8161,N_8224);
and U8594 (N_8594,N_8232,N_8129);
nor U8595 (N_8595,N_8292,N_8000);
and U8596 (N_8596,N_8337,N_8417);
nand U8597 (N_8597,N_8033,N_8090);
nor U8598 (N_8598,N_8050,N_8136);
and U8599 (N_8599,N_8266,N_8047);
and U8600 (N_8600,N_8385,N_8126);
and U8601 (N_8601,N_8035,N_8254);
and U8602 (N_8602,N_8310,N_8303);
or U8603 (N_8603,N_8239,N_8199);
and U8604 (N_8604,N_8024,N_8469);
nor U8605 (N_8605,N_8179,N_8370);
or U8606 (N_8606,N_8361,N_8109);
nand U8607 (N_8607,N_8253,N_8439);
and U8608 (N_8608,N_8209,N_8356);
and U8609 (N_8609,N_8188,N_8360);
and U8610 (N_8610,N_8055,N_8276);
nor U8611 (N_8611,N_8449,N_8241);
nand U8612 (N_8612,N_8240,N_8012);
nand U8613 (N_8613,N_8499,N_8383);
or U8614 (N_8614,N_8485,N_8214);
xor U8615 (N_8615,N_8133,N_8314);
nor U8616 (N_8616,N_8187,N_8219);
and U8617 (N_8617,N_8236,N_8374);
nor U8618 (N_8618,N_8247,N_8367);
and U8619 (N_8619,N_8327,N_8125);
nand U8620 (N_8620,N_8416,N_8172);
or U8621 (N_8621,N_8225,N_8423);
and U8622 (N_8622,N_8407,N_8169);
or U8623 (N_8623,N_8420,N_8221);
or U8624 (N_8624,N_8031,N_8252);
nor U8625 (N_8625,N_8456,N_8363);
xnor U8626 (N_8626,N_8085,N_8233);
nand U8627 (N_8627,N_8350,N_8111);
and U8628 (N_8628,N_8117,N_8057);
nor U8629 (N_8629,N_8486,N_8039);
nor U8630 (N_8630,N_8077,N_8230);
and U8631 (N_8631,N_8068,N_8316);
or U8632 (N_8632,N_8332,N_8193);
and U8633 (N_8633,N_8245,N_8298);
or U8634 (N_8634,N_8301,N_8168);
nand U8635 (N_8635,N_8305,N_8098);
nand U8636 (N_8636,N_8453,N_8280);
nor U8637 (N_8637,N_8140,N_8428);
and U8638 (N_8638,N_8418,N_8008);
and U8639 (N_8639,N_8237,N_8246);
nand U8640 (N_8640,N_8167,N_8378);
or U8641 (N_8641,N_8045,N_8195);
nor U8642 (N_8642,N_8405,N_8152);
or U8643 (N_8643,N_8402,N_8460);
or U8644 (N_8644,N_8468,N_8281);
or U8645 (N_8645,N_8461,N_8306);
or U8646 (N_8646,N_8344,N_8183);
and U8647 (N_8647,N_8157,N_8341);
nor U8648 (N_8648,N_8056,N_8399);
or U8649 (N_8649,N_8135,N_8054);
nand U8650 (N_8650,N_8401,N_8078);
and U8651 (N_8651,N_8032,N_8271);
and U8652 (N_8652,N_8471,N_8146);
nor U8653 (N_8653,N_8415,N_8020);
nor U8654 (N_8654,N_8434,N_8329);
nand U8655 (N_8655,N_8429,N_8048);
and U8656 (N_8656,N_8005,N_8249);
or U8657 (N_8657,N_8444,N_8339);
and U8658 (N_8658,N_8487,N_8044);
nor U8659 (N_8659,N_8006,N_8102);
and U8660 (N_8660,N_8153,N_8437);
nand U8661 (N_8661,N_8261,N_8483);
nor U8662 (N_8662,N_8441,N_8440);
and U8663 (N_8663,N_8272,N_8060);
nand U8664 (N_8664,N_8051,N_8481);
nand U8665 (N_8665,N_8071,N_8053);
and U8666 (N_8666,N_8011,N_8491);
xnor U8667 (N_8667,N_8497,N_8176);
nor U8668 (N_8668,N_8093,N_8289);
and U8669 (N_8669,N_8269,N_8204);
or U8670 (N_8670,N_8328,N_8287);
nor U8671 (N_8671,N_8208,N_8173);
and U8672 (N_8672,N_8477,N_8397);
nor U8673 (N_8673,N_8163,N_8036);
or U8674 (N_8674,N_8025,N_8380);
nand U8675 (N_8675,N_8108,N_8088);
nand U8676 (N_8676,N_8192,N_8283);
nand U8677 (N_8677,N_8189,N_8203);
xnor U8678 (N_8678,N_8436,N_8320);
nand U8679 (N_8679,N_8234,N_8274);
nand U8680 (N_8680,N_8143,N_8160);
or U8681 (N_8681,N_8258,N_8411);
xnor U8682 (N_8682,N_8259,N_8227);
and U8683 (N_8683,N_8489,N_8074);
or U8684 (N_8684,N_8115,N_8422);
nor U8685 (N_8685,N_8243,N_8263);
and U8686 (N_8686,N_8345,N_8141);
or U8687 (N_8687,N_8070,N_8113);
nand U8688 (N_8688,N_8336,N_8299);
nand U8689 (N_8689,N_8326,N_8061);
nand U8690 (N_8690,N_8386,N_8130);
or U8691 (N_8691,N_8285,N_8447);
or U8692 (N_8692,N_8002,N_8081);
nor U8693 (N_8693,N_8318,N_8211);
and U8694 (N_8694,N_8282,N_8275);
and U8695 (N_8695,N_8409,N_8038);
and U8696 (N_8696,N_8073,N_8279);
and U8697 (N_8697,N_8207,N_8079);
nand U8698 (N_8698,N_8457,N_8016);
nand U8699 (N_8699,N_8262,N_8451);
nor U8700 (N_8700,N_8099,N_8116);
xor U8701 (N_8701,N_8097,N_8302);
nor U8702 (N_8702,N_8174,N_8371);
nand U8703 (N_8703,N_8493,N_8009);
nand U8704 (N_8704,N_8424,N_8121);
nor U8705 (N_8705,N_8127,N_8366);
nand U8706 (N_8706,N_8171,N_8412);
and U8707 (N_8707,N_8194,N_8100);
nor U8708 (N_8708,N_8333,N_8389);
xnor U8709 (N_8709,N_8228,N_8037);
or U8710 (N_8710,N_8427,N_8348);
and U8711 (N_8711,N_8030,N_8382);
and U8712 (N_8712,N_8122,N_8435);
nor U8713 (N_8713,N_8395,N_8181);
and U8714 (N_8714,N_8354,N_8484);
nor U8715 (N_8715,N_8107,N_8200);
nand U8716 (N_8716,N_8396,N_8433);
and U8717 (N_8717,N_8479,N_8346);
nand U8718 (N_8718,N_8091,N_8123);
and U8719 (N_8719,N_8159,N_8394);
nand U8720 (N_8720,N_8321,N_8334);
nor U8721 (N_8721,N_8106,N_8375);
nor U8722 (N_8722,N_8164,N_8248);
or U8723 (N_8723,N_8180,N_8205);
nand U8724 (N_8724,N_8017,N_8270);
nor U8725 (N_8725,N_8379,N_8351);
and U8726 (N_8726,N_8080,N_8216);
or U8727 (N_8727,N_8467,N_8007);
and U8728 (N_8728,N_8010,N_8210);
and U8729 (N_8729,N_8490,N_8410);
nand U8730 (N_8730,N_8128,N_8406);
and U8731 (N_8731,N_8277,N_8082);
nand U8732 (N_8732,N_8492,N_8250);
nor U8733 (N_8733,N_8304,N_8089);
and U8734 (N_8734,N_8027,N_8144);
nand U8735 (N_8735,N_8482,N_8498);
and U8736 (N_8736,N_8365,N_8156);
nand U8737 (N_8737,N_8043,N_8450);
or U8738 (N_8738,N_8432,N_8072);
or U8739 (N_8739,N_8297,N_8413);
nor U8740 (N_8740,N_8260,N_8154);
or U8741 (N_8741,N_8222,N_8307);
or U8742 (N_8742,N_8165,N_8338);
and U8743 (N_8743,N_8134,N_8464);
or U8744 (N_8744,N_8430,N_8472);
nand U8745 (N_8745,N_8065,N_8353);
or U8746 (N_8746,N_8034,N_8325);
xnor U8747 (N_8747,N_8343,N_8372);
and U8748 (N_8748,N_8324,N_8145);
and U8749 (N_8749,N_8142,N_8331);
nand U8750 (N_8750,N_8416,N_8478);
or U8751 (N_8751,N_8014,N_8131);
and U8752 (N_8752,N_8001,N_8320);
nor U8753 (N_8753,N_8239,N_8392);
nor U8754 (N_8754,N_8455,N_8071);
or U8755 (N_8755,N_8008,N_8269);
or U8756 (N_8756,N_8169,N_8276);
and U8757 (N_8757,N_8236,N_8036);
nor U8758 (N_8758,N_8018,N_8477);
nor U8759 (N_8759,N_8022,N_8177);
nor U8760 (N_8760,N_8491,N_8100);
and U8761 (N_8761,N_8207,N_8190);
or U8762 (N_8762,N_8067,N_8116);
or U8763 (N_8763,N_8066,N_8492);
and U8764 (N_8764,N_8074,N_8325);
and U8765 (N_8765,N_8116,N_8353);
and U8766 (N_8766,N_8425,N_8238);
nor U8767 (N_8767,N_8470,N_8285);
or U8768 (N_8768,N_8306,N_8413);
nor U8769 (N_8769,N_8388,N_8496);
nor U8770 (N_8770,N_8082,N_8309);
and U8771 (N_8771,N_8079,N_8305);
and U8772 (N_8772,N_8430,N_8224);
and U8773 (N_8773,N_8068,N_8286);
and U8774 (N_8774,N_8096,N_8359);
nor U8775 (N_8775,N_8169,N_8285);
nor U8776 (N_8776,N_8347,N_8330);
and U8777 (N_8777,N_8467,N_8457);
or U8778 (N_8778,N_8100,N_8049);
and U8779 (N_8779,N_8492,N_8015);
and U8780 (N_8780,N_8064,N_8263);
and U8781 (N_8781,N_8315,N_8345);
and U8782 (N_8782,N_8271,N_8357);
nor U8783 (N_8783,N_8049,N_8076);
and U8784 (N_8784,N_8204,N_8187);
or U8785 (N_8785,N_8173,N_8062);
nor U8786 (N_8786,N_8228,N_8435);
and U8787 (N_8787,N_8430,N_8499);
nand U8788 (N_8788,N_8360,N_8298);
and U8789 (N_8789,N_8235,N_8254);
nand U8790 (N_8790,N_8251,N_8111);
and U8791 (N_8791,N_8414,N_8435);
or U8792 (N_8792,N_8130,N_8323);
nand U8793 (N_8793,N_8436,N_8061);
and U8794 (N_8794,N_8467,N_8030);
nand U8795 (N_8795,N_8210,N_8140);
nand U8796 (N_8796,N_8036,N_8337);
nand U8797 (N_8797,N_8054,N_8028);
and U8798 (N_8798,N_8151,N_8187);
nand U8799 (N_8799,N_8220,N_8327);
nand U8800 (N_8800,N_8014,N_8130);
and U8801 (N_8801,N_8237,N_8263);
nand U8802 (N_8802,N_8339,N_8043);
or U8803 (N_8803,N_8028,N_8384);
nor U8804 (N_8804,N_8388,N_8407);
nor U8805 (N_8805,N_8144,N_8428);
or U8806 (N_8806,N_8294,N_8414);
or U8807 (N_8807,N_8106,N_8289);
or U8808 (N_8808,N_8180,N_8281);
and U8809 (N_8809,N_8219,N_8407);
nand U8810 (N_8810,N_8066,N_8138);
or U8811 (N_8811,N_8009,N_8177);
nand U8812 (N_8812,N_8204,N_8296);
or U8813 (N_8813,N_8313,N_8266);
nor U8814 (N_8814,N_8227,N_8300);
nand U8815 (N_8815,N_8202,N_8028);
nor U8816 (N_8816,N_8435,N_8493);
or U8817 (N_8817,N_8415,N_8170);
and U8818 (N_8818,N_8307,N_8071);
and U8819 (N_8819,N_8383,N_8325);
or U8820 (N_8820,N_8447,N_8221);
xnor U8821 (N_8821,N_8134,N_8181);
nor U8822 (N_8822,N_8239,N_8221);
nor U8823 (N_8823,N_8191,N_8361);
and U8824 (N_8824,N_8397,N_8289);
or U8825 (N_8825,N_8301,N_8326);
nor U8826 (N_8826,N_8465,N_8094);
nand U8827 (N_8827,N_8200,N_8051);
nor U8828 (N_8828,N_8168,N_8340);
nand U8829 (N_8829,N_8318,N_8411);
and U8830 (N_8830,N_8360,N_8259);
and U8831 (N_8831,N_8494,N_8024);
nor U8832 (N_8832,N_8202,N_8313);
and U8833 (N_8833,N_8066,N_8070);
or U8834 (N_8834,N_8241,N_8376);
or U8835 (N_8835,N_8050,N_8278);
or U8836 (N_8836,N_8407,N_8253);
nor U8837 (N_8837,N_8400,N_8034);
nor U8838 (N_8838,N_8144,N_8283);
nand U8839 (N_8839,N_8120,N_8029);
nand U8840 (N_8840,N_8217,N_8054);
nand U8841 (N_8841,N_8081,N_8083);
nand U8842 (N_8842,N_8190,N_8174);
or U8843 (N_8843,N_8128,N_8309);
and U8844 (N_8844,N_8457,N_8113);
nand U8845 (N_8845,N_8117,N_8191);
xor U8846 (N_8846,N_8294,N_8377);
nand U8847 (N_8847,N_8023,N_8333);
and U8848 (N_8848,N_8297,N_8016);
and U8849 (N_8849,N_8073,N_8161);
and U8850 (N_8850,N_8459,N_8439);
xor U8851 (N_8851,N_8131,N_8163);
nor U8852 (N_8852,N_8098,N_8343);
or U8853 (N_8853,N_8109,N_8272);
or U8854 (N_8854,N_8186,N_8345);
or U8855 (N_8855,N_8190,N_8133);
and U8856 (N_8856,N_8070,N_8454);
nand U8857 (N_8857,N_8099,N_8459);
nand U8858 (N_8858,N_8455,N_8142);
nand U8859 (N_8859,N_8283,N_8257);
nand U8860 (N_8860,N_8203,N_8052);
and U8861 (N_8861,N_8483,N_8006);
or U8862 (N_8862,N_8303,N_8337);
nand U8863 (N_8863,N_8422,N_8338);
and U8864 (N_8864,N_8139,N_8255);
xnor U8865 (N_8865,N_8440,N_8358);
nand U8866 (N_8866,N_8235,N_8304);
nand U8867 (N_8867,N_8000,N_8276);
nand U8868 (N_8868,N_8445,N_8098);
and U8869 (N_8869,N_8447,N_8269);
nand U8870 (N_8870,N_8022,N_8087);
or U8871 (N_8871,N_8275,N_8303);
nand U8872 (N_8872,N_8260,N_8101);
or U8873 (N_8873,N_8121,N_8202);
nor U8874 (N_8874,N_8072,N_8293);
and U8875 (N_8875,N_8066,N_8456);
and U8876 (N_8876,N_8106,N_8223);
and U8877 (N_8877,N_8046,N_8398);
nor U8878 (N_8878,N_8376,N_8294);
or U8879 (N_8879,N_8269,N_8340);
and U8880 (N_8880,N_8188,N_8042);
nor U8881 (N_8881,N_8128,N_8271);
nor U8882 (N_8882,N_8470,N_8489);
and U8883 (N_8883,N_8041,N_8115);
nor U8884 (N_8884,N_8426,N_8433);
and U8885 (N_8885,N_8421,N_8303);
or U8886 (N_8886,N_8395,N_8333);
nand U8887 (N_8887,N_8041,N_8111);
or U8888 (N_8888,N_8301,N_8402);
nand U8889 (N_8889,N_8013,N_8453);
nor U8890 (N_8890,N_8438,N_8309);
nor U8891 (N_8891,N_8061,N_8275);
or U8892 (N_8892,N_8188,N_8090);
nand U8893 (N_8893,N_8154,N_8078);
nor U8894 (N_8894,N_8431,N_8373);
nand U8895 (N_8895,N_8125,N_8292);
or U8896 (N_8896,N_8211,N_8488);
and U8897 (N_8897,N_8386,N_8369);
nor U8898 (N_8898,N_8124,N_8372);
and U8899 (N_8899,N_8000,N_8185);
or U8900 (N_8900,N_8351,N_8334);
nand U8901 (N_8901,N_8190,N_8343);
or U8902 (N_8902,N_8389,N_8454);
and U8903 (N_8903,N_8136,N_8177);
and U8904 (N_8904,N_8136,N_8405);
or U8905 (N_8905,N_8219,N_8220);
or U8906 (N_8906,N_8239,N_8378);
nor U8907 (N_8907,N_8297,N_8005);
nor U8908 (N_8908,N_8211,N_8281);
or U8909 (N_8909,N_8004,N_8341);
nor U8910 (N_8910,N_8488,N_8470);
and U8911 (N_8911,N_8272,N_8072);
and U8912 (N_8912,N_8204,N_8117);
nor U8913 (N_8913,N_8010,N_8309);
nor U8914 (N_8914,N_8289,N_8440);
or U8915 (N_8915,N_8036,N_8074);
nand U8916 (N_8916,N_8395,N_8049);
xor U8917 (N_8917,N_8035,N_8058);
and U8918 (N_8918,N_8348,N_8396);
nand U8919 (N_8919,N_8487,N_8187);
nor U8920 (N_8920,N_8228,N_8314);
or U8921 (N_8921,N_8088,N_8408);
nand U8922 (N_8922,N_8294,N_8270);
nor U8923 (N_8923,N_8443,N_8173);
or U8924 (N_8924,N_8237,N_8042);
nor U8925 (N_8925,N_8162,N_8155);
nor U8926 (N_8926,N_8461,N_8015);
nor U8927 (N_8927,N_8024,N_8280);
and U8928 (N_8928,N_8279,N_8181);
nand U8929 (N_8929,N_8168,N_8329);
and U8930 (N_8930,N_8136,N_8489);
or U8931 (N_8931,N_8285,N_8293);
nor U8932 (N_8932,N_8011,N_8047);
or U8933 (N_8933,N_8159,N_8077);
and U8934 (N_8934,N_8419,N_8206);
nor U8935 (N_8935,N_8494,N_8168);
nor U8936 (N_8936,N_8364,N_8034);
nor U8937 (N_8937,N_8081,N_8080);
or U8938 (N_8938,N_8093,N_8285);
nand U8939 (N_8939,N_8380,N_8400);
nand U8940 (N_8940,N_8262,N_8182);
xnor U8941 (N_8941,N_8329,N_8095);
nor U8942 (N_8942,N_8395,N_8002);
nand U8943 (N_8943,N_8334,N_8456);
nand U8944 (N_8944,N_8422,N_8212);
nand U8945 (N_8945,N_8432,N_8341);
or U8946 (N_8946,N_8096,N_8335);
nor U8947 (N_8947,N_8396,N_8222);
nand U8948 (N_8948,N_8429,N_8184);
nand U8949 (N_8949,N_8049,N_8320);
nor U8950 (N_8950,N_8257,N_8431);
nor U8951 (N_8951,N_8041,N_8200);
nor U8952 (N_8952,N_8146,N_8309);
nor U8953 (N_8953,N_8082,N_8171);
or U8954 (N_8954,N_8257,N_8235);
nand U8955 (N_8955,N_8041,N_8432);
nor U8956 (N_8956,N_8100,N_8313);
or U8957 (N_8957,N_8273,N_8351);
and U8958 (N_8958,N_8212,N_8305);
nand U8959 (N_8959,N_8002,N_8440);
and U8960 (N_8960,N_8151,N_8172);
nand U8961 (N_8961,N_8427,N_8209);
or U8962 (N_8962,N_8177,N_8377);
nor U8963 (N_8963,N_8091,N_8368);
and U8964 (N_8964,N_8018,N_8407);
nor U8965 (N_8965,N_8228,N_8200);
nor U8966 (N_8966,N_8085,N_8228);
or U8967 (N_8967,N_8174,N_8096);
xor U8968 (N_8968,N_8419,N_8144);
and U8969 (N_8969,N_8080,N_8375);
or U8970 (N_8970,N_8199,N_8263);
or U8971 (N_8971,N_8273,N_8134);
or U8972 (N_8972,N_8129,N_8024);
nand U8973 (N_8973,N_8292,N_8265);
or U8974 (N_8974,N_8468,N_8186);
nor U8975 (N_8975,N_8057,N_8110);
and U8976 (N_8976,N_8205,N_8298);
or U8977 (N_8977,N_8384,N_8484);
nand U8978 (N_8978,N_8088,N_8437);
and U8979 (N_8979,N_8040,N_8097);
and U8980 (N_8980,N_8195,N_8036);
and U8981 (N_8981,N_8022,N_8435);
nor U8982 (N_8982,N_8277,N_8107);
and U8983 (N_8983,N_8448,N_8107);
nor U8984 (N_8984,N_8000,N_8062);
nor U8985 (N_8985,N_8047,N_8403);
nor U8986 (N_8986,N_8030,N_8092);
nor U8987 (N_8987,N_8150,N_8072);
nand U8988 (N_8988,N_8240,N_8087);
or U8989 (N_8989,N_8207,N_8231);
nand U8990 (N_8990,N_8466,N_8233);
and U8991 (N_8991,N_8000,N_8213);
nor U8992 (N_8992,N_8278,N_8450);
and U8993 (N_8993,N_8129,N_8272);
and U8994 (N_8994,N_8420,N_8242);
nor U8995 (N_8995,N_8288,N_8492);
and U8996 (N_8996,N_8269,N_8012);
nand U8997 (N_8997,N_8047,N_8010);
nor U8998 (N_8998,N_8260,N_8354);
nand U8999 (N_8999,N_8011,N_8252);
or U9000 (N_9000,N_8519,N_8982);
nor U9001 (N_9001,N_8994,N_8739);
nor U9002 (N_9002,N_8993,N_8949);
and U9003 (N_9003,N_8680,N_8538);
and U9004 (N_9004,N_8805,N_8533);
and U9005 (N_9005,N_8692,N_8797);
nand U9006 (N_9006,N_8687,N_8572);
nand U9007 (N_9007,N_8975,N_8978);
nor U9008 (N_9008,N_8907,N_8838);
nor U9009 (N_9009,N_8844,N_8900);
nor U9010 (N_9010,N_8537,N_8985);
nand U9011 (N_9011,N_8540,N_8914);
nor U9012 (N_9012,N_8999,N_8765);
nand U9013 (N_9013,N_8862,N_8883);
and U9014 (N_9014,N_8918,N_8749);
nor U9015 (N_9015,N_8700,N_8876);
nand U9016 (N_9016,N_8929,N_8968);
or U9017 (N_9017,N_8758,N_8814);
and U9018 (N_9018,N_8576,N_8516);
nor U9019 (N_9019,N_8926,N_8770);
nor U9020 (N_9020,N_8995,N_8954);
nor U9021 (N_9021,N_8512,N_8768);
or U9022 (N_9022,N_8694,N_8553);
or U9023 (N_9023,N_8984,N_8565);
or U9024 (N_9024,N_8650,N_8901);
nor U9025 (N_9025,N_8950,N_8745);
nand U9026 (N_9026,N_8584,N_8769);
or U9027 (N_9027,N_8737,N_8953);
nand U9028 (N_9028,N_8971,N_8808);
and U9029 (N_9029,N_8956,N_8849);
nand U9030 (N_9030,N_8571,N_8924);
and U9031 (N_9031,N_8515,N_8885);
nand U9032 (N_9032,N_8855,N_8659);
nand U9033 (N_9033,N_8788,N_8641);
and U9034 (N_9034,N_8580,N_8532);
nand U9035 (N_9035,N_8631,N_8558);
or U9036 (N_9036,N_8563,N_8922);
nor U9037 (N_9037,N_8836,N_8939);
nor U9038 (N_9038,N_8996,N_8964);
and U9039 (N_9039,N_8736,N_8643);
nor U9040 (N_9040,N_8630,N_8807);
and U9041 (N_9041,N_8931,N_8709);
and U9042 (N_9042,N_8664,N_8754);
nand U9043 (N_9043,N_8948,N_8895);
or U9044 (N_9044,N_8637,N_8607);
and U9045 (N_9045,N_8791,N_8987);
nor U9046 (N_9046,N_8670,N_8930);
and U9047 (N_9047,N_8545,N_8891);
nand U9048 (N_9048,N_8644,N_8564);
and U9049 (N_9049,N_8861,N_8937);
and U9050 (N_9050,N_8958,N_8748);
nand U9051 (N_9051,N_8648,N_8854);
or U9052 (N_9052,N_8925,N_8916);
or U9053 (N_9053,N_8685,N_8821);
or U9054 (N_9054,N_8899,N_8646);
and U9055 (N_9055,N_8866,N_8542);
nand U9056 (N_9056,N_8662,N_8718);
xnor U9057 (N_9057,N_8973,N_8729);
nand U9058 (N_9058,N_8860,N_8610);
or U9059 (N_9059,N_8823,N_8760);
nor U9060 (N_9060,N_8708,N_8853);
nand U9061 (N_9061,N_8597,N_8651);
or U9062 (N_9062,N_8536,N_8998);
or U9063 (N_9063,N_8503,N_8611);
or U9064 (N_9064,N_8738,N_8882);
or U9065 (N_9065,N_8772,N_8813);
nand U9066 (N_9066,N_8828,N_8714);
or U9067 (N_9067,N_8915,N_8573);
nand U9068 (N_9068,N_8893,N_8568);
and U9069 (N_9069,N_8586,N_8863);
nand U9070 (N_9070,N_8867,N_8661);
nor U9071 (N_9071,N_8645,N_8566);
nor U9072 (N_9072,N_8608,N_8983);
or U9073 (N_9073,N_8609,N_8835);
nor U9074 (N_9074,N_8510,N_8858);
and U9075 (N_9075,N_8679,N_8970);
and U9076 (N_9076,N_8604,N_8703);
or U9077 (N_9077,N_8908,N_8777);
and U9078 (N_9078,N_8546,N_8539);
nand U9079 (N_9079,N_8657,N_8906);
nand U9080 (N_9080,N_8992,N_8957);
and U9081 (N_9081,N_8656,N_8621);
nor U9082 (N_9082,N_8980,N_8795);
nor U9083 (N_9083,N_8549,N_8790);
and U9084 (N_9084,N_8658,N_8603);
nand U9085 (N_9085,N_8582,N_8744);
and U9086 (N_9086,N_8733,N_8585);
nand U9087 (N_9087,N_8668,N_8763);
nor U9088 (N_9088,N_8859,N_8691);
and U9089 (N_9089,N_8640,N_8903);
nand U9090 (N_9090,N_8889,N_8674);
nand U9091 (N_9091,N_8806,N_8706);
nor U9092 (N_9092,N_8921,N_8633);
nand U9093 (N_9093,N_8846,N_8874);
or U9094 (N_9094,N_8775,N_8897);
nand U9095 (N_9095,N_8726,N_8857);
and U9096 (N_9096,N_8653,N_8776);
and U9097 (N_9097,N_8960,N_8872);
nand U9098 (N_9098,N_8551,N_8870);
nor U9099 (N_9099,N_8979,N_8827);
nand U9100 (N_9100,N_8881,N_8675);
nand U9101 (N_9101,N_8552,N_8887);
and U9102 (N_9102,N_8731,N_8762);
nor U9103 (N_9103,N_8505,N_8577);
nor U9104 (N_9104,N_8911,N_8928);
and U9105 (N_9105,N_8719,N_8845);
nor U9106 (N_9106,N_8833,N_8689);
nand U9107 (N_9107,N_8638,N_8819);
or U9108 (N_9108,N_8841,N_8941);
and U9109 (N_9109,N_8636,N_8544);
and U9110 (N_9110,N_8716,N_8773);
nor U9111 (N_9111,N_8753,N_8528);
or U9112 (N_9112,N_8779,N_8919);
and U9113 (N_9113,N_8826,N_8757);
or U9114 (N_9114,N_8781,N_8710);
nand U9115 (N_9115,N_8963,N_8942);
nor U9116 (N_9116,N_8832,N_8780);
nand U9117 (N_9117,N_8940,N_8743);
nand U9118 (N_9118,N_8751,N_8880);
xnor U9119 (N_9119,N_8965,N_8851);
and U9120 (N_9120,N_8829,N_8686);
nand U9121 (N_9121,N_8717,N_8783);
nand U9122 (N_9122,N_8816,N_8683);
nand U9123 (N_9123,N_8628,N_8842);
nor U9124 (N_9124,N_8624,N_8917);
or U9125 (N_9125,N_8688,N_8831);
or U9126 (N_9126,N_8594,N_8713);
or U9127 (N_9127,N_8562,N_8910);
and U9128 (N_9128,N_8678,N_8852);
nand U9129 (N_9129,N_8892,N_8684);
nor U9130 (N_9130,N_8725,N_8521);
nand U9131 (N_9131,N_8967,N_8878);
or U9132 (N_9132,N_8839,N_8974);
nor U9133 (N_9133,N_8531,N_8811);
or U9134 (N_9134,N_8732,N_8701);
nand U9135 (N_9135,N_8825,N_8802);
nor U9136 (N_9136,N_8600,N_8879);
and U9137 (N_9137,N_8561,N_8720);
and U9138 (N_9138,N_8612,N_8617);
nor U9139 (N_9139,N_8752,N_8579);
or U9140 (N_9140,N_8848,N_8567);
nor U9141 (N_9141,N_8856,N_8548);
nor U9142 (N_9142,N_8663,N_8715);
and U9143 (N_9143,N_8933,N_8649);
or U9144 (N_9144,N_8778,N_8988);
and U9145 (N_9145,N_8547,N_8771);
nand U9146 (N_9146,N_8509,N_8697);
and U9147 (N_9147,N_8898,N_8952);
nor U9148 (N_9148,N_8875,N_8599);
nand U9149 (N_9149,N_8755,N_8793);
and U9150 (N_9150,N_8690,N_8969);
nand U9151 (N_9151,N_8810,N_8578);
and U9152 (N_9152,N_8834,N_8696);
nor U9153 (N_9153,N_8747,N_8590);
or U9154 (N_9154,N_8750,N_8961);
or U9155 (N_9155,N_8935,N_8629);
nor U9156 (N_9156,N_8740,N_8976);
nor U9157 (N_9157,N_8837,N_8947);
nand U9158 (N_9158,N_8886,N_8620);
nor U9159 (N_9159,N_8705,N_8587);
or U9160 (N_9160,N_8809,N_8932);
and U9161 (N_9161,N_8523,N_8818);
xor U9162 (N_9162,N_8575,N_8583);
nor U9163 (N_9163,N_8525,N_8873);
nand U9164 (N_9164,N_8824,N_8774);
nor U9165 (N_9165,N_8966,N_8759);
nor U9166 (N_9166,N_8535,N_8981);
nor U9167 (N_9167,N_8634,N_8888);
nor U9168 (N_9168,N_8938,N_8746);
and U9169 (N_9169,N_8792,N_8642);
or U9170 (N_9170,N_8934,N_8991);
or U9171 (N_9171,N_8560,N_8682);
nor U9172 (N_9172,N_8517,N_8506);
nor U9173 (N_9173,N_8677,N_8787);
nor U9174 (N_9174,N_8728,N_8799);
or U9175 (N_9175,N_8555,N_8527);
and U9176 (N_9176,N_8524,N_8672);
nor U9177 (N_9177,N_8785,N_8526);
or U9178 (N_9178,N_8789,N_8800);
nand U9179 (N_9179,N_8616,N_8959);
and U9180 (N_9180,N_8977,N_8518);
and U9181 (N_9181,N_8817,N_8711);
nand U9182 (N_9182,N_8522,N_8721);
nor U9183 (N_9183,N_8511,N_8830);
nand U9184 (N_9184,N_8596,N_8735);
or U9185 (N_9185,N_8798,N_8786);
nor U9186 (N_9186,N_8615,N_8623);
nor U9187 (N_9187,N_8727,N_8507);
nand U9188 (N_9188,N_8554,N_8550);
and U9189 (N_9189,N_8944,N_8588);
nand U9190 (N_9190,N_8822,N_8767);
and U9191 (N_9191,N_8520,N_8734);
nand U9192 (N_9192,N_8592,N_8632);
nor U9193 (N_9193,N_8595,N_8660);
and U9194 (N_9194,N_8766,N_8556);
or U9195 (N_9195,N_8500,N_8671);
and U9196 (N_9196,N_8655,N_8529);
nand U9197 (N_9197,N_8951,N_8943);
and U9198 (N_9198,N_8912,N_8639);
nand U9199 (N_9199,N_8896,N_8782);
or U9200 (N_9200,N_8847,N_8724);
or U9201 (N_9201,N_8865,N_8756);
xnor U9202 (N_9202,N_8581,N_8986);
or U9203 (N_9203,N_8614,N_8635);
nor U9204 (N_9204,N_8804,N_8574);
and U9205 (N_9205,N_8955,N_8619);
nor U9206 (N_9206,N_8902,N_8626);
and U9207 (N_9207,N_8815,N_8894);
nand U9208 (N_9208,N_8723,N_8869);
nor U9209 (N_9209,N_8764,N_8606);
nand U9210 (N_9210,N_8702,N_8840);
nand U9211 (N_9211,N_8654,N_8598);
or U9212 (N_9212,N_8864,N_8508);
nand U9213 (N_9213,N_8707,N_8534);
and U9214 (N_9214,N_8559,N_8890);
nand U9215 (N_9215,N_8920,N_8681);
nand U9216 (N_9216,N_8936,N_8652);
or U9217 (N_9217,N_8905,N_8820);
or U9218 (N_9218,N_8673,N_8990);
nor U9219 (N_9219,N_8923,N_8794);
or U9220 (N_9220,N_8543,N_8741);
nand U9221 (N_9221,N_8667,N_8502);
or U9222 (N_9222,N_8627,N_8695);
nor U9223 (N_9223,N_8593,N_8843);
or U9224 (N_9224,N_8945,N_8812);
nand U9225 (N_9225,N_8504,N_8784);
and U9226 (N_9226,N_8676,N_8850);
nor U9227 (N_9227,N_8803,N_8946);
and U9228 (N_9228,N_8962,N_8699);
or U9229 (N_9229,N_8722,N_8570);
nor U9230 (N_9230,N_8589,N_8557);
nand U9231 (N_9231,N_8602,N_8613);
nor U9232 (N_9232,N_8927,N_8904);
nor U9233 (N_9233,N_8877,N_8665);
nand U9234 (N_9234,N_8972,N_8730);
nand U9235 (N_9235,N_8513,N_8989);
or U9236 (N_9236,N_8647,N_8625);
xnor U9237 (N_9237,N_8997,N_8796);
nand U9238 (N_9238,N_8591,N_8501);
and U9239 (N_9239,N_8666,N_8530);
nand U9240 (N_9240,N_8712,N_8622);
and U9241 (N_9241,N_8541,N_8909);
or U9242 (N_9242,N_8698,N_8601);
nand U9243 (N_9243,N_8871,N_8669);
and U9244 (N_9244,N_8605,N_8761);
nor U9245 (N_9245,N_8868,N_8569);
or U9246 (N_9246,N_8693,N_8514);
or U9247 (N_9247,N_8742,N_8801);
and U9248 (N_9248,N_8913,N_8704);
and U9249 (N_9249,N_8884,N_8618);
and U9250 (N_9250,N_8994,N_8934);
and U9251 (N_9251,N_8992,N_8947);
and U9252 (N_9252,N_8624,N_8501);
nand U9253 (N_9253,N_8817,N_8513);
and U9254 (N_9254,N_8878,N_8728);
nor U9255 (N_9255,N_8767,N_8645);
or U9256 (N_9256,N_8969,N_8588);
nor U9257 (N_9257,N_8702,N_8651);
nand U9258 (N_9258,N_8520,N_8999);
or U9259 (N_9259,N_8729,N_8841);
and U9260 (N_9260,N_8616,N_8707);
nor U9261 (N_9261,N_8544,N_8978);
and U9262 (N_9262,N_8864,N_8557);
nand U9263 (N_9263,N_8619,N_8839);
or U9264 (N_9264,N_8581,N_8842);
nand U9265 (N_9265,N_8590,N_8662);
nand U9266 (N_9266,N_8535,N_8589);
nand U9267 (N_9267,N_8975,N_8601);
or U9268 (N_9268,N_8542,N_8686);
or U9269 (N_9269,N_8500,N_8773);
or U9270 (N_9270,N_8805,N_8645);
nor U9271 (N_9271,N_8629,N_8906);
nor U9272 (N_9272,N_8611,N_8786);
xnor U9273 (N_9273,N_8626,N_8832);
or U9274 (N_9274,N_8769,N_8784);
xnor U9275 (N_9275,N_8670,N_8634);
nand U9276 (N_9276,N_8812,N_8642);
or U9277 (N_9277,N_8500,N_8626);
nor U9278 (N_9278,N_8978,N_8655);
nand U9279 (N_9279,N_8954,N_8710);
xnor U9280 (N_9280,N_8912,N_8962);
nand U9281 (N_9281,N_8536,N_8877);
and U9282 (N_9282,N_8792,N_8564);
and U9283 (N_9283,N_8666,N_8726);
or U9284 (N_9284,N_8794,N_8980);
nor U9285 (N_9285,N_8706,N_8781);
nor U9286 (N_9286,N_8874,N_8818);
nand U9287 (N_9287,N_8681,N_8936);
and U9288 (N_9288,N_8801,N_8577);
nor U9289 (N_9289,N_8664,N_8637);
nor U9290 (N_9290,N_8755,N_8738);
and U9291 (N_9291,N_8963,N_8958);
nand U9292 (N_9292,N_8885,N_8661);
and U9293 (N_9293,N_8502,N_8611);
nand U9294 (N_9294,N_8984,N_8549);
and U9295 (N_9295,N_8715,N_8775);
nand U9296 (N_9296,N_8608,N_8798);
or U9297 (N_9297,N_8936,N_8507);
and U9298 (N_9298,N_8895,N_8788);
or U9299 (N_9299,N_8624,N_8945);
nand U9300 (N_9300,N_8594,N_8710);
nand U9301 (N_9301,N_8920,N_8817);
nand U9302 (N_9302,N_8898,N_8777);
nor U9303 (N_9303,N_8560,N_8993);
nor U9304 (N_9304,N_8554,N_8882);
xor U9305 (N_9305,N_8742,N_8695);
nor U9306 (N_9306,N_8721,N_8753);
nand U9307 (N_9307,N_8951,N_8568);
nor U9308 (N_9308,N_8680,N_8548);
and U9309 (N_9309,N_8728,N_8755);
nor U9310 (N_9310,N_8693,N_8568);
or U9311 (N_9311,N_8902,N_8699);
nor U9312 (N_9312,N_8597,N_8826);
and U9313 (N_9313,N_8826,N_8825);
and U9314 (N_9314,N_8749,N_8630);
and U9315 (N_9315,N_8950,N_8957);
nand U9316 (N_9316,N_8582,N_8960);
or U9317 (N_9317,N_8649,N_8554);
or U9318 (N_9318,N_8781,N_8504);
nand U9319 (N_9319,N_8999,N_8518);
and U9320 (N_9320,N_8691,N_8698);
nor U9321 (N_9321,N_8814,N_8997);
and U9322 (N_9322,N_8779,N_8884);
and U9323 (N_9323,N_8793,N_8746);
nand U9324 (N_9324,N_8546,N_8715);
nor U9325 (N_9325,N_8679,N_8878);
or U9326 (N_9326,N_8931,N_8894);
nor U9327 (N_9327,N_8855,N_8895);
nand U9328 (N_9328,N_8773,N_8664);
nand U9329 (N_9329,N_8559,N_8995);
nand U9330 (N_9330,N_8515,N_8997);
and U9331 (N_9331,N_8525,N_8999);
xnor U9332 (N_9332,N_8814,N_8787);
and U9333 (N_9333,N_8969,N_8550);
nor U9334 (N_9334,N_8846,N_8528);
nor U9335 (N_9335,N_8564,N_8691);
and U9336 (N_9336,N_8988,N_8780);
nor U9337 (N_9337,N_8724,N_8869);
nand U9338 (N_9338,N_8932,N_8704);
nand U9339 (N_9339,N_8517,N_8575);
nand U9340 (N_9340,N_8632,N_8870);
nor U9341 (N_9341,N_8571,N_8765);
or U9342 (N_9342,N_8845,N_8809);
nand U9343 (N_9343,N_8642,N_8817);
nand U9344 (N_9344,N_8643,N_8794);
nand U9345 (N_9345,N_8855,N_8789);
nor U9346 (N_9346,N_8595,N_8969);
and U9347 (N_9347,N_8964,N_8766);
nor U9348 (N_9348,N_8966,N_8603);
nand U9349 (N_9349,N_8685,N_8512);
and U9350 (N_9350,N_8533,N_8887);
and U9351 (N_9351,N_8935,N_8688);
nor U9352 (N_9352,N_8774,N_8949);
nor U9353 (N_9353,N_8967,N_8882);
nand U9354 (N_9354,N_8760,N_8697);
or U9355 (N_9355,N_8764,N_8549);
nand U9356 (N_9356,N_8916,N_8744);
nor U9357 (N_9357,N_8586,N_8870);
nand U9358 (N_9358,N_8577,N_8696);
nand U9359 (N_9359,N_8939,N_8888);
or U9360 (N_9360,N_8661,N_8738);
nor U9361 (N_9361,N_8675,N_8949);
nand U9362 (N_9362,N_8749,N_8923);
nand U9363 (N_9363,N_8988,N_8881);
nor U9364 (N_9364,N_8738,N_8624);
nor U9365 (N_9365,N_8619,N_8539);
nor U9366 (N_9366,N_8559,N_8521);
or U9367 (N_9367,N_8827,N_8508);
and U9368 (N_9368,N_8816,N_8736);
and U9369 (N_9369,N_8910,N_8789);
and U9370 (N_9370,N_8804,N_8625);
or U9371 (N_9371,N_8752,N_8956);
nand U9372 (N_9372,N_8712,N_8921);
and U9373 (N_9373,N_8774,N_8910);
nand U9374 (N_9374,N_8822,N_8970);
nand U9375 (N_9375,N_8995,N_8700);
and U9376 (N_9376,N_8898,N_8984);
or U9377 (N_9377,N_8858,N_8951);
nand U9378 (N_9378,N_8840,N_8583);
and U9379 (N_9379,N_8986,N_8586);
nand U9380 (N_9380,N_8740,N_8861);
nand U9381 (N_9381,N_8588,N_8668);
or U9382 (N_9382,N_8650,N_8811);
and U9383 (N_9383,N_8810,N_8933);
and U9384 (N_9384,N_8631,N_8821);
and U9385 (N_9385,N_8872,N_8515);
nor U9386 (N_9386,N_8520,N_8709);
or U9387 (N_9387,N_8556,N_8820);
or U9388 (N_9388,N_8725,N_8990);
nor U9389 (N_9389,N_8555,N_8740);
nor U9390 (N_9390,N_8709,N_8919);
nor U9391 (N_9391,N_8819,N_8864);
nor U9392 (N_9392,N_8591,N_8734);
nand U9393 (N_9393,N_8728,N_8637);
nand U9394 (N_9394,N_8982,N_8708);
nor U9395 (N_9395,N_8951,N_8696);
or U9396 (N_9396,N_8885,N_8595);
nand U9397 (N_9397,N_8581,N_8863);
nor U9398 (N_9398,N_8516,N_8934);
nor U9399 (N_9399,N_8908,N_8715);
and U9400 (N_9400,N_8842,N_8736);
and U9401 (N_9401,N_8909,N_8651);
or U9402 (N_9402,N_8997,N_8731);
nand U9403 (N_9403,N_8708,N_8781);
and U9404 (N_9404,N_8987,N_8836);
and U9405 (N_9405,N_8991,N_8683);
and U9406 (N_9406,N_8956,N_8841);
and U9407 (N_9407,N_8761,N_8839);
xnor U9408 (N_9408,N_8978,N_8763);
or U9409 (N_9409,N_8888,N_8752);
or U9410 (N_9410,N_8898,N_8753);
nor U9411 (N_9411,N_8925,N_8735);
nor U9412 (N_9412,N_8778,N_8965);
or U9413 (N_9413,N_8810,N_8851);
nand U9414 (N_9414,N_8851,N_8778);
nor U9415 (N_9415,N_8816,N_8738);
nand U9416 (N_9416,N_8546,N_8563);
or U9417 (N_9417,N_8909,N_8716);
nor U9418 (N_9418,N_8516,N_8946);
or U9419 (N_9419,N_8881,N_8714);
or U9420 (N_9420,N_8639,N_8975);
nor U9421 (N_9421,N_8844,N_8586);
nor U9422 (N_9422,N_8784,N_8604);
nor U9423 (N_9423,N_8836,N_8849);
nor U9424 (N_9424,N_8713,N_8808);
or U9425 (N_9425,N_8600,N_8748);
nand U9426 (N_9426,N_8670,N_8520);
and U9427 (N_9427,N_8876,N_8517);
nor U9428 (N_9428,N_8545,N_8635);
or U9429 (N_9429,N_8977,N_8906);
nand U9430 (N_9430,N_8621,N_8794);
or U9431 (N_9431,N_8903,N_8637);
nor U9432 (N_9432,N_8968,N_8625);
nand U9433 (N_9433,N_8597,N_8787);
nand U9434 (N_9434,N_8863,N_8664);
or U9435 (N_9435,N_8653,N_8505);
nor U9436 (N_9436,N_8740,N_8985);
nand U9437 (N_9437,N_8654,N_8702);
nand U9438 (N_9438,N_8578,N_8527);
and U9439 (N_9439,N_8645,N_8680);
nand U9440 (N_9440,N_8945,N_8930);
nand U9441 (N_9441,N_8842,N_8752);
and U9442 (N_9442,N_8912,N_8928);
or U9443 (N_9443,N_8910,N_8746);
and U9444 (N_9444,N_8906,N_8776);
nand U9445 (N_9445,N_8952,N_8980);
and U9446 (N_9446,N_8605,N_8721);
nand U9447 (N_9447,N_8881,N_8862);
nand U9448 (N_9448,N_8728,N_8555);
and U9449 (N_9449,N_8656,N_8920);
and U9450 (N_9450,N_8879,N_8631);
nor U9451 (N_9451,N_8591,N_8882);
and U9452 (N_9452,N_8718,N_8819);
nand U9453 (N_9453,N_8516,N_8978);
or U9454 (N_9454,N_8761,N_8613);
nand U9455 (N_9455,N_8821,N_8694);
and U9456 (N_9456,N_8777,N_8769);
or U9457 (N_9457,N_8534,N_8948);
or U9458 (N_9458,N_8916,N_8516);
and U9459 (N_9459,N_8971,N_8877);
nand U9460 (N_9460,N_8947,N_8650);
or U9461 (N_9461,N_8909,N_8602);
nor U9462 (N_9462,N_8593,N_8634);
and U9463 (N_9463,N_8777,N_8770);
and U9464 (N_9464,N_8874,N_8841);
nand U9465 (N_9465,N_8837,N_8940);
nand U9466 (N_9466,N_8902,N_8849);
and U9467 (N_9467,N_8881,N_8706);
or U9468 (N_9468,N_8566,N_8738);
nor U9469 (N_9469,N_8994,N_8999);
and U9470 (N_9470,N_8866,N_8608);
nor U9471 (N_9471,N_8586,N_8747);
and U9472 (N_9472,N_8934,N_8834);
nand U9473 (N_9473,N_8684,N_8623);
and U9474 (N_9474,N_8703,N_8501);
nand U9475 (N_9475,N_8991,N_8983);
or U9476 (N_9476,N_8755,N_8913);
nand U9477 (N_9477,N_8691,N_8648);
and U9478 (N_9478,N_8869,N_8810);
nor U9479 (N_9479,N_8552,N_8650);
nand U9480 (N_9480,N_8868,N_8955);
and U9481 (N_9481,N_8953,N_8614);
nor U9482 (N_9482,N_8976,N_8658);
nand U9483 (N_9483,N_8615,N_8863);
or U9484 (N_9484,N_8661,N_8978);
and U9485 (N_9485,N_8558,N_8510);
or U9486 (N_9486,N_8860,N_8809);
or U9487 (N_9487,N_8578,N_8693);
or U9488 (N_9488,N_8640,N_8688);
or U9489 (N_9489,N_8718,N_8836);
or U9490 (N_9490,N_8962,N_8707);
or U9491 (N_9491,N_8523,N_8857);
nor U9492 (N_9492,N_8706,N_8577);
xnor U9493 (N_9493,N_8775,N_8656);
nor U9494 (N_9494,N_8648,N_8997);
nand U9495 (N_9495,N_8724,N_8866);
and U9496 (N_9496,N_8598,N_8967);
nand U9497 (N_9497,N_8506,N_8546);
and U9498 (N_9498,N_8517,N_8847);
nor U9499 (N_9499,N_8597,N_8864);
or U9500 (N_9500,N_9489,N_9429);
or U9501 (N_9501,N_9089,N_9474);
nor U9502 (N_9502,N_9209,N_9044);
nor U9503 (N_9503,N_9085,N_9081);
or U9504 (N_9504,N_9002,N_9494);
and U9505 (N_9505,N_9203,N_9420);
nand U9506 (N_9506,N_9094,N_9330);
nand U9507 (N_9507,N_9374,N_9376);
and U9508 (N_9508,N_9234,N_9445);
nor U9509 (N_9509,N_9274,N_9497);
xnor U9510 (N_9510,N_9174,N_9096);
nand U9511 (N_9511,N_9216,N_9242);
and U9512 (N_9512,N_9390,N_9295);
nor U9513 (N_9513,N_9286,N_9208);
nor U9514 (N_9514,N_9112,N_9326);
nor U9515 (N_9515,N_9364,N_9181);
and U9516 (N_9516,N_9224,N_9443);
and U9517 (N_9517,N_9073,N_9438);
or U9518 (N_9518,N_9090,N_9289);
or U9519 (N_9519,N_9393,N_9460);
and U9520 (N_9520,N_9177,N_9426);
and U9521 (N_9521,N_9206,N_9187);
nor U9522 (N_9522,N_9037,N_9389);
and U9523 (N_9523,N_9010,N_9086);
nand U9524 (N_9524,N_9023,N_9196);
nand U9525 (N_9525,N_9465,N_9457);
nor U9526 (N_9526,N_9146,N_9225);
or U9527 (N_9527,N_9228,N_9396);
nor U9528 (N_9528,N_9333,N_9188);
or U9529 (N_9529,N_9098,N_9257);
nand U9530 (N_9530,N_9031,N_9113);
nand U9531 (N_9531,N_9323,N_9373);
and U9532 (N_9532,N_9012,N_9276);
nand U9533 (N_9533,N_9487,N_9329);
xor U9534 (N_9534,N_9210,N_9264);
nand U9535 (N_9535,N_9418,N_9381);
nand U9536 (N_9536,N_9054,N_9045);
and U9537 (N_9537,N_9104,N_9256);
nand U9538 (N_9538,N_9442,N_9356);
nor U9539 (N_9539,N_9353,N_9130);
nand U9540 (N_9540,N_9214,N_9284);
or U9541 (N_9541,N_9265,N_9447);
nand U9542 (N_9542,N_9229,N_9278);
nand U9543 (N_9543,N_9122,N_9009);
and U9544 (N_9544,N_9360,N_9307);
nor U9545 (N_9545,N_9271,N_9392);
nor U9546 (N_9546,N_9036,N_9022);
nor U9547 (N_9547,N_9431,N_9472);
or U9548 (N_9548,N_9111,N_9316);
nand U9549 (N_9549,N_9170,N_9064);
nor U9550 (N_9550,N_9499,N_9127);
nand U9551 (N_9551,N_9154,N_9239);
or U9552 (N_9552,N_9145,N_9056);
or U9553 (N_9553,N_9369,N_9118);
and U9554 (N_9554,N_9491,N_9101);
nand U9555 (N_9555,N_9144,N_9245);
nor U9556 (N_9556,N_9133,N_9226);
nand U9557 (N_9557,N_9252,N_9412);
nor U9558 (N_9558,N_9057,N_9071);
and U9559 (N_9559,N_9117,N_9195);
or U9560 (N_9560,N_9476,N_9379);
nor U9561 (N_9561,N_9223,N_9268);
and U9562 (N_9562,N_9190,N_9046);
nor U9563 (N_9563,N_9424,N_9299);
and U9564 (N_9564,N_9281,N_9346);
and U9565 (N_9565,N_9151,N_9291);
xnor U9566 (N_9566,N_9018,N_9027);
xnor U9567 (N_9567,N_9157,N_9495);
nand U9568 (N_9568,N_9490,N_9213);
nor U9569 (N_9569,N_9074,N_9033);
nand U9570 (N_9570,N_9132,N_9449);
nor U9571 (N_9571,N_9029,N_9298);
nand U9572 (N_9572,N_9266,N_9032);
and U9573 (N_9573,N_9082,N_9158);
or U9574 (N_9574,N_9425,N_9315);
and U9575 (N_9575,N_9149,N_9125);
nand U9576 (N_9576,N_9019,N_9391);
or U9577 (N_9577,N_9419,N_9070);
and U9578 (N_9578,N_9231,N_9128);
nand U9579 (N_9579,N_9302,N_9183);
nand U9580 (N_9580,N_9131,N_9484);
and U9581 (N_9581,N_9359,N_9279);
nand U9582 (N_9582,N_9290,N_9338);
or U9583 (N_9583,N_9218,N_9382);
nand U9584 (N_9584,N_9087,N_9446);
and U9585 (N_9585,N_9479,N_9292);
and U9586 (N_9586,N_9314,N_9088);
or U9587 (N_9587,N_9380,N_9141);
and U9588 (N_9588,N_9212,N_9428);
nor U9589 (N_9589,N_9237,N_9017);
xor U9590 (N_9590,N_9365,N_9304);
or U9591 (N_9591,N_9232,N_9435);
nor U9592 (N_9592,N_9439,N_9058);
nor U9593 (N_9593,N_9053,N_9186);
nand U9594 (N_9594,N_9093,N_9403);
or U9595 (N_9595,N_9349,N_9282);
nand U9596 (N_9596,N_9025,N_9475);
and U9597 (N_9597,N_9341,N_9191);
and U9598 (N_9598,N_9319,N_9189);
and U9599 (N_9599,N_9202,N_9395);
nor U9600 (N_9600,N_9034,N_9411);
and U9601 (N_9601,N_9005,N_9318);
nand U9602 (N_9602,N_9253,N_9312);
or U9603 (N_9603,N_9347,N_9417);
and U9604 (N_9604,N_9115,N_9003);
nand U9605 (N_9605,N_9423,N_9059);
nand U9606 (N_9606,N_9168,N_9311);
and U9607 (N_9607,N_9348,N_9357);
nand U9608 (N_9608,N_9105,N_9397);
or U9609 (N_9609,N_9272,N_9211);
and U9610 (N_9610,N_9296,N_9467);
and U9611 (N_9611,N_9452,N_9163);
nand U9612 (N_9612,N_9076,N_9135);
nand U9613 (N_9613,N_9325,N_9416);
nand U9614 (N_9614,N_9477,N_9481);
nand U9615 (N_9615,N_9173,N_9159);
nand U9616 (N_9616,N_9335,N_9126);
and U9617 (N_9617,N_9028,N_9204);
nor U9618 (N_9618,N_9107,N_9180);
nor U9619 (N_9619,N_9062,N_9421);
and U9620 (N_9620,N_9124,N_9148);
or U9621 (N_9621,N_9167,N_9109);
nand U9622 (N_9622,N_9102,N_9184);
or U9623 (N_9623,N_9415,N_9493);
or U9624 (N_9624,N_9337,N_9176);
or U9625 (N_9625,N_9331,N_9235);
and U9626 (N_9626,N_9249,N_9197);
or U9627 (N_9627,N_9116,N_9079);
nor U9628 (N_9628,N_9041,N_9440);
nor U9629 (N_9629,N_9134,N_9459);
or U9630 (N_9630,N_9138,N_9372);
or U9631 (N_9631,N_9466,N_9358);
and U9632 (N_9632,N_9297,N_9354);
nor U9633 (N_9633,N_9065,N_9377);
nor U9634 (N_9634,N_9014,N_9336);
and U9635 (N_9635,N_9114,N_9166);
and U9636 (N_9636,N_9024,N_9273);
nand U9637 (N_9637,N_9285,N_9280);
nand U9638 (N_9638,N_9498,N_9456);
and U9639 (N_9639,N_9039,N_9251);
and U9640 (N_9640,N_9152,N_9207);
and U9641 (N_9641,N_9258,N_9080);
nor U9642 (N_9642,N_9370,N_9201);
and U9643 (N_9643,N_9436,N_9077);
nand U9644 (N_9644,N_9355,N_9006);
or U9645 (N_9645,N_9063,N_9048);
nor U9646 (N_9646,N_9255,N_9488);
nand U9647 (N_9647,N_9066,N_9451);
nand U9648 (N_9648,N_9000,N_9454);
nor U9649 (N_9649,N_9156,N_9486);
or U9650 (N_9650,N_9362,N_9342);
nor U9651 (N_9651,N_9496,N_9378);
and U9652 (N_9652,N_9406,N_9461);
and U9653 (N_9653,N_9328,N_9471);
nand U9654 (N_9654,N_9061,N_9055);
or U9655 (N_9655,N_9433,N_9069);
nand U9656 (N_9656,N_9480,N_9227);
and U9657 (N_9657,N_9339,N_9247);
xnor U9658 (N_9658,N_9343,N_9453);
nor U9659 (N_9659,N_9040,N_9143);
nor U9660 (N_9660,N_9404,N_9222);
nand U9661 (N_9661,N_9482,N_9261);
nand U9662 (N_9662,N_9269,N_9084);
and U9663 (N_9663,N_9473,N_9468);
and U9664 (N_9664,N_9244,N_9147);
or U9665 (N_9665,N_9007,N_9260);
or U9666 (N_9666,N_9463,N_9016);
and U9667 (N_9667,N_9165,N_9434);
and U9668 (N_9668,N_9388,N_9215);
and U9669 (N_9669,N_9368,N_9240);
or U9670 (N_9670,N_9198,N_9363);
nand U9671 (N_9671,N_9178,N_9169);
nor U9672 (N_9672,N_9366,N_9413);
and U9673 (N_9673,N_9175,N_9427);
nand U9674 (N_9674,N_9386,N_9092);
nor U9675 (N_9675,N_9004,N_9345);
xnor U9676 (N_9676,N_9309,N_9437);
nor U9677 (N_9677,N_9052,N_9095);
nor U9678 (N_9678,N_9485,N_9038);
or U9679 (N_9679,N_9294,N_9430);
and U9680 (N_9680,N_9327,N_9230);
and U9681 (N_9681,N_9020,N_9217);
nor U9682 (N_9682,N_9091,N_9120);
nor U9683 (N_9683,N_9097,N_9350);
nand U9684 (N_9684,N_9008,N_9030);
nor U9685 (N_9685,N_9469,N_9385);
or U9686 (N_9686,N_9361,N_9409);
nor U9687 (N_9687,N_9241,N_9047);
nand U9688 (N_9688,N_9283,N_9317);
xor U9689 (N_9689,N_9246,N_9121);
or U9690 (N_9690,N_9137,N_9262);
and U9691 (N_9691,N_9321,N_9001);
nor U9692 (N_9692,N_9219,N_9136);
xor U9693 (N_9693,N_9155,N_9248);
or U9694 (N_9694,N_9060,N_9313);
nand U9695 (N_9695,N_9194,N_9103);
and U9696 (N_9696,N_9172,N_9332);
or U9697 (N_9697,N_9351,N_9171);
and U9698 (N_9698,N_9287,N_9123);
or U9699 (N_9699,N_9049,N_9402);
and U9700 (N_9700,N_9051,N_9387);
and U9701 (N_9701,N_9305,N_9205);
and U9702 (N_9702,N_9042,N_9455);
nor U9703 (N_9703,N_9384,N_9250);
nor U9704 (N_9704,N_9015,N_9043);
nor U9705 (N_9705,N_9310,N_9221);
and U9706 (N_9706,N_9021,N_9450);
nor U9707 (N_9707,N_9199,N_9078);
and U9708 (N_9708,N_9410,N_9236);
and U9709 (N_9709,N_9407,N_9129);
nand U9710 (N_9710,N_9013,N_9142);
and U9711 (N_9711,N_9394,N_9324);
or U9712 (N_9712,N_9026,N_9448);
and U9713 (N_9713,N_9153,N_9140);
nor U9714 (N_9714,N_9344,N_9259);
and U9715 (N_9715,N_9422,N_9139);
nor U9716 (N_9716,N_9306,N_9301);
nand U9717 (N_9717,N_9099,N_9400);
nand U9718 (N_9718,N_9414,N_9200);
and U9719 (N_9719,N_9320,N_9160);
nand U9720 (N_9720,N_9185,N_9408);
nor U9721 (N_9721,N_9100,N_9263);
xnor U9722 (N_9722,N_9270,N_9288);
and U9723 (N_9723,N_9444,N_9110);
xor U9724 (N_9724,N_9182,N_9322);
or U9725 (N_9725,N_9164,N_9106);
and U9726 (N_9726,N_9068,N_9119);
and U9727 (N_9727,N_9367,N_9193);
or U9728 (N_9728,N_9483,N_9308);
or U9729 (N_9729,N_9050,N_9192);
and U9730 (N_9730,N_9478,N_9401);
xnor U9731 (N_9731,N_9075,N_9300);
nor U9732 (N_9732,N_9220,N_9162);
nor U9733 (N_9733,N_9462,N_9067);
nand U9734 (N_9734,N_9035,N_9293);
or U9735 (N_9735,N_9432,N_9243);
nor U9736 (N_9736,N_9072,N_9405);
or U9737 (N_9737,N_9340,N_9150);
nand U9738 (N_9738,N_9275,N_9254);
nor U9739 (N_9739,N_9371,N_9233);
nand U9740 (N_9740,N_9470,N_9161);
or U9741 (N_9741,N_9399,N_9267);
and U9742 (N_9742,N_9303,N_9375);
nor U9743 (N_9743,N_9398,N_9334);
nand U9744 (N_9744,N_9238,N_9441);
nand U9745 (N_9745,N_9108,N_9464);
or U9746 (N_9746,N_9083,N_9352);
nand U9747 (N_9747,N_9492,N_9458);
nor U9748 (N_9748,N_9179,N_9277);
and U9749 (N_9749,N_9011,N_9383);
xnor U9750 (N_9750,N_9252,N_9240);
nor U9751 (N_9751,N_9003,N_9117);
nor U9752 (N_9752,N_9026,N_9073);
and U9753 (N_9753,N_9151,N_9025);
nand U9754 (N_9754,N_9105,N_9435);
and U9755 (N_9755,N_9025,N_9340);
or U9756 (N_9756,N_9120,N_9439);
and U9757 (N_9757,N_9224,N_9017);
and U9758 (N_9758,N_9053,N_9147);
or U9759 (N_9759,N_9062,N_9435);
or U9760 (N_9760,N_9331,N_9329);
or U9761 (N_9761,N_9490,N_9233);
nand U9762 (N_9762,N_9096,N_9086);
and U9763 (N_9763,N_9328,N_9100);
nor U9764 (N_9764,N_9003,N_9337);
or U9765 (N_9765,N_9079,N_9387);
nand U9766 (N_9766,N_9309,N_9490);
or U9767 (N_9767,N_9483,N_9281);
or U9768 (N_9768,N_9444,N_9405);
nor U9769 (N_9769,N_9380,N_9230);
or U9770 (N_9770,N_9321,N_9250);
or U9771 (N_9771,N_9258,N_9260);
or U9772 (N_9772,N_9052,N_9279);
or U9773 (N_9773,N_9164,N_9473);
or U9774 (N_9774,N_9442,N_9359);
or U9775 (N_9775,N_9184,N_9318);
or U9776 (N_9776,N_9334,N_9248);
and U9777 (N_9777,N_9327,N_9460);
nand U9778 (N_9778,N_9014,N_9030);
nand U9779 (N_9779,N_9414,N_9425);
or U9780 (N_9780,N_9059,N_9188);
nand U9781 (N_9781,N_9199,N_9364);
nor U9782 (N_9782,N_9182,N_9302);
nand U9783 (N_9783,N_9206,N_9339);
or U9784 (N_9784,N_9250,N_9288);
and U9785 (N_9785,N_9371,N_9297);
nand U9786 (N_9786,N_9465,N_9150);
and U9787 (N_9787,N_9307,N_9339);
and U9788 (N_9788,N_9006,N_9329);
nor U9789 (N_9789,N_9046,N_9144);
or U9790 (N_9790,N_9327,N_9160);
nor U9791 (N_9791,N_9374,N_9360);
or U9792 (N_9792,N_9305,N_9373);
nand U9793 (N_9793,N_9497,N_9037);
and U9794 (N_9794,N_9302,N_9144);
nand U9795 (N_9795,N_9385,N_9347);
nor U9796 (N_9796,N_9252,N_9392);
and U9797 (N_9797,N_9491,N_9020);
nor U9798 (N_9798,N_9194,N_9091);
and U9799 (N_9799,N_9045,N_9302);
nand U9800 (N_9800,N_9190,N_9102);
nor U9801 (N_9801,N_9089,N_9459);
nand U9802 (N_9802,N_9224,N_9244);
nor U9803 (N_9803,N_9079,N_9321);
nor U9804 (N_9804,N_9077,N_9081);
nor U9805 (N_9805,N_9439,N_9297);
and U9806 (N_9806,N_9129,N_9274);
and U9807 (N_9807,N_9118,N_9212);
nand U9808 (N_9808,N_9000,N_9085);
and U9809 (N_9809,N_9274,N_9373);
nor U9810 (N_9810,N_9312,N_9202);
nor U9811 (N_9811,N_9349,N_9471);
and U9812 (N_9812,N_9499,N_9086);
nand U9813 (N_9813,N_9299,N_9129);
nor U9814 (N_9814,N_9441,N_9205);
nor U9815 (N_9815,N_9296,N_9086);
nand U9816 (N_9816,N_9416,N_9459);
and U9817 (N_9817,N_9236,N_9139);
and U9818 (N_9818,N_9133,N_9147);
nand U9819 (N_9819,N_9173,N_9233);
or U9820 (N_9820,N_9022,N_9130);
nor U9821 (N_9821,N_9169,N_9166);
nand U9822 (N_9822,N_9288,N_9463);
nor U9823 (N_9823,N_9019,N_9241);
or U9824 (N_9824,N_9347,N_9047);
or U9825 (N_9825,N_9148,N_9366);
and U9826 (N_9826,N_9382,N_9471);
nand U9827 (N_9827,N_9470,N_9473);
nand U9828 (N_9828,N_9263,N_9385);
xnor U9829 (N_9829,N_9289,N_9403);
and U9830 (N_9830,N_9119,N_9400);
xnor U9831 (N_9831,N_9459,N_9160);
or U9832 (N_9832,N_9252,N_9372);
and U9833 (N_9833,N_9256,N_9426);
or U9834 (N_9834,N_9438,N_9057);
nor U9835 (N_9835,N_9108,N_9103);
nor U9836 (N_9836,N_9010,N_9483);
and U9837 (N_9837,N_9365,N_9182);
or U9838 (N_9838,N_9442,N_9184);
nand U9839 (N_9839,N_9188,N_9401);
or U9840 (N_9840,N_9052,N_9441);
nand U9841 (N_9841,N_9208,N_9424);
nor U9842 (N_9842,N_9049,N_9115);
or U9843 (N_9843,N_9345,N_9431);
nor U9844 (N_9844,N_9077,N_9340);
nor U9845 (N_9845,N_9475,N_9039);
nand U9846 (N_9846,N_9442,N_9252);
nand U9847 (N_9847,N_9320,N_9063);
nand U9848 (N_9848,N_9163,N_9410);
nor U9849 (N_9849,N_9389,N_9358);
or U9850 (N_9850,N_9499,N_9410);
or U9851 (N_9851,N_9367,N_9185);
or U9852 (N_9852,N_9173,N_9402);
and U9853 (N_9853,N_9160,N_9205);
nand U9854 (N_9854,N_9285,N_9174);
or U9855 (N_9855,N_9163,N_9023);
xor U9856 (N_9856,N_9408,N_9274);
or U9857 (N_9857,N_9223,N_9120);
nor U9858 (N_9858,N_9296,N_9375);
nand U9859 (N_9859,N_9134,N_9380);
and U9860 (N_9860,N_9222,N_9291);
nand U9861 (N_9861,N_9234,N_9403);
nor U9862 (N_9862,N_9468,N_9108);
and U9863 (N_9863,N_9416,N_9498);
nand U9864 (N_9864,N_9211,N_9268);
or U9865 (N_9865,N_9054,N_9455);
nand U9866 (N_9866,N_9131,N_9197);
nor U9867 (N_9867,N_9002,N_9446);
nand U9868 (N_9868,N_9400,N_9003);
nand U9869 (N_9869,N_9038,N_9209);
nand U9870 (N_9870,N_9209,N_9402);
nor U9871 (N_9871,N_9445,N_9451);
nand U9872 (N_9872,N_9411,N_9109);
nand U9873 (N_9873,N_9267,N_9198);
nor U9874 (N_9874,N_9472,N_9328);
nand U9875 (N_9875,N_9060,N_9196);
nor U9876 (N_9876,N_9420,N_9169);
or U9877 (N_9877,N_9014,N_9230);
nand U9878 (N_9878,N_9016,N_9400);
nand U9879 (N_9879,N_9197,N_9145);
or U9880 (N_9880,N_9396,N_9301);
nand U9881 (N_9881,N_9375,N_9130);
xnor U9882 (N_9882,N_9285,N_9128);
or U9883 (N_9883,N_9133,N_9243);
nor U9884 (N_9884,N_9435,N_9147);
nand U9885 (N_9885,N_9341,N_9112);
or U9886 (N_9886,N_9403,N_9266);
nor U9887 (N_9887,N_9141,N_9281);
or U9888 (N_9888,N_9408,N_9153);
nor U9889 (N_9889,N_9464,N_9273);
nand U9890 (N_9890,N_9286,N_9361);
nor U9891 (N_9891,N_9016,N_9329);
or U9892 (N_9892,N_9228,N_9104);
nand U9893 (N_9893,N_9306,N_9221);
and U9894 (N_9894,N_9178,N_9298);
or U9895 (N_9895,N_9409,N_9097);
nor U9896 (N_9896,N_9484,N_9108);
or U9897 (N_9897,N_9449,N_9302);
nor U9898 (N_9898,N_9042,N_9479);
nor U9899 (N_9899,N_9434,N_9450);
nand U9900 (N_9900,N_9213,N_9479);
nand U9901 (N_9901,N_9298,N_9496);
xnor U9902 (N_9902,N_9128,N_9173);
or U9903 (N_9903,N_9347,N_9187);
nor U9904 (N_9904,N_9052,N_9001);
or U9905 (N_9905,N_9466,N_9149);
nand U9906 (N_9906,N_9212,N_9341);
or U9907 (N_9907,N_9466,N_9229);
and U9908 (N_9908,N_9151,N_9332);
and U9909 (N_9909,N_9344,N_9069);
or U9910 (N_9910,N_9234,N_9094);
nor U9911 (N_9911,N_9365,N_9138);
or U9912 (N_9912,N_9014,N_9431);
or U9913 (N_9913,N_9229,N_9422);
and U9914 (N_9914,N_9437,N_9486);
nor U9915 (N_9915,N_9365,N_9206);
and U9916 (N_9916,N_9266,N_9227);
or U9917 (N_9917,N_9457,N_9420);
and U9918 (N_9918,N_9125,N_9380);
nand U9919 (N_9919,N_9216,N_9277);
nor U9920 (N_9920,N_9078,N_9155);
and U9921 (N_9921,N_9002,N_9357);
or U9922 (N_9922,N_9471,N_9478);
or U9923 (N_9923,N_9383,N_9092);
nand U9924 (N_9924,N_9006,N_9129);
or U9925 (N_9925,N_9058,N_9271);
or U9926 (N_9926,N_9459,N_9187);
nand U9927 (N_9927,N_9168,N_9147);
nand U9928 (N_9928,N_9444,N_9203);
or U9929 (N_9929,N_9041,N_9456);
and U9930 (N_9930,N_9007,N_9138);
nor U9931 (N_9931,N_9388,N_9309);
or U9932 (N_9932,N_9205,N_9015);
nand U9933 (N_9933,N_9462,N_9468);
or U9934 (N_9934,N_9071,N_9009);
nor U9935 (N_9935,N_9162,N_9484);
nand U9936 (N_9936,N_9283,N_9058);
nand U9937 (N_9937,N_9261,N_9344);
nor U9938 (N_9938,N_9255,N_9205);
or U9939 (N_9939,N_9224,N_9491);
nand U9940 (N_9940,N_9082,N_9026);
nor U9941 (N_9941,N_9335,N_9487);
nand U9942 (N_9942,N_9352,N_9051);
nand U9943 (N_9943,N_9063,N_9065);
nand U9944 (N_9944,N_9179,N_9460);
nor U9945 (N_9945,N_9107,N_9305);
nand U9946 (N_9946,N_9271,N_9255);
and U9947 (N_9947,N_9399,N_9220);
nor U9948 (N_9948,N_9254,N_9223);
and U9949 (N_9949,N_9366,N_9035);
nor U9950 (N_9950,N_9068,N_9490);
or U9951 (N_9951,N_9212,N_9435);
or U9952 (N_9952,N_9477,N_9409);
xnor U9953 (N_9953,N_9260,N_9309);
nor U9954 (N_9954,N_9173,N_9063);
nor U9955 (N_9955,N_9122,N_9269);
xor U9956 (N_9956,N_9069,N_9161);
nand U9957 (N_9957,N_9363,N_9013);
and U9958 (N_9958,N_9235,N_9147);
or U9959 (N_9959,N_9022,N_9000);
or U9960 (N_9960,N_9409,N_9349);
or U9961 (N_9961,N_9457,N_9350);
nand U9962 (N_9962,N_9167,N_9460);
or U9963 (N_9963,N_9198,N_9356);
or U9964 (N_9964,N_9443,N_9285);
and U9965 (N_9965,N_9422,N_9002);
nand U9966 (N_9966,N_9458,N_9209);
nor U9967 (N_9967,N_9134,N_9429);
or U9968 (N_9968,N_9240,N_9426);
and U9969 (N_9969,N_9306,N_9005);
nor U9970 (N_9970,N_9242,N_9090);
nand U9971 (N_9971,N_9387,N_9435);
or U9972 (N_9972,N_9239,N_9301);
nand U9973 (N_9973,N_9013,N_9125);
and U9974 (N_9974,N_9037,N_9320);
or U9975 (N_9975,N_9218,N_9030);
and U9976 (N_9976,N_9001,N_9409);
nor U9977 (N_9977,N_9123,N_9303);
or U9978 (N_9978,N_9314,N_9082);
and U9979 (N_9979,N_9248,N_9416);
or U9980 (N_9980,N_9090,N_9305);
nor U9981 (N_9981,N_9281,N_9487);
nor U9982 (N_9982,N_9060,N_9341);
nor U9983 (N_9983,N_9162,N_9111);
or U9984 (N_9984,N_9070,N_9204);
nor U9985 (N_9985,N_9441,N_9028);
nor U9986 (N_9986,N_9039,N_9189);
nor U9987 (N_9987,N_9062,N_9445);
nand U9988 (N_9988,N_9119,N_9299);
nand U9989 (N_9989,N_9454,N_9387);
nand U9990 (N_9990,N_9155,N_9137);
or U9991 (N_9991,N_9149,N_9380);
xnor U9992 (N_9992,N_9328,N_9047);
and U9993 (N_9993,N_9073,N_9297);
or U9994 (N_9994,N_9452,N_9012);
xnor U9995 (N_9995,N_9350,N_9311);
nor U9996 (N_9996,N_9358,N_9237);
or U9997 (N_9997,N_9440,N_9214);
and U9998 (N_9998,N_9041,N_9230);
nor U9999 (N_9999,N_9413,N_9345);
nand UO_0 (O_0,N_9778,N_9860);
or UO_1 (O_1,N_9582,N_9996);
nand UO_2 (O_2,N_9522,N_9746);
nor UO_3 (O_3,N_9580,N_9764);
or UO_4 (O_4,N_9867,N_9788);
or UO_5 (O_5,N_9562,N_9804);
and UO_6 (O_6,N_9636,N_9849);
and UO_7 (O_7,N_9674,N_9631);
or UO_8 (O_8,N_9870,N_9981);
nor UO_9 (O_9,N_9808,N_9779);
and UO_10 (O_10,N_9713,N_9783);
nor UO_11 (O_11,N_9814,N_9898);
or UO_12 (O_12,N_9581,N_9982);
nor UO_13 (O_13,N_9977,N_9663);
nor UO_14 (O_14,N_9927,N_9610);
or UO_15 (O_15,N_9979,N_9551);
or UO_16 (O_16,N_9645,N_9865);
or UO_17 (O_17,N_9875,N_9703);
and UO_18 (O_18,N_9584,N_9708);
nand UO_19 (O_19,N_9727,N_9920);
and UO_20 (O_20,N_9847,N_9595);
nor UO_21 (O_21,N_9940,N_9975);
or UO_22 (O_22,N_9662,N_9993);
or UO_23 (O_23,N_9791,N_9838);
nor UO_24 (O_24,N_9845,N_9655);
or UO_25 (O_25,N_9650,N_9987);
nor UO_26 (O_26,N_9682,N_9776);
or UO_27 (O_27,N_9629,N_9574);
and UO_28 (O_28,N_9583,N_9864);
nand UO_29 (O_29,N_9770,N_9564);
and UO_30 (O_30,N_9895,N_9863);
nor UO_31 (O_31,N_9908,N_9614);
and UO_32 (O_32,N_9578,N_9911);
or UO_33 (O_33,N_9876,N_9789);
and UO_34 (O_34,N_9586,N_9974);
nor UO_35 (O_35,N_9724,N_9843);
nand UO_36 (O_36,N_9677,N_9577);
nor UO_37 (O_37,N_9740,N_9762);
and UO_38 (O_38,N_9566,N_9968);
nor UO_39 (O_39,N_9602,N_9837);
nor UO_40 (O_40,N_9589,N_9971);
or UO_41 (O_41,N_9914,N_9731);
nor UO_42 (O_42,N_9687,N_9633);
nor UO_43 (O_43,N_9561,N_9873);
and UO_44 (O_44,N_9763,N_9518);
nand UO_45 (O_45,N_9997,N_9649);
nor UO_46 (O_46,N_9548,N_9652);
nand UO_47 (O_47,N_9509,N_9596);
or UO_48 (O_48,N_9954,N_9739);
or UO_49 (O_49,N_9533,N_9866);
or UO_50 (O_50,N_9805,N_9760);
nand UO_51 (O_51,N_9976,N_9790);
nor UO_52 (O_52,N_9513,N_9918);
and UO_53 (O_53,N_9820,N_9716);
and UO_54 (O_54,N_9872,N_9736);
and UO_55 (O_55,N_9786,N_9528);
or UO_56 (O_56,N_9912,N_9666);
xnor UO_57 (O_57,N_9698,N_9671);
and UO_58 (O_58,N_9714,N_9903);
or UO_59 (O_59,N_9989,N_9693);
nand UO_60 (O_60,N_9951,N_9516);
nand UO_61 (O_61,N_9759,N_9742);
or UO_62 (O_62,N_9905,N_9973);
and UO_63 (O_63,N_9619,N_9505);
and UO_64 (O_64,N_9824,N_9777);
and UO_65 (O_65,N_9750,N_9544);
nor UO_66 (O_66,N_9709,N_9882);
or UO_67 (O_67,N_9868,N_9711);
or UO_68 (O_68,N_9521,N_9816);
or UO_69 (O_69,N_9801,N_9780);
or UO_70 (O_70,N_9621,N_9542);
or UO_71 (O_71,N_9678,N_9541);
and UO_72 (O_72,N_9956,N_9807);
nand UO_73 (O_73,N_9710,N_9720);
or UO_74 (O_74,N_9980,N_9902);
nor UO_75 (O_75,N_9794,N_9952);
and UO_76 (O_76,N_9827,N_9565);
nand UO_77 (O_77,N_9923,N_9921);
and UO_78 (O_78,N_9726,N_9963);
and UO_79 (O_79,N_9901,N_9692);
nor UO_80 (O_80,N_9928,N_9628);
and UO_81 (O_81,N_9833,N_9948);
or UO_82 (O_82,N_9506,N_9514);
or UO_83 (O_83,N_9925,N_9620);
or UO_84 (O_84,N_9959,N_9657);
and UO_85 (O_85,N_9571,N_9815);
and UO_86 (O_86,N_9665,N_9729);
nor UO_87 (O_87,N_9758,N_9861);
and UO_88 (O_88,N_9730,N_9653);
and UO_89 (O_89,N_9785,N_9524);
or UO_90 (O_90,N_9719,N_9737);
nand UO_91 (O_91,N_9941,N_9936);
nor UO_92 (O_92,N_9638,N_9688);
or UO_93 (O_93,N_9747,N_9855);
or UO_94 (O_94,N_9879,N_9915);
and UO_95 (O_95,N_9717,N_9884);
nand UO_96 (O_96,N_9543,N_9897);
and UO_97 (O_97,N_9673,N_9818);
nor UO_98 (O_98,N_9825,N_9691);
or UO_99 (O_99,N_9643,N_9696);
nor UO_100 (O_100,N_9699,N_9797);
nor UO_101 (O_101,N_9569,N_9632);
and UO_102 (O_102,N_9906,N_9819);
or UO_103 (O_103,N_9723,N_9994);
and UO_104 (O_104,N_9817,N_9961);
and UO_105 (O_105,N_9531,N_9627);
nor UO_106 (O_106,N_9811,N_9637);
nand UO_107 (O_107,N_9686,N_9896);
nor UO_108 (O_108,N_9555,N_9715);
or UO_109 (O_109,N_9587,N_9608);
nand UO_110 (O_110,N_9784,N_9641);
nor UO_111 (O_111,N_9556,N_9676);
or UO_112 (O_112,N_9613,N_9831);
nand UO_113 (O_113,N_9766,N_9839);
or UO_114 (O_114,N_9768,N_9782);
or UO_115 (O_115,N_9851,N_9751);
and UO_116 (O_116,N_9557,N_9532);
or UO_117 (O_117,N_9943,N_9697);
or UO_118 (O_118,N_9950,N_9878);
nand UO_119 (O_119,N_9567,N_9651);
or UO_120 (O_120,N_9536,N_9597);
and UO_121 (O_121,N_9683,N_9519);
nand UO_122 (O_122,N_9721,N_9656);
and UO_123 (O_123,N_9738,N_9933);
and UO_124 (O_124,N_9880,N_9771);
nor UO_125 (O_125,N_9741,N_9892);
nand UO_126 (O_126,N_9605,N_9835);
and UO_127 (O_127,N_9874,N_9559);
nor UO_128 (O_128,N_9648,N_9848);
or UO_129 (O_129,N_9917,N_9732);
or UO_130 (O_130,N_9856,N_9995);
nor UO_131 (O_131,N_9972,N_9558);
and UO_132 (O_132,N_9909,N_9773);
or UO_133 (O_133,N_9886,N_9850);
and UO_134 (O_134,N_9826,N_9796);
or UO_135 (O_135,N_9667,N_9588);
nor UO_136 (O_136,N_9871,N_9767);
or UO_137 (O_137,N_9593,N_9953);
nor UO_138 (O_138,N_9931,N_9834);
or UO_139 (O_139,N_9803,N_9579);
and UO_140 (O_140,N_9822,N_9769);
nand UO_141 (O_141,N_9765,N_9828);
and UO_142 (O_142,N_9842,N_9735);
xnor UO_143 (O_143,N_9781,N_9992);
nand UO_144 (O_144,N_9609,N_9603);
or UO_145 (O_145,N_9590,N_9965);
nor UO_146 (O_146,N_9660,N_9836);
nor UO_147 (O_147,N_9700,N_9949);
or UO_148 (O_148,N_9707,N_9932);
or UO_149 (O_149,N_9757,N_9946);
nand UO_150 (O_150,N_9670,N_9535);
and UO_151 (O_151,N_9907,N_9685);
and UO_152 (O_152,N_9576,N_9575);
nor UO_153 (O_153,N_9787,N_9545);
nor UO_154 (O_154,N_9538,N_9572);
xnor UO_155 (O_155,N_9598,N_9681);
xnor UO_156 (O_156,N_9958,N_9922);
and UO_157 (O_157,N_9552,N_9560);
nand UO_158 (O_158,N_9844,N_9623);
nand UO_159 (O_159,N_9664,N_9942);
nor UO_160 (O_160,N_9625,N_9859);
and UO_161 (O_161,N_9793,N_9890);
or UO_162 (O_162,N_9969,N_9606);
nand UO_163 (O_163,N_9617,N_9527);
and UO_164 (O_164,N_9702,N_9858);
nor UO_165 (O_165,N_9540,N_9743);
nand UO_166 (O_166,N_9728,N_9599);
nor UO_167 (O_167,N_9924,N_9978);
nor UO_168 (O_168,N_9600,N_9744);
nand UO_169 (O_169,N_9615,N_9935);
xor UO_170 (O_170,N_9661,N_9887);
nor UO_171 (O_171,N_9601,N_9930);
nand UO_172 (O_172,N_9675,N_9704);
and UO_173 (O_173,N_9694,N_9510);
and UO_174 (O_174,N_9523,N_9534);
or UO_175 (O_175,N_9689,N_9998);
nand UO_176 (O_176,N_9550,N_9984);
nand UO_177 (O_177,N_9611,N_9517);
nand UO_178 (O_178,N_9883,N_9756);
nor UO_179 (O_179,N_9926,N_9985);
and UO_180 (O_180,N_9955,N_9646);
or UO_181 (O_181,N_9624,N_9734);
or UO_182 (O_182,N_9592,N_9829);
nor UO_183 (O_183,N_9669,N_9983);
or UO_184 (O_184,N_9899,N_9604);
xnor UO_185 (O_185,N_9916,N_9841);
or UO_186 (O_186,N_9919,N_9626);
and UO_187 (O_187,N_9647,N_9622);
or UO_188 (O_188,N_9634,N_9888);
nand UO_189 (O_189,N_9795,N_9701);
nor UO_190 (O_190,N_9725,N_9680);
and UO_191 (O_191,N_9549,N_9511);
and UO_192 (O_192,N_9640,N_9846);
nor UO_193 (O_193,N_9722,N_9806);
and UO_194 (O_194,N_9754,N_9900);
and UO_195 (O_195,N_9658,N_9752);
nor UO_196 (O_196,N_9853,N_9947);
nor UO_197 (O_197,N_9684,N_9672);
nor UO_198 (O_198,N_9991,N_9644);
nor UO_199 (O_199,N_9999,N_9934);
and UO_200 (O_200,N_9547,N_9712);
nand UO_201 (O_201,N_9563,N_9945);
nand UO_202 (O_202,N_9986,N_9862);
nand UO_203 (O_203,N_9799,N_9990);
nor UO_204 (O_204,N_9594,N_9706);
xnor UO_205 (O_205,N_9966,N_9939);
and UO_206 (O_206,N_9618,N_9570);
and UO_207 (O_207,N_9537,N_9668);
nand UO_208 (O_208,N_9967,N_9554);
nor UO_209 (O_209,N_9830,N_9970);
nand UO_210 (O_210,N_9772,N_9512);
or UO_211 (O_211,N_9659,N_9755);
and UO_212 (O_212,N_9840,N_9573);
or UO_213 (O_213,N_9508,N_9893);
and UO_214 (O_214,N_9809,N_9526);
and UO_215 (O_215,N_9904,N_9775);
or UO_216 (O_216,N_9635,N_9501);
and UO_217 (O_217,N_9823,N_9503);
and UO_218 (O_218,N_9962,N_9642);
nor UO_219 (O_219,N_9733,N_9500);
and UO_220 (O_220,N_9869,N_9553);
or UO_221 (O_221,N_9695,N_9894);
nand UO_222 (O_222,N_9529,N_9891);
nor UO_223 (O_223,N_9539,N_9913);
nor UO_224 (O_224,N_9938,N_9679);
nor UO_225 (O_225,N_9802,N_9964);
nor UO_226 (O_226,N_9585,N_9929);
nor UO_227 (O_227,N_9530,N_9612);
or UO_228 (O_228,N_9718,N_9944);
and UO_229 (O_229,N_9854,N_9813);
and UO_230 (O_230,N_9568,N_9591);
nor UO_231 (O_231,N_9988,N_9748);
and UO_232 (O_232,N_9937,N_9877);
and UO_233 (O_233,N_9852,N_9821);
nor UO_234 (O_234,N_9798,N_9630);
nand UO_235 (O_235,N_9810,N_9515);
nor UO_236 (O_236,N_9881,N_9857);
nor UO_237 (O_237,N_9753,N_9800);
nand UO_238 (O_238,N_9607,N_9792);
or UO_239 (O_239,N_9885,N_9690);
and UO_240 (O_240,N_9502,N_9749);
or UO_241 (O_241,N_9774,N_9960);
and UO_242 (O_242,N_9832,N_9546);
and UO_243 (O_243,N_9889,N_9654);
and UO_244 (O_244,N_9507,N_9616);
or UO_245 (O_245,N_9812,N_9520);
nor UO_246 (O_246,N_9639,N_9705);
nand UO_247 (O_247,N_9761,N_9957);
nor UO_248 (O_248,N_9910,N_9504);
nand UO_249 (O_249,N_9525,N_9745);
xnor UO_250 (O_250,N_9631,N_9945);
and UO_251 (O_251,N_9692,N_9765);
nor UO_252 (O_252,N_9993,N_9561);
and UO_253 (O_253,N_9558,N_9881);
and UO_254 (O_254,N_9944,N_9526);
nor UO_255 (O_255,N_9867,N_9786);
nand UO_256 (O_256,N_9677,N_9761);
or UO_257 (O_257,N_9895,N_9515);
nor UO_258 (O_258,N_9681,N_9893);
nor UO_259 (O_259,N_9829,N_9812);
or UO_260 (O_260,N_9997,N_9523);
nand UO_261 (O_261,N_9634,N_9543);
nand UO_262 (O_262,N_9808,N_9580);
nand UO_263 (O_263,N_9924,N_9799);
nand UO_264 (O_264,N_9716,N_9527);
and UO_265 (O_265,N_9837,N_9802);
xnor UO_266 (O_266,N_9874,N_9919);
xnor UO_267 (O_267,N_9628,N_9621);
nor UO_268 (O_268,N_9768,N_9776);
nor UO_269 (O_269,N_9848,N_9940);
or UO_270 (O_270,N_9567,N_9873);
or UO_271 (O_271,N_9819,N_9920);
nor UO_272 (O_272,N_9790,N_9641);
and UO_273 (O_273,N_9799,N_9928);
nand UO_274 (O_274,N_9788,N_9888);
nor UO_275 (O_275,N_9790,N_9918);
and UO_276 (O_276,N_9597,N_9545);
or UO_277 (O_277,N_9779,N_9885);
nor UO_278 (O_278,N_9575,N_9620);
nor UO_279 (O_279,N_9982,N_9920);
nand UO_280 (O_280,N_9994,N_9998);
nor UO_281 (O_281,N_9919,N_9902);
nor UO_282 (O_282,N_9630,N_9889);
and UO_283 (O_283,N_9720,N_9834);
nand UO_284 (O_284,N_9650,N_9571);
nand UO_285 (O_285,N_9652,N_9898);
nor UO_286 (O_286,N_9998,N_9852);
or UO_287 (O_287,N_9897,N_9668);
nor UO_288 (O_288,N_9863,N_9534);
and UO_289 (O_289,N_9583,N_9717);
or UO_290 (O_290,N_9527,N_9644);
nor UO_291 (O_291,N_9879,N_9531);
or UO_292 (O_292,N_9968,N_9765);
xnor UO_293 (O_293,N_9528,N_9568);
and UO_294 (O_294,N_9753,N_9600);
or UO_295 (O_295,N_9600,N_9819);
and UO_296 (O_296,N_9663,N_9789);
nand UO_297 (O_297,N_9688,N_9899);
nand UO_298 (O_298,N_9606,N_9929);
nor UO_299 (O_299,N_9658,N_9919);
nand UO_300 (O_300,N_9651,N_9656);
nor UO_301 (O_301,N_9943,N_9634);
nor UO_302 (O_302,N_9628,N_9812);
or UO_303 (O_303,N_9871,N_9583);
or UO_304 (O_304,N_9646,N_9712);
nand UO_305 (O_305,N_9637,N_9914);
or UO_306 (O_306,N_9697,N_9599);
nand UO_307 (O_307,N_9760,N_9563);
or UO_308 (O_308,N_9507,N_9735);
and UO_309 (O_309,N_9612,N_9742);
nand UO_310 (O_310,N_9957,N_9796);
nand UO_311 (O_311,N_9585,N_9919);
nor UO_312 (O_312,N_9990,N_9674);
nand UO_313 (O_313,N_9904,N_9743);
and UO_314 (O_314,N_9631,N_9827);
or UO_315 (O_315,N_9714,N_9524);
nand UO_316 (O_316,N_9649,N_9903);
nand UO_317 (O_317,N_9873,N_9885);
or UO_318 (O_318,N_9569,N_9717);
and UO_319 (O_319,N_9932,N_9770);
or UO_320 (O_320,N_9885,N_9808);
nand UO_321 (O_321,N_9677,N_9810);
or UO_322 (O_322,N_9671,N_9591);
and UO_323 (O_323,N_9559,N_9756);
nand UO_324 (O_324,N_9668,N_9921);
or UO_325 (O_325,N_9548,N_9800);
nor UO_326 (O_326,N_9698,N_9918);
nor UO_327 (O_327,N_9905,N_9963);
nand UO_328 (O_328,N_9800,N_9871);
or UO_329 (O_329,N_9877,N_9795);
or UO_330 (O_330,N_9717,N_9518);
or UO_331 (O_331,N_9654,N_9752);
nand UO_332 (O_332,N_9933,N_9971);
nand UO_333 (O_333,N_9892,N_9607);
nand UO_334 (O_334,N_9992,N_9871);
nor UO_335 (O_335,N_9702,N_9751);
or UO_336 (O_336,N_9696,N_9927);
nor UO_337 (O_337,N_9926,N_9776);
or UO_338 (O_338,N_9824,N_9662);
nor UO_339 (O_339,N_9578,N_9765);
or UO_340 (O_340,N_9831,N_9808);
or UO_341 (O_341,N_9857,N_9621);
nand UO_342 (O_342,N_9528,N_9565);
and UO_343 (O_343,N_9541,N_9942);
or UO_344 (O_344,N_9516,N_9897);
and UO_345 (O_345,N_9981,N_9899);
and UO_346 (O_346,N_9654,N_9609);
nand UO_347 (O_347,N_9530,N_9778);
nand UO_348 (O_348,N_9791,N_9557);
and UO_349 (O_349,N_9711,N_9565);
and UO_350 (O_350,N_9850,N_9732);
nor UO_351 (O_351,N_9960,N_9919);
or UO_352 (O_352,N_9597,N_9576);
nor UO_353 (O_353,N_9589,N_9595);
and UO_354 (O_354,N_9654,N_9993);
or UO_355 (O_355,N_9801,N_9640);
nand UO_356 (O_356,N_9844,N_9831);
and UO_357 (O_357,N_9901,N_9783);
nand UO_358 (O_358,N_9788,N_9989);
nor UO_359 (O_359,N_9592,N_9542);
or UO_360 (O_360,N_9621,N_9915);
nor UO_361 (O_361,N_9601,N_9899);
nand UO_362 (O_362,N_9809,N_9777);
nand UO_363 (O_363,N_9501,N_9590);
or UO_364 (O_364,N_9799,N_9593);
and UO_365 (O_365,N_9660,N_9672);
and UO_366 (O_366,N_9700,N_9511);
or UO_367 (O_367,N_9807,N_9706);
or UO_368 (O_368,N_9935,N_9763);
nand UO_369 (O_369,N_9617,N_9514);
nand UO_370 (O_370,N_9863,N_9828);
nand UO_371 (O_371,N_9886,N_9685);
nor UO_372 (O_372,N_9910,N_9963);
nor UO_373 (O_373,N_9846,N_9916);
or UO_374 (O_374,N_9942,N_9728);
and UO_375 (O_375,N_9707,N_9988);
nor UO_376 (O_376,N_9962,N_9807);
or UO_377 (O_377,N_9831,N_9829);
and UO_378 (O_378,N_9533,N_9752);
nor UO_379 (O_379,N_9958,N_9583);
nand UO_380 (O_380,N_9694,N_9631);
nor UO_381 (O_381,N_9635,N_9965);
and UO_382 (O_382,N_9623,N_9610);
or UO_383 (O_383,N_9966,N_9918);
nor UO_384 (O_384,N_9779,N_9985);
and UO_385 (O_385,N_9877,N_9575);
nand UO_386 (O_386,N_9918,N_9991);
and UO_387 (O_387,N_9934,N_9507);
or UO_388 (O_388,N_9992,N_9941);
and UO_389 (O_389,N_9973,N_9641);
nor UO_390 (O_390,N_9537,N_9809);
xnor UO_391 (O_391,N_9562,N_9731);
or UO_392 (O_392,N_9625,N_9614);
nand UO_393 (O_393,N_9582,N_9680);
or UO_394 (O_394,N_9515,N_9743);
or UO_395 (O_395,N_9581,N_9754);
and UO_396 (O_396,N_9528,N_9843);
or UO_397 (O_397,N_9669,N_9849);
nand UO_398 (O_398,N_9830,N_9566);
or UO_399 (O_399,N_9909,N_9795);
or UO_400 (O_400,N_9813,N_9740);
and UO_401 (O_401,N_9986,N_9824);
nor UO_402 (O_402,N_9743,N_9684);
or UO_403 (O_403,N_9731,N_9679);
and UO_404 (O_404,N_9743,N_9840);
nand UO_405 (O_405,N_9988,N_9612);
nor UO_406 (O_406,N_9500,N_9644);
nor UO_407 (O_407,N_9575,N_9536);
nand UO_408 (O_408,N_9973,N_9543);
nor UO_409 (O_409,N_9700,N_9802);
xor UO_410 (O_410,N_9891,N_9840);
and UO_411 (O_411,N_9994,N_9798);
or UO_412 (O_412,N_9570,N_9590);
or UO_413 (O_413,N_9737,N_9554);
or UO_414 (O_414,N_9573,N_9597);
or UO_415 (O_415,N_9853,N_9944);
nor UO_416 (O_416,N_9828,N_9978);
nor UO_417 (O_417,N_9758,N_9970);
or UO_418 (O_418,N_9804,N_9629);
and UO_419 (O_419,N_9543,N_9903);
or UO_420 (O_420,N_9895,N_9707);
nand UO_421 (O_421,N_9915,N_9726);
and UO_422 (O_422,N_9684,N_9903);
nor UO_423 (O_423,N_9756,N_9609);
nor UO_424 (O_424,N_9606,N_9932);
or UO_425 (O_425,N_9622,N_9796);
nand UO_426 (O_426,N_9729,N_9935);
and UO_427 (O_427,N_9983,N_9500);
and UO_428 (O_428,N_9548,N_9799);
or UO_429 (O_429,N_9944,N_9726);
and UO_430 (O_430,N_9814,N_9741);
nor UO_431 (O_431,N_9632,N_9930);
nor UO_432 (O_432,N_9767,N_9759);
and UO_433 (O_433,N_9762,N_9712);
xor UO_434 (O_434,N_9646,N_9666);
nor UO_435 (O_435,N_9719,N_9545);
or UO_436 (O_436,N_9644,N_9836);
xor UO_437 (O_437,N_9553,N_9529);
nor UO_438 (O_438,N_9659,N_9739);
and UO_439 (O_439,N_9555,N_9503);
nand UO_440 (O_440,N_9607,N_9899);
and UO_441 (O_441,N_9956,N_9563);
nor UO_442 (O_442,N_9960,N_9595);
and UO_443 (O_443,N_9667,N_9992);
nor UO_444 (O_444,N_9617,N_9735);
or UO_445 (O_445,N_9643,N_9644);
and UO_446 (O_446,N_9646,N_9815);
or UO_447 (O_447,N_9760,N_9782);
and UO_448 (O_448,N_9521,N_9877);
and UO_449 (O_449,N_9785,N_9897);
and UO_450 (O_450,N_9695,N_9978);
or UO_451 (O_451,N_9516,N_9641);
or UO_452 (O_452,N_9847,N_9625);
or UO_453 (O_453,N_9644,N_9609);
nor UO_454 (O_454,N_9914,N_9811);
and UO_455 (O_455,N_9902,N_9527);
and UO_456 (O_456,N_9616,N_9728);
nand UO_457 (O_457,N_9529,N_9551);
or UO_458 (O_458,N_9512,N_9844);
nand UO_459 (O_459,N_9875,N_9583);
or UO_460 (O_460,N_9857,N_9576);
or UO_461 (O_461,N_9518,N_9653);
and UO_462 (O_462,N_9660,N_9776);
or UO_463 (O_463,N_9821,N_9702);
nor UO_464 (O_464,N_9970,N_9912);
nand UO_465 (O_465,N_9804,N_9995);
nand UO_466 (O_466,N_9898,N_9659);
nor UO_467 (O_467,N_9830,N_9773);
nor UO_468 (O_468,N_9534,N_9869);
and UO_469 (O_469,N_9635,N_9801);
nand UO_470 (O_470,N_9698,N_9894);
nand UO_471 (O_471,N_9599,N_9802);
nand UO_472 (O_472,N_9871,N_9512);
and UO_473 (O_473,N_9771,N_9562);
nand UO_474 (O_474,N_9725,N_9909);
nand UO_475 (O_475,N_9899,N_9599);
and UO_476 (O_476,N_9703,N_9755);
nor UO_477 (O_477,N_9912,N_9793);
nand UO_478 (O_478,N_9919,N_9853);
nor UO_479 (O_479,N_9976,N_9524);
or UO_480 (O_480,N_9623,N_9516);
nor UO_481 (O_481,N_9601,N_9922);
nor UO_482 (O_482,N_9988,N_9657);
nand UO_483 (O_483,N_9794,N_9698);
or UO_484 (O_484,N_9960,N_9540);
and UO_485 (O_485,N_9778,N_9993);
nor UO_486 (O_486,N_9840,N_9953);
nand UO_487 (O_487,N_9974,N_9568);
nand UO_488 (O_488,N_9601,N_9595);
or UO_489 (O_489,N_9758,N_9713);
nand UO_490 (O_490,N_9561,N_9617);
and UO_491 (O_491,N_9691,N_9530);
nand UO_492 (O_492,N_9543,N_9947);
nor UO_493 (O_493,N_9590,N_9822);
or UO_494 (O_494,N_9894,N_9534);
nor UO_495 (O_495,N_9849,N_9692);
nand UO_496 (O_496,N_9507,N_9823);
and UO_497 (O_497,N_9706,N_9841);
and UO_498 (O_498,N_9529,N_9851);
nand UO_499 (O_499,N_9762,N_9643);
and UO_500 (O_500,N_9886,N_9557);
nor UO_501 (O_501,N_9661,N_9602);
and UO_502 (O_502,N_9844,N_9892);
and UO_503 (O_503,N_9748,N_9608);
and UO_504 (O_504,N_9772,N_9983);
xnor UO_505 (O_505,N_9595,N_9796);
and UO_506 (O_506,N_9645,N_9953);
nor UO_507 (O_507,N_9734,N_9716);
and UO_508 (O_508,N_9509,N_9941);
nor UO_509 (O_509,N_9565,N_9622);
or UO_510 (O_510,N_9642,N_9779);
or UO_511 (O_511,N_9619,N_9604);
and UO_512 (O_512,N_9518,N_9738);
nand UO_513 (O_513,N_9732,N_9787);
and UO_514 (O_514,N_9555,N_9737);
and UO_515 (O_515,N_9714,N_9844);
nor UO_516 (O_516,N_9912,N_9925);
and UO_517 (O_517,N_9942,N_9946);
and UO_518 (O_518,N_9959,N_9779);
nor UO_519 (O_519,N_9772,N_9778);
nand UO_520 (O_520,N_9941,N_9837);
nor UO_521 (O_521,N_9972,N_9836);
or UO_522 (O_522,N_9547,N_9646);
nand UO_523 (O_523,N_9944,N_9597);
nor UO_524 (O_524,N_9820,N_9707);
and UO_525 (O_525,N_9625,N_9722);
or UO_526 (O_526,N_9707,N_9734);
and UO_527 (O_527,N_9807,N_9500);
nor UO_528 (O_528,N_9736,N_9758);
or UO_529 (O_529,N_9835,N_9593);
or UO_530 (O_530,N_9809,N_9503);
nor UO_531 (O_531,N_9631,N_9543);
or UO_532 (O_532,N_9540,N_9708);
nor UO_533 (O_533,N_9599,N_9849);
nor UO_534 (O_534,N_9922,N_9884);
nor UO_535 (O_535,N_9954,N_9946);
and UO_536 (O_536,N_9885,N_9544);
nand UO_537 (O_537,N_9651,N_9591);
nor UO_538 (O_538,N_9568,N_9959);
and UO_539 (O_539,N_9537,N_9787);
nand UO_540 (O_540,N_9923,N_9521);
or UO_541 (O_541,N_9523,N_9598);
nor UO_542 (O_542,N_9815,N_9955);
nand UO_543 (O_543,N_9965,N_9510);
nand UO_544 (O_544,N_9830,N_9760);
xor UO_545 (O_545,N_9751,N_9503);
nor UO_546 (O_546,N_9555,N_9606);
and UO_547 (O_547,N_9743,N_9770);
nand UO_548 (O_548,N_9568,N_9744);
or UO_549 (O_549,N_9615,N_9769);
nand UO_550 (O_550,N_9680,N_9942);
and UO_551 (O_551,N_9617,N_9535);
nor UO_552 (O_552,N_9794,N_9685);
and UO_553 (O_553,N_9501,N_9869);
nor UO_554 (O_554,N_9875,N_9945);
and UO_555 (O_555,N_9670,N_9920);
or UO_556 (O_556,N_9916,N_9631);
nor UO_557 (O_557,N_9701,N_9773);
nand UO_558 (O_558,N_9589,N_9869);
nor UO_559 (O_559,N_9547,N_9997);
and UO_560 (O_560,N_9845,N_9887);
nand UO_561 (O_561,N_9827,N_9552);
or UO_562 (O_562,N_9864,N_9681);
and UO_563 (O_563,N_9527,N_9983);
nor UO_564 (O_564,N_9732,N_9884);
or UO_565 (O_565,N_9895,N_9872);
and UO_566 (O_566,N_9680,N_9803);
or UO_567 (O_567,N_9934,N_9627);
nand UO_568 (O_568,N_9932,N_9754);
nor UO_569 (O_569,N_9687,N_9745);
nor UO_570 (O_570,N_9872,N_9909);
or UO_571 (O_571,N_9645,N_9599);
and UO_572 (O_572,N_9924,N_9632);
or UO_573 (O_573,N_9577,N_9607);
nand UO_574 (O_574,N_9626,N_9644);
nand UO_575 (O_575,N_9920,N_9915);
nor UO_576 (O_576,N_9807,N_9715);
nand UO_577 (O_577,N_9500,N_9954);
nor UO_578 (O_578,N_9727,N_9587);
nand UO_579 (O_579,N_9979,N_9605);
xnor UO_580 (O_580,N_9761,N_9655);
or UO_581 (O_581,N_9670,N_9694);
nand UO_582 (O_582,N_9931,N_9568);
nand UO_583 (O_583,N_9957,N_9894);
or UO_584 (O_584,N_9617,N_9625);
nand UO_585 (O_585,N_9893,N_9630);
and UO_586 (O_586,N_9971,N_9562);
nand UO_587 (O_587,N_9916,N_9792);
or UO_588 (O_588,N_9606,N_9624);
nand UO_589 (O_589,N_9922,N_9597);
nand UO_590 (O_590,N_9663,N_9657);
nor UO_591 (O_591,N_9948,N_9564);
and UO_592 (O_592,N_9524,N_9596);
or UO_593 (O_593,N_9997,N_9515);
or UO_594 (O_594,N_9883,N_9989);
and UO_595 (O_595,N_9755,N_9660);
or UO_596 (O_596,N_9749,N_9955);
nor UO_597 (O_597,N_9661,N_9501);
and UO_598 (O_598,N_9768,N_9668);
xor UO_599 (O_599,N_9604,N_9875);
nand UO_600 (O_600,N_9535,N_9913);
nand UO_601 (O_601,N_9579,N_9895);
or UO_602 (O_602,N_9937,N_9979);
nand UO_603 (O_603,N_9600,N_9525);
and UO_604 (O_604,N_9600,N_9913);
nor UO_605 (O_605,N_9849,N_9550);
nand UO_606 (O_606,N_9826,N_9704);
or UO_607 (O_607,N_9975,N_9648);
nor UO_608 (O_608,N_9554,N_9522);
or UO_609 (O_609,N_9587,N_9643);
and UO_610 (O_610,N_9589,N_9875);
nand UO_611 (O_611,N_9860,N_9610);
and UO_612 (O_612,N_9693,N_9751);
or UO_613 (O_613,N_9991,N_9579);
and UO_614 (O_614,N_9650,N_9621);
nor UO_615 (O_615,N_9540,N_9942);
or UO_616 (O_616,N_9514,N_9603);
nand UO_617 (O_617,N_9506,N_9630);
and UO_618 (O_618,N_9646,N_9618);
or UO_619 (O_619,N_9736,N_9812);
or UO_620 (O_620,N_9679,N_9828);
xor UO_621 (O_621,N_9876,N_9681);
and UO_622 (O_622,N_9661,N_9618);
nand UO_623 (O_623,N_9566,N_9530);
and UO_624 (O_624,N_9854,N_9785);
or UO_625 (O_625,N_9901,N_9976);
nor UO_626 (O_626,N_9971,N_9795);
nor UO_627 (O_627,N_9514,N_9685);
or UO_628 (O_628,N_9745,N_9651);
and UO_629 (O_629,N_9525,N_9828);
nor UO_630 (O_630,N_9853,N_9585);
and UO_631 (O_631,N_9928,N_9543);
nand UO_632 (O_632,N_9918,N_9875);
nand UO_633 (O_633,N_9959,N_9671);
or UO_634 (O_634,N_9554,N_9500);
nand UO_635 (O_635,N_9874,N_9803);
and UO_636 (O_636,N_9528,N_9779);
or UO_637 (O_637,N_9937,N_9689);
nand UO_638 (O_638,N_9653,N_9785);
or UO_639 (O_639,N_9858,N_9547);
nor UO_640 (O_640,N_9748,N_9755);
nor UO_641 (O_641,N_9547,N_9797);
or UO_642 (O_642,N_9521,N_9976);
nor UO_643 (O_643,N_9850,N_9685);
nand UO_644 (O_644,N_9642,N_9502);
and UO_645 (O_645,N_9889,N_9881);
and UO_646 (O_646,N_9966,N_9983);
nand UO_647 (O_647,N_9643,N_9943);
or UO_648 (O_648,N_9627,N_9769);
nor UO_649 (O_649,N_9941,N_9507);
and UO_650 (O_650,N_9995,N_9616);
nand UO_651 (O_651,N_9862,N_9599);
and UO_652 (O_652,N_9803,N_9885);
and UO_653 (O_653,N_9624,N_9787);
nand UO_654 (O_654,N_9734,N_9569);
nand UO_655 (O_655,N_9848,N_9546);
and UO_656 (O_656,N_9797,N_9579);
and UO_657 (O_657,N_9638,N_9530);
nand UO_658 (O_658,N_9999,N_9908);
nor UO_659 (O_659,N_9526,N_9671);
nand UO_660 (O_660,N_9919,N_9848);
or UO_661 (O_661,N_9908,N_9959);
and UO_662 (O_662,N_9642,N_9948);
xor UO_663 (O_663,N_9690,N_9658);
nor UO_664 (O_664,N_9680,N_9696);
and UO_665 (O_665,N_9522,N_9997);
and UO_666 (O_666,N_9896,N_9965);
and UO_667 (O_667,N_9609,N_9750);
nand UO_668 (O_668,N_9673,N_9712);
and UO_669 (O_669,N_9552,N_9561);
nor UO_670 (O_670,N_9512,N_9823);
nor UO_671 (O_671,N_9755,N_9732);
or UO_672 (O_672,N_9534,N_9788);
nand UO_673 (O_673,N_9862,N_9671);
and UO_674 (O_674,N_9946,N_9879);
and UO_675 (O_675,N_9694,N_9924);
and UO_676 (O_676,N_9566,N_9760);
nor UO_677 (O_677,N_9799,N_9979);
nand UO_678 (O_678,N_9868,N_9540);
or UO_679 (O_679,N_9570,N_9868);
nor UO_680 (O_680,N_9936,N_9766);
nand UO_681 (O_681,N_9800,N_9661);
or UO_682 (O_682,N_9588,N_9851);
or UO_683 (O_683,N_9732,N_9643);
nor UO_684 (O_684,N_9767,N_9507);
nand UO_685 (O_685,N_9678,N_9957);
nand UO_686 (O_686,N_9569,N_9519);
nand UO_687 (O_687,N_9711,N_9629);
and UO_688 (O_688,N_9893,N_9763);
or UO_689 (O_689,N_9768,N_9713);
or UO_690 (O_690,N_9934,N_9621);
and UO_691 (O_691,N_9591,N_9719);
and UO_692 (O_692,N_9668,N_9562);
nor UO_693 (O_693,N_9929,N_9858);
and UO_694 (O_694,N_9754,N_9767);
nor UO_695 (O_695,N_9535,N_9669);
nand UO_696 (O_696,N_9920,N_9934);
nor UO_697 (O_697,N_9864,N_9632);
nor UO_698 (O_698,N_9809,N_9508);
nor UO_699 (O_699,N_9987,N_9503);
nand UO_700 (O_700,N_9971,N_9968);
or UO_701 (O_701,N_9514,N_9573);
nor UO_702 (O_702,N_9674,N_9519);
nand UO_703 (O_703,N_9901,N_9581);
and UO_704 (O_704,N_9612,N_9706);
nand UO_705 (O_705,N_9590,N_9675);
or UO_706 (O_706,N_9682,N_9858);
or UO_707 (O_707,N_9870,N_9884);
and UO_708 (O_708,N_9689,N_9722);
and UO_709 (O_709,N_9901,N_9832);
xnor UO_710 (O_710,N_9644,N_9931);
nor UO_711 (O_711,N_9871,N_9539);
nor UO_712 (O_712,N_9672,N_9810);
and UO_713 (O_713,N_9861,N_9826);
or UO_714 (O_714,N_9970,N_9770);
nand UO_715 (O_715,N_9676,N_9982);
nor UO_716 (O_716,N_9845,N_9583);
nor UO_717 (O_717,N_9867,N_9644);
and UO_718 (O_718,N_9801,N_9695);
or UO_719 (O_719,N_9504,N_9872);
nor UO_720 (O_720,N_9959,N_9590);
or UO_721 (O_721,N_9527,N_9940);
or UO_722 (O_722,N_9622,N_9545);
nor UO_723 (O_723,N_9834,N_9957);
nor UO_724 (O_724,N_9887,N_9608);
nor UO_725 (O_725,N_9975,N_9647);
nand UO_726 (O_726,N_9608,N_9997);
xnor UO_727 (O_727,N_9635,N_9975);
or UO_728 (O_728,N_9937,N_9623);
xnor UO_729 (O_729,N_9605,N_9597);
and UO_730 (O_730,N_9760,N_9749);
or UO_731 (O_731,N_9697,N_9800);
or UO_732 (O_732,N_9945,N_9747);
nand UO_733 (O_733,N_9655,N_9868);
xor UO_734 (O_734,N_9897,N_9504);
nand UO_735 (O_735,N_9872,N_9573);
nor UO_736 (O_736,N_9996,N_9796);
nor UO_737 (O_737,N_9853,N_9651);
nor UO_738 (O_738,N_9878,N_9826);
nor UO_739 (O_739,N_9796,N_9608);
nor UO_740 (O_740,N_9503,N_9996);
or UO_741 (O_741,N_9957,N_9905);
nand UO_742 (O_742,N_9872,N_9992);
and UO_743 (O_743,N_9579,N_9877);
nor UO_744 (O_744,N_9600,N_9793);
and UO_745 (O_745,N_9537,N_9522);
nor UO_746 (O_746,N_9613,N_9854);
and UO_747 (O_747,N_9752,N_9885);
and UO_748 (O_748,N_9514,N_9893);
and UO_749 (O_749,N_9726,N_9730);
or UO_750 (O_750,N_9639,N_9794);
and UO_751 (O_751,N_9729,N_9606);
and UO_752 (O_752,N_9863,N_9777);
and UO_753 (O_753,N_9780,N_9637);
and UO_754 (O_754,N_9836,N_9942);
nand UO_755 (O_755,N_9808,N_9951);
and UO_756 (O_756,N_9501,N_9927);
and UO_757 (O_757,N_9700,N_9554);
nand UO_758 (O_758,N_9800,N_9821);
and UO_759 (O_759,N_9738,N_9677);
nand UO_760 (O_760,N_9636,N_9844);
or UO_761 (O_761,N_9996,N_9574);
nor UO_762 (O_762,N_9794,N_9594);
nor UO_763 (O_763,N_9991,N_9590);
nor UO_764 (O_764,N_9693,N_9776);
nand UO_765 (O_765,N_9753,N_9792);
nand UO_766 (O_766,N_9621,N_9879);
nor UO_767 (O_767,N_9902,N_9609);
and UO_768 (O_768,N_9783,N_9642);
or UO_769 (O_769,N_9911,N_9700);
or UO_770 (O_770,N_9774,N_9724);
or UO_771 (O_771,N_9747,N_9670);
nor UO_772 (O_772,N_9563,N_9684);
or UO_773 (O_773,N_9553,N_9796);
or UO_774 (O_774,N_9571,N_9758);
nor UO_775 (O_775,N_9956,N_9707);
nand UO_776 (O_776,N_9628,N_9906);
or UO_777 (O_777,N_9950,N_9517);
nand UO_778 (O_778,N_9729,N_9828);
nor UO_779 (O_779,N_9863,N_9869);
nand UO_780 (O_780,N_9742,N_9730);
nand UO_781 (O_781,N_9591,N_9855);
or UO_782 (O_782,N_9714,N_9817);
nor UO_783 (O_783,N_9524,N_9817);
nor UO_784 (O_784,N_9691,N_9980);
or UO_785 (O_785,N_9820,N_9850);
nand UO_786 (O_786,N_9677,N_9972);
nand UO_787 (O_787,N_9858,N_9574);
and UO_788 (O_788,N_9570,N_9611);
nor UO_789 (O_789,N_9606,N_9877);
and UO_790 (O_790,N_9554,N_9817);
nand UO_791 (O_791,N_9925,N_9507);
or UO_792 (O_792,N_9626,N_9675);
or UO_793 (O_793,N_9666,N_9941);
and UO_794 (O_794,N_9828,N_9596);
xnor UO_795 (O_795,N_9930,N_9876);
nor UO_796 (O_796,N_9594,N_9740);
or UO_797 (O_797,N_9957,N_9780);
or UO_798 (O_798,N_9677,N_9546);
or UO_799 (O_799,N_9725,N_9528);
or UO_800 (O_800,N_9759,N_9717);
and UO_801 (O_801,N_9961,N_9972);
nand UO_802 (O_802,N_9898,N_9789);
nor UO_803 (O_803,N_9809,N_9586);
nor UO_804 (O_804,N_9646,N_9874);
nand UO_805 (O_805,N_9959,N_9825);
or UO_806 (O_806,N_9851,N_9914);
nand UO_807 (O_807,N_9785,N_9879);
and UO_808 (O_808,N_9843,N_9864);
and UO_809 (O_809,N_9700,N_9814);
and UO_810 (O_810,N_9970,N_9882);
nor UO_811 (O_811,N_9509,N_9929);
nand UO_812 (O_812,N_9981,N_9997);
nand UO_813 (O_813,N_9704,N_9871);
and UO_814 (O_814,N_9796,N_9877);
nor UO_815 (O_815,N_9994,N_9815);
nor UO_816 (O_816,N_9516,N_9534);
nand UO_817 (O_817,N_9796,N_9984);
and UO_818 (O_818,N_9614,N_9751);
nand UO_819 (O_819,N_9843,N_9703);
nor UO_820 (O_820,N_9588,N_9749);
and UO_821 (O_821,N_9699,N_9936);
xnor UO_822 (O_822,N_9771,N_9660);
and UO_823 (O_823,N_9530,N_9619);
or UO_824 (O_824,N_9866,N_9995);
nor UO_825 (O_825,N_9837,N_9649);
and UO_826 (O_826,N_9709,N_9632);
or UO_827 (O_827,N_9982,N_9577);
xnor UO_828 (O_828,N_9802,N_9926);
and UO_829 (O_829,N_9699,N_9741);
nor UO_830 (O_830,N_9502,N_9727);
nand UO_831 (O_831,N_9591,N_9975);
and UO_832 (O_832,N_9530,N_9660);
nor UO_833 (O_833,N_9997,N_9734);
and UO_834 (O_834,N_9853,N_9906);
or UO_835 (O_835,N_9760,N_9647);
or UO_836 (O_836,N_9851,N_9691);
and UO_837 (O_837,N_9972,N_9997);
or UO_838 (O_838,N_9880,N_9879);
and UO_839 (O_839,N_9843,N_9573);
and UO_840 (O_840,N_9794,N_9650);
nand UO_841 (O_841,N_9888,N_9839);
nor UO_842 (O_842,N_9656,N_9641);
and UO_843 (O_843,N_9665,N_9732);
nor UO_844 (O_844,N_9805,N_9748);
and UO_845 (O_845,N_9564,N_9640);
nand UO_846 (O_846,N_9756,N_9565);
nand UO_847 (O_847,N_9773,N_9646);
and UO_848 (O_848,N_9509,N_9618);
or UO_849 (O_849,N_9604,N_9665);
nand UO_850 (O_850,N_9534,N_9636);
and UO_851 (O_851,N_9733,N_9678);
nor UO_852 (O_852,N_9543,N_9938);
xnor UO_853 (O_853,N_9831,N_9761);
and UO_854 (O_854,N_9854,N_9819);
nor UO_855 (O_855,N_9787,N_9611);
or UO_856 (O_856,N_9973,N_9718);
nor UO_857 (O_857,N_9581,N_9574);
and UO_858 (O_858,N_9915,N_9849);
or UO_859 (O_859,N_9738,N_9607);
nand UO_860 (O_860,N_9881,N_9535);
nor UO_861 (O_861,N_9934,N_9516);
nor UO_862 (O_862,N_9931,N_9915);
nand UO_863 (O_863,N_9857,N_9751);
and UO_864 (O_864,N_9996,N_9547);
xnor UO_865 (O_865,N_9749,N_9910);
and UO_866 (O_866,N_9691,N_9810);
and UO_867 (O_867,N_9812,N_9503);
xnor UO_868 (O_868,N_9634,N_9673);
or UO_869 (O_869,N_9632,N_9590);
and UO_870 (O_870,N_9972,N_9675);
nand UO_871 (O_871,N_9990,N_9657);
nor UO_872 (O_872,N_9833,N_9897);
nor UO_873 (O_873,N_9995,N_9854);
nor UO_874 (O_874,N_9696,N_9901);
and UO_875 (O_875,N_9652,N_9601);
nand UO_876 (O_876,N_9804,N_9630);
and UO_877 (O_877,N_9589,N_9732);
or UO_878 (O_878,N_9936,N_9870);
nand UO_879 (O_879,N_9761,N_9909);
nor UO_880 (O_880,N_9653,N_9981);
nor UO_881 (O_881,N_9759,N_9600);
xor UO_882 (O_882,N_9596,N_9547);
and UO_883 (O_883,N_9717,N_9970);
nand UO_884 (O_884,N_9978,N_9960);
nand UO_885 (O_885,N_9942,N_9536);
nor UO_886 (O_886,N_9531,N_9733);
or UO_887 (O_887,N_9548,N_9659);
nor UO_888 (O_888,N_9525,N_9626);
nand UO_889 (O_889,N_9841,N_9911);
and UO_890 (O_890,N_9659,N_9751);
or UO_891 (O_891,N_9552,N_9900);
nand UO_892 (O_892,N_9909,N_9691);
xnor UO_893 (O_893,N_9851,N_9592);
or UO_894 (O_894,N_9775,N_9931);
nor UO_895 (O_895,N_9938,N_9768);
or UO_896 (O_896,N_9861,N_9569);
or UO_897 (O_897,N_9796,N_9857);
nand UO_898 (O_898,N_9641,N_9587);
or UO_899 (O_899,N_9786,N_9872);
nor UO_900 (O_900,N_9665,N_9922);
nor UO_901 (O_901,N_9788,N_9941);
nand UO_902 (O_902,N_9963,N_9528);
nand UO_903 (O_903,N_9751,N_9968);
or UO_904 (O_904,N_9526,N_9957);
nor UO_905 (O_905,N_9897,N_9644);
or UO_906 (O_906,N_9572,N_9713);
and UO_907 (O_907,N_9848,N_9676);
nor UO_908 (O_908,N_9851,N_9548);
or UO_909 (O_909,N_9848,N_9635);
and UO_910 (O_910,N_9845,N_9854);
or UO_911 (O_911,N_9716,N_9686);
or UO_912 (O_912,N_9822,N_9763);
nor UO_913 (O_913,N_9586,N_9752);
nor UO_914 (O_914,N_9760,N_9900);
nand UO_915 (O_915,N_9810,N_9909);
nor UO_916 (O_916,N_9961,N_9871);
and UO_917 (O_917,N_9935,N_9873);
nor UO_918 (O_918,N_9935,N_9811);
or UO_919 (O_919,N_9880,N_9677);
and UO_920 (O_920,N_9618,N_9734);
nand UO_921 (O_921,N_9998,N_9770);
nor UO_922 (O_922,N_9932,N_9546);
or UO_923 (O_923,N_9674,N_9865);
or UO_924 (O_924,N_9613,N_9575);
and UO_925 (O_925,N_9822,N_9616);
or UO_926 (O_926,N_9810,N_9791);
nand UO_927 (O_927,N_9533,N_9575);
or UO_928 (O_928,N_9773,N_9785);
nor UO_929 (O_929,N_9586,N_9987);
nand UO_930 (O_930,N_9671,N_9938);
nand UO_931 (O_931,N_9552,N_9670);
or UO_932 (O_932,N_9552,N_9651);
or UO_933 (O_933,N_9981,N_9920);
or UO_934 (O_934,N_9523,N_9706);
or UO_935 (O_935,N_9974,N_9787);
or UO_936 (O_936,N_9873,N_9502);
nor UO_937 (O_937,N_9972,N_9766);
nor UO_938 (O_938,N_9731,N_9629);
and UO_939 (O_939,N_9553,N_9530);
nand UO_940 (O_940,N_9588,N_9857);
or UO_941 (O_941,N_9816,N_9833);
nor UO_942 (O_942,N_9561,N_9910);
nor UO_943 (O_943,N_9790,N_9982);
or UO_944 (O_944,N_9623,N_9747);
and UO_945 (O_945,N_9541,N_9634);
nor UO_946 (O_946,N_9698,N_9833);
nor UO_947 (O_947,N_9660,N_9570);
nor UO_948 (O_948,N_9561,N_9522);
and UO_949 (O_949,N_9873,N_9697);
nor UO_950 (O_950,N_9831,N_9868);
and UO_951 (O_951,N_9613,N_9524);
or UO_952 (O_952,N_9853,N_9971);
or UO_953 (O_953,N_9682,N_9715);
and UO_954 (O_954,N_9915,N_9938);
nand UO_955 (O_955,N_9843,N_9638);
or UO_956 (O_956,N_9724,N_9885);
nor UO_957 (O_957,N_9977,N_9587);
or UO_958 (O_958,N_9676,N_9726);
nand UO_959 (O_959,N_9874,N_9846);
nand UO_960 (O_960,N_9884,N_9593);
nor UO_961 (O_961,N_9727,N_9774);
nand UO_962 (O_962,N_9674,N_9822);
nor UO_963 (O_963,N_9844,N_9580);
or UO_964 (O_964,N_9980,N_9953);
or UO_965 (O_965,N_9708,N_9754);
or UO_966 (O_966,N_9678,N_9641);
nand UO_967 (O_967,N_9696,N_9684);
or UO_968 (O_968,N_9846,N_9929);
nor UO_969 (O_969,N_9795,N_9874);
and UO_970 (O_970,N_9915,N_9599);
or UO_971 (O_971,N_9600,N_9846);
nand UO_972 (O_972,N_9926,N_9755);
and UO_973 (O_973,N_9973,N_9654);
nand UO_974 (O_974,N_9572,N_9994);
nor UO_975 (O_975,N_9638,N_9996);
nand UO_976 (O_976,N_9557,N_9822);
or UO_977 (O_977,N_9987,N_9720);
nand UO_978 (O_978,N_9870,N_9951);
nor UO_979 (O_979,N_9749,N_9825);
or UO_980 (O_980,N_9855,N_9607);
nor UO_981 (O_981,N_9741,N_9851);
nand UO_982 (O_982,N_9705,N_9854);
or UO_983 (O_983,N_9611,N_9550);
nand UO_984 (O_984,N_9711,N_9975);
nand UO_985 (O_985,N_9624,N_9537);
or UO_986 (O_986,N_9815,N_9518);
nand UO_987 (O_987,N_9524,N_9535);
nand UO_988 (O_988,N_9666,N_9781);
and UO_989 (O_989,N_9666,N_9546);
nor UO_990 (O_990,N_9754,N_9753);
or UO_991 (O_991,N_9609,N_9652);
or UO_992 (O_992,N_9545,N_9974);
nor UO_993 (O_993,N_9643,N_9989);
nand UO_994 (O_994,N_9681,N_9971);
nor UO_995 (O_995,N_9799,N_9598);
or UO_996 (O_996,N_9657,N_9518);
and UO_997 (O_997,N_9672,N_9803);
or UO_998 (O_998,N_9953,N_9638);
nand UO_999 (O_999,N_9542,N_9856);
nor UO_1000 (O_1000,N_9825,N_9842);
or UO_1001 (O_1001,N_9997,N_9948);
and UO_1002 (O_1002,N_9658,N_9784);
nor UO_1003 (O_1003,N_9699,N_9844);
nand UO_1004 (O_1004,N_9743,N_9585);
or UO_1005 (O_1005,N_9897,N_9847);
nor UO_1006 (O_1006,N_9635,N_9511);
or UO_1007 (O_1007,N_9504,N_9636);
nor UO_1008 (O_1008,N_9925,N_9768);
nor UO_1009 (O_1009,N_9773,N_9783);
or UO_1010 (O_1010,N_9970,N_9872);
nor UO_1011 (O_1011,N_9965,N_9759);
nor UO_1012 (O_1012,N_9877,N_9907);
nor UO_1013 (O_1013,N_9781,N_9725);
nand UO_1014 (O_1014,N_9621,N_9653);
nand UO_1015 (O_1015,N_9537,N_9954);
or UO_1016 (O_1016,N_9549,N_9703);
nand UO_1017 (O_1017,N_9618,N_9836);
nand UO_1018 (O_1018,N_9750,N_9818);
or UO_1019 (O_1019,N_9637,N_9925);
nor UO_1020 (O_1020,N_9874,N_9680);
nand UO_1021 (O_1021,N_9566,N_9538);
and UO_1022 (O_1022,N_9624,N_9747);
or UO_1023 (O_1023,N_9529,N_9547);
nand UO_1024 (O_1024,N_9899,N_9987);
and UO_1025 (O_1025,N_9936,N_9871);
nor UO_1026 (O_1026,N_9960,N_9787);
nand UO_1027 (O_1027,N_9906,N_9948);
nand UO_1028 (O_1028,N_9903,N_9730);
nor UO_1029 (O_1029,N_9770,N_9860);
nand UO_1030 (O_1030,N_9937,N_9666);
and UO_1031 (O_1031,N_9500,N_9795);
and UO_1032 (O_1032,N_9986,N_9846);
nor UO_1033 (O_1033,N_9760,N_9931);
nor UO_1034 (O_1034,N_9814,N_9669);
nand UO_1035 (O_1035,N_9971,N_9716);
nor UO_1036 (O_1036,N_9798,N_9960);
or UO_1037 (O_1037,N_9662,N_9527);
or UO_1038 (O_1038,N_9832,N_9913);
or UO_1039 (O_1039,N_9937,N_9578);
xnor UO_1040 (O_1040,N_9655,N_9695);
nand UO_1041 (O_1041,N_9983,N_9852);
xnor UO_1042 (O_1042,N_9602,N_9610);
nor UO_1043 (O_1043,N_9912,N_9957);
nor UO_1044 (O_1044,N_9974,N_9516);
xnor UO_1045 (O_1045,N_9959,N_9943);
xor UO_1046 (O_1046,N_9525,N_9888);
or UO_1047 (O_1047,N_9861,N_9820);
and UO_1048 (O_1048,N_9569,N_9719);
or UO_1049 (O_1049,N_9934,N_9909);
nor UO_1050 (O_1050,N_9644,N_9894);
nor UO_1051 (O_1051,N_9970,N_9723);
and UO_1052 (O_1052,N_9996,N_9656);
nor UO_1053 (O_1053,N_9900,N_9896);
or UO_1054 (O_1054,N_9997,N_9840);
and UO_1055 (O_1055,N_9950,N_9524);
nor UO_1056 (O_1056,N_9862,N_9600);
nand UO_1057 (O_1057,N_9504,N_9573);
nor UO_1058 (O_1058,N_9686,N_9706);
or UO_1059 (O_1059,N_9615,N_9919);
nand UO_1060 (O_1060,N_9764,N_9759);
nor UO_1061 (O_1061,N_9818,N_9633);
nor UO_1062 (O_1062,N_9896,N_9553);
nor UO_1063 (O_1063,N_9594,N_9806);
or UO_1064 (O_1064,N_9633,N_9653);
nor UO_1065 (O_1065,N_9604,N_9631);
nand UO_1066 (O_1066,N_9690,N_9675);
nand UO_1067 (O_1067,N_9720,N_9995);
and UO_1068 (O_1068,N_9741,N_9743);
xor UO_1069 (O_1069,N_9732,N_9603);
or UO_1070 (O_1070,N_9561,N_9974);
or UO_1071 (O_1071,N_9565,N_9566);
nor UO_1072 (O_1072,N_9830,N_9570);
nor UO_1073 (O_1073,N_9687,N_9678);
nand UO_1074 (O_1074,N_9912,N_9980);
or UO_1075 (O_1075,N_9632,N_9746);
or UO_1076 (O_1076,N_9608,N_9504);
and UO_1077 (O_1077,N_9718,N_9641);
and UO_1078 (O_1078,N_9517,N_9576);
nor UO_1079 (O_1079,N_9546,N_9678);
nor UO_1080 (O_1080,N_9987,N_9873);
or UO_1081 (O_1081,N_9723,N_9886);
nand UO_1082 (O_1082,N_9721,N_9646);
or UO_1083 (O_1083,N_9646,N_9785);
and UO_1084 (O_1084,N_9500,N_9783);
or UO_1085 (O_1085,N_9803,N_9891);
and UO_1086 (O_1086,N_9757,N_9604);
nor UO_1087 (O_1087,N_9796,N_9513);
or UO_1088 (O_1088,N_9998,N_9913);
nor UO_1089 (O_1089,N_9687,N_9945);
nor UO_1090 (O_1090,N_9848,N_9609);
nand UO_1091 (O_1091,N_9844,N_9579);
or UO_1092 (O_1092,N_9738,N_9829);
and UO_1093 (O_1093,N_9935,N_9522);
nor UO_1094 (O_1094,N_9861,N_9917);
nor UO_1095 (O_1095,N_9879,N_9847);
nand UO_1096 (O_1096,N_9716,N_9646);
nor UO_1097 (O_1097,N_9885,N_9970);
and UO_1098 (O_1098,N_9784,N_9775);
or UO_1099 (O_1099,N_9745,N_9844);
nand UO_1100 (O_1100,N_9572,N_9563);
or UO_1101 (O_1101,N_9626,N_9595);
nand UO_1102 (O_1102,N_9716,N_9596);
or UO_1103 (O_1103,N_9818,N_9885);
nand UO_1104 (O_1104,N_9900,N_9871);
or UO_1105 (O_1105,N_9502,N_9800);
nor UO_1106 (O_1106,N_9955,N_9745);
nand UO_1107 (O_1107,N_9586,N_9827);
xor UO_1108 (O_1108,N_9514,N_9501);
nand UO_1109 (O_1109,N_9761,N_9501);
nand UO_1110 (O_1110,N_9867,N_9559);
and UO_1111 (O_1111,N_9521,N_9625);
or UO_1112 (O_1112,N_9663,N_9874);
or UO_1113 (O_1113,N_9761,N_9764);
and UO_1114 (O_1114,N_9630,N_9788);
and UO_1115 (O_1115,N_9953,N_9539);
and UO_1116 (O_1116,N_9998,N_9991);
or UO_1117 (O_1117,N_9642,N_9883);
or UO_1118 (O_1118,N_9778,N_9888);
nand UO_1119 (O_1119,N_9509,N_9820);
or UO_1120 (O_1120,N_9939,N_9564);
and UO_1121 (O_1121,N_9641,N_9991);
or UO_1122 (O_1122,N_9813,N_9925);
xor UO_1123 (O_1123,N_9597,N_9772);
and UO_1124 (O_1124,N_9982,N_9833);
nor UO_1125 (O_1125,N_9926,N_9902);
or UO_1126 (O_1126,N_9597,N_9585);
or UO_1127 (O_1127,N_9756,N_9804);
nand UO_1128 (O_1128,N_9825,N_9588);
or UO_1129 (O_1129,N_9977,N_9875);
nand UO_1130 (O_1130,N_9831,N_9581);
nand UO_1131 (O_1131,N_9879,N_9504);
and UO_1132 (O_1132,N_9986,N_9892);
nand UO_1133 (O_1133,N_9552,N_9592);
nand UO_1134 (O_1134,N_9524,N_9653);
and UO_1135 (O_1135,N_9867,N_9994);
and UO_1136 (O_1136,N_9941,N_9564);
nor UO_1137 (O_1137,N_9976,N_9729);
or UO_1138 (O_1138,N_9775,N_9634);
nand UO_1139 (O_1139,N_9869,N_9616);
and UO_1140 (O_1140,N_9535,N_9802);
nor UO_1141 (O_1141,N_9734,N_9960);
nor UO_1142 (O_1142,N_9758,N_9894);
or UO_1143 (O_1143,N_9822,N_9699);
and UO_1144 (O_1144,N_9641,N_9716);
or UO_1145 (O_1145,N_9988,N_9916);
nor UO_1146 (O_1146,N_9590,N_9638);
or UO_1147 (O_1147,N_9777,N_9813);
nor UO_1148 (O_1148,N_9967,N_9875);
or UO_1149 (O_1149,N_9992,N_9620);
nor UO_1150 (O_1150,N_9579,N_9806);
or UO_1151 (O_1151,N_9623,N_9742);
nand UO_1152 (O_1152,N_9836,N_9737);
and UO_1153 (O_1153,N_9978,N_9539);
or UO_1154 (O_1154,N_9604,N_9643);
nor UO_1155 (O_1155,N_9998,N_9814);
nand UO_1156 (O_1156,N_9810,N_9908);
or UO_1157 (O_1157,N_9930,N_9670);
nor UO_1158 (O_1158,N_9603,N_9879);
nand UO_1159 (O_1159,N_9902,N_9797);
or UO_1160 (O_1160,N_9874,N_9780);
and UO_1161 (O_1161,N_9821,N_9720);
and UO_1162 (O_1162,N_9729,N_9838);
or UO_1163 (O_1163,N_9634,N_9945);
and UO_1164 (O_1164,N_9863,N_9679);
and UO_1165 (O_1165,N_9870,N_9616);
nand UO_1166 (O_1166,N_9525,N_9609);
or UO_1167 (O_1167,N_9946,N_9560);
and UO_1168 (O_1168,N_9529,N_9704);
or UO_1169 (O_1169,N_9541,N_9633);
and UO_1170 (O_1170,N_9900,N_9976);
or UO_1171 (O_1171,N_9569,N_9998);
nor UO_1172 (O_1172,N_9837,N_9616);
nor UO_1173 (O_1173,N_9882,N_9924);
nor UO_1174 (O_1174,N_9737,N_9969);
nor UO_1175 (O_1175,N_9933,N_9865);
or UO_1176 (O_1176,N_9748,N_9654);
and UO_1177 (O_1177,N_9608,N_9524);
nand UO_1178 (O_1178,N_9535,N_9752);
and UO_1179 (O_1179,N_9597,N_9908);
nand UO_1180 (O_1180,N_9980,N_9856);
and UO_1181 (O_1181,N_9998,N_9714);
and UO_1182 (O_1182,N_9520,N_9519);
nand UO_1183 (O_1183,N_9782,N_9795);
xor UO_1184 (O_1184,N_9724,N_9780);
or UO_1185 (O_1185,N_9533,N_9834);
or UO_1186 (O_1186,N_9933,N_9965);
or UO_1187 (O_1187,N_9683,N_9583);
nand UO_1188 (O_1188,N_9988,N_9691);
and UO_1189 (O_1189,N_9799,N_9507);
and UO_1190 (O_1190,N_9878,N_9931);
and UO_1191 (O_1191,N_9849,N_9511);
nor UO_1192 (O_1192,N_9728,N_9655);
and UO_1193 (O_1193,N_9688,N_9868);
and UO_1194 (O_1194,N_9634,N_9832);
or UO_1195 (O_1195,N_9811,N_9506);
nor UO_1196 (O_1196,N_9854,N_9524);
nor UO_1197 (O_1197,N_9512,N_9719);
nand UO_1198 (O_1198,N_9843,N_9591);
or UO_1199 (O_1199,N_9567,N_9929);
and UO_1200 (O_1200,N_9710,N_9940);
xor UO_1201 (O_1201,N_9564,N_9626);
or UO_1202 (O_1202,N_9958,N_9752);
or UO_1203 (O_1203,N_9572,N_9887);
or UO_1204 (O_1204,N_9978,N_9799);
or UO_1205 (O_1205,N_9720,N_9733);
or UO_1206 (O_1206,N_9877,N_9751);
or UO_1207 (O_1207,N_9646,N_9797);
nand UO_1208 (O_1208,N_9668,N_9909);
or UO_1209 (O_1209,N_9803,N_9818);
nand UO_1210 (O_1210,N_9758,N_9776);
and UO_1211 (O_1211,N_9706,N_9875);
nor UO_1212 (O_1212,N_9877,N_9675);
or UO_1213 (O_1213,N_9921,N_9683);
and UO_1214 (O_1214,N_9758,N_9800);
nand UO_1215 (O_1215,N_9745,N_9521);
and UO_1216 (O_1216,N_9643,N_9973);
nor UO_1217 (O_1217,N_9960,N_9800);
and UO_1218 (O_1218,N_9820,N_9953);
and UO_1219 (O_1219,N_9526,N_9760);
or UO_1220 (O_1220,N_9736,N_9938);
or UO_1221 (O_1221,N_9839,N_9800);
or UO_1222 (O_1222,N_9615,N_9745);
or UO_1223 (O_1223,N_9775,N_9558);
xor UO_1224 (O_1224,N_9634,N_9850);
and UO_1225 (O_1225,N_9988,N_9679);
and UO_1226 (O_1226,N_9669,N_9597);
nand UO_1227 (O_1227,N_9659,N_9822);
or UO_1228 (O_1228,N_9809,N_9997);
nor UO_1229 (O_1229,N_9503,N_9628);
nand UO_1230 (O_1230,N_9900,N_9980);
nor UO_1231 (O_1231,N_9851,N_9676);
nor UO_1232 (O_1232,N_9834,N_9524);
and UO_1233 (O_1233,N_9781,N_9686);
nor UO_1234 (O_1234,N_9557,N_9824);
and UO_1235 (O_1235,N_9861,N_9859);
and UO_1236 (O_1236,N_9895,N_9815);
nand UO_1237 (O_1237,N_9718,N_9523);
and UO_1238 (O_1238,N_9569,N_9962);
or UO_1239 (O_1239,N_9597,N_9904);
nor UO_1240 (O_1240,N_9708,N_9611);
nand UO_1241 (O_1241,N_9568,N_9893);
or UO_1242 (O_1242,N_9782,N_9672);
nor UO_1243 (O_1243,N_9795,N_9503);
nor UO_1244 (O_1244,N_9886,N_9953);
or UO_1245 (O_1245,N_9503,N_9830);
or UO_1246 (O_1246,N_9861,N_9823);
nor UO_1247 (O_1247,N_9925,N_9991);
nor UO_1248 (O_1248,N_9608,N_9807);
nor UO_1249 (O_1249,N_9676,N_9611);
nor UO_1250 (O_1250,N_9905,N_9792);
or UO_1251 (O_1251,N_9753,N_9670);
nor UO_1252 (O_1252,N_9793,N_9965);
or UO_1253 (O_1253,N_9512,N_9705);
nand UO_1254 (O_1254,N_9915,N_9536);
and UO_1255 (O_1255,N_9846,N_9817);
nor UO_1256 (O_1256,N_9830,N_9671);
and UO_1257 (O_1257,N_9940,N_9648);
nand UO_1258 (O_1258,N_9741,N_9831);
nand UO_1259 (O_1259,N_9535,N_9614);
or UO_1260 (O_1260,N_9767,N_9879);
or UO_1261 (O_1261,N_9712,N_9517);
nand UO_1262 (O_1262,N_9873,N_9648);
or UO_1263 (O_1263,N_9623,N_9912);
or UO_1264 (O_1264,N_9729,N_9932);
or UO_1265 (O_1265,N_9791,N_9832);
or UO_1266 (O_1266,N_9884,N_9566);
and UO_1267 (O_1267,N_9755,N_9743);
nand UO_1268 (O_1268,N_9737,N_9768);
or UO_1269 (O_1269,N_9970,N_9659);
nand UO_1270 (O_1270,N_9711,N_9969);
nand UO_1271 (O_1271,N_9576,N_9754);
and UO_1272 (O_1272,N_9813,N_9714);
or UO_1273 (O_1273,N_9515,N_9783);
or UO_1274 (O_1274,N_9697,N_9895);
or UO_1275 (O_1275,N_9511,N_9696);
or UO_1276 (O_1276,N_9551,N_9777);
or UO_1277 (O_1277,N_9624,N_9963);
nor UO_1278 (O_1278,N_9751,N_9698);
and UO_1279 (O_1279,N_9759,N_9946);
nand UO_1280 (O_1280,N_9689,N_9885);
nand UO_1281 (O_1281,N_9598,N_9730);
or UO_1282 (O_1282,N_9973,N_9918);
nand UO_1283 (O_1283,N_9959,N_9743);
nor UO_1284 (O_1284,N_9808,N_9509);
or UO_1285 (O_1285,N_9706,N_9689);
nand UO_1286 (O_1286,N_9616,N_9774);
and UO_1287 (O_1287,N_9733,N_9832);
and UO_1288 (O_1288,N_9650,N_9593);
nand UO_1289 (O_1289,N_9704,N_9995);
nor UO_1290 (O_1290,N_9953,N_9635);
or UO_1291 (O_1291,N_9569,N_9802);
and UO_1292 (O_1292,N_9647,N_9657);
nand UO_1293 (O_1293,N_9580,N_9987);
nand UO_1294 (O_1294,N_9833,N_9569);
xnor UO_1295 (O_1295,N_9787,N_9961);
xnor UO_1296 (O_1296,N_9651,N_9863);
or UO_1297 (O_1297,N_9897,N_9917);
and UO_1298 (O_1298,N_9688,N_9682);
and UO_1299 (O_1299,N_9859,N_9663);
and UO_1300 (O_1300,N_9518,N_9844);
nor UO_1301 (O_1301,N_9602,N_9893);
and UO_1302 (O_1302,N_9819,N_9557);
nand UO_1303 (O_1303,N_9768,N_9662);
or UO_1304 (O_1304,N_9836,N_9782);
or UO_1305 (O_1305,N_9616,N_9948);
nand UO_1306 (O_1306,N_9725,N_9819);
and UO_1307 (O_1307,N_9973,N_9819);
nand UO_1308 (O_1308,N_9663,N_9745);
and UO_1309 (O_1309,N_9766,N_9772);
nand UO_1310 (O_1310,N_9861,N_9697);
and UO_1311 (O_1311,N_9976,N_9802);
and UO_1312 (O_1312,N_9678,N_9947);
or UO_1313 (O_1313,N_9672,N_9885);
and UO_1314 (O_1314,N_9964,N_9507);
and UO_1315 (O_1315,N_9911,N_9752);
or UO_1316 (O_1316,N_9727,N_9823);
and UO_1317 (O_1317,N_9527,N_9550);
or UO_1318 (O_1318,N_9628,N_9997);
or UO_1319 (O_1319,N_9896,N_9711);
and UO_1320 (O_1320,N_9738,N_9528);
nor UO_1321 (O_1321,N_9932,N_9710);
or UO_1322 (O_1322,N_9732,N_9747);
nand UO_1323 (O_1323,N_9834,N_9684);
and UO_1324 (O_1324,N_9829,N_9642);
or UO_1325 (O_1325,N_9832,N_9991);
nand UO_1326 (O_1326,N_9766,N_9629);
nor UO_1327 (O_1327,N_9612,N_9931);
and UO_1328 (O_1328,N_9986,N_9764);
or UO_1329 (O_1329,N_9746,N_9702);
nand UO_1330 (O_1330,N_9792,N_9515);
nand UO_1331 (O_1331,N_9652,N_9853);
and UO_1332 (O_1332,N_9800,N_9808);
or UO_1333 (O_1333,N_9533,N_9970);
and UO_1334 (O_1334,N_9840,N_9959);
or UO_1335 (O_1335,N_9625,N_9801);
nor UO_1336 (O_1336,N_9693,N_9558);
or UO_1337 (O_1337,N_9850,N_9750);
nor UO_1338 (O_1338,N_9763,N_9587);
and UO_1339 (O_1339,N_9505,N_9657);
and UO_1340 (O_1340,N_9599,N_9857);
and UO_1341 (O_1341,N_9598,N_9602);
nor UO_1342 (O_1342,N_9516,N_9726);
nand UO_1343 (O_1343,N_9921,N_9787);
and UO_1344 (O_1344,N_9754,N_9803);
or UO_1345 (O_1345,N_9705,N_9555);
nand UO_1346 (O_1346,N_9855,N_9980);
and UO_1347 (O_1347,N_9560,N_9770);
and UO_1348 (O_1348,N_9558,N_9743);
or UO_1349 (O_1349,N_9502,N_9541);
and UO_1350 (O_1350,N_9633,N_9521);
or UO_1351 (O_1351,N_9762,N_9558);
and UO_1352 (O_1352,N_9956,N_9905);
and UO_1353 (O_1353,N_9826,N_9939);
and UO_1354 (O_1354,N_9976,N_9538);
nand UO_1355 (O_1355,N_9539,N_9869);
nand UO_1356 (O_1356,N_9652,N_9674);
nor UO_1357 (O_1357,N_9893,N_9927);
nand UO_1358 (O_1358,N_9963,N_9659);
nand UO_1359 (O_1359,N_9634,N_9877);
or UO_1360 (O_1360,N_9794,N_9956);
nand UO_1361 (O_1361,N_9924,N_9592);
or UO_1362 (O_1362,N_9775,N_9986);
nor UO_1363 (O_1363,N_9894,N_9690);
nand UO_1364 (O_1364,N_9567,N_9909);
nor UO_1365 (O_1365,N_9917,N_9931);
and UO_1366 (O_1366,N_9896,N_9664);
and UO_1367 (O_1367,N_9766,N_9631);
nor UO_1368 (O_1368,N_9669,N_9676);
nand UO_1369 (O_1369,N_9620,N_9743);
or UO_1370 (O_1370,N_9562,N_9676);
nand UO_1371 (O_1371,N_9991,N_9750);
and UO_1372 (O_1372,N_9920,N_9893);
nor UO_1373 (O_1373,N_9860,N_9618);
or UO_1374 (O_1374,N_9542,N_9874);
nand UO_1375 (O_1375,N_9582,N_9601);
nor UO_1376 (O_1376,N_9832,N_9826);
or UO_1377 (O_1377,N_9571,N_9998);
or UO_1378 (O_1378,N_9856,N_9817);
nand UO_1379 (O_1379,N_9648,N_9962);
xnor UO_1380 (O_1380,N_9847,N_9910);
nor UO_1381 (O_1381,N_9891,N_9918);
nor UO_1382 (O_1382,N_9933,N_9709);
or UO_1383 (O_1383,N_9947,N_9552);
and UO_1384 (O_1384,N_9891,N_9600);
and UO_1385 (O_1385,N_9723,N_9636);
or UO_1386 (O_1386,N_9673,N_9566);
nand UO_1387 (O_1387,N_9895,N_9568);
nand UO_1388 (O_1388,N_9871,N_9703);
or UO_1389 (O_1389,N_9665,N_9799);
nor UO_1390 (O_1390,N_9953,N_9589);
nor UO_1391 (O_1391,N_9642,N_9969);
and UO_1392 (O_1392,N_9810,N_9767);
or UO_1393 (O_1393,N_9619,N_9630);
nor UO_1394 (O_1394,N_9805,N_9720);
or UO_1395 (O_1395,N_9858,N_9959);
or UO_1396 (O_1396,N_9769,N_9573);
nand UO_1397 (O_1397,N_9880,N_9991);
and UO_1398 (O_1398,N_9965,N_9551);
nor UO_1399 (O_1399,N_9692,N_9696);
and UO_1400 (O_1400,N_9925,N_9806);
nor UO_1401 (O_1401,N_9687,N_9671);
or UO_1402 (O_1402,N_9881,N_9901);
or UO_1403 (O_1403,N_9553,N_9773);
xor UO_1404 (O_1404,N_9886,N_9939);
or UO_1405 (O_1405,N_9683,N_9767);
or UO_1406 (O_1406,N_9969,N_9579);
nand UO_1407 (O_1407,N_9692,N_9716);
nor UO_1408 (O_1408,N_9808,N_9732);
or UO_1409 (O_1409,N_9955,N_9859);
and UO_1410 (O_1410,N_9981,N_9923);
and UO_1411 (O_1411,N_9597,N_9913);
and UO_1412 (O_1412,N_9608,N_9750);
and UO_1413 (O_1413,N_9685,N_9619);
or UO_1414 (O_1414,N_9840,N_9718);
nand UO_1415 (O_1415,N_9870,N_9785);
nor UO_1416 (O_1416,N_9648,N_9886);
nand UO_1417 (O_1417,N_9676,N_9778);
or UO_1418 (O_1418,N_9545,N_9768);
or UO_1419 (O_1419,N_9762,N_9778);
or UO_1420 (O_1420,N_9788,N_9575);
or UO_1421 (O_1421,N_9688,N_9745);
or UO_1422 (O_1422,N_9829,N_9817);
and UO_1423 (O_1423,N_9584,N_9728);
or UO_1424 (O_1424,N_9584,N_9685);
and UO_1425 (O_1425,N_9949,N_9713);
nor UO_1426 (O_1426,N_9623,N_9551);
nand UO_1427 (O_1427,N_9711,N_9633);
xor UO_1428 (O_1428,N_9850,N_9843);
nor UO_1429 (O_1429,N_9958,N_9971);
nand UO_1430 (O_1430,N_9946,N_9593);
or UO_1431 (O_1431,N_9847,N_9902);
and UO_1432 (O_1432,N_9714,N_9652);
and UO_1433 (O_1433,N_9791,N_9522);
xnor UO_1434 (O_1434,N_9578,N_9760);
or UO_1435 (O_1435,N_9698,N_9667);
and UO_1436 (O_1436,N_9642,N_9553);
nor UO_1437 (O_1437,N_9937,N_9698);
or UO_1438 (O_1438,N_9956,N_9590);
or UO_1439 (O_1439,N_9534,N_9857);
nor UO_1440 (O_1440,N_9923,N_9626);
nand UO_1441 (O_1441,N_9646,N_9879);
nor UO_1442 (O_1442,N_9854,N_9984);
and UO_1443 (O_1443,N_9845,N_9573);
and UO_1444 (O_1444,N_9523,N_9655);
or UO_1445 (O_1445,N_9782,N_9786);
nor UO_1446 (O_1446,N_9619,N_9805);
nor UO_1447 (O_1447,N_9963,N_9596);
nand UO_1448 (O_1448,N_9992,N_9697);
nand UO_1449 (O_1449,N_9617,N_9768);
or UO_1450 (O_1450,N_9872,N_9850);
and UO_1451 (O_1451,N_9668,N_9619);
and UO_1452 (O_1452,N_9844,N_9787);
or UO_1453 (O_1453,N_9527,N_9701);
or UO_1454 (O_1454,N_9920,N_9726);
nor UO_1455 (O_1455,N_9781,N_9576);
or UO_1456 (O_1456,N_9741,N_9637);
and UO_1457 (O_1457,N_9600,N_9684);
nor UO_1458 (O_1458,N_9774,N_9933);
and UO_1459 (O_1459,N_9984,N_9786);
nand UO_1460 (O_1460,N_9832,N_9706);
or UO_1461 (O_1461,N_9922,N_9777);
nor UO_1462 (O_1462,N_9836,N_9669);
nand UO_1463 (O_1463,N_9906,N_9505);
nand UO_1464 (O_1464,N_9870,N_9778);
nor UO_1465 (O_1465,N_9859,N_9836);
nor UO_1466 (O_1466,N_9783,N_9677);
or UO_1467 (O_1467,N_9864,N_9822);
and UO_1468 (O_1468,N_9847,N_9954);
xnor UO_1469 (O_1469,N_9717,N_9516);
nand UO_1470 (O_1470,N_9576,N_9646);
and UO_1471 (O_1471,N_9607,N_9905);
or UO_1472 (O_1472,N_9509,N_9738);
or UO_1473 (O_1473,N_9586,N_9977);
or UO_1474 (O_1474,N_9775,N_9716);
nand UO_1475 (O_1475,N_9624,N_9954);
nand UO_1476 (O_1476,N_9677,N_9621);
nor UO_1477 (O_1477,N_9738,N_9539);
nor UO_1478 (O_1478,N_9758,N_9946);
nor UO_1479 (O_1479,N_9997,N_9886);
nor UO_1480 (O_1480,N_9801,N_9550);
or UO_1481 (O_1481,N_9770,N_9848);
nor UO_1482 (O_1482,N_9907,N_9636);
or UO_1483 (O_1483,N_9543,N_9729);
and UO_1484 (O_1484,N_9910,N_9527);
nor UO_1485 (O_1485,N_9692,N_9640);
and UO_1486 (O_1486,N_9577,N_9714);
xor UO_1487 (O_1487,N_9597,N_9685);
nand UO_1488 (O_1488,N_9887,N_9591);
and UO_1489 (O_1489,N_9542,N_9614);
and UO_1490 (O_1490,N_9817,N_9552);
nor UO_1491 (O_1491,N_9664,N_9749);
nor UO_1492 (O_1492,N_9753,N_9542);
nand UO_1493 (O_1493,N_9706,N_9666);
nand UO_1494 (O_1494,N_9657,N_9651);
nor UO_1495 (O_1495,N_9819,N_9812);
nor UO_1496 (O_1496,N_9771,N_9637);
and UO_1497 (O_1497,N_9947,N_9925);
or UO_1498 (O_1498,N_9505,N_9711);
nor UO_1499 (O_1499,N_9506,N_9934);
endmodule