module basic_1000_10000_1500_10_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_533,In_985);
nor U1 (N_1,In_608,In_700);
nand U2 (N_2,In_118,In_768);
or U3 (N_3,In_726,In_70);
or U4 (N_4,In_863,In_143);
and U5 (N_5,In_581,In_442);
nor U6 (N_6,In_363,In_822);
nand U7 (N_7,In_83,In_716);
nor U8 (N_8,In_163,In_114);
nand U9 (N_9,In_634,In_541);
nand U10 (N_10,In_339,In_406);
or U11 (N_11,In_825,In_529);
or U12 (N_12,In_193,In_401);
nand U13 (N_13,In_855,In_523);
nand U14 (N_14,In_928,In_174);
xnor U15 (N_15,In_667,In_140);
nor U16 (N_16,In_84,In_785);
nor U17 (N_17,In_834,In_287);
nand U18 (N_18,In_511,In_970);
nand U19 (N_19,In_666,In_777);
or U20 (N_20,In_325,In_853);
nand U21 (N_21,In_458,In_563);
nand U22 (N_22,In_448,In_914);
nand U23 (N_23,In_3,In_148);
nand U24 (N_24,In_102,In_802);
nand U25 (N_25,In_144,In_191);
nor U26 (N_26,In_490,In_595);
nand U27 (N_27,In_813,In_601);
nand U28 (N_28,In_436,In_322);
or U29 (N_29,In_285,In_43);
or U30 (N_30,In_819,In_49);
nor U31 (N_31,In_44,In_316);
and U32 (N_32,In_94,In_133);
and U33 (N_33,In_350,In_247);
or U34 (N_34,In_284,In_656);
nor U35 (N_35,In_412,In_261);
nand U36 (N_36,In_535,In_121);
nor U37 (N_37,In_223,In_924);
or U38 (N_38,In_299,In_417);
nand U39 (N_39,In_865,In_911);
nor U40 (N_40,In_784,In_388);
or U41 (N_41,In_922,In_661);
nand U42 (N_42,In_781,In_717);
or U43 (N_43,In_642,In_105);
or U44 (N_44,In_727,In_443);
and U45 (N_45,In_127,In_204);
or U46 (N_46,In_951,In_521);
and U47 (N_47,In_167,In_131);
nand U48 (N_48,In_303,In_190);
nor U49 (N_49,In_762,In_984);
and U50 (N_50,In_434,In_475);
and U51 (N_51,In_889,In_923);
nand U52 (N_52,In_444,In_969);
xor U53 (N_53,In_791,In_702);
and U54 (N_54,In_512,In_407);
nand U55 (N_55,In_237,In_671);
xnor U56 (N_56,In_230,In_126);
nor U57 (N_57,In_674,In_383);
and U58 (N_58,In_631,In_706);
nor U59 (N_59,In_35,In_931);
nand U60 (N_60,In_32,In_93);
nor U61 (N_61,In_293,In_73);
and U62 (N_62,In_829,In_108);
nor U63 (N_63,In_977,In_747);
nand U64 (N_64,In_773,In_389);
or U65 (N_65,In_275,In_856);
nor U66 (N_66,In_830,In_809);
or U67 (N_67,In_103,In_740);
xor U68 (N_68,In_846,In_867);
or U69 (N_69,In_679,In_905);
nor U70 (N_70,In_570,In_251);
or U71 (N_71,In_425,In_421);
nor U72 (N_72,In_37,In_390);
and U73 (N_73,In_882,In_898);
or U74 (N_74,In_233,In_927);
and U75 (N_75,In_146,In_359);
or U76 (N_76,In_764,In_67);
and U77 (N_77,In_268,In_173);
and U78 (N_78,In_673,In_722);
nor U79 (N_79,In_637,In_758);
nor U80 (N_80,In_348,In_151);
nand U81 (N_81,In_921,In_956);
nand U82 (N_82,In_116,In_95);
and U83 (N_83,In_866,In_286);
or U84 (N_84,In_155,In_797);
nor U85 (N_85,In_423,In_823);
or U86 (N_86,In_986,In_480);
nor U87 (N_87,In_495,In_987);
or U88 (N_88,In_714,In_918);
or U89 (N_89,In_779,In_685);
or U90 (N_90,In_254,In_119);
nand U91 (N_91,In_464,In_930);
or U92 (N_92,In_467,In_225);
nand U93 (N_93,In_583,In_302);
and U94 (N_94,In_575,In_892);
nand U95 (N_95,In_159,In_690);
nand U96 (N_96,In_368,In_451);
and U97 (N_97,In_701,In_851);
nor U98 (N_98,In_962,In_798);
nor U99 (N_99,In_912,In_399);
xnor U100 (N_100,In_418,In_818);
or U101 (N_101,In_526,In_852);
nor U102 (N_102,In_270,In_677);
and U103 (N_103,In_60,In_196);
and U104 (N_104,In_562,In_874);
or U105 (N_105,In_153,In_248);
nand U106 (N_106,In_547,In_397);
and U107 (N_107,In_184,In_670);
or U108 (N_108,In_925,In_959);
or U109 (N_109,In_371,In_698);
nor U110 (N_110,In_849,In_788);
nor U111 (N_111,In_626,In_554);
and U112 (N_112,In_705,In_946);
xnor U113 (N_113,In_457,In_172);
xor U114 (N_114,In_950,In_933);
and U115 (N_115,In_156,In_945);
nand U116 (N_116,In_440,In_327);
xnor U117 (N_117,In_646,In_619);
or U118 (N_118,In_519,In_691);
nand U119 (N_119,In_944,In_504);
nor U120 (N_120,In_422,In_952);
and U121 (N_121,In_355,In_229);
nor U122 (N_122,In_557,In_871);
and U123 (N_123,In_800,In_621);
nand U124 (N_124,In_662,In_17);
and U125 (N_125,In_139,In_415);
xnor U126 (N_126,In_364,In_873);
xnor U127 (N_127,In_978,In_639);
nand U128 (N_128,In_338,In_112);
nand U129 (N_129,In_789,In_913);
nor U130 (N_130,In_602,In_210);
xnor U131 (N_131,In_844,In_538);
and U132 (N_132,In_376,In_366);
nand U133 (N_133,In_257,In_672);
nand U134 (N_134,In_596,In_328);
nand U135 (N_135,In_697,In_265);
nor U136 (N_136,In_377,In_347);
or U137 (N_137,In_859,In_737);
xnor U138 (N_138,In_72,In_427);
and U139 (N_139,In_232,In_117);
nor U140 (N_140,In_16,In_90);
xnor U141 (N_141,In_576,In_915);
nand U142 (N_142,In_817,In_886);
nand U143 (N_143,In_729,In_298);
or U144 (N_144,In_435,In_708);
nor U145 (N_145,In_658,In_306);
and U146 (N_146,In_836,In_604);
or U147 (N_147,In_326,In_885);
nor U148 (N_148,In_28,In_288);
or U149 (N_149,In_565,In_907);
and U150 (N_150,In_782,In_719);
nand U151 (N_151,In_291,In_197);
nand U152 (N_152,In_130,In_957);
and U153 (N_153,In_409,In_568);
and U154 (N_154,In_725,In_344);
and U155 (N_155,In_982,In_999);
and U156 (N_156,In_372,In_981);
nor U157 (N_157,In_908,In_460);
nand U158 (N_158,In_361,In_175);
and U159 (N_159,In_584,In_99);
nor U160 (N_160,In_431,In_137);
or U161 (N_161,In_125,In_48);
nand U162 (N_162,In_235,In_593);
or U163 (N_163,In_168,In_842);
nand U164 (N_164,In_820,In_215);
or U165 (N_165,In_644,In_980);
nor U166 (N_166,In_553,In_75);
or U167 (N_167,In_578,In_244);
nor U168 (N_168,In_189,In_23);
and U169 (N_169,In_732,In_45);
and U170 (N_170,In_295,In_269);
nand U171 (N_171,In_976,In_241);
or U172 (N_172,In_96,In_466);
and U173 (N_173,In_113,In_157);
xnor U174 (N_174,In_315,In_122);
or U175 (N_175,In_497,In_107);
or U176 (N_176,In_653,In_824);
or U177 (N_177,In_971,In_41);
or U178 (N_178,In_815,In_531);
nor U179 (N_179,In_605,In_57);
and U180 (N_180,In_741,In_66);
nand U181 (N_181,In_854,In_461);
nand U182 (N_182,In_98,In_21);
nand U183 (N_183,In_447,In_895);
and U184 (N_184,In_939,In_365);
or U185 (N_185,In_920,In_394);
and U186 (N_186,In_180,In_899);
or U187 (N_187,In_926,In_445);
xor U188 (N_188,In_884,In_333);
nor U189 (N_189,In_577,In_381);
or U190 (N_190,In_778,In_61);
nand U191 (N_191,In_571,In_686);
nand U192 (N_192,In_810,In_510);
nand U193 (N_193,In_534,In_101);
nor U194 (N_194,In_751,In_524);
or U195 (N_195,In_185,In_280);
or U196 (N_196,In_52,In_580);
and U197 (N_197,In_947,In_478);
nand U198 (N_198,In_900,In_527);
xor U199 (N_199,In_454,In_713);
or U200 (N_200,In_242,In_532);
xor U201 (N_201,In_731,In_763);
and U202 (N_202,In_166,In_165);
and U203 (N_203,In_537,In_841);
nand U204 (N_204,In_195,In_860);
nand U205 (N_205,In_828,In_559);
and U206 (N_206,In_65,In_680);
xnor U207 (N_207,In_398,In_681);
nor U208 (N_208,In_872,In_80);
nor U209 (N_209,In_277,In_152);
or U210 (N_210,In_203,In_879);
nand U211 (N_211,In_0,In_25);
nand U212 (N_212,In_635,In_546);
or U213 (N_213,In_518,In_689);
nand U214 (N_214,In_878,In_160);
and U215 (N_215,In_276,In_134);
and U216 (N_216,In_106,In_755);
xnor U217 (N_217,In_668,In_761);
or U218 (N_218,In_181,In_753);
or U219 (N_219,In_682,In_641);
nand U220 (N_220,In_862,In_238);
or U221 (N_221,In_346,In_20);
nand U222 (N_222,In_452,In_488);
nor U223 (N_223,In_433,In_514);
or U224 (N_224,In_120,In_88);
xnor U225 (N_225,In_963,In_796);
nand U226 (N_226,In_942,In_77);
xor U227 (N_227,In_993,In_733);
nor U228 (N_228,In_588,In_224);
and U229 (N_229,In_539,In_840);
or U230 (N_230,In_356,In_266);
and U231 (N_231,In_19,In_649);
or U232 (N_232,In_470,In_728);
nand U233 (N_233,In_81,In_752);
and U234 (N_234,In_243,In_542);
xor U235 (N_235,In_786,In_730);
nor U236 (N_236,In_556,In_955);
nor U237 (N_237,In_282,In_55);
or U238 (N_238,In_463,In_861);
xnor U239 (N_239,In_551,In_386);
xor U240 (N_240,In_86,In_651);
nor U241 (N_241,In_39,In_622);
nand U242 (N_242,In_10,In_916);
nor U243 (N_243,In_100,In_735);
or U244 (N_244,In_227,In_46);
xnor U245 (N_245,In_484,In_154);
nor U246 (N_246,In_974,In_507);
and U247 (N_247,In_917,In_300);
and U248 (N_248,In_477,In_767);
or U249 (N_249,In_256,In_309);
and U250 (N_250,In_491,In_632);
nor U251 (N_251,In_178,In_489);
or U252 (N_252,In_234,In_612);
nor U253 (N_253,In_206,In_171);
nand U254 (N_254,In_663,In_648);
or U255 (N_255,In_561,In_250);
and U256 (N_256,In_188,In_618);
nand U257 (N_257,In_158,In_142);
xor U258 (N_258,In_236,In_82);
nand U259 (N_259,In_345,In_343);
and U260 (N_260,In_887,In_318);
and U261 (N_261,In_687,In_833);
nand U262 (N_262,In_79,In_506);
nor U263 (N_263,In_370,In_192);
or U264 (N_264,In_441,In_321);
nand U265 (N_265,In_274,In_793);
nor U266 (N_266,In_267,In_483);
and U267 (N_267,In_292,In_164);
or U268 (N_268,In_305,In_501);
nand U269 (N_269,In_645,In_471);
or U270 (N_270,In_948,In_749);
nand U271 (N_271,In_402,In_323);
xnor U272 (N_272,In_76,In_246);
and U273 (N_273,In_995,In_759);
or U274 (N_274,In_487,In_744);
and U275 (N_275,In_597,In_482);
and U276 (N_276,In_240,In_395);
nor U277 (N_277,In_176,In_313);
xor U278 (N_278,In_502,In_904);
and U279 (N_279,In_479,In_994);
nor U280 (N_280,In_330,In_430);
nand U281 (N_281,In_354,In_591);
nor U282 (N_282,In_474,In_432);
or U283 (N_283,In_954,In_69);
and U284 (N_284,In_807,In_249);
nor U285 (N_285,In_770,In_515);
xnor U286 (N_286,In_704,In_972);
nand U287 (N_287,In_426,In_26);
nor U288 (N_288,In_410,In_965);
or U289 (N_289,In_869,In_614);
nor U290 (N_290,In_226,In_929);
nand U291 (N_291,In_647,In_765);
nor U292 (N_292,In_54,In_297);
nor U293 (N_293,In_940,In_549);
and U294 (N_294,In_396,In_179);
nand U295 (N_295,In_989,In_801);
or U296 (N_296,In_736,In_391);
and U297 (N_297,In_845,In_848);
nor U298 (N_298,In_462,In_997);
nor U299 (N_299,In_992,In_745);
nand U300 (N_300,In_31,In_205);
nor U301 (N_301,In_481,In_569);
and U302 (N_302,In_279,In_228);
nand U303 (N_303,In_1,In_558);
nand U304 (N_304,In_358,In_806);
nand U305 (N_305,In_312,In_91);
nand U306 (N_306,In_827,In_499);
nor U307 (N_307,In_200,In_2);
nand U308 (N_308,In_212,In_960);
nand U309 (N_309,In_281,In_494);
and U310 (N_310,In_880,In_587);
and U311 (N_311,In_858,In_572);
and U312 (N_312,In_308,In_528);
and U313 (N_313,In_718,In_403);
or U314 (N_314,In_525,In_721);
and U315 (N_315,In_966,In_803);
nand U316 (N_316,In_617,In_754);
nand U317 (N_317,In_40,In_664);
nor U318 (N_318,In_795,In_351);
nand U319 (N_319,In_564,In_493);
and U320 (N_320,In_630,In_883);
or U321 (N_321,In_162,In_465);
nand U322 (N_322,In_901,In_875);
and U323 (N_323,In_42,In_517);
nor U324 (N_324,In_253,In_574);
and U325 (N_325,In_748,In_307);
nor U326 (N_326,In_688,In_382);
nand U327 (N_327,In_961,In_22);
and U328 (N_328,In_387,In_411);
nand U329 (N_329,In_603,In_790);
nor U330 (N_330,In_897,In_620);
and U331 (N_331,In_420,In_804);
and U332 (N_332,In_566,In_473);
or U333 (N_333,In_115,In_723);
and U334 (N_334,In_336,In_278);
nor U335 (N_335,In_317,In_314);
or U336 (N_336,In_812,In_935);
nor U337 (N_337,In_374,In_509);
nor U338 (N_338,In_699,In_272);
and U339 (N_339,In_530,In_147);
and U340 (N_340,In_949,In_353);
nand U341 (N_341,In_695,In_141);
or U342 (N_342,In_202,In_216);
nand U343 (N_343,In_207,In_742);
nor U344 (N_344,In_676,In_380);
nand U345 (N_345,In_998,In_74);
nor U346 (N_346,In_683,In_6);
nor U347 (N_347,In_934,In_636);
nor U348 (N_348,In_331,In_455);
or U349 (N_349,In_341,In_104);
nor U350 (N_350,In_405,In_638);
nor U351 (N_351,In_821,In_953);
nand U352 (N_352,In_498,In_610);
nand U353 (N_353,In_349,In_832);
and U354 (N_354,In_329,In_27);
nor U355 (N_355,In_289,In_941);
xnor U356 (N_356,In_544,In_124);
nand U357 (N_357,In_675,In_369);
xnor U358 (N_358,In_335,In_89);
and U359 (N_359,In_633,In_5);
or U360 (N_360,In_772,In_585);
or U361 (N_361,In_24,In_18);
and U362 (N_362,In_453,In_332);
or U363 (N_363,In_360,In_36);
nor U364 (N_364,In_352,In_13);
nand U365 (N_365,In_734,In_63);
xor U366 (N_366,In_890,In_550);
nor U367 (N_367,In_110,In_774);
and U368 (N_368,In_492,In_598);
xor U369 (N_369,In_627,In_337);
or U370 (N_370,In_150,In_594);
and U371 (N_371,In_468,In_857);
and U372 (N_372,In_12,In_936);
nand U373 (N_373,In_792,In_47);
xor U374 (N_374,In_643,In_843);
and U375 (N_375,In_177,In_198);
or U376 (N_376,In_161,In_209);
nor U377 (N_377,In_983,In_404);
nand U378 (N_378,In_239,In_231);
nor U379 (N_379,In_222,In_252);
nor U380 (N_380,In_876,In_324);
nor U381 (N_381,In_783,In_486);
or U382 (N_382,In_438,In_59);
or U383 (N_383,In_573,In_320);
nor U384 (N_384,In_893,In_414);
nor U385 (N_385,In_709,In_847);
and U386 (N_386,In_837,In_868);
and U387 (N_387,In_259,In_283);
or U388 (N_388,In_273,In_586);
and U389 (N_389,In_654,In_424);
and U390 (N_390,In_891,In_552);
and U391 (N_391,In_606,In_449);
nor U392 (N_392,In_805,In_794);
and U393 (N_393,In_9,In_780);
or U394 (N_394,In_659,In_787);
nor U395 (N_395,In_296,In_187);
and U396 (N_396,In_92,In_301);
and U397 (N_397,In_870,In_15);
nand U398 (N_398,In_799,In_138);
or U399 (N_399,In_694,In_750);
nand U400 (N_400,In_996,In_657);
and U401 (N_401,In_684,In_712);
and U402 (N_402,In_58,In_186);
nand U403 (N_403,In_446,In_988);
nor U404 (N_404,In_567,In_811);
nand U405 (N_405,In_607,In_469);
nor U406 (N_406,In_932,In_903);
nand U407 (N_407,In_724,In_888);
nand U408 (N_408,In_500,In_29);
or U409 (N_409,In_208,In_937);
or U410 (N_410,In_496,In_145);
nor U411 (N_411,In_199,In_53);
nor U412 (N_412,In_660,In_746);
xnor U413 (N_413,In_375,In_217);
xnor U414 (N_414,In_692,In_958);
nand U415 (N_415,In_715,In_582);
or U416 (N_416,In_373,In_623);
or U417 (N_417,In_943,In_814);
or U418 (N_418,In_290,In_258);
nor U419 (N_419,In_910,In_214);
or U420 (N_420,In_545,In_560);
or U421 (N_421,In_938,In_609);
and U422 (N_422,In_294,In_262);
nand U423 (N_423,In_720,In_776);
nor U424 (N_424,In_419,In_385);
or U425 (N_425,In_964,In_816);
and U426 (N_426,In_766,In_975);
or U427 (N_427,In_808,In_743);
or U428 (N_428,In_973,In_378);
nand U429 (N_429,In_459,In_7);
nor U430 (N_430,In_835,In_864);
nand U431 (N_431,In_640,In_260);
xor U432 (N_432,In_838,In_476);
nand U433 (N_433,In_392,In_87);
nor U434 (N_434,In_194,In_472);
and U435 (N_435,In_652,In_51);
xor U436 (N_436,In_149,In_400);
and U437 (N_437,In_56,In_170);
nand U438 (N_438,In_271,In_760);
or U439 (N_439,In_678,In_428);
xnor U440 (N_440,In_38,In_221);
or U441 (N_441,In_109,In_135);
and U442 (N_442,In_30,In_429);
and U443 (N_443,In_33,In_437);
nor U444 (N_444,In_579,In_132);
or U445 (N_445,In_624,In_78);
or U446 (N_446,In_34,In_169);
xnor U447 (N_447,In_255,In_839);
or U448 (N_448,In_771,In_485);
nor U449 (N_449,In_508,In_979);
and U450 (N_450,In_757,In_555);
or U451 (N_451,In_600,In_909);
nand U452 (N_452,In_967,In_384);
and U453 (N_453,In_362,In_548);
nand U454 (N_454,In_201,In_310);
nand U455 (N_455,In_739,In_503);
or U456 (N_456,In_894,In_71);
and U457 (N_457,In_826,In_357);
nor U458 (N_458,In_613,In_881);
nor U459 (N_459,In_219,In_340);
or U460 (N_460,In_665,In_919);
nand U461 (N_461,In_128,In_218);
and U462 (N_462,In_342,In_703);
or U463 (N_463,In_379,In_906);
nor U464 (N_464,In_334,In_738);
nand U465 (N_465,In_669,In_220);
nor U466 (N_466,In_707,In_245);
nand U467 (N_467,In_616,In_456);
or U468 (N_468,In_393,In_592);
and U469 (N_469,In_50,In_756);
or U470 (N_470,In_136,In_211);
or U471 (N_471,In_4,In_590);
nand U472 (N_472,In_990,In_11);
nor U473 (N_473,In_367,In_611);
and U474 (N_474,In_516,In_628);
or U475 (N_475,In_696,In_64);
and U476 (N_476,In_85,In_693);
xor U477 (N_477,In_769,In_850);
nor U478 (N_478,In_599,In_263);
xnor U479 (N_479,In_319,In_213);
nand U480 (N_480,In_8,In_711);
or U481 (N_481,In_775,In_877);
or U482 (N_482,In_968,In_304);
and U483 (N_483,In_14,In_536);
nor U484 (N_484,In_615,In_413);
nand U485 (N_485,In_183,In_520);
xor U486 (N_486,In_540,In_991);
and U487 (N_487,In_111,In_97);
nand U488 (N_488,In_589,In_543);
nand U489 (N_489,In_902,In_625);
or U490 (N_490,In_311,In_123);
nor U491 (N_491,In_505,In_264);
xnor U492 (N_492,In_439,In_655);
nand U493 (N_493,In_896,In_182);
nor U494 (N_494,In_450,In_710);
or U495 (N_495,In_831,In_522);
and U496 (N_496,In_62,In_629);
and U497 (N_497,In_408,In_513);
or U498 (N_498,In_129,In_650);
nor U499 (N_499,In_68,In_416);
nor U500 (N_500,In_233,In_365);
or U501 (N_501,In_916,In_475);
or U502 (N_502,In_814,In_769);
nor U503 (N_503,In_431,In_522);
nand U504 (N_504,In_731,In_442);
nor U505 (N_505,In_62,In_833);
and U506 (N_506,In_308,In_400);
nor U507 (N_507,In_690,In_514);
or U508 (N_508,In_10,In_900);
and U509 (N_509,In_61,In_878);
or U510 (N_510,In_14,In_254);
and U511 (N_511,In_174,In_452);
or U512 (N_512,In_212,In_973);
nor U513 (N_513,In_376,In_14);
nor U514 (N_514,In_58,In_260);
and U515 (N_515,In_476,In_449);
or U516 (N_516,In_747,In_717);
nor U517 (N_517,In_735,In_168);
and U518 (N_518,In_920,In_852);
nand U519 (N_519,In_981,In_356);
nand U520 (N_520,In_966,In_164);
and U521 (N_521,In_880,In_515);
or U522 (N_522,In_720,In_290);
nor U523 (N_523,In_214,In_977);
and U524 (N_524,In_729,In_907);
and U525 (N_525,In_713,In_155);
nand U526 (N_526,In_893,In_816);
nand U527 (N_527,In_281,In_601);
nor U528 (N_528,In_355,In_70);
xnor U529 (N_529,In_5,In_982);
nor U530 (N_530,In_644,In_913);
nor U531 (N_531,In_433,In_428);
and U532 (N_532,In_117,In_895);
and U533 (N_533,In_795,In_872);
nand U534 (N_534,In_460,In_383);
or U535 (N_535,In_812,In_572);
or U536 (N_536,In_321,In_127);
nand U537 (N_537,In_651,In_951);
nor U538 (N_538,In_278,In_1);
nor U539 (N_539,In_627,In_363);
or U540 (N_540,In_101,In_803);
nor U541 (N_541,In_993,In_937);
and U542 (N_542,In_272,In_982);
or U543 (N_543,In_59,In_826);
nor U544 (N_544,In_58,In_102);
nor U545 (N_545,In_256,In_573);
nand U546 (N_546,In_465,In_60);
nand U547 (N_547,In_20,In_489);
nor U548 (N_548,In_251,In_813);
and U549 (N_549,In_178,In_657);
and U550 (N_550,In_957,In_377);
nand U551 (N_551,In_297,In_198);
nor U552 (N_552,In_403,In_789);
xnor U553 (N_553,In_655,In_86);
nor U554 (N_554,In_537,In_179);
xnor U555 (N_555,In_670,In_866);
xnor U556 (N_556,In_619,In_556);
or U557 (N_557,In_724,In_504);
nand U558 (N_558,In_34,In_566);
and U559 (N_559,In_928,In_251);
nor U560 (N_560,In_356,In_448);
or U561 (N_561,In_765,In_498);
and U562 (N_562,In_109,In_54);
nand U563 (N_563,In_346,In_303);
nand U564 (N_564,In_239,In_876);
and U565 (N_565,In_274,In_694);
or U566 (N_566,In_2,In_929);
xor U567 (N_567,In_956,In_724);
and U568 (N_568,In_33,In_488);
and U569 (N_569,In_293,In_8);
nor U570 (N_570,In_786,In_314);
nor U571 (N_571,In_692,In_820);
nor U572 (N_572,In_330,In_158);
nor U573 (N_573,In_428,In_193);
and U574 (N_574,In_360,In_966);
or U575 (N_575,In_646,In_294);
or U576 (N_576,In_730,In_714);
nand U577 (N_577,In_995,In_672);
nor U578 (N_578,In_171,In_384);
and U579 (N_579,In_673,In_397);
nor U580 (N_580,In_267,In_74);
nor U581 (N_581,In_268,In_829);
and U582 (N_582,In_769,In_948);
xnor U583 (N_583,In_999,In_942);
nand U584 (N_584,In_817,In_599);
and U585 (N_585,In_340,In_789);
xnor U586 (N_586,In_782,In_734);
and U587 (N_587,In_247,In_320);
nor U588 (N_588,In_134,In_8);
nor U589 (N_589,In_336,In_865);
nand U590 (N_590,In_448,In_871);
nand U591 (N_591,In_505,In_416);
nand U592 (N_592,In_753,In_556);
nand U593 (N_593,In_47,In_738);
and U594 (N_594,In_486,In_567);
and U595 (N_595,In_597,In_783);
and U596 (N_596,In_286,In_530);
xnor U597 (N_597,In_533,In_422);
or U598 (N_598,In_217,In_582);
xor U599 (N_599,In_558,In_763);
nand U600 (N_600,In_475,In_938);
nand U601 (N_601,In_980,In_277);
nand U602 (N_602,In_227,In_874);
nand U603 (N_603,In_267,In_531);
and U604 (N_604,In_449,In_940);
and U605 (N_605,In_189,In_312);
nand U606 (N_606,In_963,In_347);
nor U607 (N_607,In_724,In_641);
nor U608 (N_608,In_168,In_986);
nand U609 (N_609,In_103,In_531);
nor U610 (N_610,In_223,In_319);
nand U611 (N_611,In_326,In_586);
or U612 (N_612,In_914,In_28);
nand U613 (N_613,In_800,In_805);
nor U614 (N_614,In_127,In_178);
and U615 (N_615,In_464,In_557);
nor U616 (N_616,In_69,In_733);
and U617 (N_617,In_307,In_515);
xnor U618 (N_618,In_904,In_282);
or U619 (N_619,In_187,In_382);
nor U620 (N_620,In_566,In_576);
nor U621 (N_621,In_37,In_607);
or U622 (N_622,In_443,In_396);
nand U623 (N_623,In_389,In_739);
nand U624 (N_624,In_756,In_873);
nor U625 (N_625,In_269,In_916);
and U626 (N_626,In_632,In_526);
nand U627 (N_627,In_748,In_591);
and U628 (N_628,In_295,In_511);
and U629 (N_629,In_841,In_531);
or U630 (N_630,In_874,In_47);
nor U631 (N_631,In_486,In_813);
and U632 (N_632,In_909,In_698);
nor U633 (N_633,In_844,In_153);
nor U634 (N_634,In_534,In_930);
nor U635 (N_635,In_450,In_28);
nand U636 (N_636,In_974,In_1);
or U637 (N_637,In_425,In_257);
xnor U638 (N_638,In_908,In_854);
or U639 (N_639,In_521,In_362);
and U640 (N_640,In_869,In_941);
xor U641 (N_641,In_729,In_432);
nand U642 (N_642,In_554,In_287);
or U643 (N_643,In_219,In_191);
xnor U644 (N_644,In_846,In_353);
nand U645 (N_645,In_127,In_443);
nand U646 (N_646,In_27,In_927);
nand U647 (N_647,In_907,In_381);
nor U648 (N_648,In_457,In_831);
nor U649 (N_649,In_13,In_725);
nor U650 (N_650,In_530,In_152);
or U651 (N_651,In_233,In_596);
or U652 (N_652,In_167,In_392);
xnor U653 (N_653,In_519,In_936);
nand U654 (N_654,In_193,In_591);
or U655 (N_655,In_966,In_384);
and U656 (N_656,In_425,In_747);
nand U657 (N_657,In_346,In_541);
and U658 (N_658,In_80,In_986);
nand U659 (N_659,In_895,In_642);
xor U660 (N_660,In_443,In_124);
nand U661 (N_661,In_167,In_252);
and U662 (N_662,In_700,In_11);
nor U663 (N_663,In_238,In_660);
nand U664 (N_664,In_468,In_999);
nor U665 (N_665,In_97,In_752);
nor U666 (N_666,In_769,In_983);
or U667 (N_667,In_935,In_986);
or U668 (N_668,In_264,In_441);
nand U669 (N_669,In_537,In_87);
and U670 (N_670,In_236,In_609);
or U671 (N_671,In_133,In_163);
and U672 (N_672,In_351,In_232);
xnor U673 (N_673,In_96,In_745);
or U674 (N_674,In_134,In_696);
nor U675 (N_675,In_172,In_637);
and U676 (N_676,In_968,In_129);
and U677 (N_677,In_696,In_444);
nor U678 (N_678,In_845,In_667);
xnor U679 (N_679,In_518,In_245);
nand U680 (N_680,In_840,In_232);
nand U681 (N_681,In_514,In_369);
and U682 (N_682,In_261,In_577);
nand U683 (N_683,In_211,In_972);
nor U684 (N_684,In_358,In_89);
or U685 (N_685,In_472,In_519);
nor U686 (N_686,In_542,In_683);
and U687 (N_687,In_623,In_839);
nand U688 (N_688,In_825,In_111);
nand U689 (N_689,In_581,In_732);
nand U690 (N_690,In_347,In_289);
or U691 (N_691,In_841,In_589);
xor U692 (N_692,In_447,In_233);
and U693 (N_693,In_63,In_326);
or U694 (N_694,In_858,In_776);
nor U695 (N_695,In_118,In_202);
nor U696 (N_696,In_280,In_635);
and U697 (N_697,In_392,In_920);
nand U698 (N_698,In_122,In_285);
nor U699 (N_699,In_7,In_142);
and U700 (N_700,In_341,In_975);
nor U701 (N_701,In_935,In_101);
or U702 (N_702,In_106,In_35);
nor U703 (N_703,In_656,In_271);
nand U704 (N_704,In_181,In_676);
and U705 (N_705,In_366,In_198);
nand U706 (N_706,In_7,In_468);
and U707 (N_707,In_977,In_856);
nor U708 (N_708,In_997,In_986);
and U709 (N_709,In_893,In_188);
or U710 (N_710,In_965,In_154);
or U711 (N_711,In_802,In_21);
nor U712 (N_712,In_115,In_895);
nor U713 (N_713,In_882,In_223);
or U714 (N_714,In_362,In_146);
nor U715 (N_715,In_852,In_751);
nor U716 (N_716,In_529,In_40);
nor U717 (N_717,In_103,In_156);
nand U718 (N_718,In_422,In_615);
nor U719 (N_719,In_963,In_304);
and U720 (N_720,In_495,In_443);
nand U721 (N_721,In_347,In_664);
and U722 (N_722,In_563,In_483);
and U723 (N_723,In_761,In_170);
nor U724 (N_724,In_779,In_453);
and U725 (N_725,In_266,In_457);
and U726 (N_726,In_285,In_648);
xnor U727 (N_727,In_7,In_589);
nand U728 (N_728,In_642,In_308);
and U729 (N_729,In_599,In_369);
nor U730 (N_730,In_992,In_569);
or U731 (N_731,In_438,In_936);
and U732 (N_732,In_245,In_399);
and U733 (N_733,In_40,In_614);
nor U734 (N_734,In_614,In_336);
nor U735 (N_735,In_50,In_796);
and U736 (N_736,In_120,In_768);
nor U737 (N_737,In_376,In_142);
nor U738 (N_738,In_95,In_363);
nand U739 (N_739,In_731,In_95);
nor U740 (N_740,In_708,In_283);
nand U741 (N_741,In_351,In_989);
and U742 (N_742,In_425,In_740);
and U743 (N_743,In_244,In_368);
or U744 (N_744,In_777,In_416);
xor U745 (N_745,In_763,In_575);
nor U746 (N_746,In_90,In_43);
or U747 (N_747,In_171,In_9);
or U748 (N_748,In_743,In_689);
or U749 (N_749,In_644,In_202);
nor U750 (N_750,In_872,In_265);
nor U751 (N_751,In_336,In_21);
nand U752 (N_752,In_974,In_174);
nand U753 (N_753,In_769,In_306);
nor U754 (N_754,In_216,In_55);
nand U755 (N_755,In_807,In_891);
nand U756 (N_756,In_100,In_347);
nand U757 (N_757,In_394,In_12);
xnor U758 (N_758,In_947,In_276);
or U759 (N_759,In_502,In_62);
nor U760 (N_760,In_876,In_573);
or U761 (N_761,In_73,In_497);
or U762 (N_762,In_27,In_109);
and U763 (N_763,In_356,In_921);
nand U764 (N_764,In_522,In_261);
nand U765 (N_765,In_859,In_366);
nand U766 (N_766,In_754,In_714);
nand U767 (N_767,In_942,In_593);
nand U768 (N_768,In_303,In_568);
nor U769 (N_769,In_533,In_537);
nor U770 (N_770,In_572,In_476);
nand U771 (N_771,In_902,In_224);
xor U772 (N_772,In_709,In_202);
or U773 (N_773,In_516,In_555);
nor U774 (N_774,In_2,In_515);
nor U775 (N_775,In_537,In_575);
nor U776 (N_776,In_295,In_423);
nand U777 (N_777,In_875,In_461);
or U778 (N_778,In_92,In_424);
nor U779 (N_779,In_74,In_111);
or U780 (N_780,In_279,In_608);
nand U781 (N_781,In_500,In_469);
xnor U782 (N_782,In_232,In_948);
xor U783 (N_783,In_859,In_573);
or U784 (N_784,In_65,In_438);
nor U785 (N_785,In_442,In_995);
or U786 (N_786,In_294,In_649);
or U787 (N_787,In_244,In_702);
nand U788 (N_788,In_658,In_665);
nor U789 (N_789,In_376,In_138);
or U790 (N_790,In_590,In_737);
nor U791 (N_791,In_511,In_273);
nor U792 (N_792,In_208,In_758);
or U793 (N_793,In_756,In_512);
xnor U794 (N_794,In_299,In_407);
nor U795 (N_795,In_37,In_78);
nand U796 (N_796,In_143,In_125);
nand U797 (N_797,In_481,In_312);
nor U798 (N_798,In_136,In_909);
or U799 (N_799,In_755,In_464);
nor U800 (N_800,In_986,In_533);
xnor U801 (N_801,In_976,In_884);
or U802 (N_802,In_121,In_983);
nand U803 (N_803,In_71,In_604);
nor U804 (N_804,In_974,In_345);
or U805 (N_805,In_544,In_485);
nand U806 (N_806,In_309,In_749);
and U807 (N_807,In_277,In_311);
xor U808 (N_808,In_10,In_217);
xnor U809 (N_809,In_803,In_494);
nor U810 (N_810,In_397,In_527);
or U811 (N_811,In_483,In_703);
nor U812 (N_812,In_327,In_483);
and U813 (N_813,In_451,In_218);
or U814 (N_814,In_719,In_417);
nor U815 (N_815,In_339,In_676);
nor U816 (N_816,In_376,In_108);
nor U817 (N_817,In_651,In_124);
and U818 (N_818,In_905,In_200);
or U819 (N_819,In_848,In_646);
nand U820 (N_820,In_775,In_792);
and U821 (N_821,In_18,In_572);
and U822 (N_822,In_154,In_941);
xnor U823 (N_823,In_584,In_23);
nand U824 (N_824,In_874,In_422);
nand U825 (N_825,In_945,In_954);
or U826 (N_826,In_635,In_885);
xnor U827 (N_827,In_973,In_189);
and U828 (N_828,In_402,In_536);
nand U829 (N_829,In_736,In_909);
and U830 (N_830,In_964,In_899);
xor U831 (N_831,In_345,In_538);
or U832 (N_832,In_686,In_765);
or U833 (N_833,In_263,In_170);
nor U834 (N_834,In_703,In_806);
or U835 (N_835,In_397,In_926);
or U836 (N_836,In_831,In_426);
and U837 (N_837,In_546,In_489);
nor U838 (N_838,In_303,In_547);
nand U839 (N_839,In_688,In_278);
nor U840 (N_840,In_414,In_477);
and U841 (N_841,In_472,In_827);
and U842 (N_842,In_650,In_965);
and U843 (N_843,In_795,In_483);
nand U844 (N_844,In_210,In_166);
nand U845 (N_845,In_275,In_219);
nor U846 (N_846,In_73,In_628);
nand U847 (N_847,In_809,In_807);
and U848 (N_848,In_666,In_225);
and U849 (N_849,In_955,In_16);
or U850 (N_850,In_661,In_23);
or U851 (N_851,In_994,In_842);
nor U852 (N_852,In_287,In_330);
nand U853 (N_853,In_931,In_171);
and U854 (N_854,In_199,In_174);
xor U855 (N_855,In_230,In_321);
xor U856 (N_856,In_588,In_76);
or U857 (N_857,In_832,In_281);
nand U858 (N_858,In_947,In_436);
nor U859 (N_859,In_756,In_487);
nand U860 (N_860,In_191,In_381);
nand U861 (N_861,In_495,In_945);
nand U862 (N_862,In_263,In_58);
or U863 (N_863,In_928,In_955);
and U864 (N_864,In_909,In_164);
or U865 (N_865,In_596,In_511);
xor U866 (N_866,In_471,In_911);
nand U867 (N_867,In_53,In_220);
or U868 (N_868,In_177,In_404);
xor U869 (N_869,In_777,In_753);
nand U870 (N_870,In_796,In_459);
nand U871 (N_871,In_216,In_569);
nand U872 (N_872,In_582,In_18);
xnor U873 (N_873,In_425,In_128);
or U874 (N_874,In_511,In_200);
nor U875 (N_875,In_200,In_303);
and U876 (N_876,In_59,In_23);
xor U877 (N_877,In_816,In_579);
or U878 (N_878,In_31,In_923);
nor U879 (N_879,In_691,In_298);
nor U880 (N_880,In_497,In_31);
nor U881 (N_881,In_977,In_242);
and U882 (N_882,In_692,In_75);
and U883 (N_883,In_201,In_264);
nand U884 (N_884,In_130,In_826);
nand U885 (N_885,In_669,In_160);
xor U886 (N_886,In_406,In_25);
nand U887 (N_887,In_799,In_76);
or U888 (N_888,In_281,In_651);
nand U889 (N_889,In_824,In_773);
and U890 (N_890,In_670,In_941);
nand U891 (N_891,In_942,In_780);
and U892 (N_892,In_357,In_396);
nand U893 (N_893,In_527,In_237);
nor U894 (N_894,In_874,In_206);
and U895 (N_895,In_463,In_825);
nand U896 (N_896,In_58,In_473);
xnor U897 (N_897,In_601,In_462);
or U898 (N_898,In_127,In_459);
xnor U899 (N_899,In_36,In_639);
nor U900 (N_900,In_429,In_844);
or U901 (N_901,In_847,In_694);
and U902 (N_902,In_900,In_332);
nor U903 (N_903,In_268,In_366);
and U904 (N_904,In_909,In_969);
nor U905 (N_905,In_756,In_922);
nand U906 (N_906,In_823,In_762);
and U907 (N_907,In_511,In_21);
and U908 (N_908,In_704,In_752);
or U909 (N_909,In_319,In_879);
or U910 (N_910,In_344,In_851);
nand U911 (N_911,In_334,In_922);
and U912 (N_912,In_675,In_14);
or U913 (N_913,In_528,In_134);
or U914 (N_914,In_844,In_788);
nand U915 (N_915,In_146,In_629);
xor U916 (N_916,In_815,In_632);
or U917 (N_917,In_677,In_302);
xor U918 (N_918,In_609,In_861);
nor U919 (N_919,In_859,In_77);
nand U920 (N_920,In_789,In_763);
or U921 (N_921,In_585,In_532);
and U922 (N_922,In_934,In_669);
or U923 (N_923,In_315,In_993);
and U924 (N_924,In_615,In_368);
or U925 (N_925,In_713,In_296);
or U926 (N_926,In_996,In_274);
and U927 (N_927,In_189,In_392);
nand U928 (N_928,In_290,In_868);
xnor U929 (N_929,In_877,In_797);
nor U930 (N_930,In_621,In_3);
nor U931 (N_931,In_954,In_756);
or U932 (N_932,In_333,In_476);
or U933 (N_933,In_402,In_384);
or U934 (N_934,In_919,In_167);
nand U935 (N_935,In_184,In_883);
nor U936 (N_936,In_609,In_944);
and U937 (N_937,In_848,In_14);
and U938 (N_938,In_300,In_117);
and U939 (N_939,In_625,In_384);
or U940 (N_940,In_728,In_278);
nor U941 (N_941,In_270,In_790);
and U942 (N_942,In_898,In_839);
nor U943 (N_943,In_686,In_460);
and U944 (N_944,In_101,In_444);
or U945 (N_945,In_729,In_756);
xor U946 (N_946,In_92,In_387);
or U947 (N_947,In_511,In_808);
or U948 (N_948,In_922,In_298);
and U949 (N_949,In_544,In_701);
and U950 (N_950,In_38,In_994);
nor U951 (N_951,In_778,In_526);
nand U952 (N_952,In_29,In_582);
or U953 (N_953,In_567,In_522);
and U954 (N_954,In_466,In_200);
nand U955 (N_955,In_22,In_305);
or U956 (N_956,In_588,In_469);
nor U957 (N_957,In_490,In_735);
or U958 (N_958,In_553,In_463);
nor U959 (N_959,In_925,In_415);
or U960 (N_960,In_599,In_426);
and U961 (N_961,In_77,In_566);
nand U962 (N_962,In_320,In_647);
nor U963 (N_963,In_390,In_910);
xnor U964 (N_964,In_820,In_855);
nand U965 (N_965,In_716,In_28);
nor U966 (N_966,In_573,In_145);
nor U967 (N_967,In_940,In_867);
and U968 (N_968,In_318,In_89);
nand U969 (N_969,In_767,In_34);
and U970 (N_970,In_312,In_791);
nand U971 (N_971,In_818,In_302);
or U972 (N_972,In_214,In_246);
nor U973 (N_973,In_337,In_80);
nor U974 (N_974,In_123,In_932);
nor U975 (N_975,In_349,In_522);
or U976 (N_976,In_977,In_450);
and U977 (N_977,In_842,In_521);
or U978 (N_978,In_914,In_74);
nor U979 (N_979,In_275,In_39);
nor U980 (N_980,In_516,In_737);
and U981 (N_981,In_20,In_195);
nor U982 (N_982,In_101,In_40);
and U983 (N_983,In_412,In_14);
nor U984 (N_984,In_341,In_565);
or U985 (N_985,In_811,In_904);
or U986 (N_986,In_440,In_128);
nor U987 (N_987,In_616,In_444);
nor U988 (N_988,In_335,In_246);
nor U989 (N_989,In_256,In_101);
nand U990 (N_990,In_721,In_494);
nor U991 (N_991,In_390,In_886);
xnor U992 (N_992,In_836,In_858);
nor U993 (N_993,In_172,In_833);
nor U994 (N_994,In_591,In_625);
nand U995 (N_995,In_218,In_857);
and U996 (N_996,In_376,In_868);
xnor U997 (N_997,In_734,In_118);
or U998 (N_998,In_191,In_202);
nand U999 (N_999,In_507,In_773);
xor U1000 (N_1000,N_548,N_857);
and U1001 (N_1001,N_29,N_135);
nand U1002 (N_1002,N_56,N_73);
nand U1003 (N_1003,N_391,N_756);
nand U1004 (N_1004,N_62,N_915);
nor U1005 (N_1005,N_656,N_304);
or U1006 (N_1006,N_723,N_290);
or U1007 (N_1007,N_147,N_587);
or U1008 (N_1008,N_467,N_244);
and U1009 (N_1009,N_591,N_539);
and U1010 (N_1010,N_760,N_767);
or U1011 (N_1011,N_789,N_678);
and U1012 (N_1012,N_832,N_14);
or U1013 (N_1013,N_976,N_117);
nor U1014 (N_1014,N_178,N_521);
nor U1015 (N_1015,N_637,N_714);
or U1016 (N_1016,N_104,N_800);
nor U1017 (N_1017,N_441,N_454);
nand U1018 (N_1018,N_376,N_351);
or U1019 (N_1019,N_442,N_59);
or U1020 (N_1020,N_553,N_269);
nand U1021 (N_1021,N_863,N_680);
nand U1022 (N_1022,N_318,N_958);
nand U1023 (N_1023,N_53,N_823);
and U1024 (N_1024,N_142,N_815);
or U1025 (N_1025,N_191,N_941);
and U1026 (N_1026,N_60,N_416);
nor U1027 (N_1027,N_12,N_150);
xor U1028 (N_1028,N_664,N_72);
or U1029 (N_1029,N_717,N_49);
nand U1030 (N_1030,N_488,N_683);
nor U1031 (N_1031,N_8,N_872);
xnor U1032 (N_1032,N_759,N_295);
and U1033 (N_1033,N_813,N_795);
nor U1034 (N_1034,N_786,N_992);
or U1035 (N_1035,N_445,N_386);
or U1036 (N_1036,N_939,N_688);
and U1037 (N_1037,N_897,N_133);
nor U1038 (N_1038,N_838,N_595);
nor U1039 (N_1039,N_563,N_550);
and U1040 (N_1040,N_93,N_388);
xor U1041 (N_1041,N_564,N_906);
or U1042 (N_1042,N_528,N_115);
and U1043 (N_1043,N_124,N_741);
and U1044 (N_1044,N_242,N_275);
or U1045 (N_1045,N_537,N_729);
nand U1046 (N_1046,N_139,N_165);
and U1047 (N_1047,N_427,N_237);
nand U1048 (N_1048,N_594,N_551);
nand U1049 (N_1049,N_814,N_856);
or U1050 (N_1050,N_903,N_901);
nand U1051 (N_1051,N_109,N_77);
nand U1052 (N_1052,N_288,N_842);
nor U1053 (N_1053,N_702,N_765);
nand U1054 (N_1054,N_468,N_464);
xnor U1055 (N_1055,N_448,N_881);
and U1056 (N_1056,N_605,N_761);
nand U1057 (N_1057,N_90,N_924);
and U1058 (N_1058,N_793,N_758);
nand U1059 (N_1059,N_538,N_422);
nand U1060 (N_1060,N_598,N_990);
xor U1061 (N_1061,N_625,N_470);
or U1062 (N_1062,N_647,N_762);
nand U1063 (N_1063,N_119,N_735);
nor U1064 (N_1064,N_339,N_505);
and U1065 (N_1065,N_65,N_10);
or U1066 (N_1066,N_905,N_151);
nand U1067 (N_1067,N_263,N_884);
or U1068 (N_1068,N_390,N_533);
nor U1069 (N_1069,N_203,N_229);
or U1070 (N_1070,N_943,N_703);
or U1071 (N_1071,N_42,N_718);
nand U1072 (N_1072,N_826,N_329);
nand U1073 (N_1073,N_22,N_102);
nand U1074 (N_1074,N_619,N_541);
and U1075 (N_1075,N_774,N_788);
and U1076 (N_1076,N_525,N_849);
nand U1077 (N_1077,N_790,N_0);
and U1078 (N_1078,N_228,N_27);
and U1079 (N_1079,N_865,N_927);
and U1080 (N_1080,N_699,N_933);
and U1081 (N_1081,N_271,N_577);
xor U1082 (N_1082,N_326,N_11);
nand U1083 (N_1083,N_103,N_477);
or U1084 (N_1084,N_996,N_476);
or U1085 (N_1085,N_571,N_968);
nand U1086 (N_1086,N_300,N_404);
and U1087 (N_1087,N_163,N_211);
and U1088 (N_1088,N_320,N_149);
xnor U1089 (N_1089,N_475,N_784);
nand U1090 (N_1090,N_522,N_753);
and U1091 (N_1091,N_166,N_955);
nor U1092 (N_1092,N_155,N_372);
xor U1093 (N_1093,N_394,N_316);
or U1094 (N_1094,N_89,N_912);
nand U1095 (N_1095,N_67,N_827);
nor U1096 (N_1096,N_640,N_576);
xor U1097 (N_1097,N_169,N_183);
and U1098 (N_1098,N_37,N_164);
nand U1099 (N_1099,N_243,N_942);
nor U1100 (N_1100,N_919,N_91);
nor U1101 (N_1101,N_250,N_979);
nor U1102 (N_1102,N_689,N_172);
xnor U1103 (N_1103,N_822,N_754);
or U1104 (N_1104,N_221,N_825);
nand U1105 (N_1105,N_31,N_218);
nand U1106 (N_1106,N_214,N_978);
nand U1107 (N_1107,N_447,N_877);
nor U1108 (N_1108,N_82,N_929);
and U1109 (N_1109,N_128,N_954);
nand U1110 (N_1110,N_642,N_365);
or U1111 (N_1111,N_504,N_584);
or U1112 (N_1112,N_695,N_395);
or U1113 (N_1113,N_170,N_900);
nand U1114 (N_1114,N_239,N_397);
nand U1115 (N_1115,N_868,N_532);
nor U1116 (N_1116,N_904,N_349);
and U1117 (N_1117,N_592,N_412);
nand U1118 (N_1118,N_808,N_30);
and U1119 (N_1119,N_626,N_489);
nand U1120 (N_1120,N_146,N_371);
nand U1121 (N_1121,N_332,N_763);
and U1122 (N_1122,N_994,N_187);
and U1123 (N_1123,N_101,N_913);
or U1124 (N_1124,N_215,N_463);
xnor U1125 (N_1125,N_852,N_567);
and U1126 (N_1126,N_543,N_330);
and U1127 (N_1127,N_706,N_518);
and U1128 (N_1128,N_226,N_988);
nand U1129 (N_1129,N_141,N_662);
or U1130 (N_1130,N_616,N_583);
and U1131 (N_1131,N_742,N_682);
nor U1132 (N_1132,N_948,N_770);
nand U1133 (N_1133,N_327,N_2);
or U1134 (N_1134,N_274,N_676);
nor U1135 (N_1135,N_831,N_247);
xnor U1136 (N_1136,N_28,N_796);
and U1137 (N_1137,N_579,N_989);
nand U1138 (N_1138,N_323,N_935);
and U1139 (N_1139,N_482,N_993);
nor U1140 (N_1140,N_886,N_156);
and U1141 (N_1141,N_853,N_696);
nand U1142 (N_1142,N_552,N_861);
nand U1143 (N_1143,N_556,N_737);
and U1144 (N_1144,N_660,N_342);
xor U1145 (N_1145,N_544,N_34);
and U1146 (N_1146,N_778,N_658);
nor U1147 (N_1147,N_216,N_435);
and U1148 (N_1148,N_792,N_651);
nor U1149 (N_1149,N_783,N_32);
nand U1150 (N_1150,N_600,N_646);
and U1151 (N_1151,N_833,N_357);
nand U1152 (N_1152,N_889,N_631);
nand U1153 (N_1153,N_570,N_494);
nand U1154 (N_1154,N_190,N_712);
and U1155 (N_1155,N_107,N_423);
and U1156 (N_1156,N_782,N_478);
or U1157 (N_1157,N_455,N_217);
xor U1158 (N_1158,N_755,N_722);
xnor U1159 (N_1159,N_393,N_896);
nor U1160 (N_1160,N_991,N_959);
nor U1161 (N_1161,N_83,N_36);
nor U1162 (N_1162,N_212,N_632);
and U1163 (N_1163,N_433,N_387);
nand U1164 (N_1164,N_108,N_52);
nand U1165 (N_1165,N_286,N_284);
nor U1166 (N_1166,N_343,N_259);
nor U1167 (N_1167,N_716,N_125);
and U1168 (N_1168,N_620,N_78);
nand U1169 (N_1169,N_480,N_310);
or U1170 (N_1170,N_389,N_479);
or U1171 (N_1171,N_398,N_987);
xnor U1172 (N_1172,N_622,N_186);
nand U1173 (N_1173,N_750,N_878);
and U1174 (N_1174,N_909,N_58);
or U1175 (N_1175,N_324,N_44);
or U1176 (N_1176,N_160,N_986);
xor U1177 (N_1177,N_802,N_599);
xor U1178 (N_1178,N_947,N_697);
and U1179 (N_1179,N_261,N_402);
nor U1180 (N_1180,N_490,N_224);
nand U1181 (N_1181,N_174,N_908);
and U1182 (N_1182,N_360,N_985);
or U1183 (N_1183,N_6,N_381);
or U1184 (N_1184,N_265,N_426);
nor U1185 (N_1185,N_569,N_575);
xnor U1186 (N_1186,N_18,N_844);
nor U1187 (N_1187,N_68,N_273);
nor U1188 (N_1188,N_930,N_830);
or U1189 (N_1189,N_719,N_130);
xnor U1190 (N_1190,N_828,N_588);
and U1191 (N_1191,N_775,N_507);
nand U1192 (N_1192,N_154,N_787);
nand U1193 (N_1193,N_998,N_529);
nor U1194 (N_1194,N_366,N_510);
and U1195 (N_1195,N_473,N_196);
nand U1196 (N_1196,N_781,N_33);
and U1197 (N_1197,N_354,N_806);
nor U1198 (N_1198,N_950,N_208);
nand U1199 (N_1199,N_961,N_585);
or U1200 (N_1200,N_740,N_613);
and U1201 (N_1201,N_608,N_644);
and U1202 (N_1202,N_967,N_667);
nor U1203 (N_1203,N_171,N_257);
or U1204 (N_1204,N_399,N_965);
nor U1205 (N_1205,N_421,N_361);
or U1206 (N_1206,N_440,N_565);
xnor U1207 (N_1207,N_406,N_264);
nand U1208 (N_1208,N_668,N_975);
or U1209 (N_1209,N_777,N_66);
nand U1210 (N_1210,N_966,N_715);
and U1211 (N_1211,N_841,N_629);
or U1212 (N_1212,N_276,N_951);
nand U1213 (N_1213,N_508,N_952);
xor U1214 (N_1214,N_450,N_785);
nand U1215 (N_1215,N_894,N_185);
or U1216 (N_1216,N_526,N_299);
nor U1217 (N_1217,N_430,N_859);
nor U1218 (N_1218,N_684,N_545);
nor U1219 (N_1219,N_129,N_285);
and U1220 (N_1220,N_807,N_298);
xnor U1221 (N_1221,N_283,N_341);
xor U1222 (N_1222,N_704,N_385);
nand U1223 (N_1223,N_314,N_674);
nand U1224 (N_1224,N_984,N_296);
nand U1225 (N_1225,N_818,N_400);
nand U1226 (N_1226,N_472,N_606);
nor U1227 (N_1227,N_408,N_997);
nor U1228 (N_1228,N_136,N_574);
or U1229 (N_1229,N_874,N_534);
and U1230 (N_1230,N_168,N_798);
nor U1231 (N_1231,N_921,N_213);
or U1232 (N_1232,N_752,N_309);
xnor U1233 (N_1233,N_438,N_429);
nor U1234 (N_1234,N_500,N_733);
nor U1235 (N_1235,N_971,N_615);
and U1236 (N_1236,N_418,N_691);
nand U1237 (N_1237,N_804,N_559);
xnor U1238 (N_1238,N_414,N_368);
and U1239 (N_1239,N_627,N_801);
nor U1240 (N_1240,N_514,N_636);
and U1241 (N_1241,N_157,N_817);
and U1242 (N_1242,N_493,N_439);
or U1243 (N_1243,N_337,N_13);
nor U1244 (N_1244,N_661,N_35);
nand U1245 (N_1245,N_465,N_140);
xnor U1246 (N_1246,N_883,N_223);
xnor U1247 (N_1247,N_248,N_195);
and U1248 (N_1248,N_340,N_768);
and U1249 (N_1249,N_673,N_612);
nand U1250 (N_1250,N_55,N_824);
nand U1251 (N_1251,N_653,N_969);
xnor U1252 (N_1252,N_106,N_206);
nand U1253 (N_1253,N_291,N_127);
and U1254 (N_1254,N_633,N_312);
nor U1255 (N_1255,N_855,N_654);
nand U1256 (N_1256,N_888,N_317);
nand U1257 (N_1257,N_573,N_847);
nand U1258 (N_1258,N_116,N_222);
and U1259 (N_1259,N_880,N_145);
nand U1260 (N_1260,N_603,N_837);
nand U1261 (N_1261,N_241,N_983);
or U1262 (N_1262,N_84,N_829);
or U1263 (N_1263,N_209,N_225);
nand U1264 (N_1264,N_811,N_384);
nand U1265 (N_1265,N_23,N_280);
nand U1266 (N_1266,N_483,N_512);
or U1267 (N_1267,N_444,N_428);
and U1268 (N_1268,N_363,N_932);
or U1269 (N_1269,N_301,N_374);
nor U1270 (N_1270,N_302,N_590);
nand U1271 (N_1271,N_100,N_461);
xnor U1272 (N_1272,N_893,N_410);
xnor U1273 (N_1273,N_726,N_39);
and U1274 (N_1274,N_803,N_999);
and U1275 (N_1275,N_210,N_916);
nor U1276 (N_1276,N_748,N_144);
nor U1277 (N_1277,N_303,N_415);
or U1278 (N_1278,N_546,N_848);
nand U1279 (N_1279,N_370,N_88);
nand U1280 (N_1280,N_746,N_344);
and U1281 (N_1281,N_918,N_609);
and U1282 (N_1282,N_420,N_542);
nand U1283 (N_1283,N_557,N_845);
nor U1284 (N_1284,N_621,N_405);
and U1285 (N_1285,N_663,N_252);
nand U1286 (N_1286,N_74,N_436);
and U1287 (N_1287,N_131,N_97);
nand U1288 (N_1288,N_492,N_834);
and U1289 (N_1289,N_369,N_45);
nor U1290 (N_1290,N_333,N_452);
nand U1291 (N_1291,N_294,N_7);
or U1292 (N_1292,N_474,N_460);
or U1293 (N_1293,N_75,N_352);
or U1294 (N_1294,N_835,N_64);
and U1295 (N_1295,N_356,N_535);
nor U1296 (N_1296,N_665,N_143);
and U1297 (N_1297,N_272,N_628);
and U1298 (N_1298,N_730,N_392);
and U1299 (N_1299,N_458,N_70);
and U1300 (N_1300,N_380,N_580);
and U1301 (N_1301,N_509,N_597);
nor U1302 (N_1302,N_555,N_953);
or U1303 (N_1303,N_772,N_797);
and U1304 (N_1304,N_655,N_325);
and U1305 (N_1305,N_189,N_315);
xnor U1306 (N_1306,N_527,N_353);
nand U1307 (N_1307,N_523,N_419);
nor U1308 (N_1308,N_890,N_638);
xor U1309 (N_1309,N_589,N_604);
or U1310 (N_1310,N_256,N_554);
nand U1311 (N_1311,N_926,N_558);
or U1312 (N_1312,N_87,N_974);
nand U1313 (N_1313,N_197,N_491);
or U1314 (N_1314,N_277,N_840);
and U1315 (N_1315,N_920,N_113);
or U1316 (N_1316,N_499,N_693);
nand U1317 (N_1317,N_364,N_159);
xnor U1318 (N_1318,N_610,N_724);
and U1319 (N_1319,N_94,N_530);
xor U1320 (N_1320,N_687,N_671);
nand U1321 (N_1321,N_816,N_401);
nor U1322 (N_1322,N_944,N_700);
and U1323 (N_1323,N_586,N_192);
nor U1324 (N_1324,N_9,N_858);
and U1325 (N_1325,N_182,N_17);
or U1326 (N_1326,N_679,N_396);
nand U1327 (N_1327,N_54,N_923);
or U1328 (N_1328,N_885,N_81);
and U1329 (N_1329,N_866,N_549);
xor U1330 (N_1330,N_946,N_431);
nor U1331 (N_1331,N_582,N_378);
or U1332 (N_1332,N_240,N_383);
and U1333 (N_1333,N_648,N_496);
and U1334 (N_1334,N_207,N_980);
and U1335 (N_1335,N_973,N_854);
and U1336 (N_1336,N_536,N_289);
or U1337 (N_1337,N_581,N_238);
xor U1338 (N_1338,N_134,N_268);
xor U1339 (N_1339,N_669,N_233);
and U1340 (N_1340,N_158,N_515);
or U1341 (N_1341,N_873,N_519);
xnor U1342 (N_1342,N_24,N_895);
nand U1343 (N_1343,N_345,N_359);
and U1344 (N_1344,N_805,N_956);
xor U1345 (N_1345,N_776,N_21);
nand U1346 (N_1346,N_891,N_96);
nand U1347 (N_1347,N_922,N_945);
or U1348 (N_1348,N_362,N_227);
xnor U1349 (N_1349,N_281,N_936);
xor U1350 (N_1350,N_278,N_16);
nor U1351 (N_1351,N_111,N_766);
nand U1352 (N_1352,N_307,N_293);
nor U1353 (N_1353,N_623,N_487);
nor U1354 (N_1354,N_120,N_862);
nor U1355 (N_1355,N_411,N_870);
and U1356 (N_1356,N_745,N_670);
nor U1357 (N_1357,N_614,N_1);
nand U1358 (N_1358,N_799,N_358);
or U1359 (N_1359,N_63,N_200);
or U1360 (N_1360,N_749,N_643);
or U1361 (N_1361,N_20,N_602);
and U1362 (N_1362,N_25,N_618);
and U1363 (N_1363,N_328,N_486);
and U1364 (N_1364,N_725,N_520);
nor U1365 (N_1365,N_437,N_409);
nor U1366 (N_1366,N_47,N_728);
or U1367 (N_1367,N_516,N_681);
nand U1368 (N_1368,N_173,N_506);
nor U1369 (N_1369,N_892,N_871);
nor U1370 (N_1370,N_547,N_118);
and U1371 (N_1371,N_709,N_757);
and U1372 (N_1372,N_43,N_262);
or U1373 (N_1373,N_367,N_910);
nor U1374 (N_1374,N_649,N_705);
nand U1375 (N_1375,N_132,N_972);
nor U1376 (N_1376,N_764,N_502);
or U1377 (N_1377,N_403,N_744);
or U1378 (N_1378,N_287,N_161);
nor U1379 (N_1379,N_931,N_449);
nor U1380 (N_1380,N_937,N_692);
and U1381 (N_1381,N_123,N_938);
xnor U1382 (N_1382,N_235,N_319);
nor U1383 (N_1383,N_914,N_675);
nand U1384 (N_1384,N_846,N_561);
and U1385 (N_1385,N_138,N_484);
and U1386 (N_1386,N_940,N_887);
nand U1387 (N_1387,N_666,N_607);
nor U1388 (N_1388,N_672,N_355);
and U1389 (N_1389,N_875,N_220);
nor U1390 (N_1390,N_471,N_198);
and U1391 (N_1391,N_657,N_194);
nor U1392 (N_1392,N_112,N_677);
nand U1393 (N_1393,N_266,N_346);
nor U1394 (N_1394,N_710,N_864);
and U1395 (N_1395,N_466,N_820);
nor U1396 (N_1396,N_377,N_432);
nand U1397 (N_1397,N_179,N_40);
or U1398 (N_1398,N_925,N_902);
nor U1399 (N_1399,N_560,N_611);
nand U1400 (N_1400,N_202,N_167);
and U1401 (N_1401,N_76,N_152);
and U1402 (N_1402,N_180,N_879);
or U1403 (N_1403,N_578,N_201);
nor U1404 (N_1404,N_860,N_635);
and U1405 (N_1405,N_736,N_596);
or U1406 (N_1406,N_511,N_57);
nor U1407 (N_1407,N_572,N_181);
nand U1408 (N_1408,N_524,N_517);
xnor U1409 (N_1409,N_434,N_898);
nor U1410 (N_1410,N_379,N_907);
and U1411 (N_1411,N_199,N_331);
and U1412 (N_1412,N_957,N_462);
nor U1413 (N_1413,N_685,N_251);
and U1414 (N_1414,N_964,N_634);
nor U1415 (N_1415,N_751,N_3);
and U1416 (N_1416,N_779,N_734);
and U1417 (N_1417,N_869,N_279);
xor U1418 (N_1418,N_485,N_249);
nand U1419 (N_1419,N_459,N_836);
xor U1420 (N_1420,N_105,N_26);
or U1421 (N_1421,N_469,N_949);
or U1422 (N_1422,N_46,N_446);
or U1423 (N_1423,N_456,N_443);
or U1424 (N_1424,N_773,N_690);
or U1425 (N_1425,N_92,N_720);
or U1426 (N_1426,N_50,N_601);
nand U1427 (N_1427,N_876,N_641);
xor U1428 (N_1428,N_231,N_413);
and U1429 (N_1429,N_566,N_960);
and U1430 (N_1430,N_95,N_80);
and U1431 (N_1431,N_867,N_457);
nand U1432 (N_1432,N_61,N_253);
xnor U1433 (N_1433,N_407,N_503);
and U1434 (N_1434,N_348,N_375);
or U1435 (N_1435,N_743,N_137);
or U1436 (N_1436,N_48,N_86);
nand U1437 (N_1437,N_246,N_747);
or U1438 (N_1438,N_780,N_122);
or U1439 (N_1439,N_188,N_69);
or U1440 (N_1440,N_843,N_313);
nor U1441 (N_1441,N_711,N_245);
nand U1442 (N_1442,N_267,N_562);
and U1443 (N_1443,N_321,N_513);
nor U1444 (N_1444,N_645,N_51);
and U1445 (N_1445,N_85,N_347);
nand U1446 (N_1446,N_851,N_568);
and U1447 (N_1447,N_707,N_176);
nor U1448 (N_1448,N_821,N_451);
or U1449 (N_1449,N_254,N_305);
and U1450 (N_1450,N_162,N_204);
nand U1451 (N_1451,N_686,N_497);
nand U1452 (N_1452,N_850,N_810);
nor U1453 (N_1453,N_963,N_322);
nor U1454 (N_1454,N_995,N_694);
nand U1455 (N_1455,N_713,N_652);
and U1456 (N_1456,N_977,N_540);
nand U1457 (N_1457,N_701,N_373);
nand U1458 (N_1458,N_899,N_617);
or U1459 (N_1459,N_727,N_19);
nor U1460 (N_1460,N_982,N_424);
xnor U1461 (N_1461,N_205,N_15);
nand U1462 (N_1462,N_624,N_99);
and U1463 (N_1463,N_153,N_981);
nand U1464 (N_1464,N_282,N_350);
nor U1465 (N_1465,N_148,N_481);
or U1466 (N_1466,N_839,N_501);
or U1467 (N_1467,N_98,N_819);
xnor U1468 (N_1468,N_308,N_126);
and U1469 (N_1469,N_769,N_771);
and U1470 (N_1470,N_650,N_739);
nand U1471 (N_1471,N_292,N_794);
xnor U1472 (N_1472,N_928,N_234);
and U1473 (N_1473,N_425,N_639);
and U1474 (N_1474,N_41,N_184);
and U1475 (N_1475,N_219,N_260);
nand U1476 (N_1476,N_230,N_79);
nand U1477 (N_1477,N_232,N_659);
nand U1478 (N_1478,N_708,N_738);
or U1479 (N_1479,N_177,N_382);
xnor U1480 (N_1480,N_882,N_334);
nand U1481 (N_1481,N_453,N_531);
and U1482 (N_1482,N_110,N_721);
or U1483 (N_1483,N_236,N_917);
or U1484 (N_1484,N_114,N_338);
or U1485 (N_1485,N_498,N_5);
and U1486 (N_1486,N_495,N_335);
and U1487 (N_1487,N_731,N_297);
and U1488 (N_1488,N_698,N_336);
nor U1489 (N_1489,N_258,N_630);
xnor U1490 (N_1490,N_270,N_38);
nand U1491 (N_1491,N_306,N_934);
or U1492 (N_1492,N_193,N_809);
nor U1493 (N_1493,N_593,N_121);
nand U1494 (N_1494,N_970,N_255);
nor U1495 (N_1495,N_732,N_175);
nor U1496 (N_1496,N_911,N_962);
xnor U1497 (N_1497,N_812,N_311);
or U1498 (N_1498,N_417,N_791);
and U1499 (N_1499,N_4,N_71);
and U1500 (N_1500,N_930,N_11);
nor U1501 (N_1501,N_472,N_725);
xnor U1502 (N_1502,N_374,N_45);
nand U1503 (N_1503,N_885,N_281);
and U1504 (N_1504,N_945,N_742);
nand U1505 (N_1505,N_496,N_669);
and U1506 (N_1506,N_261,N_408);
or U1507 (N_1507,N_637,N_946);
nor U1508 (N_1508,N_275,N_42);
or U1509 (N_1509,N_822,N_513);
xor U1510 (N_1510,N_699,N_51);
nand U1511 (N_1511,N_292,N_964);
nand U1512 (N_1512,N_788,N_141);
and U1513 (N_1513,N_698,N_692);
and U1514 (N_1514,N_593,N_260);
xnor U1515 (N_1515,N_84,N_116);
nand U1516 (N_1516,N_221,N_292);
nand U1517 (N_1517,N_242,N_713);
nand U1518 (N_1518,N_995,N_337);
and U1519 (N_1519,N_219,N_719);
or U1520 (N_1520,N_647,N_539);
or U1521 (N_1521,N_299,N_866);
nor U1522 (N_1522,N_258,N_773);
or U1523 (N_1523,N_341,N_266);
and U1524 (N_1524,N_846,N_99);
and U1525 (N_1525,N_249,N_623);
or U1526 (N_1526,N_78,N_47);
or U1527 (N_1527,N_261,N_339);
and U1528 (N_1528,N_141,N_490);
nand U1529 (N_1529,N_52,N_43);
nand U1530 (N_1530,N_439,N_854);
nor U1531 (N_1531,N_509,N_129);
nand U1532 (N_1532,N_448,N_239);
nand U1533 (N_1533,N_417,N_885);
nor U1534 (N_1534,N_944,N_768);
nor U1535 (N_1535,N_385,N_578);
xor U1536 (N_1536,N_281,N_471);
or U1537 (N_1537,N_283,N_154);
nand U1538 (N_1538,N_81,N_421);
and U1539 (N_1539,N_249,N_458);
nor U1540 (N_1540,N_740,N_756);
nor U1541 (N_1541,N_106,N_437);
nor U1542 (N_1542,N_118,N_636);
or U1543 (N_1543,N_506,N_451);
and U1544 (N_1544,N_701,N_858);
and U1545 (N_1545,N_621,N_846);
and U1546 (N_1546,N_662,N_980);
nor U1547 (N_1547,N_95,N_251);
nor U1548 (N_1548,N_821,N_801);
xor U1549 (N_1549,N_809,N_276);
and U1550 (N_1550,N_108,N_126);
nand U1551 (N_1551,N_12,N_334);
or U1552 (N_1552,N_281,N_323);
and U1553 (N_1553,N_282,N_935);
or U1554 (N_1554,N_912,N_54);
xor U1555 (N_1555,N_147,N_64);
and U1556 (N_1556,N_260,N_499);
nor U1557 (N_1557,N_937,N_883);
nand U1558 (N_1558,N_324,N_688);
nand U1559 (N_1559,N_338,N_873);
or U1560 (N_1560,N_683,N_556);
and U1561 (N_1561,N_341,N_387);
or U1562 (N_1562,N_824,N_10);
nor U1563 (N_1563,N_852,N_408);
nand U1564 (N_1564,N_592,N_545);
nand U1565 (N_1565,N_226,N_315);
nand U1566 (N_1566,N_673,N_107);
nor U1567 (N_1567,N_542,N_355);
or U1568 (N_1568,N_155,N_552);
nor U1569 (N_1569,N_450,N_955);
nor U1570 (N_1570,N_60,N_575);
and U1571 (N_1571,N_678,N_603);
or U1572 (N_1572,N_560,N_713);
or U1573 (N_1573,N_775,N_70);
xnor U1574 (N_1574,N_820,N_78);
and U1575 (N_1575,N_292,N_447);
and U1576 (N_1576,N_961,N_627);
or U1577 (N_1577,N_69,N_420);
and U1578 (N_1578,N_651,N_920);
nand U1579 (N_1579,N_966,N_857);
nand U1580 (N_1580,N_596,N_527);
nand U1581 (N_1581,N_958,N_933);
and U1582 (N_1582,N_904,N_253);
and U1583 (N_1583,N_263,N_585);
or U1584 (N_1584,N_733,N_344);
and U1585 (N_1585,N_101,N_432);
nand U1586 (N_1586,N_401,N_37);
nor U1587 (N_1587,N_965,N_136);
or U1588 (N_1588,N_189,N_804);
or U1589 (N_1589,N_685,N_650);
nor U1590 (N_1590,N_103,N_133);
nand U1591 (N_1591,N_516,N_952);
nand U1592 (N_1592,N_470,N_908);
nand U1593 (N_1593,N_314,N_184);
xor U1594 (N_1594,N_551,N_682);
nand U1595 (N_1595,N_555,N_119);
or U1596 (N_1596,N_495,N_863);
nand U1597 (N_1597,N_575,N_247);
and U1598 (N_1598,N_774,N_16);
or U1599 (N_1599,N_525,N_299);
nor U1600 (N_1600,N_54,N_470);
and U1601 (N_1601,N_887,N_74);
or U1602 (N_1602,N_732,N_712);
nor U1603 (N_1603,N_909,N_680);
and U1604 (N_1604,N_968,N_13);
or U1605 (N_1605,N_148,N_215);
and U1606 (N_1606,N_363,N_195);
xnor U1607 (N_1607,N_44,N_493);
nor U1608 (N_1608,N_709,N_458);
or U1609 (N_1609,N_614,N_735);
nor U1610 (N_1610,N_306,N_448);
xor U1611 (N_1611,N_64,N_920);
nor U1612 (N_1612,N_91,N_972);
nor U1613 (N_1613,N_240,N_408);
nor U1614 (N_1614,N_668,N_685);
nor U1615 (N_1615,N_170,N_5);
or U1616 (N_1616,N_262,N_152);
nor U1617 (N_1617,N_457,N_763);
or U1618 (N_1618,N_465,N_421);
or U1619 (N_1619,N_53,N_436);
or U1620 (N_1620,N_289,N_648);
or U1621 (N_1621,N_969,N_855);
or U1622 (N_1622,N_462,N_847);
nor U1623 (N_1623,N_515,N_234);
nand U1624 (N_1624,N_742,N_184);
nor U1625 (N_1625,N_618,N_595);
nand U1626 (N_1626,N_928,N_407);
nand U1627 (N_1627,N_598,N_79);
and U1628 (N_1628,N_403,N_181);
xnor U1629 (N_1629,N_777,N_203);
xor U1630 (N_1630,N_630,N_436);
nand U1631 (N_1631,N_533,N_287);
or U1632 (N_1632,N_253,N_848);
or U1633 (N_1633,N_112,N_889);
or U1634 (N_1634,N_533,N_567);
nor U1635 (N_1635,N_892,N_96);
xor U1636 (N_1636,N_402,N_731);
and U1637 (N_1637,N_817,N_991);
nand U1638 (N_1638,N_132,N_968);
or U1639 (N_1639,N_369,N_36);
or U1640 (N_1640,N_681,N_917);
nor U1641 (N_1641,N_235,N_842);
and U1642 (N_1642,N_246,N_992);
and U1643 (N_1643,N_294,N_371);
nor U1644 (N_1644,N_284,N_739);
or U1645 (N_1645,N_653,N_454);
or U1646 (N_1646,N_921,N_113);
nor U1647 (N_1647,N_231,N_903);
or U1648 (N_1648,N_708,N_180);
nand U1649 (N_1649,N_961,N_721);
xor U1650 (N_1650,N_477,N_189);
and U1651 (N_1651,N_864,N_310);
and U1652 (N_1652,N_31,N_755);
nand U1653 (N_1653,N_62,N_343);
xor U1654 (N_1654,N_540,N_32);
xnor U1655 (N_1655,N_148,N_256);
or U1656 (N_1656,N_631,N_778);
nand U1657 (N_1657,N_893,N_939);
nand U1658 (N_1658,N_176,N_368);
nand U1659 (N_1659,N_349,N_268);
xnor U1660 (N_1660,N_61,N_860);
or U1661 (N_1661,N_569,N_117);
nor U1662 (N_1662,N_591,N_199);
nand U1663 (N_1663,N_552,N_575);
or U1664 (N_1664,N_319,N_734);
xnor U1665 (N_1665,N_810,N_318);
and U1666 (N_1666,N_191,N_859);
or U1667 (N_1667,N_6,N_545);
or U1668 (N_1668,N_410,N_370);
nand U1669 (N_1669,N_985,N_770);
nor U1670 (N_1670,N_952,N_528);
or U1671 (N_1671,N_780,N_50);
nor U1672 (N_1672,N_971,N_719);
nor U1673 (N_1673,N_775,N_583);
xor U1674 (N_1674,N_656,N_238);
nand U1675 (N_1675,N_184,N_691);
nand U1676 (N_1676,N_47,N_908);
nor U1677 (N_1677,N_616,N_43);
nand U1678 (N_1678,N_111,N_209);
and U1679 (N_1679,N_853,N_573);
or U1680 (N_1680,N_262,N_242);
and U1681 (N_1681,N_898,N_922);
xnor U1682 (N_1682,N_286,N_974);
or U1683 (N_1683,N_92,N_568);
or U1684 (N_1684,N_148,N_583);
and U1685 (N_1685,N_943,N_404);
nand U1686 (N_1686,N_275,N_411);
nand U1687 (N_1687,N_292,N_928);
nor U1688 (N_1688,N_198,N_589);
nand U1689 (N_1689,N_811,N_480);
nand U1690 (N_1690,N_697,N_795);
and U1691 (N_1691,N_510,N_196);
or U1692 (N_1692,N_909,N_338);
and U1693 (N_1693,N_422,N_162);
xnor U1694 (N_1694,N_131,N_984);
xor U1695 (N_1695,N_86,N_768);
and U1696 (N_1696,N_622,N_300);
or U1697 (N_1697,N_958,N_518);
nand U1698 (N_1698,N_632,N_450);
or U1699 (N_1699,N_749,N_445);
and U1700 (N_1700,N_623,N_61);
nand U1701 (N_1701,N_117,N_340);
nor U1702 (N_1702,N_74,N_557);
and U1703 (N_1703,N_807,N_44);
nand U1704 (N_1704,N_801,N_911);
or U1705 (N_1705,N_954,N_808);
nand U1706 (N_1706,N_27,N_260);
nor U1707 (N_1707,N_43,N_732);
or U1708 (N_1708,N_979,N_283);
or U1709 (N_1709,N_17,N_871);
and U1710 (N_1710,N_823,N_593);
nand U1711 (N_1711,N_544,N_732);
or U1712 (N_1712,N_750,N_856);
and U1713 (N_1713,N_461,N_428);
nor U1714 (N_1714,N_578,N_656);
nand U1715 (N_1715,N_664,N_574);
nand U1716 (N_1716,N_971,N_273);
nor U1717 (N_1717,N_783,N_328);
nand U1718 (N_1718,N_912,N_183);
nand U1719 (N_1719,N_329,N_556);
nor U1720 (N_1720,N_561,N_520);
and U1721 (N_1721,N_382,N_256);
nand U1722 (N_1722,N_376,N_451);
or U1723 (N_1723,N_292,N_799);
nand U1724 (N_1724,N_699,N_817);
nor U1725 (N_1725,N_823,N_397);
nand U1726 (N_1726,N_614,N_434);
or U1727 (N_1727,N_838,N_604);
nand U1728 (N_1728,N_792,N_679);
or U1729 (N_1729,N_577,N_156);
and U1730 (N_1730,N_612,N_907);
or U1731 (N_1731,N_617,N_577);
xnor U1732 (N_1732,N_186,N_344);
nor U1733 (N_1733,N_57,N_829);
or U1734 (N_1734,N_117,N_874);
nand U1735 (N_1735,N_876,N_899);
nor U1736 (N_1736,N_474,N_609);
or U1737 (N_1737,N_320,N_788);
or U1738 (N_1738,N_958,N_319);
nor U1739 (N_1739,N_449,N_735);
and U1740 (N_1740,N_390,N_754);
or U1741 (N_1741,N_39,N_693);
nand U1742 (N_1742,N_146,N_63);
nand U1743 (N_1743,N_38,N_822);
and U1744 (N_1744,N_598,N_364);
nor U1745 (N_1745,N_562,N_598);
and U1746 (N_1746,N_601,N_975);
nand U1747 (N_1747,N_878,N_903);
and U1748 (N_1748,N_416,N_934);
or U1749 (N_1749,N_166,N_807);
xor U1750 (N_1750,N_125,N_832);
and U1751 (N_1751,N_971,N_787);
or U1752 (N_1752,N_113,N_574);
xor U1753 (N_1753,N_978,N_751);
and U1754 (N_1754,N_616,N_177);
nand U1755 (N_1755,N_700,N_959);
or U1756 (N_1756,N_239,N_958);
or U1757 (N_1757,N_968,N_540);
or U1758 (N_1758,N_999,N_906);
nor U1759 (N_1759,N_589,N_557);
or U1760 (N_1760,N_329,N_340);
nand U1761 (N_1761,N_299,N_749);
or U1762 (N_1762,N_653,N_259);
or U1763 (N_1763,N_477,N_524);
and U1764 (N_1764,N_28,N_928);
and U1765 (N_1765,N_809,N_405);
or U1766 (N_1766,N_746,N_686);
nor U1767 (N_1767,N_433,N_760);
xor U1768 (N_1768,N_871,N_488);
nor U1769 (N_1769,N_843,N_458);
and U1770 (N_1770,N_86,N_27);
nor U1771 (N_1771,N_530,N_272);
nand U1772 (N_1772,N_135,N_564);
nor U1773 (N_1773,N_184,N_939);
and U1774 (N_1774,N_796,N_871);
nor U1775 (N_1775,N_868,N_496);
nand U1776 (N_1776,N_873,N_69);
xor U1777 (N_1777,N_628,N_351);
nand U1778 (N_1778,N_32,N_160);
and U1779 (N_1779,N_119,N_941);
or U1780 (N_1780,N_454,N_36);
and U1781 (N_1781,N_872,N_340);
nand U1782 (N_1782,N_129,N_521);
nor U1783 (N_1783,N_891,N_149);
and U1784 (N_1784,N_528,N_472);
and U1785 (N_1785,N_942,N_18);
xor U1786 (N_1786,N_493,N_997);
nand U1787 (N_1787,N_950,N_778);
or U1788 (N_1788,N_500,N_452);
and U1789 (N_1789,N_808,N_619);
xnor U1790 (N_1790,N_439,N_343);
and U1791 (N_1791,N_775,N_231);
and U1792 (N_1792,N_533,N_763);
nor U1793 (N_1793,N_83,N_576);
nand U1794 (N_1794,N_618,N_972);
nor U1795 (N_1795,N_387,N_42);
or U1796 (N_1796,N_430,N_497);
xor U1797 (N_1797,N_71,N_986);
xnor U1798 (N_1798,N_570,N_1);
nand U1799 (N_1799,N_894,N_498);
or U1800 (N_1800,N_644,N_7);
nand U1801 (N_1801,N_904,N_277);
or U1802 (N_1802,N_505,N_566);
and U1803 (N_1803,N_370,N_810);
xor U1804 (N_1804,N_572,N_402);
nand U1805 (N_1805,N_889,N_458);
nand U1806 (N_1806,N_886,N_329);
nand U1807 (N_1807,N_691,N_760);
nand U1808 (N_1808,N_260,N_47);
nand U1809 (N_1809,N_678,N_848);
nand U1810 (N_1810,N_909,N_562);
and U1811 (N_1811,N_924,N_120);
or U1812 (N_1812,N_337,N_916);
nand U1813 (N_1813,N_725,N_942);
nand U1814 (N_1814,N_734,N_895);
or U1815 (N_1815,N_43,N_886);
and U1816 (N_1816,N_751,N_725);
or U1817 (N_1817,N_605,N_885);
or U1818 (N_1818,N_117,N_365);
or U1819 (N_1819,N_351,N_15);
and U1820 (N_1820,N_763,N_557);
and U1821 (N_1821,N_358,N_814);
and U1822 (N_1822,N_160,N_390);
nand U1823 (N_1823,N_478,N_753);
and U1824 (N_1824,N_735,N_634);
nor U1825 (N_1825,N_961,N_548);
nand U1826 (N_1826,N_594,N_870);
and U1827 (N_1827,N_274,N_63);
nand U1828 (N_1828,N_154,N_311);
nand U1829 (N_1829,N_861,N_785);
nand U1830 (N_1830,N_239,N_233);
nor U1831 (N_1831,N_956,N_759);
and U1832 (N_1832,N_442,N_191);
nand U1833 (N_1833,N_756,N_881);
and U1834 (N_1834,N_586,N_45);
nand U1835 (N_1835,N_208,N_640);
or U1836 (N_1836,N_549,N_686);
nand U1837 (N_1837,N_394,N_670);
nand U1838 (N_1838,N_559,N_168);
xor U1839 (N_1839,N_672,N_0);
or U1840 (N_1840,N_229,N_212);
and U1841 (N_1841,N_632,N_553);
nand U1842 (N_1842,N_315,N_385);
and U1843 (N_1843,N_902,N_833);
or U1844 (N_1844,N_146,N_409);
xnor U1845 (N_1845,N_919,N_158);
or U1846 (N_1846,N_841,N_943);
nor U1847 (N_1847,N_526,N_771);
and U1848 (N_1848,N_118,N_914);
nor U1849 (N_1849,N_872,N_175);
nor U1850 (N_1850,N_283,N_604);
or U1851 (N_1851,N_64,N_72);
or U1852 (N_1852,N_611,N_292);
or U1853 (N_1853,N_78,N_506);
or U1854 (N_1854,N_720,N_608);
and U1855 (N_1855,N_491,N_39);
and U1856 (N_1856,N_272,N_196);
nor U1857 (N_1857,N_236,N_771);
and U1858 (N_1858,N_387,N_201);
nand U1859 (N_1859,N_815,N_665);
xnor U1860 (N_1860,N_666,N_80);
or U1861 (N_1861,N_121,N_64);
xor U1862 (N_1862,N_326,N_437);
or U1863 (N_1863,N_520,N_1);
or U1864 (N_1864,N_457,N_849);
nor U1865 (N_1865,N_22,N_67);
nand U1866 (N_1866,N_725,N_501);
or U1867 (N_1867,N_584,N_665);
and U1868 (N_1868,N_599,N_961);
nand U1869 (N_1869,N_835,N_707);
nor U1870 (N_1870,N_956,N_197);
nor U1871 (N_1871,N_566,N_873);
xnor U1872 (N_1872,N_974,N_224);
nand U1873 (N_1873,N_262,N_618);
or U1874 (N_1874,N_446,N_387);
xnor U1875 (N_1875,N_318,N_116);
nand U1876 (N_1876,N_933,N_799);
and U1877 (N_1877,N_329,N_427);
and U1878 (N_1878,N_972,N_216);
nand U1879 (N_1879,N_866,N_385);
or U1880 (N_1880,N_49,N_627);
nand U1881 (N_1881,N_568,N_732);
and U1882 (N_1882,N_979,N_640);
or U1883 (N_1883,N_857,N_528);
or U1884 (N_1884,N_93,N_498);
nand U1885 (N_1885,N_717,N_386);
and U1886 (N_1886,N_111,N_712);
and U1887 (N_1887,N_741,N_993);
and U1888 (N_1888,N_825,N_110);
or U1889 (N_1889,N_689,N_37);
nand U1890 (N_1890,N_656,N_387);
and U1891 (N_1891,N_857,N_994);
nor U1892 (N_1892,N_135,N_500);
or U1893 (N_1893,N_401,N_418);
xnor U1894 (N_1894,N_710,N_338);
or U1895 (N_1895,N_658,N_351);
and U1896 (N_1896,N_169,N_29);
xnor U1897 (N_1897,N_500,N_756);
nand U1898 (N_1898,N_87,N_594);
and U1899 (N_1899,N_881,N_845);
xor U1900 (N_1900,N_451,N_646);
nor U1901 (N_1901,N_72,N_600);
or U1902 (N_1902,N_295,N_625);
nor U1903 (N_1903,N_616,N_755);
nand U1904 (N_1904,N_830,N_577);
and U1905 (N_1905,N_969,N_447);
and U1906 (N_1906,N_439,N_981);
and U1907 (N_1907,N_850,N_516);
and U1908 (N_1908,N_541,N_171);
or U1909 (N_1909,N_136,N_561);
or U1910 (N_1910,N_476,N_810);
nand U1911 (N_1911,N_679,N_168);
and U1912 (N_1912,N_237,N_137);
nand U1913 (N_1913,N_199,N_817);
and U1914 (N_1914,N_45,N_182);
nor U1915 (N_1915,N_452,N_376);
xor U1916 (N_1916,N_607,N_468);
nor U1917 (N_1917,N_99,N_920);
and U1918 (N_1918,N_237,N_81);
nor U1919 (N_1919,N_554,N_26);
or U1920 (N_1920,N_841,N_194);
nor U1921 (N_1921,N_609,N_112);
or U1922 (N_1922,N_56,N_668);
xor U1923 (N_1923,N_6,N_923);
nor U1924 (N_1924,N_403,N_274);
nand U1925 (N_1925,N_548,N_278);
xnor U1926 (N_1926,N_609,N_816);
nand U1927 (N_1927,N_50,N_495);
and U1928 (N_1928,N_446,N_562);
nand U1929 (N_1929,N_70,N_717);
xnor U1930 (N_1930,N_32,N_533);
and U1931 (N_1931,N_866,N_391);
nor U1932 (N_1932,N_164,N_573);
and U1933 (N_1933,N_434,N_68);
and U1934 (N_1934,N_134,N_945);
nor U1935 (N_1935,N_951,N_622);
or U1936 (N_1936,N_547,N_857);
nand U1937 (N_1937,N_653,N_797);
or U1938 (N_1938,N_114,N_854);
xnor U1939 (N_1939,N_339,N_844);
xor U1940 (N_1940,N_353,N_97);
nand U1941 (N_1941,N_138,N_44);
nor U1942 (N_1942,N_942,N_238);
nor U1943 (N_1943,N_269,N_873);
nand U1944 (N_1944,N_654,N_679);
nor U1945 (N_1945,N_904,N_224);
or U1946 (N_1946,N_961,N_808);
and U1947 (N_1947,N_940,N_470);
or U1948 (N_1948,N_642,N_643);
and U1949 (N_1949,N_417,N_373);
and U1950 (N_1950,N_545,N_891);
nand U1951 (N_1951,N_178,N_948);
or U1952 (N_1952,N_135,N_556);
and U1953 (N_1953,N_591,N_258);
nor U1954 (N_1954,N_537,N_954);
or U1955 (N_1955,N_932,N_401);
or U1956 (N_1956,N_402,N_375);
nand U1957 (N_1957,N_310,N_354);
or U1958 (N_1958,N_80,N_34);
or U1959 (N_1959,N_65,N_402);
xnor U1960 (N_1960,N_293,N_862);
and U1961 (N_1961,N_440,N_402);
xnor U1962 (N_1962,N_982,N_603);
nand U1963 (N_1963,N_172,N_596);
nand U1964 (N_1964,N_249,N_64);
and U1965 (N_1965,N_601,N_68);
nand U1966 (N_1966,N_611,N_507);
xor U1967 (N_1967,N_574,N_977);
xnor U1968 (N_1968,N_297,N_710);
nand U1969 (N_1969,N_60,N_745);
xnor U1970 (N_1970,N_722,N_144);
nand U1971 (N_1971,N_914,N_370);
xnor U1972 (N_1972,N_510,N_35);
nand U1973 (N_1973,N_989,N_157);
or U1974 (N_1974,N_415,N_917);
nand U1975 (N_1975,N_544,N_736);
or U1976 (N_1976,N_350,N_235);
nand U1977 (N_1977,N_614,N_491);
or U1978 (N_1978,N_295,N_913);
nor U1979 (N_1979,N_45,N_330);
xor U1980 (N_1980,N_260,N_293);
or U1981 (N_1981,N_730,N_539);
nor U1982 (N_1982,N_243,N_761);
nand U1983 (N_1983,N_153,N_766);
and U1984 (N_1984,N_705,N_29);
nand U1985 (N_1985,N_310,N_116);
and U1986 (N_1986,N_918,N_18);
nor U1987 (N_1987,N_297,N_951);
xnor U1988 (N_1988,N_749,N_443);
or U1989 (N_1989,N_618,N_450);
nor U1990 (N_1990,N_717,N_973);
or U1991 (N_1991,N_486,N_132);
nand U1992 (N_1992,N_762,N_223);
nand U1993 (N_1993,N_112,N_575);
and U1994 (N_1994,N_804,N_269);
nand U1995 (N_1995,N_402,N_973);
nand U1996 (N_1996,N_605,N_688);
nor U1997 (N_1997,N_361,N_934);
or U1998 (N_1998,N_194,N_368);
xnor U1999 (N_1999,N_49,N_705);
and U2000 (N_2000,N_1256,N_1208);
nor U2001 (N_2001,N_1873,N_1967);
and U2002 (N_2002,N_1022,N_1470);
and U2003 (N_2003,N_1935,N_1707);
or U2004 (N_2004,N_1765,N_1174);
or U2005 (N_2005,N_1757,N_1002);
nor U2006 (N_2006,N_1433,N_1004);
nor U2007 (N_2007,N_1098,N_1439);
or U2008 (N_2008,N_1771,N_1729);
nor U2009 (N_2009,N_1352,N_1250);
and U2010 (N_2010,N_1743,N_1849);
nand U2011 (N_2011,N_1346,N_1431);
nor U2012 (N_2012,N_1501,N_1369);
xor U2013 (N_2013,N_1750,N_1337);
xor U2014 (N_2014,N_1238,N_1906);
nand U2015 (N_2015,N_1538,N_1127);
nand U2016 (N_2016,N_1602,N_1522);
nor U2017 (N_2017,N_1770,N_1206);
nand U2018 (N_2018,N_1218,N_1491);
or U2019 (N_2019,N_1359,N_1129);
nand U2020 (N_2020,N_1136,N_1230);
and U2021 (N_2021,N_1490,N_1840);
nand U2022 (N_2022,N_1875,N_1609);
and U2023 (N_2023,N_1778,N_1973);
or U2024 (N_2024,N_1144,N_1692);
or U2025 (N_2025,N_1546,N_1674);
nor U2026 (N_2026,N_1343,N_1299);
nor U2027 (N_2027,N_1656,N_1453);
nor U2028 (N_2028,N_1495,N_1306);
nor U2029 (N_2029,N_1108,N_1442);
or U2030 (N_2030,N_1414,N_1994);
nor U2031 (N_2031,N_1619,N_1769);
xnor U2032 (N_2032,N_1310,N_1460);
and U2033 (N_2033,N_1627,N_1444);
or U2034 (N_2034,N_1662,N_1107);
nor U2035 (N_2035,N_1149,N_1412);
or U2036 (N_2036,N_1160,N_1478);
and U2037 (N_2037,N_1852,N_1457);
xor U2038 (N_2038,N_1008,N_1767);
nor U2039 (N_2039,N_1007,N_1166);
nand U2040 (N_2040,N_1341,N_1394);
or U2041 (N_2041,N_1315,N_1725);
or U2042 (N_2042,N_1361,N_1654);
and U2043 (N_2043,N_1389,N_1625);
or U2044 (N_2044,N_1279,N_1751);
or U2045 (N_2045,N_1589,N_1746);
and U2046 (N_2046,N_1465,N_1115);
xor U2047 (N_2047,N_1664,N_1438);
nor U2048 (N_2048,N_1985,N_1801);
or U2049 (N_2049,N_1698,N_1908);
and U2050 (N_2050,N_1301,N_1533);
or U2051 (N_2051,N_1871,N_1611);
and U2052 (N_2052,N_1259,N_1956);
and U2053 (N_2053,N_1917,N_1185);
xnor U2054 (N_2054,N_1190,N_1135);
or U2055 (N_2055,N_1622,N_1103);
and U2056 (N_2056,N_1752,N_1648);
nor U2057 (N_2057,N_1963,N_1387);
and U2058 (N_2058,N_1949,N_1049);
xnor U2059 (N_2059,N_1035,N_1030);
or U2060 (N_2060,N_1632,N_1061);
xnor U2061 (N_2061,N_1441,N_1362);
and U2062 (N_2062,N_1693,N_1815);
or U2063 (N_2063,N_1477,N_1584);
nor U2064 (N_2064,N_1095,N_1400);
nor U2065 (N_2065,N_1447,N_1694);
nor U2066 (N_2066,N_1506,N_1437);
xnor U2067 (N_2067,N_1381,N_1472);
and U2068 (N_2068,N_1284,N_1086);
and U2069 (N_2069,N_1317,N_1581);
nor U2070 (N_2070,N_1146,N_1088);
nor U2071 (N_2071,N_1678,N_1327);
and U2072 (N_2072,N_1946,N_1225);
nand U2073 (N_2073,N_1111,N_1630);
xnor U2074 (N_2074,N_1766,N_1948);
and U2075 (N_2075,N_1959,N_1455);
or U2076 (N_2076,N_1395,N_1021);
and U2077 (N_2077,N_1233,N_1521);
and U2078 (N_2078,N_1047,N_1684);
xor U2079 (N_2079,N_1267,N_1789);
nor U2080 (N_2080,N_1886,N_1566);
nor U2081 (N_2081,N_1154,N_1303);
or U2082 (N_2082,N_1215,N_1229);
and U2083 (N_2083,N_1704,N_1112);
nor U2084 (N_2084,N_1874,N_1645);
and U2085 (N_2085,N_1762,N_1081);
or U2086 (N_2086,N_1822,N_1682);
and U2087 (N_2087,N_1863,N_1969);
and U2088 (N_2088,N_1717,N_1050);
nor U2089 (N_2089,N_1124,N_1504);
or U2090 (N_2090,N_1554,N_1203);
or U2091 (N_2091,N_1534,N_1624);
nor U2092 (N_2092,N_1335,N_1843);
or U2093 (N_2093,N_1904,N_1170);
xnor U2094 (N_2094,N_1423,N_1205);
nor U2095 (N_2095,N_1309,N_1851);
or U2096 (N_2096,N_1888,N_1520);
nand U2097 (N_2097,N_1248,N_1527);
nand U2098 (N_2098,N_1347,N_1096);
nand U2099 (N_2099,N_1749,N_1151);
nor U2100 (N_2100,N_1861,N_1845);
and U2101 (N_2101,N_1342,N_1125);
nor U2102 (N_2102,N_1688,N_1031);
nand U2103 (N_2103,N_1812,N_1672);
and U2104 (N_2104,N_1014,N_1826);
or U2105 (N_2105,N_1100,N_1739);
nor U2106 (N_2106,N_1721,N_1823);
and U2107 (N_2107,N_1519,N_1076);
and U2108 (N_2108,N_1869,N_1194);
nand U2109 (N_2109,N_1669,N_1041);
and U2110 (N_2110,N_1025,N_1382);
nand U2111 (N_2111,N_1177,N_1407);
nand U2112 (N_2112,N_1690,N_1740);
nor U2113 (N_2113,N_1807,N_1727);
xnor U2114 (N_2114,N_1032,N_1181);
nand U2115 (N_2115,N_1759,N_1307);
nand U2116 (N_2116,N_1422,N_1418);
or U2117 (N_2117,N_1536,N_1958);
or U2118 (N_2118,N_1574,N_1859);
nand U2119 (N_2119,N_1417,N_1493);
and U2120 (N_2120,N_1514,N_1449);
and U2121 (N_2121,N_1420,N_1187);
nor U2122 (N_2122,N_1742,N_1953);
and U2123 (N_2123,N_1432,N_1910);
nor U2124 (N_2124,N_1523,N_1253);
xnor U2125 (N_2125,N_1313,N_1921);
xor U2126 (N_2126,N_1539,N_1551);
and U2127 (N_2127,N_1055,N_1251);
nor U2128 (N_2128,N_1857,N_1406);
and U2129 (N_2129,N_1265,N_1071);
nor U2130 (N_2130,N_1408,N_1780);
xor U2131 (N_2131,N_1641,N_1612);
and U2132 (N_2132,N_1350,N_1810);
xnor U2133 (N_2133,N_1776,N_1065);
or U2134 (N_2134,N_1847,N_1120);
or U2135 (N_2135,N_1800,N_1930);
nand U2136 (N_2136,N_1064,N_1126);
and U2137 (N_2137,N_1834,N_1737);
nor U2138 (N_2138,N_1487,N_1102);
and U2139 (N_2139,N_1312,N_1837);
and U2140 (N_2140,N_1858,N_1099);
nand U2141 (N_2141,N_1074,N_1063);
xnor U2142 (N_2142,N_1164,N_1458);
or U2143 (N_2143,N_1263,N_1344);
or U2144 (N_2144,N_1084,N_1020);
and U2145 (N_2145,N_1603,N_1304);
xor U2146 (N_2146,N_1123,N_1201);
and U2147 (N_2147,N_1221,N_1082);
or U2148 (N_2148,N_1282,N_1555);
or U2149 (N_2149,N_1634,N_1615);
nand U2150 (N_2150,N_1790,N_1816);
or U2151 (N_2151,N_1867,N_1223);
nand U2152 (N_2152,N_1913,N_1971);
nand U2153 (N_2153,N_1119,N_1137);
or U2154 (N_2154,N_1524,N_1349);
or U2155 (N_2155,N_1753,N_1712);
nor U2156 (N_2156,N_1665,N_1792);
nor U2157 (N_2157,N_1821,N_1791);
or U2158 (N_2158,N_1585,N_1512);
and U2159 (N_2159,N_1799,N_1195);
or U2160 (N_2160,N_1133,N_1371);
or U2161 (N_2161,N_1951,N_1802);
or U2162 (N_2162,N_1280,N_1000);
xor U2163 (N_2163,N_1475,N_1827);
nand U2164 (N_2164,N_1864,N_1782);
nand U2165 (N_2165,N_1838,N_1012);
xnor U2166 (N_2166,N_1110,N_1498);
and U2167 (N_2167,N_1582,N_1211);
or U2168 (N_2168,N_1121,N_1842);
or U2169 (N_2169,N_1924,N_1197);
and U2170 (N_2170,N_1204,N_1249);
xnor U2171 (N_2171,N_1375,N_1188);
xnor U2172 (N_2172,N_1401,N_1268);
nand U2173 (N_2173,N_1269,N_1676);
xnor U2174 (N_2174,N_1222,N_1373);
or U2175 (N_2175,N_1345,N_1945);
and U2176 (N_2176,N_1901,N_1464);
nor U2177 (N_2177,N_1097,N_1775);
or U2178 (N_2178,N_1809,N_1768);
and U2179 (N_2179,N_1954,N_1868);
and U2180 (N_2180,N_1636,N_1326);
nor U2181 (N_2181,N_1288,N_1289);
and U2182 (N_2182,N_1034,N_1606);
or U2183 (N_2183,N_1803,N_1518);
and U2184 (N_2184,N_1116,N_1547);
and U2185 (N_2185,N_1793,N_1474);
and U2186 (N_2186,N_1726,N_1605);
nor U2187 (N_2187,N_1062,N_1200);
xnor U2188 (N_2188,N_1754,N_1537);
and U2189 (N_2189,N_1033,N_1733);
nand U2190 (N_2190,N_1080,N_1159);
or U2191 (N_2191,N_1542,N_1109);
nand U2192 (N_2192,N_1923,N_1356);
nand U2193 (N_2193,N_1364,N_1811);
nand U2194 (N_2194,N_1180,N_1883);
or U2195 (N_2195,N_1243,N_1966);
or U2196 (N_2196,N_1899,N_1545);
or U2197 (N_2197,N_1586,N_1054);
xnor U2198 (N_2198,N_1644,N_1716);
nor U2199 (N_2199,N_1492,N_1940);
nor U2200 (N_2200,N_1416,N_1140);
nand U2201 (N_2201,N_1237,N_1068);
xor U2202 (N_2202,N_1597,N_1829);
nand U2203 (N_2203,N_1553,N_1427);
nand U2204 (N_2204,N_1499,N_1330);
and U2205 (N_2205,N_1515,N_1741);
or U2206 (N_2206,N_1898,N_1797);
or U2207 (N_2207,N_1189,N_1629);
nand U2208 (N_2208,N_1244,N_1885);
nand U2209 (N_2209,N_1525,N_1909);
and U2210 (N_2210,N_1747,N_1302);
or U2211 (N_2211,N_1918,N_1430);
nand U2212 (N_2212,N_1220,N_1974);
nand U2213 (N_2213,N_1059,N_1040);
and U2214 (N_2214,N_1419,N_1794);
nor U2215 (N_2215,N_1083,N_1075);
nand U2216 (N_2216,N_1718,N_1604);
nand U2217 (N_2217,N_1227,N_1278);
or U2218 (N_2218,N_1318,N_1755);
nor U2219 (N_2219,N_1657,N_1168);
nand U2220 (N_2220,N_1489,N_1053);
or U2221 (N_2221,N_1101,N_1393);
or U2222 (N_2222,N_1329,N_1198);
nor U2223 (N_2223,N_1176,N_1944);
and U2224 (N_2224,N_1667,N_1943);
and U2225 (N_2225,N_1607,N_1576);
or U2226 (N_2226,N_1919,N_1992);
and U2227 (N_2227,N_1380,N_1640);
nor U2228 (N_2228,N_1922,N_1931);
and U2229 (N_2229,N_1660,N_1179);
or U2230 (N_2230,N_1051,N_1982);
nor U2231 (N_2231,N_1436,N_1916);
and U2232 (N_2232,N_1482,N_1570);
nor U2233 (N_2233,N_1587,N_1153);
and U2234 (N_2234,N_1722,N_1865);
and U2235 (N_2235,N_1675,N_1505);
and U2236 (N_2236,N_1483,N_1714);
nand U2237 (N_2237,N_1556,N_1339);
and U2238 (N_2238,N_1563,N_1798);
xnor U2239 (N_2239,N_1503,N_1937);
xor U2240 (N_2240,N_1896,N_1736);
nor U2241 (N_2241,N_1655,N_1378);
nand U2242 (N_2242,N_1947,N_1145);
xnor U2243 (N_2243,N_1286,N_1273);
and U2244 (N_2244,N_1616,N_1333);
xor U2245 (N_2245,N_1650,N_1087);
nand U2246 (N_2246,N_1009,N_1038);
and U2247 (N_2247,N_1836,N_1724);
and U2248 (N_2248,N_1572,N_1297);
nor U2249 (N_2249,N_1900,N_1013);
and U2250 (N_2250,N_1564,N_1595);
or U2251 (N_2251,N_1132,N_1700);
nor U2252 (N_2252,N_1708,N_1405);
nor U2253 (N_2253,N_1163,N_1072);
nand U2254 (N_2254,N_1348,N_1060);
nand U2255 (N_2255,N_1999,N_1272);
nand U2256 (N_2256,N_1635,N_1252);
or U2257 (N_2257,N_1496,N_1912);
and U2258 (N_2258,N_1575,N_1452);
and U2259 (N_2259,N_1543,N_1182);
or U2260 (N_2260,N_1508,N_1321);
or U2261 (N_2261,N_1148,N_1613);
and U2262 (N_2262,N_1649,N_1036);
nor U2263 (N_2263,N_1365,N_1424);
nand U2264 (N_2264,N_1673,N_1853);
nand U2265 (N_2265,N_1332,N_1239);
xor U2266 (N_2266,N_1633,N_1480);
xor U2267 (N_2267,N_1155,N_1451);
xnor U2268 (N_2268,N_1941,N_1323);
nand U2269 (N_2269,N_1637,N_1653);
or U2270 (N_2270,N_1473,N_1274);
or U2271 (N_2271,N_1016,N_1577);
or U2272 (N_2272,N_1232,N_1774);
or U2273 (N_2273,N_1281,N_1409);
nor U2274 (N_2274,N_1411,N_1830);
nor U2275 (N_2275,N_1976,N_1738);
nor U2276 (N_2276,N_1240,N_1045);
nand U2277 (N_2277,N_1578,N_1659);
nand U2278 (N_2278,N_1705,N_1028);
and U2279 (N_2279,N_1384,N_1787);
nor U2280 (N_2280,N_1017,N_1580);
nand U2281 (N_2281,N_1157,N_1078);
or U2282 (N_2282,N_1980,N_1454);
nor U2283 (N_2283,N_1744,N_1687);
and U2284 (N_2284,N_1298,N_1397);
or U2285 (N_2285,N_1358,N_1271);
or U2286 (N_2286,N_1048,N_1434);
nand U2287 (N_2287,N_1881,N_1894);
nand U2288 (N_2288,N_1311,N_1241);
and U2289 (N_2289,N_1043,N_1996);
and U2290 (N_2290,N_1089,N_1173);
and U2291 (N_2291,N_1535,N_1890);
and U2292 (N_2292,N_1989,N_1706);
nor U2293 (N_2293,N_1510,N_1224);
or U2294 (N_2294,N_1162,N_1446);
nor U2295 (N_2295,N_1711,N_1668);
and U2296 (N_2296,N_1122,N_1820);
and U2297 (N_2297,N_1614,N_1567);
and U2298 (N_2298,N_1024,N_1010);
nor U2299 (N_2299,N_1965,N_1846);
or U2300 (N_2300,N_1351,N_1158);
nor U2301 (N_2301,N_1915,N_1530);
nor U2302 (N_2302,N_1552,N_1319);
nand U2303 (N_2303,N_1178,N_1425);
or U2304 (N_2304,N_1404,N_1236);
nand U2305 (N_2305,N_1294,N_1077);
or U2306 (N_2306,N_1219,N_1628);
and U2307 (N_2307,N_1957,N_1936);
xor U2308 (N_2308,N_1696,N_1114);
or U2309 (N_2309,N_1893,N_1494);
or U2310 (N_2310,N_1529,N_1386);
or U2311 (N_2311,N_1832,N_1476);
xor U2312 (N_2312,N_1841,N_1594);
and U2313 (N_2313,N_1817,N_1818);
xnor U2314 (N_2314,N_1328,N_1388);
or U2315 (N_2315,N_1978,N_1702);
and U2316 (N_2316,N_1283,N_1651);
nor U2317 (N_2317,N_1887,N_1399);
or U2318 (N_2318,N_1593,N_1939);
nand U2319 (N_2319,N_1322,N_1287);
or U2320 (N_2320,N_1517,N_1143);
or U2321 (N_2321,N_1764,N_1044);
and U2322 (N_2322,N_1872,N_1005);
nor U2323 (N_2323,N_1128,N_1091);
xor U2324 (N_2324,N_1292,N_1402);
nor U2325 (N_2325,N_1426,N_1715);
nand U2326 (N_2326,N_1011,N_1573);
xnor U2327 (N_2327,N_1410,N_1104);
nor U2328 (N_2328,N_1652,N_1786);
or U2329 (N_2329,N_1235,N_1903);
xor U2330 (N_2330,N_1262,N_1598);
xor U2331 (N_2331,N_1850,N_1559);
or U2332 (N_2332,N_1760,N_1689);
nor U2333 (N_2333,N_1142,N_1285);
nand U2334 (N_2334,N_1026,N_1516);
nand U2335 (N_2335,N_1316,N_1878);
or U2336 (N_2336,N_1808,N_1734);
and U2337 (N_2337,N_1877,N_1991);
and U2338 (N_2338,N_1952,N_1165);
and U2339 (N_2339,N_1968,N_1376);
nand U2340 (N_2340,N_1459,N_1257);
nor U2341 (N_2341,N_1254,N_1932);
or U2342 (N_2342,N_1709,N_1626);
or U2343 (N_2343,N_1617,N_1920);
nor U2344 (N_2344,N_1828,N_1831);
or U2345 (N_2345,N_1987,N_1497);
and U2346 (N_2346,N_1905,N_1320);
nand U2347 (N_2347,N_1370,N_1993);
nor U2348 (N_2348,N_1981,N_1147);
or U2349 (N_2349,N_1785,N_1979);
xnor U2350 (N_2350,N_1732,N_1781);
nand U2351 (N_2351,N_1368,N_1325);
xnor U2352 (N_2352,N_1367,N_1338);
and U2353 (N_2353,N_1324,N_1073);
nand U2354 (N_2354,N_1085,N_1199);
and U2355 (N_2355,N_1467,N_1977);
and U2356 (N_2356,N_1067,N_1748);
and U2357 (N_2357,N_1105,N_1548);
nand U2358 (N_2358,N_1193,N_1972);
nand U2359 (N_2359,N_1462,N_1308);
nor U2360 (N_2360,N_1879,N_1710);
nand U2361 (N_2361,N_1428,N_1509);
or U2362 (N_2362,N_1139,N_1964);
or U2363 (N_2363,N_1242,N_1621);
nor U2364 (N_2364,N_1363,N_1374);
nand U2365 (N_2365,N_1513,N_1763);
nand U2366 (N_2366,N_1046,N_1860);
or U2367 (N_2367,N_1216,N_1118);
nor U2368 (N_2368,N_1925,N_1862);
and U2369 (N_2369,N_1398,N_1579);
nor U2370 (N_2370,N_1907,N_1006);
nand U2371 (N_2371,N_1596,N_1360);
nand U2372 (N_2372,N_1150,N_1391);
nor U2373 (N_2373,N_1683,N_1599);
nor U2374 (N_2374,N_1027,N_1415);
nand U2375 (N_2375,N_1592,N_1039);
nor U2376 (N_2376,N_1463,N_1019);
or U2377 (N_2377,N_1260,N_1106);
and U2378 (N_2378,N_1531,N_1844);
nor U2379 (N_2379,N_1544,N_1680);
nor U2380 (N_2380,N_1942,N_1549);
nor U2381 (N_2381,N_1069,N_1934);
or U2382 (N_2382,N_1819,N_1113);
nor U2383 (N_2383,N_1336,N_1541);
nor U2384 (N_2384,N_1590,N_1988);
nand U2385 (N_2385,N_1353,N_1562);
nor U2386 (N_2386,N_1591,N_1421);
and U2387 (N_2387,N_1481,N_1403);
or U2388 (N_2388,N_1275,N_1167);
or U2389 (N_2389,N_1234,N_1018);
and U2390 (N_2390,N_1639,N_1507);
or U2391 (N_2391,N_1212,N_1788);
nor U2392 (N_2392,N_1600,N_1719);
nand U2393 (N_2393,N_1192,N_1003);
xnor U2394 (N_2394,N_1731,N_1138);
nor U2395 (N_2395,N_1486,N_1001);
and U2396 (N_2396,N_1565,N_1484);
and U2397 (N_2397,N_1057,N_1247);
nand U2398 (N_2398,N_1855,N_1557);
nand U2399 (N_2399,N_1997,N_1213);
nand U2400 (N_2400,N_1670,N_1784);
nor U2401 (N_2401,N_1183,N_1445);
nand U2402 (N_2402,N_1814,N_1960);
xnor U2403 (N_2403,N_1701,N_1663);
xnor U2404 (N_2404,N_1175,N_1291);
and U2405 (N_2405,N_1300,N_1052);
nand U2406 (N_2406,N_1355,N_1354);
nor U2407 (N_2407,N_1209,N_1290);
or U2408 (N_2408,N_1392,N_1270);
xnor U2409 (N_2409,N_1485,N_1526);
or U2410 (N_2410,N_1642,N_1891);
and U2411 (N_2411,N_1990,N_1671);
or U2412 (N_2412,N_1372,N_1331);
nand U2413 (N_2413,N_1488,N_1502);
or U2414 (N_2414,N_1889,N_1761);
or U2415 (N_2415,N_1647,N_1686);
nand U2416 (N_2416,N_1171,N_1561);
nor U2417 (N_2417,N_1703,N_1443);
or U2418 (N_2418,N_1277,N_1681);
or U2419 (N_2419,N_1390,N_1720);
nor U2420 (N_2420,N_1970,N_1804);
and U2421 (N_2421,N_1450,N_1079);
or U2422 (N_2422,N_1568,N_1833);
nand U2423 (N_2423,N_1479,N_1092);
xor U2424 (N_2424,N_1094,N_1246);
xnor U2425 (N_2425,N_1583,N_1466);
and U2426 (N_2426,N_1884,N_1015);
nand U2427 (N_2427,N_1914,N_1231);
and U2428 (N_2428,N_1334,N_1623);
xor U2429 (N_2429,N_1870,N_1758);
or U2430 (N_2430,N_1255,N_1848);
nand U2431 (N_2431,N_1661,N_1950);
nor U2432 (N_2432,N_1588,N_1679);
nor U2433 (N_2433,N_1245,N_1666);
nand U2434 (N_2434,N_1305,N_1902);
and U2435 (N_2435,N_1835,N_1745);
and U2436 (N_2436,N_1152,N_1995);
and U2437 (N_2437,N_1928,N_1296);
nor U2438 (N_2438,N_1723,N_1824);
xor U2439 (N_2439,N_1134,N_1897);
or U2440 (N_2440,N_1658,N_1066);
nor U2441 (N_2441,N_1610,N_1440);
nand U2442 (N_2442,N_1196,N_1984);
nand U2443 (N_2443,N_1261,N_1880);
nor U2444 (N_2444,N_1396,N_1295);
nand U2445 (N_2445,N_1184,N_1117);
and U2446 (N_2446,N_1938,N_1558);
or U2447 (N_2447,N_1207,N_1866);
or U2448 (N_2448,N_1806,N_1448);
nand U2449 (N_2449,N_1186,N_1456);
nor U2450 (N_2450,N_1461,N_1357);
or U2451 (N_2451,N_1975,N_1379);
xor U2452 (N_2452,N_1214,N_1795);
nor U2453 (N_2453,N_1813,N_1825);
nand U2454 (N_2454,N_1226,N_1856);
and U2455 (N_2455,N_1070,N_1429);
and U2456 (N_2456,N_1413,N_1699);
and U2457 (N_2457,N_1998,N_1735);
nor U2458 (N_2458,N_1773,N_1366);
nand U2459 (N_2459,N_1962,N_1156);
xnor U2460 (N_2460,N_1276,N_1340);
nor U2461 (N_2461,N_1560,N_1037);
or U2462 (N_2462,N_1500,N_1772);
nor U2463 (N_2463,N_1202,N_1228);
or U2464 (N_2464,N_1677,N_1093);
nor U2465 (N_2465,N_1550,N_1532);
xor U2466 (N_2466,N_1839,N_1695);
and U2467 (N_2467,N_1892,N_1029);
xnor U2468 (N_2468,N_1266,N_1023);
nand U2469 (N_2469,N_1796,N_1042);
nor U2470 (N_2470,N_1646,N_1933);
and U2471 (N_2471,N_1377,N_1131);
nor U2472 (N_2472,N_1090,N_1141);
nand U2473 (N_2473,N_1805,N_1697);
and U2474 (N_2474,N_1385,N_1631);
and U2475 (N_2475,N_1471,N_1961);
xor U2476 (N_2476,N_1876,N_1756);
or U2477 (N_2477,N_1638,N_1172);
nor U2478 (N_2478,N_1169,N_1293);
xnor U2479 (N_2479,N_1161,N_1058);
and U2480 (N_2480,N_1777,N_1528);
and U2481 (N_2481,N_1056,N_1468);
or U2482 (N_2482,N_1264,N_1895);
and U2483 (N_2483,N_1783,N_1191);
nor U2484 (N_2484,N_1511,N_1691);
and U2485 (N_2485,N_1469,N_1210);
nand U2486 (N_2486,N_1713,N_1728);
xnor U2487 (N_2487,N_1854,N_1620);
and U2488 (N_2488,N_1730,N_1314);
nor U2489 (N_2489,N_1618,N_1911);
nand U2490 (N_2490,N_1643,N_1435);
or U2491 (N_2491,N_1986,N_1882);
xnor U2492 (N_2492,N_1779,N_1130);
nor U2493 (N_2493,N_1383,N_1217);
nor U2494 (N_2494,N_1258,N_1983);
nand U2495 (N_2495,N_1601,N_1929);
nand U2496 (N_2496,N_1685,N_1927);
nand U2497 (N_2497,N_1955,N_1571);
nand U2498 (N_2498,N_1569,N_1926);
xor U2499 (N_2499,N_1608,N_1540);
xor U2500 (N_2500,N_1240,N_1465);
nor U2501 (N_2501,N_1411,N_1872);
nor U2502 (N_2502,N_1048,N_1987);
nor U2503 (N_2503,N_1230,N_1958);
nor U2504 (N_2504,N_1721,N_1667);
or U2505 (N_2505,N_1707,N_1517);
or U2506 (N_2506,N_1190,N_1301);
or U2507 (N_2507,N_1187,N_1326);
or U2508 (N_2508,N_1120,N_1744);
nand U2509 (N_2509,N_1759,N_1227);
or U2510 (N_2510,N_1798,N_1005);
or U2511 (N_2511,N_1529,N_1108);
nor U2512 (N_2512,N_1713,N_1016);
xor U2513 (N_2513,N_1210,N_1573);
or U2514 (N_2514,N_1034,N_1655);
nand U2515 (N_2515,N_1831,N_1326);
xor U2516 (N_2516,N_1856,N_1367);
nand U2517 (N_2517,N_1668,N_1572);
or U2518 (N_2518,N_1637,N_1205);
and U2519 (N_2519,N_1263,N_1943);
xor U2520 (N_2520,N_1170,N_1837);
nand U2521 (N_2521,N_1799,N_1722);
nor U2522 (N_2522,N_1648,N_1323);
nor U2523 (N_2523,N_1314,N_1951);
or U2524 (N_2524,N_1867,N_1911);
or U2525 (N_2525,N_1432,N_1946);
and U2526 (N_2526,N_1987,N_1761);
nor U2527 (N_2527,N_1174,N_1111);
nand U2528 (N_2528,N_1465,N_1473);
or U2529 (N_2529,N_1739,N_1069);
and U2530 (N_2530,N_1292,N_1267);
or U2531 (N_2531,N_1371,N_1395);
nor U2532 (N_2532,N_1152,N_1596);
or U2533 (N_2533,N_1668,N_1100);
and U2534 (N_2534,N_1389,N_1115);
and U2535 (N_2535,N_1703,N_1647);
or U2536 (N_2536,N_1792,N_1979);
and U2537 (N_2537,N_1016,N_1685);
xnor U2538 (N_2538,N_1105,N_1763);
nand U2539 (N_2539,N_1344,N_1712);
or U2540 (N_2540,N_1688,N_1988);
and U2541 (N_2541,N_1740,N_1866);
nand U2542 (N_2542,N_1475,N_1391);
and U2543 (N_2543,N_1977,N_1083);
nor U2544 (N_2544,N_1579,N_1176);
nand U2545 (N_2545,N_1762,N_1982);
xnor U2546 (N_2546,N_1170,N_1976);
or U2547 (N_2547,N_1950,N_1722);
and U2548 (N_2548,N_1328,N_1534);
or U2549 (N_2549,N_1243,N_1455);
or U2550 (N_2550,N_1782,N_1136);
and U2551 (N_2551,N_1634,N_1834);
and U2552 (N_2552,N_1549,N_1999);
nor U2553 (N_2553,N_1560,N_1513);
nand U2554 (N_2554,N_1059,N_1139);
and U2555 (N_2555,N_1474,N_1175);
xor U2556 (N_2556,N_1818,N_1067);
nor U2557 (N_2557,N_1095,N_1515);
or U2558 (N_2558,N_1335,N_1944);
nor U2559 (N_2559,N_1027,N_1763);
nor U2560 (N_2560,N_1430,N_1532);
nand U2561 (N_2561,N_1551,N_1062);
nor U2562 (N_2562,N_1388,N_1694);
xor U2563 (N_2563,N_1509,N_1091);
nand U2564 (N_2564,N_1158,N_1941);
nor U2565 (N_2565,N_1429,N_1647);
nand U2566 (N_2566,N_1257,N_1773);
and U2567 (N_2567,N_1976,N_1941);
xnor U2568 (N_2568,N_1220,N_1545);
or U2569 (N_2569,N_1259,N_1072);
xor U2570 (N_2570,N_1346,N_1344);
xor U2571 (N_2571,N_1639,N_1279);
nor U2572 (N_2572,N_1239,N_1536);
and U2573 (N_2573,N_1765,N_1684);
nand U2574 (N_2574,N_1940,N_1846);
nor U2575 (N_2575,N_1786,N_1137);
xnor U2576 (N_2576,N_1914,N_1504);
and U2577 (N_2577,N_1019,N_1493);
xnor U2578 (N_2578,N_1130,N_1992);
nand U2579 (N_2579,N_1527,N_1096);
nor U2580 (N_2580,N_1019,N_1104);
and U2581 (N_2581,N_1598,N_1473);
or U2582 (N_2582,N_1163,N_1862);
nand U2583 (N_2583,N_1887,N_1507);
or U2584 (N_2584,N_1971,N_1525);
and U2585 (N_2585,N_1833,N_1383);
nand U2586 (N_2586,N_1230,N_1978);
or U2587 (N_2587,N_1161,N_1614);
and U2588 (N_2588,N_1727,N_1181);
nand U2589 (N_2589,N_1747,N_1872);
nand U2590 (N_2590,N_1848,N_1720);
or U2591 (N_2591,N_1981,N_1640);
nor U2592 (N_2592,N_1394,N_1130);
and U2593 (N_2593,N_1909,N_1811);
nor U2594 (N_2594,N_1285,N_1708);
or U2595 (N_2595,N_1202,N_1854);
nor U2596 (N_2596,N_1360,N_1424);
xor U2597 (N_2597,N_1435,N_1996);
and U2598 (N_2598,N_1015,N_1858);
or U2599 (N_2599,N_1861,N_1050);
nor U2600 (N_2600,N_1099,N_1725);
nand U2601 (N_2601,N_1612,N_1234);
or U2602 (N_2602,N_1819,N_1212);
nor U2603 (N_2603,N_1319,N_1137);
and U2604 (N_2604,N_1386,N_1334);
and U2605 (N_2605,N_1160,N_1125);
or U2606 (N_2606,N_1924,N_1958);
nand U2607 (N_2607,N_1077,N_1883);
xnor U2608 (N_2608,N_1112,N_1213);
xor U2609 (N_2609,N_1564,N_1437);
xnor U2610 (N_2610,N_1740,N_1142);
nand U2611 (N_2611,N_1450,N_1447);
and U2612 (N_2612,N_1394,N_1628);
and U2613 (N_2613,N_1266,N_1619);
nor U2614 (N_2614,N_1114,N_1947);
nor U2615 (N_2615,N_1943,N_1363);
nand U2616 (N_2616,N_1612,N_1281);
xnor U2617 (N_2617,N_1854,N_1527);
nand U2618 (N_2618,N_1758,N_1410);
and U2619 (N_2619,N_1723,N_1095);
xor U2620 (N_2620,N_1706,N_1695);
and U2621 (N_2621,N_1825,N_1019);
nor U2622 (N_2622,N_1623,N_1025);
nand U2623 (N_2623,N_1811,N_1890);
and U2624 (N_2624,N_1118,N_1987);
xnor U2625 (N_2625,N_1964,N_1586);
xor U2626 (N_2626,N_1722,N_1016);
or U2627 (N_2627,N_1590,N_1212);
nor U2628 (N_2628,N_1563,N_1699);
xnor U2629 (N_2629,N_1789,N_1005);
or U2630 (N_2630,N_1749,N_1921);
xor U2631 (N_2631,N_1192,N_1963);
xor U2632 (N_2632,N_1380,N_1578);
xnor U2633 (N_2633,N_1048,N_1610);
and U2634 (N_2634,N_1602,N_1642);
xor U2635 (N_2635,N_1774,N_1443);
nor U2636 (N_2636,N_1200,N_1740);
or U2637 (N_2637,N_1499,N_1324);
and U2638 (N_2638,N_1001,N_1624);
and U2639 (N_2639,N_1996,N_1323);
and U2640 (N_2640,N_1600,N_1898);
nor U2641 (N_2641,N_1053,N_1238);
or U2642 (N_2642,N_1854,N_1520);
and U2643 (N_2643,N_1480,N_1941);
and U2644 (N_2644,N_1386,N_1548);
nor U2645 (N_2645,N_1223,N_1264);
and U2646 (N_2646,N_1180,N_1035);
nor U2647 (N_2647,N_1451,N_1312);
nand U2648 (N_2648,N_1086,N_1819);
nand U2649 (N_2649,N_1293,N_1398);
and U2650 (N_2650,N_1931,N_1762);
nor U2651 (N_2651,N_1563,N_1452);
and U2652 (N_2652,N_1071,N_1795);
xnor U2653 (N_2653,N_1876,N_1411);
nand U2654 (N_2654,N_1511,N_1800);
or U2655 (N_2655,N_1303,N_1029);
and U2656 (N_2656,N_1499,N_1125);
nor U2657 (N_2657,N_1307,N_1980);
or U2658 (N_2658,N_1664,N_1210);
or U2659 (N_2659,N_1050,N_1414);
xnor U2660 (N_2660,N_1260,N_1576);
or U2661 (N_2661,N_1150,N_1506);
xor U2662 (N_2662,N_1576,N_1773);
and U2663 (N_2663,N_1516,N_1877);
or U2664 (N_2664,N_1431,N_1881);
or U2665 (N_2665,N_1776,N_1538);
and U2666 (N_2666,N_1565,N_1642);
xor U2667 (N_2667,N_1902,N_1887);
and U2668 (N_2668,N_1988,N_1236);
nor U2669 (N_2669,N_1241,N_1011);
nand U2670 (N_2670,N_1907,N_1583);
nand U2671 (N_2671,N_1095,N_1689);
or U2672 (N_2672,N_1066,N_1309);
xor U2673 (N_2673,N_1665,N_1830);
or U2674 (N_2674,N_1349,N_1412);
or U2675 (N_2675,N_1608,N_1024);
nand U2676 (N_2676,N_1829,N_1683);
nand U2677 (N_2677,N_1307,N_1594);
nor U2678 (N_2678,N_1650,N_1661);
nand U2679 (N_2679,N_1571,N_1715);
nor U2680 (N_2680,N_1992,N_1873);
nor U2681 (N_2681,N_1073,N_1351);
nor U2682 (N_2682,N_1195,N_1845);
nand U2683 (N_2683,N_1938,N_1175);
xor U2684 (N_2684,N_1326,N_1433);
or U2685 (N_2685,N_1965,N_1851);
nand U2686 (N_2686,N_1698,N_1428);
or U2687 (N_2687,N_1776,N_1237);
nand U2688 (N_2688,N_1074,N_1278);
nand U2689 (N_2689,N_1471,N_1695);
nand U2690 (N_2690,N_1057,N_1774);
nor U2691 (N_2691,N_1573,N_1805);
nand U2692 (N_2692,N_1755,N_1107);
and U2693 (N_2693,N_1085,N_1042);
nand U2694 (N_2694,N_1601,N_1678);
nand U2695 (N_2695,N_1345,N_1750);
nand U2696 (N_2696,N_1826,N_1200);
nor U2697 (N_2697,N_1720,N_1172);
xnor U2698 (N_2698,N_1001,N_1691);
nand U2699 (N_2699,N_1037,N_1167);
xnor U2700 (N_2700,N_1253,N_1640);
nand U2701 (N_2701,N_1545,N_1020);
nand U2702 (N_2702,N_1125,N_1576);
xnor U2703 (N_2703,N_1444,N_1528);
or U2704 (N_2704,N_1785,N_1103);
and U2705 (N_2705,N_1907,N_1655);
xnor U2706 (N_2706,N_1031,N_1829);
or U2707 (N_2707,N_1043,N_1084);
and U2708 (N_2708,N_1258,N_1522);
nor U2709 (N_2709,N_1774,N_1463);
nand U2710 (N_2710,N_1488,N_1627);
xor U2711 (N_2711,N_1192,N_1527);
and U2712 (N_2712,N_1273,N_1767);
xor U2713 (N_2713,N_1590,N_1181);
or U2714 (N_2714,N_1402,N_1646);
xnor U2715 (N_2715,N_1152,N_1085);
nand U2716 (N_2716,N_1359,N_1056);
xor U2717 (N_2717,N_1622,N_1958);
or U2718 (N_2718,N_1206,N_1091);
nor U2719 (N_2719,N_1210,N_1075);
and U2720 (N_2720,N_1706,N_1749);
and U2721 (N_2721,N_1832,N_1715);
and U2722 (N_2722,N_1273,N_1029);
nor U2723 (N_2723,N_1226,N_1526);
and U2724 (N_2724,N_1720,N_1624);
and U2725 (N_2725,N_1700,N_1346);
or U2726 (N_2726,N_1391,N_1006);
xnor U2727 (N_2727,N_1337,N_1763);
or U2728 (N_2728,N_1403,N_1494);
nor U2729 (N_2729,N_1651,N_1317);
xnor U2730 (N_2730,N_1509,N_1169);
nor U2731 (N_2731,N_1161,N_1423);
xnor U2732 (N_2732,N_1158,N_1042);
nand U2733 (N_2733,N_1003,N_1580);
and U2734 (N_2734,N_1117,N_1293);
nor U2735 (N_2735,N_1844,N_1065);
nand U2736 (N_2736,N_1621,N_1081);
xnor U2737 (N_2737,N_1115,N_1930);
xnor U2738 (N_2738,N_1920,N_1625);
or U2739 (N_2739,N_1852,N_1972);
xor U2740 (N_2740,N_1375,N_1662);
nand U2741 (N_2741,N_1286,N_1957);
and U2742 (N_2742,N_1590,N_1335);
nand U2743 (N_2743,N_1216,N_1458);
nor U2744 (N_2744,N_1729,N_1827);
nand U2745 (N_2745,N_1893,N_1377);
nand U2746 (N_2746,N_1135,N_1787);
nand U2747 (N_2747,N_1548,N_1949);
and U2748 (N_2748,N_1911,N_1966);
nand U2749 (N_2749,N_1504,N_1408);
nand U2750 (N_2750,N_1702,N_1809);
or U2751 (N_2751,N_1825,N_1982);
or U2752 (N_2752,N_1999,N_1910);
and U2753 (N_2753,N_1590,N_1357);
and U2754 (N_2754,N_1342,N_1312);
nor U2755 (N_2755,N_1556,N_1330);
nand U2756 (N_2756,N_1384,N_1847);
and U2757 (N_2757,N_1296,N_1104);
or U2758 (N_2758,N_1341,N_1238);
nand U2759 (N_2759,N_1700,N_1654);
and U2760 (N_2760,N_1766,N_1730);
nor U2761 (N_2761,N_1737,N_1731);
nor U2762 (N_2762,N_1508,N_1985);
nor U2763 (N_2763,N_1080,N_1192);
nor U2764 (N_2764,N_1292,N_1509);
nand U2765 (N_2765,N_1628,N_1870);
or U2766 (N_2766,N_1771,N_1609);
nor U2767 (N_2767,N_1093,N_1199);
nand U2768 (N_2768,N_1356,N_1799);
and U2769 (N_2769,N_1779,N_1471);
or U2770 (N_2770,N_1949,N_1671);
nor U2771 (N_2771,N_1748,N_1516);
xor U2772 (N_2772,N_1550,N_1135);
xor U2773 (N_2773,N_1475,N_1351);
or U2774 (N_2774,N_1938,N_1266);
or U2775 (N_2775,N_1014,N_1047);
nor U2776 (N_2776,N_1141,N_1028);
and U2777 (N_2777,N_1723,N_1308);
nor U2778 (N_2778,N_1126,N_1754);
and U2779 (N_2779,N_1916,N_1281);
xnor U2780 (N_2780,N_1344,N_1026);
nor U2781 (N_2781,N_1574,N_1218);
or U2782 (N_2782,N_1693,N_1107);
or U2783 (N_2783,N_1089,N_1662);
or U2784 (N_2784,N_1800,N_1404);
and U2785 (N_2785,N_1225,N_1681);
or U2786 (N_2786,N_1906,N_1455);
xor U2787 (N_2787,N_1241,N_1893);
and U2788 (N_2788,N_1631,N_1623);
nand U2789 (N_2789,N_1302,N_1390);
nor U2790 (N_2790,N_1372,N_1610);
nand U2791 (N_2791,N_1349,N_1997);
and U2792 (N_2792,N_1658,N_1530);
or U2793 (N_2793,N_1174,N_1951);
xnor U2794 (N_2794,N_1853,N_1772);
and U2795 (N_2795,N_1858,N_1256);
and U2796 (N_2796,N_1208,N_1978);
and U2797 (N_2797,N_1854,N_1548);
nor U2798 (N_2798,N_1573,N_1374);
or U2799 (N_2799,N_1396,N_1592);
and U2800 (N_2800,N_1809,N_1751);
xor U2801 (N_2801,N_1366,N_1271);
or U2802 (N_2802,N_1740,N_1581);
and U2803 (N_2803,N_1971,N_1793);
xor U2804 (N_2804,N_1922,N_1722);
xor U2805 (N_2805,N_1204,N_1197);
nor U2806 (N_2806,N_1233,N_1143);
nand U2807 (N_2807,N_1006,N_1560);
and U2808 (N_2808,N_1557,N_1537);
nor U2809 (N_2809,N_1827,N_1272);
or U2810 (N_2810,N_1695,N_1147);
nand U2811 (N_2811,N_1858,N_1322);
nor U2812 (N_2812,N_1782,N_1645);
nor U2813 (N_2813,N_1626,N_1054);
nor U2814 (N_2814,N_1376,N_1853);
nand U2815 (N_2815,N_1095,N_1757);
or U2816 (N_2816,N_1061,N_1780);
nor U2817 (N_2817,N_1427,N_1504);
nor U2818 (N_2818,N_1727,N_1629);
or U2819 (N_2819,N_1444,N_1743);
and U2820 (N_2820,N_1892,N_1306);
xor U2821 (N_2821,N_1028,N_1591);
nor U2822 (N_2822,N_1991,N_1360);
nor U2823 (N_2823,N_1011,N_1064);
nor U2824 (N_2824,N_1709,N_1750);
nand U2825 (N_2825,N_1073,N_1269);
or U2826 (N_2826,N_1250,N_1133);
and U2827 (N_2827,N_1842,N_1706);
and U2828 (N_2828,N_1485,N_1127);
nand U2829 (N_2829,N_1190,N_1255);
or U2830 (N_2830,N_1567,N_1529);
nor U2831 (N_2831,N_1871,N_1161);
and U2832 (N_2832,N_1766,N_1820);
nor U2833 (N_2833,N_1087,N_1978);
and U2834 (N_2834,N_1050,N_1531);
or U2835 (N_2835,N_1703,N_1833);
nor U2836 (N_2836,N_1044,N_1721);
and U2837 (N_2837,N_1379,N_1511);
or U2838 (N_2838,N_1460,N_1042);
nand U2839 (N_2839,N_1750,N_1615);
nor U2840 (N_2840,N_1797,N_1478);
nor U2841 (N_2841,N_1107,N_1733);
nor U2842 (N_2842,N_1636,N_1620);
nor U2843 (N_2843,N_1615,N_1909);
nor U2844 (N_2844,N_1443,N_1785);
nand U2845 (N_2845,N_1148,N_1568);
and U2846 (N_2846,N_1652,N_1590);
nor U2847 (N_2847,N_1219,N_1350);
and U2848 (N_2848,N_1880,N_1041);
or U2849 (N_2849,N_1131,N_1087);
nor U2850 (N_2850,N_1507,N_1572);
nand U2851 (N_2851,N_1264,N_1289);
or U2852 (N_2852,N_1644,N_1596);
nor U2853 (N_2853,N_1817,N_1533);
or U2854 (N_2854,N_1454,N_1671);
nand U2855 (N_2855,N_1799,N_1826);
or U2856 (N_2856,N_1535,N_1693);
and U2857 (N_2857,N_1140,N_1191);
and U2858 (N_2858,N_1125,N_1187);
and U2859 (N_2859,N_1008,N_1319);
or U2860 (N_2860,N_1411,N_1796);
nand U2861 (N_2861,N_1014,N_1326);
or U2862 (N_2862,N_1802,N_1517);
or U2863 (N_2863,N_1748,N_1066);
xnor U2864 (N_2864,N_1805,N_1118);
nor U2865 (N_2865,N_1404,N_1020);
and U2866 (N_2866,N_1863,N_1077);
nor U2867 (N_2867,N_1840,N_1367);
nand U2868 (N_2868,N_1606,N_1964);
or U2869 (N_2869,N_1238,N_1892);
and U2870 (N_2870,N_1565,N_1370);
xnor U2871 (N_2871,N_1652,N_1446);
nor U2872 (N_2872,N_1332,N_1439);
nor U2873 (N_2873,N_1727,N_1154);
or U2874 (N_2874,N_1846,N_1450);
and U2875 (N_2875,N_1624,N_1082);
and U2876 (N_2876,N_1157,N_1939);
and U2877 (N_2877,N_1994,N_1479);
nand U2878 (N_2878,N_1150,N_1285);
and U2879 (N_2879,N_1649,N_1067);
or U2880 (N_2880,N_1613,N_1925);
nand U2881 (N_2881,N_1276,N_1696);
or U2882 (N_2882,N_1858,N_1248);
or U2883 (N_2883,N_1747,N_1974);
or U2884 (N_2884,N_1887,N_1826);
nor U2885 (N_2885,N_1300,N_1953);
or U2886 (N_2886,N_1040,N_1996);
and U2887 (N_2887,N_1768,N_1212);
and U2888 (N_2888,N_1794,N_1404);
and U2889 (N_2889,N_1805,N_1318);
and U2890 (N_2890,N_1801,N_1069);
nand U2891 (N_2891,N_1028,N_1664);
nor U2892 (N_2892,N_1741,N_1237);
nand U2893 (N_2893,N_1910,N_1046);
and U2894 (N_2894,N_1971,N_1298);
and U2895 (N_2895,N_1939,N_1714);
nand U2896 (N_2896,N_1185,N_1028);
or U2897 (N_2897,N_1878,N_1648);
or U2898 (N_2898,N_1843,N_1340);
nor U2899 (N_2899,N_1501,N_1142);
nand U2900 (N_2900,N_1615,N_1788);
nor U2901 (N_2901,N_1270,N_1124);
and U2902 (N_2902,N_1285,N_1858);
nand U2903 (N_2903,N_1475,N_1968);
nor U2904 (N_2904,N_1260,N_1812);
nor U2905 (N_2905,N_1555,N_1618);
nor U2906 (N_2906,N_1339,N_1003);
or U2907 (N_2907,N_1300,N_1965);
and U2908 (N_2908,N_1084,N_1210);
nand U2909 (N_2909,N_1690,N_1635);
xor U2910 (N_2910,N_1782,N_1646);
nor U2911 (N_2911,N_1172,N_1839);
and U2912 (N_2912,N_1980,N_1393);
and U2913 (N_2913,N_1812,N_1001);
nor U2914 (N_2914,N_1959,N_1648);
xnor U2915 (N_2915,N_1189,N_1863);
or U2916 (N_2916,N_1424,N_1669);
and U2917 (N_2917,N_1452,N_1510);
and U2918 (N_2918,N_1961,N_1554);
nor U2919 (N_2919,N_1290,N_1605);
nor U2920 (N_2920,N_1164,N_1661);
xnor U2921 (N_2921,N_1547,N_1866);
nand U2922 (N_2922,N_1196,N_1043);
nand U2923 (N_2923,N_1370,N_1049);
nor U2924 (N_2924,N_1016,N_1002);
nand U2925 (N_2925,N_1334,N_1792);
nand U2926 (N_2926,N_1227,N_1018);
nand U2927 (N_2927,N_1495,N_1650);
or U2928 (N_2928,N_1473,N_1353);
and U2929 (N_2929,N_1213,N_1821);
nand U2930 (N_2930,N_1576,N_1028);
and U2931 (N_2931,N_1421,N_1805);
and U2932 (N_2932,N_1529,N_1336);
nor U2933 (N_2933,N_1210,N_1747);
nor U2934 (N_2934,N_1321,N_1184);
nand U2935 (N_2935,N_1151,N_1734);
xor U2936 (N_2936,N_1303,N_1800);
xnor U2937 (N_2937,N_1317,N_1583);
nand U2938 (N_2938,N_1001,N_1080);
and U2939 (N_2939,N_1728,N_1014);
nor U2940 (N_2940,N_1459,N_1322);
nor U2941 (N_2941,N_1756,N_1680);
and U2942 (N_2942,N_1228,N_1248);
and U2943 (N_2943,N_1217,N_1896);
or U2944 (N_2944,N_1493,N_1577);
xnor U2945 (N_2945,N_1670,N_1705);
nand U2946 (N_2946,N_1518,N_1197);
or U2947 (N_2947,N_1555,N_1675);
or U2948 (N_2948,N_1332,N_1474);
and U2949 (N_2949,N_1283,N_1479);
nand U2950 (N_2950,N_1860,N_1096);
nor U2951 (N_2951,N_1959,N_1437);
nor U2952 (N_2952,N_1340,N_1123);
or U2953 (N_2953,N_1682,N_1096);
nor U2954 (N_2954,N_1033,N_1871);
or U2955 (N_2955,N_1107,N_1926);
or U2956 (N_2956,N_1370,N_1006);
and U2957 (N_2957,N_1234,N_1288);
nor U2958 (N_2958,N_1063,N_1316);
and U2959 (N_2959,N_1361,N_1767);
nor U2960 (N_2960,N_1194,N_1533);
and U2961 (N_2961,N_1183,N_1738);
nor U2962 (N_2962,N_1042,N_1861);
nor U2963 (N_2963,N_1422,N_1030);
nand U2964 (N_2964,N_1617,N_1323);
and U2965 (N_2965,N_1333,N_1460);
nor U2966 (N_2966,N_1132,N_1620);
xnor U2967 (N_2967,N_1991,N_1581);
nand U2968 (N_2968,N_1193,N_1285);
nor U2969 (N_2969,N_1420,N_1683);
or U2970 (N_2970,N_1678,N_1012);
or U2971 (N_2971,N_1747,N_1833);
nor U2972 (N_2972,N_1478,N_1198);
nand U2973 (N_2973,N_1876,N_1065);
nand U2974 (N_2974,N_1381,N_1804);
and U2975 (N_2975,N_1173,N_1324);
xor U2976 (N_2976,N_1765,N_1170);
or U2977 (N_2977,N_1294,N_1572);
nand U2978 (N_2978,N_1121,N_1682);
and U2979 (N_2979,N_1349,N_1392);
and U2980 (N_2980,N_1807,N_1720);
nand U2981 (N_2981,N_1555,N_1214);
nand U2982 (N_2982,N_1710,N_1244);
and U2983 (N_2983,N_1040,N_1354);
or U2984 (N_2984,N_1536,N_1284);
nor U2985 (N_2985,N_1549,N_1802);
and U2986 (N_2986,N_1661,N_1043);
nand U2987 (N_2987,N_1869,N_1084);
nand U2988 (N_2988,N_1694,N_1673);
nand U2989 (N_2989,N_1543,N_1153);
and U2990 (N_2990,N_1297,N_1940);
nor U2991 (N_2991,N_1597,N_1361);
or U2992 (N_2992,N_1219,N_1160);
xor U2993 (N_2993,N_1925,N_1000);
nor U2994 (N_2994,N_1909,N_1388);
nand U2995 (N_2995,N_1378,N_1715);
nor U2996 (N_2996,N_1780,N_1003);
nor U2997 (N_2997,N_1172,N_1559);
nand U2998 (N_2998,N_1211,N_1585);
and U2999 (N_2999,N_1001,N_1704);
nor U3000 (N_3000,N_2391,N_2363);
or U3001 (N_3001,N_2206,N_2491);
and U3002 (N_3002,N_2428,N_2625);
nand U3003 (N_3003,N_2186,N_2298);
and U3004 (N_3004,N_2168,N_2485);
xnor U3005 (N_3005,N_2291,N_2189);
nor U3006 (N_3006,N_2470,N_2015);
xor U3007 (N_3007,N_2576,N_2759);
or U3008 (N_3008,N_2224,N_2596);
and U3009 (N_3009,N_2593,N_2272);
and U3010 (N_3010,N_2247,N_2176);
nor U3011 (N_3011,N_2644,N_2503);
or U3012 (N_3012,N_2094,N_2058);
or U3013 (N_3013,N_2557,N_2723);
xor U3014 (N_3014,N_2336,N_2925);
nor U3015 (N_3015,N_2151,N_2267);
or U3016 (N_3016,N_2314,N_2187);
nor U3017 (N_3017,N_2829,N_2167);
nor U3018 (N_3018,N_2992,N_2139);
or U3019 (N_3019,N_2653,N_2210);
or U3020 (N_3020,N_2817,N_2463);
or U3021 (N_3021,N_2700,N_2376);
nand U3022 (N_3022,N_2136,N_2698);
and U3023 (N_3023,N_2871,N_2414);
and U3024 (N_3024,N_2431,N_2506);
and U3025 (N_3025,N_2243,N_2248);
nand U3026 (N_3026,N_2795,N_2575);
nand U3027 (N_3027,N_2872,N_2241);
or U3028 (N_3028,N_2535,N_2319);
nand U3029 (N_3029,N_2328,N_2157);
nor U3030 (N_3030,N_2201,N_2231);
or U3031 (N_3031,N_2878,N_2061);
nand U3032 (N_3032,N_2626,N_2322);
and U3033 (N_3033,N_2707,N_2837);
or U3034 (N_3034,N_2358,N_2311);
and U3035 (N_3035,N_2184,N_2156);
xor U3036 (N_3036,N_2216,N_2798);
and U3037 (N_3037,N_2558,N_2048);
nand U3038 (N_3038,N_2832,N_2235);
nor U3039 (N_3039,N_2859,N_2426);
nor U3040 (N_3040,N_2631,N_2198);
xor U3041 (N_3041,N_2359,N_2733);
nor U3042 (N_3042,N_2964,N_2988);
and U3043 (N_3043,N_2325,N_2312);
nor U3044 (N_3044,N_2573,N_2996);
and U3045 (N_3045,N_2595,N_2303);
nand U3046 (N_3046,N_2246,N_2571);
nand U3047 (N_3047,N_2137,N_2731);
or U3048 (N_3048,N_2882,N_2743);
xor U3049 (N_3049,N_2822,N_2332);
nand U3050 (N_3050,N_2831,N_2761);
nor U3051 (N_3051,N_2114,N_2676);
and U3052 (N_3052,N_2757,N_2977);
xor U3053 (N_3053,N_2038,N_2310);
nand U3054 (N_3054,N_2523,N_2824);
nand U3055 (N_3055,N_2263,N_2495);
nor U3056 (N_3056,N_2889,N_2851);
xor U3057 (N_3057,N_2835,N_2497);
nand U3058 (N_3058,N_2254,N_2300);
xor U3059 (N_3059,N_2685,N_2570);
nand U3060 (N_3060,N_2672,N_2739);
and U3061 (N_3061,N_2338,N_2869);
nand U3062 (N_3062,N_2389,N_2984);
and U3063 (N_3063,N_2409,N_2531);
and U3064 (N_3064,N_2043,N_2746);
and U3065 (N_3065,N_2906,N_2930);
or U3066 (N_3066,N_2429,N_2682);
nor U3067 (N_3067,N_2599,N_2861);
or U3068 (N_3068,N_2553,N_2732);
nor U3069 (N_3069,N_2991,N_2021);
or U3070 (N_3070,N_2126,N_2270);
nand U3071 (N_3071,N_2771,N_2987);
nor U3072 (N_3072,N_2393,N_2070);
nand U3073 (N_3073,N_2960,N_2366);
xnor U3074 (N_3074,N_2983,N_2800);
or U3075 (N_3075,N_2605,N_2350);
xnor U3076 (N_3076,N_2640,N_2727);
nand U3077 (N_3077,N_2057,N_2102);
or U3078 (N_3078,N_2666,N_2636);
nand U3079 (N_3079,N_2630,N_2180);
xnor U3080 (N_3080,N_2945,N_2153);
nor U3081 (N_3081,N_2858,N_2588);
nand U3082 (N_3082,N_2067,N_2489);
nand U3083 (N_3083,N_2624,N_2063);
xnor U3084 (N_3084,N_2117,N_2279);
and U3085 (N_3085,N_2195,N_2197);
and U3086 (N_3086,N_2000,N_2737);
nor U3087 (N_3087,N_2888,N_2074);
and U3088 (N_3088,N_2348,N_2234);
or U3089 (N_3089,N_2440,N_2213);
or U3090 (N_3090,N_2099,N_2055);
nand U3091 (N_3091,N_2637,N_2657);
xnor U3092 (N_3092,N_2401,N_2677);
and U3093 (N_3093,N_2592,N_2266);
nand U3094 (N_3094,N_2435,N_2381);
xor U3095 (N_3095,N_2935,N_2719);
nor U3096 (N_3096,N_2710,N_2540);
or U3097 (N_3097,N_2365,N_2967);
nor U3098 (N_3098,N_2649,N_2068);
or U3099 (N_3099,N_2623,N_2915);
and U3100 (N_3100,N_2205,N_2769);
nor U3101 (N_3101,N_2229,N_2430);
or U3102 (N_3102,N_2635,N_2484);
nor U3103 (N_3103,N_2768,N_2883);
xor U3104 (N_3104,N_2937,N_2375);
or U3105 (N_3105,N_2536,N_2346);
xor U3106 (N_3106,N_2678,N_2276);
and U3107 (N_3107,N_2360,N_2679);
nand U3108 (N_3108,N_2674,N_2514);
and U3109 (N_3109,N_2821,N_2308);
or U3110 (N_3110,N_2708,N_2980);
nand U3111 (N_3111,N_2131,N_2766);
and U3112 (N_3112,N_2335,N_2193);
and U3113 (N_3113,N_2403,N_2486);
nor U3114 (N_3114,N_2979,N_2842);
nand U3115 (N_3115,N_2284,N_2345);
nand U3116 (N_3116,N_2518,N_2022);
nand U3117 (N_3117,N_2212,N_2788);
or U3118 (N_3118,N_2159,N_2245);
nand U3119 (N_3119,N_2368,N_2309);
and U3120 (N_3120,N_2443,N_2493);
and U3121 (N_3121,N_2863,N_2090);
nand U3122 (N_3122,N_2482,N_2876);
or U3123 (N_3123,N_2681,N_2268);
nor U3124 (N_3124,N_2574,N_2934);
nand U3125 (N_3125,N_2447,N_2966);
nand U3126 (N_3126,N_2107,N_2778);
and U3127 (N_3127,N_2961,N_2646);
nor U3128 (N_3128,N_2549,N_2011);
nand U3129 (N_3129,N_2053,N_2958);
nand U3130 (N_3130,N_2460,N_2718);
xor U3131 (N_3131,N_2907,N_2146);
nand U3132 (N_3132,N_2620,N_2668);
or U3133 (N_3133,N_2388,N_2475);
or U3134 (N_3134,N_2647,N_2232);
nor U3135 (N_3135,N_2455,N_2548);
or U3136 (N_3136,N_2087,N_2295);
or U3137 (N_3137,N_2404,N_2294);
and U3138 (N_3138,N_2199,N_2974);
nand U3139 (N_3139,N_2610,N_2572);
xnor U3140 (N_3140,N_2149,N_2799);
xnor U3141 (N_3141,N_2249,N_2611);
nor U3142 (N_3142,N_2041,N_2116);
or U3143 (N_3143,N_2299,N_2892);
nor U3144 (N_3144,N_2713,N_2385);
and U3145 (N_3145,N_2801,N_2989);
nor U3146 (N_3146,N_2545,N_2551);
or U3147 (N_3147,N_2807,N_2814);
or U3148 (N_3148,N_2776,N_2519);
xor U3149 (N_3149,N_2877,N_2018);
and U3150 (N_3150,N_2233,N_2562);
xnor U3151 (N_3151,N_2113,N_2833);
nand U3152 (N_3152,N_2612,N_2128);
nor U3153 (N_3153,N_2533,N_2292);
nand U3154 (N_3154,N_2971,N_2926);
or U3155 (N_3155,N_2826,N_2754);
nor U3156 (N_3156,N_2777,N_2617);
and U3157 (N_3157,N_2418,N_2780);
nor U3158 (N_3158,N_2097,N_2045);
nor U3159 (N_3159,N_2394,N_2855);
or U3160 (N_3160,N_2382,N_2112);
nand U3161 (N_3161,N_2024,N_2577);
and U3162 (N_3162,N_2032,N_2690);
nor U3163 (N_3163,N_2694,N_2804);
xor U3164 (N_3164,N_2741,N_2616);
or U3165 (N_3165,N_2029,N_2101);
and U3166 (N_3166,N_2969,N_2086);
nor U3167 (N_3167,N_2717,N_2661);
nor U3168 (N_3168,N_2929,N_2257);
nand U3169 (N_3169,N_2341,N_2020);
nor U3170 (N_3170,N_2283,N_2315);
and U3171 (N_3171,N_2454,N_2367);
or U3172 (N_3172,N_2106,N_2880);
nor U3173 (N_3173,N_2902,N_2342);
and U3174 (N_3174,N_2852,N_2242);
or U3175 (N_3175,N_2501,N_2639);
and U3176 (N_3176,N_2995,N_2490);
nand U3177 (N_3177,N_2405,N_2185);
or U3178 (N_3178,N_2856,N_2480);
nand U3179 (N_3179,N_2083,N_2488);
nor U3180 (N_3180,N_2261,N_2815);
nand U3181 (N_3181,N_2377,N_2753);
or U3182 (N_3182,N_2012,N_2986);
or U3183 (N_3183,N_2450,N_2467);
nor U3184 (N_3184,N_2181,N_2673);
and U3185 (N_3185,N_2786,N_2100);
and U3186 (N_3186,N_2035,N_2357);
or U3187 (N_3187,N_2515,N_2569);
nor U3188 (N_3188,N_2508,N_2420);
xnor U3189 (N_3189,N_2158,N_2349);
or U3190 (N_3190,N_2343,N_2013);
and U3191 (N_3191,N_2092,N_2323);
or U3192 (N_3192,N_2155,N_2908);
and U3193 (N_3193,N_2699,N_2803);
xnor U3194 (N_3194,N_2913,N_2845);
xor U3195 (N_3195,N_2361,N_2237);
or U3196 (N_3196,N_2862,N_2665);
xnor U3197 (N_3197,N_2655,N_2396);
or U3198 (N_3198,N_2098,N_2287);
nor U3199 (N_3199,N_2093,N_2065);
nor U3200 (N_3200,N_2433,N_2903);
nor U3201 (N_3201,N_2684,N_2938);
nand U3202 (N_3202,N_2749,N_2884);
nor U3203 (N_3203,N_2683,N_2785);
nor U3204 (N_3204,N_2395,N_2687);
and U3205 (N_3205,N_2179,N_2281);
nor U3206 (N_3206,N_2347,N_2942);
nand U3207 (N_3207,N_2203,N_2597);
nor U3208 (N_3208,N_2161,N_2001);
and U3209 (N_3209,N_2546,N_2652);
and U3210 (N_3210,N_2949,N_2006);
and U3211 (N_3211,N_2783,N_2520);
nor U3212 (N_3212,N_2525,N_2073);
xor U3213 (N_3213,N_2010,N_2337);
or U3214 (N_3214,N_2260,N_2316);
nor U3215 (N_3215,N_2830,N_2905);
and U3216 (N_3216,N_2633,N_2096);
or U3217 (N_3217,N_2554,N_2277);
nor U3218 (N_3218,N_2479,N_2946);
and U3219 (N_3219,N_2805,N_2601);
nor U3220 (N_3220,N_2478,N_2943);
nand U3221 (N_3221,N_2129,N_2118);
and U3222 (N_3222,N_2947,N_2921);
and U3223 (N_3223,N_2274,N_2530);
nor U3224 (N_3224,N_2910,N_2072);
and U3225 (N_3225,N_2912,N_2051);
nor U3226 (N_3226,N_2148,N_2779);
or U3227 (N_3227,N_2544,N_2629);
or U3228 (N_3228,N_2005,N_2280);
or U3229 (N_3229,N_2836,N_2244);
nor U3230 (N_3230,N_2371,N_2190);
nor U3231 (N_3231,N_2772,N_2529);
or U3232 (N_3232,N_2999,N_2773);
and U3233 (N_3233,N_2033,N_2162);
nand U3234 (N_3234,N_2502,N_2787);
nor U3235 (N_3235,N_2143,N_2142);
nor U3236 (N_3236,N_2296,N_2400);
and U3237 (N_3237,N_2568,N_2030);
and U3238 (N_3238,N_2004,N_2613);
or U3239 (N_3239,N_2680,N_2221);
nor U3240 (N_3240,N_2049,N_2066);
nand U3241 (N_3241,N_2432,N_2191);
and U3242 (N_3242,N_2932,N_2793);
or U3243 (N_3243,N_2471,N_2725);
nand U3244 (N_3244,N_2751,N_2209);
nor U3245 (N_3245,N_2663,N_2056);
and U3246 (N_3246,N_2563,N_2002);
nand U3247 (N_3247,N_2386,N_2062);
nand U3248 (N_3248,N_2567,N_2164);
nor U3249 (N_3249,N_2782,N_2172);
and U3250 (N_3250,N_2696,N_2111);
or U3251 (N_3251,N_2427,N_2327);
xor U3252 (N_3252,N_2584,N_2944);
or U3253 (N_3253,N_2448,N_2973);
and U3254 (N_3254,N_2868,N_2927);
and U3255 (N_3255,N_2899,N_2196);
xnor U3256 (N_3256,N_2583,N_2522);
or U3257 (N_3257,N_2622,N_2147);
or U3258 (N_3258,N_2036,N_2524);
or U3259 (N_3259,N_2269,N_2078);
and U3260 (N_3260,N_2765,N_2370);
or U3261 (N_3261,N_2970,N_2014);
nor U3262 (N_3262,N_2105,N_2306);
and U3263 (N_3263,N_2919,N_2660);
nand U3264 (N_3264,N_2378,N_2874);
and U3265 (N_3265,N_2847,N_2556);
xor U3266 (N_3266,N_2591,N_2521);
nand U3267 (N_3267,N_2806,N_2256);
or U3268 (N_3268,N_2288,N_2103);
nor U3269 (N_3269,N_2069,N_2825);
nor U3270 (N_3270,N_2931,N_2507);
nor U3271 (N_3271,N_2658,N_2354);
xor U3272 (N_3272,N_2252,N_2981);
or U3273 (N_3273,N_2517,N_2152);
nor U3274 (N_3274,N_2009,N_2526);
nand U3275 (N_3275,N_2586,N_2924);
nand U3276 (N_3276,N_2618,N_2704);
and U3277 (N_3277,N_2474,N_2374);
or U3278 (N_3278,N_2656,N_2819);
or U3279 (N_3279,N_2461,N_2972);
nand U3280 (N_3280,N_2755,N_2671);
nand U3281 (N_3281,N_2659,N_2648);
nor U3282 (N_3282,N_2415,N_2796);
nor U3283 (N_3283,N_2603,N_2726);
nor U3284 (N_3284,N_2594,N_2140);
and U3285 (N_3285,N_2134,N_2081);
or U3286 (N_3286,N_2750,N_2615);
or U3287 (N_3287,N_2411,N_2505);
nor U3288 (N_3288,N_2820,N_2273);
or U3289 (N_3289,N_2227,N_2222);
and U3290 (N_3290,N_2692,N_2587);
and U3291 (N_3291,N_2650,N_2364);
or U3292 (N_3292,N_2604,N_2387);
nor U3293 (N_3293,N_2498,N_2566);
and U3294 (N_3294,N_2425,N_2133);
and U3295 (N_3295,N_2742,N_2438);
or U3296 (N_3296,N_2775,N_2177);
xnor U3297 (N_3297,N_2959,N_2614);
and U3298 (N_3298,N_2532,N_2564);
nor U3299 (N_3299,N_2027,N_2050);
nand U3300 (N_3300,N_2442,N_2397);
nor U3301 (N_3301,N_2468,N_2154);
nand U3302 (N_3302,N_2552,N_2642);
or U3303 (N_3303,N_2307,N_2898);
and U3304 (N_3304,N_2885,N_2866);
xnor U3305 (N_3305,N_2543,N_2781);
nor U3306 (N_3306,N_2802,N_2132);
or U3307 (N_3307,N_2080,N_2380);
nand U3308 (N_3308,N_2169,N_2954);
or U3309 (N_3309,N_2259,N_2458);
nand U3310 (N_3310,N_2900,N_2703);
nand U3311 (N_3311,N_2634,N_2638);
nor U3312 (N_3312,N_2952,N_2748);
and U3313 (N_3313,N_2774,N_2130);
or U3314 (N_3314,N_2951,N_2127);
nand U3315 (N_3315,N_2997,N_2669);
or U3316 (N_3316,N_2228,N_2079);
or U3317 (N_3317,N_2178,N_2188);
nor U3318 (N_3318,N_2728,N_2909);
and U3319 (N_3319,N_2712,N_2891);
nor U3320 (N_3320,N_2740,N_2729);
nor U3321 (N_3321,N_2922,N_2976);
nand U3322 (N_3322,N_2262,N_2645);
and U3323 (N_3323,N_2369,N_2542);
nand U3324 (N_3324,N_2251,N_2108);
and U3325 (N_3325,N_2144,N_2419);
nand U3326 (N_3326,N_2406,N_2064);
or U3327 (N_3327,N_2091,N_2894);
or U3328 (N_3328,N_2123,N_2706);
nand U3329 (N_3329,N_2606,N_2846);
nor U3330 (N_3330,N_2372,N_2844);
xor U3331 (N_3331,N_2724,N_2607);
xnor U3332 (N_3332,N_2077,N_2339);
nand U3333 (N_3333,N_2459,N_2499);
nand U3334 (N_3334,N_2095,N_2941);
nor U3335 (N_3335,N_2928,N_2745);
nand U3336 (N_3336,N_2392,N_2760);
xnor U3337 (N_3337,N_2953,N_2165);
nand U3338 (N_3338,N_2285,N_2449);
or U3339 (N_3339,N_2441,N_2265);
and U3340 (N_3340,N_2813,N_2963);
or U3341 (N_3341,N_2580,N_2709);
nor U3342 (N_3342,N_2084,N_2076);
nor U3343 (N_3343,N_2879,N_2163);
or U3344 (N_3344,N_2864,N_2686);
nand U3345 (N_3345,N_2122,N_2695);
xor U3346 (N_3346,N_2320,N_2223);
xor U3347 (N_3347,N_2715,N_2512);
and U3348 (N_3348,N_2344,N_2582);
or U3349 (N_3349,N_2956,N_2939);
xnor U3350 (N_3350,N_2561,N_2812);
and U3351 (N_3351,N_2150,N_2452);
xnor U3352 (N_3352,N_2289,N_2810);
nor U3353 (N_3353,N_2439,N_2538);
or U3354 (N_3354,N_2481,N_2840);
or U3355 (N_3355,N_2602,N_2492);
nand U3356 (N_3356,N_2326,N_2059);
nor U3357 (N_3357,N_2220,N_2664);
nand U3358 (N_3358,N_2691,N_2352);
and U3359 (N_3359,N_2434,N_2758);
nor U3360 (N_3360,N_2313,N_2258);
or U3361 (N_3361,N_2962,N_2464);
nand U3362 (N_3362,N_2194,N_2513);
nand U3363 (N_3363,N_2849,N_2735);
nor U3364 (N_3364,N_2711,N_2019);
or U3365 (N_3365,N_2071,N_2355);
nor U3366 (N_3366,N_2641,N_2867);
nor U3367 (N_3367,N_2811,N_2598);
nor U3368 (N_3368,N_2818,N_2860);
nand U3369 (N_3369,N_2330,N_2843);
and U3370 (N_3370,N_2950,N_2689);
nor U3371 (N_3371,N_2911,N_2017);
nand U3372 (N_3372,N_2457,N_2762);
or U3373 (N_3373,N_2250,N_2456);
and U3374 (N_3374,N_2379,N_2763);
and U3375 (N_3375,N_2609,N_2301);
nand U3376 (N_3376,N_2890,N_2318);
xnor U3377 (N_3377,N_2477,N_2887);
or U3378 (N_3378,N_2423,N_2218);
nand U3379 (N_3379,N_2957,N_2870);
nor U3380 (N_3380,N_2792,N_2351);
and U3381 (N_3381,N_2720,N_2895);
nand U3382 (N_3382,N_2383,N_2914);
nand U3383 (N_3383,N_2255,N_2560);
or U3384 (N_3384,N_2333,N_2736);
and U3385 (N_3385,N_2042,N_2075);
nand U3386 (N_3386,N_2444,N_2886);
nand U3387 (N_3387,N_2628,N_2756);
or U3388 (N_3388,N_2085,N_2175);
xor U3389 (N_3389,N_2412,N_2119);
and U3390 (N_3390,N_2290,N_2643);
nand U3391 (N_3391,N_2565,N_2994);
nor U3392 (N_3392,N_2025,N_2271);
and U3393 (N_3393,N_2770,N_2487);
nor U3394 (N_3394,N_2413,N_2496);
nand U3395 (N_3395,N_2236,N_2917);
nor U3396 (N_3396,N_2722,N_2896);
nand U3397 (N_3397,N_2125,N_2110);
and U3398 (N_3398,N_2916,N_2982);
xor U3399 (N_3399,N_2023,N_2559);
nor U3400 (N_3400,N_2701,N_2834);
and U3401 (N_3401,N_2621,N_2225);
nor U3402 (N_3402,N_2402,N_2923);
nand U3403 (N_3403,N_2437,N_2219);
xor U3404 (N_3404,N_2933,N_2200);
and U3405 (N_3405,N_2183,N_2693);
nand U3406 (N_3406,N_2453,N_2940);
nand U3407 (N_3407,N_2321,N_2767);
nand U3408 (N_3408,N_2476,N_2747);
nand U3409 (N_3409,N_2208,N_2124);
nor U3410 (N_3410,N_2993,N_2881);
and U3411 (N_3411,N_2721,N_2590);
xor U3412 (N_3412,N_2848,N_2238);
or U3413 (N_3413,N_2702,N_2893);
xnor U3414 (N_3414,N_2865,N_2334);
nor U3415 (N_3415,N_2034,N_2145);
or U3416 (N_3416,N_2579,N_2424);
or U3417 (N_3417,N_2230,N_2253);
nand U3418 (N_3418,N_2965,N_2465);
and U3419 (N_3419,N_2304,N_2317);
nand U3420 (N_3420,N_2264,N_2037);
nor U3421 (N_3421,N_2654,N_2857);
nor U3422 (N_3422,N_2918,N_2578);
nand U3423 (N_3423,N_2509,N_2904);
or U3424 (N_3424,N_2282,N_2662);
or U3425 (N_3425,N_2044,N_2500);
or U3426 (N_3426,N_2534,N_2998);
and U3427 (N_3427,N_2469,N_2978);
and U3428 (N_3428,N_2115,N_2293);
or U3429 (N_3429,N_2539,N_2823);
or U3430 (N_3430,N_2297,N_2302);
nor U3431 (N_3431,N_2504,N_2088);
and U3432 (N_3432,N_2714,N_2160);
xor U3433 (N_3433,N_2581,N_2331);
nor U3434 (N_3434,N_2046,N_2555);
or U3435 (N_3435,N_2275,N_2510);
nand U3436 (N_3436,N_2026,N_2240);
nor U3437 (N_3437,N_2784,N_2794);
nor U3438 (N_3438,N_2516,N_2827);
and U3439 (N_3439,N_2436,N_2166);
nand U3440 (N_3440,N_2373,N_2541);
nand U3441 (N_3441,N_2028,N_2353);
or U3442 (N_3442,N_2632,N_2651);
or U3443 (N_3443,N_2362,N_2039);
or U3444 (N_3444,N_2670,N_2171);
or U3445 (N_3445,N_2054,N_2990);
xor U3446 (N_3446,N_2838,N_2104);
and U3447 (N_3447,N_2791,N_2138);
nand U3448 (N_3448,N_2955,N_2547);
nor U3449 (N_3449,N_2003,N_2985);
nand U3450 (N_3450,N_2445,N_2528);
nand U3451 (N_3451,N_2734,N_2619);
nor U3452 (N_3452,N_2390,N_2853);
or U3453 (N_3453,N_2040,N_2550);
nand U3454 (N_3454,N_2790,N_2816);
nand U3455 (N_3455,N_2667,N_2120);
nand U3456 (N_3456,N_2089,N_2466);
nand U3457 (N_3457,N_2808,N_2410);
xor U3458 (N_3458,N_2627,N_2809);
xnor U3459 (N_3459,N_2936,N_2173);
or U3460 (N_3460,N_2416,N_2850);
and U3461 (N_3461,N_2192,N_2141);
nand U3462 (N_3462,N_2901,N_2217);
or U3463 (N_3463,N_2839,N_2211);
nand U3464 (N_3464,N_2329,N_2697);
nor U3465 (N_3465,N_2340,N_2202);
or U3466 (N_3466,N_2875,N_2174);
nand U3467 (N_3467,N_2407,N_2214);
and U3468 (N_3468,N_2109,N_2239);
or U3469 (N_3469,N_2527,N_2082);
nand U3470 (N_3470,N_2008,N_2408);
and U3471 (N_3471,N_2446,N_2483);
and U3472 (N_3472,N_2585,N_2462);
nor U3473 (N_3473,N_2215,N_2738);
nor U3474 (N_3474,N_2688,N_2511);
nor U3475 (N_3475,N_2473,N_2016);
nor U3476 (N_3476,N_2417,N_2975);
xnor U3477 (N_3477,N_2060,N_2286);
nor U3478 (N_3478,N_2472,N_2031);
or U3479 (N_3479,N_2841,N_2278);
or U3480 (N_3480,N_2052,N_2047);
or U3481 (N_3481,N_2121,N_2873);
nand U3482 (N_3482,N_2182,N_2384);
nand U3483 (N_3483,N_2744,N_2204);
nor U3484 (N_3484,N_2968,N_2828);
nor U3485 (N_3485,N_2797,N_2600);
and U3486 (N_3486,N_2356,N_2854);
or U3487 (N_3487,N_2170,N_2494);
nand U3488 (N_3488,N_2920,N_2730);
and U3489 (N_3489,N_2422,N_2675);
nor U3490 (N_3490,N_2716,N_2537);
nor U3491 (N_3491,N_2948,N_2207);
or U3492 (N_3492,N_2789,N_2421);
or U3493 (N_3493,N_2135,N_2324);
nor U3494 (N_3494,N_2305,N_2705);
or U3495 (N_3495,N_2608,N_2007);
and U3496 (N_3496,N_2399,N_2226);
nand U3497 (N_3497,N_2451,N_2589);
and U3498 (N_3498,N_2398,N_2764);
or U3499 (N_3499,N_2897,N_2752);
nor U3500 (N_3500,N_2032,N_2975);
or U3501 (N_3501,N_2738,N_2276);
and U3502 (N_3502,N_2234,N_2447);
nor U3503 (N_3503,N_2898,N_2812);
nand U3504 (N_3504,N_2044,N_2821);
nand U3505 (N_3505,N_2714,N_2475);
or U3506 (N_3506,N_2523,N_2794);
nor U3507 (N_3507,N_2371,N_2996);
nand U3508 (N_3508,N_2560,N_2850);
nand U3509 (N_3509,N_2030,N_2514);
nand U3510 (N_3510,N_2162,N_2294);
nand U3511 (N_3511,N_2001,N_2936);
and U3512 (N_3512,N_2181,N_2421);
nor U3513 (N_3513,N_2252,N_2576);
or U3514 (N_3514,N_2256,N_2378);
and U3515 (N_3515,N_2153,N_2904);
xnor U3516 (N_3516,N_2626,N_2378);
and U3517 (N_3517,N_2526,N_2212);
and U3518 (N_3518,N_2339,N_2128);
and U3519 (N_3519,N_2337,N_2928);
nand U3520 (N_3520,N_2218,N_2143);
nor U3521 (N_3521,N_2157,N_2098);
nand U3522 (N_3522,N_2864,N_2497);
or U3523 (N_3523,N_2169,N_2147);
and U3524 (N_3524,N_2106,N_2734);
and U3525 (N_3525,N_2955,N_2909);
or U3526 (N_3526,N_2848,N_2370);
or U3527 (N_3527,N_2383,N_2946);
or U3528 (N_3528,N_2957,N_2074);
and U3529 (N_3529,N_2229,N_2071);
nor U3530 (N_3530,N_2391,N_2915);
nor U3531 (N_3531,N_2861,N_2156);
nor U3532 (N_3532,N_2742,N_2227);
nand U3533 (N_3533,N_2935,N_2197);
and U3534 (N_3534,N_2523,N_2083);
and U3535 (N_3535,N_2449,N_2122);
xnor U3536 (N_3536,N_2215,N_2584);
and U3537 (N_3537,N_2047,N_2139);
or U3538 (N_3538,N_2488,N_2632);
and U3539 (N_3539,N_2320,N_2654);
nor U3540 (N_3540,N_2007,N_2651);
or U3541 (N_3541,N_2043,N_2291);
nand U3542 (N_3542,N_2193,N_2962);
and U3543 (N_3543,N_2935,N_2676);
and U3544 (N_3544,N_2325,N_2254);
and U3545 (N_3545,N_2054,N_2048);
xnor U3546 (N_3546,N_2665,N_2848);
nand U3547 (N_3547,N_2224,N_2049);
nand U3548 (N_3548,N_2391,N_2532);
nand U3549 (N_3549,N_2160,N_2838);
nand U3550 (N_3550,N_2747,N_2626);
nand U3551 (N_3551,N_2974,N_2264);
or U3552 (N_3552,N_2700,N_2844);
or U3553 (N_3553,N_2768,N_2159);
nand U3554 (N_3554,N_2933,N_2727);
or U3555 (N_3555,N_2053,N_2386);
nand U3556 (N_3556,N_2762,N_2889);
nand U3557 (N_3557,N_2205,N_2856);
and U3558 (N_3558,N_2779,N_2160);
or U3559 (N_3559,N_2948,N_2549);
xnor U3560 (N_3560,N_2861,N_2335);
nor U3561 (N_3561,N_2820,N_2139);
or U3562 (N_3562,N_2825,N_2438);
and U3563 (N_3563,N_2804,N_2070);
and U3564 (N_3564,N_2031,N_2408);
or U3565 (N_3565,N_2216,N_2641);
and U3566 (N_3566,N_2609,N_2305);
and U3567 (N_3567,N_2849,N_2844);
or U3568 (N_3568,N_2193,N_2538);
nand U3569 (N_3569,N_2523,N_2194);
nand U3570 (N_3570,N_2265,N_2694);
nand U3571 (N_3571,N_2882,N_2278);
nand U3572 (N_3572,N_2703,N_2124);
nor U3573 (N_3573,N_2880,N_2286);
nor U3574 (N_3574,N_2018,N_2936);
nand U3575 (N_3575,N_2039,N_2213);
xnor U3576 (N_3576,N_2647,N_2768);
and U3577 (N_3577,N_2623,N_2914);
nor U3578 (N_3578,N_2815,N_2823);
or U3579 (N_3579,N_2686,N_2898);
nor U3580 (N_3580,N_2024,N_2838);
and U3581 (N_3581,N_2347,N_2494);
and U3582 (N_3582,N_2635,N_2932);
nor U3583 (N_3583,N_2583,N_2638);
or U3584 (N_3584,N_2411,N_2660);
nand U3585 (N_3585,N_2502,N_2677);
nor U3586 (N_3586,N_2081,N_2524);
nor U3587 (N_3587,N_2680,N_2104);
nand U3588 (N_3588,N_2218,N_2965);
nor U3589 (N_3589,N_2384,N_2238);
nand U3590 (N_3590,N_2432,N_2395);
nand U3591 (N_3591,N_2793,N_2704);
or U3592 (N_3592,N_2415,N_2495);
nand U3593 (N_3593,N_2771,N_2891);
nor U3594 (N_3594,N_2504,N_2289);
or U3595 (N_3595,N_2388,N_2311);
nor U3596 (N_3596,N_2413,N_2523);
nand U3597 (N_3597,N_2142,N_2990);
xnor U3598 (N_3598,N_2422,N_2922);
and U3599 (N_3599,N_2959,N_2375);
or U3600 (N_3600,N_2997,N_2306);
nand U3601 (N_3601,N_2936,N_2865);
or U3602 (N_3602,N_2765,N_2005);
nor U3603 (N_3603,N_2065,N_2490);
nand U3604 (N_3604,N_2774,N_2656);
and U3605 (N_3605,N_2616,N_2977);
or U3606 (N_3606,N_2897,N_2456);
nor U3607 (N_3607,N_2570,N_2455);
nor U3608 (N_3608,N_2812,N_2780);
and U3609 (N_3609,N_2908,N_2892);
and U3610 (N_3610,N_2632,N_2669);
or U3611 (N_3611,N_2785,N_2871);
and U3612 (N_3612,N_2089,N_2204);
nor U3613 (N_3613,N_2247,N_2468);
or U3614 (N_3614,N_2748,N_2130);
and U3615 (N_3615,N_2626,N_2468);
and U3616 (N_3616,N_2706,N_2793);
xor U3617 (N_3617,N_2919,N_2215);
nand U3618 (N_3618,N_2026,N_2024);
and U3619 (N_3619,N_2395,N_2601);
nor U3620 (N_3620,N_2840,N_2663);
nor U3621 (N_3621,N_2455,N_2554);
nand U3622 (N_3622,N_2342,N_2722);
and U3623 (N_3623,N_2320,N_2171);
and U3624 (N_3624,N_2197,N_2779);
xor U3625 (N_3625,N_2091,N_2013);
nor U3626 (N_3626,N_2847,N_2517);
and U3627 (N_3627,N_2269,N_2177);
nor U3628 (N_3628,N_2639,N_2380);
or U3629 (N_3629,N_2217,N_2360);
and U3630 (N_3630,N_2741,N_2470);
or U3631 (N_3631,N_2486,N_2501);
or U3632 (N_3632,N_2430,N_2135);
nand U3633 (N_3633,N_2001,N_2136);
or U3634 (N_3634,N_2538,N_2434);
or U3635 (N_3635,N_2330,N_2902);
and U3636 (N_3636,N_2582,N_2306);
nor U3637 (N_3637,N_2138,N_2730);
and U3638 (N_3638,N_2186,N_2141);
nand U3639 (N_3639,N_2504,N_2607);
and U3640 (N_3640,N_2276,N_2760);
nand U3641 (N_3641,N_2976,N_2307);
or U3642 (N_3642,N_2223,N_2260);
and U3643 (N_3643,N_2401,N_2436);
nor U3644 (N_3644,N_2466,N_2519);
and U3645 (N_3645,N_2711,N_2225);
and U3646 (N_3646,N_2971,N_2424);
nor U3647 (N_3647,N_2741,N_2379);
and U3648 (N_3648,N_2450,N_2649);
nand U3649 (N_3649,N_2083,N_2334);
and U3650 (N_3650,N_2016,N_2812);
and U3651 (N_3651,N_2705,N_2929);
nand U3652 (N_3652,N_2621,N_2100);
and U3653 (N_3653,N_2889,N_2361);
and U3654 (N_3654,N_2995,N_2266);
or U3655 (N_3655,N_2417,N_2111);
nand U3656 (N_3656,N_2809,N_2650);
or U3657 (N_3657,N_2763,N_2548);
nor U3658 (N_3658,N_2234,N_2745);
nand U3659 (N_3659,N_2764,N_2809);
nand U3660 (N_3660,N_2069,N_2940);
and U3661 (N_3661,N_2730,N_2296);
and U3662 (N_3662,N_2946,N_2522);
and U3663 (N_3663,N_2877,N_2200);
or U3664 (N_3664,N_2832,N_2390);
nand U3665 (N_3665,N_2976,N_2303);
nand U3666 (N_3666,N_2242,N_2157);
nand U3667 (N_3667,N_2864,N_2585);
nor U3668 (N_3668,N_2842,N_2893);
nand U3669 (N_3669,N_2170,N_2437);
nand U3670 (N_3670,N_2946,N_2011);
nor U3671 (N_3671,N_2198,N_2159);
or U3672 (N_3672,N_2063,N_2996);
or U3673 (N_3673,N_2012,N_2239);
or U3674 (N_3674,N_2512,N_2613);
or U3675 (N_3675,N_2422,N_2663);
xor U3676 (N_3676,N_2761,N_2281);
xnor U3677 (N_3677,N_2383,N_2856);
nand U3678 (N_3678,N_2717,N_2076);
or U3679 (N_3679,N_2112,N_2438);
xnor U3680 (N_3680,N_2535,N_2665);
and U3681 (N_3681,N_2632,N_2025);
or U3682 (N_3682,N_2305,N_2752);
nor U3683 (N_3683,N_2171,N_2696);
or U3684 (N_3684,N_2814,N_2270);
or U3685 (N_3685,N_2894,N_2716);
or U3686 (N_3686,N_2802,N_2179);
and U3687 (N_3687,N_2619,N_2418);
or U3688 (N_3688,N_2588,N_2338);
nand U3689 (N_3689,N_2718,N_2479);
and U3690 (N_3690,N_2218,N_2402);
and U3691 (N_3691,N_2129,N_2987);
nand U3692 (N_3692,N_2320,N_2466);
and U3693 (N_3693,N_2485,N_2795);
nor U3694 (N_3694,N_2152,N_2418);
nor U3695 (N_3695,N_2707,N_2753);
xor U3696 (N_3696,N_2574,N_2213);
nand U3697 (N_3697,N_2882,N_2289);
and U3698 (N_3698,N_2107,N_2584);
nor U3699 (N_3699,N_2986,N_2163);
nor U3700 (N_3700,N_2647,N_2637);
and U3701 (N_3701,N_2168,N_2280);
nand U3702 (N_3702,N_2037,N_2570);
or U3703 (N_3703,N_2137,N_2207);
nor U3704 (N_3704,N_2871,N_2345);
nand U3705 (N_3705,N_2762,N_2216);
or U3706 (N_3706,N_2338,N_2330);
nand U3707 (N_3707,N_2447,N_2843);
xor U3708 (N_3708,N_2493,N_2107);
nand U3709 (N_3709,N_2571,N_2298);
xor U3710 (N_3710,N_2986,N_2676);
and U3711 (N_3711,N_2499,N_2057);
and U3712 (N_3712,N_2506,N_2227);
nor U3713 (N_3713,N_2710,N_2984);
nand U3714 (N_3714,N_2355,N_2278);
xor U3715 (N_3715,N_2136,N_2447);
nand U3716 (N_3716,N_2929,N_2145);
xnor U3717 (N_3717,N_2834,N_2797);
or U3718 (N_3718,N_2505,N_2521);
xnor U3719 (N_3719,N_2173,N_2201);
or U3720 (N_3720,N_2531,N_2005);
nor U3721 (N_3721,N_2375,N_2609);
nor U3722 (N_3722,N_2370,N_2182);
nor U3723 (N_3723,N_2688,N_2849);
nor U3724 (N_3724,N_2060,N_2403);
nor U3725 (N_3725,N_2652,N_2341);
xor U3726 (N_3726,N_2402,N_2583);
nor U3727 (N_3727,N_2329,N_2869);
nor U3728 (N_3728,N_2114,N_2369);
and U3729 (N_3729,N_2279,N_2740);
nor U3730 (N_3730,N_2553,N_2795);
xnor U3731 (N_3731,N_2511,N_2991);
or U3732 (N_3732,N_2478,N_2549);
nand U3733 (N_3733,N_2198,N_2849);
and U3734 (N_3734,N_2688,N_2669);
nor U3735 (N_3735,N_2771,N_2254);
nand U3736 (N_3736,N_2568,N_2840);
nand U3737 (N_3737,N_2354,N_2753);
or U3738 (N_3738,N_2968,N_2678);
nand U3739 (N_3739,N_2116,N_2409);
nor U3740 (N_3740,N_2209,N_2277);
and U3741 (N_3741,N_2829,N_2008);
nand U3742 (N_3742,N_2789,N_2159);
nor U3743 (N_3743,N_2860,N_2732);
nor U3744 (N_3744,N_2838,N_2416);
nor U3745 (N_3745,N_2041,N_2154);
nor U3746 (N_3746,N_2798,N_2056);
nor U3747 (N_3747,N_2506,N_2578);
and U3748 (N_3748,N_2440,N_2000);
nand U3749 (N_3749,N_2220,N_2116);
nor U3750 (N_3750,N_2368,N_2207);
nor U3751 (N_3751,N_2336,N_2141);
nand U3752 (N_3752,N_2389,N_2696);
nand U3753 (N_3753,N_2127,N_2633);
and U3754 (N_3754,N_2810,N_2370);
or U3755 (N_3755,N_2756,N_2072);
nor U3756 (N_3756,N_2384,N_2482);
or U3757 (N_3757,N_2162,N_2928);
nor U3758 (N_3758,N_2902,N_2854);
or U3759 (N_3759,N_2238,N_2018);
or U3760 (N_3760,N_2785,N_2185);
and U3761 (N_3761,N_2262,N_2177);
and U3762 (N_3762,N_2546,N_2333);
nor U3763 (N_3763,N_2296,N_2153);
or U3764 (N_3764,N_2875,N_2923);
nor U3765 (N_3765,N_2271,N_2850);
nor U3766 (N_3766,N_2267,N_2788);
or U3767 (N_3767,N_2778,N_2060);
and U3768 (N_3768,N_2767,N_2181);
nor U3769 (N_3769,N_2961,N_2074);
or U3770 (N_3770,N_2096,N_2343);
xor U3771 (N_3771,N_2050,N_2154);
nand U3772 (N_3772,N_2850,N_2918);
nand U3773 (N_3773,N_2096,N_2806);
nor U3774 (N_3774,N_2761,N_2775);
nand U3775 (N_3775,N_2217,N_2151);
nand U3776 (N_3776,N_2823,N_2621);
or U3777 (N_3777,N_2767,N_2779);
and U3778 (N_3778,N_2507,N_2024);
nor U3779 (N_3779,N_2065,N_2135);
nand U3780 (N_3780,N_2814,N_2336);
or U3781 (N_3781,N_2222,N_2030);
nor U3782 (N_3782,N_2958,N_2644);
xor U3783 (N_3783,N_2873,N_2062);
or U3784 (N_3784,N_2551,N_2110);
xor U3785 (N_3785,N_2213,N_2593);
nand U3786 (N_3786,N_2449,N_2730);
nor U3787 (N_3787,N_2565,N_2649);
nor U3788 (N_3788,N_2069,N_2245);
xnor U3789 (N_3789,N_2972,N_2943);
nand U3790 (N_3790,N_2084,N_2806);
or U3791 (N_3791,N_2540,N_2588);
nor U3792 (N_3792,N_2380,N_2147);
and U3793 (N_3793,N_2249,N_2601);
or U3794 (N_3794,N_2688,N_2659);
or U3795 (N_3795,N_2620,N_2207);
nor U3796 (N_3796,N_2633,N_2100);
nand U3797 (N_3797,N_2001,N_2145);
and U3798 (N_3798,N_2348,N_2022);
and U3799 (N_3799,N_2375,N_2867);
or U3800 (N_3800,N_2854,N_2880);
or U3801 (N_3801,N_2872,N_2031);
nor U3802 (N_3802,N_2094,N_2827);
or U3803 (N_3803,N_2756,N_2565);
and U3804 (N_3804,N_2838,N_2902);
xor U3805 (N_3805,N_2085,N_2702);
or U3806 (N_3806,N_2272,N_2823);
nand U3807 (N_3807,N_2356,N_2532);
and U3808 (N_3808,N_2676,N_2889);
nor U3809 (N_3809,N_2111,N_2213);
and U3810 (N_3810,N_2087,N_2780);
nand U3811 (N_3811,N_2471,N_2185);
and U3812 (N_3812,N_2714,N_2429);
xor U3813 (N_3813,N_2786,N_2141);
and U3814 (N_3814,N_2773,N_2241);
xor U3815 (N_3815,N_2172,N_2041);
xnor U3816 (N_3816,N_2359,N_2307);
or U3817 (N_3817,N_2224,N_2097);
xnor U3818 (N_3818,N_2787,N_2155);
xnor U3819 (N_3819,N_2733,N_2385);
and U3820 (N_3820,N_2695,N_2723);
nor U3821 (N_3821,N_2156,N_2942);
and U3822 (N_3822,N_2662,N_2755);
nand U3823 (N_3823,N_2477,N_2831);
and U3824 (N_3824,N_2856,N_2178);
and U3825 (N_3825,N_2368,N_2607);
nor U3826 (N_3826,N_2721,N_2786);
nand U3827 (N_3827,N_2930,N_2365);
nand U3828 (N_3828,N_2372,N_2416);
nor U3829 (N_3829,N_2489,N_2950);
and U3830 (N_3830,N_2375,N_2845);
or U3831 (N_3831,N_2868,N_2027);
and U3832 (N_3832,N_2506,N_2515);
nor U3833 (N_3833,N_2152,N_2705);
nand U3834 (N_3834,N_2825,N_2186);
nor U3835 (N_3835,N_2213,N_2632);
nand U3836 (N_3836,N_2362,N_2486);
nor U3837 (N_3837,N_2669,N_2014);
nor U3838 (N_3838,N_2249,N_2803);
and U3839 (N_3839,N_2051,N_2530);
and U3840 (N_3840,N_2744,N_2631);
nand U3841 (N_3841,N_2261,N_2930);
or U3842 (N_3842,N_2797,N_2227);
and U3843 (N_3843,N_2655,N_2725);
nor U3844 (N_3844,N_2361,N_2821);
and U3845 (N_3845,N_2177,N_2796);
or U3846 (N_3846,N_2759,N_2815);
and U3847 (N_3847,N_2594,N_2205);
nand U3848 (N_3848,N_2935,N_2771);
or U3849 (N_3849,N_2741,N_2058);
nand U3850 (N_3850,N_2277,N_2416);
and U3851 (N_3851,N_2397,N_2952);
and U3852 (N_3852,N_2321,N_2656);
or U3853 (N_3853,N_2343,N_2572);
nor U3854 (N_3854,N_2889,N_2430);
xnor U3855 (N_3855,N_2929,N_2830);
or U3856 (N_3856,N_2887,N_2667);
and U3857 (N_3857,N_2689,N_2036);
nor U3858 (N_3858,N_2160,N_2448);
nor U3859 (N_3859,N_2765,N_2324);
and U3860 (N_3860,N_2434,N_2114);
nand U3861 (N_3861,N_2980,N_2345);
and U3862 (N_3862,N_2642,N_2668);
and U3863 (N_3863,N_2690,N_2692);
nand U3864 (N_3864,N_2664,N_2332);
or U3865 (N_3865,N_2854,N_2182);
nor U3866 (N_3866,N_2759,N_2615);
nor U3867 (N_3867,N_2567,N_2120);
nand U3868 (N_3868,N_2380,N_2220);
nand U3869 (N_3869,N_2995,N_2706);
or U3870 (N_3870,N_2400,N_2647);
and U3871 (N_3871,N_2665,N_2814);
xnor U3872 (N_3872,N_2607,N_2126);
xor U3873 (N_3873,N_2358,N_2827);
nand U3874 (N_3874,N_2471,N_2172);
and U3875 (N_3875,N_2983,N_2961);
nand U3876 (N_3876,N_2778,N_2721);
nand U3877 (N_3877,N_2589,N_2769);
xnor U3878 (N_3878,N_2485,N_2309);
nand U3879 (N_3879,N_2801,N_2879);
nor U3880 (N_3880,N_2985,N_2338);
and U3881 (N_3881,N_2080,N_2798);
and U3882 (N_3882,N_2444,N_2206);
and U3883 (N_3883,N_2794,N_2336);
xnor U3884 (N_3884,N_2949,N_2813);
or U3885 (N_3885,N_2936,N_2108);
nor U3886 (N_3886,N_2819,N_2663);
nand U3887 (N_3887,N_2011,N_2194);
and U3888 (N_3888,N_2029,N_2181);
nor U3889 (N_3889,N_2108,N_2674);
nor U3890 (N_3890,N_2802,N_2294);
or U3891 (N_3891,N_2891,N_2268);
nand U3892 (N_3892,N_2170,N_2126);
xor U3893 (N_3893,N_2393,N_2866);
or U3894 (N_3894,N_2209,N_2908);
or U3895 (N_3895,N_2751,N_2084);
or U3896 (N_3896,N_2741,N_2630);
and U3897 (N_3897,N_2150,N_2768);
and U3898 (N_3898,N_2694,N_2011);
nor U3899 (N_3899,N_2338,N_2711);
and U3900 (N_3900,N_2652,N_2157);
nor U3901 (N_3901,N_2576,N_2183);
nor U3902 (N_3902,N_2059,N_2853);
nor U3903 (N_3903,N_2383,N_2656);
nand U3904 (N_3904,N_2924,N_2073);
and U3905 (N_3905,N_2556,N_2054);
nor U3906 (N_3906,N_2042,N_2824);
and U3907 (N_3907,N_2718,N_2689);
or U3908 (N_3908,N_2274,N_2181);
and U3909 (N_3909,N_2817,N_2408);
and U3910 (N_3910,N_2279,N_2771);
and U3911 (N_3911,N_2791,N_2755);
or U3912 (N_3912,N_2812,N_2161);
nor U3913 (N_3913,N_2239,N_2471);
and U3914 (N_3914,N_2769,N_2085);
nor U3915 (N_3915,N_2945,N_2946);
and U3916 (N_3916,N_2770,N_2682);
nor U3917 (N_3917,N_2393,N_2268);
or U3918 (N_3918,N_2718,N_2879);
nand U3919 (N_3919,N_2574,N_2615);
xnor U3920 (N_3920,N_2956,N_2131);
or U3921 (N_3921,N_2599,N_2062);
xor U3922 (N_3922,N_2543,N_2859);
or U3923 (N_3923,N_2796,N_2393);
or U3924 (N_3924,N_2474,N_2161);
nor U3925 (N_3925,N_2201,N_2780);
and U3926 (N_3926,N_2232,N_2172);
nor U3927 (N_3927,N_2379,N_2786);
nor U3928 (N_3928,N_2796,N_2770);
or U3929 (N_3929,N_2031,N_2065);
and U3930 (N_3930,N_2642,N_2411);
xor U3931 (N_3931,N_2769,N_2949);
nor U3932 (N_3932,N_2784,N_2002);
nand U3933 (N_3933,N_2752,N_2739);
or U3934 (N_3934,N_2449,N_2279);
nor U3935 (N_3935,N_2744,N_2808);
nor U3936 (N_3936,N_2694,N_2808);
or U3937 (N_3937,N_2677,N_2733);
nand U3938 (N_3938,N_2039,N_2196);
nand U3939 (N_3939,N_2860,N_2877);
nand U3940 (N_3940,N_2313,N_2068);
and U3941 (N_3941,N_2770,N_2296);
nor U3942 (N_3942,N_2087,N_2802);
nand U3943 (N_3943,N_2068,N_2809);
nand U3944 (N_3944,N_2002,N_2012);
nand U3945 (N_3945,N_2329,N_2788);
nor U3946 (N_3946,N_2899,N_2726);
nand U3947 (N_3947,N_2239,N_2190);
and U3948 (N_3948,N_2687,N_2388);
and U3949 (N_3949,N_2916,N_2244);
nor U3950 (N_3950,N_2871,N_2411);
and U3951 (N_3951,N_2560,N_2379);
or U3952 (N_3952,N_2805,N_2973);
and U3953 (N_3953,N_2416,N_2475);
and U3954 (N_3954,N_2446,N_2886);
nand U3955 (N_3955,N_2655,N_2979);
nand U3956 (N_3956,N_2408,N_2714);
or U3957 (N_3957,N_2444,N_2381);
or U3958 (N_3958,N_2867,N_2545);
or U3959 (N_3959,N_2673,N_2862);
xnor U3960 (N_3960,N_2610,N_2278);
nand U3961 (N_3961,N_2863,N_2776);
nand U3962 (N_3962,N_2865,N_2855);
xor U3963 (N_3963,N_2548,N_2019);
or U3964 (N_3964,N_2591,N_2715);
nand U3965 (N_3965,N_2423,N_2052);
or U3966 (N_3966,N_2717,N_2438);
nor U3967 (N_3967,N_2759,N_2627);
or U3968 (N_3968,N_2403,N_2045);
and U3969 (N_3969,N_2296,N_2583);
nor U3970 (N_3970,N_2834,N_2309);
xor U3971 (N_3971,N_2965,N_2404);
nand U3972 (N_3972,N_2956,N_2161);
nand U3973 (N_3973,N_2985,N_2644);
nand U3974 (N_3974,N_2477,N_2572);
and U3975 (N_3975,N_2169,N_2442);
nor U3976 (N_3976,N_2915,N_2533);
nor U3977 (N_3977,N_2790,N_2577);
nand U3978 (N_3978,N_2105,N_2003);
or U3979 (N_3979,N_2669,N_2382);
nor U3980 (N_3980,N_2651,N_2089);
xor U3981 (N_3981,N_2829,N_2393);
nor U3982 (N_3982,N_2348,N_2710);
and U3983 (N_3983,N_2763,N_2494);
nor U3984 (N_3984,N_2338,N_2360);
nor U3985 (N_3985,N_2844,N_2477);
or U3986 (N_3986,N_2458,N_2371);
or U3987 (N_3987,N_2135,N_2244);
nor U3988 (N_3988,N_2098,N_2207);
xor U3989 (N_3989,N_2927,N_2285);
and U3990 (N_3990,N_2341,N_2921);
nor U3991 (N_3991,N_2329,N_2670);
and U3992 (N_3992,N_2613,N_2741);
or U3993 (N_3993,N_2231,N_2770);
or U3994 (N_3994,N_2915,N_2268);
nor U3995 (N_3995,N_2332,N_2166);
nor U3996 (N_3996,N_2871,N_2981);
nand U3997 (N_3997,N_2578,N_2411);
and U3998 (N_3998,N_2859,N_2427);
nand U3999 (N_3999,N_2633,N_2119);
or U4000 (N_4000,N_3944,N_3889);
xor U4001 (N_4001,N_3192,N_3996);
nor U4002 (N_4002,N_3547,N_3954);
nor U4003 (N_4003,N_3785,N_3760);
or U4004 (N_4004,N_3541,N_3240);
and U4005 (N_4005,N_3712,N_3791);
and U4006 (N_4006,N_3136,N_3134);
nand U4007 (N_4007,N_3563,N_3465);
nand U4008 (N_4008,N_3918,N_3200);
xnor U4009 (N_4009,N_3025,N_3897);
and U4010 (N_4010,N_3925,N_3522);
or U4011 (N_4011,N_3038,N_3709);
nor U4012 (N_4012,N_3277,N_3949);
nand U4013 (N_4013,N_3969,N_3828);
nand U4014 (N_4014,N_3501,N_3135);
and U4015 (N_4015,N_3405,N_3759);
nand U4016 (N_4016,N_3885,N_3400);
nor U4017 (N_4017,N_3724,N_3109);
xor U4018 (N_4018,N_3890,N_3381);
and U4019 (N_4019,N_3372,N_3950);
and U4020 (N_4020,N_3713,N_3856);
or U4021 (N_4021,N_3325,N_3199);
nor U4022 (N_4022,N_3978,N_3887);
or U4023 (N_4023,N_3855,N_3682);
or U4024 (N_4024,N_3124,N_3018);
or U4025 (N_4025,N_3190,N_3297);
xor U4026 (N_4026,N_3171,N_3590);
nand U4027 (N_4027,N_3609,N_3464);
nor U4028 (N_4028,N_3274,N_3533);
or U4029 (N_4029,N_3451,N_3185);
or U4030 (N_4030,N_3482,N_3496);
nand U4031 (N_4031,N_3706,N_3387);
nand U4032 (N_4032,N_3064,N_3284);
nor U4033 (N_4033,N_3896,N_3378);
or U4034 (N_4034,N_3061,N_3304);
nor U4035 (N_4035,N_3768,N_3193);
and U4036 (N_4036,N_3567,N_3060);
nor U4037 (N_4037,N_3101,N_3253);
and U4038 (N_4038,N_3529,N_3764);
and U4039 (N_4039,N_3259,N_3014);
nor U4040 (N_4040,N_3086,N_3396);
nor U4041 (N_4041,N_3234,N_3801);
nor U4042 (N_4042,N_3227,N_3849);
or U4043 (N_4043,N_3099,N_3532);
or U4044 (N_4044,N_3265,N_3915);
and U4045 (N_4045,N_3539,N_3467);
nor U4046 (N_4046,N_3556,N_3043);
and U4047 (N_4047,N_3231,N_3758);
nand U4048 (N_4048,N_3137,N_3080);
nor U4049 (N_4049,N_3814,N_3865);
nor U4050 (N_4050,N_3521,N_3557);
and U4051 (N_4051,N_3312,N_3302);
nor U4052 (N_4052,N_3543,N_3347);
nor U4053 (N_4053,N_3797,N_3870);
nand U4054 (N_4054,N_3667,N_3775);
nand U4055 (N_4055,N_3275,N_3412);
xnor U4056 (N_4056,N_3631,N_3421);
and U4057 (N_4057,N_3119,N_3391);
or U4058 (N_4058,N_3219,N_3177);
or U4059 (N_4059,N_3348,N_3009);
nor U4060 (N_4060,N_3030,N_3360);
or U4061 (N_4061,N_3685,N_3019);
or U4062 (N_4062,N_3049,N_3242);
xnor U4063 (N_4063,N_3359,N_3409);
xnor U4064 (N_4064,N_3904,N_3401);
or U4065 (N_4065,N_3224,N_3504);
and U4066 (N_4066,N_3763,N_3634);
or U4067 (N_4067,N_3702,N_3938);
and U4068 (N_4068,N_3746,N_3001);
and U4069 (N_4069,N_3975,N_3537);
nor U4070 (N_4070,N_3620,N_3053);
nor U4071 (N_4071,N_3819,N_3926);
or U4072 (N_4072,N_3373,N_3735);
nor U4073 (N_4073,N_3542,N_3357);
nor U4074 (N_4074,N_3477,N_3612);
and U4075 (N_4075,N_3248,N_3050);
or U4076 (N_4076,N_3204,N_3241);
nor U4077 (N_4077,N_3509,N_3784);
or U4078 (N_4078,N_3292,N_3494);
nor U4079 (N_4079,N_3168,N_3438);
nor U4080 (N_4080,N_3389,N_3638);
nand U4081 (N_4081,N_3349,N_3629);
nor U4082 (N_4082,N_3106,N_3803);
nand U4083 (N_4083,N_3850,N_3102);
and U4084 (N_4084,N_3796,N_3771);
or U4085 (N_4085,N_3573,N_3930);
nor U4086 (N_4086,N_3643,N_3042);
or U4087 (N_4087,N_3316,N_3600);
or U4088 (N_4088,N_3914,N_3144);
nor U4089 (N_4089,N_3225,N_3603);
nand U4090 (N_4090,N_3447,N_3490);
nor U4091 (N_4091,N_3344,N_3187);
and U4092 (N_4092,N_3617,N_3008);
xor U4093 (N_4093,N_3103,N_3805);
or U4094 (N_4094,N_3485,N_3321);
xnor U4095 (N_4095,N_3569,N_3689);
nor U4096 (N_4096,N_3059,N_3720);
nand U4097 (N_4097,N_3630,N_3082);
nor U4098 (N_4098,N_3153,N_3941);
or U4099 (N_4099,N_3305,N_3880);
nand U4100 (N_4100,N_3829,N_3523);
nor U4101 (N_4101,N_3395,N_3728);
and U4102 (N_4102,N_3211,N_3363);
or U4103 (N_4103,N_3096,N_3005);
nor U4104 (N_4104,N_3595,N_3318);
nand U4105 (N_4105,N_3752,N_3633);
and U4106 (N_4106,N_3139,N_3761);
nand U4107 (N_4107,N_3650,N_3962);
or U4108 (N_4108,N_3141,N_3430);
and U4109 (N_4109,N_3085,N_3794);
and U4110 (N_4110,N_3879,N_3597);
nor U4111 (N_4111,N_3466,N_3236);
nand U4112 (N_4112,N_3841,N_3959);
and U4113 (N_4113,N_3252,N_3498);
or U4114 (N_4114,N_3118,N_3860);
nand U4115 (N_4115,N_3123,N_3847);
nor U4116 (N_4116,N_3753,N_3964);
and U4117 (N_4117,N_3779,N_3218);
nor U4118 (N_4118,N_3152,N_3448);
nor U4119 (N_4119,N_3007,N_3672);
or U4120 (N_4120,N_3489,N_3770);
nor U4121 (N_4121,N_3296,N_3436);
nand U4122 (N_4122,N_3486,N_3356);
xnor U4123 (N_4123,N_3756,N_3881);
nand U4124 (N_4124,N_3546,N_3121);
and U4125 (N_4125,N_3966,N_3151);
nand U4126 (N_4126,N_3974,N_3361);
and U4127 (N_4127,N_3655,N_3181);
and U4128 (N_4128,N_3116,N_3868);
nor U4129 (N_4129,N_3524,N_3016);
nor U4130 (N_4130,N_3488,N_3766);
xnor U4131 (N_4131,N_3992,N_3876);
xor U4132 (N_4132,N_3149,N_3867);
or U4133 (N_4133,N_3342,N_3510);
nor U4134 (N_4134,N_3044,N_3100);
nand U4135 (N_4135,N_3223,N_3769);
nor U4136 (N_4136,N_3972,N_3422);
xnor U4137 (N_4137,N_3800,N_3472);
and U4138 (N_4138,N_3194,N_3145);
xnor U4139 (N_4139,N_3767,N_3861);
nor U4140 (N_4140,N_3632,N_3163);
and U4141 (N_4141,N_3207,N_3502);
nor U4142 (N_4142,N_3783,N_3201);
and U4143 (N_4143,N_3550,N_3062);
xor U4144 (N_4144,N_3343,N_3704);
nand U4145 (N_4145,N_3948,N_3257);
or U4146 (N_4146,N_3452,N_3947);
xor U4147 (N_4147,N_3983,N_3439);
nor U4148 (N_4148,N_3802,N_3538);
nand U4149 (N_4149,N_3815,N_3913);
xor U4150 (N_4150,N_3246,N_3984);
nand U4151 (N_4151,N_3455,N_3507);
nor U4152 (N_4152,N_3513,N_3916);
xnor U4153 (N_4153,N_3084,N_3694);
and U4154 (N_4154,N_3751,N_3536);
nand U4155 (N_4155,N_3491,N_3888);
and U4156 (N_4156,N_3492,N_3776);
nand U4157 (N_4157,N_3970,N_3046);
or U4158 (N_4158,N_3433,N_3744);
nand U4159 (N_4159,N_3671,N_3923);
nand U4160 (N_4160,N_3040,N_3982);
xor U4161 (N_4161,N_3055,N_3935);
or U4162 (N_4162,N_3125,N_3745);
and U4163 (N_4163,N_3262,N_3777);
nor U4164 (N_4164,N_3045,N_3379);
nor U4165 (N_4165,N_3514,N_3127);
nor U4166 (N_4166,N_3355,N_3731);
or U4167 (N_4167,N_3585,N_3213);
or U4168 (N_4168,N_3495,N_3812);
and U4169 (N_4169,N_3107,N_3786);
nand U4170 (N_4170,N_3138,N_3933);
and U4171 (N_4171,N_3673,N_3251);
or U4172 (N_4172,N_3503,N_3002);
or U4173 (N_4173,N_3220,N_3471);
nor U4174 (N_4174,N_3010,N_3073);
or U4175 (N_4175,N_3303,N_3233);
nor U4176 (N_4176,N_3150,N_3416);
nor U4177 (N_4177,N_3155,N_3353);
nand U4178 (N_4178,N_3454,N_3475);
or U4179 (N_4179,N_3813,N_3376);
and U4180 (N_4180,N_3352,N_3266);
nor U4181 (N_4181,N_3574,N_3140);
and U4182 (N_4182,N_3039,N_3268);
nand U4183 (N_4183,N_3858,N_3540);
and U4184 (N_4184,N_3057,N_3269);
or U4185 (N_4185,N_3512,N_3029);
nor U4186 (N_4186,N_3608,N_3877);
and U4187 (N_4187,N_3826,N_3095);
or U4188 (N_4188,N_3075,N_3657);
nor U4189 (N_4189,N_3216,N_3000);
and U4190 (N_4190,N_3698,N_3903);
nor U4191 (N_4191,N_3725,N_3535);
or U4192 (N_4192,N_3651,N_3956);
and U4193 (N_4193,N_3239,N_3210);
nor U4194 (N_4194,N_3300,N_3998);
nand U4195 (N_4195,N_3179,N_3517);
or U4196 (N_4196,N_3559,N_3399);
and U4197 (N_4197,N_3505,N_3474);
or U4198 (N_4198,N_3660,N_3738);
nor U4199 (N_4199,N_3161,N_3639);
nand U4200 (N_4200,N_3159,N_3957);
xor U4201 (N_4201,N_3074,N_3782);
and U4202 (N_4202,N_3202,N_3684);
nand U4203 (N_4203,N_3696,N_3825);
or U4204 (N_4204,N_3048,N_3866);
nand U4205 (N_4205,N_3607,N_3058);
nand U4206 (N_4206,N_3129,N_3324);
and U4207 (N_4207,N_3079,N_3111);
and U4208 (N_4208,N_3531,N_3027);
and U4209 (N_4209,N_3308,N_3368);
nand U4210 (N_4210,N_3205,N_3988);
nand U4211 (N_4211,N_3656,N_3332);
or U4212 (N_4212,N_3250,N_3051);
or U4213 (N_4213,N_3928,N_3747);
xor U4214 (N_4214,N_3716,N_3328);
nand U4215 (N_4215,N_3967,N_3664);
and U4216 (N_4216,N_3895,N_3034);
and U4217 (N_4217,N_3424,N_3024);
xor U4218 (N_4218,N_3593,N_3162);
and U4219 (N_4219,N_3549,N_3417);
or U4220 (N_4220,N_3874,N_3461);
nand U4221 (N_4221,N_3288,N_3968);
nor U4222 (N_4222,N_3670,N_3640);
and U4223 (N_4223,N_3852,N_3271);
nand U4224 (N_4224,N_3428,N_3339);
nor U4225 (N_4225,N_3217,N_3555);
and U4226 (N_4226,N_3568,N_3104);
or U4227 (N_4227,N_3626,N_3221);
nor U4228 (N_4228,N_3483,N_3208);
or U4229 (N_4229,N_3781,N_3649);
or U4230 (N_4230,N_3936,N_3133);
nand U4231 (N_4231,N_3445,N_3203);
nor U4232 (N_4232,N_3798,N_3911);
nor U4233 (N_4233,N_3098,N_3666);
nand U4234 (N_4234,N_3884,N_3619);
nand U4235 (N_4235,N_3307,N_3054);
nand U4236 (N_4236,N_3859,N_3661);
nor U4237 (N_4237,N_3037,N_3088);
nor U4238 (N_4238,N_3375,N_3601);
and U4239 (N_4239,N_3922,N_3249);
nand U4240 (N_4240,N_3367,N_3799);
and U4241 (N_4241,N_3699,N_3830);
or U4242 (N_4242,N_3420,N_3069);
xnor U4243 (N_4243,N_3319,N_3165);
nand U4244 (N_4244,N_3806,N_3762);
xor U4245 (N_4245,N_3929,N_3157);
or U4246 (N_4246,N_3989,N_3299);
and U4247 (N_4247,N_3519,N_3668);
nand U4248 (N_4248,N_3708,N_3460);
and U4249 (N_4249,N_3117,N_3662);
nor U4250 (N_4250,N_3792,N_3579);
or U4251 (N_4251,N_3390,N_3456);
or U4252 (N_4252,N_3337,N_3435);
xnor U4253 (N_4253,N_3077,N_3026);
nor U4254 (N_4254,N_3446,N_3571);
or U4255 (N_4255,N_3818,N_3330);
or U4256 (N_4256,N_3642,N_3329);
nand U4257 (N_4257,N_3473,N_3370);
xor U4258 (N_4258,N_3680,N_3089);
or U4259 (N_4259,N_3908,N_3953);
or U4260 (N_4260,N_3015,N_3173);
nand U4261 (N_4261,N_3614,N_3900);
nor U4262 (N_4262,N_3919,N_3743);
or U4263 (N_4263,N_3833,N_3222);
or U4264 (N_4264,N_3028,N_3577);
nand U4265 (N_4265,N_3591,N_3552);
and U4266 (N_4266,N_3920,N_3710);
xnor U4267 (N_4267,N_3602,N_3065);
or U4268 (N_4268,N_3354,N_3824);
nor U4269 (N_4269,N_3291,N_3973);
and U4270 (N_4270,N_3875,N_3912);
nand U4271 (N_4271,N_3226,N_3398);
or U4272 (N_4272,N_3723,N_3737);
xnor U4273 (N_4273,N_3857,N_3156);
nor U4274 (N_4274,N_3658,N_3838);
and U4275 (N_4275,N_3130,N_3939);
or U4276 (N_4276,N_3063,N_3429);
xor U4277 (N_4277,N_3835,N_3851);
xnor U4278 (N_4278,N_3081,N_3917);
nand U4279 (N_4279,N_3839,N_3122);
or U4280 (N_4280,N_3176,N_3963);
nor U4281 (N_4281,N_3440,N_3976);
or U4282 (N_4282,N_3148,N_3613);
and U4283 (N_4283,N_3289,N_3182);
xor U4284 (N_4284,N_3545,N_3644);
nand U4285 (N_4285,N_3693,N_3663);
and U4286 (N_4286,N_3506,N_3290);
nand U4287 (N_4287,N_3722,N_3114);
and U4288 (N_4288,N_3645,N_3235);
and U4289 (N_4289,N_3434,N_3309);
nand U4290 (N_4290,N_3615,N_3022);
or U4291 (N_4291,N_3484,N_3554);
or U4292 (N_4292,N_3618,N_3237);
or U4293 (N_4293,N_3413,N_3817);
nand U4294 (N_4294,N_3611,N_3115);
xor U4295 (N_4295,N_3047,N_3515);
or U4296 (N_4296,N_3703,N_3788);
or U4297 (N_4297,N_3891,N_3654);
or U4298 (N_4298,N_3254,N_3131);
and U4299 (N_4299,N_3286,N_3596);
nand U4300 (N_4300,N_3346,N_3997);
and U4301 (N_4301,N_3311,N_3604);
nand U4302 (N_4302,N_3285,N_3843);
or U4303 (N_4303,N_3993,N_3091);
nand U4304 (N_4304,N_3278,N_3273);
and U4305 (N_4305,N_3906,N_3909);
xnor U4306 (N_4306,N_3755,N_3527);
nand U4307 (N_4307,N_3358,N_3772);
or U4308 (N_4308,N_3132,N_3493);
or U4309 (N_4309,N_3822,N_3006);
xnor U4310 (N_4310,N_3985,N_3943);
or U4311 (N_4311,N_3842,N_3481);
nor U4312 (N_4312,N_3675,N_3083);
or U4313 (N_4313,N_3314,N_3711);
nand U4314 (N_4314,N_3478,N_3071);
and U4315 (N_4315,N_3598,N_3012);
and U4316 (N_4316,N_3374,N_3191);
or U4317 (N_4317,N_3076,N_3659);
or U4318 (N_4318,N_3572,N_3740);
and U4319 (N_4319,N_3036,N_3816);
nor U4320 (N_4320,N_3653,N_3566);
or U4321 (N_4321,N_3470,N_3587);
nand U4322 (N_4322,N_3317,N_3393);
nor U4323 (N_4323,N_3905,N_3279);
nand U4324 (N_4324,N_3691,N_3586);
and U4325 (N_4325,N_3092,N_3748);
xor U4326 (N_4326,N_3683,N_3754);
nor U4327 (N_4327,N_3707,N_3576);
and U4328 (N_4328,N_3789,N_3459);
nor U4329 (N_4329,N_3369,N_3994);
and U4330 (N_4330,N_3831,N_3195);
xor U4331 (N_4331,N_3690,N_3678);
nand U4332 (N_4332,N_3588,N_3212);
xor U4333 (N_4333,N_3174,N_3003);
nand U4334 (N_4334,N_3322,N_3366);
and U4335 (N_4335,N_3741,N_3610);
nand U4336 (N_4336,N_3726,N_3031);
and U4337 (N_4337,N_3561,N_3415);
and U4338 (N_4338,N_3564,N_3158);
nor U4339 (N_4339,N_3108,N_3320);
nand U4340 (N_4340,N_3589,N_3719);
nand U4341 (N_4341,N_3910,N_3450);
nor U4342 (N_4342,N_3298,N_3844);
nand U4343 (N_4343,N_3810,N_3377);
and U4344 (N_4344,N_3261,N_3907);
or U4345 (N_4345,N_3872,N_3423);
nor U4346 (N_4346,N_3511,N_3469);
nor U4347 (N_4347,N_3727,N_3625);
and U4348 (N_4348,N_3848,N_3977);
xor U4349 (N_4349,N_3739,N_3147);
and U4350 (N_4350,N_3990,N_3499);
and U4351 (N_4351,N_3110,N_3442);
and U4352 (N_4352,N_3999,N_3583);
or U4353 (N_4353,N_3468,N_3067);
nor U4354 (N_4354,N_3697,N_3169);
or U4355 (N_4355,N_3313,N_3804);
or U4356 (N_4356,N_3232,N_3773);
nand U4357 (N_4357,N_3364,N_3636);
nand U4358 (N_4358,N_3351,N_3862);
or U4359 (N_4359,N_3899,N_3394);
xnor U4360 (N_4360,N_3705,N_3384);
nand U4361 (N_4361,N_3827,N_3004);
or U4362 (N_4362,N_3945,N_3293);
and U4363 (N_4363,N_3677,N_3411);
nor U4364 (N_4364,N_3942,N_3525);
or U4365 (N_4365,N_3853,N_3560);
nor U4366 (N_4366,N_3627,N_3154);
and U4367 (N_4367,N_3338,N_3732);
and U4368 (N_4368,N_3334,N_3443);
nor U4369 (N_4369,N_3624,N_3981);
xnor U4370 (N_4370,N_3404,N_3457);
nand U4371 (N_4371,N_3834,N_3243);
or U4372 (N_4372,N_3570,N_3476);
nor U4373 (N_4373,N_3898,N_3184);
nand U4374 (N_4374,N_3635,N_3845);
nand U4375 (N_4375,N_3701,N_3458);
and U4376 (N_4376,N_3894,N_3534);
or U4377 (N_4377,N_3017,N_3143);
and U4378 (N_4378,N_3365,N_3164);
nand U4379 (N_4379,N_3808,N_3955);
nor U4380 (N_4380,N_3120,N_3392);
xnor U4381 (N_4381,N_3175,N_3991);
and U4382 (N_4382,N_3196,N_3960);
and U4383 (N_4383,N_3616,N_3979);
or U4384 (N_4384,N_3530,N_3385);
xnor U4385 (N_4385,N_3883,N_3315);
nand U4386 (N_4386,N_3528,N_3951);
nor U4387 (N_4387,N_3410,N_3362);
and U4388 (N_4388,N_3688,N_3052);
and U4389 (N_4389,N_3652,N_3382);
nor U4390 (N_4390,N_3444,N_3295);
nand U4391 (N_4391,N_3715,N_3987);
and U4392 (N_4392,N_3733,N_3160);
and U4393 (N_4393,N_3245,N_3331);
nand U4394 (N_4394,N_3840,N_3934);
or U4395 (N_4395,N_3070,N_3787);
nand U4396 (N_4396,N_3749,N_3270);
nand U4397 (N_4397,N_3345,N_3425);
nor U4398 (N_4398,N_3508,N_3790);
xor U4399 (N_4399,N_3820,N_3255);
nand U4400 (N_4400,N_3282,N_3878);
nand U4401 (N_4401,N_3700,N_3695);
and U4402 (N_4402,N_3449,N_3686);
or U4403 (N_4403,N_3674,N_3341);
xnor U4404 (N_4404,N_3562,N_3692);
xor U4405 (N_4405,N_3821,N_3648);
xor U4406 (N_4406,N_3582,N_3407);
or U4407 (N_4407,N_3869,N_3170);
or U4408 (N_4408,N_3441,N_3462);
and U4409 (N_4409,N_3995,N_3628);
nand U4410 (N_4410,N_3621,N_3599);
or U4411 (N_4411,N_3260,N_3729);
nand U4412 (N_4412,N_3340,N_3742);
xnor U4413 (N_4413,N_3426,N_3553);
nor U4414 (N_4414,N_3020,N_3244);
nor U4415 (N_4415,N_3453,N_3066);
nor U4416 (N_4416,N_3846,N_3924);
nor U4417 (N_4417,N_3350,N_3606);
or U4418 (N_4418,N_3669,N_3778);
nor U4419 (N_4419,N_3500,N_3952);
nor U4420 (N_4420,N_3078,N_3971);
xor U4421 (N_4421,N_3837,N_3718);
nor U4422 (N_4422,N_3836,N_3605);
xnor U4423 (N_4423,N_3097,N_3780);
nor U4424 (N_4424,N_3397,N_3487);
nor U4425 (N_4425,N_3437,N_3310);
and U4426 (N_4426,N_3230,N_3301);
nor U4427 (N_4427,N_3811,N_3188);
nor U4428 (N_4428,N_3750,N_3765);
or U4429 (N_4429,N_3823,N_3276);
or U4430 (N_4430,N_3565,N_3093);
nor U4431 (N_4431,N_3258,N_3105);
xor U4432 (N_4432,N_3166,N_3383);
nor U4433 (N_4433,N_3056,N_3637);
and U4434 (N_4434,N_3902,N_3209);
or U4435 (N_4435,N_3526,N_3371);
nand U4436 (N_4436,N_3544,N_3714);
and U4437 (N_4437,N_3113,N_3730);
xor U4438 (N_4438,N_3641,N_3665);
xnor U4439 (N_4439,N_3335,N_3263);
nand U4440 (N_4440,N_3734,N_3035);
and U4441 (N_4441,N_3578,N_3551);
xor U4442 (N_4442,N_3418,N_3336);
and U4443 (N_4443,N_3594,N_3189);
nor U4444 (N_4444,N_3087,N_3832);
or U4445 (N_4445,N_3272,N_3592);
xnor U4446 (N_4446,N_3326,N_3264);
or U4447 (N_4447,N_3229,N_3516);
nor U4448 (N_4448,N_3146,N_3558);
and U4449 (N_4449,N_3402,N_3721);
and U4450 (N_4450,N_3893,N_3901);
and U4451 (N_4451,N_3921,N_3927);
or U4452 (N_4452,N_3306,N_3873);
and U4453 (N_4453,N_3623,N_3167);
and U4454 (N_4454,N_3965,N_3520);
nand U4455 (N_4455,N_3882,N_3807);
nand U4456 (N_4456,N_3283,N_3333);
nand U4457 (N_4457,N_3932,N_3403);
or U4458 (N_4458,N_3432,N_3215);
or U4459 (N_4459,N_3480,N_3958);
or U4460 (N_4460,N_3575,N_3681);
xor U4461 (N_4461,N_3041,N_3774);
nor U4462 (N_4462,N_3622,N_3183);
or U4463 (N_4463,N_3580,N_3946);
or U4464 (N_4464,N_3267,N_3679);
and U4465 (N_4465,N_3198,N_3406);
nand U4466 (N_4466,N_3736,N_3238);
and U4467 (N_4467,N_3793,N_3548);
and U4468 (N_4468,N_3795,N_3871);
and U4469 (N_4469,N_3986,N_3419);
xnor U4470 (N_4470,N_3646,N_3937);
nor U4471 (N_4471,N_3126,N_3427);
and U4472 (N_4472,N_3584,N_3180);
xor U4473 (N_4473,N_3072,N_3886);
nor U4474 (N_4474,N_3931,N_3256);
and U4475 (N_4475,N_3033,N_3287);
nor U4476 (N_4476,N_3128,N_3388);
or U4477 (N_4477,N_3228,N_3214);
nor U4478 (N_4478,N_3479,N_3961);
nand U4479 (N_4479,N_3380,N_3408);
nor U4480 (N_4480,N_3178,N_3980);
and U4481 (N_4481,N_3172,N_3864);
nand U4482 (N_4482,N_3247,N_3281);
nor U4483 (N_4483,N_3647,N_3717);
or U4484 (N_4484,N_3327,N_3581);
and U4485 (N_4485,N_3068,N_3021);
xor U4486 (N_4486,N_3090,N_3863);
xor U4487 (N_4487,N_3023,N_3809);
and U4488 (N_4488,N_3414,N_3094);
nor U4489 (N_4489,N_3431,N_3186);
or U4490 (N_4490,N_3687,N_3386);
nand U4491 (N_4491,N_3940,N_3463);
or U4492 (N_4492,N_3013,N_3280);
xnor U4493 (N_4493,N_3497,N_3112);
xnor U4494 (N_4494,N_3323,N_3518);
nor U4495 (N_4495,N_3011,N_3032);
or U4496 (N_4496,N_3676,N_3892);
nor U4497 (N_4497,N_3757,N_3854);
nor U4498 (N_4498,N_3197,N_3142);
nand U4499 (N_4499,N_3294,N_3206);
and U4500 (N_4500,N_3622,N_3538);
or U4501 (N_4501,N_3771,N_3753);
or U4502 (N_4502,N_3574,N_3459);
nand U4503 (N_4503,N_3651,N_3112);
xor U4504 (N_4504,N_3832,N_3300);
or U4505 (N_4505,N_3368,N_3552);
and U4506 (N_4506,N_3358,N_3444);
and U4507 (N_4507,N_3604,N_3510);
or U4508 (N_4508,N_3946,N_3083);
and U4509 (N_4509,N_3324,N_3467);
or U4510 (N_4510,N_3177,N_3855);
or U4511 (N_4511,N_3507,N_3395);
nor U4512 (N_4512,N_3217,N_3423);
or U4513 (N_4513,N_3330,N_3787);
nor U4514 (N_4514,N_3514,N_3551);
nand U4515 (N_4515,N_3832,N_3607);
nand U4516 (N_4516,N_3340,N_3849);
or U4517 (N_4517,N_3006,N_3173);
or U4518 (N_4518,N_3196,N_3648);
or U4519 (N_4519,N_3905,N_3704);
xnor U4520 (N_4520,N_3628,N_3656);
nor U4521 (N_4521,N_3704,N_3577);
and U4522 (N_4522,N_3613,N_3716);
or U4523 (N_4523,N_3808,N_3329);
nor U4524 (N_4524,N_3847,N_3098);
or U4525 (N_4525,N_3099,N_3220);
nor U4526 (N_4526,N_3232,N_3373);
and U4527 (N_4527,N_3995,N_3973);
nor U4528 (N_4528,N_3059,N_3793);
nand U4529 (N_4529,N_3526,N_3363);
and U4530 (N_4530,N_3336,N_3937);
xor U4531 (N_4531,N_3337,N_3814);
nand U4532 (N_4532,N_3812,N_3846);
xnor U4533 (N_4533,N_3728,N_3712);
or U4534 (N_4534,N_3334,N_3889);
or U4535 (N_4535,N_3318,N_3321);
xnor U4536 (N_4536,N_3134,N_3782);
and U4537 (N_4537,N_3829,N_3091);
or U4538 (N_4538,N_3524,N_3653);
nor U4539 (N_4539,N_3277,N_3096);
and U4540 (N_4540,N_3868,N_3424);
and U4541 (N_4541,N_3528,N_3091);
or U4542 (N_4542,N_3080,N_3730);
nor U4543 (N_4543,N_3923,N_3866);
nand U4544 (N_4544,N_3683,N_3579);
or U4545 (N_4545,N_3852,N_3011);
nand U4546 (N_4546,N_3200,N_3527);
or U4547 (N_4547,N_3581,N_3144);
and U4548 (N_4548,N_3197,N_3637);
nand U4549 (N_4549,N_3778,N_3500);
or U4550 (N_4550,N_3420,N_3594);
nor U4551 (N_4551,N_3888,N_3504);
xnor U4552 (N_4552,N_3155,N_3364);
nor U4553 (N_4553,N_3223,N_3997);
nand U4554 (N_4554,N_3135,N_3979);
nand U4555 (N_4555,N_3431,N_3882);
nand U4556 (N_4556,N_3140,N_3370);
xnor U4557 (N_4557,N_3025,N_3654);
nand U4558 (N_4558,N_3624,N_3742);
or U4559 (N_4559,N_3487,N_3951);
nand U4560 (N_4560,N_3786,N_3205);
xnor U4561 (N_4561,N_3335,N_3501);
nor U4562 (N_4562,N_3674,N_3468);
nor U4563 (N_4563,N_3013,N_3035);
nor U4564 (N_4564,N_3401,N_3877);
and U4565 (N_4565,N_3649,N_3325);
nand U4566 (N_4566,N_3616,N_3342);
nor U4567 (N_4567,N_3454,N_3810);
or U4568 (N_4568,N_3937,N_3835);
nand U4569 (N_4569,N_3923,N_3889);
and U4570 (N_4570,N_3139,N_3507);
nand U4571 (N_4571,N_3529,N_3976);
and U4572 (N_4572,N_3610,N_3439);
nand U4573 (N_4573,N_3917,N_3343);
or U4574 (N_4574,N_3770,N_3961);
and U4575 (N_4575,N_3083,N_3823);
nor U4576 (N_4576,N_3908,N_3565);
and U4577 (N_4577,N_3258,N_3754);
and U4578 (N_4578,N_3996,N_3249);
or U4579 (N_4579,N_3477,N_3757);
nand U4580 (N_4580,N_3540,N_3890);
nor U4581 (N_4581,N_3408,N_3199);
nand U4582 (N_4582,N_3269,N_3080);
or U4583 (N_4583,N_3657,N_3432);
or U4584 (N_4584,N_3887,N_3851);
or U4585 (N_4585,N_3161,N_3055);
or U4586 (N_4586,N_3488,N_3840);
nand U4587 (N_4587,N_3541,N_3250);
and U4588 (N_4588,N_3114,N_3767);
nand U4589 (N_4589,N_3392,N_3416);
nor U4590 (N_4590,N_3943,N_3912);
nor U4591 (N_4591,N_3779,N_3513);
or U4592 (N_4592,N_3102,N_3735);
or U4593 (N_4593,N_3223,N_3452);
and U4594 (N_4594,N_3699,N_3736);
nand U4595 (N_4595,N_3879,N_3905);
or U4596 (N_4596,N_3521,N_3073);
or U4597 (N_4597,N_3778,N_3975);
or U4598 (N_4598,N_3428,N_3742);
nand U4599 (N_4599,N_3408,N_3048);
nand U4600 (N_4600,N_3980,N_3326);
nand U4601 (N_4601,N_3305,N_3942);
or U4602 (N_4602,N_3638,N_3479);
nor U4603 (N_4603,N_3474,N_3976);
nor U4604 (N_4604,N_3020,N_3280);
or U4605 (N_4605,N_3190,N_3784);
nand U4606 (N_4606,N_3108,N_3814);
nor U4607 (N_4607,N_3351,N_3003);
nand U4608 (N_4608,N_3505,N_3999);
nor U4609 (N_4609,N_3522,N_3053);
or U4610 (N_4610,N_3947,N_3342);
nor U4611 (N_4611,N_3920,N_3489);
nor U4612 (N_4612,N_3748,N_3583);
or U4613 (N_4613,N_3890,N_3883);
or U4614 (N_4614,N_3123,N_3589);
and U4615 (N_4615,N_3590,N_3179);
nor U4616 (N_4616,N_3293,N_3354);
nor U4617 (N_4617,N_3953,N_3346);
nand U4618 (N_4618,N_3659,N_3965);
nor U4619 (N_4619,N_3482,N_3837);
or U4620 (N_4620,N_3322,N_3408);
or U4621 (N_4621,N_3037,N_3308);
nor U4622 (N_4622,N_3762,N_3373);
nor U4623 (N_4623,N_3406,N_3718);
nor U4624 (N_4624,N_3102,N_3440);
nand U4625 (N_4625,N_3100,N_3517);
nor U4626 (N_4626,N_3222,N_3976);
and U4627 (N_4627,N_3194,N_3391);
nor U4628 (N_4628,N_3995,N_3593);
nand U4629 (N_4629,N_3843,N_3906);
nand U4630 (N_4630,N_3544,N_3359);
nor U4631 (N_4631,N_3398,N_3127);
nor U4632 (N_4632,N_3504,N_3191);
nand U4633 (N_4633,N_3122,N_3636);
nand U4634 (N_4634,N_3843,N_3336);
nor U4635 (N_4635,N_3869,N_3564);
nand U4636 (N_4636,N_3717,N_3710);
nor U4637 (N_4637,N_3632,N_3011);
xor U4638 (N_4638,N_3992,N_3610);
nor U4639 (N_4639,N_3436,N_3509);
xnor U4640 (N_4640,N_3365,N_3348);
xnor U4641 (N_4641,N_3336,N_3389);
nor U4642 (N_4642,N_3882,N_3360);
nand U4643 (N_4643,N_3793,N_3833);
or U4644 (N_4644,N_3758,N_3458);
nand U4645 (N_4645,N_3036,N_3039);
or U4646 (N_4646,N_3952,N_3019);
or U4647 (N_4647,N_3964,N_3507);
and U4648 (N_4648,N_3783,N_3090);
and U4649 (N_4649,N_3653,N_3862);
nor U4650 (N_4650,N_3950,N_3967);
and U4651 (N_4651,N_3427,N_3876);
or U4652 (N_4652,N_3266,N_3947);
and U4653 (N_4653,N_3572,N_3709);
or U4654 (N_4654,N_3473,N_3826);
nand U4655 (N_4655,N_3132,N_3637);
xnor U4656 (N_4656,N_3816,N_3338);
and U4657 (N_4657,N_3179,N_3239);
xor U4658 (N_4658,N_3433,N_3939);
or U4659 (N_4659,N_3845,N_3019);
or U4660 (N_4660,N_3531,N_3748);
xor U4661 (N_4661,N_3038,N_3831);
nor U4662 (N_4662,N_3366,N_3555);
nor U4663 (N_4663,N_3068,N_3440);
or U4664 (N_4664,N_3001,N_3604);
nor U4665 (N_4665,N_3510,N_3196);
and U4666 (N_4666,N_3250,N_3977);
nor U4667 (N_4667,N_3998,N_3727);
xnor U4668 (N_4668,N_3912,N_3876);
xor U4669 (N_4669,N_3971,N_3123);
nand U4670 (N_4670,N_3766,N_3818);
and U4671 (N_4671,N_3797,N_3004);
or U4672 (N_4672,N_3647,N_3640);
or U4673 (N_4673,N_3361,N_3876);
nand U4674 (N_4674,N_3412,N_3187);
or U4675 (N_4675,N_3527,N_3343);
and U4676 (N_4676,N_3089,N_3021);
and U4677 (N_4677,N_3085,N_3555);
nor U4678 (N_4678,N_3440,N_3279);
or U4679 (N_4679,N_3459,N_3576);
and U4680 (N_4680,N_3801,N_3857);
xnor U4681 (N_4681,N_3682,N_3600);
and U4682 (N_4682,N_3035,N_3709);
nand U4683 (N_4683,N_3579,N_3696);
and U4684 (N_4684,N_3476,N_3664);
nor U4685 (N_4685,N_3516,N_3175);
and U4686 (N_4686,N_3373,N_3241);
and U4687 (N_4687,N_3155,N_3519);
and U4688 (N_4688,N_3529,N_3162);
nor U4689 (N_4689,N_3206,N_3506);
and U4690 (N_4690,N_3792,N_3392);
or U4691 (N_4691,N_3180,N_3258);
nand U4692 (N_4692,N_3389,N_3606);
and U4693 (N_4693,N_3090,N_3546);
nor U4694 (N_4694,N_3454,N_3728);
and U4695 (N_4695,N_3900,N_3535);
and U4696 (N_4696,N_3454,N_3546);
nor U4697 (N_4697,N_3094,N_3022);
nor U4698 (N_4698,N_3335,N_3422);
nand U4699 (N_4699,N_3937,N_3363);
or U4700 (N_4700,N_3631,N_3735);
nor U4701 (N_4701,N_3082,N_3538);
and U4702 (N_4702,N_3771,N_3694);
or U4703 (N_4703,N_3728,N_3272);
and U4704 (N_4704,N_3270,N_3148);
nand U4705 (N_4705,N_3319,N_3677);
or U4706 (N_4706,N_3838,N_3247);
and U4707 (N_4707,N_3396,N_3553);
or U4708 (N_4708,N_3791,N_3268);
nand U4709 (N_4709,N_3054,N_3711);
nor U4710 (N_4710,N_3687,N_3911);
nor U4711 (N_4711,N_3365,N_3595);
nor U4712 (N_4712,N_3944,N_3632);
nor U4713 (N_4713,N_3151,N_3771);
nor U4714 (N_4714,N_3495,N_3378);
nor U4715 (N_4715,N_3056,N_3785);
and U4716 (N_4716,N_3945,N_3440);
nor U4717 (N_4717,N_3809,N_3451);
nor U4718 (N_4718,N_3618,N_3529);
or U4719 (N_4719,N_3923,N_3711);
xnor U4720 (N_4720,N_3919,N_3595);
and U4721 (N_4721,N_3595,N_3035);
nand U4722 (N_4722,N_3248,N_3306);
xnor U4723 (N_4723,N_3921,N_3335);
nor U4724 (N_4724,N_3022,N_3199);
or U4725 (N_4725,N_3817,N_3984);
and U4726 (N_4726,N_3235,N_3695);
nand U4727 (N_4727,N_3610,N_3783);
nor U4728 (N_4728,N_3681,N_3196);
xor U4729 (N_4729,N_3199,N_3519);
nand U4730 (N_4730,N_3921,N_3030);
nand U4731 (N_4731,N_3985,N_3952);
or U4732 (N_4732,N_3107,N_3468);
or U4733 (N_4733,N_3283,N_3852);
nand U4734 (N_4734,N_3855,N_3976);
and U4735 (N_4735,N_3296,N_3284);
nor U4736 (N_4736,N_3524,N_3060);
xor U4737 (N_4737,N_3440,N_3151);
and U4738 (N_4738,N_3392,N_3408);
nand U4739 (N_4739,N_3137,N_3208);
or U4740 (N_4740,N_3408,N_3488);
nor U4741 (N_4741,N_3656,N_3536);
and U4742 (N_4742,N_3007,N_3425);
nor U4743 (N_4743,N_3518,N_3883);
nand U4744 (N_4744,N_3034,N_3452);
or U4745 (N_4745,N_3055,N_3238);
or U4746 (N_4746,N_3791,N_3227);
and U4747 (N_4747,N_3870,N_3008);
nor U4748 (N_4748,N_3319,N_3820);
nand U4749 (N_4749,N_3839,N_3825);
nand U4750 (N_4750,N_3341,N_3232);
nor U4751 (N_4751,N_3560,N_3646);
or U4752 (N_4752,N_3249,N_3631);
nor U4753 (N_4753,N_3261,N_3024);
nand U4754 (N_4754,N_3886,N_3516);
and U4755 (N_4755,N_3260,N_3562);
or U4756 (N_4756,N_3432,N_3092);
and U4757 (N_4757,N_3109,N_3712);
nand U4758 (N_4758,N_3553,N_3737);
nor U4759 (N_4759,N_3289,N_3203);
and U4760 (N_4760,N_3781,N_3800);
xor U4761 (N_4761,N_3735,N_3662);
and U4762 (N_4762,N_3040,N_3073);
nand U4763 (N_4763,N_3944,N_3356);
or U4764 (N_4764,N_3737,N_3950);
nand U4765 (N_4765,N_3681,N_3144);
nand U4766 (N_4766,N_3974,N_3531);
nor U4767 (N_4767,N_3221,N_3832);
nor U4768 (N_4768,N_3744,N_3769);
or U4769 (N_4769,N_3272,N_3111);
nand U4770 (N_4770,N_3200,N_3007);
and U4771 (N_4771,N_3668,N_3497);
nand U4772 (N_4772,N_3876,N_3246);
and U4773 (N_4773,N_3347,N_3544);
nor U4774 (N_4774,N_3490,N_3225);
or U4775 (N_4775,N_3446,N_3643);
nor U4776 (N_4776,N_3780,N_3623);
and U4777 (N_4777,N_3545,N_3180);
nand U4778 (N_4778,N_3088,N_3972);
and U4779 (N_4779,N_3051,N_3461);
and U4780 (N_4780,N_3218,N_3673);
nand U4781 (N_4781,N_3340,N_3422);
xnor U4782 (N_4782,N_3490,N_3906);
nand U4783 (N_4783,N_3595,N_3607);
nand U4784 (N_4784,N_3708,N_3149);
xor U4785 (N_4785,N_3315,N_3932);
or U4786 (N_4786,N_3067,N_3213);
nor U4787 (N_4787,N_3062,N_3109);
or U4788 (N_4788,N_3784,N_3847);
xnor U4789 (N_4789,N_3222,N_3575);
nand U4790 (N_4790,N_3858,N_3061);
xor U4791 (N_4791,N_3249,N_3395);
nand U4792 (N_4792,N_3147,N_3305);
nor U4793 (N_4793,N_3713,N_3964);
and U4794 (N_4794,N_3345,N_3408);
nand U4795 (N_4795,N_3346,N_3239);
nand U4796 (N_4796,N_3265,N_3933);
and U4797 (N_4797,N_3377,N_3841);
nand U4798 (N_4798,N_3886,N_3027);
nor U4799 (N_4799,N_3839,N_3402);
and U4800 (N_4800,N_3079,N_3178);
nand U4801 (N_4801,N_3748,N_3281);
and U4802 (N_4802,N_3347,N_3091);
and U4803 (N_4803,N_3606,N_3904);
nand U4804 (N_4804,N_3507,N_3756);
or U4805 (N_4805,N_3214,N_3206);
or U4806 (N_4806,N_3179,N_3599);
nand U4807 (N_4807,N_3592,N_3265);
and U4808 (N_4808,N_3732,N_3606);
nor U4809 (N_4809,N_3697,N_3892);
and U4810 (N_4810,N_3909,N_3527);
nor U4811 (N_4811,N_3657,N_3253);
and U4812 (N_4812,N_3841,N_3941);
nor U4813 (N_4813,N_3575,N_3249);
nor U4814 (N_4814,N_3139,N_3482);
nor U4815 (N_4815,N_3517,N_3519);
xnor U4816 (N_4816,N_3364,N_3297);
or U4817 (N_4817,N_3681,N_3250);
nand U4818 (N_4818,N_3168,N_3905);
or U4819 (N_4819,N_3115,N_3776);
nand U4820 (N_4820,N_3855,N_3077);
nor U4821 (N_4821,N_3001,N_3206);
or U4822 (N_4822,N_3667,N_3176);
or U4823 (N_4823,N_3410,N_3177);
nand U4824 (N_4824,N_3560,N_3758);
nand U4825 (N_4825,N_3629,N_3121);
nor U4826 (N_4826,N_3133,N_3992);
and U4827 (N_4827,N_3374,N_3728);
and U4828 (N_4828,N_3757,N_3781);
nor U4829 (N_4829,N_3115,N_3481);
nand U4830 (N_4830,N_3626,N_3492);
nor U4831 (N_4831,N_3503,N_3593);
or U4832 (N_4832,N_3388,N_3416);
nand U4833 (N_4833,N_3637,N_3737);
nor U4834 (N_4834,N_3268,N_3618);
or U4835 (N_4835,N_3736,N_3830);
nand U4836 (N_4836,N_3467,N_3843);
or U4837 (N_4837,N_3509,N_3687);
and U4838 (N_4838,N_3173,N_3728);
nand U4839 (N_4839,N_3727,N_3986);
or U4840 (N_4840,N_3304,N_3928);
nor U4841 (N_4841,N_3314,N_3996);
nor U4842 (N_4842,N_3988,N_3235);
xor U4843 (N_4843,N_3356,N_3537);
nand U4844 (N_4844,N_3756,N_3853);
nand U4845 (N_4845,N_3356,N_3706);
nor U4846 (N_4846,N_3468,N_3087);
nor U4847 (N_4847,N_3271,N_3399);
nand U4848 (N_4848,N_3899,N_3360);
nand U4849 (N_4849,N_3915,N_3091);
nand U4850 (N_4850,N_3715,N_3831);
nor U4851 (N_4851,N_3636,N_3160);
nand U4852 (N_4852,N_3119,N_3051);
and U4853 (N_4853,N_3493,N_3979);
nor U4854 (N_4854,N_3119,N_3486);
nand U4855 (N_4855,N_3559,N_3924);
nor U4856 (N_4856,N_3675,N_3949);
and U4857 (N_4857,N_3798,N_3207);
nand U4858 (N_4858,N_3292,N_3989);
nor U4859 (N_4859,N_3120,N_3236);
nor U4860 (N_4860,N_3660,N_3605);
and U4861 (N_4861,N_3420,N_3559);
nand U4862 (N_4862,N_3328,N_3685);
or U4863 (N_4863,N_3296,N_3339);
and U4864 (N_4864,N_3937,N_3829);
nand U4865 (N_4865,N_3359,N_3749);
nor U4866 (N_4866,N_3865,N_3540);
nor U4867 (N_4867,N_3808,N_3506);
and U4868 (N_4868,N_3522,N_3169);
and U4869 (N_4869,N_3212,N_3778);
and U4870 (N_4870,N_3206,N_3059);
nor U4871 (N_4871,N_3456,N_3315);
or U4872 (N_4872,N_3674,N_3193);
nor U4873 (N_4873,N_3849,N_3796);
or U4874 (N_4874,N_3790,N_3674);
or U4875 (N_4875,N_3173,N_3267);
and U4876 (N_4876,N_3360,N_3487);
nor U4877 (N_4877,N_3335,N_3757);
nand U4878 (N_4878,N_3724,N_3561);
and U4879 (N_4879,N_3309,N_3527);
nand U4880 (N_4880,N_3278,N_3934);
nand U4881 (N_4881,N_3931,N_3583);
nor U4882 (N_4882,N_3649,N_3557);
nand U4883 (N_4883,N_3392,N_3311);
nor U4884 (N_4884,N_3786,N_3665);
and U4885 (N_4885,N_3738,N_3597);
nand U4886 (N_4886,N_3399,N_3792);
and U4887 (N_4887,N_3132,N_3128);
and U4888 (N_4888,N_3728,N_3133);
and U4889 (N_4889,N_3095,N_3510);
and U4890 (N_4890,N_3631,N_3155);
nor U4891 (N_4891,N_3992,N_3092);
and U4892 (N_4892,N_3688,N_3615);
nor U4893 (N_4893,N_3029,N_3137);
xnor U4894 (N_4894,N_3945,N_3566);
nand U4895 (N_4895,N_3733,N_3866);
or U4896 (N_4896,N_3411,N_3451);
nand U4897 (N_4897,N_3365,N_3908);
or U4898 (N_4898,N_3631,N_3808);
nand U4899 (N_4899,N_3030,N_3302);
nand U4900 (N_4900,N_3906,N_3917);
and U4901 (N_4901,N_3786,N_3224);
or U4902 (N_4902,N_3964,N_3505);
nor U4903 (N_4903,N_3815,N_3383);
nor U4904 (N_4904,N_3467,N_3566);
nand U4905 (N_4905,N_3769,N_3447);
nor U4906 (N_4906,N_3284,N_3134);
or U4907 (N_4907,N_3866,N_3629);
and U4908 (N_4908,N_3032,N_3668);
nor U4909 (N_4909,N_3628,N_3209);
or U4910 (N_4910,N_3120,N_3504);
or U4911 (N_4911,N_3642,N_3614);
nand U4912 (N_4912,N_3264,N_3687);
nor U4913 (N_4913,N_3227,N_3411);
or U4914 (N_4914,N_3248,N_3857);
or U4915 (N_4915,N_3463,N_3583);
and U4916 (N_4916,N_3800,N_3288);
nand U4917 (N_4917,N_3190,N_3300);
nor U4918 (N_4918,N_3151,N_3377);
xnor U4919 (N_4919,N_3505,N_3704);
or U4920 (N_4920,N_3074,N_3896);
and U4921 (N_4921,N_3553,N_3491);
xor U4922 (N_4922,N_3523,N_3456);
and U4923 (N_4923,N_3204,N_3260);
nand U4924 (N_4924,N_3055,N_3024);
nor U4925 (N_4925,N_3467,N_3803);
nand U4926 (N_4926,N_3487,N_3735);
xnor U4927 (N_4927,N_3353,N_3053);
nand U4928 (N_4928,N_3179,N_3367);
nand U4929 (N_4929,N_3095,N_3847);
and U4930 (N_4930,N_3617,N_3879);
nand U4931 (N_4931,N_3228,N_3339);
nor U4932 (N_4932,N_3401,N_3719);
or U4933 (N_4933,N_3621,N_3830);
nor U4934 (N_4934,N_3659,N_3708);
nor U4935 (N_4935,N_3560,N_3574);
nand U4936 (N_4936,N_3212,N_3187);
and U4937 (N_4937,N_3319,N_3292);
nand U4938 (N_4938,N_3644,N_3224);
nor U4939 (N_4939,N_3400,N_3571);
or U4940 (N_4940,N_3060,N_3219);
or U4941 (N_4941,N_3623,N_3871);
or U4942 (N_4942,N_3457,N_3794);
nor U4943 (N_4943,N_3168,N_3329);
xnor U4944 (N_4944,N_3579,N_3200);
nor U4945 (N_4945,N_3621,N_3739);
nand U4946 (N_4946,N_3180,N_3321);
nor U4947 (N_4947,N_3826,N_3504);
nand U4948 (N_4948,N_3898,N_3422);
or U4949 (N_4949,N_3238,N_3784);
nand U4950 (N_4950,N_3476,N_3638);
and U4951 (N_4951,N_3906,N_3255);
xnor U4952 (N_4952,N_3453,N_3838);
or U4953 (N_4953,N_3541,N_3512);
and U4954 (N_4954,N_3874,N_3039);
or U4955 (N_4955,N_3597,N_3096);
nand U4956 (N_4956,N_3088,N_3100);
and U4957 (N_4957,N_3157,N_3489);
nand U4958 (N_4958,N_3960,N_3308);
or U4959 (N_4959,N_3124,N_3976);
and U4960 (N_4960,N_3311,N_3530);
nand U4961 (N_4961,N_3220,N_3656);
nand U4962 (N_4962,N_3035,N_3112);
nand U4963 (N_4963,N_3477,N_3835);
or U4964 (N_4964,N_3402,N_3715);
xor U4965 (N_4965,N_3611,N_3641);
nand U4966 (N_4966,N_3181,N_3815);
or U4967 (N_4967,N_3972,N_3905);
or U4968 (N_4968,N_3930,N_3975);
nor U4969 (N_4969,N_3776,N_3533);
and U4970 (N_4970,N_3703,N_3159);
nand U4971 (N_4971,N_3962,N_3688);
nand U4972 (N_4972,N_3394,N_3927);
or U4973 (N_4973,N_3172,N_3224);
and U4974 (N_4974,N_3165,N_3485);
nand U4975 (N_4975,N_3090,N_3562);
or U4976 (N_4976,N_3665,N_3911);
nand U4977 (N_4977,N_3740,N_3260);
and U4978 (N_4978,N_3117,N_3896);
nor U4979 (N_4979,N_3304,N_3276);
nand U4980 (N_4980,N_3145,N_3128);
or U4981 (N_4981,N_3848,N_3945);
nor U4982 (N_4982,N_3224,N_3902);
xor U4983 (N_4983,N_3221,N_3100);
nand U4984 (N_4984,N_3187,N_3664);
xor U4985 (N_4985,N_3309,N_3506);
or U4986 (N_4986,N_3663,N_3057);
or U4987 (N_4987,N_3698,N_3519);
or U4988 (N_4988,N_3046,N_3567);
or U4989 (N_4989,N_3737,N_3308);
nand U4990 (N_4990,N_3072,N_3906);
nand U4991 (N_4991,N_3779,N_3950);
or U4992 (N_4992,N_3562,N_3902);
and U4993 (N_4993,N_3019,N_3282);
and U4994 (N_4994,N_3291,N_3356);
or U4995 (N_4995,N_3713,N_3196);
or U4996 (N_4996,N_3352,N_3922);
xor U4997 (N_4997,N_3111,N_3825);
or U4998 (N_4998,N_3661,N_3828);
and U4999 (N_4999,N_3865,N_3124);
or U5000 (N_5000,N_4011,N_4192);
or U5001 (N_5001,N_4881,N_4986);
nand U5002 (N_5002,N_4898,N_4727);
nand U5003 (N_5003,N_4020,N_4263);
and U5004 (N_5004,N_4870,N_4350);
nor U5005 (N_5005,N_4184,N_4850);
and U5006 (N_5006,N_4536,N_4674);
or U5007 (N_5007,N_4864,N_4512);
nor U5008 (N_5008,N_4501,N_4089);
and U5009 (N_5009,N_4498,N_4387);
nor U5010 (N_5010,N_4960,N_4289);
nor U5011 (N_5011,N_4481,N_4801);
and U5012 (N_5012,N_4516,N_4343);
nor U5013 (N_5013,N_4310,N_4836);
and U5014 (N_5014,N_4629,N_4706);
nor U5015 (N_5015,N_4726,N_4084);
and U5016 (N_5016,N_4781,N_4635);
or U5017 (N_5017,N_4433,N_4002);
nand U5018 (N_5018,N_4332,N_4539);
nor U5019 (N_5019,N_4693,N_4487);
or U5020 (N_5020,N_4579,N_4718);
and U5021 (N_5021,N_4054,N_4141);
or U5022 (N_5022,N_4630,N_4111);
or U5023 (N_5023,N_4030,N_4157);
nand U5024 (N_5024,N_4071,N_4307);
and U5025 (N_5025,N_4440,N_4928);
nor U5026 (N_5026,N_4599,N_4722);
nor U5027 (N_5027,N_4747,N_4117);
and U5028 (N_5028,N_4919,N_4892);
nand U5029 (N_5029,N_4428,N_4740);
or U5030 (N_5030,N_4255,N_4240);
and U5031 (N_5031,N_4026,N_4772);
or U5032 (N_5032,N_4499,N_4340);
nand U5033 (N_5033,N_4195,N_4637);
nor U5034 (N_5034,N_4092,N_4225);
or U5035 (N_5035,N_4865,N_4839);
nor U5036 (N_5036,N_4979,N_4602);
nor U5037 (N_5037,N_4473,N_4384);
or U5038 (N_5038,N_4010,N_4641);
nand U5039 (N_5039,N_4562,N_4634);
or U5040 (N_5040,N_4330,N_4743);
or U5041 (N_5041,N_4181,N_4770);
nor U5042 (N_5042,N_4404,N_4708);
nand U5043 (N_5043,N_4155,N_4085);
and U5044 (N_5044,N_4873,N_4578);
and U5045 (N_5045,N_4577,N_4122);
and U5046 (N_5046,N_4866,N_4761);
nand U5047 (N_5047,N_4994,N_4265);
and U5048 (N_5048,N_4282,N_4006);
xnor U5049 (N_5049,N_4720,N_4052);
xor U5050 (N_5050,N_4197,N_4570);
nor U5051 (N_5051,N_4165,N_4750);
or U5052 (N_5052,N_4259,N_4206);
and U5053 (N_5053,N_4547,N_4738);
or U5054 (N_5054,N_4956,N_4057);
and U5055 (N_5055,N_4502,N_4521);
nor U5056 (N_5056,N_4477,N_4749);
nand U5057 (N_5057,N_4863,N_4083);
nor U5058 (N_5058,N_4619,N_4372);
and U5059 (N_5059,N_4902,N_4403);
or U5060 (N_5060,N_4786,N_4779);
nand U5061 (N_5061,N_4078,N_4453);
nor U5062 (N_5062,N_4860,N_4788);
xor U5063 (N_5063,N_4491,N_4804);
or U5064 (N_5064,N_4542,N_4731);
or U5065 (N_5065,N_4716,N_4508);
or U5066 (N_5066,N_4912,N_4303);
nand U5067 (N_5067,N_4436,N_4245);
and U5068 (N_5068,N_4742,N_4612);
and U5069 (N_5069,N_4696,N_4368);
or U5070 (N_5070,N_4402,N_4909);
and U5071 (N_5071,N_4435,N_4035);
nand U5072 (N_5072,N_4686,N_4322);
nand U5073 (N_5073,N_4479,N_4586);
nor U5074 (N_5074,N_4583,N_4555);
or U5075 (N_5075,N_4982,N_4766);
and U5076 (N_5076,N_4201,N_4519);
nand U5077 (N_5077,N_4047,N_4906);
or U5078 (N_5078,N_4998,N_4464);
or U5079 (N_5079,N_4831,N_4894);
or U5080 (N_5080,N_4358,N_4389);
or U5081 (N_5081,N_4013,N_4224);
nor U5082 (N_5082,N_4449,N_4018);
nor U5083 (N_5083,N_4137,N_4971);
and U5084 (N_5084,N_4534,N_4463);
or U5085 (N_5085,N_4659,N_4689);
nor U5086 (N_5086,N_4613,N_4700);
xnor U5087 (N_5087,N_4895,N_4807);
and U5088 (N_5088,N_4569,N_4532);
and U5089 (N_5089,N_4136,N_4896);
nor U5090 (N_5090,N_4441,N_4952);
nand U5091 (N_5091,N_4407,N_4151);
and U5092 (N_5092,N_4735,N_4269);
nand U5093 (N_5093,N_4628,N_4390);
xor U5094 (N_5094,N_4995,N_4120);
and U5095 (N_5095,N_4210,N_4905);
nand U5096 (N_5096,N_4848,N_4765);
nor U5097 (N_5097,N_4760,N_4872);
and U5098 (N_5098,N_4036,N_4106);
nand U5099 (N_5099,N_4150,N_4654);
and U5100 (N_5100,N_4987,N_4661);
or U5101 (N_5101,N_4060,N_4230);
and U5102 (N_5102,N_4710,N_4672);
nor U5103 (N_5103,N_4764,N_4203);
xor U5104 (N_5104,N_4143,N_4156);
and U5105 (N_5105,N_4645,N_4056);
xor U5106 (N_5106,N_4335,N_4194);
or U5107 (N_5107,N_4783,N_4129);
and U5108 (N_5108,N_4300,N_4997);
or U5109 (N_5109,N_4219,N_4044);
nor U5110 (N_5110,N_4623,N_4116);
nand U5111 (N_5111,N_4782,N_4746);
or U5112 (N_5112,N_4684,N_4878);
and U5113 (N_5113,N_4585,N_4851);
and U5114 (N_5114,N_4533,N_4290);
or U5115 (N_5115,N_4298,N_4955);
and U5116 (N_5116,N_4703,N_4546);
or U5117 (N_5117,N_4027,N_4879);
nand U5118 (N_5118,N_4355,N_4093);
and U5119 (N_5119,N_4171,N_4843);
or U5120 (N_5120,N_4345,N_4077);
or U5121 (N_5121,N_4317,N_4600);
or U5122 (N_5122,N_4875,N_4581);
or U5123 (N_5123,N_4490,N_4597);
nand U5124 (N_5124,N_4816,N_4888);
and U5125 (N_5125,N_4837,N_4560);
and U5126 (N_5126,N_4552,N_4275);
xnor U5127 (N_5127,N_4636,N_4520);
and U5128 (N_5128,N_4469,N_4958);
nor U5129 (N_5129,N_4386,N_4103);
and U5130 (N_5130,N_4899,N_4671);
nor U5131 (N_5131,N_4347,N_4304);
and U5132 (N_5132,N_4177,N_4741);
nor U5133 (N_5133,N_4426,N_4271);
nor U5134 (N_5134,N_4395,N_4468);
nor U5135 (N_5135,N_4796,N_4144);
nand U5136 (N_5136,N_4179,N_4063);
or U5137 (N_5137,N_4311,N_4214);
and U5138 (N_5138,N_4438,N_4256);
or U5139 (N_5139,N_4734,N_4705);
nor U5140 (N_5140,N_4187,N_4154);
or U5141 (N_5141,N_4405,N_4470);
xnor U5142 (N_5142,N_4467,N_4970);
and U5143 (N_5143,N_4251,N_4076);
or U5144 (N_5144,N_4889,N_4457);
or U5145 (N_5145,N_4797,N_4833);
nor U5146 (N_5146,N_4711,N_4417);
nand U5147 (N_5147,N_4363,N_4416);
nand U5148 (N_5148,N_4717,N_4545);
nor U5149 (N_5149,N_4697,N_4528);
or U5150 (N_5150,N_4244,N_4461);
nand U5151 (N_5151,N_4495,N_4131);
nor U5152 (N_5152,N_4795,N_4305);
nor U5153 (N_5153,N_4945,N_4608);
or U5154 (N_5154,N_4531,N_4236);
nor U5155 (N_5155,N_4411,N_4066);
nand U5156 (N_5156,N_4062,N_4663);
nor U5157 (N_5157,N_4984,N_4789);
xor U5158 (N_5158,N_4721,N_4125);
nand U5159 (N_5159,N_4991,N_4687);
or U5160 (N_5160,N_4406,N_4302);
nor U5161 (N_5161,N_4321,N_4961);
nand U5162 (N_5162,N_4949,N_4965);
and U5163 (N_5163,N_4174,N_4603);
or U5164 (N_5164,N_4168,N_4723);
or U5165 (N_5165,N_4517,N_4660);
or U5166 (N_5166,N_4664,N_4124);
or U5167 (N_5167,N_4415,N_4065);
nand U5168 (N_5168,N_4218,N_4840);
nor U5169 (N_5169,N_4105,N_4568);
or U5170 (N_5170,N_4480,N_4421);
and U5171 (N_5171,N_4922,N_4972);
nand U5172 (N_5172,N_4513,N_4252);
or U5173 (N_5173,N_4088,N_4525);
nand U5174 (N_5174,N_4080,N_4079);
nor U5175 (N_5175,N_4353,N_4178);
and U5176 (N_5176,N_4200,N_4262);
and U5177 (N_5177,N_4459,N_4698);
or U5178 (N_5178,N_4454,N_4338);
xor U5179 (N_5179,N_4408,N_4934);
and U5180 (N_5180,N_4932,N_4937);
nand U5181 (N_5181,N_4926,N_4294);
nor U5182 (N_5182,N_4704,N_4605);
and U5183 (N_5183,N_4769,N_4334);
and U5184 (N_5184,N_4130,N_4073);
xor U5185 (N_5185,N_4028,N_4299);
nand U5186 (N_5186,N_4170,N_4064);
nand U5187 (N_5187,N_4683,N_4427);
or U5188 (N_5188,N_4025,N_4553);
nand U5189 (N_5189,N_4382,N_4486);
nor U5190 (N_5190,N_4694,N_4448);
nor U5191 (N_5191,N_4884,N_4900);
or U5192 (N_5192,N_4148,N_4633);
or U5193 (N_5193,N_4974,N_4903);
or U5194 (N_5194,N_4524,N_4337);
or U5195 (N_5195,N_4444,N_4847);
or U5196 (N_5196,N_4814,N_4400);
or U5197 (N_5197,N_4145,N_4152);
nand U5198 (N_5198,N_4183,N_4114);
nor U5199 (N_5199,N_4515,N_4316);
nor U5200 (N_5200,N_4050,N_4069);
nand U5201 (N_5201,N_4915,N_4792);
xor U5202 (N_5202,N_4754,N_4466);
nand U5203 (N_5203,N_4943,N_4679);
and U5204 (N_5204,N_4587,N_4166);
nor U5205 (N_5205,N_4544,N_4068);
and U5206 (N_5206,N_4649,N_4655);
or U5207 (N_5207,N_4996,N_4451);
and U5208 (N_5208,N_4622,N_4159);
and U5209 (N_5209,N_4993,N_4591);
and U5210 (N_5210,N_4045,N_4284);
and U5211 (N_5211,N_4505,N_4673);
or U5212 (N_5212,N_4431,N_4090);
and U5213 (N_5213,N_4383,N_4015);
and U5214 (N_5214,N_4901,N_4005);
nand U5215 (N_5215,N_4360,N_4859);
and U5216 (N_5216,N_4162,N_4046);
xor U5217 (N_5217,N_4618,N_4685);
and U5218 (N_5218,N_4173,N_4930);
nand U5219 (N_5219,N_4980,N_4295);
nand U5220 (N_5220,N_4670,N_4112);
and U5221 (N_5221,N_4308,N_4222);
or U5222 (N_5222,N_4753,N_4456);
nand U5223 (N_5223,N_4589,N_4551);
nand U5224 (N_5224,N_4108,N_4042);
nor U5225 (N_5225,N_4647,N_4333);
or U5226 (N_5226,N_4209,N_4110);
xnor U5227 (N_5227,N_4215,N_4667);
nor U5228 (N_5228,N_4627,N_4917);
xnor U5229 (N_5229,N_4399,N_4817);
nor U5230 (N_5230,N_4810,N_4235);
nor U5231 (N_5231,N_4351,N_4526);
and U5232 (N_5232,N_4541,N_4575);
nand U5233 (N_5233,N_4580,N_4959);
and U5234 (N_5234,N_4558,N_4756);
and U5235 (N_5235,N_4656,N_4730);
nor U5236 (N_5236,N_4616,N_4055);
nand U5237 (N_5237,N_4999,N_4274);
or U5238 (N_5238,N_4095,N_4429);
or U5239 (N_5239,N_4008,N_4410);
nor U5240 (N_5240,N_4356,N_4852);
or U5241 (N_5241,N_4301,N_4361);
nand U5242 (N_5242,N_4794,N_4279);
nor U5243 (N_5243,N_4554,N_4931);
and U5244 (N_5244,N_4500,N_4669);
nand U5245 (N_5245,N_4614,N_4253);
and U5246 (N_5246,N_4666,N_4824);
and U5247 (N_5247,N_4283,N_4983);
nor U5248 (N_5248,N_4014,N_4072);
nor U5249 (N_5249,N_4232,N_4439);
nand U5250 (N_5250,N_4733,N_4682);
or U5251 (N_5251,N_4530,N_4450);
nor U5252 (N_5252,N_4344,N_4856);
and U5253 (N_5253,N_4818,N_4196);
and U5254 (N_5254,N_4887,N_4370);
nor U5255 (N_5255,N_4348,N_4815);
or U5256 (N_5256,N_4913,N_4313);
or U5257 (N_5257,N_4947,N_4728);
or U5258 (N_5258,N_4808,N_4571);
nor U5259 (N_5259,N_4594,N_4364);
nor U5260 (N_5260,N_4771,N_4950);
xnor U5261 (N_5261,N_4180,N_4805);
or U5262 (N_5262,N_4186,N_4610);
or U5263 (N_5263,N_4153,N_4037);
nor U5264 (N_5264,N_4445,N_4973);
nor U5265 (N_5265,N_4869,N_4662);
nor U5266 (N_5266,N_4237,N_4584);
nand U5267 (N_5267,N_4446,N_4396);
nand U5268 (N_5268,N_4657,N_4273);
or U5269 (N_5269,N_4841,N_4161);
or U5270 (N_5270,N_4424,N_4329);
nand U5271 (N_5271,N_4167,N_4548);
nand U5272 (N_5272,N_4043,N_4202);
or U5273 (N_5273,N_4853,N_4504);
xnor U5274 (N_5274,N_4988,N_4285);
nor U5275 (N_5275,N_4927,N_4458);
or U5276 (N_5276,N_4871,N_4744);
or U5277 (N_5277,N_4009,N_4094);
and U5278 (N_5278,N_4207,N_4632);
and U5279 (N_5279,N_4455,N_4774);
xor U5280 (N_5280,N_4688,N_4990);
and U5281 (N_5281,N_4297,N_4572);
nor U5282 (N_5282,N_4425,N_4211);
and U5283 (N_5283,N_4739,N_4217);
nand U5284 (N_5284,N_4529,N_4509);
nor U5285 (N_5285,N_4346,N_4208);
nor U5286 (N_5286,N_4714,N_4326);
and U5287 (N_5287,N_4376,N_4462);
or U5288 (N_5288,N_4296,N_4392);
nor U5289 (N_5289,N_4590,N_4118);
and U5290 (N_5290,N_4827,N_4198);
or U5291 (N_5291,N_4022,N_4910);
and U5292 (N_5292,N_4737,N_4767);
and U5293 (N_5293,N_4437,N_4857);
or U5294 (N_5294,N_4147,N_4024);
xor U5295 (N_5295,N_4061,N_4938);
and U5296 (N_5296,N_4272,N_4642);
nand U5297 (N_5297,N_4725,N_4388);
nor U5298 (N_5298,N_4104,N_4327);
or U5299 (N_5299,N_4081,N_4366);
nor U5300 (N_5300,N_4842,N_4434);
nor U5301 (N_5301,N_4966,N_4646);
nor U5302 (N_5302,N_4699,N_4748);
nand U5303 (N_5303,N_4371,N_4012);
nand U5304 (N_5304,N_4191,N_4653);
xnor U5305 (N_5305,N_4963,N_4397);
nor U5306 (N_5306,N_4595,N_4331);
and U5307 (N_5307,N_4835,N_4258);
nand U5308 (N_5308,N_4709,N_4452);
and U5309 (N_5309,N_4288,N_4625);
nand U5310 (N_5310,N_4886,N_4212);
and U5311 (N_5311,N_4598,N_4806);
nand U5312 (N_5312,N_4086,N_4380);
nor U5313 (N_5313,N_4342,N_4527);
and U5314 (N_5314,N_4862,N_4163);
xor U5315 (N_5315,N_4430,N_4574);
nor U5316 (N_5316,N_4139,N_4820);
xnor U5317 (N_5317,N_4476,N_4119);
xor U5318 (N_5318,N_4375,N_4241);
nor U5319 (N_5319,N_4315,N_4828);
nor U5320 (N_5320,N_4049,N_4609);
or U5321 (N_5321,N_4695,N_4443);
nor U5322 (N_5322,N_4149,N_4442);
nor U5323 (N_5323,N_4229,N_4292);
nor U5324 (N_5324,N_4422,N_4854);
or U5325 (N_5325,N_4306,N_4017);
and U5326 (N_5326,N_4040,N_4496);
nand U5327 (N_5327,N_4099,N_4164);
and U5328 (N_5328,N_4755,N_4096);
nand U5329 (N_5329,N_4277,N_4732);
and U5330 (N_5330,N_4098,N_4626);
and U5331 (N_5331,N_4650,N_4893);
nand U5332 (N_5332,N_4234,N_4556);
nand U5333 (N_5333,N_4812,N_4838);
and U5334 (N_5334,N_4260,N_4328);
nand U5335 (N_5335,N_4447,N_4354);
nand U5336 (N_5336,N_4923,N_4377);
or U5337 (N_5337,N_4518,N_4822);
nand U5338 (N_5338,N_4675,N_4032);
xnor U5339 (N_5339,N_4140,N_4787);
nor U5340 (N_5340,N_4713,N_4751);
or U5341 (N_5341,N_4549,N_4257);
or U5342 (N_5342,N_4097,N_4051);
nand U5343 (N_5343,N_4221,N_4891);
or U5344 (N_5344,N_4715,N_4855);
nor U5345 (N_5345,N_4543,N_4778);
nor U5346 (N_5346,N_4921,N_4123);
nand U5347 (N_5347,N_4780,N_4784);
nand U5348 (N_5348,N_4320,N_4904);
nand U5349 (N_5349,N_4975,N_4540);
or U5350 (N_5350,N_4908,N_4877);
xnor U5351 (N_5351,N_4776,N_4185);
nor U5352 (N_5352,N_4176,N_4712);
and U5353 (N_5353,N_4385,N_4911);
and U5354 (N_5354,N_4977,N_4160);
nor U5355 (N_5355,N_4668,N_4373);
or U5356 (N_5356,N_4325,N_4621);
nor U5357 (N_5357,N_4882,N_4418);
and U5358 (N_5358,N_4398,N_4620);
or U5359 (N_5359,N_4825,N_4216);
xnor U5360 (N_5360,N_4369,N_4199);
nor U5361 (N_5361,N_4193,N_4341);
nand U5362 (N_5362,N_4034,N_4803);
nor U5363 (N_5363,N_4953,N_4261);
or U5364 (N_5364,N_4019,N_4918);
nor U5365 (N_5365,N_4511,N_4550);
nor U5366 (N_5366,N_4367,N_4362);
xnor U5367 (N_5367,N_4967,N_4231);
nand U5368 (N_5368,N_4278,N_4314);
and U5369 (N_5369,N_4482,N_4916);
xnor U5370 (N_5370,N_4107,N_4565);
nor U5371 (N_5371,N_4640,N_4601);
nand U5372 (N_5372,N_4175,N_4799);
nor U5373 (N_5373,N_4133,N_4409);
or U5374 (N_5374,N_4791,N_4226);
nor U5375 (N_5375,N_4115,N_4651);
nor U5376 (N_5376,N_4567,N_4826);
or U5377 (N_5377,N_4091,N_4954);
nor U5378 (N_5378,N_4243,N_4293);
or U5379 (N_5379,N_4576,N_4239);
nand U5380 (N_5380,N_4758,N_4537);
nor U5381 (N_5381,N_4678,N_4264);
nor U5382 (N_5382,N_4109,N_4414);
nor U5383 (N_5383,N_4978,N_4652);
and U5384 (N_5384,N_4522,N_4004);
nor U5385 (N_5385,N_4510,N_4844);
or U5386 (N_5386,N_4033,N_4793);
or U5387 (N_5387,N_4981,N_4082);
nand U5388 (N_5388,N_4102,N_4939);
and U5389 (N_5389,N_4053,N_4607);
nor U5390 (N_5390,N_4503,N_4920);
or U5391 (N_5391,N_4413,N_4359);
nor U5392 (N_5392,N_4132,N_4126);
nor U5393 (N_5393,N_4615,N_4867);
nand U5394 (N_5394,N_4336,N_4475);
or U5395 (N_5395,N_4763,N_4883);
nand U5396 (N_5396,N_4819,N_4190);
or U5397 (N_5397,N_4701,N_4204);
nor U5398 (N_5398,N_4003,N_4777);
or U5399 (N_5399,N_4489,N_4559);
and U5400 (N_5400,N_4058,N_4617);
nand U5401 (N_5401,N_4691,N_4485);
nor U5402 (N_5402,N_4420,N_4472);
nand U5403 (N_5403,N_4067,N_4573);
or U5404 (N_5404,N_4985,N_4432);
or U5405 (N_5405,N_4007,N_4287);
nand U5406 (N_5406,N_4205,N_4000);
nor U5407 (N_5407,N_4270,N_4412);
nor U5408 (N_5408,N_4323,N_4665);
nor U5409 (N_5409,N_4291,N_4557);
nand U5410 (N_5410,N_4266,N_4798);
nand U5411 (N_5411,N_4648,N_4757);
and U5412 (N_5412,N_4729,N_4381);
or U5413 (N_5413,N_4039,N_4514);
nand U5414 (N_5414,N_4592,N_4924);
nor U5415 (N_5415,N_4379,N_4561);
nor U5416 (N_5416,N_4134,N_4493);
nor U5417 (N_5417,N_4228,N_4929);
or U5418 (N_5418,N_4507,N_4658);
nor U5419 (N_5419,N_4624,N_4318);
nand U5420 (N_5420,N_4989,N_4074);
or U5421 (N_5421,N_4339,N_4100);
nand U5422 (N_5422,N_4811,N_4745);
or U5423 (N_5423,N_4566,N_4773);
or U5424 (N_5424,N_4478,N_4227);
and U5425 (N_5425,N_4849,N_4775);
and U5426 (N_5426,N_4638,N_4936);
nor U5427 (N_5427,N_4254,N_4135);
xnor U5428 (N_5428,N_4246,N_4823);
and U5429 (N_5429,N_4643,N_4604);
or U5430 (N_5430,N_4169,N_4942);
nand U5431 (N_5431,N_4564,N_4535);
and U5432 (N_5432,N_4897,N_4846);
or U5433 (N_5433,N_4752,N_4087);
and U5434 (N_5434,N_4031,N_4868);
and U5435 (N_5435,N_4680,N_4719);
or U5436 (N_5436,N_4702,N_4631);
nor U5437 (N_5437,N_4059,N_4834);
nand U5438 (N_5438,N_4250,N_4021);
nor U5439 (N_5439,N_4378,N_4127);
or U5440 (N_5440,N_4692,N_4121);
and U5441 (N_5441,N_4940,N_4038);
nand U5442 (N_5442,N_4484,N_4276);
nor U5443 (N_5443,N_4324,N_4312);
nand U5444 (N_5444,N_4223,N_4001);
and U5445 (N_5445,N_4474,N_4724);
xnor U5446 (N_5446,N_4785,N_4401);
xnor U5447 (N_5447,N_4933,N_4821);
nand U5448 (N_5448,N_4874,N_4041);
xnor U5449 (N_5449,N_4267,N_4914);
nor U5450 (N_5450,N_4596,N_4423);
xor U5451 (N_5451,N_4172,N_4220);
nand U5452 (N_5452,N_4248,N_4497);
xnor U5453 (N_5453,N_4182,N_4070);
or U5454 (N_5454,N_4677,N_4813);
xor U5455 (N_5455,N_4880,N_4858);
or U5456 (N_5456,N_4016,N_4349);
or U5457 (N_5457,N_4861,N_4365);
or U5458 (N_5458,N_4189,N_4465);
nand U5459 (N_5459,N_4113,N_4506);
nand U5460 (N_5460,N_4492,N_4023);
and U5461 (N_5461,N_4249,N_4969);
nor U5462 (N_5462,N_4941,N_4676);
nand U5463 (N_5463,N_4606,N_4736);
nor U5464 (N_5464,N_4048,N_4247);
nor U5465 (N_5465,N_4890,N_4962);
and U5466 (N_5466,N_4281,N_4563);
or U5467 (N_5467,N_4393,N_4391);
nand U5468 (N_5468,N_4588,N_4968);
nand U5469 (N_5469,N_4523,N_4582);
or U5470 (N_5470,N_4946,N_4876);
nand U5471 (N_5471,N_4829,N_4142);
xor U5472 (N_5472,N_4158,N_4944);
or U5473 (N_5473,N_4075,N_4809);
or U5474 (N_5474,N_4483,N_4494);
and U5475 (N_5475,N_4188,N_4925);
nor U5476 (N_5476,N_4885,N_4611);
nor U5477 (N_5477,N_4790,N_4976);
or U5478 (N_5478,N_4681,N_4029);
nand U5479 (N_5479,N_4957,N_4309);
nor U5480 (N_5480,N_4707,N_4460);
or U5481 (N_5481,N_4762,N_4280);
or U5482 (N_5482,N_4286,N_4845);
xor U5483 (N_5483,N_4768,N_4101);
nor U5484 (N_5484,N_4593,N_4538);
nand U5485 (N_5485,N_4233,N_4242);
and U5486 (N_5486,N_4951,N_4832);
and U5487 (N_5487,N_4357,N_4146);
nor U5488 (N_5488,N_4319,N_4907);
or U5489 (N_5489,N_4268,N_4639);
or U5490 (N_5490,N_4471,N_4948);
and U5491 (N_5491,N_4374,N_4800);
and U5492 (N_5492,N_4644,N_4138);
or U5493 (N_5493,N_4419,N_4759);
xor U5494 (N_5494,N_4488,N_4690);
nor U5495 (N_5495,N_4964,N_4802);
nor U5496 (N_5496,N_4992,N_4830);
nor U5497 (N_5497,N_4352,N_4238);
or U5498 (N_5498,N_4935,N_4128);
nand U5499 (N_5499,N_4394,N_4213);
nor U5500 (N_5500,N_4292,N_4662);
and U5501 (N_5501,N_4956,N_4071);
nand U5502 (N_5502,N_4610,N_4532);
xor U5503 (N_5503,N_4358,N_4143);
nand U5504 (N_5504,N_4243,N_4026);
nand U5505 (N_5505,N_4202,N_4643);
nand U5506 (N_5506,N_4737,N_4153);
and U5507 (N_5507,N_4618,N_4869);
or U5508 (N_5508,N_4680,N_4897);
nor U5509 (N_5509,N_4703,N_4146);
or U5510 (N_5510,N_4367,N_4677);
or U5511 (N_5511,N_4104,N_4850);
and U5512 (N_5512,N_4218,N_4134);
nor U5513 (N_5513,N_4888,N_4291);
and U5514 (N_5514,N_4834,N_4772);
or U5515 (N_5515,N_4719,N_4424);
and U5516 (N_5516,N_4434,N_4978);
or U5517 (N_5517,N_4956,N_4123);
or U5518 (N_5518,N_4394,N_4309);
and U5519 (N_5519,N_4305,N_4771);
and U5520 (N_5520,N_4305,N_4183);
or U5521 (N_5521,N_4199,N_4893);
nor U5522 (N_5522,N_4809,N_4022);
or U5523 (N_5523,N_4795,N_4828);
nor U5524 (N_5524,N_4797,N_4364);
xnor U5525 (N_5525,N_4684,N_4940);
or U5526 (N_5526,N_4513,N_4212);
or U5527 (N_5527,N_4142,N_4162);
and U5528 (N_5528,N_4505,N_4209);
nor U5529 (N_5529,N_4402,N_4498);
nor U5530 (N_5530,N_4961,N_4122);
or U5531 (N_5531,N_4388,N_4802);
and U5532 (N_5532,N_4942,N_4903);
or U5533 (N_5533,N_4992,N_4667);
and U5534 (N_5534,N_4736,N_4388);
or U5535 (N_5535,N_4630,N_4531);
nand U5536 (N_5536,N_4339,N_4760);
nor U5537 (N_5537,N_4130,N_4820);
nand U5538 (N_5538,N_4334,N_4672);
nor U5539 (N_5539,N_4954,N_4933);
nand U5540 (N_5540,N_4863,N_4994);
xnor U5541 (N_5541,N_4714,N_4459);
and U5542 (N_5542,N_4678,N_4055);
nor U5543 (N_5543,N_4441,N_4615);
nand U5544 (N_5544,N_4293,N_4069);
or U5545 (N_5545,N_4349,N_4323);
or U5546 (N_5546,N_4313,N_4856);
or U5547 (N_5547,N_4771,N_4979);
and U5548 (N_5548,N_4811,N_4796);
and U5549 (N_5549,N_4449,N_4007);
nor U5550 (N_5550,N_4472,N_4905);
nand U5551 (N_5551,N_4088,N_4567);
nand U5552 (N_5552,N_4577,N_4442);
nor U5553 (N_5553,N_4624,N_4605);
and U5554 (N_5554,N_4656,N_4407);
and U5555 (N_5555,N_4275,N_4943);
nor U5556 (N_5556,N_4125,N_4491);
nor U5557 (N_5557,N_4615,N_4328);
and U5558 (N_5558,N_4841,N_4317);
xnor U5559 (N_5559,N_4384,N_4374);
nand U5560 (N_5560,N_4276,N_4880);
or U5561 (N_5561,N_4784,N_4493);
nand U5562 (N_5562,N_4277,N_4924);
or U5563 (N_5563,N_4209,N_4367);
nor U5564 (N_5564,N_4026,N_4512);
and U5565 (N_5565,N_4892,N_4872);
nand U5566 (N_5566,N_4983,N_4835);
nand U5567 (N_5567,N_4745,N_4096);
or U5568 (N_5568,N_4441,N_4857);
nor U5569 (N_5569,N_4578,N_4075);
nor U5570 (N_5570,N_4241,N_4320);
nand U5571 (N_5571,N_4424,N_4278);
nor U5572 (N_5572,N_4130,N_4558);
nand U5573 (N_5573,N_4990,N_4137);
and U5574 (N_5574,N_4794,N_4899);
and U5575 (N_5575,N_4202,N_4549);
or U5576 (N_5576,N_4629,N_4582);
nor U5577 (N_5577,N_4959,N_4751);
or U5578 (N_5578,N_4647,N_4771);
xor U5579 (N_5579,N_4365,N_4759);
or U5580 (N_5580,N_4152,N_4009);
or U5581 (N_5581,N_4293,N_4736);
and U5582 (N_5582,N_4909,N_4606);
nor U5583 (N_5583,N_4099,N_4245);
or U5584 (N_5584,N_4680,N_4141);
or U5585 (N_5585,N_4838,N_4659);
and U5586 (N_5586,N_4003,N_4882);
and U5587 (N_5587,N_4532,N_4757);
nand U5588 (N_5588,N_4278,N_4426);
nand U5589 (N_5589,N_4956,N_4181);
nand U5590 (N_5590,N_4885,N_4684);
xor U5591 (N_5591,N_4566,N_4138);
or U5592 (N_5592,N_4240,N_4918);
nor U5593 (N_5593,N_4052,N_4862);
and U5594 (N_5594,N_4514,N_4723);
nand U5595 (N_5595,N_4845,N_4715);
and U5596 (N_5596,N_4997,N_4279);
and U5597 (N_5597,N_4066,N_4555);
nand U5598 (N_5598,N_4712,N_4557);
and U5599 (N_5599,N_4985,N_4063);
or U5600 (N_5600,N_4279,N_4349);
and U5601 (N_5601,N_4172,N_4411);
or U5602 (N_5602,N_4623,N_4774);
nand U5603 (N_5603,N_4849,N_4435);
and U5604 (N_5604,N_4319,N_4760);
nor U5605 (N_5605,N_4851,N_4934);
or U5606 (N_5606,N_4864,N_4853);
nand U5607 (N_5607,N_4544,N_4677);
nor U5608 (N_5608,N_4833,N_4300);
nor U5609 (N_5609,N_4831,N_4120);
or U5610 (N_5610,N_4093,N_4157);
nand U5611 (N_5611,N_4731,N_4726);
nor U5612 (N_5612,N_4164,N_4171);
nor U5613 (N_5613,N_4052,N_4378);
and U5614 (N_5614,N_4096,N_4452);
nor U5615 (N_5615,N_4956,N_4315);
or U5616 (N_5616,N_4527,N_4714);
and U5617 (N_5617,N_4808,N_4382);
xnor U5618 (N_5618,N_4491,N_4446);
or U5619 (N_5619,N_4403,N_4752);
nor U5620 (N_5620,N_4598,N_4422);
and U5621 (N_5621,N_4134,N_4405);
or U5622 (N_5622,N_4246,N_4764);
nor U5623 (N_5623,N_4014,N_4877);
nand U5624 (N_5624,N_4067,N_4047);
nor U5625 (N_5625,N_4814,N_4197);
and U5626 (N_5626,N_4195,N_4646);
nand U5627 (N_5627,N_4449,N_4059);
xor U5628 (N_5628,N_4138,N_4951);
and U5629 (N_5629,N_4089,N_4511);
or U5630 (N_5630,N_4479,N_4104);
or U5631 (N_5631,N_4255,N_4719);
xnor U5632 (N_5632,N_4916,N_4227);
and U5633 (N_5633,N_4338,N_4110);
xnor U5634 (N_5634,N_4251,N_4077);
nand U5635 (N_5635,N_4150,N_4448);
nand U5636 (N_5636,N_4401,N_4709);
xor U5637 (N_5637,N_4230,N_4108);
and U5638 (N_5638,N_4326,N_4402);
and U5639 (N_5639,N_4684,N_4994);
nand U5640 (N_5640,N_4215,N_4424);
and U5641 (N_5641,N_4952,N_4083);
nand U5642 (N_5642,N_4403,N_4255);
nand U5643 (N_5643,N_4523,N_4305);
xnor U5644 (N_5644,N_4393,N_4405);
nand U5645 (N_5645,N_4381,N_4290);
and U5646 (N_5646,N_4234,N_4757);
or U5647 (N_5647,N_4415,N_4420);
or U5648 (N_5648,N_4497,N_4757);
xnor U5649 (N_5649,N_4102,N_4335);
and U5650 (N_5650,N_4081,N_4567);
xor U5651 (N_5651,N_4316,N_4347);
and U5652 (N_5652,N_4254,N_4370);
and U5653 (N_5653,N_4818,N_4279);
and U5654 (N_5654,N_4648,N_4616);
and U5655 (N_5655,N_4902,N_4319);
nor U5656 (N_5656,N_4227,N_4131);
nor U5657 (N_5657,N_4444,N_4370);
nand U5658 (N_5658,N_4768,N_4911);
or U5659 (N_5659,N_4216,N_4569);
nand U5660 (N_5660,N_4556,N_4947);
and U5661 (N_5661,N_4374,N_4695);
or U5662 (N_5662,N_4669,N_4021);
nor U5663 (N_5663,N_4816,N_4299);
and U5664 (N_5664,N_4095,N_4599);
and U5665 (N_5665,N_4413,N_4577);
nor U5666 (N_5666,N_4199,N_4356);
nor U5667 (N_5667,N_4145,N_4066);
nand U5668 (N_5668,N_4277,N_4313);
nand U5669 (N_5669,N_4584,N_4947);
and U5670 (N_5670,N_4620,N_4833);
or U5671 (N_5671,N_4974,N_4584);
and U5672 (N_5672,N_4861,N_4402);
nor U5673 (N_5673,N_4236,N_4590);
nand U5674 (N_5674,N_4187,N_4944);
nand U5675 (N_5675,N_4916,N_4172);
nor U5676 (N_5676,N_4046,N_4411);
nor U5677 (N_5677,N_4955,N_4489);
nor U5678 (N_5678,N_4709,N_4257);
xor U5679 (N_5679,N_4510,N_4646);
nor U5680 (N_5680,N_4947,N_4161);
nand U5681 (N_5681,N_4020,N_4135);
or U5682 (N_5682,N_4021,N_4216);
nor U5683 (N_5683,N_4460,N_4124);
nor U5684 (N_5684,N_4174,N_4960);
nor U5685 (N_5685,N_4989,N_4189);
nor U5686 (N_5686,N_4770,N_4615);
or U5687 (N_5687,N_4756,N_4195);
nor U5688 (N_5688,N_4511,N_4514);
nand U5689 (N_5689,N_4562,N_4075);
nand U5690 (N_5690,N_4144,N_4700);
nor U5691 (N_5691,N_4291,N_4708);
and U5692 (N_5692,N_4695,N_4827);
nand U5693 (N_5693,N_4724,N_4855);
nor U5694 (N_5694,N_4450,N_4782);
nor U5695 (N_5695,N_4008,N_4535);
nand U5696 (N_5696,N_4310,N_4054);
nor U5697 (N_5697,N_4729,N_4831);
and U5698 (N_5698,N_4406,N_4135);
and U5699 (N_5699,N_4295,N_4092);
nand U5700 (N_5700,N_4136,N_4367);
and U5701 (N_5701,N_4325,N_4423);
nor U5702 (N_5702,N_4846,N_4717);
and U5703 (N_5703,N_4435,N_4257);
nor U5704 (N_5704,N_4356,N_4181);
or U5705 (N_5705,N_4607,N_4161);
and U5706 (N_5706,N_4255,N_4739);
or U5707 (N_5707,N_4928,N_4611);
nor U5708 (N_5708,N_4601,N_4492);
nor U5709 (N_5709,N_4978,N_4571);
nor U5710 (N_5710,N_4272,N_4247);
nand U5711 (N_5711,N_4061,N_4480);
nor U5712 (N_5712,N_4523,N_4830);
nor U5713 (N_5713,N_4995,N_4617);
nand U5714 (N_5714,N_4296,N_4408);
and U5715 (N_5715,N_4379,N_4088);
and U5716 (N_5716,N_4597,N_4376);
and U5717 (N_5717,N_4619,N_4564);
nand U5718 (N_5718,N_4495,N_4496);
and U5719 (N_5719,N_4897,N_4373);
or U5720 (N_5720,N_4996,N_4575);
and U5721 (N_5721,N_4525,N_4937);
nand U5722 (N_5722,N_4227,N_4475);
or U5723 (N_5723,N_4082,N_4218);
xor U5724 (N_5724,N_4727,N_4433);
and U5725 (N_5725,N_4470,N_4113);
nand U5726 (N_5726,N_4634,N_4986);
nor U5727 (N_5727,N_4077,N_4566);
nand U5728 (N_5728,N_4353,N_4528);
or U5729 (N_5729,N_4751,N_4012);
nand U5730 (N_5730,N_4459,N_4760);
and U5731 (N_5731,N_4320,N_4513);
nor U5732 (N_5732,N_4166,N_4100);
nand U5733 (N_5733,N_4508,N_4711);
and U5734 (N_5734,N_4070,N_4591);
nand U5735 (N_5735,N_4399,N_4059);
nor U5736 (N_5736,N_4754,N_4860);
nand U5737 (N_5737,N_4269,N_4903);
nor U5738 (N_5738,N_4643,N_4805);
xnor U5739 (N_5739,N_4205,N_4162);
nand U5740 (N_5740,N_4527,N_4362);
or U5741 (N_5741,N_4654,N_4053);
nor U5742 (N_5742,N_4461,N_4039);
or U5743 (N_5743,N_4341,N_4684);
or U5744 (N_5744,N_4825,N_4477);
nor U5745 (N_5745,N_4698,N_4603);
nor U5746 (N_5746,N_4123,N_4222);
and U5747 (N_5747,N_4147,N_4356);
nor U5748 (N_5748,N_4136,N_4670);
xor U5749 (N_5749,N_4543,N_4720);
nor U5750 (N_5750,N_4833,N_4329);
nor U5751 (N_5751,N_4399,N_4278);
or U5752 (N_5752,N_4807,N_4186);
nor U5753 (N_5753,N_4649,N_4824);
nand U5754 (N_5754,N_4712,N_4874);
xor U5755 (N_5755,N_4987,N_4424);
and U5756 (N_5756,N_4958,N_4386);
xor U5757 (N_5757,N_4430,N_4078);
or U5758 (N_5758,N_4230,N_4307);
nand U5759 (N_5759,N_4207,N_4129);
nor U5760 (N_5760,N_4116,N_4544);
nor U5761 (N_5761,N_4374,N_4757);
and U5762 (N_5762,N_4902,N_4960);
nand U5763 (N_5763,N_4886,N_4258);
or U5764 (N_5764,N_4832,N_4496);
and U5765 (N_5765,N_4717,N_4654);
nor U5766 (N_5766,N_4181,N_4863);
nor U5767 (N_5767,N_4585,N_4287);
xnor U5768 (N_5768,N_4421,N_4553);
nor U5769 (N_5769,N_4295,N_4126);
nand U5770 (N_5770,N_4892,N_4721);
xor U5771 (N_5771,N_4583,N_4778);
xnor U5772 (N_5772,N_4556,N_4682);
and U5773 (N_5773,N_4004,N_4354);
nor U5774 (N_5774,N_4444,N_4054);
xnor U5775 (N_5775,N_4424,N_4342);
nand U5776 (N_5776,N_4286,N_4079);
nand U5777 (N_5777,N_4458,N_4054);
nor U5778 (N_5778,N_4745,N_4784);
nand U5779 (N_5779,N_4334,N_4468);
nor U5780 (N_5780,N_4488,N_4011);
and U5781 (N_5781,N_4838,N_4896);
or U5782 (N_5782,N_4837,N_4194);
nand U5783 (N_5783,N_4294,N_4060);
and U5784 (N_5784,N_4972,N_4182);
and U5785 (N_5785,N_4036,N_4566);
nor U5786 (N_5786,N_4260,N_4152);
nand U5787 (N_5787,N_4730,N_4874);
xor U5788 (N_5788,N_4506,N_4368);
nand U5789 (N_5789,N_4949,N_4183);
nand U5790 (N_5790,N_4699,N_4866);
or U5791 (N_5791,N_4538,N_4950);
and U5792 (N_5792,N_4993,N_4814);
nor U5793 (N_5793,N_4010,N_4517);
or U5794 (N_5794,N_4525,N_4215);
xnor U5795 (N_5795,N_4491,N_4921);
and U5796 (N_5796,N_4357,N_4133);
or U5797 (N_5797,N_4965,N_4586);
nor U5798 (N_5798,N_4808,N_4341);
nor U5799 (N_5799,N_4469,N_4503);
nor U5800 (N_5800,N_4137,N_4082);
or U5801 (N_5801,N_4698,N_4393);
and U5802 (N_5802,N_4792,N_4961);
and U5803 (N_5803,N_4254,N_4256);
nand U5804 (N_5804,N_4215,N_4085);
and U5805 (N_5805,N_4222,N_4294);
nor U5806 (N_5806,N_4026,N_4275);
and U5807 (N_5807,N_4319,N_4574);
or U5808 (N_5808,N_4302,N_4514);
nor U5809 (N_5809,N_4331,N_4749);
nand U5810 (N_5810,N_4349,N_4783);
nand U5811 (N_5811,N_4612,N_4392);
nand U5812 (N_5812,N_4061,N_4227);
or U5813 (N_5813,N_4877,N_4588);
or U5814 (N_5814,N_4231,N_4352);
and U5815 (N_5815,N_4835,N_4097);
or U5816 (N_5816,N_4088,N_4808);
nor U5817 (N_5817,N_4591,N_4657);
xor U5818 (N_5818,N_4858,N_4395);
nor U5819 (N_5819,N_4871,N_4202);
nand U5820 (N_5820,N_4871,N_4345);
xnor U5821 (N_5821,N_4428,N_4555);
and U5822 (N_5822,N_4637,N_4127);
and U5823 (N_5823,N_4963,N_4859);
or U5824 (N_5824,N_4684,N_4947);
or U5825 (N_5825,N_4084,N_4508);
or U5826 (N_5826,N_4142,N_4388);
xnor U5827 (N_5827,N_4266,N_4116);
xor U5828 (N_5828,N_4819,N_4129);
xnor U5829 (N_5829,N_4261,N_4297);
nor U5830 (N_5830,N_4034,N_4237);
xor U5831 (N_5831,N_4778,N_4196);
nor U5832 (N_5832,N_4345,N_4004);
or U5833 (N_5833,N_4437,N_4131);
nand U5834 (N_5834,N_4491,N_4150);
or U5835 (N_5835,N_4679,N_4325);
nand U5836 (N_5836,N_4556,N_4304);
nor U5837 (N_5837,N_4496,N_4528);
nand U5838 (N_5838,N_4894,N_4867);
nor U5839 (N_5839,N_4239,N_4826);
nor U5840 (N_5840,N_4326,N_4054);
nand U5841 (N_5841,N_4453,N_4903);
and U5842 (N_5842,N_4711,N_4973);
xnor U5843 (N_5843,N_4926,N_4341);
nor U5844 (N_5844,N_4066,N_4904);
or U5845 (N_5845,N_4025,N_4516);
nand U5846 (N_5846,N_4125,N_4260);
nand U5847 (N_5847,N_4838,N_4121);
and U5848 (N_5848,N_4242,N_4123);
nor U5849 (N_5849,N_4108,N_4082);
and U5850 (N_5850,N_4027,N_4472);
or U5851 (N_5851,N_4491,N_4937);
and U5852 (N_5852,N_4607,N_4627);
or U5853 (N_5853,N_4472,N_4986);
or U5854 (N_5854,N_4359,N_4935);
nand U5855 (N_5855,N_4270,N_4867);
or U5856 (N_5856,N_4085,N_4283);
nor U5857 (N_5857,N_4022,N_4715);
xor U5858 (N_5858,N_4575,N_4854);
nand U5859 (N_5859,N_4866,N_4521);
or U5860 (N_5860,N_4402,N_4698);
or U5861 (N_5861,N_4746,N_4540);
nor U5862 (N_5862,N_4771,N_4086);
and U5863 (N_5863,N_4547,N_4834);
nor U5864 (N_5864,N_4990,N_4249);
and U5865 (N_5865,N_4468,N_4503);
nand U5866 (N_5866,N_4354,N_4612);
nand U5867 (N_5867,N_4776,N_4467);
and U5868 (N_5868,N_4473,N_4328);
xor U5869 (N_5869,N_4806,N_4883);
and U5870 (N_5870,N_4151,N_4640);
nor U5871 (N_5871,N_4993,N_4462);
nor U5872 (N_5872,N_4327,N_4652);
and U5873 (N_5873,N_4708,N_4102);
nor U5874 (N_5874,N_4372,N_4122);
xor U5875 (N_5875,N_4703,N_4899);
and U5876 (N_5876,N_4531,N_4814);
or U5877 (N_5877,N_4764,N_4648);
nor U5878 (N_5878,N_4683,N_4017);
nor U5879 (N_5879,N_4057,N_4718);
nor U5880 (N_5880,N_4351,N_4514);
nand U5881 (N_5881,N_4820,N_4982);
and U5882 (N_5882,N_4919,N_4253);
nand U5883 (N_5883,N_4043,N_4416);
nand U5884 (N_5884,N_4381,N_4917);
or U5885 (N_5885,N_4166,N_4011);
or U5886 (N_5886,N_4671,N_4762);
or U5887 (N_5887,N_4260,N_4032);
nand U5888 (N_5888,N_4370,N_4670);
and U5889 (N_5889,N_4017,N_4751);
nand U5890 (N_5890,N_4923,N_4694);
and U5891 (N_5891,N_4281,N_4988);
or U5892 (N_5892,N_4532,N_4108);
or U5893 (N_5893,N_4260,N_4985);
nand U5894 (N_5894,N_4797,N_4931);
or U5895 (N_5895,N_4944,N_4737);
or U5896 (N_5896,N_4052,N_4438);
xor U5897 (N_5897,N_4685,N_4861);
or U5898 (N_5898,N_4618,N_4483);
and U5899 (N_5899,N_4371,N_4399);
nor U5900 (N_5900,N_4248,N_4984);
and U5901 (N_5901,N_4718,N_4880);
and U5902 (N_5902,N_4798,N_4175);
nor U5903 (N_5903,N_4329,N_4503);
xnor U5904 (N_5904,N_4437,N_4137);
nor U5905 (N_5905,N_4617,N_4997);
nor U5906 (N_5906,N_4544,N_4501);
and U5907 (N_5907,N_4569,N_4169);
or U5908 (N_5908,N_4240,N_4067);
and U5909 (N_5909,N_4710,N_4728);
nand U5910 (N_5910,N_4014,N_4289);
and U5911 (N_5911,N_4249,N_4589);
and U5912 (N_5912,N_4150,N_4821);
nand U5913 (N_5913,N_4798,N_4532);
nand U5914 (N_5914,N_4929,N_4882);
nor U5915 (N_5915,N_4131,N_4511);
and U5916 (N_5916,N_4707,N_4497);
or U5917 (N_5917,N_4381,N_4667);
xor U5918 (N_5918,N_4734,N_4455);
xor U5919 (N_5919,N_4076,N_4573);
and U5920 (N_5920,N_4145,N_4394);
nand U5921 (N_5921,N_4917,N_4527);
nor U5922 (N_5922,N_4754,N_4969);
or U5923 (N_5923,N_4035,N_4735);
and U5924 (N_5924,N_4286,N_4383);
or U5925 (N_5925,N_4697,N_4097);
nand U5926 (N_5926,N_4990,N_4360);
nand U5927 (N_5927,N_4008,N_4583);
nand U5928 (N_5928,N_4168,N_4380);
nor U5929 (N_5929,N_4057,N_4427);
nand U5930 (N_5930,N_4600,N_4592);
xor U5931 (N_5931,N_4032,N_4698);
and U5932 (N_5932,N_4060,N_4613);
xnor U5933 (N_5933,N_4779,N_4735);
xor U5934 (N_5934,N_4330,N_4067);
nand U5935 (N_5935,N_4882,N_4562);
and U5936 (N_5936,N_4246,N_4684);
and U5937 (N_5937,N_4554,N_4877);
xnor U5938 (N_5938,N_4615,N_4960);
nand U5939 (N_5939,N_4892,N_4085);
and U5940 (N_5940,N_4586,N_4735);
and U5941 (N_5941,N_4014,N_4201);
or U5942 (N_5942,N_4436,N_4336);
or U5943 (N_5943,N_4860,N_4603);
or U5944 (N_5944,N_4009,N_4061);
nand U5945 (N_5945,N_4474,N_4089);
or U5946 (N_5946,N_4452,N_4859);
or U5947 (N_5947,N_4397,N_4667);
nor U5948 (N_5948,N_4204,N_4868);
nor U5949 (N_5949,N_4247,N_4269);
nand U5950 (N_5950,N_4294,N_4036);
and U5951 (N_5951,N_4297,N_4844);
and U5952 (N_5952,N_4614,N_4193);
or U5953 (N_5953,N_4467,N_4594);
nor U5954 (N_5954,N_4979,N_4480);
and U5955 (N_5955,N_4903,N_4247);
nand U5956 (N_5956,N_4923,N_4713);
nand U5957 (N_5957,N_4616,N_4421);
or U5958 (N_5958,N_4576,N_4574);
nand U5959 (N_5959,N_4278,N_4623);
or U5960 (N_5960,N_4272,N_4456);
or U5961 (N_5961,N_4227,N_4560);
or U5962 (N_5962,N_4058,N_4049);
and U5963 (N_5963,N_4617,N_4133);
or U5964 (N_5964,N_4330,N_4339);
or U5965 (N_5965,N_4026,N_4826);
or U5966 (N_5966,N_4557,N_4370);
nor U5967 (N_5967,N_4693,N_4661);
and U5968 (N_5968,N_4476,N_4985);
nor U5969 (N_5969,N_4790,N_4486);
xnor U5970 (N_5970,N_4093,N_4696);
nor U5971 (N_5971,N_4553,N_4306);
and U5972 (N_5972,N_4557,N_4261);
xnor U5973 (N_5973,N_4078,N_4054);
and U5974 (N_5974,N_4758,N_4293);
or U5975 (N_5975,N_4512,N_4396);
or U5976 (N_5976,N_4239,N_4080);
or U5977 (N_5977,N_4138,N_4662);
and U5978 (N_5978,N_4368,N_4551);
nand U5979 (N_5979,N_4229,N_4555);
and U5980 (N_5980,N_4190,N_4697);
xnor U5981 (N_5981,N_4868,N_4257);
nor U5982 (N_5982,N_4743,N_4144);
and U5983 (N_5983,N_4716,N_4146);
or U5984 (N_5984,N_4432,N_4508);
nor U5985 (N_5985,N_4525,N_4482);
and U5986 (N_5986,N_4025,N_4730);
xor U5987 (N_5987,N_4633,N_4259);
or U5988 (N_5988,N_4009,N_4135);
nor U5989 (N_5989,N_4772,N_4960);
nor U5990 (N_5990,N_4603,N_4554);
nor U5991 (N_5991,N_4248,N_4457);
or U5992 (N_5992,N_4732,N_4249);
nor U5993 (N_5993,N_4708,N_4630);
and U5994 (N_5994,N_4440,N_4790);
and U5995 (N_5995,N_4218,N_4708);
or U5996 (N_5996,N_4705,N_4585);
nand U5997 (N_5997,N_4499,N_4873);
and U5998 (N_5998,N_4227,N_4315);
and U5999 (N_5999,N_4820,N_4882);
nor U6000 (N_6000,N_5545,N_5989);
nor U6001 (N_6001,N_5039,N_5296);
nand U6002 (N_6002,N_5065,N_5647);
and U6003 (N_6003,N_5575,N_5873);
xnor U6004 (N_6004,N_5045,N_5083);
nand U6005 (N_6005,N_5210,N_5872);
xnor U6006 (N_6006,N_5659,N_5132);
xor U6007 (N_6007,N_5156,N_5202);
or U6008 (N_6008,N_5828,N_5255);
xnor U6009 (N_6009,N_5500,N_5302);
nor U6010 (N_6010,N_5108,N_5766);
or U6011 (N_6011,N_5152,N_5022);
or U6012 (N_6012,N_5008,N_5295);
nand U6013 (N_6013,N_5087,N_5637);
xor U6014 (N_6014,N_5369,N_5301);
or U6015 (N_6015,N_5898,N_5436);
nand U6016 (N_6016,N_5116,N_5126);
and U6017 (N_6017,N_5394,N_5829);
or U6018 (N_6018,N_5053,N_5088);
nand U6019 (N_6019,N_5100,N_5891);
xor U6020 (N_6020,N_5485,N_5908);
and U6021 (N_6021,N_5334,N_5316);
xor U6022 (N_6022,N_5502,N_5358);
nand U6023 (N_6023,N_5398,N_5158);
or U6024 (N_6024,N_5818,N_5609);
nor U6025 (N_6025,N_5760,N_5952);
or U6026 (N_6026,N_5694,N_5017);
nor U6027 (N_6027,N_5538,N_5486);
and U6028 (N_6028,N_5598,N_5174);
or U6029 (N_6029,N_5875,N_5115);
nor U6030 (N_6030,N_5527,N_5804);
and U6031 (N_6031,N_5374,N_5874);
nand U6032 (N_6032,N_5733,N_5880);
or U6033 (N_6033,N_5676,N_5988);
or U6034 (N_6034,N_5376,N_5762);
xor U6035 (N_6035,N_5916,N_5712);
or U6036 (N_6036,N_5550,N_5761);
and U6037 (N_6037,N_5275,N_5863);
or U6038 (N_6038,N_5458,N_5680);
xor U6039 (N_6039,N_5972,N_5672);
or U6040 (N_6040,N_5936,N_5404);
or U6041 (N_6041,N_5477,N_5077);
and U6042 (N_6042,N_5469,N_5367);
xnor U6043 (N_6043,N_5529,N_5014);
and U6044 (N_6044,N_5998,N_5810);
xor U6045 (N_6045,N_5879,N_5127);
nor U6046 (N_6046,N_5385,N_5582);
and U6047 (N_6047,N_5101,N_5870);
or U6048 (N_6048,N_5889,N_5573);
or U6049 (N_6049,N_5270,N_5516);
or U6050 (N_6050,N_5885,N_5262);
nand U6051 (N_6051,N_5946,N_5758);
xnor U6052 (N_6052,N_5211,N_5608);
and U6053 (N_6053,N_5589,N_5024);
xor U6054 (N_6054,N_5695,N_5504);
nand U6055 (N_6055,N_5777,N_5491);
nand U6056 (N_6056,N_5806,N_5556);
nand U6057 (N_6057,N_5452,N_5093);
and U6058 (N_6058,N_5876,N_5652);
and U6059 (N_6059,N_5416,N_5624);
and U6060 (N_6060,N_5945,N_5483);
or U6061 (N_6061,N_5434,N_5382);
or U6062 (N_6062,N_5217,N_5537);
nor U6063 (N_6063,N_5744,N_5714);
and U6064 (N_6064,N_5172,N_5613);
nand U6065 (N_6065,N_5058,N_5786);
or U6066 (N_6066,N_5449,N_5525);
nor U6067 (N_6067,N_5599,N_5431);
nand U6068 (N_6068,N_5967,N_5727);
and U6069 (N_6069,N_5759,N_5897);
nand U6070 (N_6070,N_5182,N_5283);
and U6071 (N_6071,N_5159,N_5413);
and U6072 (N_6072,N_5441,N_5932);
or U6073 (N_6073,N_5464,N_5845);
and U6074 (N_6074,N_5682,N_5837);
xor U6075 (N_6075,N_5277,N_5164);
nand U6076 (N_6076,N_5492,N_5512);
and U6077 (N_6077,N_5754,N_5992);
nand U6078 (N_6078,N_5388,N_5420);
and U6079 (N_6079,N_5995,N_5004);
nor U6080 (N_6080,N_5300,N_5197);
nand U6081 (N_6081,N_5196,N_5639);
xnor U6082 (N_6082,N_5463,N_5604);
xnor U6083 (N_6083,N_5042,N_5403);
nand U6084 (N_6084,N_5969,N_5662);
and U6085 (N_6085,N_5980,N_5240);
and U6086 (N_6086,N_5025,N_5865);
or U6087 (N_6087,N_5813,N_5585);
or U6088 (N_6088,N_5543,N_5185);
nand U6089 (N_6089,N_5113,N_5503);
or U6090 (N_6090,N_5161,N_5553);
nand U6091 (N_6091,N_5232,N_5086);
or U6092 (N_6092,N_5052,N_5352);
xnor U6093 (N_6093,N_5143,N_5827);
nor U6094 (N_6094,N_5982,N_5072);
or U6095 (N_6095,N_5106,N_5227);
or U6096 (N_6096,N_5489,N_5931);
nor U6097 (N_6097,N_5219,N_5805);
xnor U6098 (N_6098,N_5142,N_5443);
nor U6099 (N_6099,N_5993,N_5447);
and U6100 (N_6100,N_5842,N_5344);
nor U6101 (N_6101,N_5298,N_5321);
nand U6102 (N_6102,N_5666,N_5005);
nor U6103 (N_6103,N_5594,N_5834);
nor U6104 (N_6104,N_5702,N_5364);
xnor U6105 (N_6105,N_5281,N_5203);
nor U6106 (N_6106,N_5124,N_5038);
xor U6107 (N_6107,N_5269,N_5168);
nor U6108 (N_6108,N_5332,N_5866);
nand U6109 (N_6109,N_5139,N_5610);
and U6110 (N_6110,N_5985,N_5986);
and U6111 (N_6111,N_5186,N_5401);
or U6112 (N_6112,N_5470,N_5170);
or U6113 (N_6113,N_5214,N_5763);
or U6114 (N_6114,N_5001,N_5011);
and U6115 (N_6115,N_5596,N_5569);
or U6116 (N_6116,N_5435,N_5707);
and U6117 (N_6117,N_5696,N_5723);
nor U6118 (N_6118,N_5944,N_5307);
or U6119 (N_6119,N_5264,N_5822);
and U6120 (N_6120,N_5069,N_5780);
xor U6121 (N_6121,N_5246,N_5788);
nor U6122 (N_6122,N_5207,N_5465);
xor U6123 (N_6123,N_5824,N_5311);
or U6124 (N_6124,N_5631,N_5261);
nor U6125 (N_6125,N_5542,N_5429);
or U6126 (N_6126,N_5427,N_5071);
nand U6127 (N_6127,N_5131,N_5122);
and U6128 (N_6128,N_5007,N_5798);
or U6129 (N_6129,N_5169,N_5488);
or U6130 (N_6130,N_5239,N_5773);
nand U6131 (N_6131,N_5657,N_5724);
and U6132 (N_6132,N_5082,N_5817);
nor U6133 (N_6133,N_5700,N_5109);
nand U6134 (N_6134,N_5271,N_5858);
xor U6135 (N_6135,N_5628,N_5848);
or U6136 (N_6136,N_5366,N_5384);
xnor U6137 (N_6137,N_5336,N_5918);
nor U6138 (N_6138,N_5233,N_5578);
nor U6139 (N_6139,N_5851,N_5854);
or U6140 (N_6140,N_5319,N_5655);
xor U6141 (N_6141,N_5493,N_5481);
and U6142 (N_6142,N_5948,N_5941);
nand U6143 (N_6143,N_5559,N_5654);
nor U6144 (N_6144,N_5000,N_5642);
xnor U6145 (N_6145,N_5424,N_5593);
and U6146 (N_6146,N_5426,N_5446);
nand U6147 (N_6147,N_5351,N_5286);
and U6148 (N_6148,N_5141,N_5835);
nor U6149 (N_6149,N_5526,N_5949);
nor U6150 (N_6150,N_5860,N_5965);
nor U6151 (N_6151,N_5976,N_5297);
nor U6152 (N_6152,N_5480,N_5510);
nand U6153 (N_6153,N_5135,N_5970);
nand U6154 (N_6154,N_5354,N_5035);
nand U6155 (N_6155,N_5140,N_5641);
nand U6156 (N_6156,N_5368,N_5062);
or U6157 (N_6157,N_5670,N_5231);
nand U6158 (N_6158,N_5074,N_5797);
nand U6159 (N_6159,N_5268,N_5815);
nor U6160 (N_6160,N_5840,N_5034);
nand U6161 (N_6161,N_5428,N_5939);
or U6162 (N_6162,N_5318,N_5868);
or U6163 (N_6163,N_5922,N_5392);
or U6164 (N_6164,N_5414,N_5685);
nand U6165 (N_6165,N_5557,N_5807);
nor U6166 (N_6166,N_5563,N_5341);
or U6167 (N_6167,N_5450,N_5893);
and U6168 (N_6168,N_5630,N_5611);
nor U6169 (N_6169,N_5208,N_5079);
nor U6170 (N_6170,N_5479,N_5096);
or U6171 (N_6171,N_5558,N_5357);
or U6172 (N_6172,N_5323,N_5471);
xor U6173 (N_6173,N_5044,N_5439);
and U6174 (N_6174,N_5864,N_5279);
and U6175 (N_6175,N_5617,N_5406);
and U6176 (N_6176,N_5451,N_5548);
nor U6177 (N_6177,N_5244,N_5956);
nand U6178 (N_6178,N_5583,N_5390);
or U6179 (N_6179,N_5473,N_5950);
nand U6180 (N_6180,N_5725,N_5770);
or U6181 (N_6181,N_5343,N_5935);
nand U6182 (N_6182,N_5484,N_5595);
nor U6183 (N_6183,N_5112,N_5783);
or U6184 (N_6184,N_5110,N_5372);
or U6185 (N_6185,N_5934,N_5900);
nor U6186 (N_6186,N_5460,N_5187);
nand U6187 (N_6187,N_5160,N_5789);
or U6188 (N_6188,N_5119,N_5561);
or U6189 (N_6189,N_5509,N_5991);
and U6190 (N_6190,N_5066,N_5448);
and U6191 (N_6191,N_5117,N_5644);
or U6192 (N_6192,N_5816,N_5792);
xnor U6193 (N_6193,N_5650,N_5528);
nor U6194 (N_6194,N_5686,N_5658);
nor U6195 (N_6195,N_5205,N_5199);
and U6196 (N_6196,N_5524,N_5955);
and U6197 (N_6197,N_5123,N_5060);
or U6198 (N_6198,N_5974,N_5303);
and U6199 (N_6199,N_5960,N_5314);
or U6200 (N_6200,N_5811,N_5511);
or U6201 (N_6201,N_5507,N_5825);
or U6202 (N_6202,N_5252,N_5943);
xor U6203 (N_6203,N_5907,N_5085);
nor U6204 (N_6204,N_5328,N_5966);
and U6205 (N_6205,N_5619,N_5091);
nor U6206 (N_6206,N_5013,N_5289);
or U6207 (N_6207,N_5084,N_5983);
nand U6208 (N_6208,N_5353,N_5395);
nor U6209 (N_6209,N_5692,N_5615);
nand U6210 (N_6210,N_5250,N_5517);
nand U6211 (N_6211,N_5348,N_5892);
or U6212 (N_6212,N_5664,N_5153);
and U6213 (N_6213,N_5740,N_5016);
nor U6214 (N_6214,N_5688,N_5911);
xnor U6215 (N_6215,N_5968,N_5535);
or U6216 (N_6216,N_5570,N_5691);
nor U6217 (N_6217,N_5601,N_5444);
or U6218 (N_6218,N_5412,N_5154);
or U6219 (N_6219,N_5961,N_5812);
or U6220 (N_6220,N_5309,N_5393);
nor U6221 (N_6221,N_5979,N_5947);
or U6222 (N_6222,N_5743,N_5146);
xor U6223 (N_6223,N_5803,N_5081);
and U6224 (N_6224,N_5386,N_5549);
nand U6225 (N_6225,N_5746,N_5705);
and U6226 (N_6226,N_5661,N_5994);
or U6227 (N_6227,N_5793,N_5587);
and U6228 (N_6228,N_5750,N_5973);
nor U6229 (N_6229,N_5605,N_5711);
nor U6230 (N_6230,N_5335,N_5304);
and U6231 (N_6231,N_5814,N_5389);
and U6232 (N_6232,N_5718,N_5057);
xor U6233 (N_6233,N_5090,N_5363);
and U6234 (N_6234,N_5775,N_5346);
nor U6235 (N_6235,N_5247,N_5399);
nand U6236 (N_6236,N_5177,N_5467);
or U6237 (N_6237,N_5166,N_5667);
xor U6238 (N_6238,N_5098,N_5753);
or U6239 (N_6239,N_5468,N_5248);
nand U6240 (N_6240,N_5663,N_5047);
nor U6241 (N_6241,N_5534,N_5306);
xor U6242 (N_6242,N_5099,N_5713);
nor U6243 (N_6243,N_5536,N_5926);
nor U6244 (N_6244,N_5669,N_5462);
nand U6245 (N_6245,N_5522,N_5523);
nand U6246 (N_6246,N_5736,N_5791);
and U6247 (N_6247,N_5590,N_5033);
nor U6248 (N_6248,N_5929,N_5405);
nor U6249 (N_6249,N_5129,N_5597);
nor U6250 (N_6250,N_5653,N_5906);
nand U6251 (N_6251,N_5322,N_5681);
and U6252 (N_6252,N_5173,N_5704);
xor U6253 (N_6253,N_5826,N_5472);
and U6254 (N_6254,N_5576,N_5496);
and U6255 (N_6255,N_5719,N_5337);
and U6256 (N_6256,N_5012,N_5795);
and U6257 (N_6257,N_5540,N_5331);
nand U6258 (N_6258,N_5189,N_5506);
and U6259 (N_6259,N_5338,N_5915);
nor U6260 (N_6260,N_5820,N_5380);
nor U6261 (N_6261,N_5254,N_5138);
nand U6262 (N_6262,N_5317,N_5417);
nor U6263 (N_6263,N_5032,N_5877);
and U6264 (N_6264,N_5379,N_5291);
nand U6265 (N_6265,N_5194,N_5285);
xor U6266 (N_6266,N_5292,N_5720);
nand U6267 (N_6267,N_5329,N_5019);
or U6268 (N_6268,N_5241,N_5562);
xor U6269 (N_6269,N_5716,N_5027);
nor U6270 (N_6270,N_5018,N_5310);
nand U6271 (N_6271,N_5155,N_5768);
xor U6272 (N_6272,N_5678,N_5373);
nor U6273 (N_6273,N_5103,N_5381);
and U6274 (N_6274,N_5784,N_5913);
nand U6275 (N_6275,N_5176,N_5061);
nor U6276 (N_6276,N_5499,N_5180);
nor U6277 (N_6277,N_5130,N_5128);
and U6278 (N_6278,N_5769,N_5881);
or U6279 (N_6279,N_5201,N_5717);
or U6280 (N_6280,N_5819,N_5709);
or U6281 (N_6281,N_5067,N_5895);
and U6282 (N_6282,N_5163,N_5095);
or U6283 (N_6283,N_5050,N_5755);
or U6284 (N_6284,N_5555,N_5422);
and U6285 (N_6285,N_5799,N_5320);
or U6286 (N_6286,N_5178,N_5251);
nor U6287 (N_6287,N_5150,N_5305);
xnor U6288 (N_6288,N_5411,N_5673);
or U6289 (N_6289,N_5097,N_5779);
nor U6290 (N_6290,N_5263,N_5752);
and U6291 (N_6291,N_5706,N_5102);
nand U6292 (N_6292,N_5914,N_5294);
and U6293 (N_6293,N_5359,N_5757);
and U6294 (N_6294,N_5518,N_5635);
and U6295 (N_6295,N_5508,N_5764);
nor U6296 (N_6296,N_5697,N_5782);
nor U6297 (N_6297,N_5776,N_5839);
and U6298 (N_6298,N_5574,N_5930);
or U6299 (N_6299,N_5572,N_5505);
nand U6300 (N_6300,N_5882,N_5886);
nor U6301 (N_6301,N_5687,N_5342);
xnor U6302 (N_6302,N_5772,N_5094);
nor U6303 (N_6303,N_5721,N_5482);
and U6304 (N_6304,N_5888,N_5532);
nand U6305 (N_6305,N_5977,N_5076);
or U6306 (N_6306,N_5220,N_5188);
or U6307 (N_6307,N_5919,N_5756);
nor U6308 (N_6308,N_5588,N_5841);
nand U6309 (N_6309,N_5212,N_5409);
or U6310 (N_6310,N_5925,N_5501);
or U6311 (N_6311,N_5747,N_5036);
or U6312 (N_6312,N_5771,N_5355);
nor U6313 (N_6313,N_5902,N_5010);
nand U6314 (N_6314,N_5984,N_5433);
nor U6315 (N_6315,N_5903,N_5148);
nor U6316 (N_6316,N_5387,N_5075);
nor U6317 (N_6317,N_5046,N_5461);
nor U6318 (N_6318,N_5415,N_5288);
and U6319 (N_6319,N_5040,N_5551);
and U6320 (N_6320,N_5831,N_5715);
nand U6321 (N_6321,N_5498,N_5147);
or U6322 (N_6322,N_5190,N_5937);
nor U6323 (N_6323,N_5282,N_5396);
or U6324 (N_6324,N_5636,N_5923);
xnor U6325 (N_6325,N_5136,N_5204);
nand U6326 (N_6326,N_5849,N_5996);
nor U6327 (N_6327,N_5371,N_5584);
nand U6328 (N_6328,N_5894,N_5568);
or U6329 (N_6329,N_5571,N_5333);
nand U6330 (N_6330,N_5869,N_5266);
nand U6331 (N_6331,N_5738,N_5515);
nand U6332 (N_6332,N_5445,N_5603);
or U6333 (N_6333,N_5229,N_5632);
and U6334 (N_6334,N_5978,N_5226);
xnor U6335 (N_6335,N_5361,N_5209);
nand U6336 (N_6336,N_5037,N_5326);
nor U6337 (N_6337,N_5808,N_5253);
nor U6338 (N_6338,N_5735,N_5475);
and U6339 (N_6339,N_5728,N_5003);
xor U6340 (N_6340,N_5802,N_5238);
nand U6341 (N_6341,N_5698,N_5221);
nor U6342 (N_6342,N_5377,N_5265);
and U6343 (N_6343,N_5618,N_5887);
or U6344 (N_6344,N_5092,N_5951);
nand U6345 (N_6345,N_5577,N_5175);
nor U6346 (N_6346,N_5623,N_5620);
xor U6347 (N_6347,N_5063,N_5833);
nor U6348 (N_6348,N_5015,N_5519);
xnor U6349 (N_6349,N_5459,N_5726);
or U6350 (N_6350,N_5999,N_5048);
and U6351 (N_6351,N_5181,N_5162);
nand U6352 (N_6352,N_5684,N_5963);
nand U6353 (N_6353,N_5896,N_5378);
nand U6354 (N_6354,N_5616,N_5104);
nand U6355 (N_6355,N_5683,N_5213);
or U6356 (N_6356,N_5218,N_5474);
or U6357 (N_6357,N_5838,N_5645);
xor U6358 (N_6358,N_5689,N_5054);
or U6359 (N_6359,N_5455,N_5237);
xnor U6360 (N_6360,N_5494,N_5612);
xnor U6361 (N_6361,N_5677,N_5442);
or U6362 (N_6362,N_5668,N_5224);
nor U6363 (N_6363,N_5990,N_5339);
or U6364 (N_6364,N_5179,N_5850);
xnor U6365 (N_6365,N_5308,N_5809);
nor U6366 (N_6366,N_5137,N_5068);
or U6367 (N_6367,N_5049,N_5051);
or U6368 (N_6368,N_5729,N_5064);
nor U6369 (N_6369,N_5749,N_5546);
nand U6370 (N_6370,N_5638,N_5745);
nand U6371 (N_6371,N_5924,N_5794);
xor U6372 (N_6372,N_5671,N_5293);
nor U6373 (N_6373,N_5586,N_5591);
or U6374 (N_6374,N_5391,N_5890);
nand U6375 (N_6375,N_5114,N_5345);
or U6376 (N_6376,N_5859,N_5272);
and U6377 (N_6377,N_5454,N_5778);
or U6378 (N_6378,N_5975,N_5222);
nand U6379 (N_6379,N_5765,N_5002);
xor U6380 (N_6380,N_5330,N_5656);
nor U6381 (N_6381,N_5634,N_5497);
nand U6382 (N_6382,N_5312,N_5144);
nor U6383 (N_6383,N_5847,N_5080);
and U6384 (N_6384,N_5958,N_5324);
nor U6385 (N_6385,N_5120,N_5901);
nor U6386 (N_6386,N_5495,N_5862);
or U6387 (N_6387,N_5513,N_5767);
nor U6388 (N_6388,N_5009,N_5260);
or U6389 (N_6389,N_5235,N_5157);
nand U6390 (N_6390,N_5626,N_5751);
nand U6391 (N_6391,N_5402,N_5453);
or U6392 (N_6392,N_5739,N_5478);
nor U6393 (N_6393,N_5029,N_5910);
or U6394 (N_6394,N_5927,N_5737);
or U6395 (N_6395,N_5622,N_5206);
nor U6396 (N_6396,N_5151,N_5423);
nand U6397 (N_6397,N_5884,N_5846);
nand U6398 (N_6398,N_5230,N_5006);
and U6399 (N_6399,N_5940,N_5383);
nand U6400 (N_6400,N_5649,N_5942);
nor U6401 (N_6401,N_5781,N_5962);
nand U6402 (N_6402,N_5957,N_5920);
nor U6403 (N_6403,N_5933,N_5184);
or U6404 (N_6404,N_5690,N_5325);
or U6405 (N_6405,N_5362,N_5432);
or U6406 (N_6406,N_5350,N_5917);
nand U6407 (N_6407,N_5710,N_5349);
and U6408 (N_6408,N_5476,N_5273);
nor U6409 (N_6409,N_5964,N_5228);
nand U6410 (N_6410,N_5056,N_5836);
nor U6411 (N_6411,N_5953,N_5857);
nor U6412 (N_6412,N_5853,N_5021);
nand U6413 (N_6413,N_5356,N_5111);
nor U6414 (N_6414,N_5938,N_5340);
nor U6415 (N_6415,N_5198,N_5397);
xnor U6416 (N_6416,N_5365,N_5679);
and U6417 (N_6417,N_5871,N_5200);
nor U6418 (N_6418,N_5133,N_5245);
nand U6419 (N_6419,N_5419,N_5215);
nand U6420 (N_6420,N_5375,N_5959);
nor U6421 (N_6421,N_5801,N_5565);
xor U6422 (N_6422,N_5466,N_5708);
or U6423 (N_6423,N_5370,N_5912);
nand U6424 (N_6424,N_5257,N_5665);
or U6425 (N_6425,N_5734,N_5055);
nor U6426 (N_6426,N_5242,N_5790);
xnor U6427 (N_6427,N_5832,N_5742);
and U6428 (N_6428,N_5438,N_5701);
or U6429 (N_6429,N_5287,N_5675);
or U6430 (N_6430,N_5089,N_5059);
nand U6431 (N_6431,N_5487,N_5078);
nand U6432 (N_6432,N_5430,N_5703);
or U6433 (N_6433,N_5928,N_5579);
nor U6434 (N_6434,N_5315,N_5073);
nand U6435 (N_6435,N_5347,N_5730);
nor U6436 (N_6436,N_5830,N_5149);
nor U6437 (N_6437,N_5627,N_5566);
or U6438 (N_6438,N_5225,N_5787);
nor U6439 (N_6439,N_5023,N_5276);
or U6440 (N_6440,N_5861,N_5852);
nor U6441 (N_6441,N_5541,N_5410);
or U6442 (N_6442,N_5785,N_5284);
nand U6443 (N_6443,N_5674,N_5651);
xor U6444 (N_6444,N_5621,N_5606);
and U6445 (N_6445,N_5560,N_5552);
nand U6446 (N_6446,N_5105,N_5490);
nand U6447 (N_6447,N_5521,N_5121);
nor U6448 (N_6448,N_5193,N_5192);
xor U6449 (N_6449,N_5625,N_5554);
or U6450 (N_6450,N_5531,N_5125);
and U6451 (N_6451,N_5418,N_5020);
nor U6452 (N_6452,N_5183,N_5171);
nand U6453 (N_6453,N_5564,N_5514);
xnor U6454 (N_6454,N_5258,N_5425);
or U6455 (N_6455,N_5437,N_5165);
xor U6456 (N_6456,N_5823,N_5290);
nor U6457 (N_6457,N_5299,N_5741);
and U6458 (N_6458,N_5070,N_5167);
or U6459 (N_6459,N_5134,N_5581);
or U6460 (N_6460,N_5580,N_5774);
nor U6461 (N_6461,N_5732,N_5456);
or U6462 (N_6462,N_5267,N_5646);
or U6463 (N_6463,N_5195,N_5904);
nor U6464 (N_6464,N_5614,N_5280);
nor U6465 (N_6465,N_5234,N_5748);
nand U6466 (N_6466,N_5028,N_5660);
nor U6467 (N_6467,N_5592,N_5278);
or U6468 (N_6468,N_5643,N_5256);
nand U6469 (N_6469,N_5699,N_5457);
nand U6470 (N_6470,N_5800,N_5031);
or U6471 (N_6471,N_5360,N_5600);
nor U6472 (N_6472,N_5633,N_5856);
nor U6473 (N_6473,N_5407,N_5987);
nor U6474 (N_6474,N_5145,N_5981);
nand U6475 (N_6475,N_5216,N_5693);
nand U6476 (N_6476,N_5921,N_5030);
nand U6477 (N_6477,N_5533,N_5629);
xor U6478 (N_6478,N_5883,N_5421);
nor U6479 (N_6479,N_5313,N_5259);
and U6480 (N_6480,N_5547,N_5236);
xor U6481 (N_6481,N_5843,N_5878);
nand U6482 (N_6482,N_5722,N_5867);
or U6483 (N_6483,N_5327,N_5107);
or U6484 (N_6484,N_5041,N_5899);
nor U6485 (N_6485,N_5520,N_5408);
and U6486 (N_6486,N_5544,N_5043);
or U6487 (N_6487,N_5026,N_5530);
and U6488 (N_6488,N_5821,N_5118);
and U6489 (N_6489,N_5997,N_5191);
nand U6490 (N_6490,N_5223,N_5440);
nor U6491 (N_6491,N_5855,N_5905);
nand U6492 (N_6492,N_5796,N_5274);
and U6493 (N_6493,N_5971,N_5539);
or U6494 (N_6494,N_5249,N_5731);
nand U6495 (N_6495,N_5400,N_5602);
or U6496 (N_6496,N_5648,N_5909);
and U6497 (N_6497,N_5844,N_5243);
xnor U6498 (N_6498,N_5567,N_5640);
and U6499 (N_6499,N_5954,N_5607);
nor U6500 (N_6500,N_5419,N_5646);
nor U6501 (N_6501,N_5921,N_5519);
xor U6502 (N_6502,N_5479,N_5371);
nand U6503 (N_6503,N_5853,N_5334);
and U6504 (N_6504,N_5182,N_5329);
or U6505 (N_6505,N_5916,N_5245);
nand U6506 (N_6506,N_5219,N_5423);
nand U6507 (N_6507,N_5495,N_5405);
xnor U6508 (N_6508,N_5427,N_5925);
and U6509 (N_6509,N_5747,N_5498);
and U6510 (N_6510,N_5383,N_5025);
or U6511 (N_6511,N_5525,N_5500);
xor U6512 (N_6512,N_5774,N_5592);
or U6513 (N_6513,N_5379,N_5149);
and U6514 (N_6514,N_5688,N_5056);
nor U6515 (N_6515,N_5910,N_5228);
nand U6516 (N_6516,N_5318,N_5748);
nor U6517 (N_6517,N_5999,N_5363);
or U6518 (N_6518,N_5643,N_5383);
nor U6519 (N_6519,N_5050,N_5905);
or U6520 (N_6520,N_5237,N_5266);
or U6521 (N_6521,N_5850,N_5886);
nor U6522 (N_6522,N_5060,N_5715);
and U6523 (N_6523,N_5290,N_5438);
nor U6524 (N_6524,N_5849,N_5454);
nand U6525 (N_6525,N_5359,N_5604);
xor U6526 (N_6526,N_5539,N_5255);
nand U6527 (N_6527,N_5555,N_5900);
nand U6528 (N_6528,N_5519,N_5406);
or U6529 (N_6529,N_5180,N_5896);
nor U6530 (N_6530,N_5287,N_5714);
nor U6531 (N_6531,N_5161,N_5610);
xnor U6532 (N_6532,N_5022,N_5829);
xnor U6533 (N_6533,N_5032,N_5523);
and U6534 (N_6534,N_5707,N_5361);
or U6535 (N_6535,N_5025,N_5220);
xnor U6536 (N_6536,N_5439,N_5982);
nand U6537 (N_6537,N_5323,N_5631);
nor U6538 (N_6538,N_5400,N_5229);
nand U6539 (N_6539,N_5215,N_5696);
or U6540 (N_6540,N_5779,N_5844);
or U6541 (N_6541,N_5407,N_5653);
nor U6542 (N_6542,N_5407,N_5105);
or U6543 (N_6543,N_5687,N_5688);
and U6544 (N_6544,N_5375,N_5565);
nand U6545 (N_6545,N_5331,N_5486);
nand U6546 (N_6546,N_5956,N_5231);
xnor U6547 (N_6547,N_5705,N_5337);
xor U6548 (N_6548,N_5438,N_5066);
and U6549 (N_6549,N_5489,N_5406);
or U6550 (N_6550,N_5523,N_5331);
or U6551 (N_6551,N_5062,N_5850);
or U6552 (N_6552,N_5611,N_5134);
nor U6553 (N_6553,N_5498,N_5586);
and U6554 (N_6554,N_5260,N_5807);
and U6555 (N_6555,N_5748,N_5541);
xor U6556 (N_6556,N_5073,N_5957);
nor U6557 (N_6557,N_5255,N_5904);
or U6558 (N_6558,N_5914,N_5389);
xor U6559 (N_6559,N_5353,N_5770);
nand U6560 (N_6560,N_5617,N_5456);
and U6561 (N_6561,N_5869,N_5291);
or U6562 (N_6562,N_5141,N_5696);
or U6563 (N_6563,N_5751,N_5337);
nand U6564 (N_6564,N_5800,N_5357);
nand U6565 (N_6565,N_5892,N_5063);
nand U6566 (N_6566,N_5926,N_5391);
xnor U6567 (N_6567,N_5572,N_5106);
and U6568 (N_6568,N_5785,N_5279);
nand U6569 (N_6569,N_5585,N_5794);
nand U6570 (N_6570,N_5816,N_5413);
nand U6571 (N_6571,N_5882,N_5436);
or U6572 (N_6572,N_5288,N_5948);
xnor U6573 (N_6573,N_5941,N_5504);
nor U6574 (N_6574,N_5997,N_5048);
nand U6575 (N_6575,N_5545,N_5067);
or U6576 (N_6576,N_5902,N_5768);
nand U6577 (N_6577,N_5761,N_5082);
and U6578 (N_6578,N_5896,N_5971);
nand U6579 (N_6579,N_5900,N_5090);
nor U6580 (N_6580,N_5460,N_5723);
nor U6581 (N_6581,N_5337,N_5021);
xor U6582 (N_6582,N_5421,N_5720);
nand U6583 (N_6583,N_5983,N_5967);
or U6584 (N_6584,N_5889,N_5996);
nand U6585 (N_6585,N_5962,N_5130);
nand U6586 (N_6586,N_5958,N_5529);
nor U6587 (N_6587,N_5636,N_5011);
and U6588 (N_6588,N_5576,N_5057);
and U6589 (N_6589,N_5942,N_5151);
or U6590 (N_6590,N_5944,N_5387);
and U6591 (N_6591,N_5610,N_5708);
or U6592 (N_6592,N_5026,N_5186);
nand U6593 (N_6593,N_5227,N_5389);
or U6594 (N_6594,N_5700,N_5043);
or U6595 (N_6595,N_5667,N_5914);
and U6596 (N_6596,N_5170,N_5280);
or U6597 (N_6597,N_5806,N_5199);
and U6598 (N_6598,N_5156,N_5472);
or U6599 (N_6599,N_5418,N_5902);
nor U6600 (N_6600,N_5311,N_5590);
xor U6601 (N_6601,N_5735,N_5015);
nand U6602 (N_6602,N_5550,N_5628);
or U6603 (N_6603,N_5666,N_5281);
or U6604 (N_6604,N_5883,N_5367);
nand U6605 (N_6605,N_5314,N_5600);
and U6606 (N_6606,N_5316,N_5745);
nor U6607 (N_6607,N_5296,N_5490);
xnor U6608 (N_6608,N_5578,N_5066);
nor U6609 (N_6609,N_5401,N_5397);
nor U6610 (N_6610,N_5659,N_5123);
nor U6611 (N_6611,N_5251,N_5290);
nor U6612 (N_6612,N_5360,N_5837);
nor U6613 (N_6613,N_5311,N_5481);
xor U6614 (N_6614,N_5242,N_5032);
and U6615 (N_6615,N_5198,N_5516);
xor U6616 (N_6616,N_5005,N_5682);
and U6617 (N_6617,N_5496,N_5126);
and U6618 (N_6618,N_5969,N_5268);
and U6619 (N_6619,N_5669,N_5112);
or U6620 (N_6620,N_5695,N_5854);
xnor U6621 (N_6621,N_5746,N_5210);
nor U6622 (N_6622,N_5933,N_5862);
nor U6623 (N_6623,N_5220,N_5621);
nand U6624 (N_6624,N_5890,N_5528);
nor U6625 (N_6625,N_5450,N_5159);
nor U6626 (N_6626,N_5581,N_5841);
nand U6627 (N_6627,N_5552,N_5647);
nand U6628 (N_6628,N_5973,N_5383);
or U6629 (N_6629,N_5699,N_5711);
nor U6630 (N_6630,N_5978,N_5358);
nand U6631 (N_6631,N_5403,N_5916);
and U6632 (N_6632,N_5195,N_5163);
nor U6633 (N_6633,N_5677,N_5544);
nand U6634 (N_6634,N_5765,N_5256);
nand U6635 (N_6635,N_5148,N_5719);
nor U6636 (N_6636,N_5256,N_5523);
and U6637 (N_6637,N_5377,N_5708);
nand U6638 (N_6638,N_5939,N_5192);
or U6639 (N_6639,N_5678,N_5795);
nor U6640 (N_6640,N_5812,N_5062);
and U6641 (N_6641,N_5103,N_5073);
nand U6642 (N_6642,N_5849,N_5165);
and U6643 (N_6643,N_5128,N_5807);
and U6644 (N_6644,N_5038,N_5421);
nor U6645 (N_6645,N_5411,N_5004);
xnor U6646 (N_6646,N_5265,N_5216);
nor U6647 (N_6647,N_5622,N_5906);
and U6648 (N_6648,N_5582,N_5556);
xnor U6649 (N_6649,N_5355,N_5327);
nand U6650 (N_6650,N_5423,N_5230);
or U6651 (N_6651,N_5893,N_5552);
and U6652 (N_6652,N_5942,N_5842);
nor U6653 (N_6653,N_5168,N_5932);
xor U6654 (N_6654,N_5859,N_5023);
or U6655 (N_6655,N_5121,N_5084);
and U6656 (N_6656,N_5120,N_5379);
and U6657 (N_6657,N_5959,N_5990);
and U6658 (N_6658,N_5935,N_5102);
and U6659 (N_6659,N_5402,N_5086);
or U6660 (N_6660,N_5104,N_5207);
nand U6661 (N_6661,N_5765,N_5100);
xor U6662 (N_6662,N_5083,N_5644);
or U6663 (N_6663,N_5046,N_5491);
xnor U6664 (N_6664,N_5614,N_5089);
and U6665 (N_6665,N_5336,N_5294);
or U6666 (N_6666,N_5793,N_5620);
nor U6667 (N_6667,N_5638,N_5208);
nor U6668 (N_6668,N_5036,N_5399);
or U6669 (N_6669,N_5650,N_5955);
xnor U6670 (N_6670,N_5265,N_5665);
and U6671 (N_6671,N_5815,N_5059);
or U6672 (N_6672,N_5695,N_5626);
nand U6673 (N_6673,N_5392,N_5432);
and U6674 (N_6674,N_5911,N_5313);
or U6675 (N_6675,N_5918,N_5436);
and U6676 (N_6676,N_5312,N_5446);
nor U6677 (N_6677,N_5499,N_5146);
or U6678 (N_6678,N_5074,N_5282);
nor U6679 (N_6679,N_5502,N_5096);
and U6680 (N_6680,N_5829,N_5501);
nand U6681 (N_6681,N_5443,N_5922);
nand U6682 (N_6682,N_5486,N_5337);
or U6683 (N_6683,N_5967,N_5387);
xnor U6684 (N_6684,N_5742,N_5595);
or U6685 (N_6685,N_5278,N_5264);
nor U6686 (N_6686,N_5641,N_5174);
or U6687 (N_6687,N_5237,N_5465);
and U6688 (N_6688,N_5379,N_5760);
and U6689 (N_6689,N_5355,N_5661);
nor U6690 (N_6690,N_5121,N_5353);
nand U6691 (N_6691,N_5672,N_5454);
nand U6692 (N_6692,N_5777,N_5369);
xnor U6693 (N_6693,N_5835,N_5081);
nor U6694 (N_6694,N_5958,N_5960);
or U6695 (N_6695,N_5499,N_5653);
or U6696 (N_6696,N_5578,N_5306);
nand U6697 (N_6697,N_5240,N_5120);
or U6698 (N_6698,N_5984,N_5482);
and U6699 (N_6699,N_5406,N_5858);
and U6700 (N_6700,N_5363,N_5151);
nand U6701 (N_6701,N_5747,N_5042);
nand U6702 (N_6702,N_5249,N_5696);
and U6703 (N_6703,N_5121,N_5130);
and U6704 (N_6704,N_5614,N_5827);
nor U6705 (N_6705,N_5338,N_5822);
xor U6706 (N_6706,N_5448,N_5263);
xor U6707 (N_6707,N_5266,N_5134);
nor U6708 (N_6708,N_5846,N_5107);
nor U6709 (N_6709,N_5400,N_5890);
or U6710 (N_6710,N_5723,N_5412);
nor U6711 (N_6711,N_5007,N_5510);
or U6712 (N_6712,N_5599,N_5280);
or U6713 (N_6713,N_5295,N_5968);
and U6714 (N_6714,N_5329,N_5745);
or U6715 (N_6715,N_5167,N_5703);
and U6716 (N_6716,N_5202,N_5382);
and U6717 (N_6717,N_5205,N_5425);
and U6718 (N_6718,N_5585,N_5115);
and U6719 (N_6719,N_5362,N_5961);
and U6720 (N_6720,N_5108,N_5926);
or U6721 (N_6721,N_5588,N_5217);
or U6722 (N_6722,N_5868,N_5634);
nor U6723 (N_6723,N_5748,N_5034);
nand U6724 (N_6724,N_5861,N_5931);
xnor U6725 (N_6725,N_5055,N_5311);
nor U6726 (N_6726,N_5997,N_5271);
nand U6727 (N_6727,N_5033,N_5342);
or U6728 (N_6728,N_5315,N_5147);
xor U6729 (N_6729,N_5030,N_5514);
xnor U6730 (N_6730,N_5735,N_5329);
and U6731 (N_6731,N_5731,N_5741);
and U6732 (N_6732,N_5701,N_5525);
nand U6733 (N_6733,N_5741,N_5380);
and U6734 (N_6734,N_5060,N_5400);
nand U6735 (N_6735,N_5515,N_5664);
nand U6736 (N_6736,N_5140,N_5256);
nand U6737 (N_6737,N_5338,N_5485);
or U6738 (N_6738,N_5109,N_5769);
or U6739 (N_6739,N_5482,N_5168);
and U6740 (N_6740,N_5525,N_5442);
or U6741 (N_6741,N_5180,N_5186);
and U6742 (N_6742,N_5747,N_5585);
nor U6743 (N_6743,N_5730,N_5414);
or U6744 (N_6744,N_5904,N_5889);
nand U6745 (N_6745,N_5130,N_5861);
nand U6746 (N_6746,N_5830,N_5127);
or U6747 (N_6747,N_5264,N_5943);
xor U6748 (N_6748,N_5884,N_5499);
and U6749 (N_6749,N_5465,N_5325);
and U6750 (N_6750,N_5418,N_5054);
or U6751 (N_6751,N_5358,N_5725);
nand U6752 (N_6752,N_5262,N_5093);
nand U6753 (N_6753,N_5068,N_5498);
and U6754 (N_6754,N_5070,N_5485);
or U6755 (N_6755,N_5544,N_5698);
or U6756 (N_6756,N_5158,N_5804);
nor U6757 (N_6757,N_5354,N_5248);
nand U6758 (N_6758,N_5742,N_5913);
nor U6759 (N_6759,N_5914,N_5938);
xnor U6760 (N_6760,N_5122,N_5436);
or U6761 (N_6761,N_5037,N_5176);
nor U6762 (N_6762,N_5722,N_5780);
or U6763 (N_6763,N_5105,N_5917);
xor U6764 (N_6764,N_5621,N_5643);
nand U6765 (N_6765,N_5145,N_5287);
nand U6766 (N_6766,N_5886,N_5488);
or U6767 (N_6767,N_5144,N_5197);
nor U6768 (N_6768,N_5484,N_5667);
nor U6769 (N_6769,N_5010,N_5988);
and U6770 (N_6770,N_5609,N_5969);
and U6771 (N_6771,N_5321,N_5124);
nor U6772 (N_6772,N_5001,N_5768);
nand U6773 (N_6773,N_5058,N_5633);
nand U6774 (N_6774,N_5488,N_5687);
or U6775 (N_6775,N_5953,N_5305);
xnor U6776 (N_6776,N_5203,N_5236);
and U6777 (N_6777,N_5426,N_5805);
nor U6778 (N_6778,N_5563,N_5360);
nor U6779 (N_6779,N_5946,N_5793);
nand U6780 (N_6780,N_5660,N_5649);
nand U6781 (N_6781,N_5460,N_5865);
nor U6782 (N_6782,N_5253,N_5274);
nand U6783 (N_6783,N_5314,N_5790);
nor U6784 (N_6784,N_5216,N_5440);
nand U6785 (N_6785,N_5753,N_5631);
nand U6786 (N_6786,N_5697,N_5151);
and U6787 (N_6787,N_5957,N_5841);
nor U6788 (N_6788,N_5070,N_5127);
or U6789 (N_6789,N_5012,N_5387);
nand U6790 (N_6790,N_5936,N_5784);
nand U6791 (N_6791,N_5390,N_5031);
or U6792 (N_6792,N_5935,N_5790);
and U6793 (N_6793,N_5931,N_5556);
nor U6794 (N_6794,N_5168,N_5899);
nor U6795 (N_6795,N_5505,N_5804);
nor U6796 (N_6796,N_5799,N_5534);
nand U6797 (N_6797,N_5710,N_5612);
nand U6798 (N_6798,N_5193,N_5794);
and U6799 (N_6799,N_5367,N_5993);
nor U6800 (N_6800,N_5997,N_5496);
or U6801 (N_6801,N_5657,N_5580);
and U6802 (N_6802,N_5481,N_5033);
or U6803 (N_6803,N_5990,N_5907);
nand U6804 (N_6804,N_5155,N_5629);
xor U6805 (N_6805,N_5077,N_5103);
nor U6806 (N_6806,N_5965,N_5725);
and U6807 (N_6807,N_5055,N_5497);
or U6808 (N_6808,N_5700,N_5976);
nor U6809 (N_6809,N_5258,N_5203);
and U6810 (N_6810,N_5145,N_5599);
or U6811 (N_6811,N_5607,N_5485);
or U6812 (N_6812,N_5760,N_5402);
nor U6813 (N_6813,N_5050,N_5754);
nor U6814 (N_6814,N_5282,N_5979);
nand U6815 (N_6815,N_5951,N_5416);
and U6816 (N_6816,N_5921,N_5781);
nor U6817 (N_6817,N_5123,N_5412);
nand U6818 (N_6818,N_5069,N_5054);
and U6819 (N_6819,N_5924,N_5144);
nor U6820 (N_6820,N_5588,N_5540);
nor U6821 (N_6821,N_5808,N_5505);
or U6822 (N_6822,N_5981,N_5897);
nor U6823 (N_6823,N_5560,N_5946);
or U6824 (N_6824,N_5507,N_5177);
and U6825 (N_6825,N_5103,N_5224);
nand U6826 (N_6826,N_5499,N_5275);
or U6827 (N_6827,N_5854,N_5460);
nand U6828 (N_6828,N_5047,N_5988);
or U6829 (N_6829,N_5800,N_5831);
nand U6830 (N_6830,N_5379,N_5709);
or U6831 (N_6831,N_5203,N_5668);
and U6832 (N_6832,N_5988,N_5774);
xor U6833 (N_6833,N_5249,N_5146);
nor U6834 (N_6834,N_5775,N_5180);
nor U6835 (N_6835,N_5018,N_5740);
or U6836 (N_6836,N_5562,N_5186);
nand U6837 (N_6837,N_5153,N_5123);
nor U6838 (N_6838,N_5862,N_5222);
or U6839 (N_6839,N_5813,N_5466);
or U6840 (N_6840,N_5743,N_5085);
nand U6841 (N_6841,N_5159,N_5051);
and U6842 (N_6842,N_5368,N_5016);
nand U6843 (N_6843,N_5989,N_5002);
nor U6844 (N_6844,N_5708,N_5822);
and U6845 (N_6845,N_5023,N_5073);
nor U6846 (N_6846,N_5133,N_5287);
nand U6847 (N_6847,N_5389,N_5428);
and U6848 (N_6848,N_5629,N_5752);
and U6849 (N_6849,N_5463,N_5588);
nand U6850 (N_6850,N_5586,N_5833);
nor U6851 (N_6851,N_5387,N_5689);
or U6852 (N_6852,N_5483,N_5058);
or U6853 (N_6853,N_5687,N_5107);
nor U6854 (N_6854,N_5323,N_5926);
and U6855 (N_6855,N_5214,N_5089);
or U6856 (N_6856,N_5533,N_5236);
nand U6857 (N_6857,N_5106,N_5031);
nand U6858 (N_6858,N_5382,N_5578);
nor U6859 (N_6859,N_5313,N_5116);
and U6860 (N_6860,N_5572,N_5097);
and U6861 (N_6861,N_5213,N_5157);
and U6862 (N_6862,N_5985,N_5414);
nand U6863 (N_6863,N_5638,N_5520);
and U6864 (N_6864,N_5488,N_5402);
and U6865 (N_6865,N_5648,N_5253);
nand U6866 (N_6866,N_5794,N_5120);
nor U6867 (N_6867,N_5677,N_5821);
nand U6868 (N_6868,N_5949,N_5438);
nand U6869 (N_6869,N_5876,N_5487);
nand U6870 (N_6870,N_5798,N_5646);
and U6871 (N_6871,N_5713,N_5170);
xnor U6872 (N_6872,N_5707,N_5157);
and U6873 (N_6873,N_5008,N_5141);
or U6874 (N_6874,N_5127,N_5252);
and U6875 (N_6875,N_5742,N_5131);
nand U6876 (N_6876,N_5250,N_5652);
nand U6877 (N_6877,N_5690,N_5410);
nor U6878 (N_6878,N_5178,N_5361);
nor U6879 (N_6879,N_5570,N_5407);
and U6880 (N_6880,N_5059,N_5601);
nor U6881 (N_6881,N_5556,N_5647);
xor U6882 (N_6882,N_5998,N_5671);
or U6883 (N_6883,N_5914,N_5182);
or U6884 (N_6884,N_5421,N_5396);
and U6885 (N_6885,N_5801,N_5833);
nand U6886 (N_6886,N_5158,N_5751);
nand U6887 (N_6887,N_5487,N_5039);
nand U6888 (N_6888,N_5702,N_5495);
nand U6889 (N_6889,N_5804,N_5602);
nand U6890 (N_6890,N_5040,N_5001);
or U6891 (N_6891,N_5032,N_5764);
or U6892 (N_6892,N_5440,N_5877);
nor U6893 (N_6893,N_5689,N_5031);
nand U6894 (N_6894,N_5897,N_5139);
and U6895 (N_6895,N_5972,N_5325);
or U6896 (N_6896,N_5376,N_5042);
xor U6897 (N_6897,N_5613,N_5201);
or U6898 (N_6898,N_5486,N_5788);
and U6899 (N_6899,N_5914,N_5878);
or U6900 (N_6900,N_5406,N_5570);
or U6901 (N_6901,N_5309,N_5569);
and U6902 (N_6902,N_5371,N_5660);
nor U6903 (N_6903,N_5645,N_5277);
and U6904 (N_6904,N_5524,N_5929);
xor U6905 (N_6905,N_5148,N_5293);
or U6906 (N_6906,N_5527,N_5753);
xor U6907 (N_6907,N_5238,N_5792);
nand U6908 (N_6908,N_5914,N_5519);
nand U6909 (N_6909,N_5633,N_5834);
nor U6910 (N_6910,N_5351,N_5671);
nor U6911 (N_6911,N_5509,N_5867);
nand U6912 (N_6912,N_5410,N_5177);
xnor U6913 (N_6913,N_5208,N_5328);
or U6914 (N_6914,N_5201,N_5886);
or U6915 (N_6915,N_5877,N_5052);
nor U6916 (N_6916,N_5151,N_5691);
and U6917 (N_6917,N_5474,N_5442);
nand U6918 (N_6918,N_5161,N_5171);
nor U6919 (N_6919,N_5591,N_5533);
and U6920 (N_6920,N_5184,N_5345);
nor U6921 (N_6921,N_5755,N_5639);
xnor U6922 (N_6922,N_5414,N_5064);
or U6923 (N_6923,N_5277,N_5414);
xor U6924 (N_6924,N_5937,N_5804);
nand U6925 (N_6925,N_5656,N_5463);
and U6926 (N_6926,N_5686,N_5913);
or U6927 (N_6927,N_5053,N_5204);
or U6928 (N_6928,N_5867,N_5456);
and U6929 (N_6929,N_5858,N_5703);
and U6930 (N_6930,N_5205,N_5082);
nand U6931 (N_6931,N_5151,N_5885);
nor U6932 (N_6932,N_5570,N_5463);
nor U6933 (N_6933,N_5824,N_5723);
nor U6934 (N_6934,N_5852,N_5152);
nor U6935 (N_6935,N_5286,N_5999);
and U6936 (N_6936,N_5002,N_5474);
nand U6937 (N_6937,N_5475,N_5086);
nor U6938 (N_6938,N_5603,N_5348);
nor U6939 (N_6939,N_5398,N_5714);
nor U6940 (N_6940,N_5595,N_5691);
or U6941 (N_6941,N_5426,N_5214);
and U6942 (N_6942,N_5147,N_5023);
nor U6943 (N_6943,N_5755,N_5336);
and U6944 (N_6944,N_5366,N_5967);
and U6945 (N_6945,N_5943,N_5119);
or U6946 (N_6946,N_5799,N_5301);
nor U6947 (N_6947,N_5172,N_5897);
and U6948 (N_6948,N_5761,N_5645);
or U6949 (N_6949,N_5664,N_5132);
and U6950 (N_6950,N_5666,N_5806);
and U6951 (N_6951,N_5298,N_5907);
nor U6952 (N_6952,N_5395,N_5138);
nor U6953 (N_6953,N_5842,N_5323);
nor U6954 (N_6954,N_5637,N_5458);
or U6955 (N_6955,N_5477,N_5384);
or U6956 (N_6956,N_5609,N_5106);
nand U6957 (N_6957,N_5982,N_5237);
or U6958 (N_6958,N_5121,N_5345);
and U6959 (N_6959,N_5074,N_5842);
nand U6960 (N_6960,N_5794,N_5232);
and U6961 (N_6961,N_5604,N_5266);
xor U6962 (N_6962,N_5977,N_5644);
and U6963 (N_6963,N_5002,N_5917);
xor U6964 (N_6964,N_5272,N_5741);
and U6965 (N_6965,N_5629,N_5379);
nand U6966 (N_6966,N_5237,N_5416);
nor U6967 (N_6967,N_5616,N_5570);
or U6968 (N_6968,N_5657,N_5465);
or U6969 (N_6969,N_5472,N_5595);
and U6970 (N_6970,N_5403,N_5177);
nand U6971 (N_6971,N_5023,N_5706);
nor U6972 (N_6972,N_5464,N_5923);
or U6973 (N_6973,N_5770,N_5548);
nand U6974 (N_6974,N_5093,N_5265);
nand U6975 (N_6975,N_5330,N_5907);
nor U6976 (N_6976,N_5703,N_5394);
nand U6977 (N_6977,N_5043,N_5238);
nand U6978 (N_6978,N_5935,N_5983);
or U6979 (N_6979,N_5240,N_5230);
or U6980 (N_6980,N_5775,N_5736);
and U6981 (N_6981,N_5744,N_5632);
or U6982 (N_6982,N_5685,N_5181);
nand U6983 (N_6983,N_5395,N_5394);
or U6984 (N_6984,N_5208,N_5950);
nor U6985 (N_6985,N_5658,N_5682);
nand U6986 (N_6986,N_5645,N_5795);
or U6987 (N_6987,N_5997,N_5160);
nand U6988 (N_6988,N_5540,N_5340);
and U6989 (N_6989,N_5039,N_5948);
xnor U6990 (N_6990,N_5986,N_5928);
nor U6991 (N_6991,N_5929,N_5044);
nor U6992 (N_6992,N_5797,N_5355);
or U6993 (N_6993,N_5648,N_5058);
nor U6994 (N_6994,N_5019,N_5441);
and U6995 (N_6995,N_5636,N_5918);
and U6996 (N_6996,N_5611,N_5741);
nand U6997 (N_6997,N_5443,N_5478);
or U6998 (N_6998,N_5319,N_5202);
nor U6999 (N_6999,N_5167,N_5785);
nor U7000 (N_7000,N_6652,N_6417);
and U7001 (N_7001,N_6781,N_6901);
or U7002 (N_7002,N_6984,N_6041);
or U7003 (N_7003,N_6076,N_6713);
nand U7004 (N_7004,N_6599,N_6560);
nand U7005 (N_7005,N_6738,N_6936);
or U7006 (N_7006,N_6403,N_6411);
and U7007 (N_7007,N_6635,N_6211);
and U7008 (N_7008,N_6267,N_6844);
and U7009 (N_7009,N_6911,N_6078);
nor U7010 (N_7010,N_6780,N_6768);
or U7011 (N_7011,N_6261,N_6239);
and U7012 (N_7012,N_6064,N_6005);
or U7013 (N_7013,N_6576,N_6173);
or U7014 (N_7014,N_6703,N_6996);
nand U7015 (N_7015,N_6837,N_6312);
nor U7016 (N_7016,N_6235,N_6744);
nand U7017 (N_7017,N_6386,N_6721);
nor U7018 (N_7018,N_6546,N_6185);
and U7019 (N_7019,N_6096,N_6465);
nand U7020 (N_7020,N_6052,N_6718);
nand U7021 (N_7021,N_6704,N_6279);
nor U7022 (N_7022,N_6973,N_6583);
nor U7023 (N_7023,N_6522,N_6907);
nor U7024 (N_7024,N_6342,N_6841);
and U7025 (N_7025,N_6653,N_6506);
nor U7026 (N_7026,N_6071,N_6266);
xnor U7027 (N_7027,N_6799,N_6863);
and U7028 (N_7028,N_6087,N_6997);
and U7029 (N_7029,N_6253,N_6352);
nand U7030 (N_7030,N_6600,N_6004);
and U7031 (N_7031,N_6949,N_6036);
nand U7032 (N_7032,N_6413,N_6529);
nand U7033 (N_7033,N_6823,N_6150);
nor U7034 (N_7034,N_6124,N_6487);
nor U7035 (N_7035,N_6976,N_6785);
nand U7036 (N_7036,N_6451,N_6471);
nand U7037 (N_7037,N_6903,N_6545);
or U7038 (N_7038,N_6439,N_6942);
nand U7039 (N_7039,N_6251,N_6387);
or U7040 (N_7040,N_6783,N_6670);
and U7041 (N_7041,N_6460,N_6500);
or U7042 (N_7042,N_6532,N_6572);
nor U7043 (N_7043,N_6050,N_6526);
nand U7044 (N_7044,N_6601,N_6515);
nand U7045 (N_7045,N_6429,N_6832);
or U7046 (N_7046,N_6369,N_6330);
and U7047 (N_7047,N_6639,N_6126);
nor U7048 (N_7048,N_6569,N_6328);
or U7049 (N_7049,N_6158,N_6497);
xnor U7050 (N_7050,N_6750,N_6264);
nor U7051 (N_7051,N_6905,N_6656);
or U7052 (N_7052,N_6365,N_6385);
or U7053 (N_7053,N_6876,N_6646);
or U7054 (N_7054,N_6461,N_6118);
or U7055 (N_7055,N_6018,N_6691);
or U7056 (N_7056,N_6080,N_6383);
nand U7057 (N_7057,N_6134,N_6906);
xor U7058 (N_7058,N_6618,N_6673);
nand U7059 (N_7059,N_6496,N_6394);
or U7060 (N_7060,N_6516,N_6489);
nor U7061 (N_7061,N_6669,N_6100);
or U7062 (N_7062,N_6751,N_6433);
or U7063 (N_7063,N_6298,N_6986);
xnor U7064 (N_7064,N_6829,N_6504);
nand U7065 (N_7065,N_6000,N_6699);
xor U7066 (N_7066,N_6320,N_6553);
xor U7067 (N_7067,N_6313,N_6414);
nor U7068 (N_7068,N_6854,N_6067);
or U7069 (N_7069,N_6478,N_6148);
and U7070 (N_7070,N_6357,N_6376);
nand U7071 (N_7071,N_6399,N_6493);
nor U7072 (N_7072,N_6458,N_6082);
nor U7073 (N_7073,N_6775,N_6486);
nand U7074 (N_7074,N_6182,N_6727);
or U7075 (N_7075,N_6959,N_6645);
and U7076 (N_7076,N_6834,N_6390);
and U7077 (N_7077,N_6739,N_6175);
nand U7078 (N_7078,N_6530,N_6157);
nor U7079 (N_7079,N_6250,N_6366);
nand U7080 (N_7080,N_6445,N_6167);
xnor U7081 (N_7081,N_6620,N_6517);
nand U7082 (N_7082,N_6715,N_6069);
nand U7083 (N_7083,N_6737,N_6068);
or U7084 (N_7084,N_6058,N_6539);
xnor U7085 (N_7085,N_6866,N_6318);
and U7086 (N_7086,N_6482,N_6345);
or U7087 (N_7087,N_6634,N_6382);
or U7088 (N_7088,N_6722,N_6073);
nor U7089 (N_7089,N_6314,N_6109);
nand U7090 (N_7090,N_6305,N_6442);
or U7091 (N_7091,N_6547,N_6895);
and U7092 (N_7092,N_6197,N_6575);
xnor U7093 (N_7093,N_6501,N_6131);
nor U7094 (N_7094,N_6363,N_6117);
nand U7095 (N_7095,N_6725,N_6144);
nor U7096 (N_7096,N_6924,N_6355);
nand U7097 (N_7097,N_6128,N_6452);
xnor U7098 (N_7098,N_6025,N_6945);
nand U7099 (N_7099,N_6753,N_6955);
or U7100 (N_7100,N_6218,N_6360);
and U7101 (N_7101,N_6650,N_6479);
nand U7102 (N_7102,N_6825,N_6999);
xnor U7103 (N_7103,N_6663,N_6558);
or U7104 (N_7104,N_6215,N_6213);
and U7105 (N_7105,N_6473,N_6970);
or U7106 (N_7106,N_6858,N_6059);
or U7107 (N_7107,N_6440,N_6586);
and U7108 (N_7108,N_6711,N_6541);
nand U7109 (N_7109,N_6935,N_6544);
or U7110 (N_7110,N_6710,N_6095);
xor U7111 (N_7111,N_6946,N_6856);
nand U7112 (N_7112,N_6054,N_6728);
nor U7113 (N_7113,N_6820,N_6874);
nand U7114 (N_7114,N_6772,N_6523);
or U7115 (N_7115,N_6922,N_6824);
nor U7116 (N_7116,N_6633,N_6003);
and U7117 (N_7117,N_6706,N_6099);
and U7118 (N_7118,N_6591,N_6480);
and U7119 (N_7119,N_6717,N_6662);
or U7120 (N_7120,N_6286,N_6685);
nand U7121 (N_7121,N_6241,N_6975);
xor U7122 (N_7122,N_6759,N_6938);
and U7123 (N_7123,N_6154,N_6643);
and U7124 (N_7124,N_6757,N_6971);
nor U7125 (N_7125,N_6426,N_6072);
nor U7126 (N_7126,N_6106,N_6503);
xor U7127 (N_7127,N_6288,N_6779);
or U7128 (N_7128,N_6990,N_6720);
nand U7129 (N_7129,N_6612,N_6980);
nor U7130 (N_7130,N_6246,N_6038);
and U7131 (N_7131,N_6393,N_6991);
nand U7132 (N_7132,N_6092,N_6227);
nand U7133 (N_7133,N_6192,N_6778);
or U7134 (N_7134,N_6133,N_6269);
nand U7135 (N_7135,N_6336,N_6333);
nand U7136 (N_7136,N_6848,N_6375);
nor U7137 (N_7137,N_6556,N_6577);
nor U7138 (N_7138,N_6915,N_6033);
or U7139 (N_7139,N_6398,N_6467);
or U7140 (N_7140,N_6459,N_6654);
nor U7141 (N_7141,N_6629,N_6542);
nand U7142 (N_7142,N_6939,N_6693);
and U7143 (N_7143,N_6047,N_6354);
xor U7144 (N_7144,N_6581,N_6761);
or U7145 (N_7145,N_6512,N_6450);
nor U7146 (N_7146,N_6243,N_6389);
nand U7147 (N_7147,N_6189,N_6667);
nor U7148 (N_7148,N_6859,N_6130);
and U7149 (N_7149,N_6093,N_6332);
nand U7150 (N_7150,N_6794,N_6217);
nor U7151 (N_7151,N_6819,N_6969);
nor U7152 (N_7152,N_6448,N_6037);
or U7153 (N_7153,N_6831,N_6540);
xor U7154 (N_7154,N_6344,N_6659);
nand U7155 (N_7155,N_6381,N_6712);
nor U7156 (N_7156,N_6488,N_6733);
nor U7157 (N_7157,N_6747,N_6514);
or U7158 (N_7158,N_6034,N_6579);
nand U7159 (N_7159,N_6896,N_6680);
and U7160 (N_7160,N_6214,N_6878);
or U7161 (N_7161,N_6568,N_6867);
nand U7162 (N_7162,N_6176,N_6690);
nand U7163 (N_7163,N_6110,N_6210);
nor U7164 (N_7164,N_6937,N_6104);
xnor U7165 (N_7165,N_6983,N_6362);
and U7166 (N_7166,N_6260,N_6828);
nand U7167 (N_7167,N_6807,N_6965);
and U7168 (N_7168,N_6309,N_6637);
or U7169 (N_7169,N_6605,N_6584);
and U7170 (N_7170,N_6833,N_6315);
and U7171 (N_7171,N_6022,N_6055);
nand U7172 (N_7172,N_6368,N_6338);
and U7173 (N_7173,N_6276,N_6894);
nor U7174 (N_7174,N_6017,N_6035);
nand U7175 (N_7175,N_6233,N_6339);
and U7176 (N_7176,N_6364,N_6709);
and U7177 (N_7177,N_6578,N_6244);
nand U7178 (N_7178,N_6190,N_6630);
xnor U7179 (N_7179,N_6769,N_6608);
nor U7180 (N_7180,N_6358,N_6206);
nand U7181 (N_7181,N_6498,N_6257);
or U7182 (N_7182,N_6049,N_6655);
or U7183 (N_7183,N_6060,N_6884);
nor U7184 (N_7184,N_6468,N_6573);
nand U7185 (N_7185,N_6282,N_6446);
nand U7186 (N_7186,N_6648,N_6081);
or U7187 (N_7187,N_6934,N_6262);
and U7188 (N_7188,N_6111,N_6145);
and U7189 (N_7189,N_6495,N_6208);
nand U7190 (N_7190,N_6283,N_6258);
nor U7191 (N_7191,N_6843,N_6582);
or U7192 (N_7192,N_6377,N_6762);
nand U7193 (N_7193,N_6928,N_6774);
nand U7194 (N_7194,N_6388,N_6948);
nand U7195 (N_7195,N_6873,N_6585);
and U7196 (N_7196,N_6507,N_6030);
and U7197 (N_7197,N_6765,N_6888);
nand U7198 (N_7198,N_6287,N_6085);
nor U7199 (N_7199,N_6510,N_6566);
and U7200 (N_7200,N_6617,N_6324);
nor U7201 (N_7201,N_6658,N_6773);
nor U7202 (N_7202,N_6379,N_6252);
or U7203 (N_7203,N_6861,N_6743);
nor U7204 (N_7204,N_6056,N_6201);
and U7205 (N_7205,N_6550,N_6155);
nand U7206 (N_7206,N_6527,N_6303);
nor U7207 (N_7207,N_6914,N_6864);
and U7208 (N_7208,N_6805,N_6631);
nand U7209 (N_7209,N_6020,N_6533);
or U7210 (N_7210,N_6679,N_6995);
or U7211 (N_7211,N_6668,N_6340);
nor U7212 (N_7212,N_6474,N_6229);
xnor U7213 (N_7213,N_6660,N_6453);
xnor U7214 (N_7214,N_6490,N_6319);
or U7215 (N_7215,N_6869,N_6163);
nor U7216 (N_7216,N_6200,N_6125);
and U7217 (N_7217,N_6694,N_6323);
or U7218 (N_7218,N_6846,N_6808);
and U7219 (N_7219,N_6817,N_6065);
and U7220 (N_7220,N_6664,N_6224);
nor U7221 (N_7221,N_6135,N_6477);
nor U7222 (N_7222,N_6108,N_6361);
xnor U7223 (N_7223,N_6793,N_6367);
and U7224 (N_7224,N_6528,N_6821);
xor U7225 (N_7225,N_6875,N_6010);
or U7226 (N_7226,N_6800,N_6304);
nand U7227 (N_7227,N_6053,N_6031);
nor U7228 (N_7228,N_6950,N_6812);
nor U7229 (N_7229,N_6961,N_6008);
nor U7230 (N_7230,N_6032,N_6316);
and U7231 (N_7231,N_6137,N_6787);
nand U7232 (N_7232,N_6610,N_6933);
and U7233 (N_7233,N_6505,N_6089);
and U7234 (N_7234,N_6188,N_6177);
or U7235 (N_7235,N_6920,N_6966);
nand U7236 (N_7236,N_6732,N_6062);
nor U7237 (N_7237,N_6968,N_6682);
and U7238 (N_7238,N_6293,N_6771);
xor U7239 (N_7239,N_6166,N_6026);
or U7240 (N_7240,N_6770,N_6044);
and U7241 (N_7241,N_6788,N_6116);
or U7242 (N_7242,N_6149,N_6327);
nor U7243 (N_7243,N_6202,N_6007);
nor U7244 (N_7244,N_6492,N_6066);
nand U7245 (N_7245,N_6219,N_6756);
or U7246 (N_7246,N_6941,N_6730);
nor U7247 (N_7247,N_6359,N_6695);
and U7248 (N_7248,N_6535,N_6334);
nand U7249 (N_7249,N_6816,N_6248);
nand U7250 (N_7250,N_6625,N_6310);
or U7251 (N_7251,N_6964,N_6434);
or U7252 (N_7252,N_6886,N_6736);
xnor U7253 (N_7253,N_6294,N_6119);
and U7254 (N_7254,N_6122,N_6892);
and U7255 (N_7255,N_6697,N_6839);
and U7256 (N_7256,N_6230,N_6749);
or U7257 (N_7257,N_6755,N_6272);
nand U7258 (N_7258,N_6838,N_6792);
nand U7259 (N_7259,N_6475,N_6666);
or U7260 (N_7260,N_6724,N_6300);
or U7261 (N_7261,N_6212,N_6207);
and U7262 (N_7262,N_6129,N_6347);
nand U7263 (N_7263,N_6814,N_6604);
and U7264 (N_7264,N_6183,N_6661);
nor U7265 (N_7265,N_6107,N_6204);
nand U7266 (N_7266,N_6019,N_6603);
nand U7267 (N_7267,N_6223,N_6337);
xnor U7268 (N_7268,N_6299,N_6373);
or U7269 (N_7269,N_6596,N_6297);
nor U7270 (N_7270,N_6256,N_6904);
nor U7271 (N_7271,N_6979,N_6407);
and U7272 (N_7272,N_6021,N_6548);
xnor U7273 (N_7273,N_6317,N_6589);
nand U7274 (N_7274,N_6987,N_6142);
nand U7275 (N_7275,N_6193,N_6882);
xor U7276 (N_7276,N_6335,N_6513);
nand U7277 (N_7277,N_6090,N_6370);
xnor U7278 (N_7278,N_6236,N_6992);
and U7279 (N_7279,N_6430,N_6077);
nor U7280 (N_7280,N_6619,N_6952);
or U7281 (N_7281,N_6804,N_6380);
nand U7282 (N_7282,N_6857,N_6395);
and U7283 (N_7283,N_6259,N_6567);
nand U7284 (N_7284,N_6196,N_6621);
nand U7285 (N_7285,N_6242,N_6571);
nand U7286 (N_7286,N_6203,N_6143);
or U7287 (N_7287,N_6245,N_6156);
nor U7288 (N_7288,N_6416,N_6168);
or U7289 (N_7289,N_6632,N_6280);
or U7290 (N_7290,N_6674,N_6371);
nor U7291 (N_7291,N_6470,N_6404);
nor U7292 (N_7292,N_6348,N_6301);
and U7293 (N_7293,N_6758,N_6097);
nand U7294 (N_7294,N_6726,N_6891);
and U7295 (N_7295,N_6870,N_6963);
nor U7296 (N_7296,N_6723,N_6902);
and U7297 (N_7297,N_6187,N_6165);
or U7298 (N_7298,N_6701,N_6782);
nor U7299 (N_7299,N_6321,N_6102);
nand U7300 (N_7300,N_6484,N_6275);
or U7301 (N_7301,N_6748,N_6642);
xnor U7302 (N_7302,N_6161,N_6588);
nor U7303 (N_7303,N_6784,N_6678);
or U7304 (N_7304,N_6651,N_6349);
nor U7305 (N_7305,N_6178,N_6469);
and U7306 (N_7306,N_6538,N_6466);
nor U7307 (N_7307,N_6595,N_6626);
and U7308 (N_7308,N_6565,N_6850);
xnor U7309 (N_7309,N_6016,N_6221);
nand U7310 (N_7310,N_6836,N_6692);
and U7311 (N_7311,N_6326,N_6464);
or U7312 (N_7312,N_6993,N_6960);
nor U7313 (N_7313,N_6754,N_6557);
nand U7314 (N_7314,N_6198,N_6141);
nand U7315 (N_7315,N_6594,N_6628);
nor U7316 (N_7316,N_6046,N_6291);
or U7317 (N_7317,N_6638,N_6735);
nand U7318 (N_7318,N_6974,N_6931);
and U7319 (N_7319,N_6890,N_6872);
nand U7320 (N_7320,N_6397,N_6428);
or U7321 (N_7321,N_6534,N_6574);
nand U7322 (N_7322,N_6249,N_6006);
or U7323 (N_7323,N_6402,N_6222);
and U7324 (N_7324,N_6688,N_6270);
and U7325 (N_7325,N_6423,N_6714);
and U7326 (N_7326,N_6234,N_6597);
nand U7327 (N_7327,N_6418,N_6278);
nor U7328 (N_7328,N_6013,N_6444);
nand U7329 (N_7329,N_6855,N_6432);
nand U7330 (N_7330,N_6623,N_6520);
or U7331 (N_7331,N_6921,N_6481);
or U7332 (N_7332,N_6883,N_6263);
or U7333 (N_7333,N_6994,N_6563);
nor U7334 (N_7334,N_6958,N_6048);
nand U7335 (N_7335,N_6273,N_6818);
nand U7336 (N_7336,N_6255,N_6042);
and U7337 (N_7337,N_6123,N_6494);
or U7338 (N_7338,N_6554,N_6412);
xnor U7339 (N_7339,N_6845,N_6179);
xnor U7340 (N_7340,N_6985,N_6307);
or U7341 (N_7341,N_6622,N_6978);
nor U7342 (N_7342,N_6777,N_6091);
nand U7343 (N_7343,N_6981,N_6681);
nand U7344 (N_7344,N_6502,N_6609);
or U7345 (N_7345,N_6796,N_6372);
nand U7346 (N_7346,N_6811,N_6640);
xnor U7347 (N_7347,N_6893,N_6741);
nor U7348 (N_7348,N_6088,N_6014);
or U7349 (N_7349,N_6598,N_6562);
and U7350 (N_7350,N_6075,N_6051);
and U7351 (N_7351,N_6815,N_6734);
and U7352 (N_7352,N_6209,N_6422);
and U7353 (N_7353,N_6665,N_6083);
nor U7354 (N_7354,N_6265,N_6687);
xnor U7355 (N_7355,N_6405,N_6136);
nor U7356 (N_7356,N_6602,N_6731);
or U7357 (N_7357,N_6636,N_6940);
or U7358 (N_7358,N_6677,N_6519);
nor U7359 (N_7359,N_6039,N_6181);
or U7360 (N_7360,N_6400,N_6801);
and U7361 (N_7361,N_6476,N_6392);
nor U7362 (N_7362,N_6180,N_6454);
or U7363 (N_7363,N_6308,N_6790);
nor U7364 (N_7364,N_6061,N_6764);
xnor U7365 (N_7365,N_6644,N_6592);
nand U7366 (N_7366,N_6795,N_6977);
nor U7367 (N_7367,N_6898,N_6094);
xnor U7368 (N_7368,N_6611,N_6485);
nor U7369 (N_7369,N_6237,N_6555);
or U7370 (N_7370,N_6729,N_6170);
xor U7371 (N_7371,N_6740,N_6536);
or U7372 (N_7372,N_6913,N_6015);
nand U7373 (N_7373,N_6951,N_6849);
or U7374 (N_7374,N_6009,N_6707);
nor U7375 (N_7375,N_6254,N_6284);
nor U7376 (N_7376,N_6027,N_6549);
nor U7377 (N_7377,N_6274,N_6767);
xor U7378 (N_7378,N_6391,N_6868);
and U7379 (N_7379,N_6409,N_6908);
nand U7380 (N_7380,N_6871,N_6716);
xnor U7381 (N_7381,N_6164,N_6115);
or U7382 (N_7382,N_6689,N_6835);
or U7383 (N_7383,N_6881,N_6760);
or U7384 (N_7384,N_6879,N_6923);
or U7385 (N_7385,N_6809,N_6865);
nor U7386 (N_7386,N_6172,N_6063);
or U7387 (N_7387,N_6810,N_6561);
or U7388 (N_7388,N_6043,N_6509);
nand U7389 (N_7389,N_6463,N_6943);
nand U7390 (N_7390,N_6281,N_6910);
or U7391 (N_7391,N_6146,N_6708);
xnor U7392 (N_7392,N_6847,N_6607);
and U7393 (N_7393,N_6401,N_6989);
or U7394 (N_7394,N_6803,N_6045);
nand U7395 (N_7395,N_6916,N_6700);
nor U7396 (N_7396,N_6472,N_6427);
or U7397 (N_7397,N_6606,N_6786);
nor U7398 (N_7398,N_6216,N_6559);
nor U7399 (N_7399,N_6240,N_6954);
and U7400 (N_7400,N_6415,N_6613);
or U7401 (N_7401,N_6551,N_6001);
or U7402 (N_7402,N_6296,N_6184);
and U7403 (N_7403,N_6086,N_6079);
and U7404 (N_7404,N_6311,N_6152);
xnor U7405 (N_7405,N_6830,N_6351);
and U7406 (N_7406,N_6587,N_6114);
or U7407 (N_7407,N_6331,N_6462);
or U7408 (N_7408,N_6295,N_6424);
xnor U7409 (N_7409,N_6531,N_6615);
and U7410 (N_7410,N_6231,N_6499);
nor U7411 (N_7411,N_6437,N_6268);
and U7412 (N_7412,N_6683,N_6797);
nand U7413 (N_7413,N_6671,N_6926);
nor U7414 (N_7414,N_6491,N_6153);
and U7415 (N_7415,N_6441,N_6447);
nor U7416 (N_7416,N_6057,N_6012);
nor U7417 (N_7417,N_6378,N_6228);
xor U7418 (N_7418,N_6002,N_6356);
nand U7419 (N_7419,N_6616,N_6806);
nand U7420 (N_7420,N_6912,N_6151);
and U7421 (N_7421,N_6084,N_6160);
xor U7422 (N_7422,N_6169,N_6552);
xor U7423 (N_7423,N_6277,N_6862);
and U7424 (N_7424,N_6396,N_6802);
or U7425 (N_7425,N_6853,N_6647);
nor U7426 (N_7426,N_6346,N_6238);
nor U7427 (N_7427,N_6826,N_6247);
xor U7428 (N_7428,N_6947,N_6029);
nor U7429 (N_7429,N_6763,N_6988);
nor U7430 (N_7430,N_6457,N_6614);
or U7431 (N_7431,N_6408,N_6719);
or U7432 (N_7432,N_6852,N_6840);
and U7433 (N_7433,N_6953,N_6776);
or U7434 (N_7434,N_6483,N_6887);
xnor U7435 (N_7435,N_6885,N_6860);
or U7436 (N_7436,N_6120,N_6162);
and U7437 (N_7437,N_6851,N_6420);
or U7438 (N_7438,N_6580,N_6742);
and U7439 (N_7439,N_6350,N_6325);
and U7440 (N_7440,N_6220,N_6406);
or U7441 (N_7441,N_6232,N_6702);
and U7442 (N_7442,N_6105,N_6525);
and U7443 (N_7443,N_6624,N_6956);
nand U7444 (N_7444,N_6127,N_6113);
or U7445 (N_7445,N_6132,N_6880);
or U7446 (N_7446,N_6746,N_6570);
nor U7447 (N_7447,N_6302,N_6998);
nor U7448 (N_7448,N_6900,N_6186);
and U7449 (N_7449,N_6174,N_6925);
or U7450 (N_7450,N_6112,N_6419);
nand U7451 (N_7451,N_6842,N_6384);
or U7452 (N_7452,N_6827,N_6967);
nor U7453 (N_7453,N_6023,N_6341);
nor U7454 (N_7454,N_6139,N_6138);
and U7455 (N_7455,N_6909,N_6813);
nand U7456 (N_7456,N_6225,N_6147);
or U7457 (N_7457,N_6011,N_6897);
or U7458 (N_7458,N_6929,N_6918);
and U7459 (N_7459,N_6199,N_6766);
nand U7460 (N_7460,N_6537,N_6329);
nand U7461 (N_7461,N_6285,N_6657);
nand U7462 (N_7462,N_6028,N_6449);
nor U7463 (N_7463,N_6289,N_6438);
and U7464 (N_7464,N_6957,N_6074);
nor U7465 (N_7465,N_6518,N_6972);
and U7466 (N_7466,N_6226,N_6421);
or U7467 (N_7467,N_6789,N_6930);
and U7468 (N_7468,N_6752,N_6455);
or U7469 (N_7469,N_6944,N_6962);
and U7470 (N_7470,N_6684,N_6171);
or U7471 (N_7471,N_6698,N_6374);
nor U7472 (N_7472,N_6343,N_6521);
and U7473 (N_7473,N_6040,N_6676);
nand U7474 (N_7474,N_6098,N_6410);
nor U7475 (N_7475,N_6435,N_6205);
nand U7476 (N_7476,N_6436,N_6641);
nor U7477 (N_7477,N_6899,N_6191);
nor U7478 (N_7478,N_6696,N_6791);
nand U7479 (N_7479,N_6070,N_6443);
and U7480 (N_7480,N_6194,N_6798);
or U7481 (N_7481,N_6917,N_6431);
xnor U7482 (N_7482,N_6121,N_6140);
or U7483 (N_7483,N_6705,N_6675);
and U7484 (N_7484,N_6590,N_6543);
or U7485 (N_7485,N_6508,N_6456);
nor U7486 (N_7486,N_6524,N_6024);
nor U7487 (N_7487,N_6627,N_6195);
or U7488 (N_7488,N_6101,N_6877);
nand U7489 (N_7489,N_6686,N_6564);
or U7490 (N_7490,N_6822,N_6322);
nand U7491 (N_7491,N_6927,N_6982);
nor U7492 (N_7492,N_6672,N_6511);
nand U7493 (N_7493,N_6306,N_6932);
nand U7494 (N_7494,N_6889,N_6103);
nand U7495 (N_7495,N_6353,N_6745);
nor U7496 (N_7496,N_6919,N_6159);
and U7497 (N_7497,N_6290,N_6649);
nor U7498 (N_7498,N_6292,N_6593);
nor U7499 (N_7499,N_6425,N_6271);
or U7500 (N_7500,N_6174,N_6307);
or U7501 (N_7501,N_6743,N_6900);
or U7502 (N_7502,N_6688,N_6392);
nor U7503 (N_7503,N_6888,N_6240);
nand U7504 (N_7504,N_6356,N_6560);
xor U7505 (N_7505,N_6864,N_6835);
and U7506 (N_7506,N_6853,N_6224);
nor U7507 (N_7507,N_6721,N_6115);
xnor U7508 (N_7508,N_6549,N_6075);
or U7509 (N_7509,N_6640,N_6190);
nor U7510 (N_7510,N_6610,N_6030);
nand U7511 (N_7511,N_6710,N_6270);
or U7512 (N_7512,N_6539,N_6217);
and U7513 (N_7513,N_6506,N_6500);
xor U7514 (N_7514,N_6976,N_6873);
and U7515 (N_7515,N_6460,N_6904);
nor U7516 (N_7516,N_6597,N_6706);
and U7517 (N_7517,N_6700,N_6084);
xor U7518 (N_7518,N_6229,N_6647);
xor U7519 (N_7519,N_6897,N_6099);
nand U7520 (N_7520,N_6592,N_6447);
nor U7521 (N_7521,N_6456,N_6578);
nand U7522 (N_7522,N_6911,N_6616);
or U7523 (N_7523,N_6435,N_6243);
and U7524 (N_7524,N_6277,N_6834);
nand U7525 (N_7525,N_6161,N_6511);
nor U7526 (N_7526,N_6532,N_6443);
nor U7527 (N_7527,N_6613,N_6167);
or U7528 (N_7528,N_6136,N_6667);
xor U7529 (N_7529,N_6077,N_6084);
nor U7530 (N_7530,N_6968,N_6907);
and U7531 (N_7531,N_6729,N_6882);
xnor U7532 (N_7532,N_6331,N_6639);
nor U7533 (N_7533,N_6360,N_6859);
and U7534 (N_7534,N_6750,N_6935);
or U7535 (N_7535,N_6025,N_6774);
or U7536 (N_7536,N_6928,N_6944);
nand U7537 (N_7537,N_6508,N_6273);
and U7538 (N_7538,N_6222,N_6484);
nand U7539 (N_7539,N_6152,N_6381);
nor U7540 (N_7540,N_6032,N_6386);
and U7541 (N_7541,N_6161,N_6399);
nor U7542 (N_7542,N_6505,N_6044);
nand U7543 (N_7543,N_6317,N_6488);
or U7544 (N_7544,N_6496,N_6123);
or U7545 (N_7545,N_6560,N_6981);
or U7546 (N_7546,N_6920,N_6460);
and U7547 (N_7547,N_6157,N_6930);
and U7548 (N_7548,N_6088,N_6104);
or U7549 (N_7549,N_6655,N_6209);
and U7550 (N_7550,N_6996,N_6722);
nand U7551 (N_7551,N_6799,N_6655);
or U7552 (N_7552,N_6253,N_6930);
and U7553 (N_7553,N_6033,N_6276);
nor U7554 (N_7554,N_6798,N_6839);
and U7555 (N_7555,N_6019,N_6582);
nand U7556 (N_7556,N_6524,N_6341);
nor U7557 (N_7557,N_6400,N_6943);
nand U7558 (N_7558,N_6825,N_6485);
nor U7559 (N_7559,N_6054,N_6193);
nor U7560 (N_7560,N_6287,N_6503);
and U7561 (N_7561,N_6078,N_6353);
nor U7562 (N_7562,N_6863,N_6735);
nand U7563 (N_7563,N_6490,N_6932);
and U7564 (N_7564,N_6915,N_6532);
nand U7565 (N_7565,N_6201,N_6549);
and U7566 (N_7566,N_6138,N_6500);
or U7567 (N_7567,N_6210,N_6018);
or U7568 (N_7568,N_6719,N_6940);
or U7569 (N_7569,N_6034,N_6969);
and U7570 (N_7570,N_6015,N_6589);
or U7571 (N_7571,N_6304,N_6793);
and U7572 (N_7572,N_6755,N_6349);
nand U7573 (N_7573,N_6851,N_6239);
nor U7574 (N_7574,N_6647,N_6924);
nand U7575 (N_7575,N_6800,N_6145);
nor U7576 (N_7576,N_6581,N_6697);
and U7577 (N_7577,N_6781,N_6080);
nor U7578 (N_7578,N_6559,N_6467);
nor U7579 (N_7579,N_6706,N_6196);
xor U7580 (N_7580,N_6332,N_6890);
nor U7581 (N_7581,N_6126,N_6629);
nor U7582 (N_7582,N_6735,N_6092);
and U7583 (N_7583,N_6608,N_6549);
or U7584 (N_7584,N_6895,N_6562);
nand U7585 (N_7585,N_6102,N_6682);
nor U7586 (N_7586,N_6176,N_6234);
or U7587 (N_7587,N_6748,N_6769);
nand U7588 (N_7588,N_6119,N_6616);
or U7589 (N_7589,N_6351,N_6757);
nand U7590 (N_7590,N_6510,N_6693);
and U7591 (N_7591,N_6586,N_6836);
nand U7592 (N_7592,N_6212,N_6831);
or U7593 (N_7593,N_6453,N_6008);
or U7594 (N_7594,N_6261,N_6976);
or U7595 (N_7595,N_6123,N_6828);
nor U7596 (N_7596,N_6547,N_6495);
nor U7597 (N_7597,N_6189,N_6096);
xor U7598 (N_7598,N_6327,N_6123);
or U7599 (N_7599,N_6401,N_6631);
or U7600 (N_7600,N_6305,N_6791);
nor U7601 (N_7601,N_6677,N_6359);
and U7602 (N_7602,N_6256,N_6678);
xnor U7603 (N_7603,N_6417,N_6460);
nor U7604 (N_7604,N_6826,N_6804);
xor U7605 (N_7605,N_6636,N_6770);
nor U7606 (N_7606,N_6790,N_6515);
or U7607 (N_7607,N_6513,N_6730);
nand U7608 (N_7608,N_6559,N_6502);
and U7609 (N_7609,N_6071,N_6440);
nand U7610 (N_7610,N_6220,N_6753);
and U7611 (N_7611,N_6141,N_6818);
and U7612 (N_7612,N_6166,N_6959);
or U7613 (N_7613,N_6459,N_6477);
xor U7614 (N_7614,N_6604,N_6571);
nor U7615 (N_7615,N_6789,N_6476);
nor U7616 (N_7616,N_6654,N_6139);
or U7617 (N_7617,N_6728,N_6015);
nor U7618 (N_7618,N_6474,N_6645);
nor U7619 (N_7619,N_6439,N_6613);
or U7620 (N_7620,N_6634,N_6331);
xor U7621 (N_7621,N_6643,N_6786);
nor U7622 (N_7622,N_6666,N_6448);
nand U7623 (N_7623,N_6560,N_6069);
or U7624 (N_7624,N_6448,N_6510);
and U7625 (N_7625,N_6244,N_6155);
nand U7626 (N_7626,N_6926,N_6186);
nand U7627 (N_7627,N_6852,N_6766);
and U7628 (N_7628,N_6189,N_6611);
nand U7629 (N_7629,N_6758,N_6545);
xor U7630 (N_7630,N_6858,N_6077);
nor U7631 (N_7631,N_6188,N_6226);
or U7632 (N_7632,N_6251,N_6613);
xor U7633 (N_7633,N_6221,N_6787);
nand U7634 (N_7634,N_6108,N_6914);
and U7635 (N_7635,N_6590,N_6467);
and U7636 (N_7636,N_6641,N_6084);
nand U7637 (N_7637,N_6780,N_6486);
xor U7638 (N_7638,N_6856,N_6027);
or U7639 (N_7639,N_6525,N_6001);
or U7640 (N_7640,N_6612,N_6445);
nand U7641 (N_7641,N_6807,N_6244);
and U7642 (N_7642,N_6064,N_6008);
or U7643 (N_7643,N_6379,N_6160);
xor U7644 (N_7644,N_6133,N_6652);
and U7645 (N_7645,N_6346,N_6040);
nand U7646 (N_7646,N_6591,N_6103);
xnor U7647 (N_7647,N_6942,N_6472);
nand U7648 (N_7648,N_6854,N_6781);
or U7649 (N_7649,N_6347,N_6122);
and U7650 (N_7650,N_6825,N_6867);
or U7651 (N_7651,N_6727,N_6173);
nand U7652 (N_7652,N_6698,N_6426);
and U7653 (N_7653,N_6223,N_6620);
xor U7654 (N_7654,N_6224,N_6815);
or U7655 (N_7655,N_6049,N_6740);
or U7656 (N_7656,N_6440,N_6181);
and U7657 (N_7657,N_6120,N_6294);
nand U7658 (N_7658,N_6109,N_6106);
xnor U7659 (N_7659,N_6514,N_6768);
and U7660 (N_7660,N_6577,N_6371);
or U7661 (N_7661,N_6962,N_6091);
nand U7662 (N_7662,N_6955,N_6244);
and U7663 (N_7663,N_6497,N_6003);
nor U7664 (N_7664,N_6157,N_6024);
nand U7665 (N_7665,N_6441,N_6304);
or U7666 (N_7666,N_6455,N_6775);
and U7667 (N_7667,N_6872,N_6653);
or U7668 (N_7668,N_6024,N_6245);
nor U7669 (N_7669,N_6229,N_6127);
and U7670 (N_7670,N_6362,N_6894);
nor U7671 (N_7671,N_6614,N_6191);
nand U7672 (N_7672,N_6126,N_6163);
nand U7673 (N_7673,N_6446,N_6674);
and U7674 (N_7674,N_6180,N_6874);
or U7675 (N_7675,N_6105,N_6799);
nor U7676 (N_7676,N_6970,N_6508);
nor U7677 (N_7677,N_6319,N_6444);
nor U7678 (N_7678,N_6566,N_6097);
nor U7679 (N_7679,N_6842,N_6164);
nand U7680 (N_7680,N_6806,N_6329);
nand U7681 (N_7681,N_6324,N_6044);
or U7682 (N_7682,N_6680,N_6173);
nand U7683 (N_7683,N_6075,N_6039);
and U7684 (N_7684,N_6766,N_6848);
or U7685 (N_7685,N_6203,N_6735);
nand U7686 (N_7686,N_6467,N_6509);
or U7687 (N_7687,N_6500,N_6793);
and U7688 (N_7688,N_6707,N_6794);
or U7689 (N_7689,N_6577,N_6883);
nand U7690 (N_7690,N_6666,N_6446);
or U7691 (N_7691,N_6217,N_6563);
nand U7692 (N_7692,N_6624,N_6211);
nand U7693 (N_7693,N_6485,N_6324);
or U7694 (N_7694,N_6068,N_6656);
and U7695 (N_7695,N_6758,N_6973);
nor U7696 (N_7696,N_6943,N_6254);
and U7697 (N_7697,N_6636,N_6130);
xnor U7698 (N_7698,N_6433,N_6361);
and U7699 (N_7699,N_6464,N_6764);
and U7700 (N_7700,N_6362,N_6554);
or U7701 (N_7701,N_6110,N_6102);
nand U7702 (N_7702,N_6243,N_6544);
or U7703 (N_7703,N_6901,N_6358);
nor U7704 (N_7704,N_6577,N_6422);
and U7705 (N_7705,N_6349,N_6774);
and U7706 (N_7706,N_6189,N_6923);
or U7707 (N_7707,N_6110,N_6903);
nor U7708 (N_7708,N_6947,N_6724);
xnor U7709 (N_7709,N_6302,N_6352);
and U7710 (N_7710,N_6866,N_6303);
and U7711 (N_7711,N_6653,N_6369);
or U7712 (N_7712,N_6959,N_6888);
nand U7713 (N_7713,N_6644,N_6456);
or U7714 (N_7714,N_6134,N_6734);
xnor U7715 (N_7715,N_6962,N_6371);
or U7716 (N_7716,N_6523,N_6055);
and U7717 (N_7717,N_6798,N_6819);
nand U7718 (N_7718,N_6197,N_6967);
and U7719 (N_7719,N_6367,N_6741);
or U7720 (N_7720,N_6490,N_6083);
and U7721 (N_7721,N_6542,N_6345);
and U7722 (N_7722,N_6488,N_6853);
nand U7723 (N_7723,N_6360,N_6619);
or U7724 (N_7724,N_6810,N_6979);
or U7725 (N_7725,N_6439,N_6135);
or U7726 (N_7726,N_6283,N_6189);
and U7727 (N_7727,N_6506,N_6634);
nor U7728 (N_7728,N_6619,N_6486);
nand U7729 (N_7729,N_6331,N_6759);
and U7730 (N_7730,N_6874,N_6655);
nand U7731 (N_7731,N_6383,N_6573);
nand U7732 (N_7732,N_6370,N_6212);
nand U7733 (N_7733,N_6646,N_6544);
nor U7734 (N_7734,N_6415,N_6059);
nand U7735 (N_7735,N_6432,N_6898);
or U7736 (N_7736,N_6302,N_6508);
nand U7737 (N_7737,N_6155,N_6307);
nor U7738 (N_7738,N_6414,N_6381);
or U7739 (N_7739,N_6770,N_6465);
or U7740 (N_7740,N_6796,N_6982);
xor U7741 (N_7741,N_6970,N_6281);
nand U7742 (N_7742,N_6688,N_6560);
nand U7743 (N_7743,N_6817,N_6452);
nand U7744 (N_7744,N_6331,N_6293);
or U7745 (N_7745,N_6443,N_6359);
nand U7746 (N_7746,N_6094,N_6991);
nor U7747 (N_7747,N_6177,N_6563);
or U7748 (N_7748,N_6696,N_6924);
and U7749 (N_7749,N_6325,N_6560);
xor U7750 (N_7750,N_6909,N_6505);
and U7751 (N_7751,N_6548,N_6811);
or U7752 (N_7752,N_6902,N_6491);
nand U7753 (N_7753,N_6016,N_6661);
or U7754 (N_7754,N_6887,N_6950);
or U7755 (N_7755,N_6419,N_6409);
and U7756 (N_7756,N_6016,N_6789);
xnor U7757 (N_7757,N_6064,N_6442);
or U7758 (N_7758,N_6131,N_6712);
and U7759 (N_7759,N_6200,N_6985);
nand U7760 (N_7760,N_6445,N_6808);
nand U7761 (N_7761,N_6825,N_6823);
or U7762 (N_7762,N_6510,N_6315);
nor U7763 (N_7763,N_6235,N_6499);
nand U7764 (N_7764,N_6205,N_6876);
and U7765 (N_7765,N_6684,N_6103);
nor U7766 (N_7766,N_6723,N_6855);
and U7767 (N_7767,N_6741,N_6522);
nand U7768 (N_7768,N_6829,N_6737);
nor U7769 (N_7769,N_6168,N_6734);
nand U7770 (N_7770,N_6074,N_6793);
nand U7771 (N_7771,N_6322,N_6508);
nand U7772 (N_7772,N_6527,N_6082);
and U7773 (N_7773,N_6672,N_6700);
nand U7774 (N_7774,N_6868,N_6763);
nand U7775 (N_7775,N_6336,N_6582);
and U7776 (N_7776,N_6453,N_6253);
nor U7777 (N_7777,N_6289,N_6834);
and U7778 (N_7778,N_6772,N_6109);
nand U7779 (N_7779,N_6710,N_6545);
nor U7780 (N_7780,N_6884,N_6930);
or U7781 (N_7781,N_6775,N_6211);
nand U7782 (N_7782,N_6067,N_6385);
or U7783 (N_7783,N_6781,N_6265);
xnor U7784 (N_7784,N_6975,N_6394);
nand U7785 (N_7785,N_6660,N_6535);
nand U7786 (N_7786,N_6888,N_6642);
nand U7787 (N_7787,N_6324,N_6064);
nand U7788 (N_7788,N_6722,N_6542);
nor U7789 (N_7789,N_6060,N_6088);
and U7790 (N_7790,N_6371,N_6305);
nand U7791 (N_7791,N_6117,N_6195);
or U7792 (N_7792,N_6995,N_6361);
or U7793 (N_7793,N_6534,N_6041);
nand U7794 (N_7794,N_6265,N_6585);
and U7795 (N_7795,N_6672,N_6231);
nand U7796 (N_7796,N_6682,N_6128);
and U7797 (N_7797,N_6196,N_6069);
nor U7798 (N_7798,N_6466,N_6005);
and U7799 (N_7799,N_6824,N_6084);
nand U7800 (N_7800,N_6948,N_6063);
nor U7801 (N_7801,N_6862,N_6806);
and U7802 (N_7802,N_6548,N_6386);
nor U7803 (N_7803,N_6403,N_6471);
nand U7804 (N_7804,N_6779,N_6068);
or U7805 (N_7805,N_6405,N_6356);
nor U7806 (N_7806,N_6808,N_6983);
nor U7807 (N_7807,N_6785,N_6258);
nand U7808 (N_7808,N_6656,N_6803);
and U7809 (N_7809,N_6164,N_6341);
nor U7810 (N_7810,N_6621,N_6012);
nor U7811 (N_7811,N_6545,N_6895);
and U7812 (N_7812,N_6640,N_6551);
nor U7813 (N_7813,N_6476,N_6850);
and U7814 (N_7814,N_6385,N_6480);
or U7815 (N_7815,N_6984,N_6581);
and U7816 (N_7816,N_6777,N_6148);
or U7817 (N_7817,N_6685,N_6986);
nor U7818 (N_7818,N_6310,N_6481);
nand U7819 (N_7819,N_6554,N_6858);
nor U7820 (N_7820,N_6678,N_6302);
or U7821 (N_7821,N_6072,N_6943);
and U7822 (N_7822,N_6399,N_6580);
xor U7823 (N_7823,N_6283,N_6374);
and U7824 (N_7824,N_6108,N_6390);
and U7825 (N_7825,N_6914,N_6840);
nor U7826 (N_7826,N_6061,N_6003);
and U7827 (N_7827,N_6459,N_6823);
or U7828 (N_7828,N_6233,N_6877);
nand U7829 (N_7829,N_6545,N_6480);
nor U7830 (N_7830,N_6114,N_6072);
or U7831 (N_7831,N_6193,N_6766);
or U7832 (N_7832,N_6355,N_6235);
xnor U7833 (N_7833,N_6808,N_6434);
and U7834 (N_7834,N_6222,N_6531);
nor U7835 (N_7835,N_6870,N_6030);
nand U7836 (N_7836,N_6177,N_6210);
nor U7837 (N_7837,N_6451,N_6375);
nand U7838 (N_7838,N_6838,N_6230);
and U7839 (N_7839,N_6100,N_6044);
and U7840 (N_7840,N_6354,N_6835);
or U7841 (N_7841,N_6964,N_6623);
nand U7842 (N_7842,N_6728,N_6378);
and U7843 (N_7843,N_6009,N_6672);
and U7844 (N_7844,N_6459,N_6137);
or U7845 (N_7845,N_6312,N_6239);
xnor U7846 (N_7846,N_6389,N_6267);
or U7847 (N_7847,N_6992,N_6253);
or U7848 (N_7848,N_6528,N_6333);
and U7849 (N_7849,N_6690,N_6301);
nor U7850 (N_7850,N_6819,N_6073);
xnor U7851 (N_7851,N_6226,N_6859);
nand U7852 (N_7852,N_6581,N_6221);
nand U7853 (N_7853,N_6389,N_6534);
and U7854 (N_7854,N_6437,N_6840);
nor U7855 (N_7855,N_6189,N_6481);
nand U7856 (N_7856,N_6029,N_6034);
or U7857 (N_7857,N_6311,N_6902);
or U7858 (N_7858,N_6417,N_6717);
or U7859 (N_7859,N_6181,N_6838);
nand U7860 (N_7860,N_6234,N_6282);
xnor U7861 (N_7861,N_6255,N_6697);
xor U7862 (N_7862,N_6089,N_6673);
or U7863 (N_7863,N_6444,N_6336);
nand U7864 (N_7864,N_6721,N_6010);
and U7865 (N_7865,N_6781,N_6354);
and U7866 (N_7866,N_6961,N_6012);
nor U7867 (N_7867,N_6463,N_6839);
nand U7868 (N_7868,N_6861,N_6039);
or U7869 (N_7869,N_6529,N_6294);
xor U7870 (N_7870,N_6462,N_6999);
nand U7871 (N_7871,N_6190,N_6646);
nor U7872 (N_7872,N_6915,N_6034);
or U7873 (N_7873,N_6261,N_6264);
or U7874 (N_7874,N_6103,N_6791);
nand U7875 (N_7875,N_6827,N_6127);
and U7876 (N_7876,N_6874,N_6511);
and U7877 (N_7877,N_6300,N_6063);
and U7878 (N_7878,N_6455,N_6125);
nor U7879 (N_7879,N_6799,N_6782);
xnor U7880 (N_7880,N_6166,N_6035);
or U7881 (N_7881,N_6235,N_6238);
nand U7882 (N_7882,N_6132,N_6759);
and U7883 (N_7883,N_6978,N_6069);
nand U7884 (N_7884,N_6241,N_6722);
nand U7885 (N_7885,N_6881,N_6880);
xnor U7886 (N_7886,N_6569,N_6874);
nand U7887 (N_7887,N_6762,N_6225);
or U7888 (N_7888,N_6772,N_6128);
or U7889 (N_7889,N_6552,N_6816);
and U7890 (N_7890,N_6387,N_6639);
nand U7891 (N_7891,N_6399,N_6818);
nor U7892 (N_7892,N_6656,N_6011);
xor U7893 (N_7893,N_6417,N_6701);
and U7894 (N_7894,N_6805,N_6335);
or U7895 (N_7895,N_6701,N_6256);
or U7896 (N_7896,N_6283,N_6938);
xnor U7897 (N_7897,N_6421,N_6766);
or U7898 (N_7898,N_6130,N_6110);
and U7899 (N_7899,N_6203,N_6417);
and U7900 (N_7900,N_6710,N_6633);
or U7901 (N_7901,N_6447,N_6241);
or U7902 (N_7902,N_6976,N_6274);
and U7903 (N_7903,N_6029,N_6890);
and U7904 (N_7904,N_6777,N_6412);
and U7905 (N_7905,N_6531,N_6390);
and U7906 (N_7906,N_6667,N_6161);
nand U7907 (N_7907,N_6956,N_6391);
or U7908 (N_7908,N_6727,N_6869);
nand U7909 (N_7909,N_6713,N_6436);
xnor U7910 (N_7910,N_6475,N_6424);
nand U7911 (N_7911,N_6626,N_6374);
or U7912 (N_7912,N_6440,N_6725);
nor U7913 (N_7913,N_6175,N_6253);
nor U7914 (N_7914,N_6635,N_6032);
nor U7915 (N_7915,N_6839,N_6319);
nor U7916 (N_7916,N_6093,N_6756);
or U7917 (N_7917,N_6722,N_6134);
nand U7918 (N_7918,N_6577,N_6229);
nor U7919 (N_7919,N_6521,N_6611);
and U7920 (N_7920,N_6678,N_6175);
or U7921 (N_7921,N_6053,N_6366);
and U7922 (N_7922,N_6289,N_6005);
and U7923 (N_7923,N_6892,N_6203);
nand U7924 (N_7924,N_6902,N_6014);
nand U7925 (N_7925,N_6697,N_6668);
or U7926 (N_7926,N_6512,N_6141);
and U7927 (N_7927,N_6208,N_6287);
nor U7928 (N_7928,N_6181,N_6958);
and U7929 (N_7929,N_6449,N_6544);
and U7930 (N_7930,N_6435,N_6977);
nor U7931 (N_7931,N_6191,N_6126);
nand U7932 (N_7932,N_6061,N_6493);
nand U7933 (N_7933,N_6238,N_6654);
or U7934 (N_7934,N_6614,N_6343);
nand U7935 (N_7935,N_6999,N_6135);
nor U7936 (N_7936,N_6360,N_6539);
or U7937 (N_7937,N_6055,N_6988);
xnor U7938 (N_7938,N_6487,N_6377);
nand U7939 (N_7939,N_6783,N_6846);
or U7940 (N_7940,N_6399,N_6642);
nor U7941 (N_7941,N_6839,N_6723);
or U7942 (N_7942,N_6703,N_6746);
nand U7943 (N_7943,N_6527,N_6210);
nand U7944 (N_7944,N_6789,N_6242);
nor U7945 (N_7945,N_6050,N_6529);
or U7946 (N_7946,N_6966,N_6744);
xor U7947 (N_7947,N_6113,N_6195);
xnor U7948 (N_7948,N_6116,N_6728);
nor U7949 (N_7949,N_6703,N_6515);
nor U7950 (N_7950,N_6115,N_6626);
xnor U7951 (N_7951,N_6488,N_6204);
xor U7952 (N_7952,N_6167,N_6088);
and U7953 (N_7953,N_6710,N_6729);
and U7954 (N_7954,N_6454,N_6477);
and U7955 (N_7955,N_6435,N_6839);
or U7956 (N_7956,N_6577,N_6640);
and U7957 (N_7957,N_6338,N_6464);
or U7958 (N_7958,N_6979,N_6726);
or U7959 (N_7959,N_6742,N_6774);
nand U7960 (N_7960,N_6295,N_6580);
xor U7961 (N_7961,N_6924,N_6015);
and U7962 (N_7962,N_6337,N_6347);
and U7963 (N_7963,N_6854,N_6168);
and U7964 (N_7964,N_6817,N_6558);
nand U7965 (N_7965,N_6380,N_6586);
or U7966 (N_7966,N_6336,N_6274);
and U7967 (N_7967,N_6559,N_6919);
and U7968 (N_7968,N_6742,N_6487);
nand U7969 (N_7969,N_6600,N_6937);
nor U7970 (N_7970,N_6420,N_6498);
nand U7971 (N_7971,N_6543,N_6651);
xnor U7972 (N_7972,N_6119,N_6284);
and U7973 (N_7973,N_6265,N_6166);
xnor U7974 (N_7974,N_6110,N_6333);
and U7975 (N_7975,N_6962,N_6007);
and U7976 (N_7976,N_6731,N_6947);
and U7977 (N_7977,N_6162,N_6860);
or U7978 (N_7978,N_6149,N_6070);
nor U7979 (N_7979,N_6822,N_6229);
xor U7980 (N_7980,N_6683,N_6866);
nand U7981 (N_7981,N_6881,N_6214);
and U7982 (N_7982,N_6827,N_6504);
nand U7983 (N_7983,N_6355,N_6018);
and U7984 (N_7984,N_6225,N_6445);
nand U7985 (N_7985,N_6106,N_6451);
xnor U7986 (N_7986,N_6042,N_6144);
xor U7987 (N_7987,N_6829,N_6079);
or U7988 (N_7988,N_6474,N_6057);
nor U7989 (N_7989,N_6855,N_6285);
nor U7990 (N_7990,N_6863,N_6917);
nand U7991 (N_7991,N_6116,N_6907);
or U7992 (N_7992,N_6084,N_6003);
or U7993 (N_7993,N_6897,N_6455);
or U7994 (N_7994,N_6015,N_6997);
and U7995 (N_7995,N_6208,N_6693);
or U7996 (N_7996,N_6359,N_6140);
nor U7997 (N_7997,N_6952,N_6751);
or U7998 (N_7998,N_6992,N_6821);
and U7999 (N_7999,N_6668,N_6894);
xnor U8000 (N_8000,N_7507,N_7167);
nor U8001 (N_8001,N_7951,N_7378);
nand U8002 (N_8002,N_7882,N_7393);
nand U8003 (N_8003,N_7346,N_7548);
nor U8004 (N_8004,N_7120,N_7181);
and U8005 (N_8005,N_7783,N_7028);
and U8006 (N_8006,N_7675,N_7004);
and U8007 (N_8007,N_7281,N_7743);
nor U8008 (N_8008,N_7283,N_7449);
nor U8009 (N_8009,N_7118,N_7288);
nor U8010 (N_8010,N_7170,N_7553);
nor U8011 (N_8011,N_7960,N_7849);
nand U8012 (N_8012,N_7663,N_7726);
xor U8013 (N_8013,N_7855,N_7116);
nand U8014 (N_8014,N_7987,N_7072);
xor U8015 (N_8015,N_7404,N_7224);
nand U8016 (N_8016,N_7262,N_7479);
nand U8017 (N_8017,N_7308,N_7785);
nand U8018 (N_8018,N_7727,N_7935);
nor U8019 (N_8019,N_7434,N_7566);
nand U8020 (N_8020,N_7252,N_7477);
nand U8021 (N_8021,N_7606,N_7319);
and U8022 (N_8022,N_7327,N_7917);
nor U8023 (N_8023,N_7988,N_7561);
xor U8024 (N_8024,N_7840,N_7552);
and U8025 (N_8025,N_7919,N_7054);
and U8026 (N_8026,N_7801,N_7196);
and U8027 (N_8027,N_7233,N_7356);
nor U8028 (N_8028,N_7459,N_7753);
or U8029 (N_8029,N_7842,N_7257);
nand U8030 (N_8030,N_7610,N_7789);
and U8031 (N_8031,N_7518,N_7201);
nor U8032 (N_8032,N_7683,N_7469);
or U8033 (N_8033,N_7556,N_7089);
or U8034 (N_8034,N_7210,N_7739);
nor U8035 (N_8035,N_7289,N_7202);
or U8036 (N_8036,N_7578,N_7784);
nor U8037 (N_8037,N_7057,N_7885);
nor U8038 (N_8038,N_7109,N_7395);
and U8039 (N_8039,N_7482,N_7156);
xnor U8040 (N_8040,N_7749,N_7690);
and U8041 (N_8041,N_7423,N_7208);
and U8042 (N_8042,N_7284,N_7833);
nor U8043 (N_8043,N_7936,N_7446);
nor U8044 (N_8044,N_7557,N_7030);
and U8045 (N_8045,N_7523,N_7586);
nand U8046 (N_8046,N_7192,N_7154);
nand U8047 (N_8047,N_7033,N_7629);
nand U8048 (N_8048,N_7517,N_7326);
and U8049 (N_8049,N_7144,N_7648);
and U8050 (N_8050,N_7619,N_7817);
or U8051 (N_8051,N_7755,N_7843);
nand U8052 (N_8052,N_7155,N_7480);
or U8053 (N_8053,N_7896,N_7915);
nand U8054 (N_8054,N_7153,N_7379);
or U8055 (N_8055,N_7246,N_7145);
and U8056 (N_8056,N_7824,N_7363);
nor U8057 (N_8057,N_7130,N_7105);
nor U8058 (N_8058,N_7403,N_7978);
nor U8059 (N_8059,N_7137,N_7168);
nor U8060 (N_8060,N_7044,N_7362);
nor U8061 (N_8061,N_7377,N_7001);
and U8062 (N_8062,N_7983,N_7803);
nand U8063 (N_8063,N_7686,N_7741);
xnor U8064 (N_8064,N_7601,N_7331);
nor U8065 (N_8065,N_7721,N_7138);
and U8066 (N_8066,N_7856,N_7002);
xor U8067 (N_8067,N_7699,N_7024);
and U8068 (N_8068,N_7938,N_7544);
or U8069 (N_8069,N_7330,N_7188);
or U8070 (N_8070,N_7035,N_7515);
nor U8071 (N_8071,N_7952,N_7055);
or U8072 (N_8072,N_7441,N_7143);
or U8073 (N_8073,N_7348,N_7718);
nand U8074 (N_8074,N_7668,N_7345);
nand U8075 (N_8075,N_7414,N_7643);
and U8076 (N_8076,N_7191,N_7198);
nor U8077 (N_8077,N_7660,N_7111);
and U8078 (N_8078,N_7813,N_7861);
or U8079 (N_8079,N_7209,N_7332);
nor U8080 (N_8080,N_7897,N_7872);
or U8081 (N_8081,N_7231,N_7802);
xnor U8082 (N_8082,N_7923,N_7133);
or U8083 (N_8083,N_7826,N_7751);
nor U8084 (N_8084,N_7452,N_7505);
or U8085 (N_8085,N_7436,N_7835);
xnor U8086 (N_8086,N_7081,N_7406);
or U8087 (N_8087,N_7779,N_7074);
nand U8088 (N_8088,N_7195,N_7169);
xnor U8089 (N_8089,N_7763,N_7388);
and U8090 (N_8090,N_7239,N_7943);
nor U8091 (N_8091,N_7053,N_7493);
or U8092 (N_8092,N_7747,N_7485);
xnor U8093 (N_8093,N_7806,N_7720);
nand U8094 (N_8094,N_7086,N_7647);
and U8095 (N_8095,N_7732,N_7029);
xnor U8096 (N_8096,N_7772,N_7961);
and U8097 (N_8097,N_7719,N_7017);
and U8098 (N_8098,N_7254,N_7757);
nand U8099 (N_8099,N_7618,N_7337);
or U8100 (N_8100,N_7582,N_7863);
or U8101 (N_8101,N_7904,N_7091);
nand U8102 (N_8102,N_7980,N_7008);
nor U8103 (N_8103,N_7929,N_7574);
nor U8104 (N_8104,N_7588,N_7812);
and U8105 (N_8105,N_7103,N_7365);
and U8106 (N_8106,N_7309,N_7922);
or U8107 (N_8107,N_7685,N_7124);
nand U8108 (N_8108,N_7948,N_7134);
nor U8109 (N_8109,N_7598,N_7958);
and U8110 (N_8110,N_7429,N_7394);
and U8111 (N_8111,N_7914,N_7359);
nand U8112 (N_8112,N_7247,N_7005);
and U8113 (N_8113,N_7075,N_7099);
nand U8114 (N_8114,N_7298,N_7009);
and U8115 (N_8115,N_7818,N_7616);
nand U8116 (N_8116,N_7318,N_7748);
nor U8117 (N_8117,N_7814,N_7650);
and U8118 (N_8118,N_7524,N_7768);
nor U8119 (N_8119,N_7995,N_7771);
nand U8120 (N_8120,N_7859,N_7569);
xnor U8121 (N_8121,N_7368,N_7628);
nand U8122 (N_8122,N_7034,N_7585);
nand U8123 (N_8123,N_7085,N_7642);
and U8124 (N_8124,N_7678,N_7049);
or U8125 (N_8125,N_7496,N_7228);
or U8126 (N_8126,N_7846,N_7399);
xnor U8127 (N_8127,N_7364,N_7697);
and U8128 (N_8128,N_7920,N_7632);
or U8129 (N_8129,N_7096,N_7537);
and U8130 (N_8130,N_7232,N_7221);
nand U8131 (N_8131,N_7163,N_7871);
nand U8132 (N_8132,N_7680,N_7993);
nor U8133 (N_8133,N_7571,N_7682);
nor U8134 (N_8134,N_7060,N_7945);
or U8135 (N_8135,N_7038,N_7750);
xnor U8136 (N_8136,N_7724,N_7893);
and U8137 (N_8137,N_7305,N_7862);
nand U8138 (N_8138,N_7531,N_7249);
xor U8139 (N_8139,N_7702,N_7455);
xnor U8140 (N_8140,N_7870,N_7745);
xnor U8141 (N_8141,N_7592,N_7177);
nand U8142 (N_8142,N_7982,N_7850);
xnor U8143 (N_8143,N_7800,N_7770);
nor U8144 (N_8144,N_7694,N_7953);
and U8145 (N_8145,N_7339,N_7707);
or U8146 (N_8146,N_7046,N_7189);
nor U8147 (N_8147,N_7067,N_7905);
nor U8148 (N_8148,N_7860,N_7821);
nor U8149 (N_8149,N_7389,N_7401);
or U8150 (N_8150,N_7928,N_7303);
or U8151 (N_8151,N_7278,N_7639);
nor U8152 (N_8152,N_7659,N_7672);
and U8153 (N_8153,N_7733,N_7324);
nor U8154 (N_8154,N_7158,N_7061);
and U8155 (N_8155,N_7558,N_7218);
nand U8156 (N_8156,N_7612,N_7413);
nor U8157 (N_8157,N_7023,N_7152);
nand U8158 (N_8158,N_7355,N_7123);
nand U8159 (N_8159,N_7489,N_7693);
and U8160 (N_8160,N_7119,N_7594);
nor U8161 (N_8161,N_7658,N_7015);
and U8162 (N_8162,N_7581,N_7142);
and U8163 (N_8163,N_7966,N_7357);
nand U8164 (N_8164,N_7754,N_7907);
nor U8165 (N_8165,N_7827,N_7347);
and U8166 (N_8166,N_7613,N_7090);
nand U8167 (N_8167,N_7596,N_7227);
nor U8168 (N_8168,N_7725,N_7443);
and U8169 (N_8169,N_7799,N_7352);
nor U8170 (N_8170,N_7621,N_7723);
nor U8171 (N_8171,N_7466,N_7106);
or U8172 (N_8172,N_7780,N_7161);
nor U8173 (N_8173,N_7492,N_7662);
xor U8174 (N_8174,N_7657,N_7491);
or U8175 (N_8175,N_7398,N_7323);
or U8176 (N_8176,N_7992,N_7104);
and U8177 (N_8177,N_7756,N_7059);
and U8178 (N_8178,N_7165,N_7782);
nor U8179 (N_8179,N_7912,N_7937);
and U8180 (N_8180,N_7121,N_7867);
nand U8181 (N_8181,N_7730,N_7036);
nand U8182 (N_8182,N_7516,N_7708);
or U8183 (N_8183,N_7101,N_7869);
or U8184 (N_8184,N_7962,N_7473);
xor U8185 (N_8185,N_7635,N_7894);
nand U8186 (N_8186,N_7568,N_7955);
nand U8187 (N_8187,N_7243,N_7888);
nand U8188 (N_8188,N_7972,N_7875);
nor U8189 (N_8189,N_7865,N_7590);
and U8190 (N_8190,N_7458,N_7230);
nand U8191 (N_8191,N_7792,N_7385);
and U8192 (N_8192,N_7440,N_7409);
nor U8193 (N_8193,N_7013,N_7020);
nand U8194 (N_8194,N_7216,N_7173);
xor U8195 (N_8195,N_7149,N_7025);
or U8196 (N_8196,N_7942,N_7847);
nor U8197 (N_8197,N_7302,N_7903);
xor U8198 (N_8198,N_7819,N_7194);
or U8199 (N_8199,N_7710,N_7217);
xnor U8200 (N_8200,N_7714,N_7380);
xor U8201 (N_8201,N_7712,N_7047);
xnor U8202 (N_8202,N_7175,N_7190);
xor U8203 (N_8203,N_7640,N_7563);
nor U8204 (N_8204,N_7212,N_7127);
or U8205 (N_8205,N_7110,N_7831);
or U8206 (N_8206,N_7361,N_7384);
xnor U8207 (N_8207,N_7372,N_7226);
nor U8208 (N_8208,N_7963,N_7665);
or U8209 (N_8209,N_7066,N_7971);
or U8210 (N_8210,N_7711,N_7911);
or U8211 (N_8211,N_7615,N_7270);
nor U8212 (N_8212,N_7624,N_7497);
xor U8213 (N_8213,N_7798,N_7898);
or U8214 (N_8214,N_7369,N_7397);
and U8215 (N_8215,N_7607,N_7019);
xnor U8216 (N_8216,N_7215,N_7206);
or U8217 (N_8217,N_7744,N_7391);
xor U8218 (N_8218,N_7087,N_7554);
or U8219 (N_8219,N_7631,N_7630);
xor U8220 (N_8220,N_7830,N_7451);
nor U8221 (N_8221,N_7265,N_7781);
and U8222 (N_8222,N_7010,N_7462);
and U8223 (N_8223,N_7453,N_7437);
and U8224 (N_8224,N_7884,N_7713);
or U8225 (N_8225,N_7535,N_7486);
and U8226 (N_8226,N_7128,N_7716);
nand U8227 (N_8227,N_7921,N_7135);
and U8228 (N_8228,N_7320,N_7287);
or U8229 (N_8229,N_7698,N_7979);
nor U8230 (N_8230,N_7522,N_7509);
nand U8231 (N_8231,N_7811,N_7545);
nor U8232 (N_8232,N_7828,N_7845);
nor U8233 (N_8233,N_7511,N_7787);
nor U8234 (N_8234,N_7197,N_7649);
nor U8235 (N_8235,N_7696,N_7494);
nand U8236 (N_8236,N_7073,N_7609);
nand U8237 (N_8237,N_7570,N_7521);
and U8238 (N_8238,N_7102,N_7573);
and U8239 (N_8239,N_7392,N_7341);
or U8240 (N_8240,N_7674,N_7200);
xor U8241 (N_8241,N_7400,N_7562);
and U8242 (N_8242,N_7311,N_7475);
or U8243 (N_8243,N_7874,N_7031);
or U8244 (N_8244,N_7541,N_7816);
nor U8245 (N_8245,N_7108,N_7931);
or U8246 (N_8246,N_7261,N_7184);
nor U8247 (N_8247,N_7051,N_7185);
nor U8248 (N_8248,N_7868,N_7676);
and U8249 (N_8249,N_7706,N_7762);
xnor U8250 (N_8250,N_7530,N_7402);
and U8251 (N_8251,N_7390,N_7836);
nor U8252 (N_8252,N_7131,N_7350);
or U8253 (N_8253,N_7589,N_7709);
nand U8254 (N_8254,N_7236,N_7795);
or U8255 (N_8255,N_7513,N_7333);
nor U8256 (N_8256,N_7959,N_7605);
and U8257 (N_8257,N_7366,N_7746);
nand U8258 (N_8258,N_7508,N_7974);
nand U8259 (N_8259,N_7584,N_7947);
nor U8260 (N_8260,N_7758,N_7367);
nor U8261 (N_8261,N_7839,N_7307);
or U8262 (N_8262,N_7576,N_7299);
nand U8263 (N_8263,N_7048,N_7250);
nor U8264 (N_8264,N_7891,N_7503);
nor U8265 (N_8265,N_7889,N_7731);
nand U8266 (N_8266,N_7622,N_7916);
or U8267 (N_8267,N_7176,N_7256);
or U8268 (N_8268,N_7810,N_7740);
nor U8269 (N_8269,N_7941,N_7500);
and U8270 (N_8270,N_7269,N_7300);
or U8271 (N_8271,N_7994,N_7141);
and U8272 (N_8272,N_7428,N_7444);
nand U8273 (N_8273,N_7910,N_7258);
nand U8274 (N_8274,N_7241,N_7673);
or U8275 (N_8275,N_7041,N_7358);
and U8276 (N_8276,N_7292,N_7572);
xor U8277 (N_8277,N_7179,N_7229);
nand U8278 (N_8278,N_7895,N_7114);
and U8279 (N_8279,N_7408,N_7906);
nor U8280 (N_8280,N_7052,N_7877);
or U8281 (N_8281,N_7722,N_7312);
nor U8282 (N_8282,N_7924,N_7166);
and U8283 (N_8283,N_7238,N_7483);
nor U8284 (N_8284,N_7335,N_7704);
and U8285 (N_8285,N_7656,N_7774);
or U8286 (N_8286,N_7881,N_7769);
or U8287 (N_8287,N_7207,N_7234);
nand U8288 (N_8288,N_7815,N_7764);
or U8289 (N_8289,N_7100,N_7555);
or U8290 (N_8290,N_7543,N_7790);
and U8291 (N_8291,N_7536,N_7652);
or U8292 (N_8292,N_7506,N_7064);
nor U8293 (N_8293,N_7421,N_7975);
nand U8294 (N_8294,N_7538,N_7684);
nand U8295 (N_8295,N_7286,N_7671);
xor U8296 (N_8296,N_7878,N_7012);
nand U8297 (N_8297,N_7000,N_7834);
or U8298 (N_8298,N_7575,N_7290);
or U8299 (N_8299,N_7094,N_7759);
nor U8300 (N_8300,N_7248,N_7285);
nand U8301 (N_8301,N_7396,N_7510);
or U8302 (N_8302,N_7418,N_7688);
xor U8303 (N_8303,N_7083,N_7183);
or U8304 (N_8304,N_7797,N_7260);
and U8305 (N_8305,N_7641,N_7180);
or U8306 (N_8306,N_7954,N_7301);
nor U8307 (N_8307,N_7514,N_7251);
or U8308 (N_8308,N_7587,N_7525);
nor U8309 (N_8309,N_7864,N_7646);
or U8310 (N_8310,N_7266,N_7767);
nand U8311 (N_8311,N_7848,N_7140);
nor U8312 (N_8312,N_7334,N_7148);
or U8313 (N_8313,N_7752,N_7040);
nor U8314 (N_8314,N_7687,N_7844);
or U8315 (N_8315,N_7014,N_7417);
nor U8316 (N_8316,N_7463,N_7115);
nor U8317 (N_8317,N_7042,N_7807);
xnor U8318 (N_8318,N_7472,N_7328);
nand U8319 (N_8319,N_7419,N_7296);
and U8320 (N_8320,N_7532,N_7879);
xor U8321 (N_8321,N_7913,N_7625);
or U8322 (N_8322,N_7321,N_7484);
nor U8323 (N_8323,N_7620,N_7794);
or U8324 (N_8324,N_7203,N_7433);
or U8325 (N_8325,N_7039,N_7273);
or U8326 (N_8326,N_7126,N_7985);
nand U8327 (N_8327,N_7591,N_7549);
nor U8328 (N_8328,N_7435,N_7223);
or U8329 (N_8329,N_7129,N_7735);
or U8330 (N_8330,N_7317,N_7310);
and U8331 (N_8331,N_7032,N_7018);
nand U8332 (N_8332,N_7011,N_7991);
and U8333 (N_8333,N_7851,N_7354);
and U8334 (N_8334,N_7426,N_7946);
nand U8335 (N_8335,N_7715,N_7737);
or U8336 (N_8336,N_7742,N_7661);
or U8337 (N_8337,N_7003,N_7351);
nand U8338 (N_8338,N_7957,N_7465);
xnor U8339 (N_8339,N_7069,N_7495);
or U8340 (N_8340,N_7279,N_7139);
nand U8341 (N_8341,N_7939,N_7095);
or U8342 (N_8342,N_7965,N_7222);
or U8343 (N_8343,N_7211,N_7079);
or U8344 (N_8344,N_7450,N_7823);
nor U8345 (N_8345,N_7186,N_7930);
and U8346 (N_8346,N_7386,N_7411);
and U8347 (N_8347,N_7567,N_7078);
and U8348 (N_8348,N_7374,N_7007);
or U8349 (N_8349,N_7457,N_7478);
or U8350 (N_8350,N_7021,N_7604);
nand U8351 (N_8351,N_7677,N_7313);
and U8352 (N_8352,N_7529,N_7542);
or U8353 (N_8353,N_7022,N_7276);
and U8354 (N_8354,N_7220,N_7205);
nor U8355 (N_8355,N_7773,N_7527);
nand U8356 (N_8356,N_7634,N_7490);
nand U8357 (N_8357,N_7984,N_7858);
or U8358 (N_8358,N_7268,N_7277);
nand U8359 (N_8359,N_7460,N_7376);
and U8360 (N_8360,N_7692,N_7342);
xnor U8361 (N_8361,N_7820,N_7970);
xor U8362 (N_8362,N_7550,N_7832);
and U8363 (N_8363,N_7540,N_7944);
and U8364 (N_8364,N_7439,N_7125);
nand U8365 (N_8365,N_7245,N_7777);
or U8366 (N_8366,N_7445,N_7499);
nand U8367 (N_8367,N_7695,N_7967);
nor U8368 (N_8368,N_7071,N_7968);
and U8369 (N_8369,N_7886,N_7442);
or U8370 (N_8370,N_7371,N_7255);
nor U8371 (N_8371,N_7214,N_7796);
nor U8372 (N_8372,N_7043,N_7876);
or U8373 (N_8373,N_7461,N_7172);
nand U8374 (N_8374,N_7887,N_7097);
nor U8375 (N_8375,N_7880,N_7599);
nand U8376 (N_8376,N_7274,N_7178);
or U8377 (N_8377,N_7271,N_7112);
and U8378 (N_8378,N_7242,N_7295);
nor U8379 (N_8379,N_7431,N_7297);
xor U8380 (N_8380,N_7805,N_7853);
nand U8381 (N_8381,N_7565,N_7653);
or U8382 (N_8382,N_7873,N_7107);
xor U8383 (N_8383,N_7058,N_7579);
and U8384 (N_8384,N_7088,N_7092);
nand U8385 (N_8385,N_7825,N_7852);
or U8386 (N_8386,N_7808,N_7070);
nor U8387 (N_8387,N_7933,N_7997);
or U8388 (N_8388,N_7412,N_7171);
and U8389 (N_8389,N_7998,N_7076);
nand U8390 (N_8390,N_7340,N_7927);
or U8391 (N_8391,N_7304,N_7338);
or U8392 (N_8392,N_7026,N_7528);
xnor U8393 (N_8393,N_7822,N_7892);
nand U8394 (N_8394,N_7539,N_7559);
xor U8395 (N_8395,N_7560,N_7432);
xor U8396 (N_8396,N_7577,N_7909);
and U8397 (N_8397,N_7456,N_7204);
or U8398 (N_8398,N_7387,N_7608);
nor U8399 (N_8399,N_7883,N_7322);
or U8400 (N_8400,N_7809,N_7705);
xnor U8401 (N_8401,N_7240,N_7375);
nor U8402 (N_8402,N_7761,N_7275);
nand U8403 (N_8403,N_7866,N_7996);
nand U8404 (N_8404,N_7027,N_7160);
xnor U8405 (N_8405,N_7890,N_7117);
nor U8406 (N_8406,N_7681,N_7602);
or U8407 (N_8407,N_7969,N_7738);
and U8408 (N_8408,N_7199,N_7551);
and U8409 (N_8409,N_7150,N_7857);
or U8410 (N_8410,N_7977,N_7651);
nor U8411 (N_8411,N_7990,N_7837);
nor U8412 (N_8412,N_7068,N_7564);
or U8413 (N_8413,N_7050,N_7416);
or U8414 (N_8414,N_7595,N_7316);
and U8415 (N_8415,N_7056,N_7934);
nor U8416 (N_8416,N_7213,N_7989);
and U8417 (N_8417,N_7136,N_7430);
and U8418 (N_8418,N_7425,N_7925);
or U8419 (N_8419,N_7468,N_7065);
or U8420 (N_8420,N_7077,N_7981);
nand U8421 (N_8421,N_7282,N_7793);
nor U8422 (N_8422,N_7546,N_7410);
nor U8423 (N_8423,N_7617,N_7644);
or U8424 (N_8424,N_7519,N_7264);
xor U8425 (N_8425,N_7600,N_7336);
xnor U8426 (N_8426,N_7918,N_7382);
nand U8427 (N_8427,N_7901,N_7164);
nand U8428 (N_8428,N_7329,N_7765);
and U8429 (N_8429,N_7438,N_7623);
or U8430 (N_8430,N_7778,N_7315);
xnor U8431 (N_8431,N_7237,N_7926);
and U8432 (N_8432,N_7314,N_7999);
and U8433 (N_8433,N_7383,N_7098);
and U8434 (N_8434,N_7940,N_7964);
nand U8435 (N_8435,N_7728,N_7689);
and U8436 (N_8436,N_7679,N_7045);
and U8437 (N_8437,N_7691,N_7084);
or U8438 (N_8438,N_7280,N_7471);
nor U8439 (N_8439,N_7187,N_7580);
nor U8440 (N_8440,N_7294,N_7788);
nand U8441 (N_8441,N_7082,N_7306);
nor U8442 (N_8442,N_7786,N_7583);
and U8443 (N_8443,N_7267,N_7841);
or U8444 (N_8444,N_7775,N_7791);
nor U8445 (N_8445,N_7766,N_7146);
or U8446 (N_8446,N_7244,N_7534);
nand U8447 (N_8447,N_7415,N_7006);
or U8448 (N_8448,N_7474,N_7407);
nand U8449 (N_8449,N_7464,N_7932);
or U8450 (N_8450,N_7701,N_7908);
and U8451 (N_8451,N_7501,N_7829);
nand U8452 (N_8452,N_7636,N_7487);
or U8453 (N_8453,N_7986,N_7593);
nor U8454 (N_8454,N_7729,N_7654);
and U8455 (N_8455,N_7405,N_7902);
or U8456 (N_8456,N_7467,N_7424);
or U8457 (N_8457,N_7498,N_7700);
and U8458 (N_8458,N_7122,N_7037);
nor U8459 (N_8459,N_7151,N_7633);
nor U8460 (N_8460,N_7597,N_7637);
or U8461 (N_8461,N_7420,N_7353);
and U8462 (N_8462,N_7225,N_7488);
or U8463 (N_8463,N_7838,N_7147);
or U8464 (N_8464,N_7533,N_7804);
and U8465 (N_8465,N_7062,N_7504);
and U8466 (N_8466,N_7272,N_7080);
nand U8467 (N_8467,N_7481,N_7447);
or U8468 (N_8468,N_7626,N_7664);
and U8469 (N_8469,N_7476,N_7162);
nand U8470 (N_8470,N_7899,N_7360);
and U8471 (N_8471,N_7666,N_7427);
or U8472 (N_8472,N_7159,N_7854);
or U8473 (N_8473,N_7370,N_7614);
nand U8474 (N_8474,N_7293,N_7182);
and U8475 (N_8475,N_7655,N_7512);
or U8476 (N_8476,N_7063,N_7373);
or U8477 (N_8477,N_7776,N_7193);
or U8478 (N_8478,N_7603,N_7669);
or U8479 (N_8479,N_7422,N_7547);
or U8480 (N_8480,N_7950,N_7470);
nor U8481 (N_8481,N_7645,N_7736);
and U8482 (N_8482,N_7976,N_7627);
or U8483 (N_8483,N_7325,N_7526);
nor U8484 (N_8484,N_7949,N_7157);
nor U8485 (N_8485,N_7638,N_7520);
nor U8486 (N_8486,N_7016,N_7502);
nor U8487 (N_8487,N_7253,N_7093);
or U8488 (N_8488,N_7174,N_7703);
or U8489 (N_8489,N_7291,N_7448);
and U8490 (N_8490,N_7454,N_7900);
nor U8491 (N_8491,N_7973,N_7132);
nand U8492 (N_8492,N_7344,N_7219);
nor U8493 (N_8493,N_7235,N_7956);
xor U8494 (N_8494,N_7343,N_7349);
nor U8495 (N_8495,N_7113,N_7259);
and U8496 (N_8496,N_7263,N_7667);
or U8497 (N_8497,N_7670,N_7717);
nor U8498 (N_8498,N_7734,N_7381);
nor U8499 (N_8499,N_7760,N_7611);
or U8500 (N_8500,N_7533,N_7727);
nor U8501 (N_8501,N_7908,N_7919);
nand U8502 (N_8502,N_7639,N_7944);
and U8503 (N_8503,N_7873,N_7620);
and U8504 (N_8504,N_7327,N_7379);
nor U8505 (N_8505,N_7155,N_7013);
nand U8506 (N_8506,N_7039,N_7916);
and U8507 (N_8507,N_7350,N_7963);
or U8508 (N_8508,N_7568,N_7052);
nand U8509 (N_8509,N_7589,N_7214);
and U8510 (N_8510,N_7472,N_7199);
and U8511 (N_8511,N_7243,N_7669);
and U8512 (N_8512,N_7062,N_7974);
or U8513 (N_8513,N_7323,N_7842);
nor U8514 (N_8514,N_7053,N_7164);
and U8515 (N_8515,N_7192,N_7437);
and U8516 (N_8516,N_7752,N_7102);
xnor U8517 (N_8517,N_7175,N_7440);
xnor U8518 (N_8518,N_7335,N_7369);
nor U8519 (N_8519,N_7308,N_7258);
and U8520 (N_8520,N_7990,N_7080);
and U8521 (N_8521,N_7374,N_7172);
nand U8522 (N_8522,N_7664,N_7635);
nor U8523 (N_8523,N_7401,N_7928);
nand U8524 (N_8524,N_7120,N_7990);
or U8525 (N_8525,N_7149,N_7736);
nand U8526 (N_8526,N_7389,N_7387);
and U8527 (N_8527,N_7934,N_7914);
nor U8528 (N_8528,N_7943,N_7464);
xor U8529 (N_8529,N_7901,N_7290);
and U8530 (N_8530,N_7699,N_7266);
or U8531 (N_8531,N_7235,N_7762);
and U8532 (N_8532,N_7721,N_7871);
nor U8533 (N_8533,N_7969,N_7965);
nor U8534 (N_8534,N_7959,N_7587);
nand U8535 (N_8535,N_7407,N_7430);
nor U8536 (N_8536,N_7721,N_7276);
nand U8537 (N_8537,N_7716,N_7045);
xnor U8538 (N_8538,N_7429,N_7580);
nor U8539 (N_8539,N_7396,N_7257);
nand U8540 (N_8540,N_7100,N_7663);
and U8541 (N_8541,N_7279,N_7148);
nand U8542 (N_8542,N_7046,N_7123);
xor U8543 (N_8543,N_7818,N_7231);
and U8544 (N_8544,N_7774,N_7572);
or U8545 (N_8545,N_7922,N_7218);
or U8546 (N_8546,N_7217,N_7719);
or U8547 (N_8547,N_7779,N_7263);
nor U8548 (N_8548,N_7738,N_7008);
or U8549 (N_8549,N_7040,N_7618);
or U8550 (N_8550,N_7795,N_7763);
xor U8551 (N_8551,N_7219,N_7548);
nor U8552 (N_8552,N_7466,N_7648);
and U8553 (N_8553,N_7877,N_7567);
or U8554 (N_8554,N_7214,N_7848);
and U8555 (N_8555,N_7456,N_7522);
or U8556 (N_8556,N_7290,N_7615);
and U8557 (N_8557,N_7489,N_7721);
nand U8558 (N_8558,N_7741,N_7320);
and U8559 (N_8559,N_7914,N_7383);
or U8560 (N_8560,N_7170,N_7745);
and U8561 (N_8561,N_7060,N_7062);
and U8562 (N_8562,N_7339,N_7365);
and U8563 (N_8563,N_7126,N_7544);
and U8564 (N_8564,N_7980,N_7201);
and U8565 (N_8565,N_7014,N_7310);
nand U8566 (N_8566,N_7153,N_7189);
nor U8567 (N_8567,N_7892,N_7940);
nor U8568 (N_8568,N_7305,N_7028);
nor U8569 (N_8569,N_7668,N_7939);
or U8570 (N_8570,N_7284,N_7030);
nand U8571 (N_8571,N_7320,N_7780);
and U8572 (N_8572,N_7206,N_7809);
nand U8573 (N_8573,N_7364,N_7329);
nand U8574 (N_8574,N_7367,N_7041);
xor U8575 (N_8575,N_7118,N_7760);
or U8576 (N_8576,N_7879,N_7749);
nor U8577 (N_8577,N_7987,N_7780);
nor U8578 (N_8578,N_7237,N_7816);
nand U8579 (N_8579,N_7914,N_7196);
or U8580 (N_8580,N_7906,N_7009);
or U8581 (N_8581,N_7577,N_7595);
and U8582 (N_8582,N_7231,N_7035);
nor U8583 (N_8583,N_7093,N_7476);
nor U8584 (N_8584,N_7660,N_7761);
or U8585 (N_8585,N_7593,N_7715);
nor U8586 (N_8586,N_7783,N_7619);
and U8587 (N_8587,N_7244,N_7167);
nand U8588 (N_8588,N_7147,N_7066);
or U8589 (N_8589,N_7554,N_7003);
nor U8590 (N_8590,N_7466,N_7404);
nand U8591 (N_8591,N_7496,N_7247);
nor U8592 (N_8592,N_7277,N_7477);
xnor U8593 (N_8593,N_7481,N_7253);
xnor U8594 (N_8594,N_7774,N_7349);
or U8595 (N_8595,N_7338,N_7400);
nor U8596 (N_8596,N_7617,N_7245);
or U8597 (N_8597,N_7558,N_7633);
xor U8598 (N_8598,N_7835,N_7420);
nor U8599 (N_8599,N_7444,N_7721);
nand U8600 (N_8600,N_7248,N_7943);
or U8601 (N_8601,N_7369,N_7509);
nand U8602 (N_8602,N_7753,N_7550);
or U8603 (N_8603,N_7769,N_7620);
nand U8604 (N_8604,N_7647,N_7110);
xnor U8605 (N_8605,N_7765,N_7730);
or U8606 (N_8606,N_7726,N_7188);
or U8607 (N_8607,N_7246,N_7009);
or U8608 (N_8608,N_7865,N_7775);
nor U8609 (N_8609,N_7862,N_7818);
or U8610 (N_8610,N_7710,N_7009);
nor U8611 (N_8611,N_7444,N_7395);
nand U8612 (N_8612,N_7603,N_7474);
nand U8613 (N_8613,N_7148,N_7122);
or U8614 (N_8614,N_7013,N_7691);
or U8615 (N_8615,N_7797,N_7775);
or U8616 (N_8616,N_7922,N_7873);
nand U8617 (N_8617,N_7034,N_7434);
and U8618 (N_8618,N_7233,N_7232);
nand U8619 (N_8619,N_7278,N_7083);
or U8620 (N_8620,N_7581,N_7415);
or U8621 (N_8621,N_7238,N_7242);
nand U8622 (N_8622,N_7000,N_7508);
or U8623 (N_8623,N_7722,N_7095);
nand U8624 (N_8624,N_7907,N_7422);
xnor U8625 (N_8625,N_7020,N_7963);
nand U8626 (N_8626,N_7215,N_7343);
nand U8627 (N_8627,N_7761,N_7219);
xor U8628 (N_8628,N_7496,N_7889);
nor U8629 (N_8629,N_7615,N_7449);
and U8630 (N_8630,N_7605,N_7663);
nand U8631 (N_8631,N_7264,N_7294);
xor U8632 (N_8632,N_7850,N_7851);
or U8633 (N_8633,N_7580,N_7570);
and U8634 (N_8634,N_7708,N_7293);
nor U8635 (N_8635,N_7643,N_7201);
and U8636 (N_8636,N_7339,N_7513);
or U8637 (N_8637,N_7648,N_7791);
and U8638 (N_8638,N_7383,N_7246);
or U8639 (N_8639,N_7865,N_7302);
nor U8640 (N_8640,N_7243,N_7748);
and U8641 (N_8641,N_7959,N_7449);
nor U8642 (N_8642,N_7110,N_7720);
nor U8643 (N_8643,N_7412,N_7701);
nor U8644 (N_8644,N_7300,N_7671);
xnor U8645 (N_8645,N_7742,N_7986);
nor U8646 (N_8646,N_7318,N_7792);
or U8647 (N_8647,N_7698,N_7165);
nand U8648 (N_8648,N_7129,N_7038);
and U8649 (N_8649,N_7594,N_7300);
or U8650 (N_8650,N_7838,N_7925);
nor U8651 (N_8651,N_7684,N_7342);
and U8652 (N_8652,N_7579,N_7357);
or U8653 (N_8653,N_7608,N_7838);
nand U8654 (N_8654,N_7039,N_7921);
or U8655 (N_8655,N_7053,N_7621);
or U8656 (N_8656,N_7780,N_7458);
and U8657 (N_8657,N_7213,N_7302);
xnor U8658 (N_8658,N_7930,N_7605);
or U8659 (N_8659,N_7625,N_7585);
nor U8660 (N_8660,N_7533,N_7132);
or U8661 (N_8661,N_7663,N_7986);
nand U8662 (N_8662,N_7625,N_7992);
or U8663 (N_8663,N_7545,N_7043);
nand U8664 (N_8664,N_7514,N_7550);
nand U8665 (N_8665,N_7563,N_7301);
nand U8666 (N_8666,N_7004,N_7164);
nor U8667 (N_8667,N_7075,N_7290);
and U8668 (N_8668,N_7830,N_7374);
nor U8669 (N_8669,N_7498,N_7108);
and U8670 (N_8670,N_7448,N_7572);
nand U8671 (N_8671,N_7848,N_7694);
or U8672 (N_8672,N_7941,N_7055);
and U8673 (N_8673,N_7353,N_7398);
xor U8674 (N_8674,N_7616,N_7038);
nor U8675 (N_8675,N_7099,N_7316);
and U8676 (N_8676,N_7977,N_7700);
nor U8677 (N_8677,N_7067,N_7148);
xor U8678 (N_8678,N_7181,N_7639);
nor U8679 (N_8679,N_7074,N_7392);
nand U8680 (N_8680,N_7147,N_7819);
nand U8681 (N_8681,N_7021,N_7007);
and U8682 (N_8682,N_7873,N_7026);
or U8683 (N_8683,N_7392,N_7460);
nor U8684 (N_8684,N_7996,N_7573);
and U8685 (N_8685,N_7276,N_7677);
nor U8686 (N_8686,N_7479,N_7859);
or U8687 (N_8687,N_7825,N_7986);
nor U8688 (N_8688,N_7684,N_7554);
nand U8689 (N_8689,N_7821,N_7577);
or U8690 (N_8690,N_7150,N_7584);
or U8691 (N_8691,N_7923,N_7013);
and U8692 (N_8692,N_7447,N_7529);
and U8693 (N_8693,N_7824,N_7409);
nand U8694 (N_8694,N_7233,N_7162);
and U8695 (N_8695,N_7119,N_7919);
nor U8696 (N_8696,N_7502,N_7568);
nor U8697 (N_8697,N_7655,N_7206);
and U8698 (N_8698,N_7109,N_7580);
or U8699 (N_8699,N_7684,N_7842);
and U8700 (N_8700,N_7777,N_7731);
and U8701 (N_8701,N_7596,N_7399);
nand U8702 (N_8702,N_7886,N_7342);
and U8703 (N_8703,N_7087,N_7343);
or U8704 (N_8704,N_7329,N_7898);
and U8705 (N_8705,N_7794,N_7105);
xnor U8706 (N_8706,N_7798,N_7723);
or U8707 (N_8707,N_7660,N_7311);
and U8708 (N_8708,N_7762,N_7910);
or U8709 (N_8709,N_7376,N_7903);
xnor U8710 (N_8710,N_7415,N_7180);
and U8711 (N_8711,N_7953,N_7066);
nand U8712 (N_8712,N_7974,N_7540);
and U8713 (N_8713,N_7318,N_7172);
nor U8714 (N_8714,N_7515,N_7590);
or U8715 (N_8715,N_7382,N_7786);
nand U8716 (N_8716,N_7446,N_7210);
or U8717 (N_8717,N_7752,N_7420);
and U8718 (N_8718,N_7459,N_7331);
nor U8719 (N_8719,N_7599,N_7846);
and U8720 (N_8720,N_7986,N_7527);
xor U8721 (N_8721,N_7018,N_7906);
nand U8722 (N_8722,N_7978,N_7353);
or U8723 (N_8723,N_7262,N_7125);
nand U8724 (N_8724,N_7271,N_7188);
and U8725 (N_8725,N_7731,N_7122);
nor U8726 (N_8726,N_7139,N_7016);
xnor U8727 (N_8727,N_7335,N_7875);
or U8728 (N_8728,N_7322,N_7473);
nor U8729 (N_8729,N_7914,N_7040);
or U8730 (N_8730,N_7975,N_7701);
nand U8731 (N_8731,N_7554,N_7558);
and U8732 (N_8732,N_7170,N_7497);
nor U8733 (N_8733,N_7976,N_7705);
or U8734 (N_8734,N_7544,N_7943);
nor U8735 (N_8735,N_7798,N_7173);
nor U8736 (N_8736,N_7305,N_7600);
and U8737 (N_8737,N_7432,N_7540);
xnor U8738 (N_8738,N_7013,N_7274);
or U8739 (N_8739,N_7436,N_7465);
and U8740 (N_8740,N_7329,N_7365);
xor U8741 (N_8741,N_7397,N_7948);
and U8742 (N_8742,N_7490,N_7195);
and U8743 (N_8743,N_7822,N_7472);
and U8744 (N_8744,N_7824,N_7107);
nor U8745 (N_8745,N_7531,N_7094);
and U8746 (N_8746,N_7684,N_7474);
or U8747 (N_8747,N_7265,N_7494);
xnor U8748 (N_8748,N_7108,N_7059);
nor U8749 (N_8749,N_7649,N_7055);
and U8750 (N_8750,N_7343,N_7445);
nor U8751 (N_8751,N_7054,N_7584);
and U8752 (N_8752,N_7406,N_7416);
nor U8753 (N_8753,N_7898,N_7928);
nor U8754 (N_8754,N_7372,N_7179);
nor U8755 (N_8755,N_7528,N_7032);
or U8756 (N_8756,N_7691,N_7032);
nor U8757 (N_8757,N_7722,N_7410);
and U8758 (N_8758,N_7120,N_7790);
nand U8759 (N_8759,N_7048,N_7462);
nor U8760 (N_8760,N_7299,N_7443);
and U8761 (N_8761,N_7647,N_7103);
and U8762 (N_8762,N_7501,N_7435);
nand U8763 (N_8763,N_7823,N_7254);
xnor U8764 (N_8764,N_7291,N_7358);
nand U8765 (N_8765,N_7504,N_7851);
nor U8766 (N_8766,N_7270,N_7429);
and U8767 (N_8767,N_7150,N_7634);
or U8768 (N_8768,N_7889,N_7720);
and U8769 (N_8769,N_7274,N_7714);
xnor U8770 (N_8770,N_7927,N_7103);
nand U8771 (N_8771,N_7541,N_7020);
xnor U8772 (N_8772,N_7801,N_7452);
nand U8773 (N_8773,N_7272,N_7857);
nor U8774 (N_8774,N_7522,N_7612);
or U8775 (N_8775,N_7490,N_7933);
xor U8776 (N_8776,N_7700,N_7310);
and U8777 (N_8777,N_7388,N_7058);
or U8778 (N_8778,N_7500,N_7781);
xnor U8779 (N_8779,N_7563,N_7925);
nor U8780 (N_8780,N_7604,N_7919);
and U8781 (N_8781,N_7517,N_7475);
xor U8782 (N_8782,N_7416,N_7546);
nor U8783 (N_8783,N_7956,N_7193);
and U8784 (N_8784,N_7923,N_7710);
nor U8785 (N_8785,N_7642,N_7666);
xor U8786 (N_8786,N_7247,N_7429);
nor U8787 (N_8787,N_7420,N_7205);
and U8788 (N_8788,N_7013,N_7356);
nand U8789 (N_8789,N_7601,N_7253);
xnor U8790 (N_8790,N_7977,N_7300);
and U8791 (N_8791,N_7756,N_7136);
nor U8792 (N_8792,N_7398,N_7604);
nor U8793 (N_8793,N_7034,N_7802);
nor U8794 (N_8794,N_7562,N_7956);
and U8795 (N_8795,N_7142,N_7224);
nor U8796 (N_8796,N_7384,N_7432);
and U8797 (N_8797,N_7863,N_7832);
and U8798 (N_8798,N_7399,N_7484);
or U8799 (N_8799,N_7537,N_7562);
and U8800 (N_8800,N_7294,N_7047);
nor U8801 (N_8801,N_7530,N_7875);
or U8802 (N_8802,N_7536,N_7184);
and U8803 (N_8803,N_7118,N_7733);
nor U8804 (N_8804,N_7257,N_7429);
nor U8805 (N_8805,N_7752,N_7798);
and U8806 (N_8806,N_7386,N_7795);
and U8807 (N_8807,N_7689,N_7489);
nand U8808 (N_8808,N_7164,N_7130);
nand U8809 (N_8809,N_7124,N_7415);
nand U8810 (N_8810,N_7176,N_7575);
and U8811 (N_8811,N_7816,N_7759);
nor U8812 (N_8812,N_7727,N_7142);
nor U8813 (N_8813,N_7849,N_7182);
or U8814 (N_8814,N_7149,N_7104);
nor U8815 (N_8815,N_7339,N_7419);
nand U8816 (N_8816,N_7872,N_7562);
and U8817 (N_8817,N_7160,N_7564);
nand U8818 (N_8818,N_7874,N_7781);
nand U8819 (N_8819,N_7022,N_7155);
nor U8820 (N_8820,N_7605,N_7861);
nor U8821 (N_8821,N_7832,N_7104);
nor U8822 (N_8822,N_7635,N_7587);
and U8823 (N_8823,N_7822,N_7929);
and U8824 (N_8824,N_7755,N_7803);
or U8825 (N_8825,N_7166,N_7626);
nand U8826 (N_8826,N_7290,N_7136);
nor U8827 (N_8827,N_7445,N_7200);
nor U8828 (N_8828,N_7047,N_7741);
nand U8829 (N_8829,N_7975,N_7722);
nor U8830 (N_8830,N_7214,N_7647);
or U8831 (N_8831,N_7572,N_7633);
nor U8832 (N_8832,N_7681,N_7974);
nand U8833 (N_8833,N_7475,N_7805);
or U8834 (N_8834,N_7641,N_7657);
and U8835 (N_8835,N_7521,N_7667);
and U8836 (N_8836,N_7687,N_7314);
or U8837 (N_8837,N_7760,N_7789);
or U8838 (N_8838,N_7029,N_7544);
xnor U8839 (N_8839,N_7072,N_7351);
nor U8840 (N_8840,N_7172,N_7972);
nor U8841 (N_8841,N_7917,N_7350);
nand U8842 (N_8842,N_7471,N_7239);
and U8843 (N_8843,N_7232,N_7900);
nor U8844 (N_8844,N_7446,N_7770);
xor U8845 (N_8845,N_7245,N_7740);
or U8846 (N_8846,N_7454,N_7218);
or U8847 (N_8847,N_7227,N_7852);
xor U8848 (N_8848,N_7921,N_7656);
nor U8849 (N_8849,N_7657,N_7211);
or U8850 (N_8850,N_7743,N_7879);
nand U8851 (N_8851,N_7772,N_7868);
nand U8852 (N_8852,N_7170,N_7742);
nor U8853 (N_8853,N_7101,N_7721);
nand U8854 (N_8854,N_7544,N_7139);
and U8855 (N_8855,N_7368,N_7534);
nand U8856 (N_8856,N_7099,N_7409);
nand U8857 (N_8857,N_7327,N_7301);
nor U8858 (N_8858,N_7720,N_7028);
nand U8859 (N_8859,N_7235,N_7772);
or U8860 (N_8860,N_7596,N_7824);
and U8861 (N_8861,N_7514,N_7696);
and U8862 (N_8862,N_7307,N_7466);
nor U8863 (N_8863,N_7607,N_7972);
nand U8864 (N_8864,N_7181,N_7842);
nor U8865 (N_8865,N_7929,N_7527);
nand U8866 (N_8866,N_7107,N_7129);
or U8867 (N_8867,N_7561,N_7688);
nor U8868 (N_8868,N_7937,N_7021);
and U8869 (N_8869,N_7837,N_7822);
xnor U8870 (N_8870,N_7847,N_7913);
nand U8871 (N_8871,N_7980,N_7910);
nand U8872 (N_8872,N_7747,N_7994);
nand U8873 (N_8873,N_7340,N_7901);
or U8874 (N_8874,N_7148,N_7566);
or U8875 (N_8875,N_7733,N_7663);
or U8876 (N_8876,N_7744,N_7877);
xor U8877 (N_8877,N_7685,N_7167);
and U8878 (N_8878,N_7825,N_7916);
and U8879 (N_8879,N_7807,N_7323);
or U8880 (N_8880,N_7275,N_7833);
nor U8881 (N_8881,N_7025,N_7800);
or U8882 (N_8882,N_7036,N_7323);
and U8883 (N_8883,N_7598,N_7584);
or U8884 (N_8884,N_7570,N_7950);
nor U8885 (N_8885,N_7868,N_7298);
and U8886 (N_8886,N_7576,N_7830);
and U8887 (N_8887,N_7261,N_7642);
or U8888 (N_8888,N_7811,N_7494);
or U8889 (N_8889,N_7042,N_7521);
or U8890 (N_8890,N_7109,N_7519);
or U8891 (N_8891,N_7671,N_7042);
nor U8892 (N_8892,N_7818,N_7279);
nand U8893 (N_8893,N_7464,N_7845);
nor U8894 (N_8894,N_7873,N_7929);
xor U8895 (N_8895,N_7896,N_7357);
nand U8896 (N_8896,N_7336,N_7194);
or U8897 (N_8897,N_7859,N_7163);
and U8898 (N_8898,N_7385,N_7168);
and U8899 (N_8899,N_7940,N_7677);
nor U8900 (N_8900,N_7827,N_7205);
nand U8901 (N_8901,N_7628,N_7394);
nand U8902 (N_8902,N_7473,N_7655);
or U8903 (N_8903,N_7910,N_7387);
or U8904 (N_8904,N_7537,N_7508);
nand U8905 (N_8905,N_7239,N_7718);
nand U8906 (N_8906,N_7800,N_7413);
or U8907 (N_8907,N_7055,N_7506);
or U8908 (N_8908,N_7511,N_7780);
and U8909 (N_8909,N_7827,N_7935);
nor U8910 (N_8910,N_7138,N_7458);
and U8911 (N_8911,N_7683,N_7876);
nand U8912 (N_8912,N_7483,N_7740);
nor U8913 (N_8913,N_7316,N_7729);
xor U8914 (N_8914,N_7372,N_7005);
nand U8915 (N_8915,N_7314,N_7686);
and U8916 (N_8916,N_7009,N_7474);
and U8917 (N_8917,N_7628,N_7811);
or U8918 (N_8918,N_7688,N_7150);
nor U8919 (N_8919,N_7826,N_7721);
nand U8920 (N_8920,N_7580,N_7647);
or U8921 (N_8921,N_7524,N_7737);
and U8922 (N_8922,N_7984,N_7919);
xor U8923 (N_8923,N_7334,N_7809);
nand U8924 (N_8924,N_7174,N_7948);
and U8925 (N_8925,N_7145,N_7808);
nand U8926 (N_8926,N_7384,N_7455);
nand U8927 (N_8927,N_7039,N_7929);
or U8928 (N_8928,N_7392,N_7277);
nor U8929 (N_8929,N_7115,N_7446);
or U8930 (N_8930,N_7225,N_7567);
or U8931 (N_8931,N_7269,N_7615);
nand U8932 (N_8932,N_7824,N_7334);
nor U8933 (N_8933,N_7915,N_7969);
nand U8934 (N_8934,N_7175,N_7084);
nand U8935 (N_8935,N_7749,N_7837);
nand U8936 (N_8936,N_7752,N_7415);
nand U8937 (N_8937,N_7346,N_7375);
nand U8938 (N_8938,N_7460,N_7754);
or U8939 (N_8939,N_7674,N_7924);
and U8940 (N_8940,N_7611,N_7035);
and U8941 (N_8941,N_7568,N_7981);
or U8942 (N_8942,N_7292,N_7642);
and U8943 (N_8943,N_7903,N_7984);
nand U8944 (N_8944,N_7988,N_7043);
and U8945 (N_8945,N_7266,N_7023);
or U8946 (N_8946,N_7542,N_7972);
and U8947 (N_8947,N_7846,N_7625);
nand U8948 (N_8948,N_7102,N_7032);
nor U8949 (N_8949,N_7959,N_7565);
nand U8950 (N_8950,N_7692,N_7232);
or U8951 (N_8951,N_7716,N_7419);
or U8952 (N_8952,N_7027,N_7786);
or U8953 (N_8953,N_7082,N_7507);
nor U8954 (N_8954,N_7415,N_7610);
nand U8955 (N_8955,N_7352,N_7264);
xnor U8956 (N_8956,N_7007,N_7542);
or U8957 (N_8957,N_7522,N_7942);
or U8958 (N_8958,N_7774,N_7457);
and U8959 (N_8959,N_7025,N_7335);
nand U8960 (N_8960,N_7499,N_7254);
nor U8961 (N_8961,N_7668,N_7285);
nand U8962 (N_8962,N_7979,N_7481);
nand U8963 (N_8963,N_7967,N_7714);
and U8964 (N_8964,N_7438,N_7861);
nor U8965 (N_8965,N_7061,N_7146);
and U8966 (N_8966,N_7040,N_7765);
and U8967 (N_8967,N_7831,N_7739);
xnor U8968 (N_8968,N_7757,N_7444);
and U8969 (N_8969,N_7588,N_7620);
nor U8970 (N_8970,N_7064,N_7382);
nand U8971 (N_8971,N_7574,N_7500);
and U8972 (N_8972,N_7382,N_7532);
nand U8973 (N_8973,N_7380,N_7412);
and U8974 (N_8974,N_7286,N_7012);
and U8975 (N_8975,N_7897,N_7018);
and U8976 (N_8976,N_7449,N_7890);
nor U8977 (N_8977,N_7263,N_7266);
nand U8978 (N_8978,N_7795,N_7558);
and U8979 (N_8979,N_7559,N_7445);
and U8980 (N_8980,N_7357,N_7704);
nand U8981 (N_8981,N_7961,N_7343);
nand U8982 (N_8982,N_7708,N_7409);
or U8983 (N_8983,N_7103,N_7646);
and U8984 (N_8984,N_7503,N_7890);
or U8985 (N_8985,N_7866,N_7136);
and U8986 (N_8986,N_7701,N_7835);
nand U8987 (N_8987,N_7125,N_7286);
and U8988 (N_8988,N_7165,N_7293);
or U8989 (N_8989,N_7029,N_7010);
nand U8990 (N_8990,N_7345,N_7615);
nor U8991 (N_8991,N_7911,N_7100);
nand U8992 (N_8992,N_7077,N_7809);
nor U8993 (N_8993,N_7480,N_7516);
or U8994 (N_8994,N_7625,N_7776);
and U8995 (N_8995,N_7788,N_7016);
and U8996 (N_8996,N_7133,N_7010);
and U8997 (N_8997,N_7626,N_7859);
or U8998 (N_8998,N_7331,N_7637);
nor U8999 (N_8999,N_7084,N_7627);
and U9000 (N_9000,N_8721,N_8607);
and U9001 (N_9001,N_8844,N_8812);
and U9002 (N_9002,N_8738,N_8839);
and U9003 (N_9003,N_8060,N_8313);
and U9004 (N_9004,N_8637,N_8981);
nand U9005 (N_9005,N_8535,N_8476);
nand U9006 (N_9006,N_8337,N_8222);
and U9007 (N_9007,N_8995,N_8118);
or U9008 (N_9008,N_8251,N_8132);
nand U9009 (N_9009,N_8010,N_8623);
or U9010 (N_9010,N_8194,N_8460);
and U9011 (N_9011,N_8207,N_8979);
and U9012 (N_9012,N_8485,N_8774);
or U9013 (N_9013,N_8677,N_8098);
or U9014 (N_9014,N_8329,N_8365);
nor U9015 (N_9015,N_8937,N_8177);
and U9016 (N_9016,N_8508,N_8260);
nand U9017 (N_9017,N_8775,N_8644);
and U9018 (N_9018,N_8241,N_8656);
nand U9019 (N_9019,N_8032,N_8291);
nand U9020 (N_9020,N_8269,N_8568);
and U9021 (N_9021,N_8469,N_8717);
nor U9022 (N_9022,N_8157,N_8396);
nor U9023 (N_9023,N_8608,N_8987);
nand U9024 (N_9024,N_8148,N_8788);
and U9025 (N_9025,N_8511,N_8614);
nor U9026 (N_9026,N_8997,N_8128);
nor U9027 (N_9027,N_8831,N_8658);
or U9028 (N_9028,N_8472,N_8802);
and U9029 (N_9029,N_8362,N_8678);
or U9030 (N_9030,N_8080,N_8785);
nand U9031 (N_9031,N_8626,N_8601);
xor U9032 (N_9032,N_8254,N_8704);
and U9033 (N_9033,N_8849,N_8063);
and U9034 (N_9034,N_8418,N_8583);
nand U9035 (N_9035,N_8851,N_8605);
nand U9036 (N_9036,N_8682,N_8896);
xor U9037 (N_9037,N_8808,N_8070);
nor U9038 (N_9038,N_8150,N_8083);
and U9039 (N_9039,N_8398,N_8187);
or U9040 (N_9040,N_8878,N_8527);
and U9041 (N_9041,N_8518,N_8430);
or U9042 (N_9042,N_8293,N_8263);
nor U9043 (N_9043,N_8184,N_8671);
and U9044 (N_9044,N_8914,N_8611);
or U9045 (N_9045,N_8809,N_8110);
or U9046 (N_9046,N_8211,N_8749);
or U9047 (N_9047,N_8922,N_8127);
xnor U9048 (N_9048,N_8426,N_8821);
xnor U9049 (N_9049,N_8624,N_8765);
nand U9050 (N_9050,N_8636,N_8968);
nor U9051 (N_9051,N_8019,N_8027);
xor U9052 (N_9052,N_8546,N_8415);
xnor U9053 (N_9053,N_8510,N_8570);
nand U9054 (N_9054,N_8845,N_8784);
nand U9055 (N_9055,N_8331,N_8308);
nor U9056 (N_9056,N_8431,N_8227);
or U9057 (N_9057,N_8092,N_8627);
xor U9058 (N_9058,N_8755,N_8996);
xnor U9059 (N_9059,N_8304,N_8631);
nor U9060 (N_9060,N_8742,N_8971);
and U9061 (N_9061,N_8911,N_8370);
nand U9062 (N_9062,N_8531,N_8423);
or U9063 (N_9063,N_8692,N_8635);
and U9064 (N_9064,N_8154,N_8200);
xor U9065 (N_9065,N_8035,N_8892);
and U9066 (N_9066,N_8556,N_8554);
and U9067 (N_9067,N_8314,N_8078);
xor U9068 (N_9068,N_8284,N_8970);
xnor U9069 (N_9069,N_8593,N_8377);
or U9070 (N_9070,N_8223,N_8838);
nor U9071 (N_9071,N_8668,N_8203);
xor U9072 (N_9072,N_8847,N_8158);
nand U9073 (N_9073,N_8218,N_8443);
or U9074 (N_9074,N_8512,N_8901);
or U9075 (N_9075,N_8822,N_8862);
or U9076 (N_9076,N_8082,N_8836);
and U9077 (N_9077,N_8024,N_8983);
nor U9078 (N_9078,N_8800,N_8230);
or U9079 (N_9079,N_8694,N_8909);
and U9080 (N_9080,N_8735,N_8366);
or U9081 (N_9081,N_8830,N_8869);
or U9082 (N_9082,N_8523,N_8950);
nand U9083 (N_9083,N_8445,N_8016);
nor U9084 (N_9084,N_8501,N_8872);
nor U9085 (N_9085,N_8720,N_8375);
and U9086 (N_9086,N_8710,N_8382);
nor U9087 (N_9087,N_8632,N_8724);
and U9088 (N_9088,N_8274,N_8205);
or U9089 (N_9089,N_8815,N_8214);
nor U9090 (N_9090,N_8948,N_8934);
nor U9091 (N_9091,N_8436,N_8379);
and U9092 (N_9092,N_8565,N_8974);
and U9093 (N_9093,N_8544,N_8347);
nand U9094 (N_9094,N_8022,N_8339);
nor U9095 (N_9095,N_8093,N_8966);
and U9096 (N_9096,N_8236,N_8285);
nand U9097 (N_9097,N_8116,N_8622);
nand U9098 (N_9098,N_8219,N_8867);
nand U9099 (N_9099,N_8621,N_8225);
nor U9100 (N_9100,N_8180,N_8553);
nor U9101 (N_9101,N_8868,N_8718);
nand U9102 (N_9102,N_8843,N_8936);
or U9103 (N_9103,N_8770,N_8924);
nand U9104 (N_9104,N_8425,N_8006);
nand U9105 (N_9105,N_8345,N_8505);
nor U9106 (N_9106,N_8902,N_8279);
or U9107 (N_9107,N_8256,N_8871);
and U9108 (N_9108,N_8952,N_8708);
or U9109 (N_9109,N_8108,N_8343);
nand U9110 (N_9110,N_8548,N_8332);
and U9111 (N_9111,N_8486,N_8638);
or U9112 (N_9112,N_8450,N_8072);
nor U9113 (N_9113,N_8360,N_8889);
or U9114 (N_9114,N_8575,N_8156);
or U9115 (N_9115,N_8283,N_8563);
nor U9116 (N_9116,N_8944,N_8767);
nand U9117 (N_9117,N_8569,N_8245);
or U9118 (N_9118,N_8048,N_8517);
nor U9119 (N_9119,N_8780,N_8615);
or U9120 (N_9120,N_8487,N_8349);
or U9121 (N_9121,N_8552,N_8617);
nand U9122 (N_9122,N_8539,N_8679);
or U9123 (N_9123,N_8811,N_8792);
and U9124 (N_9124,N_8044,N_8810);
nand U9125 (N_9125,N_8497,N_8310);
nand U9126 (N_9126,N_8424,N_8904);
xor U9127 (N_9127,N_8324,N_8005);
nand U9128 (N_9128,N_8479,N_8237);
nor U9129 (N_9129,N_8170,N_8858);
nand U9130 (N_9130,N_8100,N_8707);
nand U9131 (N_9131,N_8965,N_8993);
xnor U9132 (N_9132,N_8919,N_8797);
or U9133 (N_9133,N_8212,N_8600);
and U9134 (N_9134,N_8796,N_8561);
or U9135 (N_9135,N_8726,N_8165);
and U9136 (N_9136,N_8325,N_8482);
and U9137 (N_9137,N_8330,N_8294);
or U9138 (N_9138,N_8891,N_8490);
nor U9139 (N_9139,N_8368,N_8232);
xnor U9140 (N_9140,N_8021,N_8265);
or U9141 (N_9141,N_8786,N_8799);
or U9142 (N_9142,N_8238,N_8887);
and U9143 (N_9143,N_8988,N_8103);
nor U9144 (N_9144,N_8580,N_8860);
nand U9145 (N_9145,N_8258,N_8085);
or U9146 (N_9146,N_8712,N_8828);
or U9147 (N_9147,N_8524,N_8586);
or U9148 (N_9148,N_8541,N_8327);
nor U9149 (N_9149,N_8758,N_8226);
or U9150 (N_9150,N_8953,N_8827);
or U9151 (N_9151,N_8233,N_8558);
nand U9152 (N_9152,N_8719,N_8664);
and U9153 (N_9153,N_8645,N_8018);
nor U9154 (N_9154,N_8587,N_8163);
xnor U9155 (N_9155,N_8597,N_8940);
or U9156 (N_9156,N_8807,N_8776);
nor U9157 (N_9157,N_8540,N_8102);
and U9158 (N_9158,N_8649,N_8179);
or U9159 (N_9159,N_8787,N_8897);
or U9160 (N_9160,N_8301,N_8782);
nor U9161 (N_9161,N_8040,N_8903);
or U9162 (N_9162,N_8943,N_8647);
xnor U9163 (N_9163,N_8946,N_8959);
nor U9164 (N_9164,N_8528,N_8521);
or U9165 (N_9165,N_8120,N_8606);
nand U9166 (N_9166,N_8957,N_8088);
nand U9167 (N_9167,N_8857,N_8651);
or U9168 (N_9168,N_8852,N_8898);
xor U9169 (N_9169,N_8772,N_8646);
nor U9170 (N_9170,N_8160,N_8696);
or U9171 (N_9171,N_8198,N_8178);
and U9172 (N_9172,N_8151,N_8659);
nand U9173 (N_9173,N_8727,N_8101);
or U9174 (N_9174,N_8094,N_8318);
or U9175 (N_9175,N_8706,N_8434);
nand U9176 (N_9176,N_8444,N_8967);
and U9177 (N_9177,N_8550,N_8465);
and U9178 (N_9178,N_8419,N_8058);
and U9179 (N_9179,N_8795,N_8473);
nor U9180 (N_9180,N_8817,N_8954);
nor U9181 (N_9181,N_8842,N_8062);
nand U9182 (N_9182,N_8763,N_8984);
nand U9183 (N_9183,N_8920,N_8306);
nand U9184 (N_9184,N_8364,N_8246);
nand U9185 (N_9185,N_8801,N_8240);
and U9186 (N_9186,N_8300,N_8516);
or U9187 (N_9187,N_8725,N_8562);
or U9188 (N_9188,N_8750,N_8991);
nand U9189 (N_9189,N_8863,N_8989);
or U9190 (N_9190,N_8504,N_8939);
nand U9191 (N_9191,N_8388,N_8043);
and U9192 (N_9192,N_8267,N_8147);
and U9193 (N_9193,N_8009,N_8392);
nor U9194 (N_9194,N_8275,N_8894);
nor U9195 (N_9195,N_8104,N_8047);
and U9196 (N_9196,N_8594,N_8503);
or U9197 (N_9197,N_8174,N_8395);
nand U9198 (N_9198,N_8340,N_8754);
and U9199 (N_9199,N_8917,N_8598);
or U9200 (N_9200,N_8357,N_8777);
or U9201 (N_9201,N_8081,N_8689);
or U9202 (N_9202,N_8250,N_8768);
nand U9203 (N_9203,N_8826,N_8816);
xor U9204 (N_9204,N_8404,N_8276);
xor U9205 (N_9205,N_8814,N_8564);
nor U9206 (N_9206,N_8938,N_8945);
and U9207 (N_9207,N_8239,N_8335);
nor U9208 (N_9208,N_8217,N_8411);
nand U9209 (N_9209,N_8462,N_8282);
xnor U9210 (N_9210,N_8176,N_8819);
and U9211 (N_9211,N_8653,N_8931);
and U9212 (N_9212,N_8056,N_8429);
xor U9213 (N_9213,N_8271,N_8206);
or U9214 (N_9214,N_8481,N_8321);
or U9215 (N_9215,N_8378,N_8942);
and U9216 (N_9216,N_8790,N_8123);
and U9217 (N_9217,N_8029,N_8353);
xor U9218 (N_9218,N_8351,N_8915);
and U9219 (N_9219,N_8661,N_8168);
or U9220 (N_9220,N_8138,N_8041);
nor U9221 (N_9221,N_8383,N_8280);
and U9222 (N_9222,N_8264,N_8855);
or U9223 (N_9223,N_8399,N_8574);
nor U9224 (N_9224,N_8309,N_8705);
or U9225 (N_9225,N_8014,N_8665);
or U9226 (N_9226,N_8262,N_8963);
or U9227 (N_9227,N_8397,N_8925);
or U9228 (N_9228,N_8144,N_8055);
nor U9229 (N_9229,N_8195,N_8125);
nand U9230 (N_9230,N_8990,N_8446);
or U9231 (N_9231,N_8259,N_8739);
and U9232 (N_9232,N_8017,N_8305);
nor U9233 (N_9233,N_8380,N_8875);
and U9234 (N_9234,N_8013,N_8912);
xor U9235 (N_9235,N_8393,N_8498);
nor U9236 (N_9236,N_8759,N_8352);
nand U9237 (N_9237,N_8474,N_8648);
and U9238 (N_9238,N_8683,N_8728);
nor U9239 (N_9239,N_8525,N_8723);
and U9240 (N_9240,N_8432,N_8734);
xor U9241 (N_9241,N_8930,N_8804);
nand U9242 (N_9242,N_8573,N_8949);
or U9243 (N_9243,N_8654,N_8191);
nand U9244 (N_9244,N_8192,N_8255);
nand U9245 (N_9245,N_8249,N_8348);
nor U9246 (N_9246,N_8338,N_8376);
and U9247 (N_9247,N_8421,N_8893);
xnor U9248 (N_9248,N_8117,N_8403);
or U9249 (N_9249,N_8449,N_8509);
nor U9250 (N_9250,N_8407,N_8344);
nor U9251 (N_9251,N_8303,N_8175);
nand U9252 (N_9252,N_8038,N_8779);
or U9253 (N_9253,N_8825,N_8015);
xor U9254 (N_9254,N_8698,N_8493);
nor U9255 (N_9255,N_8890,N_8538);
or U9256 (N_9256,N_8112,N_8273);
and U9257 (N_9257,N_8662,N_8134);
or U9258 (N_9258,N_8410,N_8181);
nor U9259 (N_9259,N_8322,N_8935);
and U9260 (N_9260,N_8628,N_8655);
xor U9261 (N_9261,N_8798,N_8408);
and U9262 (N_9262,N_8409,N_8532);
nor U9263 (N_9263,N_8141,N_8559);
and U9264 (N_9264,N_8173,N_8813);
nand U9265 (N_9265,N_8064,N_8715);
nor U9266 (N_9266,N_8923,N_8882);
nand U9267 (N_9267,N_8488,N_8975);
nand U9268 (N_9268,N_8270,N_8876);
and U9269 (N_9269,N_8500,N_8086);
xor U9270 (N_9270,N_8560,N_8302);
nand U9271 (N_9271,N_8139,N_8595);
or U9272 (N_9272,N_8806,N_8278);
nor U9273 (N_9273,N_8188,N_8769);
nand U9274 (N_9274,N_8316,N_8296);
nand U9275 (N_9275,N_8602,N_8166);
nor U9276 (N_9276,N_8859,N_8204);
nor U9277 (N_9277,N_8685,N_8761);
nand U9278 (N_9278,N_8506,N_8248);
or U9279 (N_9279,N_8536,N_8545);
or U9280 (N_9280,N_8167,N_8549);
nor U9281 (N_9281,N_8475,N_8591);
nor U9282 (N_9282,N_8612,N_8744);
and U9283 (N_9283,N_8557,N_8438);
xor U9284 (N_9284,N_8292,N_8287);
nand U9285 (N_9285,N_8592,N_8703);
and U9286 (N_9286,N_8835,N_8652);
nand U9287 (N_9287,N_8840,N_8442);
nor U9288 (N_9288,N_8389,N_8215);
or U9289 (N_9289,N_8642,N_8109);
nand U9290 (N_9290,N_8958,N_8873);
nand U9291 (N_9291,N_8133,N_8566);
nor U9292 (N_9292,N_8386,N_8477);
nor U9293 (N_9293,N_8046,N_8663);
and U9294 (N_9294,N_8781,N_8803);
nand U9295 (N_9295,N_8709,N_8733);
xor U9296 (N_9296,N_8956,N_8268);
nand U9297 (N_9297,N_8091,N_8417);
or U9298 (N_9298,N_8846,N_8201);
xor U9299 (N_9299,N_8420,N_8307);
and U9300 (N_9300,N_8319,N_8427);
nor U9301 (N_9301,N_8964,N_8590);
or U9302 (N_9302,N_8381,N_8722);
or U9303 (N_9303,N_8688,N_8588);
nor U9304 (N_9304,N_8613,N_8731);
nor U9305 (N_9305,N_8618,N_8695);
xor U9306 (N_9306,N_8115,N_8752);
xnor U9307 (N_9307,N_8850,N_8002);
or U9308 (N_9308,N_8037,N_8281);
nor U9309 (N_9309,N_8910,N_8567);
or U9310 (N_9310,N_8272,N_8519);
or U9311 (N_9311,N_8576,N_8326);
nand U9312 (N_9312,N_8106,N_8155);
nor U9313 (N_9313,N_8162,N_8572);
nand U9314 (N_9314,N_8643,N_8582);
nor U9315 (N_9315,N_8484,N_8589);
nand U9316 (N_9316,N_8084,N_8253);
and U9317 (N_9317,N_8089,N_8702);
nor U9318 (N_9318,N_8447,N_8247);
or U9319 (N_9319,N_8216,N_8478);
nand U9320 (N_9320,N_8153,N_8145);
nor U9321 (N_9321,N_8657,N_8456);
or U9322 (N_9322,N_8122,N_8394);
nor U9323 (N_9323,N_8356,N_8142);
and U9324 (N_9324,N_8457,N_8143);
nor U9325 (N_9325,N_8341,N_8471);
or U9326 (N_9326,N_8877,N_8277);
and U9327 (N_9327,N_8992,N_8824);
nand U9328 (N_9328,N_8669,N_8753);
and U9329 (N_9329,N_8140,N_8054);
or U9330 (N_9330,N_8961,N_8629);
nor U9331 (N_9331,N_8745,N_8856);
or U9332 (N_9332,N_8113,N_8416);
and U9333 (N_9333,N_8320,N_8985);
and U9334 (N_9334,N_8164,N_8794);
xor U9335 (N_9335,N_8412,N_8866);
and U9336 (N_9336,N_8978,N_8619);
or U9337 (N_9337,N_8202,N_8350);
nor U9338 (N_9338,N_8077,N_8371);
or U9339 (N_9339,N_8757,N_8491);
or U9340 (N_9340,N_8713,N_8577);
nor U9341 (N_9341,N_8050,N_8542);
nand U9342 (N_9342,N_8252,N_8700);
nand U9343 (N_9343,N_8905,N_8534);
nor U9344 (N_9344,N_8052,N_8973);
nor U9345 (N_9345,N_8448,N_8955);
or U9346 (N_9346,N_8039,N_8899);
and U9347 (N_9347,N_8455,N_8099);
nor U9348 (N_9348,N_8641,N_8065);
or U9349 (N_9349,N_8960,N_8468);
xor U9350 (N_9350,N_8980,N_8049);
or U9351 (N_9351,N_8414,N_8428);
nand U9352 (N_9352,N_8895,N_8159);
or U9353 (N_9353,N_8927,N_8243);
and U9354 (N_9354,N_8823,N_8684);
or U9355 (N_9355,N_8833,N_8079);
or U9356 (N_9356,N_8235,N_8075);
and U9357 (N_9357,N_8829,N_8069);
or U9358 (N_9358,N_8470,N_8461);
nor U9359 (N_9359,N_8121,N_8464);
nand U9360 (N_9360,N_8437,N_8913);
nand U9361 (N_9361,N_8068,N_8131);
nand U9362 (N_9362,N_8007,N_8762);
nand U9363 (N_9363,N_8401,N_8391);
nor U9364 (N_9364,N_8640,N_8169);
xor U9365 (N_9365,N_8533,N_8756);
nor U9366 (N_9366,N_8452,N_8633);
nor U9367 (N_9367,N_8076,N_8818);
or U9368 (N_9368,N_8136,N_8670);
and U9369 (N_9369,N_8189,N_8361);
nand U9370 (N_9370,N_8224,N_8030);
xnor U9371 (N_9371,N_8172,N_8660);
and U9372 (N_9372,N_8489,N_8832);
or U9373 (N_9373,N_8837,N_8854);
and U9374 (N_9374,N_8231,N_8466);
or U9375 (N_9375,N_8119,N_8515);
nand U9376 (N_9376,N_8881,N_8579);
nor U9377 (N_9377,N_8290,N_8439);
nand U9378 (N_9378,N_8221,N_8028);
nand U9379 (N_9379,N_8625,N_8467);
nor U9380 (N_9380,N_8373,N_8000);
or U9381 (N_9381,N_8741,N_8921);
nor U9382 (N_9382,N_8374,N_8011);
nand U9383 (N_9383,N_8061,N_8666);
nand U9384 (N_9384,N_8096,N_8884);
or U9385 (N_9385,N_8747,N_8982);
and U9386 (N_9386,N_8208,N_8422);
or U9387 (N_9387,N_8585,N_8716);
nor U9388 (N_9388,N_8495,N_8609);
nor U9389 (N_9389,N_8480,N_8193);
and U9390 (N_9390,N_8969,N_8513);
nand U9391 (N_9391,N_8701,N_8630);
and U9392 (N_9392,N_8929,N_8196);
or U9393 (N_9393,N_8778,N_8135);
nor U9394 (N_9394,N_8947,N_8105);
or U9395 (N_9395,N_8051,N_8740);
and U9396 (N_9396,N_8674,N_8530);
nand U9397 (N_9397,N_8385,N_8494);
or U9398 (N_9398,N_8182,N_8916);
nor U9399 (N_9399,N_8673,N_8026);
or U9400 (N_9400,N_8976,N_8888);
or U9401 (N_9401,N_8751,N_8732);
nand U9402 (N_9402,N_8130,N_8186);
or U9403 (N_9403,N_8526,N_8667);
nor U9404 (N_9404,N_8650,N_8358);
nor U9405 (N_9405,N_8286,N_8289);
xor U9406 (N_9406,N_8095,N_8853);
nand U9407 (N_9407,N_8675,N_8315);
xnor U9408 (N_9408,N_8152,N_8620);
or U9409 (N_9409,N_8680,N_8584);
and U9410 (N_9410,N_8886,N_8972);
or U9411 (N_9411,N_8311,N_8336);
nand U9412 (N_9412,N_8406,N_8610);
nand U9413 (N_9413,N_8020,N_8359);
and U9414 (N_9414,N_8220,N_8023);
nor U9415 (N_9415,N_8507,N_8793);
xnor U9416 (N_9416,N_8743,N_8323);
xor U9417 (N_9417,N_8616,N_8870);
nand U9418 (N_9418,N_8190,N_8229);
and U9419 (N_9419,N_8543,N_8864);
xnor U9420 (N_9420,N_8413,N_8736);
and U9421 (N_9421,N_8547,N_8057);
and U9422 (N_9422,N_8841,N_8451);
and U9423 (N_9423,N_8676,N_8071);
nor U9424 (N_9424,N_8791,N_8228);
nand U9425 (N_9425,N_8257,N_8499);
nand U9426 (N_9426,N_8124,N_8333);
and U9427 (N_9427,N_8346,N_8492);
or U9428 (N_9428,N_8687,N_8789);
nor U9429 (N_9429,N_8928,N_8483);
nor U9430 (N_9430,N_8977,N_8213);
nand U9431 (N_9431,N_8234,N_8604);
and U9432 (N_9432,N_8907,N_8578);
or U9433 (N_9433,N_8209,N_8129);
xnor U9434 (N_9434,N_8312,N_8161);
and U9435 (N_9435,N_8885,N_8001);
or U9436 (N_9436,N_8690,N_8355);
or U9437 (N_9437,N_8402,N_8185);
nor U9438 (N_9438,N_8299,N_8691);
and U9439 (N_9439,N_8634,N_8555);
nand U9440 (N_9440,N_8522,N_8760);
or U9441 (N_9441,N_8025,N_8107);
or U9442 (N_9442,N_8087,N_8261);
nor U9443 (N_9443,N_8714,N_8440);
or U9444 (N_9444,N_8454,N_8746);
nor U9445 (N_9445,N_8879,N_8861);
nor U9446 (N_9446,N_8441,N_8183);
nand U9447 (N_9447,N_8639,N_8244);
and U9448 (N_9448,N_8328,N_8697);
nand U9449 (N_9449,N_8369,N_8199);
nor U9450 (N_9450,N_8453,N_8603);
xnor U9451 (N_9451,N_8906,N_8367);
nand U9452 (N_9452,N_8405,N_8883);
or U9453 (N_9453,N_8400,N_8693);
nand U9454 (N_9454,N_8210,N_8334);
and U9455 (N_9455,N_8711,N_8146);
nor U9456 (N_9456,N_8372,N_8880);
nand U9457 (N_9457,N_8596,N_8003);
or U9458 (N_9458,N_8387,N_8520);
xor U9459 (N_9459,N_8834,N_8171);
nor U9460 (N_9460,N_8197,N_8073);
nor U9461 (N_9461,N_8908,N_8433);
or U9462 (N_9462,N_8045,N_8496);
nand U9463 (N_9463,N_8034,N_8012);
or U9464 (N_9464,N_8149,N_8999);
nor U9465 (N_9465,N_8941,N_8900);
or U9466 (N_9466,N_8242,N_8317);
and U9467 (N_9467,N_8004,N_8137);
and U9468 (N_9468,N_8295,N_8551);
nand U9469 (N_9469,N_8042,N_8699);
nor U9470 (N_9470,N_8031,N_8266);
nor U9471 (N_9471,N_8036,N_8059);
or U9472 (N_9472,N_8926,N_8067);
nor U9473 (N_9473,N_8599,N_8994);
nand U9474 (N_9474,N_8288,N_8918);
and U9475 (N_9475,N_8298,N_8463);
or U9476 (N_9476,N_8363,N_8033);
nor U9477 (N_9477,N_8771,N_8773);
or U9478 (N_9478,N_8537,N_8932);
nor U9479 (N_9479,N_8730,N_8053);
nor U9480 (N_9480,N_8514,N_8998);
and U9481 (N_9481,N_8097,N_8342);
or U9482 (N_9482,N_8384,N_8111);
or U9483 (N_9483,N_8008,N_8962);
nor U9484 (N_9484,N_8764,N_8848);
and U9485 (N_9485,N_8581,N_8435);
nor U9486 (N_9486,N_8459,N_8114);
or U9487 (N_9487,N_8951,N_8390);
nand U9488 (N_9488,N_8090,N_8529);
xor U9489 (N_9489,N_8783,N_8986);
or U9490 (N_9490,N_8074,N_8686);
and U9491 (N_9491,N_8354,N_8820);
nand U9492 (N_9492,N_8502,N_8458);
and U9493 (N_9493,N_8066,N_8126);
nor U9494 (N_9494,N_8748,N_8297);
nand U9495 (N_9495,N_8571,N_8874);
nand U9496 (N_9496,N_8805,N_8672);
and U9497 (N_9497,N_8681,N_8933);
nand U9498 (N_9498,N_8729,N_8737);
nand U9499 (N_9499,N_8766,N_8865);
and U9500 (N_9500,N_8923,N_8863);
and U9501 (N_9501,N_8857,N_8731);
nand U9502 (N_9502,N_8281,N_8454);
and U9503 (N_9503,N_8543,N_8328);
nand U9504 (N_9504,N_8555,N_8961);
and U9505 (N_9505,N_8115,N_8355);
nand U9506 (N_9506,N_8900,N_8372);
nand U9507 (N_9507,N_8432,N_8874);
and U9508 (N_9508,N_8616,N_8222);
or U9509 (N_9509,N_8822,N_8123);
nand U9510 (N_9510,N_8666,N_8783);
nand U9511 (N_9511,N_8764,N_8438);
nor U9512 (N_9512,N_8435,N_8788);
nand U9513 (N_9513,N_8425,N_8287);
and U9514 (N_9514,N_8576,N_8374);
nor U9515 (N_9515,N_8520,N_8474);
nor U9516 (N_9516,N_8826,N_8336);
or U9517 (N_9517,N_8459,N_8241);
xor U9518 (N_9518,N_8851,N_8654);
and U9519 (N_9519,N_8139,N_8953);
and U9520 (N_9520,N_8480,N_8282);
or U9521 (N_9521,N_8095,N_8492);
or U9522 (N_9522,N_8410,N_8385);
or U9523 (N_9523,N_8870,N_8318);
nand U9524 (N_9524,N_8317,N_8938);
nand U9525 (N_9525,N_8433,N_8524);
nand U9526 (N_9526,N_8770,N_8463);
xnor U9527 (N_9527,N_8861,N_8636);
and U9528 (N_9528,N_8091,N_8671);
and U9529 (N_9529,N_8483,N_8904);
or U9530 (N_9530,N_8357,N_8058);
and U9531 (N_9531,N_8893,N_8807);
xnor U9532 (N_9532,N_8060,N_8055);
and U9533 (N_9533,N_8970,N_8511);
and U9534 (N_9534,N_8431,N_8758);
xnor U9535 (N_9535,N_8074,N_8694);
or U9536 (N_9536,N_8544,N_8734);
or U9537 (N_9537,N_8908,N_8154);
nor U9538 (N_9538,N_8800,N_8126);
nor U9539 (N_9539,N_8746,N_8598);
or U9540 (N_9540,N_8476,N_8993);
or U9541 (N_9541,N_8064,N_8652);
nor U9542 (N_9542,N_8596,N_8114);
or U9543 (N_9543,N_8063,N_8816);
xnor U9544 (N_9544,N_8628,N_8443);
xnor U9545 (N_9545,N_8078,N_8594);
and U9546 (N_9546,N_8132,N_8598);
nor U9547 (N_9547,N_8400,N_8855);
xor U9548 (N_9548,N_8762,N_8607);
nand U9549 (N_9549,N_8385,N_8313);
nor U9550 (N_9550,N_8179,N_8102);
or U9551 (N_9551,N_8182,N_8840);
and U9552 (N_9552,N_8870,N_8093);
and U9553 (N_9553,N_8029,N_8601);
nand U9554 (N_9554,N_8066,N_8994);
xor U9555 (N_9555,N_8495,N_8361);
and U9556 (N_9556,N_8400,N_8023);
or U9557 (N_9557,N_8579,N_8602);
or U9558 (N_9558,N_8735,N_8147);
and U9559 (N_9559,N_8559,N_8695);
and U9560 (N_9560,N_8402,N_8598);
xnor U9561 (N_9561,N_8797,N_8188);
nand U9562 (N_9562,N_8581,N_8305);
nor U9563 (N_9563,N_8921,N_8824);
nor U9564 (N_9564,N_8379,N_8463);
or U9565 (N_9565,N_8304,N_8994);
and U9566 (N_9566,N_8136,N_8091);
nor U9567 (N_9567,N_8744,N_8681);
or U9568 (N_9568,N_8903,N_8518);
nor U9569 (N_9569,N_8535,N_8486);
nand U9570 (N_9570,N_8189,N_8073);
xnor U9571 (N_9571,N_8433,N_8373);
nand U9572 (N_9572,N_8203,N_8865);
nor U9573 (N_9573,N_8568,N_8778);
nor U9574 (N_9574,N_8876,N_8300);
nand U9575 (N_9575,N_8205,N_8095);
and U9576 (N_9576,N_8873,N_8961);
or U9577 (N_9577,N_8608,N_8994);
nand U9578 (N_9578,N_8874,N_8834);
nand U9579 (N_9579,N_8109,N_8668);
and U9580 (N_9580,N_8690,N_8134);
nor U9581 (N_9581,N_8607,N_8723);
nand U9582 (N_9582,N_8115,N_8859);
or U9583 (N_9583,N_8136,N_8348);
nand U9584 (N_9584,N_8777,N_8196);
or U9585 (N_9585,N_8319,N_8067);
nand U9586 (N_9586,N_8124,N_8306);
or U9587 (N_9587,N_8396,N_8382);
or U9588 (N_9588,N_8320,N_8640);
nor U9589 (N_9589,N_8022,N_8101);
and U9590 (N_9590,N_8927,N_8761);
nor U9591 (N_9591,N_8667,N_8309);
and U9592 (N_9592,N_8934,N_8967);
nand U9593 (N_9593,N_8505,N_8331);
or U9594 (N_9594,N_8347,N_8253);
or U9595 (N_9595,N_8706,N_8982);
nor U9596 (N_9596,N_8840,N_8430);
nor U9597 (N_9597,N_8302,N_8555);
nor U9598 (N_9598,N_8249,N_8204);
nor U9599 (N_9599,N_8639,N_8293);
nor U9600 (N_9600,N_8277,N_8973);
nor U9601 (N_9601,N_8957,N_8832);
nor U9602 (N_9602,N_8378,N_8375);
nor U9603 (N_9603,N_8922,N_8536);
or U9604 (N_9604,N_8452,N_8908);
nor U9605 (N_9605,N_8691,N_8449);
nand U9606 (N_9606,N_8159,N_8725);
and U9607 (N_9607,N_8177,N_8665);
nand U9608 (N_9608,N_8184,N_8971);
xnor U9609 (N_9609,N_8917,N_8781);
or U9610 (N_9610,N_8497,N_8763);
nor U9611 (N_9611,N_8918,N_8974);
and U9612 (N_9612,N_8207,N_8420);
nor U9613 (N_9613,N_8736,N_8981);
nand U9614 (N_9614,N_8220,N_8066);
nand U9615 (N_9615,N_8872,N_8271);
or U9616 (N_9616,N_8003,N_8047);
and U9617 (N_9617,N_8622,N_8606);
nand U9618 (N_9618,N_8551,N_8807);
nor U9619 (N_9619,N_8613,N_8915);
and U9620 (N_9620,N_8550,N_8237);
nand U9621 (N_9621,N_8714,N_8358);
or U9622 (N_9622,N_8228,N_8279);
nand U9623 (N_9623,N_8246,N_8297);
xor U9624 (N_9624,N_8785,N_8044);
nand U9625 (N_9625,N_8739,N_8829);
or U9626 (N_9626,N_8424,N_8262);
nor U9627 (N_9627,N_8559,N_8932);
or U9628 (N_9628,N_8679,N_8838);
nor U9629 (N_9629,N_8779,N_8700);
nand U9630 (N_9630,N_8033,N_8326);
and U9631 (N_9631,N_8472,N_8907);
nand U9632 (N_9632,N_8423,N_8271);
nand U9633 (N_9633,N_8904,N_8371);
and U9634 (N_9634,N_8900,N_8192);
xnor U9635 (N_9635,N_8917,N_8018);
nor U9636 (N_9636,N_8088,N_8116);
nand U9637 (N_9637,N_8103,N_8807);
or U9638 (N_9638,N_8263,N_8873);
or U9639 (N_9639,N_8398,N_8572);
or U9640 (N_9640,N_8709,N_8679);
nand U9641 (N_9641,N_8111,N_8031);
nor U9642 (N_9642,N_8650,N_8563);
nor U9643 (N_9643,N_8061,N_8146);
xnor U9644 (N_9644,N_8573,N_8900);
nand U9645 (N_9645,N_8714,N_8545);
nor U9646 (N_9646,N_8237,N_8742);
or U9647 (N_9647,N_8432,N_8229);
or U9648 (N_9648,N_8292,N_8364);
nor U9649 (N_9649,N_8837,N_8512);
nand U9650 (N_9650,N_8632,N_8535);
nand U9651 (N_9651,N_8345,N_8012);
nor U9652 (N_9652,N_8818,N_8417);
nand U9653 (N_9653,N_8490,N_8631);
and U9654 (N_9654,N_8786,N_8475);
and U9655 (N_9655,N_8760,N_8444);
nor U9656 (N_9656,N_8435,N_8733);
nand U9657 (N_9657,N_8744,N_8664);
and U9658 (N_9658,N_8609,N_8345);
or U9659 (N_9659,N_8239,N_8636);
nand U9660 (N_9660,N_8353,N_8909);
and U9661 (N_9661,N_8174,N_8544);
nor U9662 (N_9662,N_8565,N_8381);
nor U9663 (N_9663,N_8441,N_8603);
and U9664 (N_9664,N_8595,N_8730);
nor U9665 (N_9665,N_8149,N_8389);
nand U9666 (N_9666,N_8122,N_8500);
nand U9667 (N_9667,N_8571,N_8009);
and U9668 (N_9668,N_8515,N_8478);
nor U9669 (N_9669,N_8957,N_8546);
nor U9670 (N_9670,N_8271,N_8325);
xor U9671 (N_9671,N_8573,N_8745);
nor U9672 (N_9672,N_8966,N_8645);
and U9673 (N_9673,N_8853,N_8561);
and U9674 (N_9674,N_8441,N_8515);
and U9675 (N_9675,N_8444,N_8752);
and U9676 (N_9676,N_8154,N_8143);
or U9677 (N_9677,N_8202,N_8849);
and U9678 (N_9678,N_8083,N_8364);
nor U9679 (N_9679,N_8245,N_8300);
and U9680 (N_9680,N_8095,N_8308);
xnor U9681 (N_9681,N_8688,N_8630);
or U9682 (N_9682,N_8427,N_8989);
and U9683 (N_9683,N_8559,N_8321);
or U9684 (N_9684,N_8738,N_8179);
nand U9685 (N_9685,N_8902,N_8395);
nand U9686 (N_9686,N_8483,N_8222);
and U9687 (N_9687,N_8523,N_8602);
nor U9688 (N_9688,N_8039,N_8806);
nor U9689 (N_9689,N_8806,N_8082);
nand U9690 (N_9690,N_8846,N_8024);
or U9691 (N_9691,N_8166,N_8635);
nand U9692 (N_9692,N_8169,N_8518);
xor U9693 (N_9693,N_8377,N_8574);
nand U9694 (N_9694,N_8397,N_8580);
and U9695 (N_9695,N_8311,N_8570);
and U9696 (N_9696,N_8308,N_8588);
nand U9697 (N_9697,N_8939,N_8105);
or U9698 (N_9698,N_8553,N_8240);
and U9699 (N_9699,N_8026,N_8547);
and U9700 (N_9700,N_8941,N_8366);
nor U9701 (N_9701,N_8989,N_8394);
nor U9702 (N_9702,N_8314,N_8597);
nor U9703 (N_9703,N_8213,N_8582);
nor U9704 (N_9704,N_8666,N_8089);
nand U9705 (N_9705,N_8366,N_8352);
nand U9706 (N_9706,N_8426,N_8176);
nor U9707 (N_9707,N_8378,N_8062);
nand U9708 (N_9708,N_8489,N_8902);
or U9709 (N_9709,N_8793,N_8393);
xnor U9710 (N_9710,N_8436,N_8615);
xnor U9711 (N_9711,N_8940,N_8915);
nor U9712 (N_9712,N_8996,N_8137);
and U9713 (N_9713,N_8895,N_8480);
and U9714 (N_9714,N_8544,N_8965);
nor U9715 (N_9715,N_8284,N_8561);
and U9716 (N_9716,N_8035,N_8595);
xor U9717 (N_9717,N_8350,N_8505);
and U9718 (N_9718,N_8617,N_8346);
and U9719 (N_9719,N_8858,N_8359);
nor U9720 (N_9720,N_8877,N_8079);
nor U9721 (N_9721,N_8251,N_8910);
and U9722 (N_9722,N_8730,N_8408);
xnor U9723 (N_9723,N_8187,N_8311);
nor U9724 (N_9724,N_8884,N_8656);
or U9725 (N_9725,N_8536,N_8312);
nor U9726 (N_9726,N_8038,N_8655);
xor U9727 (N_9727,N_8600,N_8763);
and U9728 (N_9728,N_8155,N_8327);
or U9729 (N_9729,N_8990,N_8613);
nor U9730 (N_9730,N_8858,N_8673);
nand U9731 (N_9731,N_8217,N_8387);
or U9732 (N_9732,N_8843,N_8571);
nand U9733 (N_9733,N_8274,N_8661);
nand U9734 (N_9734,N_8755,N_8014);
nand U9735 (N_9735,N_8337,N_8126);
nand U9736 (N_9736,N_8544,N_8389);
and U9737 (N_9737,N_8412,N_8213);
nor U9738 (N_9738,N_8441,N_8381);
nor U9739 (N_9739,N_8093,N_8216);
and U9740 (N_9740,N_8068,N_8004);
nand U9741 (N_9741,N_8337,N_8046);
nand U9742 (N_9742,N_8368,N_8573);
and U9743 (N_9743,N_8083,N_8331);
nand U9744 (N_9744,N_8656,N_8049);
and U9745 (N_9745,N_8067,N_8043);
nor U9746 (N_9746,N_8977,N_8834);
xnor U9747 (N_9747,N_8622,N_8118);
nor U9748 (N_9748,N_8555,N_8725);
or U9749 (N_9749,N_8168,N_8782);
and U9750 (N_9750,N_8085,N_8374);
nor U9751 (N_9751,N_8589,N_8846);
and U9752 (N_9752,N_8156,N_8453);
or U9753 (N_9753,N_8024,N_8961);
and U9754 (N_9754,N_8537,N_8091);
nor U9755 (N_9755,N_8217,N_8416);
or U9756 (N_9756,N_8536,N_8054);
and U9757 (N_9757,N_8725,N_8376);
nor U9758 (N_9758,N_8171,N_8869);
or U9759 (N_9759,N_8784,N_8588);
nor U9760 (N_9760,N_8967,N_8746);
nor U9761 (N_9761,N_8953,N_8713);
or U9762 (N_9762,N_8437,N_8125);
and U9763 (N_9763,N_8738,N_8818);
or U9764 (N_9764,N_8695,N_8004);
nand U9765 (N_9765,N_8285,N_8713);
nor U9766 (N_9766,N_8269,N_8157);
nor U9767 (N_9767,N_8825,N_8937);
or U9768 (N_9768,N_8681,N_8774);
or U9769 (N_9769,N_8753,N_8678);
nor U9770 (N_9770,N_8904,N_8985);
nand U9771 (N_9771,N_8843,N_8382);
and U9772 (N_9772,N_8679,N_8581);
nand U9773 (N_9773,N_8876,N_8093);
or U9774 (N_9774,N_8601,N_8480);
nor U9775 (N_9775,N_8709,N_8553);
nand U9776 (N_9776,N_8307,N_8632);
xor U9777 (N_9777,N_8573,N_8952);
and U9778 (N_9778,N_8877,N_8306);
nand U9779 (N_9779,N_8236,N_8681);
or U9780 (N_9780,N_8601,N_8813);
xor U9781 (N_9781,N_8617,N_8399);
nor U9782 (N_9782,N_8457,N_8377);
or U9783 (N_9783,N_8867,N_8473);
nor U9784 (N_9784,N_8901,N_8070);
or U9785 (N_9785,N_8278,N_8044);
nand U9786 (N_9786,N_8547,N_8584);
and U9787 (N_9787,N_8062,N_8259);
nand U9788 (N_9788,N_8485,N_8066);
xnor U9789 (N_9789,N_8353,N_8344);
and U9790 (N_9790,N_8954,N_8028);
nor U9791 (N_9791,N_8898,N_8801);
nor U9792 (N_9792,N_8242,N_8988);
nor U9793 (N_9793,N_8674,N_8968);
or U9794 (N_9794,N_8391,N_8793);
and U9795 (N_9795,N_8527,N_8194);
nor U9796 (N_9796,N_8892,N_8459);
nand U9797 (N_9797,N_8385,N_8406);
nor U9798 (N_9798,N_8713,N_8164);
nor U9799 (N_9799,N_8366,N_8039);
nand U9800 (N_9800,N_8543,N_8248);
or U9801 (N_9801,N_8308,N_8708);
and U9802 (N_9802,N_8470,N_8242);
nor U9803 (N_9803,N_8614,N_8507);
and U9804 (N_9804,N_8925,N_8430);
and U9805 (N_9805,N_8365,N_8520);
or U9806 (N_9806,N_8765,N_8241);
xor U9807 (N_9807,N_8847,N_8169);
xor U9808 (N_9808,N_8308,N_8741);
nand U9809 (N_9809,N_8213,N_8345);
or U9810 (N_9810,N_8974,N_8819);
nand U9811 (N_9811,N_8727,N_8093);
and U9812 (N_9812,N_8389,N_8911);
nor U9813 (N_9813,N_8198,N_8125);
or U9814 (N_9814,N_8572,N_8274);
nor U9815 (N_9815,N_8355,N_8973);
and U9816 (N_9816,N_8747,N_8858);
and U9817 (N_9817,N_8037,N_8706);
nand U9818 (N_9818,N_8975,N_8047);
nor U9819 (N_9819,N_8057,N_8726);
nor U9820 (N_9820,N_8366,N_8755);
or U9821 (N_9821,N_8005,N_8961);
nor U9822 (N_9822,N_8733,N_8583);
and U9823 (N_9823,N_8859,N_8310);
nor U9824 (N_9824,N_8202,N_8037);
nand U9825 (N_9825,N_8387,N_8137);
xor U9826 (N_9826,N_8154,N_8471);
and U9827 (N_9827,N_8216,N_8413);
nor U9828 (N_9828,N_8917,N_8656);
and U9829 (N_9829,N_8528,N_8774);
nand U9830 (N_9830,N_8066,N_8217);
or U9831 (N_9831,N_8221,N_8001);
nand U9832 (N_9832,N_8160,N_8562);
and U9833 (N_9833,N_8713,N_8645);
nand U9834 (N_9834,N_8624,N_8180);
nor U9835 (N_9835,N_8841,N_8488);
and U9836 (N_9836,N_8651,N_8324);
or U9837 (N_9837,N_8725,N_8495);
nand U9838 (N_9838,N_8914,N_8973);
nand U9839 (N_9839,N_8084,N_8798);
or U9840 (N_9840,N_8273,N_8691);
and U9841 (N_9841,N_8682,N_8762);
xnor U9842 (N_9842,N_8104,N_8061);
or U9843 (N_9843,N_8810,N_8554);
or U9844 (N_9844,N_8166,N_8554);
and U9845 (N_9845,N_8956,N_8963);
nand U9846 (N_9846,N_8733,N_8020);
and U9847 (N_9847,N_8725,N_8585);
and U9848 (N_9848,N_8476,N_8664);
or U9849 (N_9849,N_8298,N_8194);
and U9850 (N_9850,N_8053,N_8427);
xor U9851 (N_9851,N_8647,N_8106);
nand U9852 (N_9852,N_8338,N_8128);
nand U9853 (N_9853,N_8236,N_8322);
nand U9854 (N_9854,N_8530,N_8113);
or U9855 (N_9855,N_8602,N_8365);
nor U9856 (N_9856,N_8448,N_8015);
nor U9857 (N_9857,N_8903,N_8437);
and U9858 (N_9858,N_8724,N_8668);
nor U9859 (N_9859,N_8854,N_8481);
nor U9860 (N_9860,N_8619,N_8108);
nor U9861 (N_9861,N_8044,N_8682);
xnor U9862 (N_9862,N_8616,N_8090);
or U9863 (N_9863,N_8444,N_8120);
nand U9864 (N_9864,N_8995,N_8879);
xnor U9865 (N_9865,N_8533,N_8164);
nor U9866 (N_9866,N_8974,N_8355);
nand U9867 (N_9867,N_8057,N_8280);
nand U9868 (N_9868,N_8005,N_8686);
xnor U9869 (N_9869,N_8128,N_8819);
nand U9870 (N_9870,N_8245,N_8054);
nor U9871 (N_9871,N_8189,N_8278);
and U9872 (N_9872,N_8979,N_8792);
or U9873 (N_9873,N_8971,N_8596);
nor U9874 (N_9874,N_8423,N_8109);
and U9875 (N_9875,N_8501,N_8395);
nand U9876 (N_9876,N_8611,N_8898);
nand U9877 (N_9877,N_8215,N_8296);
and U9878 (N_9878,N_8635,N_8934);
or U9879 (N_9879,N_8983,N_8497);
and U9880 (N_9880,N_8174,N_8789);
and U9881 (N_9881,N_8144,N_8506);
and U9882 (N_9882,N_8578,N_8613);
and U9883 (N_9883,N_8476,N_8061);
nand U9884 (N_9884,N_8988,N_8105);
and U9885 (N_9885,N_8141,N_8935);
nor U9886 (N_9886,N_8842,N_8789);
or U9887 (N_9887,N_8712,N_8897);
and U9888 (N_9888,N_8875,N_8478);
or U9889 (N_9889,N_8614,N_8008);
nand U9890 (N_9890,N_8523,N_8135);
and U9891 (N_9891,N_8291,N_8847);
nand U9892 (N_9892,N_8866,N_8497);
and U9893 (N_9893,N_8214,N_8595);
or U9894 (N_9894,N_8046,N_8585);
nand U9895 (N_9895,N_8181,N_8357);
and U9896 (N_9896,N_8724,N_8156);
or U9897 (N_9897,N_8703,N_8387);
nor U9898 (N_9898,N_8930,N_8602);
xnor U9899 (N_9899,N_8292,N_8298);
and U9900 (N_9900,N_8988,N_8655);
and U9901 (N_9901,N_8389,N_8379);
or U9902 (N_9902,N_8533,N_8451);
xor U9903 (N_9903,N_8117,N_8806);
or U9904 (N_9904,N_8302,N_8181);
or U9905 (N_9905,N_8867,N_8974);
and U9906 (N_9906,N_8053,N_8657);
nand U9907 (N_9907,N_8331,N_8882);
or U9908 (N_9908,N_8709,N_8159);
nand U9909 (N_9909,N_8898,N_8790);
or U9910 (N_9910,N_8803,N_8736);
or U9911 (N_9911,N_8688,N_8966);
nand U9912 (N_9912,N_8039,N_8560);
nand U9913 (N_9913,N_8937,N_8527);
nor U9914 (N_9914,N_8331,N_8220);
nor U9915 (N_9915,N_8225,N_8973);
nand U9916 (N_9916,N_8394,N_8222);
xnor U9917 (N_9917,N_8532,N_8399);
nand U9918 (N_9918,N_8861,N_8543);
nor U9919 (N_9919,N_8584,N_8148);
and U9920 (N_9920,N_8001,N_8350);
xnor U9921 (N_9921,N_8985,N_8038);
and U9922 (N_9922,N_8607,N_8437);
and U9923 (N_9923,N_8502,N_8550);
and U9924 (N_9924,N_8055,N_8198);
nand U9925 (N_9925,N_8791,N_8736);
and U9926 (N_9926,N_8569,N_8865);
nor U9927 (N_9927,N_8994,N_8773);
nor U9928 (N_9928,N_8646,N_8927);
or U9929 (N_9929,N_8504,N_8069);
nand U9930 (N_9930,N_8701,N_8602);
nor U9931 (N_9931,N_8508,N_8897);
nor U9932 (N_9932,N_8150,N_8971);
and U9933 (N_9933,N_8824,N_8388);
or U9934 (N_9934,N_8065,N_8723);
nand U9935 (N_9935,N_8706,N_8735);
and U9936 (N_9936,N_8574,N_8566);
and U9937 (N_9937,N_8841,N_8232);
xnor U9938 (N_9938,N_8824,N_8547);
or U9939 (N_9939,N_8755,N_8074);
or U9940 (N_9940,N_8016,N_8496);
and U9941 (N_9941,N_8595,N_8106);
xor U9942 (N_9942,N_8896,N_8153);
or U9943 (N_9943,N_8198,N_8879);
or U9944 (N_9944,N_8252,N_8429);
and U9945 (N_9945,N_8818,N_8500);
or U9946 (N_9946,N_8453,N_8429);
or U9947 (N_9947,N_8431,N_8888);
and U9948 (N_9948,N_8961,N_8437);
or U9949 (N_9949,N_8854,N_8610);
or U9950 (N_9950,N_8739,N_8135);
or U9951 (N_9951,N_8357,N_8258);
nand U9952 (N_9952,N_8048,N_8749);
and U9953 (N_9953,N_8688,N_8683);
nor U9954 (N_9954,N_8480,N_8772);
nor U9955 (N_9955,N_8873,N_8217);
or U9956 (N_9956,N_8776,N_8304);
nand U9957 (N_9957,N_8817,N_8071);
nor U9958 (N_9958,N_8069,N_8111);
nor U9959 (N_9959,N_8634,N_8866);
and U9960 (N_9960,N_8754,N_8825);
and U9961 (N_9961,N_8160,N_8922);
xnor U9962 (N_9962,N_8128,N_8943);
or U9963 (N_9963,N_8058,N_8807);
or U9964 (N_9964,N_8352,N_8806);
nand U9965 (N_9965,N_8564,N_8551);
and U9966 (N_9966,N_8925,N_8917);
and U9967 (N_9967,N_8869,N_8982);
nand U9968 (N_9968,N_8475,N_8370);
or U9969 (N_9969,N_8688,N_8821);
nor U9970 (N_9970,N_8627,N_8657);
nor U9971 (N_9971,N_8198,N_8826);
nand U9972 (N_9972,N_8099,N_8333);
nor U9973 (N_9973,N_8190,N_8116);
nor U9974 (N_9974,N_8306,N_8154);
nand U9975 (N_9975,N_8693,N_8103);
and U9976 (N_9976,N_8526,N_8406);
nand U9977 (N_9977,N_8111,N_8011);
nand U9978 (N_9978,N_8597,N_8041);
and U9979 (N_9979,N_8514,N_8627);
or U9980 (N_9980,N_8052,N_8389);
and U9981 (N_9981,N_8944,N_8887);
nor U9982 (N_9982,N_8174,N_8163);
xnor U9983 (N_9983,N_8944,N_8884);
nand U9984 (N_9984,N_8617,N_8314);
or U9985 (N_9985,N_8538,N_8448);
nand U9986 (N_9986,N_8171,N_8463);
nor U9987 (N_9987,N_8906,N_8792);
nand U9988 (N_9988,N_8111,N_8432);
xor U9989 (N_9989,N_8836,N_8736);
or U9990 (N_9990,N_8433,N_8985);
nor U9991 (N_9991,N_8847,N_8313);
nor U9992 (N_9992,N_8415,N_8088);
nor U9993 (N_9993,N_8791,N_8658);
or U9994 (N_9994,N_8175,N_8004);
nor U9995 (N_9995,N_8823,N_8596);
nor U9996 (N_9996,N_8631,N_8052);
or U9997 (N_9997,N_8040,N_8397);
and U9998 (N_9998,N_8011,N_8449);
and U9999 (N_9999,N_8788,N_8983);
nand UO_0 (O_0,N_9029,N_9264);
nor UO_1 (O_1,N_9026,N_9866);
or UO_2 (O_2,N_9142,N_9967);
or UO_3 (O_3,N_9711,N_9310);
nand UO_4 (O_4,N_9621,N_9020);
nor UO_5 (O_5,N_9609,N_9728);
nand UO_6 (O_6,N_9038,N_9601);
nor UO_7 (O_7,N_9856,N_9002);
nand UO_8 (O_8,N_9559,N_9778);
xnor UO_9 (O_9,N_9780,N_9137);
xor UO_10 (O_10,N_9753,N_9152);
and UO_11 (O_11,N_9391,N_9108);
and UO_12 (O_12,N_9755,N_9471);
nor UO_13 (O_13,N_9763,N_9915);
or UO_14 (O_14,N_9092,N_9881);
or UO_15 (O_15,N_9147,N_9999);
or UO_16 (O_16,N_9634,N_9258);
nand UO_17 (O_17,N_9416,N_9618);
nor UO_18 (O_18,N_9082,N_9031);
nor UO_19 (O_19,N_9454,N_9675);
or UO_20 (O_20,N_9143,N_9247);
and UO_21 (O_21,N_9931,N_9328);
or UO_22 (O_22,N_9470,N_9798);
and UO_23 (O_23,N_9629,N_9498);
and UO_24 (O_24,N_9012,N_9420);
nand UO_25 (O_25,N_9380,N_9864);
xor UO_26 (O_26,N_9637,N_9397);
and UO_27 (O_27,N_9648,N_9669);
or UO_28 (O_28,N_9992,N_9684);
nand UO_29 (O_29,N_9099,N_9894);
nor UO_30 (O_30,N_9890,N_9001);
xnor UO_31 (O_31,N_9878,N_9988);
nor UO_32 (O_32,N_9412,N_9117);
nand UO_33 (O_33,N_9487,N_9510);
nand UO_34 (O_34,N_9751,N_9485);
or UO_35 (O_35,N_9549,N_9954);
and UO_36 (O_36,N_9814,N_9696);
and UO_37 (O_37,N_9209,N_9922);
nand UO_38 (O_38,N_9379,N_9333);
nor UO_39 (O_39,N_9784,N_9960);
nor UO_40 (O_40,N_9278,N_9052);
and UO_41 (O_41,N_9032,N_9804);
nand UO_42 (O_42,N_9821,N_9500);
nor UO_43 (O_43,N_9886,N_9920);
or UO_44 (O_44,N_9522,N_9065);
nor UO_45 (O_45,N_9961,N_9795);
nand UO_46 (O_46,N_9885,N_9519);
nor UO_47 (O_47,N_9847,N_9906);
and UO_48 (O_48,N_9055,N_9749);
nor UO_49 (O_49,N_9912,N_9168);
and UO_50 (O_50,N_9913,N_9187);
nor UO_51 (O_51,N_9255,N_9827);
nor UO_52 (O_52,N_9641,N_9647);
or UO_53 (O_53,N_9970,N_9895);
nand UO_54 (O_54,N_9315,N_9517);
or UO_55 (O_55,N_9323,N_9865);
nand UO_56 (O_56,N_9893,N_9724);
nor UO_57 (O_57,N_9713,N_9857);
nand UO_58 (O_58,N_9456,N_9443);
or UO_59 (O_59,N_9750,N_9721);
nor UO_60 (O_60,N_9241,N_9617);
xnor UO_61 (O_61,N_9119,N_9439);
nand UO_62 (O_62,N_9263,N_9844);
nor UO_63 (O_63,N_9146,N_9574);
and UO_64 (O_64,N_9271,N_9321);
or UO_65 (O_65,N_9158,N_9593);
or UO_66 (O_66,N_9174,N_9056);
nor UO_67 (O_67,N_9446,N_9435);
or UO_68 (O_68,N_9688,N_9624);
xor UO_69 (O_69,N_9178,N_9937);
xor UO_70 (O_70,N_9276,N_9503);
nor UO_71 (O_71,N_9171,N_9126);
nor UO_72 (O_72,N_9006,N_9058);
and UO_73 (O_73,N_9793,N_9909);
and UO_74 (O_74,N_9025,N_9434);
or UO_75 (O_75,N_9741,N_9662);
nand UO_76 (O_76,N_9576,N_9338);
xor UO_77 (O_77,N_9562,N_9855);
or UO_78 (O_78,N_9692,N_9017);
xnor UO_79 (O_79,N_9768,N_9156);
and UO_80 (O_80,N_9800,N_9473);
or UO_81 (O_81,N_9375,N_9650);
or UO_82 (O_82,N_9387,N_9910);
and UO_83 (O_83,N_9404,N_9494);
or UO_84 (O_84,N_9794,N_9395);
or UO_85 (O_85,N_9851,N_9513);
xnor UO_86 (O_86,N_9488,N_9744);
nand UO_87 (O_87,N_9016,N_9054);
xor UO_88 (O_88,N_9845,N_9983);
nor UO_89 (O_89,N_9709,N_9578);
and UO_90 (O_90,N_9125,N_9467);
nand UO_91 (O_91,N_9537,N_9401);
xor UO_92 (O_92,N_9291,N_9093);
nor UO_93 (O_93,N_9548,N_9036);
nand UO_94 (O_94,N_9840,N_9437);
or UO_95 (O_95,N_9973,N_9293);
or UO_96 (O_96,N_9616,N_9767);
or UO_97 (O_97,N_9850,N_9468);
nand UO_98 (O_98,N_9072,N_9431);
xnor UO_99 (O_99,N_9925,N_9674);
nand UO_100 (O_100,N_9859,N_9600);
xnor UO_101 (O_101,N_9378,N_9237);
nand UO_102 (O_102,N_9489,N_9832);
nor UO_103 (O_103,N_9927,N_9120);
or UO_104 (O_104,N_9421,N_9346);
or UO_105 (O_105,N_9889,N_9694);
nor UO_106 (O_106,N_9207,N_9245);
nand UO_107 (O_107,N_9875,N_9114);
and UO_108 (O_108,N_9294,N_9341);
nand UO_109 (O_109,N_9729,N_9136);
nand UO_110 (O_110,N_9971,N_9936);
and UO_111 (O_111,N_9560,N_9105);
and UO_112 (O_112,N_9884,N_9951);
xnor UO_113 (O_113,N_9332,N_9279);
nand UO_114 (O_114,N_9415,N_9861);
and UO_115 (O_115,N_9660,N_9450);
nand UO_116 (O_116,N_9004,N_9789);
or UO_117 (O_117,N_9769,N_9993);
and UO_118 (O_118,N_9631,N_9196);
and UO_119 (O_119,N_9710,N_9632);
xor UO_120 (O_120,N_9705,N_9934);
xor UO_121 (O_121,N_9259,N_9563);
nand UO_122 (O_122,N_9852,N_9235);
nor UO_123 (O_123,N_9290,N_9281);
nand UO_124 (O_124,N_9250,N_9667);
or UO_125 (O_125,N_9273,N_9796);
xnor UO_126 (O_126,N_9256,N_9656);
and UO_127 (O_127,N_9356,N_9981);
or UO_128 (O_128,N_9022,N_9722);
or UO_129 (O_129,N_9687,N_9766);
nand UO_130 (O_130,N_9530,N_9217);
nand UO_131 (O_131,N_9015,N_9862);
xnor UO_132 (O_132,N_9540,N_9314);
and UO_133 (O_133,N_9797,N_9090);
nand UO_134 (O_134,N_9475,N_9203);
and UO_135 (O_135,N_9402,N_9324);
or UO_136 (O_136,N_9063,N_9413);
nor UO_137 (O_137,N_9045,N_9773);
and UO_138 (O_138,N_9484,N_9752);
or UO_139 (O_139,N_9996,N_9892);
and UO_140 (O_140,N_9502,N_9130);
xnor UO_141 (O_141,N_9390,N_9389);
or UO_142 (O_142,N_9206,N_9677);
and UO_143 (O_143,N_9010,N_9896);
nand UO_144 (O_144,N_9730,N_9699);
and UO_145 (O_145,N_9633,N_9451);
xnor UO_146 (O_146,N_9067,N_9940);
and UO_147 (O_147,N_9027,N_9115);
nor UO_148 (O_148,N_9811,N_9614);
and UO_149 (O_149,N_9316,N_9939);
and UO_150 (O_150,N_9670,N_9715);
and UO_151 (O_151,N_9625,N_9101);
and UO_152 (O_152,N_9620,N_9095);
nand UO_153 (O_153,N_9430,N_9700);
xnor UO_154 (O_154,N_9400,N_9693);
nor UO_155 (O_155,N_9266,N_9159);
nand UO_156 (O_156,N_9636,N_9702);
nand UO_157 (O_157,N_9239,N_9643);
nand UO_158 (O_158,N_9304,N_9745);
and UO_159 (O_159,N_9311,N_9664);
nor UO_160 (O_160,N_9268,N_9057);
nand UO_161 (O_161,N_9571,N_9331);
or UO_162 (O_162,N_9364,N_9816);
nor UO_163 (O_163,N_9596,N_9841);
and UO_164 (O_164,N_9373,N_9867);
and UO_165 (O_165,N_9193,N_9757);
and UO_166 (O_166,N_9444,N_9575);
nand UO_167 (O_167,N_9077,N_9371);
or UO_168 (O_168,N_9595,N_9976);
and UO_169 (O_169,N_9551,N_9772);
and UO_170 (O_170,N_9528,N_9417);
nor UO_171 (O_171,N_9050,N_9949);
and UO_172 (O_172,N_9732,N_9251);
xor UO_173 (O_173,N_9573,N_9097);
nor UO_174 (O_174,N_9904,N_9781);
xor UO_175 (O_175,N_9465,N_9176);
nor UO_176 (O_176,N_9787,N_9626);
and UO_177 (O_177,N_9288,N_9139);
nand UO_178 (O_178,N_9535,N_9081);
xnor UO_179 (O_179,N_9428,N_9829);
and UO_180 (O_180,N_9028,N_9466);
or UO_181 (O_181,N_9929,N_9948);
nand UO_182 (O_182,N_9189,N_9384);
xor UO_183 (O_183,N_9989,N_9381);
or UO_184 (O_184,N_9926,N_9822);
or UO_185 (O_185,N_9007,N_9561);
and UO_186 (O_186,N_9403,N_9672);
nand UO_187 (O_187,N_9162,N_9376);
nor UO_188 (O_188,N_9083,N_9828);
or UO_189 (O_189,N_9123,N_9018);
and UO_190 (O_190,N_9351,N_9570);
nand UO_191 (O_191,N_9938,N_9112);
nor UO_192 (O_192,N_9111,N_9785);
nor UO_193 (O_193,N_9349,N_9572);
or UO_194 (O_194,N_9270,N_9908);
and UO_195 (O_195,N_9707,N_9813);
and UO_196 (O_196,N_9935,N_9405);
nand UO_197 (O_197,N_9833,N_9900);
or UO_198 (O_198,N_9374,N_9586);
and UO_199 (O_199,N_9429,N_9598);
xnor UO_200 (O_200,N_9902,N_9021);
or UO_201 (O_201,N_9542,N_9098);
nor UO_202 (O_202,N_9229,N_9830);
or UO_203 (O_203,N_9491,N_9367);
and UO_204 (O_204,N_9952,N_9887);
nor UO_205 (O_205,N_9966,N_9504);
or UO_206 (O_206,N_9262,N_9213);
or UO_207 (O_207,N_9088,N_9984);
xor UO_208 (O_208,N_9424,N_9658);
nand UO_209 (O_209,N_9426,N_9602);
or UO_210 (O_210,N_9792,N_9044);
or UO_211 (O_211,N_9612,N_9197);
and UO_212 (O_212,N_9652,N_9708);
or UO_213 (O_213,N_9605,N_9226);
or UO_214 (O_214,N_9599,N_9300);
xor UO_215 (O_215,N_9717,N_9326);
xnor UO_216 (O_216,N_9546,N_9898);
nand UO_217 (O_217,N_9165,N_9307);
xnor UO_218 (O_218,N_9282,N_9761);
nand UO_219 (O_219,N_9921,N_9169);
and UO_220 (O_220,N_9383,N_9306);
xor UO_221 (O_221,N_9253,N_9348);
or UO_222 (O_222,N_9950,N_9799);
nand UO_223 (O_223,N_9716,N_9518);
or UO_224 (O_224,N_9547,N_9303);
nor UO_225 (O_225,N_9232,N_9916);
and UO_226 (O_226,N_9355,N_9127);
nand UO_227 (O_227,N_9140,N_9014);
nor UO_228 (O_228,N_9297,N_9287);
nor UO_229 (O_229,N_9877,N_9492);
xor UO_230 (O_230,N_9144,N_9339);
or UO_231 (O_231,N_9541,N_9682);
nor UO_232 (O_232,N_9410,N_9972);
nor UO_233 (O_233,N_9582,N_9726);
nand UO_234 (O_234,N_9298,N_9776);
xnor UO_235 (O_235,N_9539,N_9627);
or UO_236 (O_236,N_9604,N_9924);
and UO_237 (O_237,N_9758,N_9527);
or UO_238 (O_238,N_9953,N_9863);
or UO_239 (O_239,N_9039,N_9414);
and UO_240 (O_240,N_9116,N_9739);
nor UO_241 (O_241,N_9037,N_9923);
nand UO_242 (O_242,N_9132,N_9153);
nor UO_243 (O_243,N_9515,N_9727);
xor UO_244 (O_244,N_9478,N_9087);
xor UO_245 (O_245,N_9385,N_9242);
or UO_246 (O_246,N_9657,N_9812);
or UO_247 (O_247,N_9735,N_9370);
xor UO_248 (O_248,N_9665,N_9536);
or UO_249 (O_249,N_9396,N_9842);
or UO_250 (O_250,N_9393,N_9577);
nor UO_251 (O_251,N_9318,N_9345);
nor UO_252 (O_252,N_9200,N_9228);
and UO_253 (O_253,N_9779,N_9107);
nor UO_254 (O_254,N_9483,N_9312);
or UO_255 (O_255,N_9289,N_9230);
nand UO_256 (O_256,N_9149,N_9918);
nand UO_257 (O_257,N_9532,N_9872);
and UO_258 (O_258,N_9096,N_9283);
or UO_259 (O_259,N_9422,N_9649);
and UO_260 (O_260,N_9868,N_9071);
or UO_261 (O_261,N_9583,N_9580);
nor UO_262 (O_262,N_9630,N_9978);
nand UO_263 (O_263,N_9337,N_9810);
or UO_264 (O_264,N_9914,N_9516);
nand UO_265 (O_265,N_9034,N_9858);
and UO_266 (O_266,N_9698,N_9085);
nand UO_267 (O_267,N_9676,N_9073);
nor UO_268 (O_268,N_9399,N_9286);
nor UO_269 (O_269,N_9673,N_9458);
nor UO_270 (O_270,N_9740,N_9825);
or UO_271 (O_271,N_9334,N_9216);
or UO_272 (O_272,N_9305,N_9481);
nand UO_273 (O_273,N_9181,N_9243);
nand UO_274 (O_274,N_9357,N_9873);
xor UO_275 (O_275,N_9584,N_9445);
nand UO_276 (O_276,N_9308,N_9899);
or UO_277 (O_277,N_9344,N_9313);
and UO_278 (O_278,N_9254,N_9457);
and UO_279 (O_279,N_9322,N_9319);
or UO_280 (O_280,N_9668,N_9023);
nand UO_281 (O_281,N_9267,N_9359);
nor UO_282 (O_282,N_9452,N_9459);
or UO_283 (O_283,N_9809,N_9738);
nand UO_284 (O_284,N_9442,N_9392);
nand UO_285 (O_285,N_9423,N_9671);
nor UO_286 (O_286,N_9060,N_9244);
nor UO_287 (O_287,N_9161,N_9957);
or UO_288 (O_288,N_9712,N_9969);
or UO_289 (O_289,N_9198,N_9523);
xnor UO_290 (O_290,N_9691,N_9008);
nand UO_291 (O_291,N_9104,N_9946);
or UO_292 (O_292,N_9526,N_9432);
nand UO_293 (O_293,N_9447,N_9277);
nand UO_294 (O_294,N_9703,N_9365);
and UO_295 (O_295,N_9803,N_9581);
and UO_296 (O_296,N_9843,N_9167);
xnor UO_297 (O_297,N_9188,N_9565);
nand UO_298 (O_298,N_9645,N_9854);
and UO_299 (O_299,N_9538,N_9463);
xnor UO_300 (O_300,N_9907,N_9497);
and UO_301 (O_301,N_9880,N_9100);
nand UO_302 (O_302,N_9495,N_9275);
or UO_303 (O_303,N_9760,N_9968);
nand UO_304 (O_304,N_9074,N_9553);
nor UO_305 (O_305,N_9474,N_9075);
nand UO_306 (O_306,N_9690,N_9141);
and UO_307 (O_307,N_9603,N_9109);
and UO_308 (O_308,N_9566,N_9876);
or UO_309 (O_309,N_9388,N_9905);
or UO_310 (O_310,N_9009,N_9272);
xor UO_311 (O_311,N_9157,N_9240);
and UO_312 (O_312,N_9639,N_9476);
xnor UO_313 (O_313,N_9680,N_9733);
or UO_314 (O_314,N_9089,N_9587);
or UO_315 (O_315,N_9743,N_9980);
xnor UO_316 (O_316,N_9932,N_9003);
or UO_317 (O_317,N_9041,N_9987);
or UO_318 (O_318,N_9408,N_9122);
nand UO_319 (O_319,N_9653,N_9086);
nand UO_320 (O_320,N_9640,N_9219);
nor UO_321 (O_321,N_9166,N_9775);
or UO_322 (O_322,N_9265,N_9771);
and UO_323 (O_323,N_9945,N_9335);
nor UO_324 (O_324,N_9661,N_9815);
or UO_325 (O_325,N_9871,N_9131);
or UO_326 (O_326,N_9479,N_9774);
or UO_327 (O_327,N_9742,N_9129);
and UO_328 (O_328,N_9106,N_9959);
and UO_329 (O_329,N_9808,N_9802);
nor UO_330 (O_330,N_9078,N_9790);
or UO_331 (O_331,N_9508,N_9301);
or UO_332 (O_332,N_9461,N_9544);
xnor UO_333 (O_333,N_9246,N_9568);
or UO_334 (O_334,N_9706,N_9782);
and UO_335 (O_335,N_9579,N_9685);
nand UO_336 (O_336,N_9531,N_9164);
nor UO_337 (O_337,N_9046,N_9236);
nor UO_338 (O_338,N_9534,N_9511);
nand UO_339 (O_339,N_9982,N_9076);
and UO_340 (O_340,N_9731,N_9848);
nand UO_341 (O_341,N_9084,N_9869);
and UO_342 (O_342,N_9663,N_9411);
nand UO_343 (O_343,N_9192,N_9962);
and UO_344 (O_344,N_9977,N_9897);
and UO_345 (O_345,N_9499,N_9590);
xnor UO_346 (O_346,N_9195,N_9352);
nand UO_347 (O_347,N_9524,N_9386);
and UO_348 (O_348,N_9666,N_9678);
xor UO_349 (O_349,N_9817,N_9933);
or UO_350 (O_350,N_9901,N_9557);
nor UO_351 (O_351,N_9175,N_9831);
or UO_352 (O_352,N_9134,N_9234);
or UO_353 (O_353,N_9490,N_9295);
or UO_354 (O_354,N_9805,N_9062);
nor UO_355 (O_355,N_9550,N_9719);
or UO_356 (O_356,N_9501,N_9151);
nand UO_357 (O_357,N_9190,N_9788);
xor UO_358 (O_358,N_9118,N_9113);
nand UO_359 (O_359,N_9419,N_9718);
and UO_360 (O_360,N_9362,N_9834);
and UO_361 (O_361,N_9043,N_9589);
nor UO_362 (O_362,N_9183,N_9124);
and UO_363 (O_363,N_9194,N_9150);
and UO_364 (O_364,N_9512,N_9746);
and UO_365 (O_365,N_9882,N_9928);
xnor UO_366 (O_366,N_9138,N_9042);
or UO_367 (O_367,N_9606,N_9154);
or UO_368 (O_368,N_9436,N_9836);
nand UO_369 (O_369,N_9615,N_9238);
nand UO_370 (O_370,N_9644,N_9091);
and UO_371 (O_371,N_9064,N_9069);
xnor UO_372 (O_372,N_9398,N_9610);
and UO_373 (O_373,N_9608,N_9363);
and UO_374 (O_374,N_9651,N_9704);
and UO_375 (O_375,N_9051,N_9448);
or UO_376 (O_376,N_9180,N_9853);
and UO_377 (O_377,N_9533,N_9818);
or UO_378 (O_378,N_9019,N_9177);
nor UO_379 (O_379,N_9035,N_9655);
or UO_380 (O_380,N_9786,N_9720);
or UO_381 (O_381,N_9681,N_9472);
or UO_382 (O_382,N_9292,N_9965);
and UO_383 (O_383,N_9879,N_9891);
nor UO_384 (O_384,N_9133,N_9947);
xnor UO_385 (O_385,N_9280,N_9225);
nand UO_386 (O_386,N_9974,N_9358);
or UO_387 (O_387,N_9942,N_9911);
and UO_388 (O_388,N_9068,N_9588);
nand UO_389 (O_389,N_9455,N_9211);
nand UO_390 (O_390,N_9425,N_9135);
xnor UO_391 (O_391,N_9903,N_9683);
and UO_392 (O_392,N_9284,N_9888);
nor UO_393 (O_393,N_9343,N_9317);
nand UO_394 (O_394,N_9201,N_9350);
nor UO_395 (O_395,N_9756,N_9529);
or UO_396 (O_396,N_9342,N_9061);
and UO_397 (O_397,N_9736,N_9214);
nand UO_398 (O_398,N_9994,N_9714);
nor UO_399 (O_399,N_9233,N_9199);
nor UO_400 (O_400,N_9460,N_9000);
nor UO_401 (O_401,N_9642,N_9496);
or UO_402 (O_402,N_9231,N_9347);
and UO_403 (O_403,N_9179,N_9441);
or UO_404 (O_404,N_9520,N_9525);
nand UO_405 (O_405,N_9368,N_9985);
nand UO_406 (O_406,N_9361,N_9257);
nor UO_407 (O_407,N_9543,N_9820);
nand UO_408 (O_408,N_9309,N_9734);
and UO_409 (O_409,N_9269,N_9611);
nor UO_410 (O_410,N_9372,N_9597);
nand UO_411 (O_411,N_9070,N_9964);
nand UO_412 (O_412,N_9747,N_9202);
or UO_413 (O_413,N_9155,N_9623);
xor UO_414 (O_414,N_9215,N_9695);
nor UO_415 (O_415,N_9659,N_9184);
and UO_416 (O_416,N_9569,N_9205);
nand UO_417 (O_417,N_9591,N_9160);
and UO_418 (O_418,N_9066,N_9944);
nor UO_419 (O_419,N_9382,N_9210);
nand UO_420 (O_420,N_9427,N_9482);
and UO_421 (O_421,N_9366,N_9930);
and UO_422 (O_422,N_9329,N_9185);
and UO_423 (O_423,N_9990,N_9837);
and UO_424 (O_424,N_9819,N_9220);
or UO_425 (O_425,N_9564,N_9592);
xnor UO_426 (O_426,N_9594,N_9013);
nor UO_427 (O_427,N_9493,N_9170);
and UO_428 (O_428,N_9725,N_9221);
nand UO_429 (O_429,N_9145,N_9261);
xor UO_430 (O_430,N_9919,N_9218);
xnor UO_431 (O_431,N_9182,N_9340);
nand UO_432 (O_432,N_9754,N_9613);
and UO_433 (O_433,N_9191,N_9701);
or UO_434 (O_434,N_9212,N_9801);
nor UO_435 (O_435,N_9679,N_9148);
or UO_436 (O_436,N_9325,N_9506);
nand UO_437 (O_437,N_9554,N_9330);
xnor UO_438 (O_438,N_9369,N_9354);
nor UO_439 (O_439,N_9998,N_9480);
nor UO_440 (O_440,N_9204,N_9839);
or UO_441 (O_441,N_9469,N_9477);
or UO_442 (O_442,N_9285,N_9824);
or UO_443 (O_443,N_9791,N_9723);
nand UO_444 (O_444,N_9173,N_9505);
and UO_445 (O_445,N_9619,N_9011);
xor UO_446 (O_446,N_9110,N_9509);
or UO_447 (O_447,N_9737,N_9975);
xnor UO_448 (O_448,N_9486,N_9521);
and UO_449 (O_449,N_9208,N_9860);
nor UO_450 (O_450,N_9053,N_9943);
or UO_451 (O_451,N_9260,N_9048);
or UO_452 (O_452,N_9585,N_9849);
xnor UO_453 (O_453,N_9030,N_9222);
xnor UO_454 (O_454,N_9024,N_9555);
nor UO_455 (O_455,N_9759,N_9628);
nand UO_456 (O_456,N_9622,N_9835);
xnor UO_457 (O_457,N_9320,N_9102);
nand UO_458 (O_458,N_9047,N_9080);
and UO_459 (O_459,N_9697,N_9689);
and UO_460 (O_460,N_9360,N_9377);
or UO_461 (O_461,N_9163,N_9449);
nor UO_462 (O_462,N_9224,N_9552);
xor UO_463 (O_463,N_9995,N_9248);
nand UO_464 (O_464,N_9353,N_9991);
nand UO_465 (O_465,N_9186,N_9327);
nor UO_466 (O_466,N_9252,N_9846);
nand UO_467 (O_467,N_9997,N_9986);
or UO_468 (O_468,N_9764,N_9545);
or UO_469 (O_469,N_9963,N_9956);
xnor UO_470 (O_470,N_9917,N_9433);
or UO_471 (O_471,N_9223,N_9005);
nor UO_472 (O_472,N_9059,N_9040);
xnor UO_473 (O_473,N_9409,N_9955);
xor UO_474 (O_474,N_9299,N_9826);
and UO_475 (O_475,N_9638,N_9121);
or UO_476 (O_476,N_9783,N_9249);
nand UO_477 (O_477,N_9128,N_9103);
or UO_478 (O_478,N_9838,N_9806);
and UO_479 (O_479,N_9394,N_9646);
nand UO_480 (O_480,N_9336,N_9777);
nor UO_481 (O_481,N_9438,N_9654);
or UO_482 (O_482,N_9958,N_9765);
nand UO_483 (O_483,N_9418,N_9635);
nor UO_484 (O_484,N_9507,N_9686);
and UO_485 (O_485,N_9440,N_9941);
nor UO_486 (O_486,N_9407,N_9453);
or UO_487 (O_487,N_9874,N_9274);
and UO_488 (O_488,N_9807,N_9823);
or UO_489 (O_489,N_9770,N_9464);
xor UO_490 (O_490,N_9870,N_9748);
xor UO_491 (O_491,N_9172,N_9979);
or UO_492 (O_492,N_9049,N_9514);
and UO_493 (O_493,N_9033,N_9302);
nor UO_494 (O_494,N_9094,N_9079);
or UO_495 (O_495,N_9607,N_9406);
or UO_496 (O_496,N_9296,N_9883);
xor UO_497 (O_497,N_9227,N_9762);
xor UO_498 (O_498,N_9462,N_9567);
or UO_499 (O_499,N_9558,N_9556);
nor UO_500 (O_500,N_9719,N_9516);
and UO_501 (O_501,N_9403,N_9997);
xnor UO_502 (O_502,N_9780,N_9265);
xor UO_503 (O_503,N_9153,N_9804);
and UO_504 (O_504,N_9072,N_9125);
xor UO_505 (O_505,N_9178,N_9814);
or UO_506 (O_506,N_9616,N_9013);
and UO_507 (O_507,N_9264,N_9880);
nand UO_508 (O_508,N_9041,N_9702);
or UO_509 (O_509,N_9933,N_9940);
nor UO_510 (O_510,N_9651,N_9117);
xnor UO_511 (O_511,N_9672,N_9392);
or UO_512 (O_512,N_9682,N_9478);
nand UO_513 (O_513,N_9926,N_9374);
or UO_514 (O_514,N_9975,N_9167);
or UO_515 (O_515,N_9581,N_9201);
nor UO_516 (O_516,N_9020,N_9780);
and UO_517 (O_517,N_9268,N_9824);
xnor UO_518 (O_518,N_9458,N_9626);
or UO_519 (O_519,N_9191,N_9525);
nor UO_520 (O_520,N_9672,N_9810);
or UO_521 (O_521,N_9308,N_9499);
nor UO_522 (O_522,N_9369,N_9295);
nand UO_523 (O_523,N_9376,N_9398);
or UO_524 (O_524,N_9600,N_9109);
nor UO_525 (O_525,N_9263,N_9900);
nor UO_526 (O_526,N_9534,N_9540);
or UO_527 (O_527,N_9970,N_9552);
nor UO_528 (O_528,N_9562,N_9233);
nand UO_529 (O_529,N_9953,N_9944);
nand UO_530 (O_530,N_9449,N_9876);
nor UO_531 (O_531,N_9933,N_9582);
or UO_532 (O_532,N_9726,N_9959);
xnor UO_533 (O_533,N_9556,N_9915);
and UO_534 (O_534,N_9282,N_9597);
and UO_535 (O_535,N_9677,N_9704);
and UO_536 (O_536,N_9387,N_9005);
xor UO_537 (O_537,N_9036,N_9451);
and UO_538 (O_538,N_9922,N_9294);
and UO_539 (O_539,N_9539,N_9021);
nor UO_540 (O_540,N_9266,N_9010);
nand UO_541 (O_541,N_9167,N_9519);
nand UO_542 (O_542,N_9630,N_9941);
nor UO_543 (O_543,N_9372,N_9699);
nor UO_544 (O_544,N_9382,N_9493);
and UO_545 (O_545,N_9752,N_9679);
nand UO_546 (O_546,N_9203,N_9723);
and UO_547 (O_547,N_9024,N_9627);
or UO_548 (O_548,N_9692,N_9336);
nor UO_549 (O_549,N_9855,N_9269);
nor UO_550 (O_550,N_9919,N_9817);
nor UO_551 (O_551,N_9243,N_9620);
nand UO_552 (O_552,N_9194,N_9226);
nor UO_553 (O_553,N_9264,N_9553);
nor UO_554 (O_554,N_9740,N_9377);
and UO_555 (O_555,N_9967,N_9672);
or UO_556 (O_556,N_9653,N_9699);
nand UO_557 (O_557,N_9429,N_9444);
nor UO_558 (O_558,N_9480,N_9915);
and UO_559 (O_559,N_9277,N_9070);
nand UO_560 (O_560,N_9060,N_9002);
or UO_561 (O_561,N_9170,N_9253);
xor UO_562 (O_562,N_9873,N_9117);
and UO_563 (O_563,N_9600,N_9601);
nand UO_564 (O_564,N_9889,N_9424);
or UO_565 (O_565,N_9977,N_9416);
and UO_566 (O_566,N_9805,N_9553);
nor UO_567 (O_567,N_9976,N_9361);
nor UO_568 (O_568,N_9415,N_9656);
or UO_569 (O_569,N_9578,N_9206);
xnor UO_570 (O_570,N_9673,N_9053);
and UO_571 (O_571,N_9427,N_9688);
nand UO_572 (O_572,N_9856,N_9936);
nand UO_573 (O_573,N_9245,N_9517);
or UO_574 (O_574,N_9438,N_9911);
nand UO_575 (O_575,N_9005,N_9529);
or UO_576 (O_576,N_9324,N_9950);
nand UO_577 (O_577,N_9610,N_9966);
xor UO_578 (O_578,N_9364,N_9611);
nor UO_579 (O_579,N_9562,N_9384);
nand UO_580 (O_580,N_9740,N_9077);
nand UO_581 (O_581,N_9610,N_9938);
and UO_582 (O_582,N_9647,N_9891);
xor UO_583 (O_583,N_9536,N_9332);
and UO_584 (O_584,N_9815,N_9190);
or UO_585 (O_585,N_9058,N_9994);
nor UO_586 (O_586,N_9945,N_9232);
nor UO_587 (O_587,N_9474,N_9318);
or UO_588 (O_588,N_9554,N_9660);
and UO_589 (O_589,N_9147,N_9983);
nor UO_590 (O_590,N_9359,N_9667);
nor UO_591 (O_591,N_9305,N_9988);
nand UO_592 (O_592,N_9916,N_9017);
or UO_593 (O_593,N_9557,N_9142);
xnor UO_594 (O_594,N_9692,N_9624);
and UO_595 (O_595,N_9779,N_9658);
or UO_596 (O_596,N_9297,N_9798);
nor UO_597 (O_597,N_9507,N_9023);
or UO_598 (O_598,N_9840,N_9297);
nand UO_599 (O_599,N_9295,N_9935);
or UO_600 (O_600,N_9854,N_9780);
nor UO_601 (O_601,N_9794,N_9077);
nand UO_602 (O_602,N_9186,N_9819);
or UO_603 (O_603,N_9228,N_9208);
nand UO_604 (O_604,N_9729,N_9408);
nand UO_605 (O_605,N_9457,N_9635);
and UO_606 (O_606,N_9859,N_9136);
nor UO_607 (O_607,N_9985,N_9231);
nor UO_608 (O_608,N_9694,N_9905);
or UO_609 (O_609,N_9218,N_9041);
nor UO_610 (O_610,N_9530,N_9435);
and UO_611 (O_611,N_9154,N_9766);
nand UO_612 (O_612,N_9282,N_9100);
nor UO_613 (O_613,N_9881,N_9446);
nand UO_614 (O_614,N_9511,N_9684);
and UO_615 (O_615,N_9527,N_9374);
or UO_616 (O_616,N_9005,N_9573);
or UO_617 (O_617,N_9750,N_9000);
and UO_618 (O_618,N_9230,N_9638);
and UO_619 (O_619,N_9008,N_9341);
or UO_620 (O_620,N_9442,N_9634);
and UO_621 (O_621,N_9453,N_9692);
and UO_622 (O_622,N_9804,N_9668);
and UO_623 (O_623,N_9394,N_9044);
or UO_624 (O_624,N_9562,N_9580);
nand UO_625 (O_625,N_9679,N_9941);
nand UO_626 (O_626,N_9791,N_9389);
or UO_627 (O_627,N_9172,N_9994);
and UO_628 (O_628,N_9369,N_9550);
nand UO_629 (O_629,N_9393,N_9952);
nor UO_630 (O_630,N_9682,N_9220);
xnor UO_631 (O_631,N_9419,N_9179);
xnor UO_632 (O_632,N_9305,N_9314);
or UO_633 (O_633,N_9711,N_9641);
xor UO_634 (O_634,N_9567,N_9593);
nor UO_635 (O_635,N_9997,N_9184);
nor UO_636 (O_636,N_9462,N_9116);
nor UO_637 (O_637,N_9088,N_9728);
xnor UO_638 (O_638,N_9911,N_9944);
or UO_639 (O_639,N_9411,N_9201);
and UO_640 (O_640,N_9920,N_9187);
nand UO_641 (O_641,N_9521,N_9854);
and UO_642 (O_642,N_9692,N_9055);
and UO_643 (O_643,N_9109,N_9792);
or UO_644 (O_644,N_9597,N_9030);
nor UO_645 (O_645,N_9253,N_9758);
nor UO_646 (O_646,N_9924,N_9401);
nor UO_647 (O_647,N_9096,N_9819);
xnor UO_648 (O_648,N_9804,N_9490);
or UO_649 (O_649,N_9431,N_9383);
nor UO_650 (O_650,N_9887,N_9697);
nand UO_651 (O_651,N_9853,N_9157);
nand UO_652 (O_652,N_9253,N_9965);
nor UO_653 (O_653,N_9919,N_9357);
or UO_654 (O_654,N_9889,N_9224);
nor UO_655 (O_655,N_9088,N_9160);
and UO_656 (O_656,N_9845,N_9595);
and UO_657 (O_657,N_9313,N_9986);
nand UO_658 (O_658,N_9704,N_9779);
nor UO_659 (O_659,N_9367,N_9802);
nor UO_660 (O_660,N_9309,N_9661);
nand UO_661 (O_661,N_9324,N_9975);
and UO_662 (O_662,N_9361,N_9674);
nor UO_663 (O_663,N_9608,N_9401);
xor UO_664 (O_664,N_9797,N_9346);
or UO_665 (O_665,N_9266,N_9443);
xor UO_666 (O_666,N_9180,N_9864);
and UO_667 (O_667,N_9536,N_9159);
xor UO_668 (O_668,N_9153,N_9067);
nor UO_669 (O_669,N_9191,N_9531);
or UO_670 (O_670,N_9810,N_9399);
nand UO_671 (O_671,N_9069,N_9276);
nor UO_672 (O_672,N_9093,N_9958);
nand UO_673 (O_673,N_9296,N_9096);
xor UO_674 (O_674,N_9396,N_9964);
nor UO_675 (O_675,N_9804,N_9370);
and UO_676 (O_676,N_9716,N_9423);
and UO_677 (O_677,N_9266,N_9196);
nor UO_678 (O_678,N_9835,N_9368);
or UO_679 (O_679,N_9514,N_9775);
nand UO_680 (O_680,N_9447,N_9563);
nand UO_681 (O_681,N_9584,N_9730);
and UO_682 (O_682,N_9694,N_9256);
or UO_683 (O_683,N_9004,N_9699);
and UO_684 (O_684,N_9744,N_9945);
and UO_685 (O_685,N_9710,N_9925);
and UO_686 (O_686,N_9060,N_9907);
nor UO_687 (O_687,N_9426,N_9621);
and UO_688 (O_688,N_9229,N_9700);
or UO_689 (O_689,N_9755,N_9617);
nand UO_690 (O_690,N_9472,N_9178);
nor UO_691 (O_691,N_9436,N_9827);
or UO_692 (O_692,N_9651,N_9329);
xnor UO_693 (O_693,N_9587,N_9884);
nor UO_694 (O_694,N_9211,N_9188);
nor UO_695 (O_695,N_9381,N_9973);
nor UO_696 (O_696,N_9920,N_9239);
and UO_697 (O_697,N_9443,N_9613);
nand UO_698 (O_698,N_9098,N_9404);
xor UO_699 (O_699,N_9592,N_9693);
and UO_700 (O_700,N_9573,N_9819);
nand UO_701 (O_701,N_9126,N_9883);
xor UO_702 (O_702,N_9277,N_9255);
and UO_703 (O_703,N_9678,N_9203);
and UO_704 (O_704,N_9424,N_9952);
nor UO_705 (O_705,N_9423,N_9338);
or UO_706 (O_706,N_9441,N_9575);
or UO_707 (O_707,N_9258,N_9018);
nand UO_708 (O_708,N_9939,N_9580);
or UO_709 (O_709,N_9529,N_9613);
nand UO_710 (O_710,N_9114,N_9294);
or UO_711 (O_711,N_9545,N_9619);
and UO_712 (O_712,N_9465,N_9688);
and UO_713 (O_713,N_9419,N_9248);
or UO_714 (O_714,N_9168,N_9596);
xor UO_715 (O_715,N_9757,N_9488);
nor UO_716 (O_716,N_9059,N_9054);
and UO_717 (O_717,N_9015,N_9870);
and UO_718 (O_718,N_9970,N_9640);
and UO_719 (O_719,N_9667,N_9718);
nand UO_720 (O_720,N_9360,N_9317);
and UO_721 (O_721,N_9208,N_9214);
nor UO_722 (O_722,N_9642,N_9650);
nand UO_723 (O_723,N_9911,N_9506);
nand UO_724 (O_724,N_9858,N_9951);
nand UO_725 (O_725,N_9499,N_9372);
or UO_726 (O_726,N_9980,N_9016);
and UO_727 (O_727,N_9922,N_9698);
or UO_728 (O_728,N_9968,N_9069);
or UO_729 (O_729,N_9192,N_9985);
nor UO_730 (O_730,N_9241,N_9318);
and UO_731 (O_731,N_9278,N_9344);
and UO_732 (O_732,N_9785,N_9770);
nand UO_733 (O_733,N_9943,N_9188);
and UO_734 (O_734,N_9731,N_9634);
nor UO_735 (O_735,N_9409,N_9997);
xor UO_736 (O_736,N_9241,N_9254);
and UO_737 (O_737,N_9643,N_9829);
nand UO_738 (O_738,N_9947,N_9750);
nand UO_739 (O_739,N_9883,N_9213);
xor UO_740 (O_740,N_9226,N_9946);
or UO_741 (O_741,N_9037,N_9196);
nor UO_742 (O_742,N_9952,N_9524);
and UO_743 (O_743,N_9666,N_9464);
nor UO_744 (O_744,N_9488,N_9708);
nor UO_745 (O_745,N_9703,N_9969);
or UO_746 (O_746,N_9020,N_9419);
or UO_747 (O_747,N_9728,N_9613);
nor UO_748 (O_748,N_9729,N_9405);
and UO_749 (O_749,N_9538,N_9588);
or UO_750 (O_750,N_9978,N_9761);
nand UO_751 (O_751,N_9516,N_9304);
nor UO_752 (O_752,N_9308,N_9463);
nor UO_753 (O_753,N_9690,N_9019);
nand UO_754 (O_754,N_9100,N_9030);
nand UO_755 (O_755,N_9650,N_9151);
nor UO_756 (O_756,N_9922,N_9192);
nor UO_757 (O_757,N_9605,N_9579);
xnor UO_758 (O_758,N_9909,N_9796);
or UO_759 (O_759,N_9910,N_9135);
nand UO_760 (O_760,N_9625,N_9843);
nor UO_761 (O_761,N_9334,N_9791);
or UO_762 (O_762,N_9840,N_9874);
and UO_763 (O_763,N_9400,N_9341);
nand UO_764 (O_764,N_9381,N_9023);
nand UO_765 (O_765,N_9949,N_9233);
nand UO_766 (O_766,N_9567,N_9039);
and UO_767 (O_767,N_9528,N_9215);
and UO_768 (O_768,N_9513,N_9289);
nand UO_769 (O_769,N_9684,N_9423);
nand UO_770 (O_770,N_9719,N_9372);
xnor UO_771 (O_771,N_9409,N_9728);
or UO_772 (O_772,N_9311,N_9862);
nand UO_773 (O_773,N_9173,N_9601);
or UO_774 (O_774,N_9032,N_9086);
or UO_775 (O_775,N_9795,N_9938);
or UO_776 (O_776,N_9342,N_9133);
nand UO_777 (O_777,N_9437,N_9565);
nand UO_778 (O_778,N_9220,N_9842);
nor UO_779 (O_779,N_9968,N_9136);
and UO_780 (O_780,N_9014,N_9474);
nand UO_781 (O_781,N_9486,N_9447);
nand UO_782 (O_782,N_9095,N_9331);
nor UO_783 (O_783,N_9456,N_9657);
xnor UO_784 (O_784,N_9645,N_9178);
and UO_785 (O_785,N_9456,N_9906);
nand UO_786 (O_786,N_9649,N_9209);
nor UO_787 (O_787,N_9024,N_9310);
or UO_788 (O_788,N_9053,N_9322);
or UO_789 (O_789,N_9581,N_9996);
nor UO_790 (O_790,N_9036,N_9903);
nor UO_791 (O_791,N_9169,N_9445);
nand UO_792 (O_792,N_9023,N_9679);
and UO_793 (O_793,N_9506,N_9905);
nand UO_794 (O_794,N_9617,N_9784);
or UO_795 (O_795,N_9060,N_9513);
nor UO_796 (O_796,N_9760,N_9682);
nand UO_797 (O_797,N_9600,N_9464);
or UO_798 (O_798,N_9889,N_9280);
and UO_799 (O_799,N_9368,N_9848);
or UO_800 (O_800,N_9806,N_9568);
or UO_801 (O_801,N_9070,N_9361);
nor UO_802 (O_802,N_9336,N_9617);
and UO_803 (O_803,N_9291,N_9806);
nor UO_804 (O_804,N_9986,N_9530);
or UO_805 (O_805,N_9251,N_9884);
and UO_806 (O_806,N_9066,N_9096);
nand UO_807 (O_807,N_9208,N_9988);
nor UO_808 (O_808,N_9740,N_9866);
and UO_809 (O_809,N_9211,N_9370);
xnor UO_810 (O_810,N_9855,N_9085);
nor UO_811 (O_811,N_9694,N_9397);
and UO_812 (O_812,N_9212,N_9862);
and UO_813 (O_813,N_9355,N_9319);
and UO_814 (O_814,N_9383,N_9975);
xnor UO_815 (O_815,N_9810,N_9497);
nor UO_816 (O_816,N_9065,N_9762);
nand UO_817 (O_817,N_9586,N_9406);
or UO_818 (O_818,N_9197,N_9753);
nor UO_819 (O_819,N_9046,N_9570);
nor UO_820 (O_820,N_9201,N_9554);
or UO_821 (O_821,N_9071,N_9021);
and UO_822 (O_822,N_9450,N_9434);
nor UO_823 (O_823,N_9558,N_9452);
or UO_824 (O_824,N_9803,N_9160);
xnor UO_825 (O_825,N_9650,N_9495);
nand UO_826 (O_826,N_9938,N_9804);
xnor UO_827 (O_827,N_9073,N_9856);
and UO_828 (O_828,N_9335,N_9956);
or UO_829 (O_829,N_9935,N_9421);
nor UO_830 (O_830,N_9695,N_9075);
or UO_831 (O_831,N_9705,N_9076);
nor UO_832 (O_832,N_9332,N_9693);
nor UO_833 (O_833,N_9435,N_9561);
nand UO_834 (O_834,N_9632,N_9962);
and UO_835 (O_835,N_9788,N_9204);
xor UO_836 (O_836,N_9136,N_9288);
and UO_837 (O_837,N_9251,N_9576);
and UO_838 (O_838,N_9578,N_9739);
or UO_839 (O_839,N_9629,N_9937);
nand UO_840 (O_840,N_9087,N_9928);
and UO_841 (O_841,N_9097,N_9416);
nor UO_842 (O_842,N_9862,N_9594);
or UO_843 (O_843,N_9512,N_9090);
and UO_844 (O_844,N_9762,N_9376);
and UO_845 (O_845,N_9960,N_9009);
nand UO_846 (O_846,N_9468,N_9041);
or UO_847 (O_847,N_9095,N_9098);
nand UO_848 (O_848,N_9293,N_9594);
nor UO_849 (O_849,N_9032,N_9209);
and UO_850 (O_850,N_9097,N_9753);
nor UO_851 (O_851,N_9709,N_9601);
or UO_852 (O_852,N_9797,N_9592);
and UO_853 (O_853,N_9259,N_9189);
and UO_854 (O_854,N_9590,N_9972);
nor UO_855 (O_855,N_9189,N_9355);
nand UO_856 (O_856,N_9132,N_9299);
nand UO_857 (O_857,N_9490,N_9387);
and UO_858 (O_858,N_9645,N_9637);
or UO_859 (O_859,N_9225,N_9886);
nand UO_860 (O_860,N_9046,N_9098);
or UO_861 (O_861,N_9690,N_9629);
and UO_862 (O_862,N_9777,N_9576);
or UO_863 (O_863,N_9297,N_9981);
xnor UO_864 (O_864,N_9283,N_9339);
nor UO_865 (O_865,N_9559,N_9512);
nand UO_866 (O_866,N_9255,N_9688);
nand UO_867 (O_867,N_9286,N_9010);
or UO_868 (O_868,N_9624,N_9294);
nand UO_869 (O_869,N_9028,N_9340);
and UO_870 (O_870,N_9581,N_9101);
and UO_871 (O_871,N_9129,N_9011);
nor UO_872 (O_872,N_9710,N_9329);
nand UO_873 (O_873,N_9279,N_9128);
and UO_874 (O_874,N_9091,N_9973);
and UO_875 (O_875,N_9305,N_9764);
nor UO_876 (O_876,N_9402,N_9222);
nor UO_877 (O_877,N_9823,N_9644);
or UO_878 (O_878,N_9544,N_9900);
or UO_879 (O_879,N_9826,N_9705);
xnor UO_880 (O_880,N_9736,N_9225);
nor UO_881 (O_881,N_9618,N_9386);
nor UO_882 (O_882,N_9918,N_9002);
or UO_883 (O_883,N_9080,N_9308);
and UO_884 (O_884,N_9505,N_9299);
or UO_885 (O_885,N_9611,N_9258);
or UO_886 (O_886,N_9532,N_9132);
nand UO_887 (O_887,N_9738,N_9571);
nand UO_888 (O_888,N_9012,N_9176);
nor UO_889 (O_889,N_9766,N_9790);
and UO_890 (O_890,N_9344,N_9440);
and UO_891 (O_891,N_9539,N_9933);
nand UO_892 (O_892,N_9527,N_9659);
nor UO_893 (O_893,N_9239,N_9928);
or UO_894 (O_894,N_9534,N_9799);
nor UO_895 (O_895,N_9602,N_9411);
and UO_896 (O_896,N_9508,N_9231);
nand UO_897 (O_897,N_9904,N_9682);
and UO_898 (O_898,N_9315,N_9594);
nand UO_899 (O_899,N_9065,N_9388);
nand UO_900 (O_900,N_9304,N_9483);
xor UO_901 (O_901,N_9310,N_9214);
xnor UO_902 (O_902,N_9554,N_9080);
and UO_903 (O_903,N_9081,N_9705);
and UO_904 (O_904,N_9016,N_9210);
nor UO_905 (O_905,N_9045,N_9538);
or UO_906 (O_906,N_9289,N_9044);
nand UO_907 (O_907,N_9868,N_9494);
or UO_908 (O_908,N_9081,N_9943);
nor UO_909 (O_909,N_9900,N_9648);
or UO_910 (O_910,N_9568,N_9016);
xor UO_911 (O_911,N_9727,N_9774);
or UO_912 (O_912,N_9248,N_9358);
and UO_913 (O_913,N_9209,N_9675);
nor UO_914 (O_914,N_9710,N_9878);
or UO_915 (O_915,N_9002,N_9988);
nand UO_916 (O_916,N_9805,N_9916);
nor UO_917 (O_917,N_9640,N_9902);
xnor UO_918 (O_918,N_9809,N_9743);
or UO_919 (O_919,N_9537,N_9260);
nand UO_920 (O_920,N_9319,N_9490);
or UO_921 (O_921,N_9375,N_9195);
nor UO_922 (O_922,N_9149,N_9997);
or UO_923 (O_923,N_9631,N_9071);
nor UO_924 (O_924,N_9910,N_9605);
and UO_925 (O_925,N_9936,N_9425);
and UO_926 (O_926,N_9870,N_9513);
nand UO_927 (O_927,N_9027,N_9702);
nor UO_928 (O_928,N_9327,N_9788);
and UO_929 (O_929,N_9887,N_9082);
or UO_930 (O_930,N_9939,N_9126);
or UO_931 (O_931,N_9913,N_9689);
and UO_932 (O_932,N_9588,N_9008);
nand UO_933 (O_933,N_9629,N_9953);
nand UO_934 (O_934,N_9449,N_9621);
nor UO_935 (O_935,N_9123,N_9657);
and UO_936 (O_936,N_9981,N_9495);
and UO_937 (O_937,N_9026,N_9528);
xnor UO_938 (O_938,N_9757,N_9814);
nand UO_939 (O_939,N_9384,N_9629);
nand UO_940 (O_940,N_9736,N_9830);
or UO_941 (O_941,N_9799,N_9362);
nand UO_942 (O_942,N_9415,N_9485);
nand UO_943 (O_943,N_9062,N_9361);
nand UO_944 (O_944,N_9948,N_9263);
or UO_945 (O_945,N_9975,N_9685);
nand UO_946 (O_946,N_9440,N_9178);
nand UO_947 (O_947,N_9571,N_9370);
or UO_948 (O_948,N_9895,N_9209);
nor UO_949 (O_949,N_9447,N_9582);
or UO_950 (O_950,N_9266,N_9211);
nor UO_951 (O_951,N_9881,N_9097);
and UO_952 (O_952,N_9517,N_9271);
nor UO_953 (O_953,N_9897,N_9537);
and UO_954 (O_954,N_9588,N_9233);
nand UO_955 (O_955,N_9804,N_9718);
xnor UO_956 (O_956,N_9808,N_9930);
or UO_957 (O_957,N_9769,N_9667);
and UO_958 (O_958,N_9686,N_9003);
or UO_959 (O_959,N_9551,N_9512);
and UO_960 (O_960,N_9917,N_9222);
nor UO_961 (O_961,N_9985,N_9064);
nand UO_962 (O_962,N_9295,N_9460);
nor UO_963 (O_963,N_9470,N_9780);
nand UO_964 (O_964,N_9928,N_9857);
and UO_965 (O_965,N_9576,N_9748);
nor UO_966 (O_966,N_9563,N_9371);
and UO_967 (O_967,N_9120,N_9101);
xnor UO_968 (O_968,N_9761,N_9487);
nand UO_969 (O_969,N_9523,N_9913);
or UO_970 (O_970,N_9160,N_9007);
and UO_971 (O_971,N_9412,N_9726);
and UO_972 (O_972,N_9894,N_9957);
and UO_973 (O_973,N_9808,N_9780);
or UO_974 (O_974,N_9375,N_9664);
and UO_975 (O_975,N_9760,N_9282);
nor UO_976 (O_976,N_9536,N_9047);
nand UO_977 (O_977,N_9814,N_9739);
nand UO_978 (O_978,N_9454,N_9421);
and UO_979 (O_979,N_9420,N_9041);
and UO_980 (O_980,N_9815,N_9893);
nand UO_981 (O_981,N_9039,N_9001);
or UO_982 (O_982,N_9559,N_9003);
nand UO_983 (O_983,N_9172,N_9257);
and UO_984 (O_984,N_9694,N_9747);
and UO_985 (O_985,N_9621,N_9010);
nand UO_986 (O_986,N_9913,N_9084);
xnor UO_987 (O_987,N_9339,N_9116);
nor UO_988 (O_988,N_9775,N_9842);
nand UO_989 (O_989,N_9842,N_9881);
and UO_990 (O_990,N_9599,N_9462);
nand UO_991 (O_991,N_9796,N_9034);
xor UO_992 (O_992,N_9442,N_9458);
nor UO_993 (O_993,N_9159,N_9116);
or UO_994 (O_994,N_9809,N_9658);
nand UO_995 (O_995,N_9887,N_9052);
or UO_996 (O_996,N_9523,N_9613);
nor UO_997 (O_997,N_9658,N_9320);
nor UO_998 (O_998,N_9608,N_9800);
nor UO_999 (O_999,N_9119,N_9771);
or UO_1000 (O_1000,N_9053,N_9030);
nor UO_1001 (O_1001,N_9469,N_9443);
xor UO_1002 (O_1002,N_9535,N_9936);
or UO_1003 (O_1003,N_9572,N_9218);
nand UO_1004 (O_1004,N_9343,N_9880);
or UO_1005 (O_1005,N_9167,N_9021);
nand UO_1006 (O_1006,N_9266,N_9437);
nand UO_1007 (O_1007,N_9614,N_9005);
xor UO_1008 (O_1008,N_9562,N_9427);
nor UO_1009 (O_1009,N_9568,N_9263);
nor UO_1010 (O_1010,N_9967,N_9805);
or UO_1011 (O_1011,N_9817,N_9326);
xor UO_1012 (O_1012,N_9527,N_9723);
nand UO_1013 (O_1013,N_9216,N_9305);
xor UO_1014 (O_1014,N_9462,N_9702);
or UO_1015 (O_1015,N_9153,N_9014);
or UO_1016 (O_1016,N_9683,N_9093);
nor UO_1017 (O_1017,N_9220,N_9294);
nor UO_1018 (O_1018,N_9527,N_9238);
or UO_1019 (O_1019,N_9820,N_9832);
xor UO_1020 (O_1020,N_9835,N_9643);
and UO_1021 (O_1021,N_9706,N_9892);
or UO_1022 (O_1022,N_9532,N_9156);
xnor UO_1023 (O_1023,N_9217,N_9537);
xor UO_1024 (O_1024,N_9487,N_9273);
nand UO_1025 (O_1025,N_9118,N_9071);
or UO_1026 (O_1026,N_9140,N_9793);
nand UO_1027 (O_1027,N_9467,N_9786);
or UO_1028 (O_1028,N_9257,N_9297);
nand UO_1029 (O_1029,N_9164,N_9734);
nor UO_1030 (O_1030,N_9909,N_9289);
nand UO_1031 (O_1031,N_9907,N_9051);
nand UO_1032 (O_1032,N_9118,N_9253);
nand UO_1033 (O_1033,N_9792,N_9048);
or UO_1034 (O_1034,N_9818,N_9893);
nand UO_1035 (O_1035,N_9143,N_9601);
and UO_1036 (O_1036,N_9325,N_9768);
or UO_1037 (O_1037,N_9913,N_9178);
nor UO_1038 (O_1038,N_9058,N_9918);
or UO_1039 (O_1039,N_9068,N_9983);
nor UO_1040 (O_1040,N_9590,N_9821);
nor UO_1041 (O_1041,N_9008,N_9182);
or UO_1042 (O_1042,N_9818,N_9735);
and UO_1043 (O_1043,N_9201,N_9933);
and UO_1044 (O_1044,N_9588,N_9671);
nand UO_1045 (O_1045,N_9413,N_9653);
nand UO_1046 (O_1046,N_9306,N_9724);
nand UO_1047 (O_1047,N_9804,N_9047);
nand UO_1048 (O_1048,N_9507,N_9351);
and UO_1049 (O_1049,N_9813,N_9971);
xnor UO_1050 (O_1050,N_9241,N_9656);
nor UO_1051 (O_1051,N_9109,N_9899);
xor UO_1052 (O_1052,N_9959,N_9101);
xor UO_1053 (O_1053,N_9072,N_9779);
or UO_1054 (O_1054,N_9127,N_9209);
and UO_1055 (O_1055,N_9016,N_9134);
and UO_1056 (O_1056,N_9220,N_9877);
and UO_1057 (O_1057,N_9294,N_9256);
nand UO_1058 (O_1058,N_9225,N_9376);
nand UO_1059 (O_1059,N_9977,N_9321);
or UO_1060 (O_1060,N_9061,N_9655);
and UO_1061 (O_1061,N_9567,N_9594);
xnor UO_1062 (O_1062,N_9838,N_9424);
xnor UO_1063 (O_1063,N_9489,N_9783);
xor UO_1064 (O_1064,N_9158,N_9412);
nand UO_1065 (O_1065,N_9738,N_9096);
nand UO_1066 (O_1066,N_9194,N_9031);
and UO_1067 (O_1067,N_9346,N_9748);
or UO_1068 (O_1068,N_9837,N_9590);
or UO_1069 (O_1069,N_9584,N_9305);
and UO_1070 (O_1070,N_9109,N_9547);
nand UO_1071 (O_1071,N_9913,N_9184);
nand UO_1072 (O_1072,N_9081,N_9919);
or UO_1073 (O_1073,N_9424,N_9595);
or UO_1074 (O_1074,N_9259,N_9523);
nor UO_1075 (O_1075,N_9722,N_9340);
nand UO_1076 (O_1076,N_9952,N_9438);
nand UO_1077 (O_1077,N_9993,N_9100);
xor UO_1078 (O_1078,N_9401,N_9989);
nor UO_1079 (O_1079,N_9563,N_9550);
nand UO_1080 (O_1080,N_9351,N_9677);
and UO_1081 (O_1081,N_9168,N_9165);
nand UO_1082 (O_1082,N_9357,N_9425);
or UO_1083 (O_1083,N_9638,N_9229);
or UO_1084 (O_1084,N_9273,N_9815);
and UO_1085 (O_1085,N_9702,N_9052);
and UO_1086 (O_1086,N_9882,N_9115);
nand UO_1087 (O_1087,N_9516,N_9318);
nor UO_1088 (O_1088,N_9450,N_9437);
nand UO_1089 (O_1089,N_9069,N_9733);
nand UO_1090 (O_1090,N_9299,N_9837);
nor UO_1091 (O_1091,N_9466,N_9156);
or UO_1092 (O_1092,N_9961,N_9644);
nor UO_1093 (O_1093,N_9136,N_9782);
xor UO_1094 (O_1094,N_9955,N_9473);
xor UO_1095 (O_1095,N_9350,N_9453);
nand UO_1096 (O_1096,N_9922,N_9594);
nand UO_1097 (O_1097,N_9440,N_9811);
xnor UO_1098 (O_1098,N_9764,N_9138);
nor UO_1099 (O_1099,N_9758,N_9498);
or UO_1100 (O_1100,N_9316,N_9896);
nand UO_1101 (O_1101,N_9395,N_9688);
nor UO_1102 (O_1102,N_9745,N_9446);
nand UO_1103 (O_1103,N_9705,N_9721);
nand UO_1104 (O_1104,N_9554,N_9617);
nand UO_1105 (O_1105,N_9779,N_9321);
or UO_1106 (O_1106,N_9849,N_9310);
or UO_1107 (O_1107,N_9441,N_9006);
and UO_1108 (O_1108,N_9996,N_9765);
or UO_1109 (O_1109,N_9444,N_9435);
or UO_1110 (O_1110,N_9326,N_9978);
nor UO_1111 (O_1111,N_9136,N_9978);
and UO_1112 (O_1112,N_9213,N_9111);
nand UO_1113 (O_1113,N_9437,N_9912);
or UO_1114 (O_1114,N_9634,N_9291);
nand UO_1115 (O_1115,N_9383,N_9328);
or UO_1116 (O_1116,N_9713,N_9653);
and UO_1117 (O_1117,N_9454,N_9791);
and UO_1118 (O_1118,N_9112,N_9188);
or UO_1119 (O_1119,N_9930,N_9508);
or UO_1120 (O_1120,N_9399,N_9043);
nor UO_1121 (O_1121,N_9823,N_9756);
or UO_1122 (O_1122,N_9965,N_9273);
nor UO_1123 (O_1123,N_9557,N_9908);
nand UO_1124 (O_1124,N_9325,N_9713);
xnor UO_1125 (O_1125,N_9766,N_9397);
nand UO_1126 (O_1126,N_9687,N_9713);
nand UO_1127 (O_1127,N_9425,N_9902);
nor UO_1128 (O_1128,N_9182,N_9648);
and UO_1129 (O_1129,N_9192,N_9988);
or UO_1130 (O_1130,N_9022,N_9045);
nand UO_1131 (O_1131,N_9286,N_9200);
nand UO_1132 (O_1132,N_9450,N_9248);
nand UO_1133 (O_1133,N_9486,N_9082);
or UO_1134 (O_1134,N_9605,N_9661);
and UO_1135 (O_1135,N_9763,N_9779);
and UO_1136 (O_1136,N_9337,N_9389);
xnor UO_1137 (O_1137,N_9524,N_9476);
nor UO_1138 (O_1138,N_9867,N_9393);
or UO_1139 (O_1139,N_9801,N_9428);
nor UO_1140 (O_1140,N_9901,N_9606);
xor UO_1141 (O_1141,N_9808,N_9016);
nor UO_1142 (O_1142,N_9940,N_9591);
nand UO_1143 (O_1143,N_9165,N_9430);
nor UO_1144 (O_1144,N_9958,N_9629);
or UO_1145 (O_1145,N_9066,N_9679);
nor UO_1146 (O_1146,N_9889,N_9287);
nand UO_1147 (O_1147,N_9690,N_9163);
nand UO_1148 (O_1148,N_9483,N_9992);
nand UO_1149 (O_1149,N_9352,N_9117);
and UO_1150 (O_1150,N_9530,N_9980);
nand UO_1151 (O_1151,N_9445,N_9679);
or UO_1152 (O_1152,N_9388,N_9596);
nand UO_1153 (O_1153,N_9601,N_9988);
and UO_1154 (O_1154,N_9269,N_9220);
nand UO_1155 (O_1155,N_9594,N_9241);
nor UO_1156 (O_1156,N_9792,N_9706);
nand UO_1157 (O_1157,N_9856,N_9685);
nand UO_1158 (O_1158,N_9405,N_9437);
and UO_1159 (O_1159,N_9208,N_9027);
nand UO_1160 (O_1160,N_9245,N_9812);
nor UO_1161 (O_1161,N_9738,N_9432);
nand UO_1162 (O_1162,N_9381,N_9816);
nor UO_1163 (O_1163,N_9892,N_9264);
nand UO_1164 (O_1164,N_9819,N_9493);
nand UO_1165 (O_1165,N_9102,N_9448);
nand UO_1166 (O_1166,N_9720,N_9254);
or UO_1167 (O_1167,N_9649,N_9430);
and UO_1168 (O_1168,N_9935,N_9413);
or UO_1169 (O_1169,N_9212,N_9077);
or UO_1170 (O_1170,N_9681,N_9729);
nor UO_1171 (O_1171,N_9723,N_9207);
nor UO_1172 (O_1172,N_9207,N_9773);
nor UO_1173 (O_1173,N_9001,N_9828);
or UO_1174 (O_1174,N_9013,N_9808);
nand UO_1175 (O_1175,N_9440,N_9603);
nor UO_1176 (O_1176,N_9031,N_9239);
or UO_1177 (O_1177,N_9098,N_9861);
nor UO_1178 (O_1178,N_9603,N_9608);
or UO_1179 (O_1179,N_9295,N_9173);
or UO_1180 (O_1180,N_9812,N_9174);
nor UO_1181 (O_1181,N_9977,N_9114);
or UO_1182 (O_1182,N_9714,N_9930);
nand UO_1183 (O_1183,N_9107,N_9422);
and UO_1184 (O_1184,N_9281,N_9271);
or UO_1185 (O_1185,N_9905,N_9874);
nor UO_1186 (O_1186,N_9751,N_9729);
and UO_1187 (O_1187,N_9081,N_9031);
and UO_1188 (O_1188,N_9952,N_9397);
nand UO_1189 (O_1189,N_9056,N_9466);
and UO_1190 (O_1190,N_9836,N_9348);
nand UO_1191 (O_1191,N_9558,N_9929);
nand UO_1192 (O_1192,N_9149,N_9629);
or UO_1193 (O_1193,N_9936,N_9116);
or UO_1194 (O_1194,N_9365,N_9017);
nand UO_1195 (O_1195,N_9513,N_9254);
nor UO_1196 (O_1196,N_9862,N_9707);
and UO_1197 (O_1197,N_9908,N_9609);
and UO_1198 (O_1198,N_9487,N_9291);
nand UO_1199 (O_1199,N_9454,N_9523);
and UO_1200 (O_1200,N_9818,N_9002);
nor UO_1201 (O_1201,N_9168,N_9985);
and UO_1202 (O_1202,N_9539,N_9379);
nor UO_1203 (O_1203,N_9121,N_9337);
xnor UO_1204 (O_1204,N_9073,N_9345);
nor UO_1205 (O_1205,N_9395,N_9422);
and UO_1206 (O_1206,N_9057,N_9411);
nand UO_1207 (O_1207,N_9531,N_9671);
nand UO_1208 (O_1208,N_9746,N_9382);
nor UO_1209 (O_1209,N_9398,N_9845);
nand UO_1210 (O_1210,N_9179,N_9594);
and UO_1211 (O_1211,N_9583,N_9802);
and UO_1212 (O_1212,N_9772,N_9130);
or UO_1213 (O_1213,N_9959,N_9801);
and UO_1214 (O_1214,N_9505,N_9911);
nand UO_1215 (O_1215,N_9609,N_9553);
or UO_1216 (O_1216,N_9635,N_9525);
xor UO_1217 (O_1217,N_9819,N_9102);
or UO_1218 (O_1218,N_9189,N_9184);
nor UO_1219 (O_1219,N_9318,N_9493);
or UO_1220 (O_1220,N_9597,N_9378);
and UO_1221 (O_1221,N_9457,N_9742);
nor UO_1222 (O_1222,N_9678,N_9017);
nand UO_1223 (O_1223,N_9685,N_9287);
nand UO_1224 (O_1224,N_9858,N_9350);
xor UO_1225 (O_1225,N_9035,N_9856);
and UO_1226 (O_1226,N_9620,N_9456);
nand UO_1227 (O_1227,N_9636,N_9389);
and UO_1228 (O_1228,N_9419,N_9398);
or UO_1229 (O_1229,N_9351,N_9148);
nand UO_1230 (O_1230,N_9649,N_9152);
nor UO_1231 (O_1231,N_9708,N_9723);
xor UO_1232 (O_1232,N_9920,N_9736);
nor UO_1233 (O_1233,N_9499,N_9491);
nor UO_1234 (O_1234,N_9616,N_9072);
nor UO_1235 (O_1235,N_9061,N_9617);
and UO_1236 (O_1236,N_9794,N_9194);
and UO_1237 (O_1237,N_9118,N_9265);
or UO_1238 (O_1238,N_9558,N_9742);
or UO_1239 (O_1239,N_9061,N_9159);
nand UO_1240 (O_1240,N_9091,N_9271);
nor UO_1241 (O_1241,N_9683,N_9267);
or UO_1242 (O_1242,N_9506,N_9934);
nor UO_1243 (O_1243,N_9178,N_9298);
xor UO_1244 (O_1244,N_9248,N_9965);
and UO_1245 (O_1245,N_9048,N_9907);
or UO_1246 (O_1246,N_9546,N_9244);
or UO_1247 (O_1247,N_9082,N_9440);
or UO_1248 (O_1248,N_9500,N_9921);
or UO_1249 (O_1249,N_9950,N_9897);
and UO_1250 (O_1250,N_9018,N_9701);
nor UO_1251 (O_1251,N_9185,N_9706);
nand UO_1252 (O_1252,N_9528,N_9676);
and UO_1253 (O_1253,N_9632,N_9916);
xor UO_1254 (O_1254,N_9000,N_9582);
nor UO_1255 (O_1255,N_9200,N_9346);
nor UO_1256 (O_1256,N_9965,N_9801);
and UO_1257 (O_1257,N_9774,N_9905);
nand UO_1258 (O_1258,N_9955,N_9480);
nand UO_1259 (O_1259,N_9513,N_9169);
or UO_1260 (O_1260,N_9745,N_9238);
nor UO_1261 (O_1261,N_9795,N_9498);
or UO_1262 (O_1262,N_9169,N_9175);
nand UO_1263 (O_1263,N_9679,N_9712);
or UO_1264 (O_1264,N_9526,N_9772);
and UO_1265 (O_1265,N_9572,N_9380);
nand UO_1266 (O_1266,N_9253,N_9220);
xor UO_1267 (O_1267,N_9727,N_9341);
or UO_1268 (O_1268,N_9322,N_9892);
or UO_1269 (O_1269,N_9844,N_9111);
nor UO_1270 (O_1270,N_9617,N_9645);
nand UO_1271 (O_1271,N_9799,N_9310);
nor UO_1272 (O_1272,N_9964,N_9486);
and UO_1273 (O_1273,N_9399,N_9559);
nand UO_1274 (O_1274,N_9231,N_9096);
nor UO_1275 (O_1275,N_9657,N_9581);
or UO_1276 (O_1276,N_9233,N_9354);
and UO_1277 (O_1277,N_9310,N_9136);
nand UO_1278 (O_1278,N_9654,N_9477);
nand UO_1279 (O_1279,N_9871,N_9103);
nand UO_1280 (O_1280,N_9881,N_9840);
xnor UO_1281 (O_1281,N_9168,N_9197);
and UO_1282 (O_1282,N_9673,N_9256);
or UO_1283 (O_1283,N_9898,N_9544);
and UO_1284 (O_1284,N_9325,N_9099);
nand UO_1285 (O_1285,N_9533,N_9738);
nand UO_1286 (O_1286,N_9612,N_9562);
or UO_1287 (O_1287,N_9339,N_9527);
nand UO_1288 (O_1288,N_9361,N_9795);
xnor UO_1289 (O_1289,N_9946,N_9392);
and UO_1290 (O_1290,N_9445,N_9565);
nand UO_1291 (O_1291,N_9834,N_9685);
and UO_1292 (O_1292,N_9670,N_9710);
nand UO_1293 (O_1293,N_9595,N_9629);
and UO_1294 (O_1294,N_9144,N_9736);
and UO_1295 (O_1295,N_9535,N_9779);
or UO_1296 (O_1296,N_9497,N_9286);
and UO_1297 (O_1297,N_9486,N_9606);
nand UO_1298 (O_1298,N_9710,N_9227);
xor UO_1299 (O_1299,N_9672,N_9405);
xnor UO_1300 (O_1300,N_9675,N_9255);
nand UO_1301 (O_1301,N_9505,N_9670);
xnor UO_1302 (O_1302,N_9601,N_9760);
or UO_1303 (O_1303,N_9548,N_9943);
nand UO_1304 (O_1304,N_9426,N_9180);
or UO_1305 (O_1305,N_9672,N_9760);
nand UO_1306 (O_1306,N_9257,N_9141);
nor UO_1307 (O_1307,N_9834,N_9360);
or UO_1308 (O_1308,N_9092,N_9102);
xor UO_1309 (O_1309,N_9813,N_9427);
nor UO_1310 (O_1310,N_9840,N_9657);
nor UO_1311 (O_1311,N_9893,N_9269);
or UO_1312 (O_1312,N_9695,N_9903);
nor UO_1313 (O_1313,N_9185,N_9191);
or UO_1314 (O_1314,N_9285,N_9138);
or UO_1315 (O_1315,N_9885,N_9203);
nor UO_1316 (O_1316,N_9525,N_9669);
and UO_1317 (O_1317,N_9763,N_9791);
and UO_1318 (O_1318,N_9790,N_9016);
nand UO_1319 (O_1319,N_9546,N_9904);
nor UO_1320 (O_1320,N_9300,N_9211);
or UO_1321 (O_1321,N_9421,N_9884);
or UO_1322 (O_1322,N_9083,N_9536);
nand UO_1323 (O_1323,N_9001,N_9104);
nand UO_1324 (O_1324,N_9478,N_9578);
xnor UO_1325 (O_1325,N_9988,N_9815);
or UO_1326 (O_1326,N_9098,N_9890);
or UO_1327 (O_1327,N_9397,N_9681);
nand UO_1328 (O_1328,N_9813,N_9542);
nand UO_1329 (O_1329,N_9408,N_9629);
or UO_1330 (O_1330,N_9696,N_9763);
nor UO_1331 (O_1331,N_9087,N_9789);
and UO_1332 (O_1332,N_9958,N_9254);
and UO_1333 (O_1333,N_9749,N_9936);
and UO_1334 (O_1334,N_9979,N_9576);
or UO_1335 (O_1335,N_9496,N_9516);
xor UO_1336 (O_1336,N_9794,N_9952);
xnor UO_1337 (O_1337,N_9527,N_9538);
nor UO_1338 (O_1338,N_9839,N_9688);
and UO_1339 (O_1339,N_9117,N_9852);
and UO_1340 (O_1340,N_9208,N_9138);
and UO_1341 (O_1341,N_9532,N_9735);
or UO_1342 (O_1342,N_9592,N_9388);
and UO_1343 (O_1343,N_9447,N_9949);
and UO_1344 (O_1344,N_9184,N_9882);
xor UO_1345 (O_1345,N_9713,N_9999);
or UO_1346 (O_1346,N_9623,N_9461);
xnor UO_1347 (O_1347,N_9763,N_9031);
or UO_1348 (O_1348,N_9568,N_9589);
xnor UO_1349 (O_1349,N_9499,N_9945);
xor UO_1350 (O_1350,N_9199,N_9934);
and UO_1351 (O_1351,N_9327,N_9453);
and UO_1352 (O_1352,N_9305,N_9253);
and UO_1353 (O_1353,N_9843,N_9774);
or UO_1354 (O_1354,N_9376,N_9968);
nand UO_1355 (O_1355,N_9393,N_9710);
nor UO_1356 (O_1356,N_9719,N_9390);
nor UO_1357 (O_1357,N_9593,N_9301);
nand UO_1358 (O_1358,N_9685,N_9899);
or UO_1359 (O_1359,N_9374,N_9317);
nor UO_1360 (O_1360,N_9969,N_9435);
nand UO_1361 (O_1361,N_9336,N_9129);
nor UO_1362 (O_1362,N_9766,N_9625);
nand UO_1363 (O_1363,N_9891,N_9376);
or UO_1364 (O_1364,N_9891,N_9613);
and UO_1365 (O_1365,N_9709,N_9767);
or UO_1366 (O_1366,N_9146,N_9478);
and UO_1367 (O_1367,N_9410,N_9866);
nor UO_1368 (O_1368,N_9950,N_9143);
and UO_1369 (O_1369,N_9027,N_9941);
and UO_1370 (O_1370,N_9243,N_9835);
and UO_1371 (O_1371,N_9302,N_9547);
or UO_1372 (O_1372,N_9115,N_9203);
and UO_1373 (O_1373,N_9182,N_9007);
or UO_1374 (O_1374,N_9929,N_9957);
nor UO_1375 (O_1375,N_9832,N_9434);
or UO_1376 (O_1376,N_9627,N_9052);
nand UO_1377 (O_1377,N_9839,N_9007);
or UO_1378 (O_1378,N_9891,N_9727);
and UO_1379 (O_1379,N_9553,N_9864);
and UO_1380 (O_1380,N_9841,N_9891);
nand UO_1381 (O_1381,N_9554,N_9077);
or UO_1382 (O_1382,N_9322,N_9389);
or UO_1383 (O_1383,N_9103,N_9366);
and UO_1384 (O_1384,N_9298,N_9247);
nand UO_1385 (O_1385,N_9162,N_9139);
nor UO_1386 (O_1386,N_9979,N_9470);
xor UO_1387 (O_1387,N_9523,N_9495);
nand UO_1388 (O_1388,N_9676,N_9960);
xor UO_1389 (O_1389,N_9243,N_9660);
nand UO_1390 (O_1390,N_9471,N_9147);
nor UO_1391 (O_1391,N_9589,N_9130);
nor UO_1392 (O_1392,N_9455,N_9639);
or UO_1393 (O_1393,N_9162,N_9013);
xor UO_1394 (O_1394,N_9753,N_9020);
nand UO_1395 (O_1395,N_9343,N_9278);
and UO_1396 (O_1396,N_9548,N_9018);
nor UO_1397 (O_1397,N_9136,N_9024);
and UO_1398 (O_1398,N_9528,N_9516);
nor UO_1399 (O_1399,N_9011,N_9671);
or UO_1400 (O_1400,N_9819,N_9756);
nor UO_1401 (O_1401,N_9905,N_9006);
or UO_1402 (O_1402,N_9312,N_9128);
nand UO_1403 (O_1403,N_9086,N_9503);
nor UO_1404 (O_1404,N_9847,N_9315);
or UO_1405 (O_1405,N_9721,N_9912);
nor UO_1406 (O_1406,N_9425,N_9749);
and UO_1407 (O_1407,N_9847,N_9353);
and UO_1408 (O_1408,N_9571,N_9518);
or UO_1409 (O_1409,N_9782,N_9468);
xor UO_1410 (O_1410,N_9510,N_9485);
or UO_1411 (O_1411,N_9315,N_9232);
nor UO_1412 (O_1412,N_9277,N_9138);
or UO_1413 (O_1413,N_9182,N_9814);
nand UO_1414 (O_1414,N_9368,N_9262);
xor UO_1415 (O_1415,N_9741,N_9607);
or UO_1416 (O_1416,N_9100,N_9511);
nand UO_1417 (O_1417,N_9096,N_9142);
nor UO_1418 (O_1418,N_9224,N_9291);
xnor UO_1419 (O_1419,N_9479,N_9225);
and UO_1420 (O_1420,N_9581,N_9187);
nand UO_1421 (O_1421,N_9002,N_9766);
nand UO_1422 (O_1422,N_9872,N_9999);
xnor UO_1423 (O_1423,N_9878,N_9451);
nand UO_1424 (O_1424,N_9558,N_9834);
nor UO_1425 (O_1425,N_9476,N_9762);
and UO_1426 (O_1426,N_9553,N_9904);
or UO_1427 (O_1427,N_9019,N_9317);
nand UO_1428 (O_1428,N_9542,N_9393);
and UO_1429 (O_1429,N_9097,N_9350);
nand UO_1430 (O_1430,N_9864,N_9875);
nor UO_1431 (O_1431,N_9384,N_9812);
and UO_1432 (O_1432,N_9293,N_9929);
and UO_1433 (O_1433,N_9787,N_9415);
or UO_1434 (O_1434,N_9899,N_9383);
nor UO_1435 (O_1435,N_9328,N_9199);
and UO_1436 (O_1436,N_9311,N_9657);
and UO_1437 (O_1437,N_9220,N_9709);
nor UO_1438 (O_1438,N_9906,N_9049);
or UO_1439 (O_1439,N_9257,N_9612);
or UO_1440 (O_1440,N_9912,N_9430);
nor UO_1441 (O_1441,N_9263,N_9526);
nor UO_1442 (O_1442,N_9464,N_9408);
or UO_1443 (O_1443,N_9541,N_9074);
and UO_1444 (O_1444,N_9692,N_9395);
nor UO_1445 (O_1445,N_9260,N_9671);
nand UO_1446 (O_1446,N_9515,N_9122);
nor UO_1447 (O_1447,N_9690,N_9384);
and UO_1448 (O_1448,N_9088,N_9233);
and UO_1449 (O_1449,N_9608,N_9684);
nor UO_1450 (O_1450,N_9217,N_9515);
xnor UO_1451 (O_1451,N_9618,N_9713);
nand UO_1452 (O_1452,N_9183,N_9519);
nand UO_1453 (O_1453,N_9845,N_9739);
or UO_1454 (O_1454,N_9468,N_9465);
or UO_1455 (O_1455,N_9806,N_9561);
nand UO_1456 (O_1456,N_9280,N_9207);
nor UO_1457 (O_1457,N_9167,N_9852);
nand UO_1458 (O_1458,N_9377,N_9889);
or UO_1459 (O_1459,N_9410,N_9529);
nor UO_1460 (O_1460,N_9207,N_9525);
or UO_1461 (O_1461,N_9554,N_9624);
nand UO_1462 (O_1462,N_9320,N_9183);
xnor UO_1463 (O_1463,N_9096,N_9487);
or UO_1464 (O_1464,N_9066,N_9753);
xor UO_1465 (O_1465,N_9199,N_9799);
or UO_1466 (O_1466,N_9144,N_9912);
nor UO_1467 (O_1467,N_9795,N_9633);
or UO_1468 (O_1468,N_9166,N_9486);
nand UO_1469 (O_1469,N_9711,N_9353);
nand UO_1470 (O_1470,N_9614,N_9344);
and UO_1471 (O_1471,N_9724,N_9825);
xor UO_1472 (O_1472,N_9288,N_9856);
nor UO_1473 (O_1473,N_9578,N_9547);
nor UO_1474 (O_1474,N_9520,N_9024);
and UO_1475 (O_1475,N_9864,N_9492);
xor UO_1476 (O_1476,N_9744,N_9889);
nor UO_1477 (O_1477,N_9410,N_9296);
xor UO_1478 (O_1478,N_9944,N_9983);
or UO_1479 (O_1479,N_9083,N_9567);
and UO_1480 (O_1480,N_9891,N_9333);
nand UO_1481 (O_1481,N_9921,N_9689);
or UO_1482 (O_1482,N_9949,N_9327);
nor UO_1483 (O_1483,N_9541,N_9722);
nor UO_1484 (O_1484,N_9524,N_9995);
and UO_1485 (O_1485,N_9069,N_9593);
nand UO_1486 (O_1486,N_9303,N_9798);
nor UO_1487 (O_1487,N_9989,N_9808);
and UO_1488 (O_1488,N_9668,N_9785);
or UO_1489 (O_1489,N_9761,N_9473);
nor UO_1490 (O_1490,N_9254,N_9835);
and UO_1491 (O_1491,N_9805,N_9161);
nor UO_1492 (O_1492,N_9612,N_9319);
and UO_1493 (O_1493,N_9503,N_9529);
nor UO_1494 (O_1494,N_9430,N_9761);
nand UO_1495 (O_1495,N_9576,N_9670);
and UO_1496 (O_1496,N_9074,N_9955);
and UO_1497 (O_1497,N_9460,N_9870);
or UO_1498 (O_1498,N_9540,N_9930);
xnor UO_1499 (O_1499,N_9236,N_9281);
endmodule