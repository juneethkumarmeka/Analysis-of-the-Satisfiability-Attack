module basic_500_3000_500_6_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_367,In_103);
and U1 (N_1,In_441,In_25);
nor U2 (N_2,In_323,In_224);
and U3 (N_3,In_374,In_259);
nand U4 (N_4,In_225,In_78);
and U5 (N_5,In_221,In_453);
nor U6 (N_6,In_84,In_198);
and U7 (N_7,In_286,In_394);
or U8 (N_8,In_306,In_55);
or U9 (N_9,In_112,In_419);
or U10 (N_10,In_216,In_324);
nor U11 (N_11,In_489,In_294);
nand U12 (N_12,In_219,In_98);
or U13 (N_13,In_277,In_312);
or U14 (N_14,In_465,In_138);
or U15 (N_15,In_478,In_378);
nor U16 (N_16,In_204,In_330);
nand U17 (N_17,In_411,In_336);
or U18 (N_18,In_389,In_316);
nor U19 (N_19,In_383,In_169);
nor U20 (N_20,In_194,In_406);
or U21 (N_21,In_265,In_71);
nor U22 (N_22,In_34,In_327);
and U23 (N_23,In_388,In_308);
nand U24 (N_24,In_104,In_17);
or U25 (N_25,In_409,In_43);
nor U26 (N_26,In_63,In_464);
or U27 (N_27,In_248,In_129);
and U28 (N_28,In_314,In_238);
or U29 (N_29,In_150,In_333);
nor U30 (N_30,In_479,In_253);
nand U31 (N_31,In_144,In_230);
and U32 (N_32,In_289,In_353);
or U33 (N_33,In_167,In_175);
nor U34 (N_34,In_325,In_414);
nor U35 (N_35,In_247,In_293);
or U36 (N_36,In_199,In_298);
and U37 (N_37,In_59,In_447);
or U38 (N_38,In_352,In_111);
nand U39 (N_39,In_387,In_496);
and U40 (N_40,In_126,In_183);
or U41 (N_41,In_184,In_498);
nand U42 (N_42,In_142,In_400);
nor U43 (N_43,In_354,In_313);
nand U44 (N_44,In_141,In_430);
nor U45 (N_45,In_281,In_269);
nor U46 (N_46,In_153,In_405);
nand U47 (N_47,In_245,In_468);
and U48 (N_48,In_47,In_487);
nand U49 (N_49,In_223,In_173);
or U50 (N_50,In_481,In_68);
xnor U51 (N_51,In_99,In_364);
and U52 (N_52,In_342,In_365);
and U53 (N_53,In_110,In_359);
nand U54 (N_54,In_191,In_168);
nor U55 (N_55,In_160,In_62);
nor U56 (N_56,In_392,In_339);
nand U57 (N_57,In_116,In_41);
nor U58 (N_58,In_345,In_228);
or U59 (N_59,In_85,In_195);
nand U60 (N_60,In_65,In_4);
and U61 (N_61,In_444,In_182);
nand U62 (N_62,In_19,In_48);
or U63 (N_63,In_279,In_463);
nand U64 (N_64,In_459,In_384);
nand U65 (N_65,In_192,In_482);
nand U66 (N_66,In_338,In_304);
nand U67 (N_67,In_89,In_240);
and U68 (N_68,In_369,In_318);
or U69 (N_69,In_490,In_206);
nand U70 (N_70,In_480,In_340);
and U71 (N_71,In_315,In_53);
and U72 (N_72,In_448,In_210);
nand U73 (N_73,In_474,In_51);
nand U74 (N_74,In_434,In_402);
nand U75 (N_75,In_494,In_23);
or U76 (N_76,In_207,In_390);
and U77 (N_77,In_321,In_270);
nand U78 (N_78,In_418,In_462);
and U79 (N_79,In_456,In_458);
or U80 (N_80,In_288,In_107);
and U81 (N_81,In_88,In_8);
nand U82 (N_82,In_215,In_28);
and U83 (N_83,In_93,In_473);
and U84 (N_84,In_393,In_346);
and U85 (N_85,In_70,In_258);
and U86 (N_86,In_469,In_403);
nor U87 (N_87,In_139,In_9);
nand U88 (N_88,In_421,In_334);
nor U89 (N_89,In_57,In_343);
and U90 (N_90,In_29,In_348);
nand U91 (N_91,In_125,In_328);
nand U92 (N_92,In_52,In_491);
nor U93 (N_93,In_229,In_275);
nand U94 (N_94,In_164,In_407);
or U95 (N_95,In_197,In_27);
nor U96 (N_96,In_83,In_246);
nor U97 (N_97,In_170,In_44);
or U98 (N_98,In_172,In_193);
nor U99 (N_99,In_220,In_360);
or U100 (N_100,In_307,In_202);
nor U101 (N_101,In_46,In_179);
nand U102 (N_102,In_397,In_127);
nor U103 (N_103,In_401,In_355);
and U104 (N_104,In_235,In_10);
and U105 (N_105,In_66,In_130);
and U106 (N_106,In_163,In_69);
nor U107 (N_107,In_31,In_263);
or U108 (N_108,In_96,In_470);
and U109 (N_109,In_12,In_329);
or U110 (N_110,In_212,In_35);
nor U111 (N_111,In_358,In_399);
or U112 (N_112,In_178,In_274);
nor U113 (N_113,In_267,In_292);
and U114 (N_114,In_154,In_436);
and U115 (N_115,In_427,In_331);
nor U116 (N_116,In_117,In_410);
nand U117 (N_117,In_95,In_102);
nand U118 (N_118,In_276,In_361);
nor U119 (N_119,In_227,In_255);
nand U120 (N_120,In_61,In_155);
nor U121 (N_121,In_381,In_429);
nor U122 (N_122,In_14,In_203);
nand U123 (N_123,In_305,In_7);
and U124 (N_124,In_311,In_485);
nor U125 (N_125,In_349,In_32);
nand U126 (N_126,In_49,In_291);
or U127 (N_127,In_319,In_450);
nor U128 (N_128,In_146,In_33);
and U129 (N_129,In_317,In_486);
and U130 (N_130,In_140,In_357);
nand U131 (N_131,In_426,In_493);
nand U132 (N_132,In_300,In_237);
nand U133 (N_133,In_299,In_157);
and U134 (N_134,In_92,In_213);
or U135 (N_135,In_428,In_186);
nor U136 (N_136,In_72,In_368);
or U137 (N_137,In_476,In_145);
nand U138 (N_138,In_309,In_90);
and U139 (N_139,In_424,In_297);
or U140 (N_140,In_128,In_67);
nand U141 (N_141,In_81,In_416);
nor U142 (N_142,In_454,In_467);
nor U143 (N_143,In_24,In_438);
or U144 (N_144,In_20,In_114);
or U145 (N_145,In_135,In_82);
nor U146 (N_146,In_239,In_162);
nand U147 (N_147,In_423,In_382);
or U148 (N_148,In_386,In_152);
or U149 (N_149,In_218,In_341);
and U150 (N_150,In_471,In_217);
and U151 (N_151,In_477,In_376);
and U152 (N_152,In_257,In_156);
nor U153 (N_153,In_205,In_475);
or U154 (N_154,In_133,In_15);
or U155 (N_155,In_137,In_188);
nor U156 (N_156,In_439,In_420);
nor U157 (N_157,In_18,In_60);
nand U158 (N_158,In_290,In_452);
or U159 (N_159,In_233,In_42);
nand U160 (N_160,In_296,In_422);
or U161 (N_161,In_432,In_396);
nor U162 (N_162,In_363,In_385);
nand U163 (N_163,In_30,In_58);
and U164 (N_164,In_200,In_123);
or U165 (N_165,In_379,In_234);
or U166 (N_166,In_181,In_6);
nor U167 (N_167,In_495,In_408);
or U168 (N_168,In_40,In_371);
nor U169 (N_169,In_113,In_391);
xor U170 (N_170,In_185,In_105);
nand U171 (N_171,In_16,In_301);
or U172 (N_172,In_37,In_80);
nor U173 (N_173,In_76,In_134);
or U174 (N_174,In_443,In_119);
nor U175 (N_175,In_395,In_335);
nor U176 (N_176,In_174,In_3);
nor U177 (N_177,In_149,In_50);
or U178 (N_178,In_77,In_94);
or U179 (N_179,In_497,In_54);
xnor U180 (N_180,In_446,In_254);
nor U181 (N_181,In_303,In_350);
nand U182 (N_182,In_121,In_362);
nand U183 (N_183,In_86,In_380);
nand U184 (N_184,In_320,In_375);
or U185 (N_185,In_256,In_284);
nor U186 (N_186,In_241,In_73);
nor U187 (N_187,In_122,In_0);
or U188 (N_188,In_208,In_332);
and U189 (N_189,In_242,In_131);
and U190 (N_190,In_260,In_282);
nor U191 (N_191,In_244,In_366);
nor U192 (N_192,In_449,In_177);
or U193 (N_193,In_273,In_437);
or U194 (N_194,In_252,In_124);
or U195 (N_195,In_417,In_433);
nand U196 (N_196,In_243,In_250);
and U197 (N_197,In_431,In_190);
and U198 (N_198,In_278,In_147);
or U199 (N_199,In_483,In_97);
or U200 (N_200,In_326,In_373);
or U201 (N_201,In_187,In_415);
and U202 (N_202,In_413,In_492);
or U203 (N_203,In_214,In_268);
xnor U204 (N_204,In_201,In_425);
or U205 (N_205,In_143,In_21);
and U206 (N_206,In_171,In_91);
nand U207 (N_207,In_272,In_271);
and U208 (N_208,In_232,In_158);
or U209 (N_209,In_236,In_435);
nor U210 (N_210,In_372,In_5);
nor U211 (N_211,In_226,In_75);
nand U212 (N_212,In_109,In_189);
or U213 (N_213,In_280,In_262);
nand U214 (N_214,In_26,In_472);
nand U215 (N_215,In_1,In_287);
or U216 (N_216,In_347,In_451);
and U217 (N_217,In_108,In_196);
nand U218 (N_218,In_442,In_231);
or U219 (N_219,In_266,In_412);
nand U220 (N_220,In_377,In_344);
and U221 (N_221,In_302,In_488);
and U222 (N_222,In_209,In_176);
nand U223 (N_223,In_161,In_166);
and U224 (N_224,In_22,In_222);
or U225 (N_225,In_457,In_445);
or U226 (N_226,In_148,In_211);
nor U227 (N_227,In_310,In_404);
nand U228 (N_228,In_370,In_440);
nor U229 (N_229,In_337,In_484);
and U230 (N_230,In_13,In_151);
and U231 (N_231,In_159,In_461);
or U232 (N_232,In_87,In_101);
nor U233 (N_233,In_295,In_120);
and U234 (N_234,In_106,In_64);
and U235 (N_235,In_2,In_118);
or U236 (N_236,In_264,In_115);
nor U237 (N_237,In_499,In_249);
or U238 (N_238,In_251,In_180);
and U239 (N_239,In_56,In_455);
and U240 (N_240,In_466,In_261);
or U241 (N_241,In_285,In_45);
nand U242 (N_242,In_356,In_460);
nor U243 (N_243,In_38,In_11);
nand U244 (N_244,In_351,In_136);
nor U245 (N_245,In_283,In_165);
or U246 (N_246,In_74,In_132);
xnor U247 (N_247,In_100,In_398);
nand U248 (N_248,In_36,In_322);
nand U249 (N_249,In_79,In_39);
and U250 (N_250,In_136,In_196);
or U251 (N_251,In_390,In_87);
nor U252 (N_252,In_289,In_303);
nor U253 (N_253,In_293,In_3);
or U254 (N_254,In_433,In_377);
nor U255 (N_255,In_0,In_165);
or U256 (N_256,In_306,In_290);
nor U257 (N_257,In_393,In_106);
and U258 (N_258,In_285,In_235);
nand U259 (N_259,In_492,In_147);
and U260 (N_260,In_476,In_352);
and U261 (N_261,In_374,In_449);
nor U262 (N_262,In_202,In_176);
nor U263 (N_263,In_114,In_89);
nand U264 (N_264,In_128,In_435);
nor U265 (N_265,In_269,In_3);
nor U266 (N_266,In_205,In_226);
xor U267 (N_267,In_466,In_248);
and U268 (N_268,In_342,In_113);
nand U269 (N_269,In_349,In_230);
nor U270 (N_270,In_279,In_123);
and U271 (N_271,In_61,In_73);
or U272 (N_272,In_220,In_202);
or U273 (N_273,In_147,In_365);
or U274 (N_274,In_335,In_388);
nor U275 (N_275,In_69,In_432);
nand U276 (N_276,In_136,In_315);
nor U277 (N_277,In_250,In_220);
nor U278 (N_278,In_179,In_254);
and U279 (N_279,In_29,In_38);
and U280 (N_280,In_334,In_45);
and U281 (N_281,In_275,In_350);
or U282 (N_282,In_208,In_495);
and U283 (N_283,In_339,In_15);
and U284 (N_284,In_72,In_84);
nor U285 (N_285,In_461,In_123);
nand U286 (N_286,In_57,In_262);
nand U287 (N_287,In_175,In_164);
or U288 (N_288,In_93,In_226);
and U289 (N_289,In_158,In_296);
and U290 (N_290,In_131,In_377);
and U291 (N_291,In_90,In_92);
nor U292 (N_292,In_417,In_86);
or U293 (N_293,In_317,In_330);
nor U294 (N_294,In_229,In_387);
nand U295 (N_295,In_350,In_241);
nand U296 (N_296,In_400,In_236);
or U297 (N_297,In_497,In_257);
and U298 (N_298,In_276,In_466);
or U299 (N_299,In_429,In_260);
nor U300 (N_300,In_326,In_422);
or U301 (N_301,In_249,In_264);
and U302 (N_302,In_119,In_30);
and U303 (N_303,In_278,In_395);
nor U304 (N_304,In_217,In_405);
nor U305 (N_305,In_251,In_241);
nor U306 (N_306,In_176,In_259);
or U307 (N_307,In_139,In_362);
and U308 (N_308,In_227,In_74);
or U309 (N_309,In_1,In_499);
nand U310 (N_310,In_323,In_483);
nand U311 (N_311,In_37,In_40);
nor U312 (N_312,In_153,In_110);
nor U313 (N_313,In_80,In_90);
nand U314 (N_314,In_420,In_421);
nor U315 (N_315,In_35,In_93);
nor U316 (N_316,In_167,In_339);
or U317 (N_317,In_292,In_442);
nand U318 (N_318,In_228,In_396);
nand U319 (N_319,In_194,In_266);
and U320 (N_320,In_16,In_457);
and U321 (N_321,In_337,In_91);
and U322 (N_322,In_341,In_331);
and U323 (N_323,In_349,In_82);
and U324 (N_324,In_95,In_260);
or U325 (N_325,In_354,In_146);
nor U326 (N_326,In_36,In_32);
and U327 (N_327,In_58,In_218);
and U328 (N_328,In_250,In_270);
and U329 (N_329,In_111,In_45);
nor U330 (N_330,In_240,In_192);
nor U331 (N_331,In_205,In_247);
nor U332 (N_332,In_402,In_263);
nand U333 (N_333,In_257,In_28);
and U334 (N_334,In_194,In_173);
or U335 (N_335,In_376,In_136);
nand U336 (N_336,In_286,In_407);
nor U337 (N_337,In_106,In_7);
or U338 (N_338,In_381,In_267);
or U339 (N_339,In_444,In_423);
nand U340 (N_340,In_122,In_406);
or U341 (N_341,In_212,In_480);
and U342 (N_342,In_205,In_367);
and U343 (N_343,In_55,In_71);
or U344 (N_344,In_47,In_111);
nand U345 (N_345,In_210,In_0);
nor U346 (N_346,In_351,In_45);
nand U347 (N_347,In_117,In_166);
nand U348 (N_348,In_48,In_318);
nor U349 (N_349,In_120,In_342);
or U350 (N_350,In_449,In_244);
and U351 (N_351,In_104,In_281);
or U352 (N_352,In_430,In_493);
or U353 (N_353,In_152,In_221);
or U354 (N_354,In_440,In_70);
xnor U355 (N_355,In_442,In_199);
nor U356 (N_356,In_380,In_428);
nor U357 (N_357,In_366,In_159);
nand U358 (N_358,In_190,In_189);
nor U359 (N_359,In_419,In_196);
or U360 (N_360,In_261,In_373);
or U361 (N_361,In_49,In_237);
and U362 (N_362,In_367,In_287);
nand U363 (N_363,In_136,In_12);
or U364 (N_364,In_466,In_75);
and U365 (N_365,In_221,In_10);
nand U366 (N_366,In_419,In_334);
or U367 (N_367,In_484,In_398);
or U368 (N_368,In_480,In_241);
nor U369 (N_369,In_195,In_150);
or U370 (N_370,In_122,In_140);
nand U371 (N_371,In_10,In_42);
nand U372 (N_372,In_260,In_7);
nor U373 (N_373,In_411,In_223);
nand U374 (N_374,In_22,In_469);
or U375 (N_375,In_393,In_443);
or U376 (N_376,In_133,In_310);
or U377 (N_377,In_119,In_436);
and U378 (N_378,In_338,In_252);
and U379 (N_379,In_23,In_152);
or U380 (N_380,In_330,In_36);
nand U381 (N_381,In_395,In_315);
nor U382 (N_382,In_49,In_247);
and U383 (N_383,In_154,In_159);
or U384 (N_384,In_444,In_248);
nor U385 (N_385,In_11,In_461);
and U386 (N_386,In_276,In_221);
or U387 (N_387,In_450,In_384);
or U388 (N_388,In_357,In_44);
nor U389 (N_389,In_258,In_133);
nor U390 (N_390,In_23,In_205);
nor U391 (N_391,In_341,In_84);
and U392 (N_392,In_25,In_65);
nand U393 (N_393,In_351,In_368);
or U394 (N_394,In_378,In_79);
nor U395 (N_395,In_485,In_445);
or U396 (N_396,In_482,In_410);
and U397 (N_397,In_76,In_276);
or U398 (N_398,In_454,In_272);
nor U399 (N_399,In_458,In_170);
or U400 (N_400,In_223,In_236);
nand U401 (N_401,In_349,In_335);
nor U402 (N_402,In_30,In_191);
and U403 (N_403,In_112,In_122);
nor U404 (N_404,In_362,In_135);
xor U405 (N_405,In_187,In_397);
or U406 (N_406,In_171,In_349);
and U407 (N_407,In_288,In_57);
nand U408 (N_408,In_161,In_277);
nor U409 (N_409,In_86,In_322);
xor U410 (N_410,In_394,In_269);
or U411 (N_411,In_263,In_213);
and U412 (N_412,In_348,In_391);
nor U413 (N_413,In_2,In_51);
nor U414 (N_414,In_338,In_201);
nand U415 (N_415,In_26,In_221);
and U416 (N_416,In_188,In_53);
or U417 (N_417,In_107,In_362);
nor U418 (N_418,In_215,In_135);
and U419 (N_419,In_248,In_485);
nor U420 (N_420,In_42,In_499);
nor U421 (N_421,In_68,In_48);
nor U422 (N_422,In_405,In_277);
and U423 (N_423,In_18,In_280);
and U424 (N_424,In_101,In_38);
or U425 (N_425,In_199,In_132);
nor U426 (N_426,In_127,In_71);
or U427 (N_427,In_389,In_32);
and U428 (N_428,In_371,In_97);
nand U429 (N_429,In_362,In_345);
nor U430 (N_430,In_104,In_403);
nand U431 (N_431,In_361,In_389);
nand U432 (N_432,In_386,In_94);
and U433 (N_433,In_158,In_15);
nor U434 (N_434,In_293,In_67);
nor U435 (N_435,In_216,In_277);
or U436 (N_436,In_283,In_138);
or U437 (N_437,In_69,In_255);
nand U438 (N_438,In_255,In_186);
nor U439 (N_439,In_305,In_164);
and U440 (N_440,In_176,In_255);
nand U441 (N_441,In_277,In_461);
and U442 (N_442,In_61,In_239);
and U443 (N_443,In_473,In_136);
or U444 (N_444,In_329,In_475);
nor U445 (N_445,In_371,In_210);
nor U446 (N_446,In_412,In_145);
nor U447 (N_447,In_86,In_288);
or U448 (N_448,In_81,In_401);
nand U449 (N_449,In_67,In_431);
nor U450 (N_450,In_64,In_27);
nor U451 (N_451,In_173,In_356);
and U452 (N_452,In_336,In_358);
nand U453 (N_453,In_400,In_260);
or U454 (N_454,In_12,In_457);
or U455 (N_455,In_348,In_288);
or U456 (N_456,In_411,In_364);
and U457 (N_457,In_383,In_259);
and U458 (N_458,In_378,In_437);
or U459 (N_459,In_468,In_332);
and U460 (N_460,In_342,In_272);
or U461 (N_461,In_88,In_49);
and U462 (N_462,In_253,In_225);
nand U463 (N_463,In_306,In_203);
or U464 (N_464,In_82,In_367);
or U465 (N_465,In_444,In_126);
nor U466 (N_466,In_310,In_253);
nand U467 (N_467,In_282,In_378);
or U468 (N_468,In_32,In_265);
nand U469 (N_469,In_323,In_54);
nand U470 (N_470,In_416,In_50);
or U471 (N_471,In_49,In_314);
nand U472 (N_472,In_202,In_316);
nand U473 (N_473,In_314,In_54);
nor U474 (N_474,In_230,In_195);
nand U475 (N_475,In_416,In_343);
nor U476 (N_476,In_115,In_399);
or U477 (N_477,In_335,In_445);
nor U478 (N_478,In_25,In_471);
or U479 (N_479,In_482,In_182);
and U480 (N_480,In_408,In_437);
and U481 (N_481,In_334,In_448);
and U482 (N_482,In_209,In_319);
nor U483 (N_483,In_324,In_140);
or U484 (N_484,In_294,In_283);
or U485 (N_485,In_443,In_45);
nand U486 (N_486,In_130,In_483);
or U487 (N_487,In_12,In_498);
nor U488 (N_488,In_236,In_78);
nand U489 (N_489,In_256,In_277);
or U490 (N_490,In_379,In_322);
nor U491 (N_491,In_70,In_433);
nand U492 (N_492,In_421,In_291);
nor U493 (N_493,In_273,In_467);
nand U494 (N_494,In_236,In_173);
nor U495 (N_495,In_101,In_113);
nand U496 (N_496,In_402,In_302);
or U497 (N_497,In_69,In_20);
and U498 (N_498,In_95,In_466);
nand U499 (N_499,In_186,In_113);
or U500 (N_500,N_453,N_21);
nand U501 (N_501,N_199,N_348);
nand U502 (N_502,N_256,N_143);
nand U503 (N_503,N_253,N_270);
nand U504 (N_504,N_52,N_162);
and U505 (N_505,N_221,N_167);
and U506 (N_506,N_272,N_191);
nand U507 (N_507,N_323,N_364);
nor U508 (N_508,N_249,N_118);
and U509 (N_509,N_189,N_28);
and U510 (N_510,N_466,N_154);
or U511 (N_511,N_289,N_438);
nand U512 (N_512,N_184,N_6);
or U513 (N_513,N_10,N_461);
and U514 (N_514,N_140,N_59);
nor U515 (N_515,N_193,N_48);
nor U516 (N_516,N_345,N_311);
and U517 (N_517,N_82,N_316);
nand U518 (N_518,N_245,N_42);
and U519 (N_519,N_246,N_111);
or U520 (N_520,N_57,N_196);
or U521 (N_521,N_240,N_350);
nand U522 (N_522,N_290,N_414);
nand U523 (N_523,N_116,N_460);
xnor U524 (N_524,N_370,N_150);
or U525 (N_525,N_352,N_122);
and U526 (N_526,N_479,N_343);
and U527 (N_527,N_340,N_239);
nand U528 (N_528,N_267,N_296);
nand U529 (N_529,N_477,N_424);
nand U530 (N_530,N_69,N_379);
or U531 (N_531,N_213,N_197);
nor U532 (N_532,N_12,N_102);
and U533 (N_533,N_106,N_9);
nand U534 (N_534,N_230,N_268);
or U535 (N_535,N_332,N_254);
and U536 (N_536,N_11,N_359);
nand U537 (N_537,N_277,N_74);
nand U538 (N_538,N_94,N_306);
nand U539 (N_539,N_41,N_161);
and U540 (N_540,N_470,N_223);
and U541 (N_541,N_139,N_329);
or U542 (N_542,N_131,N_297);
nor U543 (N_543,N_187,N_99);
and U544 (N_544,N_173,N_317);
nand U545 (N_545,N_462,N_412);
nor U546 (N_546,N_385,N_284);
nor U547 (N_547,N_381,N_30);
nand U548 (N_548,N_417,N_200);
nor U549 (N_549,N_91,N_2);
xor U550 (N_550,N_353,N_307);
nor U551 (N_551,N_107,N_105);
nor U552 (N_552,N_121,N_55);
nor U553 (N_553,N_115,N_32);
nand U554 (N_554,N_310,N_233);
and U555 (N_555,N_293,N_391);
and U556 (N_556,N_336,N_84);
nor U557 (N_557,N_47,N_229);
or U558 (N_558,N_67,N_228);
nand U559 (N_559,N_170,N_280);
and U560 (N_560,N_160,N_413);
or U561 (N_561,N_16,N_465);
nor U562 (N_562,N_401,N_361);
nor U563 (N_563,N_247,N_215);
nand U564 (N_564,N_279,N_400);
xor U565 (N_565,N_451,N_373);
or U566 (N_566,N_78,N_125);
xnor U567 (N_567,N_220,N_264);
nand U568 (N_568,N_34,N_185);
nor U569 (N_569,N_365,N_75);
and U570 (N_570,N_93,N_494);
nand U571 (N_571,N_367,N_302);
nand U572 (N_572,N_4,N_19);
or U573 (N_573,N_371,N_40);
nor U574 (N_574,N_375,N_252);
and U575 (N_575,N_175,N_190);
nor U576 (N_576,N_396,N_88);
or U577 (N_577,N_449,N_305);
nor U578 (N_578,N_337,N_135);
nor U579 (N_579,N_398,N_130);
or U580 (N_580,N_126,N_266);
nand U581 (N_581,N_282,N_321);
or U582 (N_582,N_467,N_114);
nor U583 (N_583,N_404,N_448);
or U584 (N_584,N_231,N_156);
and U585 (N_585,N_104,N_238);
nor U586 (N_586,N_440,N_100);
nand U587 (N_587,N_142,N_475);
nand U588 (N_588,N_444,N_258);
or U589 (N_589,N_169,N_144);
nand U590 (N_590,N_73,N_219);
or U591 (N_591,N_437,N_402);
and U592 (N_592,N_469,N_109);
nand U593 (N_593,N_368,N_410);
nor U594 (N_594,N_124,N_237);
and U595 (N_595,N_495,N_183);
nand U596 (N_596,N_455,N_320);
nand U597 (N_597,N_314,N_26);
xor U598 (N_598,N_145,N_20);
nor U599 (N_599,N_452,N_186);
or U600 (N_600,N_203,N_129);
nand U601 (N_601,N_274,N_148);
xor U602 (N_602,N_441,N_355);
nand U603 (N_603,N_342,N_351);
and U604 (N_604,N_387,N_39);
nor U605 (N_605,N_416,N_499);
nor U606 (N_606,N_374,N_294);
and U607 (N_607,N_159,N_480);
xnor U608 (N_608,N_201,N_7);
and U609 (N_609,N_79,N_210);
and U610 (N_610,N_117,N_76);
and U611 (N_611,N_383,N_35);
or U612 (N_612,N_110,N_285);
nand U613 (N_613,N_346,N_147);
and U614 (N_614,N_435,N_224);
nand U615 (N_615,N_360,N_134);
nor U616 (N_616,N_149,N_431);
nand U617 (N_617,N_308,N_113);
or U618 (N_618,N_51,N_386);
or U619 (N_619,N_474,N_292);
nor U620 (N_620,N_168,N_376);
nor U621 (N_621,N_283,N_303);
nor U622 (N_622,N_384,N_132);
nor U623 (N_623,N_439,N_457);
nand U624 (N_624,N_459,N_407);
or U625 (N_625,N_250,N_216);
or U626 (N_626,N_255,N_334);
or U627 (N_627,N_15,N_206);
xnor U628 (N_628,N_212,N_328);
and U629 (N_629,N_422,N_456);
nand U630 (N_630,N_71,N_146);
nand U631 (N_631,N_331,N_463);
nand U632 (N_632,N_176,N_56);
or U633 (N_633,N_259,N_64);
or U634 (N_634,N_366,N_300);
and U635 (N_635,N_66,N_5);
nor U636 (N_636,N_60,N_61);
nand U637 (N_637,N_464,N_86);
xor U638 (N_638,N_265,N_324);
or U639 (N_639,N_299,N_443);
nor U640 (N_640,N_13,N_486);
nor U641 (N_641,N_46,N_498);
and U642 (N_642,N_476,N_298);
nand U643 (N_643,N_442,N_338);
or U644 (N_644,N_271,N_421);
nand U645 (N_645,N_204,N_218);
nor U646 (N_646,N_242,N_138);
nand U647 (N_647,N_195,N_38);
nand U648 (N_648,N_36,N_432);
nor U649 (N_649,N_318,N_166);
nand U650 (N_650,N_3,N_411);
nor U651 (N_651,N_63,N_497);
or U652 (N_652,N_25,N_81);
nor U653 (N_653,N_313,N_488);
and U654 (N_654,N_95,N_363);
nor U655 (N_655,N_262,N_406);
and U656 (N_656,N_37,N_22);
nand U657 (N_657,N_235,N_485);
nor U658 (N_658,N_214,N_136);
or U659 (N_659,N_172,N_58);
nor U660 (N_660,N_49,N_236);
nand U661 (N_661,N_399,N_397);
and U662 (N_662,N_188,N_65);
and U663 (N_663,N_487,N_344);
nor U664 (N_664,N_127,N_244);
nand U665 (N_665,N_98,N_427);
or U666 (N_666,N_388,N_251);
nand U667 (N_667,N_18,N_426);
nor U668 (N_668,N_1,N_243);
or U669 (N_669,N_33,N_362);
or U670 (N_670,N_96,N_119);
or U671 (N_671,N_207,N_202);
and U672 (N_672,N_261,N_83);
or U673 (N_673,N_354,N_420);
and U674 (N_674,N_378,N_31);
and U675 (N_675,N_392,N_232);
nor U676 (N_676,N_70,N_403);
and U677 (N_677,N_434,N_304);
nor U678 (N_678,N_45,N_80);
or U679 (N_679,N_429,N_481);
and U680 (N_680,N_415,N_90);
nand U681 (N_681,N_430,N_209);
or U682 (N_682,N_377,N_181);
nor U683 (N_683,N_44,N_369);
nand U684 (N_684,N_205,N_85);
and U685 (N_685,N_490,N_211);
nor U686 (N_686,N_327,N_405);
and U687 (N_687,N_301,N_155);
or U688 (N_688,N_447,N_319);
and U689 (N_689,N_260,N_217);
nor U690 (N_690,N_263,N_89);
and U691 (N_691,N_483,N_0);
and U692 (N_692,N_62,N_491);
and U693 (N_693,N_315,N_77);
and U694 (N_694,N_312,N_178);
or U695 (N_695,N_182,N_395);
nand U696 (N_696,N_14,N_112);
nand U697 (N_697,N_288,N_54);
nor U698 (N_698,N_257,N_436);
and U699 (N_699,N_341,N_23);
and U700 (N_700,N_484,N_468);
nor U701 (N_701,N_408,N_380);
nor U702 (N_702,N_123,N_50);
or U703 (N_703,N_8,N_423);
nor U704 (N_704,N_241,N_339);
and U705 (N_705,N_68,N_128);
nand U706 (N_706,N_248,N_493);
and U707 (N_707,N_278,N_108);
nor U708 (N_708,N_322,N_87);
and U709 (N_709,N_287,N_291);
or U710 (N_710,N_120,N_496);
or U711 (N_711,N_372,N_389);
nand U712 (N_712,N_393,N_492);
and U713 (N_713,N_171,N_309);
or U714 (N_714,N_174,N_275);
and U715 (N_715,N_164,N_347);
nand U716 (N_716,N_409,N_433);
or U717 (N_717,N_137,N_349);
or U718 (N_718,N_222,N_92);
and U719 (N_719,N_458,N_53);
or U720 (N_720,N_234,N_97);
or U721 (N_721,N_152,N_482);
nand U722 (N_722,N_418,N_151);
and U723 (N_723,N_194,N_177);
xor U724 (N_724,N_163,N_276);
nor U725 (N_725,N_390,N_153);
or U726 (N_726,N_419,N_27);
nor U727 (N_727,N_180,N_24);
nand U728 (N_728,N_101,N_445);
nor U729 (N_729,N_43,N_17);
xor U730 (N_730,N_157,N_450);
nor U731 (N_731,N_326,N_141);
or U732 (N_732,N_269,N_446);
nor U733 (N_733,N_394,N_192);
nand U734 (N_734,N_158,N_227);
nand U735 (N_735,N_330,N_333);
nor U736 (N_736,N_358,N_478);
and U737 (N_737,N_356,N_382);
and U738 (N_738,N_29,N_133);
nor U739 (N_739,N_103,N_286);
xor U740 (N_740,N_473,N_454);
nor U741 (N_741,N_428,N_335);
and U742 (N_742,N_273,N_425);
or U743 (N_743,N_471,N_165);
nor U744 (N_744,N_325,N_226);
nand U745 (N_745,N_208,N_198);
nand U746 (N_746,N_357,N_179);
nor U747 (N_747,N_72,N_295);
or U748 (N_748,N_472,N_489);
nand U749 (N_749,N_281,N_225);
nor U750 (N_750,N_244,N_351);
and U751 (N_751,N_495,N_156);
and U752 (N_752,N_210,N_369);
nor U753 (N_753,N_325,N_149);
and U754 (N_754,N_45,N_477);
nor U755 (N_755,N_295,N_213);
or U756 (N_756,N_287,N_21);
and U757 (N_757,N_361,N_54);
or U758 (N_758,N_137,N_495);
and U759 (N_759,N_2,N_457);
and U760 (N_760,N_421,N_201);
nor U761 (N_761,N_308,N_304);
and U762 (N_762,N_420,N_485);
or U763 (N_763,N_191,N_155);
nor U764 (N_764,N_169,N_372);
nor U765 (N_765,N_31,N_241);
nand U766 (N_766,N_199,N_339);
nor U767 (N_767,N_494,N_456);
nor U768 (N_768,N_464,N_156);
or U769 (N_769,N_241,N_324);
and U770 (N_770,N_248,N_451);
nand U771 (N_771,N_262,N_428);
and U772 (N_772,N_137,N_426);
or U773 (N_773,N_372,N_152);
or U774 (N_774,N_279,N_202);
and U775 (N_775,N_232,N_19);
nand U776 (N_776,N_409,N_487);
and U777 (N_777,N_381,N_331);
and U778 (N_778,N_174,N_91);
and U779 (N_779,N_94,N_325);
xnor U780 (N_780,N_324,N_432);
nor U781 (N_781,N_366,N_155);
nor U782 (N_782,N_494,N_155);
nor U783 (N_783,N_170,N_379);
and U784 (N_784,N_132,N_174);
and U785 (N_785,N_17,N_206);
and U786 (N_786,N_172,N_369);
and U787 (N_787,N_362,N_447);
and U788 (N_788,N_378,N_362);
nand U789 (N_789,N_454,N_447);
and U790 (N_790,N_423,N_310);
and U791 (N_791,N_474,N_328);
nor U792 (N_792,N_306,N_369);
or U793 (N_793,N_291,N_263);
or U794 (N_794,N_66,N_352);
nor U795 (N_795,N_418,N_88);
nand U796 (N_796,N_217,N_9);
nor U797 (N_797,N_18,N_301);
nor U798 (N_798,N_277,N_121);
nor U799 (N_799,N_327,N_459);
nand U800 (N_800,N_243,N_275);
or U801 (N_801,N_143,N_229);
nand U802 (N_802,N_341,N_11);
nand U803 (N_803,N_443,N_87);
or U804 (N_804,N_378,N_352);
nand U805 (N_805,N_407,N_260);
or U806 (N_806,N_163,N_78);
or U807 (N_807,N_73,N_319);
and U808 (N_808,N_262,N_228);
or U809 (N_809,N_261,N_190);
nor U810 (N_810,N_62,N_168);
or U811 (N_811,N_121,N_138);
or U812 (N_812,N_2,N_380);
or U813 (N_813,N_453,N_380);
nand U814 (N_814,N_164,N_178);
nand U815 (N_815,N_492,N_29);
nor U816 (N_816,N_281,N_210);
nand U817 (N_817,N_310,N_493);
nand U818 (N_818,N_411,N_107);
nand U819 (N_819,N_101,N_388);
xnor U820 (N_820,N_303,N_12);
xnor U821 (N_821,N_274,N_134);
or U822 (N_822,N_248,N_308);
nor U823 (N_823,N_65,N_367);
and U824 (N_824,N_27,N_280);
nor U825 (N_825,N_333,N_171);
nand U826 (N_826,N_493,N_129);
and U827 (N_827,N_4,N_100);
or U828 (N_828,N_472,N_275);
or U829 (N_829,N_380,N_486);
nor U830 (N_830,N_458,N_467);
nand U831 (N_831,N_363,N_486);
nor U832 (N_832,N_328,N_426);
nand U833 (N_833,N_296,N_192);
nor U834 (N_834,N_296,N_357);
nor U835 (N_835,N_307,N_422);
nor U836 (N_836,N_416,N_306);
nor U837 (N_837,N_460,N_129);
and U838 (N_838,N_398,N_286);
nand U839 (N_839,N_296,N_123);
or U840 (N_840,N_154,N_230);
and U841 (N_841,N_174,N_217);
nand U842 (N_842,N_246,N_339);
and U843 (N_843,N_31,N_265);
and U844 (N_844,N_430,N_206);
nor U845 (N_845,N_161,N_258);
xor U846 (N_846,N_120,N_433);
and U847 (N_847,N_22,N_240);
xor U848 (N_848,N_419,N_90);
nor U849 (N_849,N_270,N_413);
nor U850 (N_850,N_226,N_453);
and U851 (N_851,N_81,N_113);
and U852 (N_852,N_379,N_190);
and U853 (N_853,N_308,N_95);
nor U854 (N_854,N_433,N_298);
and U855 (N_855,N_39,N_474);
or U856 (N_856,N_72,N_143);
nand U857 (N_857,N_203,N_464);
and U858 (N_858,N_438,N_309);
or U859 (N_859,N_34,N_44);
or U860 (N_860,N_90,N_139);
nor U861 (N_861,N_337,N_220);
and U862 (N_862,N_128,N_193);
nor U863 (N_863,N_474,N_168);
or U864 (N_864,N_156,N_466);
nand U865 (N_865,N_344,N_484);
or U866 (N_866,N_334,N_414);
nor U867 (N_867,N_91,N_342);
nor U868 (N_868,N_56,N_213);
nand U869 (N_869,N_487,N_443);
nand U870 (N_870,N_318,N_286);
and U871 (N_871,N_366,N_403);
and U872 (N_872,N_150,N_272);
nor U873 (N_873,N_100,N_458);
and U874 (N_874,N_64,N_14);
nor U875 (N_875,N_347,N_167);
or U876 (N_876,N_333,N_86);
or U877 (N_877,N_380,N_186);
and U878 (N_878,N_106,N_113);
nand U879 (N_879,N_182,N_379);
nor U880 (N_880,N_395,N_405);
and U881 (N_881,N_76,N_484);
nand U882 (N_882,N_44,N_167);
nor U883 (N_883,N_142,N_416);
or U884 (N_884,N_204,N_265);
or U885 (N_885,N_105,N_331);
xor U886 (N_886,N_457,N_201);
and U887 (N_887,N_220,N_225);
and U888 (N_888,N_486,N_495);
nand U889 (N_889,N_161,N_13);
or U890 (N_890,N_17,N_38);
and U891 (N_891,N_497,N_28);
and U892 (N_892,N_232,N_354);
or U893 (N_893,N_469,N_248);
or U894 (N_894,N_439,N_99);
nor U895 (N_895,N_195,N_135);
or U896 (N_896,N_450,N_360);
nor U897 (N_897,N_94,N_368);
nand U898 (N_898,N_395,N_32);
nor U899 (N_899,N_274,N_67);
nor U900 (N_900,N_310,N_389);
and U901 (N_901,N_111,N_303);
or U902 (N_902,N_229,N_207);
or U903 (N_903,N_34,N_191);
nor U904 (N_904,N_70,N_63);
nor U905 (N_905,N_411,N_204);
or U906 (N_906,N_78,N_17);
and U907 (N_907,N_398,N_219);
or U908 (N_908,N_410,N_103);
nor U909 (N_909,N_109,N_328);
nor U910 (N_910,N_62,N_50);
nand U911 (N_911,N_248,N_326);
nand U912 (N_912,N_57,N_389);
and U913 (N_913,N_182,N_353);
nor U914 (N_914,N_224,N_239);
nor U915 (N_915,N_71,N_26);
nor U916 (N_916,N_320,N_339);
and U917 (N_917,N_293,N_66);
or U918 (N_918,N_404,N_92);
nor U919 (N_919,N_27,N_31);
nor U920 (N_920,N_139,N_478);
nand U921 (N_921,N_85,N_121);
or U922 (N_922,N_397,N_352);
nand U923 (N_923,N_8,N_72);
nand U924 (N_924,N_301,N_468);
and U925 (N_925,N_280,N_420);
nand U926 (N_926,N_19,N_405);
or U927 (N_927,N_180,N_447);
or U928 (N_928,N_277,N_292);
nand U929 (N_929,N_386,N_354);
and U930 (N_930,N_405,N_41);
or U931 (N_931,N_379,N_119);
and U932 (N_932,N_180,N_474);
nor U933 (N_933,N_230,N_187);
or U934 (N_934,N_95,N_167);
or U935 (N_935,N_296,N_491);
and U936 (N_936,N_396,N_267);
or U937 (N_937,N_303,N_198);
nand U938 (N_938,N_315,N_200);
or U939 (N_939,N_140,N_389);
or U940 (N_940,N_255,N_464);
nand U941 (N_941,N_242,N_350);
nor U942 (N_942,N_38,N_109);
nor U943 (N_943,N_276,N_434);
nor U944 (N_944,N_83,N_482);
nor U945 (N_945,N_447,N_421);
nor U946 (N_946,N_369,N_67);
or U947 (N_947,N_476,N_295);
and U948 (N_948,N_61,N_383);
or U949 (N_949,N_410,N_369);
nor U950 (N_950,N_63,N_279);
and U951 (N_951,N_219,N_207);
nor U952 (N_952,N_241,N_244);
and U953 (N_953,N_407,N_139);
and U954 (N_954,N_162,N_55);
nand U955 (N_955,N_204,N_462);
and U956 (N_956,N_446,N_94);
nand U957 (N_957,N_362,N_131);
nand U958 (N_958,N_318,N_156);
and U959 (N_959,N_450,N_497);
and U960 (N_960,N_352,N_298);
and U961 (N_961,N_170,N_213);
or U962 (N_962,N_206,N_483);
or U963 (N_963,N_226,N_98);
nand U964 (N_964,N_443,N_356);
nand U965 (N_965,N_442,N_303);
and U966 (N_966,N_12,N_108);
and U967 (N_967,N_81,N_491);
or U968 (N_968,N_211,N_36);
and U969 (N_969,N_209,N_163);
nand U970 (N_970,N_195,N_399);
or U971 (N_971,N_147,N_138);
nor U972 (N_972,N_445,N_309);
nor U973 (N_973,N_347,N_120);
or U974 (N_974,N_16,N_161);
nor U975 (N_975,N_449,N_81);
nand U976 (N_976,N_85,N_236);
nor U977 (N_977,N_465,N_186);
and U978 (N_978,N_433,N_140);
or U979 (N_979,N_53,N_471);
and U980 (N_980,N_285,N_419);
or U981 (N_981,N_441,N_138);
or U982 (N_982,N_409,N_257);
or U983 (N_983,N_110,N_3);
nor U984 (N_984,N_458,N_238);
nor U985 (N_985,N_205,N_166);
nor U986 (N_986,N_201,N_57);
and U987 (N_987,N_154,N_99);
nor U988 (N_988,N_178,N_277);
nor U989 (N_989,N_55,N_415);
nand U990 (N_990,N_474,N_350);
and U991 (N_991,N_92,N_383);
and U992 (N_992,N_120,N_108);
nand U993 (N_993,N_315,N_372);
nor U994 (N_994,N_372,N_361);
nand U995 (N_995,N_327,N_323);
nor U996 (N_996,N_62,N_451);
nand U997 (N_997,N_125,N_481);
nand U998 (N_998,N_312,N_22);
and U999 (N_999,N_420,N_192);
nor U1000 (N_1000,N_679,N_954);
and U1001 (N_1001,N_896,N_561);
nor U1002 (N_1002,N_784,N_553);
nand U1003 (N_1003,N_835,N_732);
nand U1004 (N_1004,N_751,N_520);
nand U1005 (N_1005,N_841,N_869);
nand U1006 (N_1006,N_792,N_596);
nand U1007 (N_1007,N_539,N_535);
and U1008 (N_1008,N_863,N_965);
nand U1009 (N_1009,N_904,N_509);
nand U1010 (N_1010,N_580,N_708);
nor U1011 (N_1011,N_939,N_583);
nor U1012 (N_1012,N_955,N_952);
nand U1013 (N_1013,N_570,N_547);
nand U1014 (N_1014,N_603,N_614);
nand U1015 (N_1015,N_534,N_978);
nand U1016 (N_1016,N_824,N_943);
or U1017 (N_1017,N_971,N_789);
nand U1018 (N_1018,N_879,N_659);
xnor U1019 (N_1019,N_825,N_707);
and U1020 (N_1020,N_893,N_834);
and U1021 (N_1021,N_804,N_791);
nor U1022 (N_1022,N_586,N_909);
and U1023 (N_1023,N_611,N_917);
nor U1024 (N_1024,N_656,N_836);
nor U1025 (N_1025,N_742,N_655);
nand U1026 (N_1026,N_683,N_953);
nor U1027 (N_1027,N_860,N_832);
xnor U1028 (N_1028,N_667,N_619);
and U1029 (N_1029,N_672,N_950);
or U1030 (N_1030,N_724,N_768);
or U1031 (N_1031,N_563,N_858);
and U1032 (N_1032,N_712,N_981);
and U1033 (N_1033,N_517,N_692);
or U1034 (N_1034,N_541,N_526);
nor U1035 (N_1035,N_867,N_566);
nor U1036 (N_1036,N_865,N_786);
nor U1037 (N_1037,N_976,N_921);
and U1038 (N_1038,N_741,N_967);
nand U1039 (N_1039,N_937,N_951);
or U1040 (N_1040,N_963,N_959);
and U1041 (N_1041,N_633,N_703);
nand U1042 (N_1042,N_891,N_711);
nand U1043 (N_1043,N_555,N_653);
and U1044 (N_1044,N_793,N_890);
or U1045 (N_1045,N_723,N_531);
nor U1046 (N_1046,N_969,N_750);
nand U1047 (N_1047,N_812,N_630);
or U1048 (N_1048,N_739,N_598);
or U1049 (N_1049,N_805,N_722);
or U1050 (N_1050,N_765,N_588);
or U1051 (N_1051,N_994,N_974);
nand U1052 (N_1052,N_901,N_864);
nand U1053 (N_1053,N_878,N_601);
or U1054 (N_1054,N_887,N_859);
or U1055 (N_1055,N_519,N_648);
nor U1056 (N_1056,N_913,N_575);
nand U1057 (N_1057,N_689,N_914);
or U1058 (N_1058,N_626,N_629);
nor U1059 (N_1059,N_717,N_735);
and U1060 (N_1060,N_770,N_502);
or U1061 (N_1061,N_594,N_747);
nor U1062 (N_1062,N_844,N_899);
or U1063 (N_1063,N_787,N_513);
or U1064 (N_1064,N_918,N_622);
or U1065 (N_1065,N_565,N_966);
and U1066 (N_1066,N_837,N_745);
or U1067 (N_1067,N_938,N_688);
nand U1068 (N_1068,N_577,N_886);
nor U1069 (N_1069,N_854,N_972);
or U1070 (N_1070,N_640,N_797);
and U1071 (N_1071,N_846,N_521);
xnor U1072 (N_1072,N_856,N_884);
nand U1073 (N_1073,N_602,N_500);
xnor U1074 (N_1074,N_660,N_523);
or U1075 (N_1075,N_713,N_593);
or U1076 (N_1076,N_536,N_850);
nor U1077 (N_1077,N_801,N_961);
nand U1078 (N_1078,N_646,N_962);
nand U1079 (N_1079,N_810,N_554);
or U1080 (N_1080,N_999,N_610);
nor U1081 (N_1081,N_868,N_840);
or U1082 (N_1082,N_933,N_820);
nand U1083 (N_1083,N_649,N_729);
nor U1084 (N_1084,N_839,N_720);
or U1085 (N_1085,N_644,N_697);
nor U1086 (N_1086,N_774,N_525);
nand U1087 (N_1087,N_682,N_613);
or U1088 (N_1088,N_908,N_631);
and U1089 (N_1089,N_669,N_877);
or U1090 (N_1090,N_930,N_993);
nor U1091 (N_1091,N_743,N_727);
or U1092 (N_1092,N_785,N_942);
nor U1093 (N_1093,N_529,N_627);
or U1094 (N_1094,N_731,N_540);
nand U1095 (N_1095,N_866,N_756);
or U1096 (N_1096,N_730,N_946);
nor U1097 (N_1097,N_728,N_960);
nand U1098 (N_1098,N_748,N_816);
nand U1099 (N_1099,N_773,N_763);
nor U1100 (N_1100,N_924,N_704);
xnor U1101 (N_1101,N_690,N_737);
or U1102 (N_1102,N_826,N_615);
nand U1103 (N_1103,N_504,N_678);
nor U1104 (N_1104,N_783,N_906);
nor U1105 (N_1105,N_709,N_795);
nor U1106 (N_1106,N_503,N_935);
nor U1107 (N_1107,N_624,N_542);
nor U1108 (N_1108,N_638,N_823);
or U1109 (N_1109,N_685,N_986);
and U1110 (N_1110,N_803,N_929);
or U1111 (N_1111,N_964,N_873);
nand U1112 (N_1112,N_721,N_518);
nor U1113 (N_1113,N_579,N_932);
and U1114 (N_1114,N_842,N_754);
or U1115 (N_1115,N_632,N_515);
and U1116 (N_1116,N_661,N_550);
and U1117 (N_1117,N_771,N_802);
or U1118 (N_1118,N_777,N_944);
or U1119 (N_1119,N_919,N_949);
or U1120 (N_1120,N_853,N_818);
nor U1121 (N_1121,N_794,N_551);
or U1122 (N_1122,N_880,N_651);
or U1123 (N_1123,N_980,N_923);
or U1124 (N_1124,N_905,N_907);
and U1125 (N_1125,N_699,N_714);
nor U1126 (N_1126,N_746,N_883);
and U1127 (N_1127,N_581,N_926);
or U1128 (N_1128,N_779,N_664);
and U1129 (N_1129,N_900,N_817);
nor U1130 (N_1130,N_984,N_861);
and U1131 (N_1131,N_996,N_696);
and U1132 (N_1132,N_548,N_894);
nor U1133 (N_1133,N_670,N_920);
nand U1134 (N_1134,N_556,N_940);
nor U1135 (N_1135,N_821,N_781);
nor U1136 (N_1136,N_991,N_885);
nor U1137 (N_1137,N_569,N_616);
and U1138 (N_1138,N_645,N_505);
and U1139 (N_1139,N_617,N_589);
nand U1140 (N_1140,N_927,N_501);
nand U1141 (N_1141,N_874,N_813);
nand U1142 (N_1142,N_508,N_780);
and U1143 (N_1143,N_912,N_686);
nand U1144 (N_1144,N_665,N_985);
xnor U1145 (N_1145,N_642,N_764);
and U1146 (N_1146,N_695,N_510);
nand U1147 (N_1147,N_668,N_560);
xnor U1148 (N_1148,N_871,N_733);
nand U1149 (N_1149,N_538,N_641);
nor U1150 (N_1150,N_808,N_576);
and U1151 (N_1151,N_990,N_769);
nor U1152 (N_1152,N_778,N_989);
or U1153 (N_1153,N_574,N_691);
or U1154 (N_1154,N_571,N_968);
and U1155 (N_1155,N_544,N_736);
nand U1156 (N_1156,N_931,N_847);
or U1157 (N_1157,N_922,N_992);
nor U1158 (N_1158,N_895,N_753);
and U1159 (N_1159,N_684,N_654);
or U1160 (N_1160,N_928,N_957);
or U1161 (N_1161,N_822,N_995);
and U1162 (N_1162,N_620,N_533);
or U1163 (N_1163,N_755,N_814);
nand U1164 (N_1164,N_910,N_815);
nor U1165 (N_1165,N_752,N_693);
nor U1166 (N_1166,N_591,N_903);
and U1167 (N_1167,N_809,N_658);
nand U1168 (N_1168,N_934,N_546);
or U1169 (N_1169,N_558,N_639);
nand U1170 (N_1170,N_892,N_898);
and U1171 (N_1171,N_700,N_605);
nor U1172 (N_1172,N_681,N_872);
or U1173 (N_1173,N_543,N_979);
or U1174 (N_1174,N_911,N_652);
nor U1175 (N_1175,N_775,N_761);
nand U1176 (N_1176,N_875,N_549);
nor U1177 (N_1177,N_587,N_609);
nor U1178 (N_1178,N_915,N_608);
nand U1179 (N_1179,N_799,N_719);
or U1180 (N_1180,N_637,N_600);
xnor U1181 (N_1181,N_760,N_798);
nand U1182 (N_1182,N_862,N_947);
or U1183 (N_1183,N_582,N_857);
nor U1184 (N_1184,N_516,N_595);
or U1185 (N_1185,N_557,N_870);
or U1186 (N_1186,N_572,N_592);
nand U1187 (N_1187,N_843,N_527);
nand U1188 (N_1188,N_776,N_782);
nand U1189 (N_1189,N_807,N_522);
xor U1190 (N_1190,N_706,N_982);
nand U1191 (N_1191,N_897,N_694);
and U1192 (N_1192,N_562,N_568);
and U1193 (N_1193,N_788,N_749);
or U1194 (N_1194,N_811,N_806);
or U1195 (N_1195,N_833,N_671);
nor U1196 (N_1196,N_559,N_925);
or U1197 (N_1197,N_607,N_636);
or U1198 (N_1198,N_552,N_848);
nor U1199 (N_1199,N_590,N_941);
or U1200 (N_1200,N_882,N_772);
nand U1201 (N_1201,N_757,N_584);
nand U1202 (N_1202,N_710,N_948);
and U1203 (N_1203,N_830,N_829);
and U1204 (N_1204,N_657,N_507);
nand U1205 (N_1205,N_698,N_675);
nor U1206 (N_1206,N_734,N_511);
nor U1207 (N_1207,N_725,N_936);
or U1208 (N_1208,N_852,N_997);
and U1209 (N_1209,N_604,N_945);
and U1210 (N_1210,N_650,N_888);
nor U1211 (N_1211,N_674,N_758);
and U1212 (N_1212,N_767,N_881);
and U1213 (N_1213,N_687,N_702);
nor U1214 (N_1214,N_514,N_666);
and U1215 (N_1215,N_718,N_796);
nor U1216 (N_1216,N_977,N_628);
and U1217 (N_1217,N_987,N_889);
or U1218 (N_1218,N_530,N_744);
nand U1219 (N_1219,N_762,N_970);
nand U1220 (N_1220,N_635,N_983);
xnor U1221 (N_1221,N_599,N_738);
nand U1222 (N_1222,N_573,N_790);
nand U1223 (N_1223,N_975,N_726);
and U1224 (N_1224,N_623,N_612);
nand U1225 (N_1225,N_851,N_701);
nor U1226 (N_1226,N_537,N_876);
or U1227 (N_1227,N_828,N_621);
and U1228 (N_1228,N_827,N_973);
xor U1229 (N_1229,N_800,N_705);
nand U1230 (N_1230,N_606,N_958);
or U1231 (N_1231,N_715,N_634);
nor U1232 (N_1232,N_855,N_585);
nor U1233 (N_1233,N_578,N_662);
nor U1234 (N_1234,N_956,N_831);
nand U1235 (N_1235,N_528,N_618);
nor U1236 (N_1236,N_567,N_916);
nor U1237 (N_1237,N_998,N_845);
or U1238 (N_1238,N_647,N_506);
nor U1239 (N_1239,N_759,N_819);
and U1240 (N_1240,N_532,N_680);
and U1241 (N_1241,N_524,N_512);
or U1242 (N_1242,N_597,N_663);
or U1243 (N_1243,N_564,N_838);
nor U1244 (N_1244,N_988,N_643);
or U1245 (N_1245,N_902,N_716);
or U1246 (N_1246,N_766,N_545);
nor U1247 (N_1247,N_740,N_625);
nor U1248 (N_1248,N_673,N_676);
or U1249 (N_1249,N_677,N_849);
nor U1250 (N_1250,N_528,N_857);
and U1251 (N_1251,N_937,N_596);
and U1252 (N_1252,N_886,N_587);
nor U1253 (N_1253,N_802,N_830);
nand U1254 (N_1254,N_892,N_725);
or U1255 (N_1255,N_901,N_774);
or U1256 (N_1256,N_746,N_769);
or U1257 (N_1257,N_684,N_537);
nand U1258 (N_1258,N_862,N_599);
nand U1259 (N_1259,N_552,N_933);
nor U1260 (N_1260,N_866,N_717);
nor U1261 (N_1261,N_522,N_828);
or U1262 (N_1262,N_996,N_841);
nand U1263 (N_1263,N_546,N_815);
or U1264 (N_1264,N_674,N_593);
and U1265 (N_1265,N_942,N_921);
nor U1266 (N_1266,N_861,N_739);
and U1267 (N_1267,N_698,N_824);
or U1268 (N_1268,N_683,N_880);
and U1269 (N_1269,N_833,N_826);
or U1270 (N_1270,N_653,N_624);
or U1271 (N_1271,N_799,N_551);
or U1272 (N_1272,N_637,N_560);
xnor U1273 (N_1273,N_681,N_904);
nand U1274 (N_1274,N_771,N_789);
and U1275 (N_1275,N_826,N_893);
and U1276 (N_1276,N_987,N_522);
nor U1277 (N_1277,N_726,N_809);
or U1278 (N_1278,N_615,N_785);
or U1279 (N_1279,N_858,N_949);
and U1280 (N_1280,N_912,N_798);
nand U1281 (N_1281,N_533,N_920);
and U1282 (N_1282,N_912,N_591);
or U1283 (N_1283,N_647,N_841);
and U1284 (N_1284,N_780,N_691);
nand U1285 (N_1285,N_948,N_563);
nor U1286 (N_1286,N_581,N_746);
nor U1287 (N_1287,N_828,N_993);
nand U1288 (N_1288,N_616,N_882);
nand U1289 (N_1289,N_870,N_620);
nand U1290 (N_1290,N_878,N_961);
or U1291 (N_1291,N_766,N_653);
and U1292 (N_1292,N_564,N_881);
or U1293 (N_1293,N_858,N_847);
or U1294 (N_1294,N_930,N_842);
or U1295 (N_1295,N_687,N_554);
nand U1296 (N_1296,N_937,N_985);
xor U1297 (N_1297,N_754,N_543);
or U1298 (N_1298,N_733,N_564);
nor U1299 (N_1299,N_636,N_601);
nand U1300 (N_1300,N_533,N_806);
and U1301 (N_1301,N_745,N_724);
or U1302 (N_1302,N_927,N_896);
nor U1303 (N_1303,N_572,N_923);
nor U1304 (N_1304,N_561,N_536);
nand U1305 (N_1305,N_641,N_573);
nor U1306 (N_1306,N_705,N_515);
nand U1307 (N_1307,N_752,N_788);
nor U1308 (N_1308,N_808,N_600);
nor U1309 (N_1309,N_505,N_974);
or U1310 (N_1310,N_505,N_849);
or U1311 (N_1311,N_741,N_780);
nor U1312 (N_1312,N_908,N_663);
and U1313 (N_1313,N_879,N_881);
nor U1314 (N_1314,N_682,N_646);
nor U1315 (N_1315,N_619,N_764);
nor U1316 (N_1316,N_662,N_910);
and U1317 (N_1317,N_576,N_887);
nand U1318 (N_1318,N_553,N_524);
and U1319 (N_1319,N_590,N_687);
nor U1320 (N_1320,N_947,N_666);
and U1321 (N_1321,N_713,N_928);
nor U1322 (N_1322,N_505,N_501);
and U1323 (N_1323,N_579,N_526);
and U1324 (N_1324,N_783,N_732);
nor U1325 (N_1325,N_515,N_804);
nand U1326 (N_1326,N_680,N_548);
or U1327 (N_1327,N_620,N_570);
and U1328 (N_1328,N_537,N_602);
nand U1329 (N_1329,N_836,N_963);
nor U1330 (N_1330,N_778,N_567);
nor U1331 (N_1331,N_636,N_579);
or U1332 (N_1332,N_909,N_596);
or U1333 (N_1333,N_604,N_688);
nor U1334 (N_1334,N_721,N_886);
nand U1335 (N_1335,N_830,N_533);
nor U1336 (N_1336,N_980,N_847);
and U1337 (N_1337,N_914,N_675);
nor U1338 (N_1338,N_777,N_552);
and U1339 (N_1339,N_782,N_663);
or U1340 (N_1340,N_752,N_877);
xnor U1341 (N_1341,N_966,N_523);
or U1342 (N_1342,N_724,N_883);
xnor U1343 (N_1343,N_920,N_610);
xnor U1344 (N_1344,N_509,N_635);
nor U1345 (N_1345,N_526,N_610);
and U1346 (N_1346,N_774,N_757);
nand U1347 (N_1347,N_987,N_651);
nor U1348 (N_1348,N_521,N_592);
or U1349 (N_1349,N_711,N_991);
xor U1350 (N_1350,N_922,N_737);
nand U1351 (N_1351,N_862,N_683);
and U1352 (N_1352,N_740,N_696);
nand U1353 (N_1353,N_899,N_788);
and U1354 (N_1354,N_634,N_862);
and U1355 (N_1355,N_724,N_654);
or U1356 (N_1356,N_832,N_733);
or U1357 (N_1357,N_841,N_795);
nand U1358 (N_1358,N_673,N_544);
nand U1359 (N_1359,N_978,N_800);
and U1360 (N_1360,N_973,N_696);
nor U1361 (N_1361,N_555,N_958);
nor U1362 (N_1362,N_884,N_862);
and U1363 (N_1363,N_971,N_996);
nand U1364 (N_1364,N_934,N_626);
and U1365 (N_1365,N_797,N_703);
and U1366 (N_1366,N_886,N_888);
nand U1367 (N_1367,N_871,N_672);
nand U1368 (N_1368,N_743,N_700);
and U1369 (N_1369,N_562,N_702);
and U1370 (N_1370,N_862,N_734);
or U1371 (N_1371,N_989,N_919);
nand U1372 (N_1372,N_907,N_503);
nand U1373 (N_1373,N_553,N_562);
xnor U1374 (N_1374,N_726,N_705);
or U1375 (N_1375,N_985,N_938);
nor U1376 (N_1376,N_623,N_931);
or U1377 (N_1377,N_908,N_680);
nand U1378 (N_1378,N_880,N_576);
and U1379 (N_1379,N_648,N_655);
or U1380 (N_1380,N_898,N_738);
nor U1381 (N_1381,N_887,N_531);
or U1382 (N_1382,N_521,N_683);
and U1383 (N_1383,N_915,N_826);
nand U1384 (N_1384,N_571,N_771);
nand U1385 (N_1385,N_691,N_823);
nand U1386 (N_1386,N_533,N_642);
or U1387 (N_1387,N_721,N_967);
nand U1388 (N_1388,N_655,N_703);
and U1389 (N_1389,N_675,N_500);
or U1390 (N_1390,N_548,N_653);
and U1391 (N_1391,N_705,N_609);
or U1392 (N_1392,N_803,N_544);
or U1393 (N_1393,N_585,N_792);
or U1394 (N_1394,N_672,N_702);
and U1395 (N_1395,N_636,N_813);
and U1396 (N_1396,N_601,N_848);
and U1397 (N_1397,N_845,N_728);
nand U1398 (N_1398,N_893,N_957);
nand U1399 (N_1399,N_545,N_514);
nand U1400 (N_1400,N_936,N_813);
nor U1401 (N_1401,N_909,N_766);
and U1402 (N_1402,N_661,N_546);
nand U1403 (N_1403,N_958,N_680);
and U1404 (N_1404,N_727,N_984);
nor U1405 (N_1405,N_879,N_756);
or U1406 (N_1406,N_641,N_971);
nor U1407 (N_1407,N_597,N_600);
nor U1408 (N_1408,N_622,N_946);
and U1409 (N_1409,N_771,N_626);
and U1410 (N_1410,N_568,N_996);
nor U1411 (N_1411,N_803,N_711);
or U1412 (N_1412,N_591,N_555);
or U1413 (N_1413,N_618,N_650);
or U1414 (N_1414,N_901,N_800);
nor U1415 (N_1415,N_619,N_967);
and U1416 (N_1416,N_749,N_872);
nor U1417 (N_1417,N_975,N_819);
or U1418 (N_1418,N_694,N_585);
nand U1419 (N_1419,N_573,N_537);
nor U1420 (N_1420,N_933,N_869);
or U1421 (N_1421,N_975,N_891);
nor U1422 (N_1422,N_561,N_990);
and U1423 (N_1423,N_872,N_797);
nor U1424 (N_1424,N_708,N_833);
and U1425 (N_1425,N_820,N_741);
nor U1426 (N_1426,N_773,N_660);
and U1427 (N_1427,N_611,N_682);
or U1428 (N_1428,N_570,N_665);
or U1429 (N_1429,N_564,N_742);
nor U1430 (N_1430,N_917,N_838);
nand U1431 (N_1431,N_550,N_568);
nand U1432 (N_1432,N_962,N_560);
and U1433 (N_1433,N_983,N_587);
or U1434 (N_1434,N_773,N_570);
nand U1435 (N_1435,N_622,N_559);
nor U1436 (N_1436,N_512,N_843);
and U1437 (N_1437,N_539,N_690);
nand U1438 (N_1438,N_598,N_605);
nor U1439 (N_1439,N_834,N_969);
nand U1440 (N_1440,N_967,N_868);
and U1441 (N_1441,N_797,N_852);
nand U1442 (N_1442,N_512,N_569);
or U1443 (N_1443,N_785,N_706);
or U1444 (N_1444,N_600,N_764);
and U1445 (N_1445,N_853,N_845);
and U1446 (N_1446,N_616,N_511);
nor U1447 (N_1447,N_657,N_634);
or U1448 (N_1448,N_518,N_773);
nor U1449 (N_1449,N_630,N_922);
nor U1450 (N_1450,N_928,N_777);
nor U1451 (N_1451,N_646,N_943);
or U1452 (N_1452,N_613,N_840);
nand U1453 (N_1453,N_724,N_781);
nor U1454 (N_1454,N_892,N_714);
nand U1455 (N_1455,N_751,N_600);
nand U1456 (N_1456,N_868,N_805);
or U1457 (N_1457,N_983,N_723);
nand U1458 (N_1458,N_572,N_550);
or U1459 (N_1459,N_782,N_668);
nor U1460 (N_1460,N_557,N_705);
or U1461 (N_1461,N_507,N_581);
and U1462 (N_1462,N_944,N_612);
nor U1463 (N_1463,N_507,N_743);
nor U1464 (N_1464,N_643,N_716);
nor U1465 (N_1465,N_987,N_873);
or U1466 (N_1466,N_539,N_955);
or U1467 (N_1467,N_690,N_701);
xnor U1468 (N_1468,N_720,N_794);
nor U1469 (N_1469,N_801,N_589);
xnor U1470 (N_1470,N_533,N_843);
or U1471 (N_1471,N_937,N_563);
nor U1472 (N_1472,N_962,N_946);
and U1473 (N_1473,N_737,N_842);
nor U1474 (N_1474,N_957,N_998);
nor U1475 (N_1475,N_571,N_890);
nor U1476 (N_1476,N_855,N_832);
nand U1477 (N_1477,N_778,N_651);
nand U1478 (N_1478,N_699,N_619);
or U1479 (N_1479,N_824,N_545);
nor U1480 (N_1480,N_534,N_718);
or U1481 (N_1481,N_900,N_803);
xnor U1482 (N_1482,N_506,N_815);
and U1483 (N_1483,N_817,N_821);
nand U1484 (N_1484,N_501,N_837);
nand U1485 (N_1485,N_678,N_548);
or U1486 (N_1486,N_894,N_732);
nand U1487 (N_1487,N_874,N_859);
nor U1488 (N_1488,N_904,N_601);
or U1489 (N_1489,N_947,N_561);
nor U1490 (N_1490,N_705,N_684);
nand U1491 (N_1491,N_796,N_508);
nand U1492 (N_1492,N_631,N_811);
nand U1493 (N_1493,N_713,N_865);
or U1494 (N_1494,N_737,N_695);
nand U1495 (N_1495,N_763,N_500);
or U1496 (N_1496,N_663,N_852);
xor U1497 (N_1497,N_716,N_571);
and U1498 (N_1498,N_950,N_944);
nor U1499 (N_1499,N_902,N_621);
nor U1500 (N_1500,N_1326,N_1048);
nand U1501 (N_1501,N_1477,N_1420);
nor U1502 (N_1502,N_1120,N_1408);
or U1503 (N_1503,N_1208,N_1244);
nand U1504 (N_1504,N_1049,N_1128);
xnor U1505 (N_1505,N_1439,N_1034);
nand U1506 (N_1506,N_1228,N_1407);
nand U1507 (N_1507,N_1130,N_1322);
and U1508 (N_1508,N_1022,N_1294);
nor U1509 (N_1509,N_1398,N_1225);
or U1510 (N_1510,N_1395,N_1052);
and U1511 (N_1511,N_1112,N_1235);
nand U1512 (N_1512,N_1449,N_1129);
or U1513 (N_1513,N_1017,N_1219);
or U1514 (N_1514,N_1105,N_1153);
nor U1515 (N_1515,N_1174,N_1324);
or U1516 (N_1516,N_1156,N_1419);
and U1517 (N_1517,N_1142,N_1366);
nand U1518 (N_1518,N_1286,N_1230);
nor U1519 (N_1519,N_1269,N_1304);
nand U1520 (N_1520,N_1152,N_1328);
nand U1521 (N_1521,N_1397,N_1405);
nor U1522 (N_1522,N_1414,N_1250);
nand U1523 (N_1523,N_1470,N_1005);
nor U1524 (N_1524,N_1488,N_1224);
and U1525 (N_1525,N_1370,N_1400);
nor U1526 (N_1526,N_1147,N_1023);
nor U1527 (N_1527,N_1100,N_1499);
nand U1528 (N_1528,N_1284,N_1331);
and U1529 (N_1529,N_1191,N_1494);
nor U1530 (N_1530,N_1479,N_1095);
nor U1531 (N_1531,N_1201,N_1197);
nand U1532 (N_1532,N_1055,N_1200);
or U1533 (N_1533,N_1217,N_1061);
nor U1534 (N_1534,N_1046,N_1468);
nand U1535 (N_1535,N_1181,N_1424);
nand U1536 (N_1536,N_1173,N_1384);
or U1537 (N_1537,N_1213,N_1248);
nor U1538 (N_1538,N_1280,N_1483);
and U1539 (N_1539,N_1246,N_1388);
xnor U1540 (N_1540,N_1204,N_1391);
and U1541 (N_1541,N_1254,N_1498);
and U1542 (N_1542,N_1495,N_1166);
and U1543 (N_1543,N_1444,N_1072);
and U1544 (N_1544,N_1427,N_1068);
and U1545 (N_1545,N_1353,N_1050);
and U1546 (N_1546,N_1148,N_1183);
and U1547 (N_1547,N_1143,N_1441);
or U1548 (N_1548,N_1249,N_1110);
nor U1549 (N_1549,N_1103,N_1385);
and U1550 (N_1550,N_1306,N_1330);
and U1551 (N_1551,N_1350,N_1123);
or U1552 (N_1552,N_1389,N_1303);
and U1553 (N_1553,N_1067,N_1079);
or U1554 (N_1554,N_1188,N_1186);
or U1555 (N_1555,N_1283,N_1401);
and U1556 (N_1556,N_1274,N_1481);
nand U1557 (N_1557,N_1032,N_1360);
or U1558 (N_1558,N_1094,N_1010);
nor U1559 (N_1559,N_1027,N_1321);
nand U1560 (N_1560,N_1109,N_1457);
and U1561 (N_1561,N_1333,N_1221);
or U1562 (N_1562,N_1253,N_1346);
nand U1563 (N_1563,N_1099,N_1466);
nor U1564 (N_1564,N_1450,N_1451);
and U1565 (N_1565,N_1336,N_1258);
nand U1566 (N_1566,N_1090,N_1454);
or U1567 (N_1567,N_1164,N_1111);
nand U1568 (N_1568,N_1361,N_1382);
and U1569 (N_1569,N_1206,N_1452);
nand U1570 (N_1570,N_1476,N_1238);
or U1571 (N_1571,N_1210,N_1141);
and U1572 (N_1572,N_1209,N_1255);
or U1573 (N_1573,N_1308,N_1231);
nor U1574 (N_1574,N_1226,N_1394);
and U1575 (N_1575,N_1363,N_1045);
and U1576 (N_1576,N_1101,N_1014);
and U1577 (N_1577,N_1114,N_1106);
nand U1578 (N_1578,N_1019,N_1012);
nor U1579 (N_1579,N_1376,N_1497);
and U1580 (N_1580,N_1115,N_1198);
or U1581 (N_1581,N_1282,N_1078);
and U1582 (N_1582,N_1410,N_1338);
or U1583 (N_1583,N_1463,N_1030);
and U1584 (N_1584,N_1262,N_1136);
and U1585 (N_1585,N_1205,N_1489);
or U1586 (N_1586,N_1365,N_1337);
or U1587 (N_1587,N_1493,N_1240);
and U1588 (N_1588,N_1301,N_1381);
nor U1589 (N_1589,N_1311,N_1276);
nor U1590 (N_1590,N_1478,N_1092);
and U1591 (N_1591,N_1264,N_1437);
and U1592 (N_1592,N_1172,N_1297);
nor U1593 (N_1593,N_1473,N_1289);
nand U1594 (N_1594,N_1377,N_1039);
and U1595 (N_1595,N_1309,N_1179);
and U1596 (N_1596,N_1369,N_1257);
nand U1597 (N_1597,N_1462,N_1295);
or U1598 (N_1598,N_1480,N_1137);
nor U1599 (N_1599,N_1131,N_1448);
and U1600 (N_1600,N_1227,N_1354);
and U1601 (N_1601,N_1063,N_1455);
and U1602 (N_1602,N_1171,N_1440);
and U1603 (N_1603,N_1356,N_1281);
and U1604 (N_1604,N_1118,N_1373);
or U1605 (N_1605,N_1140,N_1059);
nand U1606 (N_1606,N_1344,N_1310);
and U1607 (N_1607,N_1178,N_1066);
and U1608 (N_1608,N_1232,N_1058);
or U1609 (N_1609,N_1203,N_1189);
or U1610 (N_1610,N_1418,N_1051);
nand U1611 (N_1611,N_1436,N_1266);
nand U1612 (N_1612,N_1475,N_1223);
nor U1613 (N_1613,N_1413,N_1315);
and U1614 (N_1614,N_1412,N_1013);
nor U1615 (N_1615,N_1177,N_1009);
or U1616 (N_1616,N_1229,N_1368);
nand U1617 (N_1617,N_1185,N_1220);
or U1618 (N_1618,N_1342,N_1265);
nor U1619 (N_1619,N_1447,N_1416);
xor U1620 (N_1620,N_1076,N_1456);
and U1621 (N_1621,N_1403,N_1287);
nor U1622 (N_1622,N_1314,N_1077);
or U1623 (N_1623,N_1458,N_1239);
nor U1624 (N_1624,N_1207,N_1187);
nor U1625 (N_1625,N_1340,N_1362);
nand U1626 (N_1626,N_1242,N_1469);
and U1627 (N_1627,N_1319,N_1411);
nand U1628 (N_1628,N_1082,N_1015);
nor U1629 (N_1629,N_1484,N_1162);
and U1630 (N_1630,N_1146,N_1351);
and U1631 (N_1631,N_1459,N_1133);
nand U1632 (N_1632,N_1093,N_1402);
nor U1633 (N_1633,N_1446,N_1091);
nor U1634 (N_1634,N_1263,N_1134);
and U1635 (N_1635,N_1432,N_1102);
xor U1636 (N_1636,N_1272,N_1065);
or U1637 (N_1637,N_1062,N_1318);
or U1638 (N_1638,N_1054,N_1145);
nand U1639 (N_1639,N_1426,N_1000);
nor U1640 (N_1640,N_1279,N_1335);
nor U1641 (N_1641,N_1374,N_1107);
and U1642 (N_1642,N_1071,N_1352);
nor U1643 (N_1643,N_1126,N_1438);
or U1644 (N_1644,N_1371,N_1378);
nor U1645 (N_1645,N_1199,N_1037);
nor U1646 (N_1646,N_1487,N_1445);
nand U1647 (N_1647,N_1087,N_1211);
and U1648 (N_1648,N_1404,N_1267);
nand U1649 (N_1649,N_1021,N_1035);
and U1650 (N_1650,N_1291,N_1430);
nor U1651 (N_1651,N_1379,N_1433);
and U1652 (N_1652,N_1288,N_1222);
and U1653 (N_1653,N_1367,N_1252);
xnor U1654 (N_1654,N_1236,N_1127);
or U1655 (N_1655,N_1421,N_1270);
and U1656 (N_1656,N_1332,N_1464);
and U1657 (N_1657,N_1159,N_1132);
nand U1658 (N_1658,N_1176,N_1165);
and U1659 (N_1659,N_1393,N_1490);
xnor U1660 (N_1660,N_1025,N_1196);
nor U1661 (N_1661,N_1001,N_1486);
nand U1662 (N_1662,N_1327,N_1167);
nand U1663 (N_1663,N_1121,N_1212);
nand U1664 (N_1664,N_1169,N_1259);
and U1665 (N_1665,N_1056,N_1496);
or U1666 (N_1666,N_1043,N_1472);
and U1667 (N_1667,N_1113,N_1074);
nor U1668 (N_1668,N_1435,N_1298);
xnor U1669 (N_1669,N_1268,N_1386);
nand U1670 (N_1670,N_1471,N_1358);
or U1671 (N_1671,N_1299,N_1083);
or U1672 (N_1672,N_1016,N_1396);
and U1673 (N_1673,N_1080,N_1415);
nand U1674 (N_1674,N_1004,N_1161);
nor U1675 (N_1675,N_1234,N_1302);
nand U1676 (N_1676,N_1069,N_1150);
xor U1677 (N_1677,N_1108,N_1215);
nor U1678 (N_1678,N_1359,N_1329);
nand U1679 (N_1679,N_1149,N_1316);
and U1680 (N_1680,N_1104,N_1122);
nor U1681 (N_1681,N_1345,N_1155);
nor U1682 (N_1682,N_1180,N_1474);
xnor U1683 (N_1683,N_1154,N_1348);
and U1684 (N_1684,N_1214,N_1117);
nor U1685 (N_1685,N_1357,N_1278);
and U1686 (N_1686,N_1116,N_1011);
and U1687 (N_1687,N_1399,N_1170);
nand U1688 (N_1688,N_1383,N_1406);
nand U1689 (N_1689,N_1081,N_1125);
nor U1690 (N_1690,N_1390,N_1057);
nor U1691 (N_1691,N_1042,N_1429);
nand U1692 (N_1692,N_1020,N_1380);
and U1693 (N_1693,N_1296,N_1372);
nor U1694 (N_1694,N_1392,N_1138);
nand U1695 (N_1695,N_1460,N_1292);
or U1696 (N_1696,N_1194,N_1467);
nor U1697 (N_1697,N_1168,N_1036);
or U1698 (N_1698,N_1325,N_1024);
and U1699 (N_1699,N_1290,N_1002);
or U1700 (N_1700,N_1422,N_1047);
and U1701 (N_1701,N_1492,N_1085);
nor U1702 (N_1702,N_1285,N_1355);
xnor U1703 (N_1703,N_1453,N_1119);
nor U1704 (N_1704,N_1086,N_1144);
nand U1705 (N_1705,N_1026,N_1060);
and U1706 (N_1706,N_1431,N_1312);
or U1707 (N_1707,N_1247,N_1293);
and U1708 (N_1708,N_1245,N_1184);
nand U1709 (N_1709,N_1097,N_1040);
and U1710 (N_1710,N_1038,N_1442);
and U1711 (N_1711,N_1157,N_1041);
nand U1712 (N_1712,N_1073,N_1028);
nand U1713 (N_1713,N_1409,N_1417);
or U1714 (N_1714,N_1428,N_1260);
or U1715 (N_1715,N_1423,N_1202);
nand U1716 (N_1716,N_1334,N_1300);
and U1717 (N_1717,N_1053,N_1313);
nor U1718 (N_1718,N_1218,N_1465);
nand U1719 (N_1719,N_1271,N_1317);
and U1720 (N_1720,N_1341,N_1064);
nor U1721 (N_1721,N_1485,N_1139);
nand U1722 (N_1722,N_1175,N_1243);
or U1723 (N_1723,N_1261,N_1135);
nor U1724 (N_1724,N_1216,N_1233);
nor U1725 (N_1725,N_1084,N_1160);
nand U1726 (N_1726,N_1029,N_1349);
or U1727 (N_1727,N_1192,N_1008);
and U1728 (N_1728,N_1007,N_1163);
nand U1729 (N_1729,N_1044,N_1098);
and U1730 (N_1730,N_1151,N_1003);
or U1731 (N_1731,N_1070,N_1237);
xnor U1732 (N_1732,N_1251,N_1339);
nor U1733 (N_1733,N_1195,N_1387);
nand U1734 (N_1734,N_1434,N_1277);
or U1735 (N_1735,N_1075,N_1088);
and U1736 (N_1736,N_1425,N_1096);
nand U1737 (N_1737,N_1461,N_1006);
xnor U1738 (N_1738,N_1305,N_1323);
or U1739 (N_1739,N_1482,N_1124);
or U1740 (N_1740,N_1241,N_1275);
xor U1741 (N_1741,N_1443,N_1273);
and U1742 (N_1742,N_1193,N_1375);
or U1743 (N_1743,N_1491,N_1182);
nor U1744 (N_1744,N_1320,N_1158);
or U1745 (N_1745,N_1033,N_1364);
nor U1746 (N_1746,N_1190,N_1256);
or U1747 (N_1747,N_1347,N_1307);
nand U1748 (N_1748,N_1089,N_1031);
and U1749 (N_1749,N_1343,N_1018);
nand U1750 (N_1750,N_1458,N_1376);
and U1751 (N_1751,N_1317,N_1154);
or U1752 (N_1752,N_1379,N_1030);
and U1753 (N_1753,N_1409,N_1167);
nor U1754 (N_1754,N_1045,N_1166);
or U1755 (N_1755,N_1036,N_1368);
nor U1756 (N_1756,N_1472,N_1101);
nand U1757 (N_1757,N_1255,N_1006);
nand U1758 (N_1758,N_1336,N_1296);
or U1759 (N_1759,N_1063,N_1094);
and U1760 (N_1760,N_1109,N_1145);
or U1761 (N_1761,N_1165,N_1436);
or U1762 (N_1762,N_1095,N_1451);
nand U1763 (N_1763,N_1302,N_1444);
and U1764 (N_1764,N_1494,N_1233);
or U1765 (N_1765,N_1008,N_1107);
nor U1766 (N_1766,N_1473,N_1090);
nand U1767 (N_1767,N_1064,N_1387);
nand U1768 (N_1768,N_1280,N_1055);
nand U1769 (N_1769,N_1106,N_1454);
and U1770 (N_1770,N_1196,N_1094);
nand U1771 (N_1771,N_1422,N_1411);
or U1772 (N_1772,N_1321,N_1156);
and U1773 (N_1773,N_1385,N_1311);
nor U1774 (N_1774,N_1076,N_1108);
or U1775 (N_1775,N_1410,N_1361);
nor U1776 (N_1776,N_1192,N_1218);
and U1777 (N_1777,N_1059,N_1064);
nand U1778 (N_1778,N_1130,N_1470);
and U1779 (N_1779,N_1202,N_1268);
nor U1780 (N_1780,N_1297,N_1259);
and U1781 (N_1781,N_1219,N_1363);
or U1782 (N_1782,N_1061,N_1159);
or U1783 (N_1783,N_1165,N_1172);
and U1784 (N_1784,N_1041,N_1084);
or U1785 (N_1785,N_1498,N_1286);
or U1786 (N_1786,N_1139,N_1114);
and U1787 (N_1787,N_1308,N_1421);
or U1788 (N_1788,N_1052,N_1204);
or U1789 (N_1789,N_1420,N_1006);
or U1790 (N_1790,N_1127,N_1026);
nor U1791 (N_1791,N_1124,N_1329);
or U1792 (N_1792,N_1248,N_1416);
or U1793 (N_1793,N_1304,N_1324);
nand U1794 (N_1794,N_1472,N_1394);
nand U1795 (N_1795,N_1368,N_1086);
nand U1796 (N_1796,N_1176,N_1091);
or U1797 (N_1797,N_1334,N_1012);
and U1798 (N_1798,N_1065,N_1429);
and U1799 (N_1799,N_1009,N_1327);
or U1800 (N_1800,N_1458,N_1346);
nor U1801 (N_1801,N_1089,N_1425);
nor U1802 (N_1802,N_1115,N_1125);
and U1803 (N_1803,N_1391,N_1449);
and U1804 (N_1804,N_1373,N_1365);
or U1805 (N_1805,N_1111,N_1095);
or U1806 (N_1806,N_1445,N_1394);
nand U1807 (N_1807,N_1251,N_1280);
nand U1808 (N_1808,N_1075,N_1031);
or U1809 (N_1809,N_1163,N_1382);
nor U1810 (N_1810,N_1056,N_1488);
nor U1811 (N_1811,N_1151,N_1276);
or U1812 (N_1812,N_1103,N_1359);
nor U1813 (N_1813,N_1235,N_1302);
nor U1814 (N_1814,N_1203,N_1108);
or U1815 (N_1815,N_1130,N_1387);
or U1816 (N_1816,N_1351,N_1115);
or U1817 (N_1817,N_1212,N_1265);
nor U1818 (N_1818,N_1176,N_1253);
and U1819 (N_1819,N_1317,N_1125);
and U1820 (N_1820,N_1251,N_1287);
and U1821 (N_1821,N_1337,N_1410);
xor U1822 (N_1822,N_1277,N_1132);
nand U1823 (N_1823,N_1473,N_1204);
nor U1824 (N_1824,N_1165,N_1423);
or U1825 (N_1825,N_1239,N_1285);
nor U1826 (N_1826,N_1453,N_1228);
and U1827 (N_1827,N_1077,N_1092);
nor U1828 (N_1828,N_1199,N_1489);
nor U1829 (N_1829,N_1497,N_1121);
nand U1830 (N_1830,N_1329,N_1114);
or U1831 (N_1831,N_1172,N_1175);
nor U1832 (N_1832,N_1452,N_1163);
nand U1833 (N_1833,N_1019,N_1116);
nand U1834 (N_1834,N_1439,N_1279);
nor U1835 (N_1835,N_1162,N_1115);
and U1836 (N_1836,N_1039,N_1213);
or U1837 (N_1837,N_1001,N_1367);
and U1838 (N_1838,N_1329,N_1158);
nor U1839 (N_1839,N_1083,N_1002);
nand U1840 (N_1840,N_1259,N_1491);
nor U1841 (N_1841,N_1422,N_1469);
or U1842 (N_1842,N_1320,N_1366);
and U1843 (N_1843,N_1363,N_1116);
nand U1844 (N_1844,N_1243,N_1236);
or U1845 (N_1845,N_1473,N_1497);
nand U1846 (N_1846,N_1499,N_1232);
or U1847 (N_1847,N_1366,N_1288);
nand U1848 (N_1848,N_1283,N_1299);
or U1849 (N_1849,N_1262,N_1061);
and U1850 (N_1850,N_1233,N_1040);
or U1851 (N_1851,N_1421,N_1094);
nand U1852 (N_1852,N_1258,N_1073);
or U1853 (N_1853,N_1131,N_1389);
and U1854 (N_1854,N_1455,N_1296);
nand U1855 (N_1855,N_1357,N_1016);
nand U1856 (N_1856,N_1295,N_1179);
nor U1857 (N_1857,N_1314,N_1248);
or U1858 (N_1858,N_1289,N_1299);
nand U1859 (N_1859,N_1117,N_1095);
nand U1860 (N_1860,N_1349,N_1423);
or U1861 (N_1861,N_1011,N_1136);
and U1862 (N_1862,N_1070,N_1076);
and U1863 (N_1863,N_1226,N_1409);
or U1864 (N_1864,N_1318,N_1228);
xnor U1865 (N_1865,N_1198,N_1325);
and U1866 (N_1866,N_1142,N_1122);
xnor U1867 (N_1867,N_1119,N_1237);
or U1868 (N_1868,N_1289,N_1195);
nor U1869 (N_1869,N_1484,N_1275);
and U1870 (N_1870,N_1386,N_1049);
and U1871 (N_1871,N_1147,N_1315);
nor U1872 (N_1872,N_1310,N_1089);
nand U1873 (N_1873,N_1407,N_1062);
and U1874 (N_1874,N_1447,N_1349);
nand U1875 (N_1875,N_1143,N_1459);
or U1876 (N_1876,N_1243,N_1248);
nand U1877 (N_1877,N_1427,N_1058);
nor U1878 (N_1878,N_1249,N_1011);
or U1879 (N_1879,N_1188,N_1367);
nor U1880 (N_1880,N_1312,N_1474);
and U1881 (N_1881,N_1498,N_1315);
or U1882 (N_1882,N_1458,N_1117);
nor U1883 (N_1883,N_1354,N_1441);
or U1884 (N_1884,N_1110,N_1021);
or U1885 (N_1885,N_1152,N_1119);
or U1886 (N_1886,N_1144,N_1319);
nor U1887 (N_1887,N_1172,N_1214);
and U1888 (N_1888,N_1173,N_1373);
nor U1889 (N_1889,N_1260,N_1237);
nor U1890 (N_1890,N_1004,N_1170);
xnor U1891 (N_1891,N_1212,N_1316);
nor U1892 (N_1892,N_1240,N_1458);
and U1893 (N_1893,N_1220,N_1012);
xor U1894 (N_1894,N_1040,N_1025);
or U1895 (N_1895,N_1174,N_1132);
nor U1896 (N_1896,N_1414,N_1477);
and U1897 (N_1897,N_1461,N_1094);
nand U1898 (N_1898,N_1129,N_1429);
and U1899 (N_1899,N_1226,N_1344);
and U1900 (N_1900,N_1131,N_1096);
nand U1901 (N_1901,N_1294,N_1055);
nand U1902 (N_1902,N_1354,N_1123);
nand U1903 (N_1903,N_1138,N_1437);
nor U1904 (N_1904,N_1041,N_1496);
or U1905 (N_1905,N_1400,N_1374);
and U1906 (N_1906,N_1459,N_1415);
nor U1907 (N_1907,N_1404,N_1279);
xnor U1908 (N_1908,N_1064,N_1294);
or U1909 (N_1909,N_1135,N_1176);
or U1910 (N_1910,N_1370,N_1287);
nand U1911 (N_1911,N_1276,N_1171);
and U1912 (N_1912,N_1308,N_1486);
and U1913 (N_1913,N_1219,N_1251);
nor U1914 (N_1914,N_1113,N_1153);
xor U1915 (N_1915,N_1281,N_1129);
nand U1916 (N_1916,N_1386,N_1355);
or U1917 (N_1917,N_1383,N_1061);
xnor U1918 (N_1918,N_1276,N_1122);
and U1919 (N_1919,N_1480,N_1385);
or U1920 (N_1920,N_1487,N_1397);
nor U1921 (N_1921,N_1490,N_1238);
nor U1922 (N_1922,N_1385,N_1118);
nor U1923 (N_1923,N_1429,N_1056);
and U1924 (N_1924,N_1003,N_1319);
nand U1925 (N_1925,N_1250,N_1445);
and U1926 (N_1926,N_1373,N_1388);
or U1927 (N_1927,N_1151,N_1374);
xnor U1928 (N_1928,N_1007,N_1296);
nand U1929 (N_1929,N_1404,N_1150);
and U1930 (N_1930,N_1143,N_1309);
nand U1931 (N_1931,N_1235,N_1206);
and U1932 (N_1932,N_1110,N_1060);
nor U1933 (N_1933,N_1411,N_1303);
and U1934 (N_1934,N_1083,N_1172);
or U1935 (N_1935,N_1155,N_1354);
or U1936 (N_1936,N_1091,N_1407);
or U1937 (N_1937,N_1495,N_1193);
and U1938 (N_1938,N_1403,N_1234);
and U1939 (N_1939,N_1028,N_1153);
or U1940 (N_1940,N_1256,N_1239);
and U1941 (N_1941,N_1146,N_1063);
nor U1942 (N_1942,N_1482,N_1226);
and U1943 (N_1943,N_1259,N_1248);
or U1944 (N_1944,N_1174,N_1451);
nor U1945 (N_1945,N_1022,N_1296);
nor U1946 (N_1946,N_1244,N_1275);
nor U1947 (N_1947,N_1256,N_1062);
nor U1948 (N_1948,N_1227,N_1234);
nand U1949 (N_1949,N_1393,N_1419);
nand U1950 (N_1950,N_1361,N_1453);
nor U1951 (N_1951,N_1226,N_1129);
or U1952 (N_1952,N_1450,N_1309);
and U1953 (N_1953,N_1109,N_1317);
and U1954 (N_1954,N_1143,N_1419);
nor U1955 (N_1955,N_1365,N_1443);
xnor U1956 (N_1956,N_1335,N_1228);
and U1957 (N_1957,N_1013,N_1096);
or U1958 (N_1958,N_1291,N_1210);
nor U1959 (N_1959,N_1424,N_1116);
or U1960 (N_1960,N_1205,N_1043);
and U1961 (N_1961,N_1254,N_1494);
nor U1962 (N_1962,N_1100,N_1025);
and U1963 (N_1963,N_1170,N_1169);
and U1964 (N_1964,N_1401,N_1036);
nand U1965 (N_1965,N_1175,N_1065);
or U1966 (N_1966,N_1149,N_1429);
nor U1967 (N_1967,N_1202,N_1464);
and U1968 (N_1968,N_1306,N_1217);
nor U1969 (N_1969,N_1397,N_1017);
and U1970 (N_1970,N_1183,N_1359);
and U1971 (N_1971,N_1254,N_1193);
and U1972 (N_1972,N_1235,N_1038);
nor U1973 (N_1973,N_1381,N_1187);
and U1974 (N_1974,N_1447,N_1311);
or U1975 (N_1975,N_1200,N_1304);
nand U1976 (N_1976,N_1485,N_1109);
or U1977 (N_1977,N_1234,N_1356);
or U1978 (N_1978,N_1010,N_1282);
nor U1979 (N_1979,N_1089,N_1190);
or U1980 (N_1980,N_1359,N_1044);
nor U1981 (N_1981,N_1393,N_1250);
xor U1982 (N_1982,N_1056,N_1171);
nor U1983 (N_1983,N_1095,N_1134);
and U1984 (N_1984,N_1082,N_1423);
and U1985 (N_1985,N_1006,N_1284);
or U1986 (N_1986,N_1033,N_1205);
nand U1987 (N_1987,N_1121,N_1226);
nand U1988 (N_1988,N_1326,N_1401);
nand U1989 (N_1989,N_1338,N_1376);
and U1990 (N_1990,N_1247,N_1087);
or U1991 (N_1991,N_1441,N_1420);
or U1992 (N_1992,N_1382,N_1431);
nand U1993 (N_1993,N_1073,N_1136);
nor U1994 (N_1994,N_1441,N_1297);
nand U1995 (N_1995,N_1314,N_1305);
nand U1996 (N_1996,N_1200,N_1137);
and U1997 (N_1997,N_1164,N_1231);
or U1998 (N_1998,N_1055,N_1140);
nand U1999 (N_1999,N_1010,N_1078);
xnor U2000 (N_2000,N_1550,N_1748);
or U2001 (N_2001,N_1588,N_1804);
and U2002 (N_2002,N_1916,N_1726);
and U2003 (N_2003,N_1913,N_1824);
and U2004 (N_2004,N_1912,N_1875);
and U2005 (N_2005,N_1898,N_1592);
nor U2006 (N_2006,N_1536,N_1854);
and U2007 (N_2007,N_1858,N_1671);
nand U2008 (N_2008,N_1821,N_1817);
and U2009 (N_2009,N_1539,N_1750);
nand U2010 (N_2010,N_1988,N_1818);
or U2011 (N_2011,N_1838,N_1754);
and U2012 (N_2012,N_1702,N_1587);
and U2013 (N_2013,N_1830,N_1582);
or U2014 (N_2014,N_1560,N_1709);
or U2015 (N_2015,N_1715,N_1865);
or U2016 (N_2016,N_1888,N_1695);
and U2017 (N_2017,N_1815,N_1674);
or U2018 (N_2018,N_1630,N_1848);
and U2019 (N_2019,N_1823,N_1891);
nand U2020 (N_2020,N_1800,N_1935);
nand U2021 (N_2021,N_1842,N_1515);
and U2022 (N_2022,N_1593,N_1977);
nand U2023 (N_2023,N_1921,N_1552);
nand U2024 (N_2024,N_1571,N_1814);
or U2025 (N_2025,N_1775,N_1732);
and U2026 (N_2026,N_1555,N_1970);
or U2027 (N_2027,N_1967,N_1701);
nor U2028 (N_2028,N_1791,N_1670);
and U2029 (N_2029,N_1603,N_1533);
nand U2030 (N_2030,N_1845,N_1855);
nor U2031 (N_2031,N_1739,N_1727);
and U2032 (N_2032,N_1554,N_1751);
and U2033 (N_2033,N_1500,N_1529);
or U2034 (N_2034,N_1857,N_1617);
or U2035 (N_2035,N_1849,N_1867);
nor U2036 (N_2036,N_1793,N_1553);
and U2037 (N_2037,N_1927,N_1955);
nor U2038 (N_2038,N_1876,N_1931);
nand U2039 (N_2039,N_1622,N_1509);
or U2040 (N_2040,N_1565,N_1983);
or U2041 (N_2041,N_1613,N_1526);
nor U2042 (N_2042,N_1658,N_1908);
nor U2043 (N_2043,N_1512,N_1558);
and U2044 (N_2044,N_1743,N_1869);
and U2045 (N_2045,N_1723,N_1822);
and U2046 (N_2046,N_1993,N_1924);
xnor U2047 (N_2047,N_1682,N_1774);
nor U2048 (N_2048,N_1930,N_1741);
and U2049 (N_2049,N_1946,N_1746);
or U2050 (N_2050,N_1675,N_1522);
nand U2051 (N_2051,N_1663,N_1659);
and U2052 (N_2052,N_1717,N_1566);
nand U2053 (N_2053,N_1907,N_1687);
or U2054 (N_2054,N_1646,N_1534);
nand U2055 (N_2055,N_1525,N_1538);
or U2056 (N_2056,N_1863,N_1541);
and U2057 (N_2057,N_1507,N_1847);
nand U2058 (N_2058,N_1795,N_1992);
nand U2059 (N_2059,N_1684,N_1713);
xor U2060 (N_2060,N_1759,N_1980);
and U2061 (N_2061,N_1974,N_1696);
nand U2062 (N_2062,N_1856,N_1742);
nor U2063 (N_2063,N_1962,N_1640);
and U2064 (N_2064,N_1610,N_1615);
nor U2065 (N_2065,N_1664,N_1794);
nand U2066 (N_2066,N_1537,N_1762);
nor U2067 (N_2067,N_1601,N_1986);
and U2068 (N_2068,N_1545,N_1634);
nand U2069 (N_2069,N_1919,N_1595);
xnor U2070 (N_2070,N_1785,N_1703);
nand U2071 (N_2071,N_1721,N_1789);
and U2072 (N_2072,N_1925,N_1656);
nand U2073 (N_2073,N_1599,N_1562);
nor U2074 (N_2074,N_1636,N_1944);
or U2075 (N_2075,N_1811,N_1638);
or U2076 (N_2076,N_1521,N_1535);
and U2077 (N_2077,N_1790,N_1990);
nand U2078 (N_2078,N_1809,N_1846);
and U2079 (N_2079,N_1514,N_1896);
nor U2080 (N_2080,N_1996,N_1761);
and U2081 (N_2081,N_1548,N_1589);
nor U2082 (N_2082,N_1997,N_1707);
nand U2083 (N_2083,N_1673,N_1681);
or U2084 (N_2084,N_1714,N_1685);
nor U2085 (N_2085,N_1755,N_1744);
and U2086 (N_2086,N_1792,N_1984);
or U2087 (N_2087,N_1731,N_1878);
or U2088 (N_2088,N_1561,N_1807);
or U2089 (N_2089,N_1958,N_1711);
and U2090 (N_2090,N_1532,N_1853);
or U2091 (N_2091,N_1773,N_1965);
and U2092 (N_2092,N_1770,N_1692);
nand U2093 (N_2093,N_1914,N_1570);
or U2094 (N_2094,N_1614,N_1704);
or U2095 (N_2095,N_1786,N_1850);
nor U2096 (N_2096,N_1519,N_1963);
nor U2097 (N_2097,N_1712,N_1578);
and U2098 (N_2098,N_1936,N_1691);
or U2099 (N_2099,N_1620,N_1629);
nor U2100 (N_2100,N_1575,N_1852);
and U2101 (N_2101,N_1666,N_1978);
nor U2102 (N_2102,N_1909,N_1543);
and U2103 (N_2103,N_1897,N_1937);
or U2104 (N_2104,N_1540,N_1635);
and U2105 (N_2105,N_1623,N_1995);
nand U2106 (N_2106,N_1667,N_1730);
nand U2107 (N_2107,N_1947,N_1662);
nor U2108 (N_2108,N_1778,N_1987);
nand U2109 (N_2109,N_1841,N_1871);
and U2110 (N_2110,N_1645,N_1951);
or U2111 (N_2111,N_1580,N_1956);
and U2112 (N_2112,N_1698,N_1994);
nor U2113 (N_2113,N_1672,N_1637);
nand U2114 (N_2114,N_1949,N_1763);
and U2115 (N_2115,N_1903,N_1665);
nand U2116 (N_2116,N_1998,N_1669);
nor U2117 (N_2117,N_1864,N_1579);
nand U2118 (N_2118,N_1598,N_1602);
nand U2119 (N_2119,N_1816,N_1834);
or U2120 (N_2120,N_1661,N_1915);
nor U2121 (N_2121,N_1973,N_1805);
and U2122 (N_2122,N_1733,N_1945);
xnor U2123 (N_2123,N_1722,N_1737);
nand U2124 (N_2124,N_1668,N_1942);
nand U2125 (N_2125,N_1939,N_1600);
nor U2126 (N_2126,N_1689,N_1966);
nand U2127 (N_2127,N_1577,N_1954);
nand U2128 (N_2128,N_1819,N_1969);
nand U2129 (N_2129,N_1872,N_1626);
nor U2130 (N_2130,N_1788,N_1950);
or U2131 (N_2131,N_1597,N_1839);
and U2132 (N_2132,N_1829,N_1836);
nor U2133 (N_2133,N_1758,N_1803);
and U2134 (N_2134,N_1928,N_1653);
xor U2135 (N_2135,N_1961,N_1679);
and U2136 (N_2136,N_1720,N_1729);
or U2137 (N_2137,N_1783,N_1837);
nand U2138 (N_2138,N_1879,N_1567);
or U2139 (N_2139,N_1503,N_1933);
nand U2140 (N_2140,N_1641,N_1972);
nor U2141 (N_2141,N_1884,N_1964);
nand U2142 (N_2142,N_1710,N_1825);
nand U2143 (N_2143,N_1893,N_1740);
nand U2144 (N_2144,N_1831,N_1616);
xnor U2145 (N_2145,N_1938,N_1941);
and U2146 (N_2146,N_1745,N_1642);
nor U2147 (N_2147,N_1756,N_1979);
or U2148 (N_2148,N_1920,N_1882);
or U2149 (N_2149,N_1886,N_1652);
and U2150 (N_2150,N_1568,N_1808);
or U2151 (N_2151,N_1621,N_1975);
nand U2152 (N_2152,N_1632,N_1678);
nand U2153 (N_2153,N_1881,N_1594);
nor U2154 (N_2154,N_1502,N_1736);
nor U2155 (N_2155,N_1757,N_1686);
and U2156 (N_2156,N_1870,N_1528);
nand U2157 (N_2157,N_1556,N_1504);
nor U2158 (N_2158,N_1700,N_1880);
nor U2159 (N_2159,N_1802,N_1851);
nor U2160 (N_2160,N_1591,N_1633);
nor U2161 (N_2161,N_1657,N_1835);
nand U2162 (N_2162,N_1799,N_1981);
nand U2163 (N_2163,N_1801,N_1953);
or U2164 (N_2164,N_1564,N_1883);
or U2165 (N_2165,N_1718,N_1612);
nand U2166 (N_2166,N_1840,N_1832);
nor U2167 (N_2167,N_1676,N_1520);
nor U2168 (N_2168,N_1868,N_1531);
nand U2169 (N_2169,N_1677,N_1508);
nand U2170 (N_2170,N_1572,N_1781);
or U2171 (N_2171,N_1971,N_1959);
or U2172 (N_2172,N_1918,N_1530);
and U2173 (N_2173,N_1826,N_1873);
nand U2174 (N_2174,N_1644,N_1890);
and U2175 (N_2175,N_1844,N_1688);
nand U2176 (N_2176,N_1929,N_1728);
nor U2177 (N_2177,N_1861,N_1753);
and U2178 (N_2178,N_1511,N_1866);
nor U2179 (N_2179,N_1833,N_1767);
nor U2180 (N_2180,N_1518,N_1654);
nand U2181 (N_2181,N_1952,N_1899);
nor U2182 (N_2182,N_1843,N_1506);
nor U2183 (N_2183,N_1862,N_1985);
or U2184 (N_2184,N_1697,N_1917);
and U2185 (N_2185,N_1889,N_1606);
nand U2186 (N_2186,N_1586,N_1501);
or U2187 (N_2187,N_1982,N_1900);
nor U2188 (N_2188,N_1694,N_1517);
and U2189 (N_2189,N_1902,N_1583);
or U2190 (N_2190,N_1922,N_1516);
and U2191 (N_2191,N_1557,N_1810);
and U2192 (N_2192,N_1574,N_1563);
nand U2193 (N_2193,N_1650,N_1649);
nand U2194 (N_2194,N_1765,N_1894);
nor U2195 (N_2195,N_1923,N_1991);
and U2196 (N_2196,N_1618,N_1784);
nand U2197 (N_2197,N_1590,N_1596);
nor U2198 (N_2198,N_1895,N_1960);
and U2199 (N_2199,N_1926,N_1934);
nor U2200 (N_2200,N_1619,N_1544);
nor U2201 (N_2201,N_1609,N_1527);
xor U2202 (N_2202,N_1628,N_1859);
nor U2203 (N_2203,N_1604,N_1510);
and U2204 (N_2204,N_1943,N_1989);
or U2205 (N_2205,N_1581,N_1542);
or U2206 (N_2206,N_1513,N_1573);
and U2207 (N_2207,N_1768,N_1608);
or U2208 (N_2208,N_1780,N_1631);
and U2209 (N_2209,N_1749,N_1877);
nor U2210 (N_2210,N_1546,N_1885);
or U2211 (N_2211,N_1576,N_1806);
nor U2212 (N_2212,N_1585,N_1820);
xnor U2213 (N_2213,N_1680,N_1932);
nand U2214 (N_2214,N_1699,N_1906);
nand U2215 (N_2215,N_1976,N_1735);
or U2216 (N_2216,N_1648,N_1505);
nand U2217 (N_2217,N_1705,N_1904);
nand U2218 (N_2218,N_1760,N_1547);
and U2219 (N_2219,N_1611,N_1968);
nor U2220 (N_2220,N_1940,N_1777);
nand U2221 (N_2221,N_1660,N_1797);
and U2222 (N_2222,N_1639,N_1887);
nand U2223 (N_2223,N_1647,N_1828);
or U2224 (N_2224,N_1771,N_1905);
and U2225 (N_2225,N_1892,N_1999);
nand U2226 (N_2226,N_1776,N_1708);
nand U2227 (N_2227,N_1706,N_1738);
xor U2228 (N_2228,N_1812,N_1911);
or U2229 (N_2229,N_1605,N_1798);
and U2230 (N_2230,N_1607,N_1910);
and U2231 (N_2231,N_1655,N_1734);
nand U2232 (N_2232,N_1769,N_1719);
and U2233 (N_2233,N_1559,N_1523);
and U2234 (N_2234,N_1549,N_1782);
nand U2235 (N_2235,N_1651,N_1779);
nand U2236 (N_2236,N_1874,N_1624);
xor U2237 (N_2237,N_1693,N_1901);
nor U2238 (N_2238,N_1948,N_1683);
nor U2239 (N_2239,N_1716,N_1551);
nor U2240 (N_2240,N_1725,N_1766);
nor U2241 (N_2241,N_1813,N_1524);
and U2242 (N_2242,N_1787,N_1772);
or U2243 (N_2243,N_1752,N_1796);
or U2244 (N_2244,N_1747,N_1724);
nand U2245 (N_2245,N_1569,N_1764);
nand U2246 (N_2246,N_1690,N_1625);
nor U2247 (N_2247,N_1827,N_1643);
and U2248 (N_2248,N_1627,N_1860);
nand U2249 (N_2249,N_1584,N_1957);
or U2250 (N_2250,N_1923,N_1999);
nand U2251 (N_2251,N_1984,N_1871);
or U2252 (N_2252,N_1919,N_1987);
nor U2253 (N_2253,N_1894,N_1809);
nor U2254 (N_2254,N_1712,N_1686);
or U2255 (N_2255,N_1945,N_1528);
or U2256 (N_2256,N_1833,N_1811);
nor U2257 (N_2257,N_1852,N_1780);
nor U2258 (N_2258,N_1759,N_1824);
or U2259 (N_2259,N_1561,N_1797);
nand U2260 (N_2260,N_1704,N_1829);
nor U2261 (N_2261,N_1915,N_1716);
or U2262 (N_2262,N_1762,N_1809);
or U2263 (N_2263,N_1794,N_1954);
or U2264 (N_2264,N_1669,N_1813);
nor U2265 (N_2265,N_1956,N_1512);
and U2266 (N_2266,N_1770,N_1788);
and U2267 (N_2267,N_1793,N_1963);
and U2268 (N_2268,N_1534,N_1975);
or U2269 (N_2269,N_1567,N_1963);
nand U2270 (N_2270,N_1717,N_1833);
nor U2271 (N_2271,N_1517,N_1530);
nor U2272 (N_2272,N_1867,N_1558);
nor U2273 (N_2273,N_1891,N_1740);
nand U2274 (N_2274,N_1529,N_1630);
and U2275 (N_2275,N_1702,N_1834);
nor U2276 (N_2276,N_1865,N_1972);
or U2277 (N_2277,N_1872,N_1592);
or U2278 (N_2278,N_1638,N_1904);
nand U2279 (N_2279,N_1982,N_1827);
nor U2280 (N_2280,N_1698,N_1903);
nand U2281 (N_2281,N_1646,N_1554);
nand U2282 (N_2282,N_1645,N_1818);
and U2283 (N_2283,N_1703,N_1909);
nor U2284 (N_2284,N_1820,N_1947);
or U2285 (N_2285,N_1508,N_1759);
or U2286 (N_2286,N_1879,N_1835);
and U2287 (N_2287,N_1510,N_1653);
nand U2288 (N_2288,N_1907,N_1810);
and U2289 (N_2289,N_1755,N_1850);
nor U2290 (N_2290,N_1800,N_1635);
nor U2291 (N_2291,N_1918,N_1913);
or U2292 (N_2292,N_1640,N_1516);
nand U2293 (N_2293,N_1698,N_1957);
nor U2294 (N_2294,N_1711,N_1964);
nand U2295 (N_2295,N_1628,N_1654);
nand U2296 (N_2296,N_1893,N_1824);
or U2297 (N_2297,N_1561,N_1638);
nor U2298 (N_2298,N_1873,N_1784);
xnor U2299 (N_2299,N_1959,N_1803);
nor U2300 (N_2300,N_1595,N_1696);
and U2301 (N_2301,N_1680,N_1997);
nor U2302 (N_2302,N_1624,N_1626);
nand U2303 (N_2303,N_1711,N_1622);
nor U2304 (N_2304,N_1563,N_1690);
nor U2305 (N_2305,N_1578,N_1511);
and U2306 (N_2306,N_1829,N_1792);
or U2307 (N_2307,N_1914,N_1948);
nor U2308 (N_2308,N_1769,N_1505);
or U2309 (N_2309,N_1650,N_1696);
and U2310 (N_2310,N_1814,N_1599);
nor U2311 (N_2311,N_1774,N_1504);
or U2312 (N_2312,N_1998,N_1868);
or U2313 (N_2313,N_1610,N_1971);
nor U2314 (N_2314,N_1719,N_1980);
and U2315 (N_2315,N_1521,N_1641);
and U2316 (N_2316,N_1836,N_1767);
xor U2317 (N_2317,N_1526,N_1906);
nand U2318 (N_2318,N_1877,N_1830);
nor U2319 (N_2319,N_1934,N_1892);
xnor U2320 (N_2320,N_1568,N_1967);
nor U2321 (N_2321,N_1537,N_1957);
nor U2322 (N_2322,N_1905,N_1948);
nand U2323 (N_2323,N_1510,N_1900);
nand U2324 (N_2324,N_1660,N_1847);
and U2325 (N_2325,N_1511,N_1801);
and U2326 (N_2326,N_1971,N_1762);
and U2327 (N_2327,N_1973,N_1759);
and U2328 (N_2328,N_1546,N_1869);
nand U2329 (N_2329,N_1806,N_1658);
and U2330 (N_2330,N_1747,N_1798);
nand U2331 (N_2331,N_1961,N_1757);
nand U2332 (N_2332,N_1592,N_1793);
nand U2333 (N_2333,N_1833,N_1843);
and U2334 (N_2334,N_1834,N_1949);
nand U2335 (N_2335,N_1998,N_1737);
nor U2336 (N_2336,N_1708,N_1843);
and U2337 (N_2337,N_1902,N_1647);
nor U2338 (N_2338,N_1747,N_1931);
or U2339 (N_2339,N_1532,N_1775);
nor U2340 (N_2340,N_1553,N_1958);
nand U2341 (N_2341,N_1737,N_1604);
and U2342 (N_2342,N_1901,N_1510);
nor U2343 (N_2343,N_1512,N_1825);
nand U2344 (N_2344,N_1861,N_1566);
xor U2345 (N_2345,N_1545,N_1883);
or U2346 (N_2346,N_1828,N_1978);
nand U2347 (N_2347,N_1633,N_1609);
nor U2348 (N_2348,N_1968,N_1681);
and U2349 (N_2349,N_1935,N_1862);
nand U2350 (N_2350,N_1681,N_1815);
nor U2351 (N_2351,N_1716,N_1506);
and U2352 (N_2352,N_1863,N_1872);
nor U2353 (N_2353,N_1846,N_1768);
nor U2354 (N_2354,N_1524,N_1522);
or U2355 (N_2355,N_1962,N_1852);
and U2356 (N_2356,N_1601,N_1632);
nor U2357 (N_2357,N_1679,N_1622);
and U2358 (N_2358,N_1948,N_1641);
nand U2359 (N_2359,N_1624,N_1839);
or U2360 (N_2360,N_1807,N_1675);
nor U2361 (N_2361,N_1539,N_1959);
nand U2362 (N_2362,N_1803,N_1642);
nor U2363 (N_2363,N_1636,N_1922);
and U2364 (N_2364,N_1861,N_1846);
nor U2365 (N_2365,N_1932,N_1625);
and U2366 (N_2366,N_1722,N_1795);
nand U2367 (N_2367,N_1503,N_1936);
nand U2368 (N_2368,N_1723,N_1926);
nor U2369 (N_2369,N_1846,N_1711);
and U2370 (N_2370,N_1516,N_1651);
nor U2371 (N_2371,N_1740,N_1647);
or U2372 (N_2372,N_1832,N_1879);
nand U2373 (N_2373,N_1895,N_1530);
nand U2374 (N_2374,N_1653,N_1682);
and U2375 (N_2375,N_1521,N_1616);
or U2376 (N_2376,N_1874,N_1593);
nor U2377 (N_2377,N_1687,N_1683);
or U2378 (N_2378,N_1881,N_1965);
and U2379 (N_2379,N_1659,N_1876);
or U2380 (N_2380,N_1854,N_1527);
and U2381 (N_2381,N_1654,N_1883);
nor U2382 (N_2382,N_1575,N_1728);
nor U2383 (N_2383,N_1780,N_1906);
and U2384 (N_2384,N_1572,N_1561);
and U2385 (N_2385,N_1939,N_1581);
and U2386 (N_2386,N_1661,N_1502);
nor U2387 (N_2387,N_1550,N_1628);
nand U2388 (N_2388,N_1515,N_1756);
and U2389 (N_2389,N_1561,N_1924);
or U2390 (N_2390,N_1830,N_1772);
nor U2391 (N_2391,N_1880,N_1681);
nand U2392 (N_2392,N_1510,N_1789);
nand U2393 (N_2393,N_1866,N_1976);
nand U2394 (N_2394,N_1877,N_1835);
nor U2395 (N_2395,N_1741,N_1791);
and U2396 (N_2396,N_1543,N_1677);
nand U2397 (N_2397,N_1835,N_1548);
and U2398 (N_2398,N_1603,N_1711);
and U2399 (N_2399,N_1541,N_1930);
or U2400 (N_2400,N_1781,N_1689);
or U2401 (N_2401,N_1807,N_1944);
and U2402 (N_2402,N_1827,N_1880);
and U2403 (N_2403,N_1696,N_1655);
and U2404 (N_2404,N_1957,N_1644);
nand U2405 (N_2405,N_1908,N_1874);
and U2406 (N_2406,N_1813,N_1970);
nand U2407 (N_2407,N_1753,N_1948);
or U2408 (N_2408,N_1584,N_1502);
and U2409 (N_2409,N_1861,N_1848);
or U2410 (N_2410,N_1580,N_1660);
and U2411 (N_2411,N_1804,N_1798);
nand U2412 (N_2412,N_1530,N_1672);
nor U2413 (N_2413,N_1654,N_1731);
and U2414 (N_2414,N_1601,N_1554);
or U2415 (N_2415,N_1908,N_1961);
or U2416 (N_2416,N_1523,N_1882);
nor U2417 (N_2417,N_1715,N_1657);
and U2418 (N_2418,N_1680,N_1974);
or U2419 (N_2419,N_1974,N_1678);
and U2420 (N_2420,N_1701,N_1914);
nor U2421 (N_2421,N_1919,N_1712);
nor U2422 (N_2422,N_1950,N_1904);
nor U2423 (N_2423,N_1625,N_1885);
xnor U2424 (N_2424,N_1688,N_1779);
or U2425 (N_2425,N_1521,N_1791);
or U2426 (N_2426,N_1823,N_1868);
nor U2427 (N_2427,N_1934,N_1831);
nor U2428 (N_2428,N_1894,N_1784);
nor U2429 (N_2429,N_1758,N_1642);
or U2430 (N_2430,N_1511,N_1829);
and U2431 (N_2431,N_1746,N_1986);
nand U2432 (N_2432,N_1915,N_1979);
or U2433 (N_2433,N_1857,N_1630);
and U2434 (N_2434,N_1679,N_1796);
and U2435 (N_2435,N_1967,N_1769);
or U2436 (N_2436,N_1947,N_1879);
or U2437 (N_2437,N_1548,N_1982);
nand U2438 (N_2438,N_1608,N_1754);
or U2439 (N_2439,N_1565,N_1643);
and U2440 (N_2440,N_1917,N_1969);
nand U2441 (N_2441,N_1729,N_1736);
nand U2442 (N_2442,N_1701,N_1693);
or U2443 (N_2443,N_1584,N_1549);
nor U2444 (N_2444,N_1528,N_1589);
or U2445 (N_2445,N_1949,N_1783);
nand U2446 (N_2446,N_1703,N_1548);
nand U2447 (N_2447,N_1719,N_1583);
nor U2448 (N_2448,N_1684,N_1580);
nor U2449 (N_2449,N_1994,N_1616);
or U2450 (N_2450,N_1535,N_1930);
nand U2451 (N_2451,N_1998,N_1703);
nor U2452 (N_2452,N_1944,N_1911);
and U2453 (N_2453,N_1628,N_1684);
nor U2454 (N_2454,N_1927,N_1733);
nor U2455 (N_2455,N_1569,N_1513);
and U2456 (N_2456,N_1506,N_1816);
nand U2457 (N_2457,N_1928,N_1778);
nand U2458 (N_2458,N_1712,N_1826);
nand U2459 (N_2459,N_1692,N_1713);
or U2460 (N_2460,N_1600,N_1715);
nand U2461 (N_2461,N_1698,N_1966);
nor U2462 (N_2462,N_1724,N_1886);
and U2463 (N_2463,N_1536,N_1962);
nor U2464 (N_2464,N_1609,N_1648);
nor U2465 (N_2465,N_1571,N_1585);
nor U2466 (N_2466,N_1545,N_1720);
or U2467 (N_2467,N_1805,N_1993);
and U2468 (N_2468,N_1644,N_1886);
nand U2469 (N_2469,N_1556,N_1623);
nor U2470 (N_2470,N_1720,N_1536);
or U2471 (N_2471,N_1766,N_1591);
and U2472 (N_2472,N_1566,N_1786);
nand U2473 (N_2473,N_1590,N_1740);
nor U2474 (N_2474,N_1652,N_1727);
nor U2475 (N_2475,N_1770,N_1544);
nor U2476 (N_2476,N_1887,N_1958);
xor U2477 (N_2477,N_1982,N_1954);
nor U2478 (N_2478,N_1637,N_1841);
nand U2479 (N_2479,N_1662,N_1838);
nand U2480 (N_2480,N_1860,N_1961);
nand U2481 (N_2481,N_1711,N_1751);
nand U2482 (N_2482,N_1804,N_1855);
xor U2483 (N_2483,N_1663,N_1817);
and U2484 (N_2484,N_1850,N_1589);
or U2485 (N_2485,N_1794,N_1638);
and U2486 (N_2486,N_1618,N_1528);
nand U2487 (N_2487,N_1545,N_1659);
or U2488 (N_2488,N_1584,N_1977);
nand U2489 (N_2489,N_1563,N_1667);
and U2490 (N_2490,N_1656,N_1746);
nor U2491 (N_2491,N_1512,N_1564);
or U2492 (N_2492,N_1801,N_1734);
nand U2493 (N_2493,N_1937,N_1955);
nand U2494 (N_2494,N_1784,N_1559);
or U2495 (N_2495,N_1591,N_1559);
and U2496 (N_2496,N_1870,N_1977);
nand U2497 (N_2497,N_1860,N_1630);
or U2498 (N_2498,N_1970,N_1670);
nor U2499 (N_2499,N_1521,N_1890);
nand U2500 (N_2500,N_2323,N_2308);
and U2501 (N_2501,N_2180,N_2147);
nand U2502 (N_2502,N_2316,N_2473);
nor U2503 (N_2503,N_2372,N_2488);
or U2504 (N_2504,N_2411,N_2437);
nand U2505 (N_2505,N_2191,N_2040);
nor U2506 (N_2506,N_2211,N_2283);
nand U2507 (N_2507,N_2182,N_2456);
nand U2508 (N_2508,N_2050,N_2342);
nand U2509 (N_2509,N_2144,N_2078);
nor U2510 (N_2510,N_2338,N_2448);
nand U2511 (N_2511,N_2371,N_2434);
nand U2512 (N_2512,N_2143,N_2068);
nor U2513 (N_2513,N_2482,N_2486);
or U2514 (N_2514,N_2370,N_2295);
and U2515 (N_2515,N_2141,N_2292);
nand U2516 (N_2516,N_2241,N_2045);
nand U2517 (N_2517,N_2362,N_2430);
nand U2518 (N_2518,N_2062,N_2226);
and U2519 (N_2519,N_2337,N_2197);
and U2520 (N_2520,N_2293,N_2190);
nand U2521 (N_2521,N_2163,N_2458);
nor U2522 (N_2522,N_2329,N_2264);
nand U2523 (N_2523,N_2457,N_2112);
nor U2524 (N_2524,N_2319,N_2101);
and U2525 (N_2525,N_2321,N_2250);
nand U2526 (N_2526,N_2441,N_2462);
nor U2527 (N_2527,N_2347,N_2069);
xnor U2528 (N_2528,N_2133,N_2297);
or U2529 (N_2529,N_2010,N_2084);
or U2530 (N_2530,N_2018,N_2234);
nor U2531 (N_2531,N_2122,N_2193);
and U2532 (N_2532,N_2432,N_2464);
nand U2533 (N_2533,N_2254,N_2386);
nor U2534 (N_2534,N_2136,N_2400);
nor U2535 (N_2535,N_2192,N_2352);
nand U2536 (N_2536,N_2108,N_2017);
and U2537 (N_2537,N_2027,N_2425);
nor U2538 (N_2538,N_2281,N_2120);
nand U2539 (N_2539,N_2067,N_2495);
or U2540 (N_2540,N_2460,N_2412);
or U2541 (N_2541,N_2313,N_2009);
nand U2542 (N_2542,N_2110,N_2255);
or U2543 (N_2543,N_2237,N_2198);
xnor U2544 (N_2544,N_2128,N_2228);
or U2545 (N_2545,N_2471,N_2334);
and U2546 (N_2546,N_2146,N_2404);
or U2547 (N_2547,N_2248,N_2238);
nor U2548 (N_2548,N_2200,N_2032);
or U2549 (N_2549,N_2099,N_2220);
or U2550 (N_2550,N_2326,N_2056);
and U2551 (N_2551,N_2157,N_2117);
nor U2552 (N_2552,N_2104,N_2037);
xnor U2553 (N_2553,N_2167,N_2043);
nor U2554 (N_2554,N_2155,N_2349);
and U2555 (N_2555,N_2214,N_2389);
xor U2556 (N_2556,N_2443,N_2127);
nor U2557 (N_2557,N_2291,N_2064);
nor U2558 (N_2558,N_2217,N_2369);
and U2559 (N_2559,N_2420,N_2407);
nand U2560 (N_2560,N_2208,N_2328);
or U2561 (N_2561,N_2435,N_2269);
nand U2562 (N_2562,N_2417,N_2089);
nand U2563 (N_2563,N_2048,N_2149);
nand U2564 (N_2564,N_2097,N_2421);
or U2565 (N_2565,N_2273,N_2001);
or U2566 (N_2566,N_2100,N_2233);
nand U2567 (N_2567,N_2205,N_2353);
nor U2568 (N_2568,N_2481,N_2339);
or U2569 (N_2569,N_2077,N_2090);
nor U2570 (N_2570,N_2185,N_2296);
nor U2571 (N_2571,N_2375,N_2487);
nand U2572 (N_2572,N_2429,N_2232);
and U2573 (N_2573,N_2106,N_2156);
or U2574 (N_2574,N_2409,N_2111);
nand U2575 (N_2575,N_2332,N_2236);
nor U2576 (N_2576,N_2301,N_2403);
and U2577 (N_2577,N_2171,N_2290);
nand U2578 (N_2578,N_2174,N_2072);
or U2579 (N_2579,N_2499,N_2472);
and U2580 (N_2580,N_2051,N_2431);
nand U2581 (N_2581,N_2229,N_2348);
nor U2582 (N_2582,N_2317,N_2414);
nand U2583 (N_2583,N_2224,N_2299);
and U2584 (N_2584,N_2307,N_2222);
nand U2585 (N_2585,N_2275,N_2195);
and U2586 (N_2586,N_2123,N_2350);
or U2587 (N_2587,N_2379,N_2014);
or U2588 (N_2588,N_2408,N_2249);
or U2589 (N_2589,N_2012,N_2245);
or U2590 (N_2590,N_2466,N_2131);
nor U2591 (N_2591,N_2116,N_2145);
or U2592 (N_2592,N_2115,N_2493);
nand U2593 (N_2593,N_2189,N_2331);
nand U2594 (N_2594,N_2169,N_2194);
nand U2595 (N_2595,N_2368,N_2327);
and U2596 (N_2596,N_2474,N_2113);
nor U2597 (N_2597,N_2497,N_2294);
or U2598 (N_2598,N_2324,N_2109);
nand U2599 (N_2599,N_2071,N_2271);
nor U2600 (N_2600,N_2315,N_2138);
and U2601 (N_2601,N_2002,N_2376);
and U2602 (N_2602,N_2346,N_2479);
nand U2603 (N_2603,N_2260,N_2074);
and U2604 (N_2604,N_2207,N_2212);
and U2605 (N_2605,N_2343,N_2385);
nand U2606 (N_2606,N_2240,N_2444);
nand U2607 (N_2607,N_2215,N_2161);
nand U2608 (N_2608,N_2134,N_2419);
nand U2609 (N_2609,N_2102,N_2498);
and U2610 (N_2610,N_2103,N_2150);
and U2611 (N_2611,N_2351,N_2399);
nor U2612 (N_2612,N_2082,N_2085);
or U2613 (N_2613,N_2398,N_2280);
or U2614 (N_2614,N_2478,N_2033);
nor U2615 (N_2615,N_2094,N_2160);
nand U2616 (N_2616,N_2243,N_2231);
nor U2617 (N_2617,N_2451,N_2366);
or U2618 (N_2618,N_2055,N_2046);
and U2619 (N_2619,N_2442,N_2312);
or U2620 (N_2620,N_2202,N_2054);
nand U2621 (N_2621,N_2279,N_2496);
nor U2622 (N_2622,N_2118,N_2476);
xor U2623 (N_2623,N_2251,N_2087);
and U2624 (N_2624,N_2186,N_2314);
or U2625 (N_2625,N_2199,N_2335);
nor U2626 (N_2626,N_2003,N_2176);
nand U2627 (N_2627,N_2107,N_2006);
nand U2628 (N_2628,N_2361,N_2091);
nor U2629 (N_2629,N_2203,N_2341);
nand U2630 (N_2630,N_2393,N_2378);
nor U2631 (N_2631,N_2344,N_2333);
or U2632 (N_2632,N_2066,N_2196);
or U2633 (N_2633,N_2079,N_2021);
or U2634 (N_2634,N_2423,N_2305);
nor U2635 (N_2635,N_2044,N_2396);
and U2636 (N_2636,N_2284,N_2410);
and U2637 (N_2637,N_2465,N_2039);
nand U2638 (N_2638,N_2105,N_2440);
nand U2639 (N_2639,N_2052,N_2153);
nor U2640 (N_2640,N_2042,N_2213);
xor U2641 (N_2641,N_2083,N_2204);
nor U2642 (N_2642,N_2183,N_2494);
nor U2643 (N_2643,N_2247,N_2360);
and U2644 (N_2644,N_2306,N_2322);
and U2645 (N_2645,N_2036,N_2135);
and U2646 (N_2646,N_2459,N_2272);
or U2647 (N_2647,N_2242,N_2380);
or U2648 (N_2648,N_2387,N_2452);
or U2649 (N_2649,N_2450,N_2166);
nor U2650 (N_2650,N_2053,N_2445);
nor U2651 (N_2651,N_2401,N_2354);
or U2652 (N_2652,N_2426,N_2300);
nor U2653 (N_2653,N_2268,N_2274);
and U2654 (N_2654,N_2216,N_2433);
nand U2655 (N_2655,N_2070,N_2173);
or U2656 (N_2656,N_2415,N_2029);
or U2657 (N_2657,N_2162,N_2019);
nor U2658 (N_2658,N_2402,N_2172);
and U2659 (N_2659,N_2165,N_2439);
nor U2660 (N_2660,N_2235,N_2034);
nor U2661 (N_2661,N_2219,N_2015);
and U2662 (N_2662,N_2463,N_2394);
nor U2663 (N_2663,N_2357,N_2179);
or U2664 (N_2664,N_2076,N_2159);
nand U2665 (N_2665,N_2073,N_2388);
nand U2666 (N_2666,N_2261,N_2096);
nor U2667 (N_2667,N_2065,N_2270);
nand U2668 (N_2668,N_2088,N_2383);
nand U2669 (N_2669,N_2230,N_2374);
and U2670 (N_2670,N_2098,N_2221);
and U2671 (N_2671,N_2020,N_2449);
nor U2672 (N_2672,N_2265,N_2125);
xnor U2673 (N_2673,N_2244,N_2038);
nor U2674 (N_2674,N_2391,N_2262);
and U2675 (N_2675,N_2310,N_2278);
nand U2676 (N_2676,N_2151,N_2483);
nand U2677 (N_2677,N_2177,N_2413);
or U2678 (N_2678,N_2225,N_2164);
and U2679 (N_2679,N_2302,N_2137);
nand U2680 (N_2680,N_2469,N_2320);
or U2681 (N_2681,N_2181,N_2158);
nor U2682 (N_2682,N_2489,N_2468);
or U2683 (N_2683,N_2142,N_2059);
nor U2684 (N_2684,N_2168,N_2218);
or U2685 (N_2685,N_2139,N_2390);
or U2686 (N_2686,N_2365,N_2028);
or U2687 (N_2687,N_2259,N_2114);
nor U2688 (N_2688,N_2454,N_2436);
nor U2689 (N_2689,N_2277,N_2359);
and U2690 (N_2690,N_2030,N_2397);
nand U2691 (N_2691,N_2311,N_2446);
nor U2692 (N_2692,N_2209,N_2406);
and U2693 (N_2693,N_2367,N_2022);
nor U2694 (N_2694,N_2057,N_2356);
nor U2695 (N_2695,N_2016,N_2382);
and U2696 (N_2696,N_2184,N_2477);
nand U2697 (N_2697,N_2095,N_2340);
nor U2698 (N_2698,N_2485,N_2336);
and U2699 (N_2699,N_2266,N_2201);
nand U2700 (N_2700,N_2256,N_2484);
and U2701 (N_2701,N_2210,N_2081);
nor U2702 (N_2702,N_2453,N_2049);
or U2703 (N_2703,N_2461,N_2154);
or U2704 (N_2704,N_2148,N_2188);
nor U2705 (N_2705,N_2035,N_2086);
or U2706 (N_2706,N_2304,N_2061);
nor U2707 (N_2707,N_2276,N_2170);
and U2708 (N_2708,N_2467,N_2000);
nor U2709 (N_2709,N_2373,N_2392);
and U2710 (N_2710,N_2206,N_2455);
nor U2711 (N_2711,N_2058,N_2345);
and U2712 (N_2712,N_2246,N_2130);
nand U2713 (N_2713,N_2025,N_2124);
nand U2714 (N_2714,N_2298,N_2416);
xnor U2715 (N_2715,N_2121,N_2258);
nand U2716 (N_2716,N_2011,N_2490);
or U2717 (N_2717,N_2063,N_2405);
and U2718 (N_2718,N_2289,N_2363);
xnor U2719 (N_2719,N_2227,N_2023);
nand U2720 (N_2720,N_2075,N_2492);
and U2721 (N_2721,N_2026,N_2093);
or U2722 (N_2722,N_2438,N_2381);
nand U2723 (N_2723,N_2126,N_2132);
nor U2724 (N_2724,N_2187,N_2152);
or U2725 (N_2725,N_2263,N_2470);
or U2726 (N_2726,N_2282,N_2007);
and U2727 (N_2727,N_2252,N_2330);
xnor U2728 (N_2728,N_2024,N_2325);
nand U2729 (N_2729,N_2080,N_2267);
and U2730 (N_2730,N_2286,N_2239);
or U2731 (N_2731,N_2178,N_2309);
or U2732 (N_2732,N_2418,N_2427);
or U2733 (N_2733,N_2480,N_2475);
nor U2734 (N_2734,N_2119,N_2288);
nand U2735 (N_2735,N_2005,N_2355);
or U2736 (N_2736,N_2257,N_2060);
or U2737 (N_2737,N_2287,N_2422);
nand U2738 (N_2738,N_2358,N_2318);
nor U2739 (N_2739,N_2253,N_2491);
or U2740 (N_2740,N_2013,N_2175);
or U2741 (N_2741,N_2008,N_2428);
and U2742 (N_2742,N_2285,N_2223);
or U2743 (N_2743,N_2303,N_2047);
or U2744 (N_2744,N_2140,N_2031);
and U2745 (N_2745,N_2424,N_2041);
or U2746 (N_2746,N_2004,N_2377);
nand U2747 (N_2747,N_2129,N_2395);
nor U2748 (N_2748,N_2384,N_2092);
nor U2749 (N_2749,N_2364,N_2447);
or U2750 (N_2750,N_2063,N_2485);
and U2751 (N_2751,N_2384,N_2393);
nand U2752 (N_2752,N_2053,N_2222);
or U2753 (N_2753,N_2093,N_2464);
nand U2754 (N_2754,N_2247,N_2371);
or U2755 (N_2755,N_2109,N_2435);
nor U2756 (N_2756,N_2355,N_2155);
and U2757 (N_2757,N_2076,N_2320);
or U2758 (N_2758,N_2415,N_2052);
nand U2759 (N_2759,N_2393,N_2422);
nand U2760 (N_2760,N_2065,N_2196);
or U2761 (N_2761,N_2192,N_2417);
nand U2762 (N_2762,N_2369,N_2200);
nand U2763 (N_2763,N_2434,N_2071);
nand U2764 (N_2764,N_2349,N_2152);
and U2765 (N_2765,N_2382,N_2184);
xor U2766 (N_2766,N_2045,N_2069);
and U2767 (N_2767,N_2264,N_2087);
nor U2768 (N_2768,N_2306,N_2384);
nand U2769 (N_2769,N_2168,N_2345);
nor U2770 (N_2770,N_2031,N_2343);
nor U2771 (N_2771,N_2304,N_2355);
or U2772 (N_2772,N_2435,N_2229);
or U2773 (N_2773,N_2024,N_2148);
or U2774 (N_2774,N_2466,N_2202);
and U2775 (N_2775,N_2103,N_2230);
nand U2776 (N_2776,N_2141,N_2296);
nor U2777 (N_2777,N_2067,N_2444);
nor U2778 (N_2778,N_2113,N_2333);
nor U2779 (N_2779,N_2297,N_2317);
and U2780 (N_2780,N_2354,N_2309);
nand U2781 (N_2781,N_2203,N_2359);
and U2782 (N_2782,N_2136,N_2200);
or U2783 (N_2783,N_2412,N_2021);
and U2784 (N_2784,N_2392,N_2045);
nand U2785 (N_2785,N_2208,N_2291);
nand U2786 (N_2786,N_2278,N_2332);
and U2787 (N_2787,N_2482,N_2234);
and U2788 (N_2788,N_2391,N_2177);
nor U2789 (N_2789,N_2008,N_2235);
or U2790 (N_2790,N_2365,N_2134);
and U2791 (N_2791,N_2480,N_2066);
nand U2792 (N_2792,N_2486,N_2310);
nor U2793 (N_2793,N_2491,N_2337);
or U2794 (N_2794,N_2234,N_2315);
nand U2795 (N_2795,N_2064,N_2112);
and U2796 (N_2796,N_2307,N_2270);
nand U2797 (N_2797,N_2119,N_2280);
nand U2798 (N_2798,N_2488,N_2202);
nand U2799 (N_2799,N_2324,N_2190);
and U2800 (N_2800,N_2203,N_2435);
nor U2801 (N_2801,N_2432,N_2185);
and U2802 (N_2802,N_2044,N_2326);
nor U2803 (N_2803,N_2047,N_2299);
nand U2804 (N_2804,N_2462,N_2080);
nand U2805 (N_2805,N_2178,N_2103);
nand U2806 (N_2806,N_2120,N_2177);
nor U2807 (N_2807,N_2095,N_2259);
and U2808 (N_2808,N_2337,N_2373);
nand U2809 (N_2809,N_2253,N_2365);
nor U2810 (N_2810,N_2191,N_2067);
nand U2811 (N_2811,N_2070,N_2385);
and U2812 (N_2812,N_2320,N_2130);
or U2813 (N_2813,N_2303,N_2446);
or U2814 (N_2814,N_2447,N_2081);
or U2815 (N_2815,N_2034,N_2465);
nor U2816 (N_2816,N_2352,N_2275);
nand U2817 (N_2817,N_2070,N_2129);
or U2818 (N_2818,N_2327,N_2169);
nor U2819 (N_2819,N_2205,N_2167);
nand U2820 (N_2820,N_2160,N_2299);
or U2821 (N_2821,N_2297,N_2267);
nor U2822 (N_2822,N_2302,N_2420);
nor U2823 (N_2823,N_2180,N_2408);
nor U2824 (N_2824,N_2403,N_2011);
and U2825 (N_2825,N_2452,N_2457);
nand U2826 (N_2826,N_2154,N_2075);
xor U2827 (N_2827,N_2187,N_2093);
and U2828 (N_2828,N_2298,N_2109);
or U2829 (N_2829,N_2100,N_2317);
xor U2830 (N_2830,N_2148,N_2047);
nor U2831 (N_2831,N_2027,N_2474);
nor U2832 (N_2832,N_2286,N_2278);
or U2833 (N_2833,N_2203,N_2382);
nand U2834 (N_2834,N_2410,N_2306);
and U2835 (N_2835,N_2497,N_2409);
and U2836 (N_2836,N_2402,N_2105);
or U2837 (N_2837,N_2199,N_2202);
and U2838 (N_2838,N_2478,N_2271);
or U2839 (N_2839,N_2065,N_2098);
or U2840 (N_2840,N_2169,N_2355);
or U2841 (N_2841,N_2150,N_2154);
nor U2842 (N_2842,N_2081,N_2317);
nand U2843 (N_2843,N_2335,N_2331);
nor U2844 (N_2844,N_2242,N_2173);
nand U2845 (N_2845,N_2384,N_2463);
or U2846 (N_2846,N_2232,N_2435);
nor U2847 (N_2847,N_2481,N_2065);
and U2848 (N_2848,N_2289,N_2279);
or U2849 (N_2849,N_2179,N_2257);
nor U2850 (N_2850,N_2476,N_2390);
nor U2851 (N_2851,N_2155,N_2012);
and U2852 (N_2852,N_2224,N_2408);
nor U2853 (N_2853,N_2316,N_2449);
and U2854 (N_2854,N_2256,N_2196);
or U2855 (N_2855,N_2153,N_2169);
and U2856 (N_2856,N_2471,N_2417);
nor U2857 (N_2857,N_2496,N_2378);
nor U2858 (N_2858,N_2302,N_2497);
nor U2859 (N_2859,N_2199,N_2116);
nor U2860 (N_2860,N_2169,N_2317);
nand U2861 (N_2861,N_2495,N_2319);
and U2862 (N_2862,N_2108,N_2275);
nand U2863 (N_2863,N_2006,N_2455);
and U2864 (N_2864,N_2333,N_2403);
and U2865 (N_2865,N_2407,N_2012);
or U2866 (N_2866,N_2101,N_2414);
or U2867 (N_2867,N_2331,N_2317);
nand U2868 (N_2868,N_2265,N_2364);
nor U2869 (N_2869,N_2330,N_2461);
and U2870 (N_2870,N_2155,N_2493);
nand U2871 (N_2871,N_2330,N_2186);
or U2872 (N_2872,N_2243,N_2189);
and U2873 (N_2873,N_2068,N_2076);
nor U2874 (N_2874,N_2480,N_2397);
and U2875 (N_2875,N_2371,N_2477);
nor U2876 (N_2876,N_2292,N_2478);
nor U2877 (N_2877,N_2371,N_2147);
nand U2878 (N_2878,N_2112,N_2453);
or U2879 (N_2879,N_2387,N_2055);
nor U2880 (N_2880,N_2459,N_2153);
and U2881 (N_2881,N_2437,N_2487);
nor U2882 (N_2882,N_2171,N_2387);
nand U2883 (N_2883,N_2074,N_2407);
nor U2884 (N_2884,N_2278,N_2256);
nor U2885 (N_2885,N_2188,N_2238);
and U2886 (N_2886,N_2370,N_2172);
or U2887 (N_2887,N_2378,N_2286);
nor U2888 (N_2888,N_2138,N_2060);
nor U2889 (N_2889,N_2191,N_2340);
and U2890 (N_2890,N_2331,N_2063);
and U2891 (N_2891,N_2498,N_2497);
nand U2892 (N_2892,N_2285,N_2204);
and U2893 (N_2893,N_2248,N_2383);
and U2894 (N_2894,N_2113,N_2139);
nor U2895 (N_2895,N_2344,N_2245);
nor U2896 (N_2896,N_2279,N_2240);
nand U2897 (N_2897,N_2108,N_2460);
nor U2898 (N_2898,N_2236,N_2246);
or U2899 (N_2899,N_2091,N_2206);
nor U2900 (N_2900,N_2080,N_2311);
nand U2901 (N_2901,N_2097,N_2221);
and U2902 (N_2902,N_2265,N_2452);
and U2903 (N_2903,N_2345,N_2412);
nand U2904 (N_2904,N_2373,N_2257);
nand U2905 (N_2905,N_2131,N_2071);
xor U2906 (N_2906,N_2269,N_2054);
and U2907 (N_2907,N_2288,N_2261);
nor U2908 (N_2908,N_2272,N_2384);
nand U2909 (N_2909,N_2057,N_2254);
nand U2910 (N_2910,N_2416,N_2000);
or U2911 (N_2911,N_2201,N_2424);
nand U2912 (N_2912,N_2150,N_2355);
or U2913 (N_2913,N_2138,N_2374);
or U2914 (N_2914,N_2013,N_2112);
nand U2915 (N_2915,N_2288,N_2321);
or U2916 (N_2916,N_2132,N_2393);
or U2917 (N_2917,N_2107,N_2337);
nor U2918 (N_2918,N_2315,N_2113);
nor U2919 (N_2919,N_2356,N_2021);
nor U2920 (N_2920,N_2420,N_2177);
nand U2921 (N_2921,N_2350,N_2301);
xnor U2922 (N_2922,N_2450,N_2373);
or U2923 (N_2923,N_2459,N_2168);
or U2924 (N_2924,N_2328,N_2133);
nand U2925 (N_2925,N_2070,N_2469);
nor U2926 (N_2926,N_2334,N_2042);
nand U2927 (N_2927,N_2220,N_2007);
and U2928 (N_2928,N_2088,N_2299);
nor U2929 (N_2929,N_2413,N_2453);
and U2930 (N_2930,N_2181,N_2018);
nand U2931 (N_2931,N_2012,N_2165);
and U2932 (N_2932,N_2260,N_2085);
nand U2933 (N_2933,N_2110,N_2383);
or U2934 (N_2934,N_2283,N_2213);
nand U2935 (N_2935,N_2263,N_2143);
nand U2936 (N_2936,N_2417,N_2279);
or U2937 (N_2937,N_2494,N_2214);
nor U2938 (N_2938,N_2480,N_2019);
nor U2939 (N_2939,N_2263,N_2306);
and U2940 (N_2940,N_2243,N_2447);
nor U2941 (N_2941,N_2251,N_2144);
nand U2942 (N_2942,N_2332,N_2395);
and U2943 (N_2943,N_2101,N_2318);
or U2944 (N_2944,N_2310,N_2164);
nor U2945 (N_2945,N_2103,N_2325);
nand U2946 (N_2946,N_2260,N_2070);
or U2947 (N_2947,N_2292,N_2325);
and U2948 (N_2948,N_2402,N_2309);
nand U2949 (N_2949,N_2362,N_2013);
nor U2950 (N_2950,N_2402,N_2461);
nand U2951 (N_2951,N_2002,N_2382);
or U2952 (N_2952,N_2390,N_2290);
xnor U2953 (N_2953,N_2188,N_2386);
nand U2954 (N_2954,N_2299,N_2487);
and U2955 (N_2955,N_2252,N_2367);
or U2956 (N_2956,N_2226,N_2033);
nor U2957 (N_2957,N_2245,N_2066);
and U2958 (N_2958,N_2028,N_2462);
or U2959 (N_2959,N_2374,N_2336);
or U2960 (N_2960,N_2452,N_2451);
nor U2961 (N_2961,N_2430,N_2014);
or U2962 (N_2962,N_2237,N_2229);
and U2963 (N_2963,N_2298,N_2026);
nor U2964 (N_2964,N_2394,N_2037);
and U2965 (N_2965,N_2286,N_2437);
nand U2966 (N_2966,N_2064,N_2129);
or U2967 (N_2967,N_2162,N_2222);
nor U2968 (N_2968,N_2352,N_2375);
or U2969 (N_2969,N_2234,N_2054);
nand U2970 (N_2970,N_2145,N_2446);
and U2971 (N_2971,N_2384,N_2235);
nor U2972 (N_2972,N_2408,N_2165);
nand U2973 (N_2973,N_2303,N_2103);
and U2974 (N_2974,N_2204,N_2172);
and U2975 (N_2975,N_2119,N_2283);
xor U2976 (N_2976,N_2172,N_2101);
and U2977 (N_2977,N_2475,N_2046);
and U2978 (N_2978,N_2028,N_2040);
nand U2979 (N_2979,N_2459,N_2070);
nor U2980 (N_2980,N_2147,N_2430);
nor U2981 (N_2981,N_2212,N_2463);
and U2982 (N_2982,N_2269,N_2251);
nor U2983 (N_2983,N_2350,N_2460);
or U2984 (N_2984,N_2024,N_2231);
xnor U2985 (N_2985,N_2256,N_2226);
or U2986 (N_2986,N_2483,N_2189);
nand U2987 (N_2987,N_2000,N_2142);
or U2988 (N_2988,N_2362,N_2131);
xnor U2989 (N_2989,N_2170,N_2137);
nor U2990 (N_2990,N_2017,N_2204);
nor U2991 (N_2991,N_2046,N_2202);
and U2992 (N_2992,N_2420,N_2272);
or U2993 (N_2993,N_2171,N_2340);
and U2994 (N_2994,N_2412,N_2157);
nand U2995 (N_2995,N_2366,N_2410);
or U2996 (N_2996,N_2155,N_2045);
nand U2997 (N_2997,N_2247,N_2396);
or U2998 (N_2998,N_2365,N_2030);
nor U2999 (N_2999,N_2437,N_2140);
or UO_0 (O_0,N_2663,N_2878);
or UO_1 (O_1,N_2879,N_2899);
xor UO_2 (O_2,N_2645,N_2537);
and UO_3 (O_3,N_2893,N_2575);
or UO_4 (O_4,N_2728,N_2802);
and UO_5 (O_5,N_2542,N_2896);
or UO_6 (O_6,N_2701,N_2884);
or UO_7 (O_7,N_2853,N_2628);
nor UO_8 (O_8,N_2909,N_2558);
xor UO_9 (O_9,N_2722,N_2664);
and UO_10 (O_10,N_2656,N_2507);
and UO_11 (O_11,N_2610,N_2887);
or UO_12 (O_12,N_2990,N_2522);
or UO_13 (O_13,N_2807,N_2587);
and UO_14 (O_14,N_2746,N_2959);
or UO_15 (O_15,N_2509,N_2543);
and UO_16 (O_16,N_2987,N_2799);
or UO_17 (O_17,N_2864,N_2854);
or UO_18 (O_18,N_2717,N_2801);
and UO_19 (O_19,N_2639,N_2911);
or UO_20 (O_20,N_2725,N_2501);
nand UO_21 (O_21,N_2905,N_2806);
or UO_22 (O_22,N_2737,N_2697);
and UO_23 (O_23,N_2805,N_2674);
nand UO_24 (O_24,N_2615,N_2828);
nand UO_25 (O_25,N_2997,N_2953);
nor UO_26 (O_26,N_2655,N_2825);
and UO_27 (O_27,N_2880,N_2779);
and UO_28 (O_28,N_2980,N_2745);
or UO_29 (O_29,N_2820,N_2998);
nand UO_30 (O_30,N_2970,N_2604);
nand UO_31 (O_31,N_2772,N_2557);
nor UO_32 (O_32,N_2597,N_2553);
or UO_33 (O_33,N_2931,N_2920);
nand UO_34 (O_34,N_2892,N_2868);
nor UO_35 (O_35,N_2752,N_2741);
and UO_36 (O_36,N_2598,N_2818);
and UO_37 (O_37,N_2533,N_2592);
or UO_38 (O_38,N_2515,N_2739);
or UO_39 (O_39,N_2771,N_2836);
xor UO_40 (O_40,N_2510,N_2840);
nand UO_41 (O_41,N_2785,N_2793);
and UO_42 (O_42,N_2653,N_2706);
nand UO_43 (O_43,N_2577,N_2894);
nor UO_44 (O_44,N_2709,N_2886);
and UO_45 (O_45,N_2762,N_2735);
nand UO_46 (O_46,N_2889,N_2885);
or UO_47 (O_47,N_2937,N_2742);
nand UO_48 (O_48,N_2776,N_2675);
or UO_49 (O_49,N_2829,N_2813);
or UO_50 (O_50,N_2559,N_2842);
nand UO_51 (O_51,N_2684,N_2971);
nor UO_52 (O_52,N_2789,N_2625);
and UO_53 (O_53,N_2599,N_2984);
or UO_54 (O_54,N_2595,N_2526);
or UO_55 (O_55,N_2750,N_2834);
or UO_56 (O_56,N_2614,N_2872);
nor UO_57 (O_57,N_2979,N_2993);
nand UO_58 (O_58,N_2651,N_2594);
or UO_59 (O_59,N_2946,N_2900);
nor UO_60 (O_60,N_2540,N_2535);
or UO_61 (O_61,N_2600,N_2570);
or UO_62 (O_62,N_2647,N_2564);
or UO_63 (O_63,N_2902,N_2539);
nor UO_64 (O_64,N_2965,N_2677);
or UO_65 (O_65,N_2988,N_2778);
nand UO_66 (O_66,N_2692,N_2826);
nand UO_67 (O_67,N_2780,N_2856);
nand UO_68 (O_68,N_2924,N_2898);
nand UO_69 (O_69,N_2744,N_2619);
nor UO_70 (O_70,N_2954,N_2612);
xor UO_71 (O_71,N_2652,N_2985);
and UO_72 (O_72,N_2643,N_2769);
nand UO_73 (O_73,N_2811,N_2624);
and UO_74 (O_74,N_2586,N_2566);
or UO_75 (O_75,N_2848,N_2732);
nand UO_76 (O_76,N_2506,N_2877);
nor UO_77 (O_77,N_2957,N_2883);
or UO_78 (O_78,N_2667,N_2605);
or UO_79 (O_79,N_2622,N_2904);
nor UO_80 (O_80,N_2636,N_2936);
and UO_81 (O_81,N_2631,N_2733);
or UO_82 (O_82,N_2723,N_2753);
or UO_83 (O_83,N_2994,N_2627);
or UO_84 (O_84,N_2915,N_2565);
nor UO_85 (O_85,N_2541,N_2916);
nor UO_86 (O_86,N_2602,N_2873);
nor UO_87 (O_87,N_2693,N_2958);
nand UO_88 (O_88,N_2797,N_2654);
and UO_89 (O_89,N_2830,N_2603);
nor UO_90 (O_90,N_2973,N_2504);
and UO_91 (O_91,N_2591,N_2907);
nor UO_92 (O_92,N_2804,N_2975);
nand UO_93 (O_93,N_2640,N_2669);
nor UO_94 (O_94,N_2500,N_2531);
nor UO_95 (O_95,N_2527,N_2869);
and UO_96 (O_96,N_2682,N_2579);
nand UO_97 (O_97,N_2688,N_2794);
and UO_98 (O_98,N_2863,N_2650);
nor UO_99 (O_99,N_2860,N_2730);
and UO_100 (O_100,N_2574,N_2562);
and UO_101 (O_101,N_2731,N_2502);
nor UO_102 (O_102,N_2724,N_2681);
xor UO_103 (O_103,N_2657,N_2641);
or UO_104 (O_104,N_2713,N_2666);
xor UO_105 (O_105,N_2928,N_2837);
nor UO_106 (O_106,N_2908,N_2788);
and UO_107 (O_107,N_2982,N_2956);
nor UO_108 (O_108,N_2630,N_2934);
and UO_109 (O_109,N_2646,N_2581);
nand UO_110 (O_110,N_2548,N_2758);
or UO_111 (O_111,N_2803,N_2607);
nand UO_112 (O_112,N_2665,N_2648);
nor UO_113 (O_113,N_2919,N_2938);
and UO_114 (O_114,N_2671,N_2759);
nand UO_115 (O_115,N_2765,N_2748);
or UO_116 (O_116,N_2791,N_2949);
or UO_117 (O_117,N_2638,N_2783);
and UO_118 (O_118,N_2544,N_2749);
xor UO_119 (O_119,N_2552,N_2699);
nand UO_120 (O_120,N_2968,N_2616);
nand UO_121 (O_121,N_2512,N_2576);
or UO_122 (O_122,N_2679,N_2550);
nand UO_123 (O_123,N_2734,N_2876);
nor UO_124 (O_124,N_2792,N_2707);
and UO_125 (O_125,N_2991,N_2538);
nand UO_126 (O_126,N_2635,N_2511);
or UO_127 (O_127,N_2881,N_2903);
nand UO_128 (O_128,N_2963,N_2514);
nor UO_129 (O_129,N_2747,N_2768);
nor UO_130 (O_130,N_2964,N_2572);
nor UO_131 (O_131,N_2534,N_2824);
or UO_132 (O_132,N_2634,N_2882);
or UO_133 (O_133,N_2672,N_2606);
and UO_134 (O_134,N_2906,N_2716);
nor UO_135 (O_135,N_2687,N_2668);
or UO_136 (O_136,N_2888,N_2922);
or UO_137 (O_137,N_2782,N_2966);
nor UO_138 (O_138,N_2832,N_2609);
or UO_139 (O_139,N_2571,N_2659);
and UO_140 (O_140,N_2798,N_2658);
or UO_141 (O_141,N_2796,N_2948);
or UO_142 (O_142,N_2582,N_2720);
or UO_143 (O_143,N_2901,N_2851);
and UO_144 (O_144,N_2821,N_2773);
and UO_145 (O_145,N_2913,N_2855);
nand UO_146 (O_146,N_2815,N_2555);
nand UO_147 (O_147,N_2736,N_2685);
or UO_148 (O_148,N_2917,N_2683);
nor UO_149 (O_149,N_2583,N_2866);
and UO_150 (O_150,N_2503,N_2947);
and UO_151 (O_151,N_2580,N_2867);
xnor UO_152 (O_152,N_2755,N_2764);
or UO_153 (O_153,N_2775,N_2740);
or UO_154 (O_154,N_2839,N_2695);
and UO_155 (O_155,N_2961,N_2766);
nand UO_156 (O_156,N_2623,N_2859);
nor UO_157 (O_157,N_2976,N_2554);
or UO_158 (O_158,N_2810,N_2560);
or UO_159 (O_159,N_2967,N_2865);
nor UO_160 (O_160,N_2974,N_2626);
nor UO_161 (O_161,N_2556,N_2814);
or UO_162 (O_162,N_2897,N_2932);
nor UO_163 (O_163,N_2589,N_2516);
and UO_164 (O_164,N_2563,N_2549);
or UO_165 (O_165,N_2875,N_2593);
nor UO_166 (O_166,N_2520,N_2649);
or UO_167 (O_167,N_2686,N_2874);
and UO_168 (O_168,N_2505,N_2710);
nor UO_169 (O_169,N_2618,N_2945);
nor UO_170 (O_170,N_2996,N_2862);
or UO_171 (O_171,N_2529,N_2847);
or UO_172 (O_172,N_2781,N_2841);
nor UO_173 (O_173,N_2524,N_2700);
or UO_174 (O_174,N_2962,N_2871);
or UO_175 (O_175,N_2738,N_2711);
and UO_176 (O_176,N_2952,N_2660);
or UO_177 (O_177,N_2673,N_2532);
nor UO_178 (O_178,N_2568,N_2999);
or UO_179 (O_179,N_2944,N_2989);
and UO_180 (O_180,N_2983,N_2525);
or UO_181 (O_181,N_2918,N_2754);
xnor UO_182 (O_182,N_2923,N_2546);
or UO_183 (O_183,N_2567,N_2819);
and UO_184 (O_184,N_2767,N_2519);
nand UO_185 (O_185,N_2513,N_2912);
nand UO_186 (O_186,N_2827,N_2995);
and UO_187 (O_187,N_2690,N_2551);
and UO_188 (O_188,N_2850,N_2981);
and UO_189 (O_189,N_2705,N_2661);
nor UO_190 (O_190,N_2670,N_2812);
and UO_191 (O_191,N_2578,N_2784);
or UO_192 (O_192,N_2942,N_2584);
and UO_193 (O_193,N_2977,N_2528);
nand UO_194 (O_194,N_2843,N_2910);
or UO_195 (O_195,N_2986,N_2530);
and UO_196 (O_196,N_2757,N_2561);
nand UO_197 (O_197,N_2676,N_2760);
or UO_198 (O_198,N_2992,N_2611);
nand UO_199 (O_199,N_2951,N_2596);
and UO_200 (O_200,N_2644,N_2617);
and UO_201 (O_201,N_2721,N_2521);
nand UO_202 (O_202,N_2930,N_2517);
and UO_203 (O_203,N_2573,N_2632);
nor UO_204 (O_204,N_2817,N_2547);
and UO_205 (O_205,N_2852,N_2523);
nand UO_206 (O_206,N_2914,N_2823);
nor UO_207 (O_207,N_2613,N_2940);
nand UO_208 (O_208,N_2629,N_2508);
nor UO_209 (O_209,N_2774,N_2743);
and UO_210 (O_210,N_2678,N_2972);
nor UO_211 (O_211,N_2763,N_2925);
or UO_212 (O_212,N_2943,N_2590);
nor UO_213 (O_213,N_2858,N_2833);
and UO_214 (O_214,N_2662,N_2691);
nand UO_215 (O_215,N_2545,N_2822);
or UO_216 (O_216,N_2835,N_2777);
and UO_217 (O_217,N_2585,N_2861);
nand UO_218 (O_218,N_2569,N_2726);
nand UO_219 (O_219,N_2857,N_2845);
nand UO_220 (O_220,N_2787,N_2809);
nor UO_221 (O_221,N_2950,N_2846);
or UO_222 (O_222,N_2933,N_2727);
or UO_223 (O_223,N_2808,N_2838);
or UO_224 (O_224,N_2929,N_2790);
nand UO_225 (O_225,N_2895,N_2712);
xor UO_226 (O_226,N_2756,N_2870);
or UO_227 (O_227,N_2770,N_2978);
and UO_228 (O_228,N_2800,N_2890);
and UO_229 (O_229,N_2718,N_2941);
xnor UO_230 (O_230,N_2729,N_2601);
nor UO_231 (O_231,N_2694,N_2751);
nand UO_232 (O_232,N_2891,N_2642);
xnor UO_233 (O_233,N_2708,N_2703);
nand UO_234 (O_234,N_2696,N_2844);
nor UO_235 (O_235,N_2620,N_2588);
nor UO_236 (O_236,N_2926,N_2621);
and UO_237 (O_237,N_2719,N_2702);
nand UO_238 (O_238,N_2969,N_2633);
nor UO_239 (O_239,N_2935,N_2960);
and UO_240 (O_240,N_2927,N_2831);
xnor UO_241 (O_241,N_2786,N_2536);
nor UO_242 (O_242,N_2698,N_2849);
nor UO_243 (O_243,N_2921,N_2704);
and UO_244 (O_244,N_2816,N_2637);
nand UO_245 (O_245,N_2939,N_2608);
and UO_246 (O_246,N_2680,N_2795);
nand UO_247 (O_247,N_2715,N_2955);
nor UO_248 (O_248,N_2689,N_2714);
or UO_249 (O_249,N_2761,N_2518);
and UO_250 (O_250,N_2656,N_2627);
or UO_251 (O_251,N_2732,N_2606);
nor UO_252 (O_252,N_2856,N_2574);
nand UO_253 (O_253,N_2698,N_2539);
or UO_254 (O_254,N_2620,N_2864);
or UO_255 (O_255,N_2704,N_2771);
nor UO_256 (O_256,N_2731,N_2952);
nand UO_257 (O_257,N_2625,N_2529);
and UO_258 (O_258,N_2610,N_2956);
nand UO_259 (O_259,N_2974,N_2625);
nor UO_260 (O_260,N_2852,N_2628);
nor UO_261 (O_261,N_2767,N_2780);
nor UO_262 (O_262,N_2885,N_2643);
or UO_263 (O_263,N_2738,N_2853);
nand UO_264 (O_264,N_2611,N_2675);
nand UO_265 (O_265,N_2506,N_2540);
nand UO_266 (O_266,N_2893,N_2967);
and UO_267 (O_267,N_2726,N_2819);
or UO_268 (O_268,N_2652,N_2603);
or UO_269 (O_269,N_2753,N_2634);
and UO_270 (O_270,N_2992,N_2856);
or UO_271 (O_271,N_2868,N_2544);
xnor UO_272 (O_272,N_2525,N_2965);
and UO_273 (O_273,N_2617,N_2819);
and UO_274 (O_274,N_2807,N_2736);
nor UO_275 (O_275,N_2939,N_2515);
nand UO_276 (O_276,N_2995,N_2703);
nand UO_277 (O_277,N_2660,N_2863);
nand UO_278 (O_278,N_2736,N_2759);
nor UO_279 (O_279,N_2876,N_2768);
xnor UO_280 (O_280,N_2710,N_2766);
and UO_281 (O_281,N_2767,N_2962);
nor UO_282 (O_282,N_2850,N_2804);
and UO_283 (O_283,N_2893,N_2811);
nor UO_284 (O_284,N_2569,N_2832);
nand UO_285 (O_285,N_2737,N_2626);
or UO_286 (O_286,N_2643,N_2851);
nor UO_287 (O_287,N_2858,N_2691);
and UO_288 (O_288,N_2673,N_2965);
and UO_289 (O_289,N_2710,N_2958);
nor UO_290 (O_290,N_2825,N_2719);
nand UO_291 (O_291,N_2696,N_2881);
nor UO_292 (O_292,N_2525,N_2548);
nor UO_293 (O_293,N_2650,N_2534);
nor UO_294 (O_294,N_2787,N_2806);
nor UO_295 (O_295,N_2793,N_2576);
or UO_296 (O_296,N_2941,N_2745);
or UO_297 (O_297,N_2824,N_2772);
nand UO_298 (O_298,N_2995,N_2778);
or UO_299 (O_299,N_2812,N_2826);
nand UO_300 (O_300,N_2755,N_2879);
or UO_301 (O_301,N_2634,N_2626);
or UO_302 (O_302,N_2829,N_2783);
and UO_303 (O_303,N_2770,N_2998);
nor UO_304 (O_304,N_2914,N_2552);
or UO_305 (O_305,N_2762,N_2817);
or UO_306 (O_306,N_2554,N_2694);
nand UO_307 (O_307,N_2979,N_2812);
and UO_308 (O_308,N_2926,N_2668);
nand UO_309 (O_309,N_2955,N_2971);
or UO_310 (O_310,N_2565,N_2824);
and UO_311 (O_311,N_2902,N_2946);
or UO_312 (O_312,N_2686,N_2945);
nor UO_313 (O_313,N_2978,N_2663);
nand UO_314 (O_314,N_2948,N_2817);
and UO_315 (O_315,N_2574,N_2694);
nor UO_316 (O_316,N_2579,N_2741);
and UO_317 (O_317,N_2542,N_2514);
nor UO_318 (O_318,N_2620,N_2836);
nor UO_319 (O_319,N_2594,N_2842);
nand UO_320 (O_320,N_2634,N_2651);
or UO_321 (O_321,N_2628,N_2568);
and UO_322 (O_322,N_2616,N_2644);
nor UO_323 (O_323,N_2634,N_2752);
nand UO_324 (O_324,N_2923,N_2718);
and UO_325 (O_325,N_2984,N_2510);
nor UO_326 (O_326,N_2797,N_2906);
nor UO_327 (O_327,N_2503,N_2663);
or UO_328 (O_328,N_2547,N_2642);
and UO_329 (O_329,N_2770,N_2821);
and UO_330 (O_330,N_2596,N_2552);
and UO_331 (O_331,N_2989,N_2600);
and UO_332 (O_332,N_2711,N_2662);
and UO_333 (O_333,N_2705,N_2919);
or UO_334 (O_334,N_2986,N_2566);
nand UO_335 (O_335,N_2689,N_2867);
nor UO_336 (O_336,N_2592,N_2847);
nor UO_337 (O_337,N_2598,N_2521);
or UO_338 (O_338,N_2966,N_2723);
or UO_339 (O_339,N_2613,N_2858);
nor UO_340 (O_340,N_2599,N_2775);
and UO_341 (O_341,N_2951,N_2843);
and UO_342 (O_342,N_2703,N_2503);
or UO_343 (O_343,N_2602,N_2968);
or UO_344 (O_344,N_2723,N_2961);
nand UO_345 (O_345,N_2511,N_2923);
nand UO_346 (O_346,N_2677,N_2644);
nor UO_347 (O_347,N_2880,N_2556);
and UO_348 (O_348,N_2789,N_2519);
and UO_349 (O_349,N_2966,N_2555);
and UO_350 (O_350,N_2641,N_2627);
xor UO_351 (O_351,N_2839,N_2794);
nor UO_352 (O_352,N_2778,N_2737);
nor UO_353 (O_353,N_2754,N_2636);
nor UO_354 (O_354,N_2557,N_2646);
nor UO_355 (O_355,N_2836,N_2640);
nor UO_356 (O_356,N_2655,N_2716);
nor UO_357 (O_357,N_2700,N_2626);
nor UO_358 (O_358,N_2522,N_2977);
or UO_359 (O_359,N_2754,N_2931);
nand UO_360 (O_360,N_2803,N_2879);
nand UO_361 (O_361,N_2744,N_2834);
and UO_362 (O_362,N_2922,N_2903);
or UO_363 (O_363,N_2778,N_2728);
nand UO_364 (O_364,N_2901,N_2596);
nor UO_365 (O_365,N_2969,N_2793);
nor UO_366 (O_366,N_2685,N_2861);
nand UO_367 (O_367,N_2941,N_2591);
nand UO_368 (O_368,N_2672,N_2900);
nor UO_369 (O_369,N_2954,N_2722);
nor UO_370 (O_370,N_2875,N_2714);
or UO_371 (O_371,N_2668,N_2893);
or UO_372 (O_372,N_2620,N_2962);
and UO_373 (O_373,N_2796,N_2505);
or UO_374 (O_374,N_2892,N_2546);
nand UO_375 (O_375,N_2580,N_2996);
or UO_376 (O_376,N_2547,N_2671);
nand UO_377 (O_377,N_2815,N_2635);
and UO_378 (O_378,N_2968,N_2649);
nand UO_379 (O_379,N_2738,N_2894);
and UO_380 (O_380,N_2507,N_2752);
nand UO_381 (O_381,N_2687,N_2680);
xnor UO_382 (O_382,N_2833,N_2652);
and UO_383 (O_383,N_2630,N_2748);
and UO_384 (O_384,N_2920,N_2903);
nor UO_385 (O_385,N_2535,N_2816);
nor UO_386 (O_386,N_2966,N_2631);
nor UO_387 (O_387,N_2651,N_2636);
nand UO_388 (O_388,N_2680,N_2532);
nor UO_389 (O_389,N_2979,N_2977);
or UO_390 (O_390,N_2941,N_2548);
nand UO_391 (O_391,N_2849,N_2876);
and UO_392 (O_392,N_2643,N_2870);
nor UO_393 (O_393,N_2608,N_2517);
and UO_394 (O_394,N_2712,N_2993);
nand UO_395 (O_395,N_2681,N_2537);
nor UO_396 (O_396,N_2681,N_2605);
nand UO_397 (O_397,N_2953,N_2579);
nor UO_398 (O_398,N_2767,N_2966);
and UO_399 (O_399,N_2667,N_2762);
and UO_400 (O_400,N_2574,N_2773);
or UO_401 (O_401,N_2809,N_2913);
or UO_402 (O_402,N_2598,N_2588);
nor UO_403 (O_403,N_2544,N_2735);
nand UO_404 (O_404,N_2508,N_2634);
or UO_405 (O_405,N_2672,N_2614);
nor UO_406 (O_406,N_2975,N_2561);
and UO_407 (O_407,N_2764,N_2509);
xnor UO_408 (O_408,N_2577,N_2545);
or UO_409 (O_409,N_2855,N_2829);
nand UO_410 (O_410,N_2887,N_2896);
nor UO_411 (O_411,N_2738,N_2709);
and UO_412 (O_412,N_2850,N_2971);
nand UO_413 (O_413,N_2562,N_2816);
or UO_414 (O_414,N_2740,N_2610);
nand UO_415 (O_415,N_2967,N_2914);
and UO_416 (O_416,N_2874,N_2707);
or UO_417 (O_417,N_2790,N_2986);
and UO_418 (O_418,N_2692,N_2815);
nand UO_419 (O_419,N_2993,N_2954);
nor UO_420 (O_420,N_2985,N_2744);
nand UO_421 (O_421,N_2878,N_2897);
nand UO_422 (O_422,N_2709,N_2662);
nand UO_423 (O_423,N_2610,N_2799);
nor UO_424 (O_424,N_2781,N_2565);
and UO_425 (O_425,N_2813,N_2902);
or UO_426 (O_426,N_2876,N_2508);
nor UO_427 (O_427,N_2897,N_2610);
nor UO_428 (O_428,N_2689,N_2799);
and UO_429 (O_429,N_2874,N_2946);
nor UO_430 (O_430,N_2934,N_2788);
nand UO_431 (O_431,N_2746,N_2881);
nor UO_432 (O_432,N_2945,N_2740);
or UO_433 (O_433,N_2551,N_2952);
nor UO_434 (O_434,N_2674,N_2529);
and UO_435 (O_435,N_2560,N_2685);
or UO_436 (O_436,N_2594,N_2644);
and UO_437 (O_437,N_2634,N_2905);
nor UO_438 (O_438,N_2610,N_2827);
nor UO_439 (O_439,N_2900,N_2595);
nand UO_440 (O_440,N_2824,N_2797);
nand UO_441 (O_441,N_2783,N_2742);
or UO_442 (O_442,N_2742,N_2573);
nor UO_443 (O_443,N_2549,N_2777);
nand UO_444 (O_444,N_2634,N_2523);
or UO_445 (O_445,N_2609,N_2815);
nor UO_446 (O_446,N_2649,N_2545);
nand UO_447 (O_447,N_2808,N_2839);
nand UO_448 (O_448,N_2602,N_2880);
nor UO_449 (O_449,N_2775,N_2846);
nand UO_450 (O_450,N_2864,N_2508);
nand UO_451 (O_451,N_2837,N_2940);
nand UO_452 (O_452,N_2980,N_2687);
or UO_453 (O_453,N_2939,N_2695);
nor UO_454 (O_454,N_2644,N_2615);
and UO_455 (O_455,N_2988,N_2605);
xor UO_456 (O_456,N_2661,N_2578);
nor UO_457 (O_457,N_2855,N_2561);
nand UO_458 (O_458,N_2535,N_2605);
or UO_459 (O_459,N_2934,N_2656);
and UO_460 (O_460,N_2930,N_2891);
nand UO_461 (O_461,N_2816,N_2895);
nand UO_462 (O_462,N_2729,N_2884);
nor UO_463 (O_463,N_2752,N_2823);
and UO_464 (O_464,N_2867,N_2895);
or UO_465 (O_465,N_2841,N_2514);
and UO_466 (O_466,N_2967,N_2942);
and UO_467 (O_467,N_2625,N_2682);
nand UO_468 (O_468,N_2639,N_2556);
nor UO_469 (O_469,N_2632,N_2758);
or UO_470 (O_470,N_2908,N_2633);
and UO_471 (O_471,N_2754,N_2829);
nor UO_472 (O_472,N_2663,N_2598);
or UO_473 (O_473,N_2693,N_2741);
nor UO_474 (O_474,N_2532,N_2679);
nor UO_475 (O_475,N_2735,N_2627);
nor UO_476 (O_476,N_2738,N_2649);
nor UO_477 (O_477,N_2880,N_2801);
nand UO_478 (O_478,N_2704,N_2642);
nand UO_479 (O_479,N_2845,N_2990);
and UO_480 (O_480,N_2954,N_2545);
nor UO_481 (O_481,N_2658,N_2926);
and UO_482 (O_482,N_2586,N_2610);
nand UO_483 (O_483,N_2943,N_2723);
or UO_484 (O_484,N_2814,N_2503);
xnor UO_485 (O_485,N_2643,N_2845);
nand UO_486 (O_486,N_2570,N_2959);
nand UO_487 (O_487,N_2800,N_2954);
nand UO_488 (O_488,N_2846,N_2704);
xor UO_489 (O_489,N_2819,N_2834);
and UO_490 (O_490,N_2767,N_2883);
nand UO_491 (O_491,N_2859,N_2592);
and UO_492 (O_492,N_2578,N_2901);
or UO_493 (O_493,N_2810,N_2695);
nand UO_494 (O_494,N_2950,N_2617);
or UO_495 (O_495,N_2839,N_2643);
nand UO_496 (O_496,N_2862,N_2800);
and UO_497 (O_497,N_2733,N_2574);
or UO_498 (O_498,N_2966,N_2863);
nand UO_499 (O_499,N_2930,N_2958);
endmodule