module basic_3000_30000_3500_15_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_2231,In_1075);
nand U1 (N_1,In_1148,In_1197);
nor U2 (N_2,In_2478,In_872);
and U3 (N_3,In_915,In_386);
nor U4 (N_4,In_1632,In_1905);
and U5 (N_5,In_2227,In_1513);
nor U6 (N_6,In_2547,In_1859);
and U7 (N_7,In_1211,In_2955);
or U8 (N_8,In_2774,In_1821);
and U9 (N_9,In_1424,In_2790);
xor U10 (N_10,In_1805,In_296);
and U11 (N_11,In_913,In_1706);
and U12 (N_12,In_470,In_2362);
xnor U13 (N_13,In_1724,In_68);
xnor U14 (N_14,In_221,In_231);
nand U15 (N_15,In_183,In_1602);
nor U16 (N_16,In_1208,In_1471);
nor U17 (N_17,In_2742,In_1642);
nand U18 (N_18,In_2730,In_808);
and U19 (N_19,In_2978,In_891);
and U20 (N_20,In_1231,In_2878);
and U21 (N_21,In_1176,In_2979);
and U22 (N_22,In_996,In_2931);
nand U23 (N_23,In_2308,In_703);
and U24 (N_24,In_869,In_1530);
nand U25 (N_25,In_342,In_2204);
xnor U26 (N_26,In_747,In_275);
nor U27 (N_27,In_790,In_1840);
xor U28 (N_28,In_518,In_2821);
nand U29 (N_29,In_1519,In_1520);
xnor U30 (N_30,In_1326,In_2030);
nor U31 (N_31,In_1159,In_2019);
and U32 (N_32,In_2634,In_2522);
xnor U33 (N_33,In_137,In_76);
nand U34 (N_34,In_1291,In_524);
xor U35 (N_35,In_361,In_1041);
and U36 (N_36,In_2565,In_2825);
or U37 (N_37,In_2364,In_2697);
and U38 (N_38,In_822,In_1031);
xor U39 (N_39,In_2018,In_2628);
or U40 (N_40,In_2964,In_2718);
nand U41 (N_41,In_2161,In_701);
nor U42 (N_42,In_2801,In_1654);
or U43 (N_43,In_477,In_2302);
nor U44 (N_44,In_1172,In_1698);
or U45 (N_45,In_962,In_1068);
nor U46 (N_46,In_1806,In_1767);
xor U47 (N_47,In_1762,In_2732);
nand U48 (N_48,In_911,In_1336);
xor U49 (N_49,In_1274,In_1449);
or U50 (N_50,In_485,In_1299);
xnor U51 (N_51,In_2463,In_947);
xnor U52 (N_52,In_1981,In_1670);
nand U53 (N_53,In_1628,In_2259);
or U54 (N_54,In_1119,In_924);
nand U55 (N_55,In_659,In_2813);
nor U56 (N_56,In_2014,In_2822);
nand U57 (N_57,In_2340,In_1349);
nand U58 (N_58,In_2960,In_2123);
and U59 (N_59,In_1120,In_1546);
nor U60 (N_60,In_2649,In_967);
nor U61 (N_61,In_298,In_2083);
and U62 (N_62,In_2304,In_1467);
or U63 (N_63,In_1376,In_159);
xnor U64 (N_64,In_1759,In_1486);
nand U65 (N_65,In_1776,In_1468);
nor U66 (N_66,In_1946,In_316);
nor U67 (N_67,In_1305,In_1807);
nand U68 (N_68,In_1224,In_305);
nor U69 (N_69,In_1774,In_673);
nor U70 (N_70,In_547,In_1972);
nand U71 (N_71,In_2301,In_2280);
and U72 (N_72,In_2562,In_88);
or U73 (N_73,In_597,In_1963);
and U74 (N_74,In_1690,In_2618);
nor U75 (N_75,In_1430,In_2802);
or U76 (N_76,In_465,In_1741);
or U77 (N_77,In_964,In_1366);
nor U78 (N_78,In_2136,In_1716);
or U79 (N_79,In_1085,In_2596);
xor U80 (N_80,In_2073,In_1769);
nor U81 (N_81,In_2558,In_579);
and U82 (N_82,In_1491,In_1130);
and U83 (N_83,In_2598,In_105);
xor U84 (N_84,In_1027,In_2629);
xnor U85 (N_85,In_1614,In_1631);
xor U86 (N_86,In_1686,In_909);
nand U87 (N_87,In_2533,In_2286);
and U88 (N_88,In_2417,In_658);
nand U89 (N_89,In_991,In_474);
xnor U90 (N_90,In_2450,In_1952);
or U91 (N_91,In_2542,In_1330);
xor U92 (N_92,In_2491,In_819);
nor U93 (N_93,In_543,In_1893);
nand U94 (N_94,In_371,In_2655);
xnor U95 (N_95,In_2705,In_152);
and U96 (N_96,In_2933,In_2470);
or U97 (N_97,In_1846,In_2451);
nor U98 (N_98,In_2111,In_2333);
or U99 (N_99,In_164,In_955);
and U100 (N_100,In_2215,In_520);
xnor U101 (N_101,In_1117,In_2074);
xor U102 (N_102,In_2919,In_635);
nand U103 (N_103,In_161,In_742);
nand U104 (N_104,In_1200,In_2371);
xnor U105 (N_105,In_904,In_2942);
xor U106 (N_106,In_834,In_1506);
nand U107 (N_107,In_1058,In_1728);
xnor U108 (N_108,In_1346,In_2159);
and U109 (N_109,In_2747,In_150);
nor U110 (N_110,In_761,In_1321);
nand U111 (N_111,In_1547,In_421);
xor U112 (N_112,In_2954,In_2999);
and U113 (N_113,In_2795,In_743);
nand U114 (N_114,In_2611,In_2508);
and U115 (N_115,In_1719,In_1787);
nand U116 (N_116,In_2109,In_2342);
or U117 (N_117,In_1599,In_1481);
and U118 (N_118,In_2462,In_2666);
nor U119 (N_119,In_1864,In_2752);
nor U120 (N_120,In_2603,In_2566);
or U121 (N_121,In_740,In_2860);
or U122 (N_122,In_339,In_2741);
xor U123 (N_123,In_2382,In_1517);
and U124 (N_124,In_2521,In_998);
nand U125 (N_125,In_2056,In_1249);
or U126 (N_126,In_1976,In_1934);
nor U127 (N_127,In_2394,In_1509);
xnor U128 (N_128,In_745,In_1906);
xor U129 (N_129,In_2973,In_2997);
and U130 (N_130,In_2791,In_682);
nor U131 (N_131,In_1405,In_2525);
and U132 (N_132,In_2314,In_1936);
and U133 (N_133,In_206,In_1312);
nand U134 (N_134,In_1635,In_1187);
or U135 (N_135,In_1514,In_1442);
nor U136 (N_136,In_782,In_2920);
nor U137 (N_137,In_1466,In_204);
or U138 (N_138,In_975,In_467);
nand U139 (N_139,In_1980,In_1993);
and U140 (N_140,In_450,In_1997);
or U141 (N_141,In_2309,In_2518);
nor U142 (N_142,In_1764,In_1371);
nand U143 (N_143,In_2429,In_1000);
and U144 (N_144,In_1182,In_595);
nand U145 (N_145,In_1017,In_2201);
xnor U146 (N_146,In_1745,In_1758);
and U147 (N_147,In_644,In_758);
or U148 (N_148,In_424,In_180);
nand U149 (N_149,In_444,In_1736);
or U150 (N_150,In_434,In_2276);
and U151 (N_151,In_1350,In_1358);
nor U152 (N_152,In_2710,In_1809);
nor U153 (N_153,In_638,In_1403);
and U154 (N_154,In_1913,In_718);
nor U155 (N_155,In_1340,In_2677);
or U156 (N_156,In_2102,In_1908);
and U157 (N_157,In_1775,In_2953);
xor U158 (N_158,In_880,In_1269);
nand U159 (N_159,In_211,In_1113);
nor U160 (N_160,In_1798,In_2077);
or U161 (N_161,In_1932,In_550);
xor U162 (N_162,In_890,In_2610);
and U163 (N_163,In_1688,In_1036);
or U164 (N_164,In_1239,In_1073);
nand U165 (N_165,In_2187,In_1475);
and U166 (N_166,In_2506,In_480);
and U167 (N_167,In_1488,In_2771);
and U168 (N_168,In_2320,In_2672);
nor U169 (N_169,In_2066,In_2530);
nor U170 (N_170,In_1048,In_1105);
xor U171 (N_171,In_1748,In_1169);
or U172 (N_172,In_959,In_1638);
xnor U173 (N_173,In_1332,In_2938);
or U174 (N_174,In_748,In_2769);
nand U175 (N_175,In_397,In_2380);
nor U176 (N_176,In_1056,In_2344);
xnor U177 (N_177,In_1396,In_2052);
nand U178 (N_178,In_1630,In_538);
nor U179 (N_179,In_28,In_1114);
and U180 (N_180,In_2626,In_1641);
xnor U181 (N_181,In_2166,In_1607);
nand U182 (N_182,In_2914,In_1751);
or U183 (N_183,In_805,In_2651);
and U184 (N_184,In_2962,In_762);
nand U185 (N_185,In_2004,In_922);
or U186 (N_186,In_912,In_288);
or U187 (N_187,In_2067,In_1598);
or U188 (N_188,In_2532,In_2162);
xnor U189 (N_189,In_885,In_1111);
or U190 (N_190,In_1718,In_2516);
and U191 (N_191,In_617,In_233);
and U192 (N_192,In_1785,In_1722);
nor U193 (N_193,In_2581,In_1334);
xnor U194 (N_194,In_496,In_2528);
xnor U195 (N_195,In_2674,In_117);
and U196 (N_196,In_777,In_2922);
nand U197 (N_197,In_753,In_2778);
nor U198 (N_198,In_741,In_446);
and U199 (N_199,In_1969,In_1689);
and U200 (N_200,In_2373,In_2070);
xor U201 (N_201,In_728,In_1498);
nor U202 (N_202,In_1203,In_136);
or U203 (N_203,In_1043,In_2623);
nand U204 (N_204,In_2828,In_879);
xnor U205 (N_205,In_2069,In_561);
xor U206 (N_206,In_1289,In_2434);
nor U207 (N_207,In_592,In_1538);
and U208 (N_208,In_2357,In_267);
xnor U209 (N_209,In_1377,In_727);
nand U210 (N_210,In_795,In_531);
or U211 (N_211,In_1081,In_2662);
xor U212 (N_212,In_2894,In_1589);
or U213 (N_213,In_951,In_1495);
nor U214 (N_214,In_1772,In_189);
nor U215 (N_215,In_2591,In_208);
or U216 (N_216,In_713,In_232);
and U217 (N_217,In_690,In_1600);
or U218 (N_218,In_209,In_1337);
nand U219 (N_219,In_1275,In_2681);
xnor U220 (N_220,In_1702,In_2189);
nor U221 (N_221,In_705,In_395);
nand U222 (N_222,In_2890,In_1878);
nand U223 (N_223,In_2195,In_436);
xnor U224 (N_224,In_1190,In_1282);
nor U225 (N_225,In_2910,In_1069);
nor U226 (N_226,In_2411,In_2269);
and U227 (N_227,In_1398,In_736);
nand U228 (N_228,In_1527,In_2176);
or U229 (N_229,In_2183,In_2337);
and U230 (N_230,In_2891,In_237);
or U231 (N_231,In_750,In_2143);
nor U232 (N_232,In_1064,In_2869);
xnor U233 (N_233,In_2459,In_1605);
xnor U234 (N_234,In_375,In_2445);
xnor U235 (N_235,In_1876,In_430);
or U236 (N_236,In_452,In_1264);
xnor U237 (N_237,In_2082,In_2881);
xnor U238 (N_238,In_2094,In_1884);
nor U239 (N_239,In_337,In_1055);
nand U240 (N_240,In_1916,In_416);
or U241 (N_241,In_400,In_2502);
or U242 (N_242,In_733,In_4);
nor U243 (N_243,In_2225,In_2967);
or U244 (N_244,In_1333,In_1929);
xor U245 (N_245,In_2693,In_799);
nor U246 (N_246,In_2900,In_1287);
and U247 (N_247,In_1300,In_1927);
or U248 (N_248,In_2266,In_103);
and U249 (N_249,In_2453,In_1158);
or U250 (N_250,In_26,In_1339);
nor U251 (N_251,In_2614,In_2602);
xnor U252 (N_252,In_1696,In_1059);
nor U253 (N_253,In_358,In_754);
or U254 (N_254,In_654,In_2652);
and U255 (N_255,In_2492,In_502);
nand U256 (N_256,In_2458,In_1975);
nand U257 (N_257,In_236,In_578);
nand U258 (N_258,In_1714,In_1425);
xor U259 (N_259,In_1889,In_1971);
xor U260 (N_260,In_789,In_958);
xnor U261 (N_261,In_1062,In_954);
and U262 (N_262,In_438,In_2907);
xor U263 (N_263,In_1107,In_141);
or U264 (N_264,In_588,In_573);
nand U265 (N_265,In_148,In_2098);
nor U266 (N_266,In_2807,In_2663);
or U267 (N_267,In_671,In_251);
or U268 (N_268,In_2939,In_2943);
or U269 (N_269,In_1462,In_1994);
or U270 (N_270,In_2986,In_1379);
xnor U271 (N_271,In_2148,In_2966);
and U272 (N_272,In_121,In_2864);
nand U273 (N_273,In_1296,In_2038);
xor U274 (N_274,In_1374,In_1892);
xor U275 (N_275,In_1178,In_2433);
nand U276 (N_276,In_1026,In_2258);
or U277 (N_277,In_1883,In_2993);
xor U278 (N_278,In_1133,In_2969);
and U279 (N_279,In_1438,In_1132);
nand U280 (N_280,In_24,In_2005);
nor U281 (N_281,In_1439,In_2703);
nor U282 (N_282,In_2023,In_262);
or U283 (N_283,In_581,In_85);
nand U284 (N_284,In_1213,In_1021);
nand U285 (N_285,In_1205,In_2589);
or U286 (N_286,In_2559,In_1955);
nor U287 (N_287,In_717,In_1770);
nand U288 (N_288,In_327,In_2386);
or U289 (N_289,In_576,In_1082);
nand U290 (N_290,In_809,In_2326);
and U291 (N_291,In_406,In_2590);
xnor U292 (N_292,In_182,In_2400);
or U293 (N_293,In_1917,In_864);
nand U294 (N_294,In_2410,In_2772);
and U295 (N_295,In_2128,In_2760);
nor U296 (N_296,In_95,In_138);
xor U297 (N_297,In_2902,In_82);
and U298 (N_298,In_490,In_609);
xnor U299 (N_299,In_1005,In_1811);
nand U300 (N_300,In_2250,In_1713);
or U301 (N_301,In_388,In_2378);
or U302 (N_302,In_557,In_1310);
nor U303 (N_303,In_1865,In_440);
and U304 (N_304,In_683,In_1726);
or U305 (N_305,In_279,In_2359);
or U306 (N_306,In_1930,In_2775);
xnor U307 (N_307,In_2288,In_1795);
nand U308 (N_308,In_1356,In_1850);
xnor U309 (N_309,In_2712,In_934);
nor U310 (N_310,In_2488,In_621);
or U311 (N_311,In_1415,In_1368);
xnor U312 (N_312,In_2534,In_422);
and U313 (N_313,In_623,In_651);
xnor U314 (N_314,In_1910,In_2105);
xnor U315 (N_315,In_1126,In_2814);
and U316 (N_316,In_2849,In_1237);
nand U317 (N_317,In_1140,In_1891);
nor U318 (N_318,In_1253,In_888);
nor U319 (N_319,In_2090,In_2156);
nor U320 (N_320,In_1739,In_1035);
nand U321 (N_321,In_1198,In_2743);
and U322 (N_322,In_501,In_2924);
nor U323 (N_323,In_1860,In_2880);
xor U324 (N_324,In_1047,In_2436);
nor U325 (N_325,In_1389,In_2116);
nor U326 (N_326,In_2345,In_771);
xnor U327 (N_327,In_2,In_1730);
nor U328 (N_328,In_1044,In_1435);
and U329 (N_329,In_1623,In_2403);
nand U330 (N_330,In_1037,In_79);
nand U331 (N_331,In_172,In_351);
and U332 (N_332,In_1327,In_2567);
nor U333 (N_333,In_2310,In_2817);
nor U334 (N_334,In_1255,In_437);
nor U335 (N_335,In_712,In_1106);
nand U336 (N_336,In_804,In_2746);
nor U337 (N_337,In_2733,In_1497);
or U338 (N_338,In_1359,In_1450);
or U339 (N_339,In_1460,In_166);
nand U340 (N_340,In_2175,In_2787);
nor U341 (N_341,In_1270,In_1818);
or U342 (N_342,In_636,In_664);
xnor U343 (N_343,In_2545,In_696);
or U344 (N_344,In_930,In_2830);
xnor U345 (N_345,In_47,In_393);
xor U346 (N_346,In_645,In_2640);
nand U347 (N_347,In_1254,In_64);
or U348 (N_348,In_1011,In_1629);
nor U349 (N_349,In_1465,In_2903);
nor U350 (N_350,In_2294,In_1067);
nor U351 (N_351,In_1025,In_2905);
and U352 (N_352,In_2899,In_1813);
xnor U353 (N_353,In_258,In_603);
and U354 (N_354,In_1028,In_514);
nand U355 (N_355,In_404,In_2202);
or U356 (N_356,In_55,In_1341);
nor U357 (N_357,In_2647,In_2923);
and U358 (N_358,In_849,In_2523);
nor U359 (N_359,In_1469,In_1445);
and U360 (N_360,In_887,In_677);
nand U361 (N_361,In_1986,In_179);
xnor U362 (N_362,In_2012,In_17);
nand U363 (N_363,In_2369,In_1476);
nor U364 (N_364,In_1347,In_1455);
and U365 (N_365,In_2812,In_2716);
or U366 (N_366,In_596,In_2694);
nand U367 (N_367,In_86,In_332);
xor U368 (N_368,In_1898,In_2298);
xor U369 (N_369,In_1784,In_2141);
nand U370 (N_370,In_1782,In_1083);
nor U371 (N_371,In_2982,In_2053);
or U372 (N_372,In_2198,In_725);
xor U373 (N_373,In_1861,In_287);
xnor U374 (N_374,In_373,In_162);
and U375 (N_375,In_442,In_60);
and U376 (N_376,In_1093,In_2509);
xor U377 (N_377,In_77,In_1227);
and U378 (N_378,In_230,In_112);
nor U379 (N_379,In_2592,In_12);
xnor U380 (N_380,In_1588,In_2476);
or U381 (N_381,In_2390,In_738);
nand U382 (N_382,In_308,In_1365);
nor U383 (N_383,In_2755,In_787);
and U384 (N_384,In_757,In_2190);
or U385 (N_385,In_1560,In_248);
or U386 (N_386,In_1153,In_2213);
or U387 (N_387,In_1053,In_1317);
nor U388 (N_388,In_261,In_1852);
or U389 (N_389,In_529,In_1240);
or U390 (N_390,In_96,In_1836);
nor U391 (N_391,In_2064,In_986);
and U392 (N_392,In_565,In_300);
xor U393 (N_393,In_2578,In_2781);
xor U394 (N_394,In_2316,In_193);
or U395 (N_395,In_2998,In_933);
and U396 (N_396,In_921,In_2852);
or U397 (N_397,In_234,In_980);
and U398 (N_398,In_91,In_1115);
and U399 (N_399,In_1219,In_1834);
nor U400 (N_400,In_2548,In_1578);
xnor U401 (N_401,In_1680,In_5);
and U402 (N_402,In_2140,In_895);
and U403 (N_403,In_527,In_626);
or U404 (N_404,In_1387,In_66);
nand U405 (N_405,In_336,In_1757);
nand U406 (N_406,In_2306,In_1516);
nand U407 (N_407,In_631,In_2834);
or U408 (N_408,In_87,In_396);
nor U409 (N_409,In_1926,In_1207);
nor U410 (N_410,In_1558,In_1223);
nand U411 (N_411,In_2181,In_1301);
xor U412 (N_412,In_134,In_2046);
and U413 (N_413,In_666,In_290);
nand U414 (N_414,In_871,In_497);
nor U415 (N_415,In_721,In_601);
nand U416 (N_416,In_220,In_1674);
xor U417 (N_417,In_1915,In_1581);
and U418 (N_418,In_2901,In_2670);
nand U419 (N_419,In_460,In_1252);
nand U420 (N_420,In_2132,In_2097);
or U421 (N_421,In_764,In_1692);
xnor U422 (N_422,In_1967,In_14);
nand U423 (N_423,In_1652,In_539);
and U424 (N_424,In_974,In_1597);
nor U425 (N_425,In_2605,In_2636);
nor U426 (N_426,In_94,In_2638);
and U427 (N_427,In_903,In_160);
and U428 (N_428,In_114,In_2058);
and U429 (N_429,In_2059,In_2701);
nor U430 (N_430,In_1961,In_1899);
nor U431 (N_431,In_1562,In_2151);
or U432 (N_432,In_1235,In_2557);
nor U433 (N_433,In_2932,In_285);
nor U434 (N_434,In_2574,In_1406);
and U435 (N_435,In_1508,In_2571);
or U436 (N_436,In_2688,In_2003);
xor U437 (N_437,In_2679,In_2290);
xor U438 (N_438,In_1982,In_1360);
and U439 (N_439,In_1186,In_2729);
or U440 (N_440,In_1956,In_1199);
nand U441 (N_441,In_2351,In_2671);
nor U442 (N_442,In_1742,In_2391);
nand U443 (N_443,In_1477,In_1595);
nand U444 (N_444,In_2720,In_2789);
and U445 (N_445,In_2503,In_1054);
nor U446 (N_446,In_2177,In_2277);
xor U447 (N_447,In_940,In_2644);
xor U448 (N_448,In_672,In_2927);
xor U449 (N_449,In_608,In_1715);
nand U450 (N_450,In_632,In_823);
nand U451 (N_451,In_73,In_1644);
nand U452 (N_452,In_1373,In_1583);
xnor U453 (N_453,In_1886,In_35);
xnor U454 (N_454,In_135,In_449);
nor U455 (N_455,In_2054,In_2112);
xnor U456 (N_456,In_500,In_2009);
nand U457 (N_457,In_532,In_1796);
nand U458 (N_458,In_366,In_1966);
xnor U459 (N_459,In_2117,In_1616);
or U460 (N_460,In_2619,In_2318);
nand U461 (N_461,In_158,In_265);
xor U462 (N_462,In_935,In_939);
xor U463 (N_463,In_276,In_1822);
and U464 (N_464,In_618,In_1364);
and U465 (N_465,In_34,In_1452);
xor U466 (N_466,In_1766,In_674);
or U467 (N_467,In_2051,In_2348);
nor U468 (N_468,In_2253,In_2908);
nor U469 (N_469,In_1734,In_313);
nor U470 (N_470,In_1651,In_1308);
and U471 (N_471,In_284,In_1669);
nor U472 (N_472,In_72,In_606);
or U473 (N_473,In_317,In_2608);
nand U474 (N_474,In_744,In_1401);
xor U475 (N_475,In_1189,In_982);
or U476 (N_476,In_1259,In_30);
or U477 (N_477,In_2803,In_1823);
nand U478 (N_478,In_1019,In_1962);
or U479 (N_479,In_2776,In_1673);
nand U480 (N_480,In_993,In_1183);
or U481 (N_481,In_2164,In_321);
nand U482 (N_482,In_1012,In_1783);
xor U483 (N_483,In_2022,In_2185);
nand U484 (N_484,In_1324,In_709);
xor U485 (N_485,In_868,In_143);
xnor U486 (N_486,In_2588,In_27);
nand U487 (N_487,In_2275,In_1426);
nor U488 (N_488,In_132,In_568);
and U489 (N_489,In_2246,In_907);
or U490 (N_490,In_2287,In_2263);
xnor U491 (N_491,In_1620,In_1525);
nand U492 (N_492,In_2515,In_210);
and U493 (N_493,In_1755,In_1165);
or U494 (N_494,In_2025,In_355);
or U495 (N_495,In_2756,In_249);
and U496 (N_496,In_2469,In_2683);
nor U497 (N_497,In_710,In_2397);
and U498 (N_498,In_478,In_1246);
and U499 (N_499,In_1896,In_1238);
nor U500 (N_500,In_471,In_1761);
xor U501 (N_501,In_1352,In_1384);
nand U502 (N_502,In_686,In_1232);
or U503 (N_503,In_2376,In_614);
nor U504 (N_504,In_312,In_2427);
or U505 (N_505,In_2209,In_1099);
xor U506 (N_506,In_250,In_2001);
or U507 (N_507,In_1076,In_1582);
xor U508 (N_508,In_900,In_2072);
nand U509 (N_509,In_2868,In_749);
nand U510 (N_510,In_1750,In_403);
nand U511 (N_511,In_905,In_113);
or U512 (N_512,In_854,In_2749);
nor U513 (N_513,In_1281,In_898);
nor U514 (N_514,In_2203,In_2871);
nor U515 (N_515,In_1166,In_1647);
nor U516 (N_516,In_2691,In_1650);
xor U517 (N_517,In_1683,In_1699);
xnor U518 (N_518,In_1890,In_780);
xor U519 (N_519,In_1612,In_1470);
or U520 (N_520,In_1038,In_806);
or U521 (N_521,In_2048,In_144);
or U522 (N_522,In_2104,In_1086);
and U523 (N_523,In_447,In_1060);
and U524 (N_524,In_752,In_1619);
nor U525 (N_525,In_1540,In_1710);
or U526 (N_526,In_562,In_1618);
nand U527 (N_527,In_656,In_821);
nand U528 (N_528,In_223,In_2544);
or U529 (N_529,In_188,In_1853);
or U530 (N_530,In_839,In_488);
xnor U531 (N_531,In_2242,In_25);
xnor U532 (N_532,In_84,In_1802);
nand U533 (N_533,In_2033,In_1351);
nand U534 (N_534,In_2637,In_2085);
nor U535 (N_535,In_2540,In_1138);
xor U536 (N_536,In_1284,In_1);
or U537 (N_537,In_2041,In_149);
nand U538 (N_538,In_192,In_580);
and U539 (N_539,In_1408,In_1895);
nor U540 (N_540,In_2205,In_2349);
xor U541 (N_541,In_1446,In_844);
nor U542 (N_542,In_2873,In_1815);
or U543 (N_543,In_2554,In_1645);
nor U544 (N_544,In_2665,In_1672);
nor U545 (N_545,In_1494,In_1256);
xor U546 (N_546,In_8,In_2045);
and U547 (N_547,In_985,In_698);
and U548 (N_548,In_505,In_2950);
and U549 (N_549,In_299,In_16);
or U550 (N_550,In_2493,In_2806);
nor U551 (N_551,In_2633,In_2184);
or U552 (N_552,In_1903,In_2443);
or U553 (N_553,In_2285,In_443);
nor U554 (N_554,In_2389,In_2233);
nor U555 (N_555,In_2042,In_289);
or U556 (N_556,In_1737,In_681);
xnor U557 (N_557,In_2200,In_1681);
or U558 (N_558,In_943,In_431);
xnor U559 (N_559,In_2381,In_1592);
nor U560 (N_560,In_2236,In_2496);
nand U561 (N_561,In_475,In_2234);
nor U562 (N_562,In_711,In_1378);
xnor U563 (N_563,In_1503,In_556);
or U564 (N_564,In_977,In_1510);
nand U565 (N_565,In_1863,In_2957);
nand U566 (N_566,In_1188,In_555);
and U567 (N_567,In_828,In_1694);
or U568 (N_568,In_1367,In_2230);
nor U569 (N_569,In_1958,In_1667);
nand U570 (N_570,In_1261,In_840);
nor U571 (N_571,In_2930,In_1409);
and U572 (N_572,In_2076,In_1279);
nand U573 (N_573,In_1727,In_763);
nand U574 (N_574,In_812,In_97);
nor U575 (N_575,In_2360,In_104);
nand U576 (N_576,In_278,In_1586);
or U577 (N_577,In_2659,In_1869);
or U578 (N_578,In_1286,In_2585);
or U579 (N_579,In_2645,In_1799);
or U580 (N_580,In_1251,In_124);
xor U581 (N_581,In_2575,In_2007);
nor U582 (N_582,In_1732,In_1381);
xnor U583 (N_583,In_1829,In_2060);
nand U584 (N_584,In_506,In_768);
xnor U585 (N_585,In_2455,In_1746);
and U586 (N_586,In_894,In_2913);
nand U587 (N_587,In_83,In_929);
nor U588 (N_588,In_319,In_2762);
xor U589 (N_589,In_90,In_2428);
and U590 (N_590,In_1687,In_2501);
and U591 (N_591,In_927,In_2917);
xnor U592 (N_592,In_2561,In_639);
nor U593 (N_593,In_1071,In_2676);
or U594 (N_594,In_2366,In_2971);
xor U595 (N_595,In_2846,In_2226);
and U596 (N_596,In_2797,In_2375);
nor U597 (N_597,In_794,In_127);
or U598 (N_598,In_2173,In_1855);
nor U599 (N_599,In_791,In_65);
xnor U600 (N_600,In_1010,In_641);
and U601 (N_601,In_850,In_1079);
or U602 (N_602,In_1234,In_1524);
or U603 (N_603,In_1747,In_2015);
and U604 (N_604,In_2800,In_2713);
nor U605 (N_605,In_1571,In_1949);
and U606 (N_606,In_1812,In_1707);
nand U607 (N_607,In_2142,In_402);
xor U608 (N_608,In_1496,In_1127);
xnor U609 (N_609,In_665,In_522);
nor U610 (N_610,In_2255,In_2991);
xnor U611 (N_611,In_2568,In_2811);
and U612 (N_612,In_634,In_269);
xnor U613 (N_613,In_2261,In_343);
and U614 (N_614,In_2553,In_1575);
or U615 (N_615,In_235,In_202);
or U616 (N_616,In_523,In_1854);
nand U617 (N_617,In_2887,In_1911);
or U618 (N_618,In_567,In_374);
nand U619 (N_619,In_1102,In_462);
and U620 (N_620,In_2265,In_2315);
or U621 (N_621,In_499,In_1192);
nand U622 (N_622,In_2121,In_2017);
or U623 (N_623,In_858,In_751);
and U624 (N_624,In_1565,In_1678);
and U625 (N_625,In_1214,In_1872);
and U626 (N_626,In_549,In_101);
nor U627 (N_627,In_226,In_843);
or U628 (N_628,In_2928,In_1098);
and U629 (N_629,In_1023,In_1649);
nor U630 (N_630,In_845,In_177);
and U631 (N_631,In_1216,In_277);
and U632 (N_632,In_1552,In_781);
or U633 (N_633,In_2099,In_2350);
or U634 (N_634,In_2055,In_106);
and U635 (N_635,In_860,In_1942);
nand U636 (N_636,In_147,In_1416);
or U637 (N_637,In_1147,In_153);
or U638 (N_638,In_2155,In_896);
xnor U639 (N_639,In_1585,In_2734);
nor U640 (N_640,In_1196,In_853);
nor U641 (N_641,In_1244,In_792);
or U642 (N_642,In_1866,In_2093);
or U643 (N_643,In_2918,In_1596);
xnor U644 (N_644,In_224,In_100);
nand U645 (N_645,In_536,In_46);
xnor U646 (N_646,In_472,In_1564);
or U647 (N_647,In_178,In_1543);
or U648 (N_648,In_197,In_700);
and U649 (N_649,In_2504,In_1263);
xnor U650 (N_650,In_2002,In_252);
and U651 (N_651,In_667,In_640);
nand U652 (N_652,In_1744,In_1451);
or U653 (N_653,In_1363,In_483);
and U654 (N_654,In_697,In_1912);
nor U655 (N_655,In_716,In_875);
or U656 (N_656,In_2984,In_678);
nand U657 (N_657,In_1325,In_1316);
nand U658 (N_658,In_2577,In_2707);
nor U659 (N_659,In_2970,In_2420);
nand U660 (N_660,In_2323,In_2642);
or U661 (N_661,In_2486,In_1171);
and U662 (N_662,In_2133,In_1267);
and U663 (N_663,In_353,In_198);
and U664 (N_664,In_2108,In_245);
nor U665 (N_665,In_625,In_2564);
or U666 (N_666,In_2243,In_2100);
nand U667 (N_667,In_1566,In_2535);
nand U668 (N_668,In_2011,In_824);
and U669 (N_669,In_2218,In_1977);
or U670 (N_670,In_2937,In_2853);
or U671 (N_671,In_32,In_1394);
and U672 (N_672,In_1362,In_1395);
nor U673 (N_673,In_563,In_1933);
nand U674 (N_674,In_2363,In_1121);
and U675 (N_675,In_2584,In_558);
and U676 (N_676,In_1827,In_2753);
nand U677 (N_677,In_1458,In_2699);
nand U678 (N_678,In_1957,In_1280);
xnor U679 (N_679,In_1801,In_1561);
nand U680 (N_680,In_802,In_1808);
xnor U681 (N_681,In_1348,In_2039);
or U682 (N_682,In_2643,In_2404);
or U683 (N_683,In_1046,In_2210);
xnor U684 (N_684,In_1422,In_1307);
nor U685 (N_685,In_1553,In_1606);
nor U686 (N_686,In_2303,In_33);
nand U687 (N_687,In_2541,In_306);
nor U688 (N_688,In_2546,In_2408);
nor U689 (N_689,In_10,In_1472);
or U690 (N_690,In_1265,In_1666);
nor U691 (N_691,In_583,In_377);
and U692 (N_692,In_2008,In_655);
xor U693 (N_693,In_2994,In_2131);
xnor U694 (N_694,In_1826,In_831);
nor U695 (N_695,In_607,In_1050);
and U696 (N_696,In_2883,In_62);
or U697 (N_697,In_272,In_1492);
and U698 (N_698,In_1793,In_1399);
and U699 (N_699,In_2452,In_199);
or U700 (N_700,In_2715,In_1633);
or U701 (N_701,In_2247,In_63);
xor U702 (N_702,In_2223,In_219);
or U703 (N_703,In_2050,In_2449);
xnor U704 (N_704,In_1459,In_662);
or U705 (N_705,In_1753,In_122);
xnor U706 (N_706,In_688,In_1995);
nor U707 (N_707,In_2402,In_2186);
nor U708 (N_708,In_1778,In_495);
nor U709 (N_709,In_1731,In_832);
and U710 (N_710,In_1505,In_171);
xor U711 (N_711,In_2788,In_979);
nor U712 (N_712,In_2840,In_2824);
and U713 (N_713,In_2088,In_1202);
nor U714 (N_714,In_577,In_2782);
or U715 (N_715,In_2152,In_304);
xor U716 (N_716,In_2139,In_2272);
nor U717 (N_717,In_1437,In_1243);
or U718 (N_718,In_1181,In_679);
nor U719 (N_719,In_2992,In_2977);
nand U720 (N_720,In_961,In_1045);
nor U721 (N_721,In_201,In_458);
and U722 (N_722,In_963,In_1786);
nor U723 (N_723,In_2823,In_1433);
nand U724 (N_724,In_125,In_2761);
nor U725 (N_725,In_1580,In_2947);
or U726 (N_726,In_2477,In_507);
or U727 (N_727,In_266,In_1154);
nor U728 (N_728,In_642,In_2495);
nand U729 (N_729,In_354,In_407);
and U730 (N_730,In_1164,In_2374);
or U731 (N_731,In_881,In_732);
xnor U732 (N_732,In_1136,In_1124);
or U733 (N_733,In_826,In_1039);
nand U734 (N_734,In_115,In_637);
nor U735 (N_735,In_123,In_2013);
or U736 (N_736,In_2167,In_38);
nand U737 (N_737,In_1412,In_2158);
or U738 (N_738,In_999,In_1570);
nor U739 (N_739,In_2475,In_2556);
nand U740 (N_740,In_1613,In_1125);
xnor U741 (N_741,In_2759,In_2862);
and U742 (N_742,In_2197,In_1100);
or U743 (N_743,In_988,In_1705);
and U744 (N_744,In_2010,In_1024);
xor U745 (N_745,In_693,In_1791);
xnor U746 (N_746,In_2606,In_994);
or U747 (N_747,In_755,In_1146);
nor U748 (N_748,In_1634,In_1603);
and U749 (N_749,In_1402,In_1382);
nor U750 (N_750,In_1868,In_1135);
nor U751 (N_751,In_2818,In_2766);
nor U752 (N_752,In_1594,In_1419);
and U753 (N_753,In_2714,In_110);
and U754 (N_754,In_2599,In_1991);
nor U755 (N_755,In_2897,In_2668);
or U756 (N_756,In_92,In_1432);
and U757 (N_757,In_240,In_1700);
nor U758 (N_758,In_841,In_1945);
xor U759 (N_759,In_1541,In_541);
or U760 (N_760,In_2047,In_1990);
nor U761 (N_761,In_2600,In_2165);
nand U762 (N_762,In_2731,In_1441);
or U763 (N_763,In_1278,In_1162);
nand U764 (N_764,In_1677,In_2987);
xnor U765 (N_765,In_2385,In_2347);
or U766 (N_766,In_582,In_50);
nand U767 (N_767,In_2934,In_2842);
or U768 (N_768,In_1271,In_2737);
nor U769 (N_769,In_2114,In_1142);
nand U770 (N_770,In_2168,In_1535);
and U771 (N_771,In_1063,In_1040);
xor U772 (N_772,In_2091,In_98);
nor U773 (N_773,In_1051,In_2935);
and U774 (N_774,In_473,In_2422);
nand U775 (N_775,In_1034,In_2157);
or U776 (N_776,In_546,In_2057);
nand U777 (N_777,In_1122,In_1078);
or U778 (N_778,In_325,In_997);
xor U779 (N_779,In_2594,In_1057);
xor U780 (N_780,In_829,In_378);
nand U781 (N_781,In_246,In_2414);
and U782 (N_782,In_2474,In_2229);
or U783 (N_783,In_1315,In_359);
xnor U784 (N_784,In_273,In_519);
and U785 (N_785,In_535,In_605);
and U786 (N_786,In_1499,In_174);
xnor U787 (N_787,In_552,In_1749);
nor U788 (N_788,In_322,In_2118);
nand U789 (N_789,In_1856,In_1311);
nor U790 (N_790,In_2354,In_2494);
and U791 (N_791,In_301,In_1417);
nand U792 (N_792,In_953,In_865);
nor U793 (N_793,In_2127,In_2169);
xor U794 (N_794,In_941,In_1218);
or U795 (N_795,In_1661,In_2773);
nor U796 (N_796,In_1548,In_1262);
xnor U797 (N_797,In_1149,In_1304);
nor U798 (N_798,In_1215,In_2738);
nand U799 (N_799,In_846,In_1572);
or U800 (N_800,In_925,In_2832);
and U801 (N_801,In_1294,In_244);
nor U802 (N_802,In_372,In_1549);
nand U803 (N_803,In_1042,In_1550);
nor U804 (N_804,In_1701,In_39);
or U805 (N_805,In_1052,In_1386);
nor U806 (N_806,In_1693,In_972);
and U807 (N_807,In_1542,In_2300);
or U808 (N_808,In_1049,In_2239);
or U809 (N_809,In_2885,In_836);
xor U810 (N_810,In_620,In_2401);
or U811 (N_811,In_1283,In_2936);
or U812 (N_812,In_454,In_509);
nor U813 (N_813,In_2517,In_2497);
xnor U814 (N_814,In_2639,In_1016);
or U815 (N_815,In_776,In_530);
nand U816 (N_816,In_1567,In_2249);
and U817 (N_817,In_566,In_1272);
or U818 (N_818,In_878,In_2081);
nand U819 (N_819,In_2192,In_2171);
and U820 (N_820,In_1970,In_2291);
and U821 (N_821,In_2423,In_173);
nor U822 (N_822,In_2866,In_412);
xor U823 (N_823,In_513,In_2489);
and U824 (N_824,In_461,In_1983);
or U825 (N_825,In_1072,In_2563);
nand U826 (N_826,In_946,In_1555);
nand U827 (N_827,In_585,In_1306);
xnor U828 (N_828,In_6,In_1875);
xnor U829 (N_829,In_1712,In_131);
or U830 (N_830,In_2827,In_2888);
and U831 (N_831,In_282,In_1529);
nor U832 (N_832,In_350,In_441);
nor U833 (N_833,In_2442,In_2361);
or U834 (N_834,In_2292,In_2327);
and U835 (N_835,In_1733,In_1444);
nand U836 (N_836,In_2122,In_1627);
nand U837 (N_837,In_15,In_2409);
nor U838 (N_838,In_2313,In_2607);
nand U839 (N_839,In_1018,In_1295);
or U840 (N_840,In_255,In_770);
xnor U841 (N_841,In_2086,In_2346);
or U842 (N_842,In_2332,In_653);
nor U843 (N_843,In_45,In_492);
and U844 (N_844,In_2049,In_2299);
nor U845 (N_845,In_247,In_1643);
xor U846 (N_846,In_1845,In_2552);
nand U847 (N_847,In_2160,In_493);
nand U848 (N_848,In_2392,In_746);
nor U849 (N_849,In_586,In_622);
nor U850 (N_850,In_783,In_2669);
and U851 (N_851,In_574,In_2876);
xor U852 (N_852,In_1919,In_2940);
nor U853 (N_853,In_1285,In_811);
and U854 (N_854,In_2355,In_194);
and U855 (N_855,In_2983,In_1141);
and U856 (N_856,In_1290,In_510);
or U857 (N_857,In_978,In_2339);
xnor U858 (N_858,In_1400,In_2370);
nor U859 (N_859,In_433,In_1803);
nand U860 (N_860,In_1923,In_2388);
nor U861 (N_861,In_1556,In_2512);
nand U862 (N_862,In_1157,In_2895);
and U863 (N_863,In_695,In_2325);
nor U864 (N_864,In_367,In_2569);
nand U865 (N_865,In_1810,In_356);
nor U866 (N_866,In_425,In_624);
xor U867 (N_867,In_818,In_796);
nor U868 (N_868,In_365,In_735);
nor U869 (N_869,In_271,In_1003);
nand U870 (N_870,In_1779,In_1909);
xnor U871 (N_871,In_2727,In_760);
and U872 (N_872,In_611,In_1447);
xor U873 (N_873,In_405,In_1537);
nor U874 (N_874,In_2473,In_1277);
nor U875 (N_875,In_2805,In_2498);
nand U876 (N_876,In_494,In_168);
and U877 (N_877,In_1703,In_58);
xnor U878 (N_878,In_584,In_335);
nand U879 (N_879,In_2273,In_2965);
and U880 (N_880,In_362,In_906);
and U881 (N_881,In_1531,In_798);
xnor U882 (N_882,In_1921,In_919);
and U883 (N_883,In_1788,In_2867);
and U884 (N_884,In_877,In_989);
nand U885 (N_885,In_901,In_292);
nor U886 (N_886,In_2284,In_2419);
xnor U887 (N_887,In_1155,In_2884);
or U888 (N_888,In_328,In_1241);
or U889 (N_889,In_960,In_1968);
xnor U890 (N_890,In_533,In_376);
and U891 (N_891,In_2170,In_1907);
xnor U892 (N_892,In_937,In_944);
nand U893 (N_893,In_486,In_2616);
nor U894 (N_894,In_1590,In_369);
nor U895 (N_895,In_435,In_1841);
nand U896 (N_896,In_928,In_349);
nand U897 (N_897,In_1574,In_965);
xor U898 (N_898,In_1087,In_2305);
nor U899 (N_899,In_2129,In_689);
nand U900 (N_900,In_2324,In_2698);
nand U901 (N_901,In_476,In_1004);
xor U902 (N_902,In_1777,In_324);
xnor U903 (N_903,In_419,In_2334);
or U904 (N_904,In_118,In_1820);
nor U905 (N_905,In_1344,In_1008);
nor U906 (N_906,In_1109,In_2431);
or U907 (N_907,In_1528,In_1610);
nor U908 (N_908,In_2282,In_2724);
xnor U909 (N_909,In_983,In_2519);
nor U910 (N_910,In_857,In_2043);
nand U911 (N_911,In_13,In_649);
xor U912 (N_912,In_54,In_950);
nor U913 (N_913,In_2722,In_119);
nor U914 (N_914,In_242,In_2831);
and U915 (N_915,In_2765,In_1611);
and U916 (N_916,In_1260,In_2576);
or U917 (N_917,In_571,In_190);
nand U918 (N_918,In_418,In_2460);
or U919 (N_919,In_1697,In_2735);
or U920 (N_920,In_293,In_1184);
nor U921 (N_921,In_213,In_615);
nand U922 (N_922,In_200,In_154);
nor U923 (N_923,In_363,In_1743);
or U924 (N_924,In_633,In_1343);
and U925 (N_925,In_326,In_1297);
nor U926 (N_926,In_1097,In_2393);
or U927 (N_927,In_1523,In_253);
xor U928 (N_928,In_2877,In_75);
nor U929 (N_929,In_2137,In_2949);
nor U930 (N_930,In_916,In_2479);
nand U931 (N_931,In_1420,In_89);
and U932 (N_932,In_1266,In_1763);
nand U933 (N_933,In_886,In_256);
and U934 (N_934,In_2471,In_2456);
nor U935 (N_935,In_415,In_348);
nor U936 (N_936,In_756,In_468);
nor U937 (N_937,In_1355,In_2601);
xor U938 (N_938,In_1185,In_2911);
xnor U939 (N_939,In_2135,In_239);
xor U940 (N_940,In_1370,In_409);
nand U941 (N_941,In_1463,In_2764);
or U942 (N_942,In_1804,In_627);
nor U943 (N_943,In_2437,In_2270);
or U944 (N_944,In_1201,In_142);
nor U945 (N_945,In_731,In_575);
xnor U946 (N_946,In_391,In_225);
or U947 (N_947,In_2178,In_417);
and U948 (N_948,In_2615,In_1939);
or U949 (N_949,In_109,In_1410);
xor U950 (N_950,In_7,In_2820);
xor U951 (N_951,In_1228,In_1077);
nand U952 (N_952,In_1877,In_1924);
nand U953 (N_953,In_2627,In_1943);
nand U954 (N_954,In_534,In_551);
nor U955 (N_955,In_1118,In_511);
or U956 (N_956,In_1960,In_691);
nand U957 (N_957,In_2035,In_2220);
nand U958 (N_958,In_867,In_855);
nor U959 (N_959,In_170,In_722);
xnor U960 (N_960,In_932,In_2916);
or U961 (N_961,In_1922,In_2365);
and U962 (N_962,In_1101,In_1870);
nor U963 (N_963,In_2179,In_1193);
xnor U964 (N_964,In_2144,In_685);
and U965 (N_965,In_1857,In_108);
xnor U966 (N_966,In_2624,In_2586);
xor U967 (N_967,In_1210,In_2024);
xnor U968 (N_968,In_2524,In_992);
xnor U969 (N_969,In_1502,In_2981);
and U970 (N_970,In_866,In_1061);
nor U971 (N_971,In_785,In_870);
nand U972 (N_972,In_52,In_243);
nor U973 (N_973,In_1156,In_1830);
nor U974 (N_974,In_1404,In_2974);
xnor U975 (N_975,In_1110,In_2426);
xor U976 (N_976,In_2330,In_2995);
and U977 (N_977,In_2819,In_1320);
and U978 (N_978,In_767,In_217);
xnor U979 (N_979,In_2744,In_2963);
nand U980 (N_980,In_2798,In_2750);
or U981 (N_981,In_851,In_807);
nand U982 (N_982,In_2650,In_2838);
or U983 (N_983,In_981,In_2898);
nand U984 (N_984,In_2975,In_2925);
nor U985 (N_985,In_827,In_2457);
xor U986 (N_986,In_2016,In_2028);
nor U987 (N_987,In_720,In_2511);
nor U988 (N_988,In_2851,In_2194);
nor U989 (N_989,In_1226,In_357);
xor U990 (N_990,In_1604,In_291);
xnor U991 (N_991,In_2036,In_11);
nor U992 (N_992,In_2816,In_2622);
xnor U993 (N_993,In_847,In_1576);
and U994 (N_994,In_1391,In_1319);
and U995 (N_995,In_176,In_2728);
nand U996 (N_996,In_2886,In_1831);
or U997 (N_997,In_81,In_910);
nand U998 (N_998,In_413,In_2483);
nor U999 (N_999,In_2279,In_2833);
or U1000 (N_1000,In_2845,In_2653);
or U1001 (N_1001,In_2829,In_2379);
and U1002 (N_1002,In_1380,In_1177);
xor U1003 (N_1003,In_1222,In_526);
or U1004 (N_1004,In_1032,In_861);
nor U1005 (N_1005,In_2872,In_1579);
and U1006 (N_1006,In_2863,In_1851);
xor U1007 (N_1007,In_2207,In_1704);
nor U1008 (N_1008,In_889,In_837);
xnor U1009 (N_1009,In_2297,In_2089);
or U1010 (N_1010,In_264,In_1242);
nor U1011 (N_1011,In_2543,In_2560);
nand U1012 (N_1012,In_222,In_459);
nor U1013 (N_1013,In_669,In_2527);
and U1014 (N_1014,In_968,In_1593);
nand U1015 (N_1015,In_852,In_2415);
and U1016 (N_1016,In_2708,In_2875);
xor U1017 (N_1017,In_1014,In_401);
nand U1018 (N_1018,In_1888,In_2154);
nor U1019 (N_1019,In_1608,In_2405);
nand U1020 (N_1020,In_71,In_2684);
and U1021 (N_1021,In_2267,In_2667);
nor U1022 (N_1022,In_2078,In_456);
and U1023 (N_1023,In_647,In_1427);
and U1024 (N_1024,In_382,In_1383);
nor U1025 (N_1025,In_1536,In_2328);
xor U1026 (N_1026,In_346,In_218);
nand U1027 (N_1027,In_1020,In_1518);
or U1028 (N_1028,In_1015,In_1123);
and U1029 (N_1029,In_2096,In_2580);
or U1030 (N_1030,In_2026,In_1790);
nand U1031 (N_1031,In_1828,In_1679);
and U1032 (N_1032,In_1103,In_205);
xnor U1033 (N_1033,In_616,In_1640);
or U1034 (N_1034,In_1655,In_1487);
nand U1035 (N_1035,In_1490,In_429);
xnor U1036 (N_1036,In_2739,In_2572);
or U1037 (N_1037,In_2188,In_385);
nand U1038 (N_1038,In_2321,In_1989);
or U1039 (N_1039,In_1941,In_2396);
or U1040 (N_1040,In_195,In_1298);
and U1041 (N_1041,In_2240,In_2657);
and U1042 (N_1042,In_2335,In_2904);
or U1043 (N_1043,In_2682,In_1313);
nand U1044 (N_1044,In_2244,In_1163);
or U1045 (N_1045,In_1944,In_2208);
and U1046 (N_1046,In_186,In_1443);
and U1047 (N_1047,In_423,In_1918);
and U1048 (N_1048,In_990,In_2095);
nand U1049 (N_1049,In_2312,In_540);
nand U1050 (N_1050,In_2138,In_726);
or U1051 (N_1051,In_280,In_2235);
nand U1052 (N_1052,In_2413,In_2780);
nand U1053 (N_1053,In_1392,In_966);
nand U1054 (N_1054,In_537,In_548);
or U1055 (N_1055,In_2850,In_1461);
nand U1056 (N_1056,In_2193,In_1848);
nor U1057 (N_1057,In_263,In_660);
and U1058 (N_1058,In_360,In_2311);
nor U1059 (N_1059,In_107,In_1473);
nor U1060 (N_1060,In_1559,In_2071);
or U1061 (N_1061,In_2654,In_797);
nor U1062 (N_1062,In_74,In_53);
or U1063 (N_1063,In_439,In_2678);
and U1064 (N_1064,In_1685,In_2736);
nand U1065 (N_1065,In_2439,In_2685);
and U1066 (N_1066,In_408,In_2020);
and U1067 (N_1067,In_1545,In_1131);
nor U1068 (N_1068,In_1195,In_2661);
and U1069 (N_1069,In_2367,In_1996);
nand U1070 (N_1070,In_842,In_2882);
and U1071 (N_1071,In_2206,In_719);
nor U1072 (N_1072,In_1953,In_2921);
nor U1073 (N_1073,In_604,In_628);
and U1074 (N_1074,In_2507,In_1361);
or U1075 (N_1075,In_931,In_553);
nand U1076 (N_1076,In_1104,In_833);
xnor U1077 (N_1077,In_1369,In_1221);
nor U1078 (N_1078,In_380,In_2809);
and U1079 (N_1079,In_2912,In_1309);
nor U1080 (N_1080,In_702,In_1245);
xor U1081 (N_1081,In_1092,In_41);
and U1082 (N_1082,In_737,In_370);
nor U1083 (N_1083,In_1657,In_498);
xnor U1084 (N_1084,In_191,In_1928);
and U1085 (N_1085,In_952,In_1331);
nand U1086 (N_1086,In_1128,In_902);
xnor U1087 (N_1087,In_2996,In_2031);
nor U1088 (N_1088,In_810,In_175);
or U1089 (N_1089,In_2130,In_2723);
nand U1090 (N_1090,In_1515,In_426);
or U1091 (N_1091,In_1303,In_2387);
and U1092 (N_1092,In_399,In_1948);
or U1093 (N_1093,In_1493,In_1268);
nand U1094 (N_1094,In_2926,In_2972);
nor U1095 (N_1095,In_260,In_2106);
nor U1096 (N_1096,In_2505,In_1288);
nand U1097 (N_1097,In_2777,In_2711);
and U1098 (N_1098,In_2034,In_2418);
or U1099 (N_1099,In_2785,In_1637);
or U1100 (N_1100,In_1091,In_1220);
nor U1101 (N_1101,In_1276,In_2352);
nand U1102 (N_1102,In_630,In_281);
and U1103 (N_1103,In_814,In_2172);
and U1104 (N_1104,In_2537,In_238);
xor U1105 (N_1105,In_1740,In_893);
nor U1106 (N_1106,In_2686,In_2843);
nor U1107 (N_1107,In_1858,In_1885);
nand U1108 (N_1108,In_389,In_1695);
nor U1109 (N_1109,In_2180,In_2040);
xor U1110 (N_1110,In_2065,In_1194);
and U1111 (N_1111,In_825,In_2254);
nor U1112 (N_1112,In_215,In_156);
and U1113 (N_1113,In_2570,In_445);
and U1114 (N_1114,In_650,In_1393);
or U1115 (N_1115,In_482,In_2000);
xor U1116 (N_1116,In_2604,In_2268);
and U1117 (N_1117,In_2826,In_1428);
or U1118 (N_1118,In_1478,In_918);
nand U1119 (N_1119,In_383,In_2597);
nor U1120 (N_1120,In_1457,In_1609);
and U1121 (N_1121,In_1691,In_2212);
and U1122 (N_1122,In_788,In_670);
and U1123 (N_1123,In_892,In_1089);
nand U1124 (N_1124,In_2238,In_724);
and U1125 (N_1125,In_1174,In_2224);
or U1126 (N_1126,In_2044,In_2841);
nor U1127 (N_1127,In_1225,In_2745);
xor U1128 (N_1128,In_1453,In_1096);
nor U1129 (N_1129,In_1901,In_2620);
nand U1130 (N_1130,In_469,In_2513);
nand U1131 (N_1131,In_2617,In_2889);
and U1132 (N_1132,In_1843,In_140);
nand U1133 (N_1133,In_2262,In_294);
nand U1134 (N_1134,In_1646,In_1738);
xor U1135 (N_1135,In_987,In_329);
xor U1136 (N_1136,In_504,In_2271);
nor U1137 (N_1137,In_19,In_2658);
and U1138 (N_1138,In_116,In_1999);
or U1139 (N_1139,In_1335,In_318);
or U1140 (N_1140,In_957,In_945);
nand U1141 (N_1141,In_2383,In_1489);
and U1142 (N_1142,In_2510,In_1029);
or U1143 (N_1143,In_309,In_102);
or U1144 (N_1144,In_730,In_917);
or U1145 (N_1145,In_1752,In_2296);
or U1146 (N_1146,In_2211,In_1002);
nor U1147 (N_1147,In_2466,In_1129);
and U1148 (N_1148,In_2726,In_2675);
nor U1149 (N_1149,In_1532,In_2989);
nor U1150 (N_1150,In_381,In_676);
or U1151 (N_1151,In_2944,In_1668);
xor U1152 (N_1152,In_2704,In_2536);
xor U1153 (N_1153,In_2283,In_663);
or U1154 (N_1154,In_1456,In_923);
nor U1155 (N_1155,In_1862,In_773);
nand U1156 (N_1156,In_2621,In_2514);
xor U1157 (N_1157,In_2951,In_1951);
xor U1158 (N_1158,In_2182,In_428);
xnor U1159 (N_1159,In_2896,In_2037);
nor U1160 (N_1160,In_2174,In_420);
nand U1161 (N_1161,In_1925,In_1675);
nor U1162 (N_1162,In_338,In_2815);
nor U1163 (N_1163,In_1482,In_1973);
and U1164 (N_1164,In_270,In_2976);
or U1165 (N_1165,In_1947,In_2980);
nand U1166 (N_1166,In_2087,In_31);
nor U1167 (N_1167,In_2700,In_2062);
and U1168 (N_1168,In_2857,In_1484);
or U1169 (N_1169,In_984,In_2664);
nor U1170 (N_1170,In_1624,In_2264);
xnor U1171 (N_1171,In_926,In_784);
nand U1172 (N_1172,In_1088,In_2395);
xor U1173 (N_1173,In_2874,In_1179);
or U1174 (N_1174,In_2368,In_2216);
and U1175 (N_1175,In_1507,In_157);
or U1176 (N_1176,In_2398,In_2196);
and U1177 (N_1177,In_1771,In_1760);
nor U1178 (N_1178,In_29,In_2706);
or U1179 (N_1179,In_2416,In_1385);
nor U1180 (N_1180,In_2499,In_414);
and U1181 (N_1181,In_908,In_128);
and U1182 (N_1182,In_1979,In_2472);
xor U1183 (N_1183,In_410,In_432);
xnor U1184 (N_1184,In_1998,In_1372);
nor U1185 (N_1185,In_544,In_2692);
and U1186 (N_1186,In_1664,In_2251);
nand U1187 (N_1187,In_1711,In_1423);
or U1188 (N_1188,In_2786,In_1839);
nand U1189 (N_1189,In_2687,In_800);
and U1190 (N_1190,In_165,In_2412);
and U1191 (N_1191,In_341,In_69);
xnor U1192 (N_1192,In_145,In_1116);
nand U1193 (N_1193,In_2956,In_1894);
xor U1194 (N_1194,In_196,In_2593);
xnor U1195 (N_1195,In_1938,In_599);
xor U1196 (N_1196,In_1411,In_1009);
or U1197 (N_1197,In_42,In_1070);
nand U1198 (N_1198,In_2958,In_786);
nor U1199 (N_1199,In_2631,In_882);
or U1200 (N_1200,In_126,In_572);
xor U1201 (N_1201,In_2861,In_1974);
and U1202 (N_1202,In_1143,In_2595);
and U1203 (N_1203,In_2808,In_1833);
xnor U1204 (N_1204,In_1954,In_1584);
nor U1205 (N_1205,In_1534,In_1842);
xnor U1206 (N_1206,In_2150,In_2779);
nand U1207 (N_1207,In_57,In_1935);
xnor U1208 (N_1208,In_600,In_2068);
nor U1209 (N_1209,In_2103,In_884);
and U1210 (N_1210,In_283,In_80);
or U1211 (N_1211,In_1030,In_21);
or U1212 (N_1212,In_1137,In_352);
and U1213 (N_1213,In_2107,In_1615);
nand U1214 (N_1214,In_1825,In_2407);
xnor U1215 (N_1215,In_2854,In_1407);
nor U1216 (N_1216,In_1065,In_184);
or U1217 (N_1217,In_2879,In_2338);
or U1218 (N_1218,In_1292,In_185);
or U1219 (N_1219,In_2444,In_1626);
xor U1220 (N_1220,In_268,In_1914);
nand U1221 (N_1221,In_1173,In_942);
nor U1222 (N_1222,In_484,In_734);
and U1223 (N_1223,In_1206,In_2424);
nand U1224 (N_1224,In_920,In_1191);
or U1225 (N_1225,In_793,In_40);
xor U1226 (N_1226,In_347,In_949);
xnor U1227 (N_1227,In_1539,In_593);
or U1228 (N_1228,In_2893,In_2113);
and U1229 (N_1229,In_2689,In_1345);
or U1230 (N_1230,In_2331,In_2232);
nor U1231 (N_1231,In_2632,In_2061);
xor U1232 (N_1232,In_398,In_813);
and U1233 (N_1233,In_739,In_512);
xnor U1234 (N_1234,In_1773,In_274);
xnor U1235 (N_1235,In_187,In_1940);
and U1236 (N_1236,In_2844,In_1573);
nand U1237 (N_1237,In_1022,In_411);
or U1238 (N_1238,In_1217,In_668);
nand U1239 (N_1239,In_2941,In_2438);
or U1240 (N_1240,In_1480,In_2490);
and U1241 (N_1241,In_591,In_1318);
xnor U1242 (N_1242,In_2848,In_2124);
nor U1243 (N_1243,In_2484,In_2237);
or U1244 (N_1244,In_394,In_1526);
nor U1245 (N_1245,In_1161,In_652);
or U1246 (N_1246,In_1388,In_2758);
xor U1247 (N_1247,In_1723,In_2032);
or U1248 (N_1248,In_838,In_648);
or U1249 (N_1249,In_859,In_2839);
nor U1250 (N_1250,In_167,In_44);
or U1251 (N_1251,In_729,In_1671);
and U1252 (N_1252,In_766,In_517);
and U1253 (N_1253,In_463,In_1464);
or U1254 (N_1254,In_2441,In_2646);
and U1255 (N_1255,In_1720,In_2260);
and U1256 (N_1256,In_856,In_2377);
and U1257 (N_1257,In_1431,In_2725);
nor U1258 (N_1258,In_2609,In_2579);
or U1259 (N_1259,In_1721,In_1837);
and U1260 (N_1260,In_2952,In_2855);
nor U1261 (N_1261,In_1985,In_9);
and U1262 (N_1262,In_2447,In_704);
nor U1263 (N_1263,In_1258,In_765);
xnor U1264 (N_1264,In_612,In_801);
nand U1265 (N_1265,In_775,In_1756);
nand U1266 (N_1266,In_1474,In_2549);
xor U1267 (N_1267,In_3,In_487);
xor U1268 (N_1268,In_1209,In_297);
nor U1269 (N_1269,In_1094,In_2906);
or U1270 (N_1270,In_1257,In_1658);
xor U1271 (N_1271,In_1601,In_1434);
nor U1272 (N_1272,In_1832,In_2836);
nor U1273 (N_1273,In_715,In_590);
nand U1274 (N_1274,In_2721,In_1413);
or U1275 (N_1275,In_1708,In_684);
xor U1276 (N_1276,In_1329,In_203);
or U1277 (N_1277,In_545,In_43);
nand U1278 (N_1278,In_2435,In_1500);
nand U1279 (N_1279,In_1168,In_2929);
xnor U1280 (N_1280,In_2163,In_310);
or U1281 (N_1281,In_914,In_973);
and U1282 (N_1282,In_2990,In_1436);
and U1283 (N_1283,In_2399,In_1273);
xor U1284 (N_1284,In_2448,In_1554);
xor U1285 (N_1285,In_387,In_1342);
and U1286 (N_1286,In_779,In_2748);
and U1287 (N_1287,In_67,In_2219);
or U1288 (N_1288,In_1483,In_2757);
or U1289 (N_1289,In_216,In_1824);
and U1290 (N_1290,In_139,In_876);
or U1291 (N_1291,In_257,In_146);
xnor U1292 (N_1292,In_334,In_2961);
nand U1293 (N_1293,In_2487,In_503);
or U1294 (N_1294,In_1080,In_2115);
nand U1295 (N_1295,In_1390,In_2421);
and U1296 (N_1296,In_214,In_2985);
nand U1297 (N_1297,In_594,In_181);
xor U1298 (N_1298,In_528,In_2793);
nand U1299 (N_1299,In_22,In_2480);
or U1300 (N_1300,In_163,In_120);
nor U1301 (N_1301,In_2968,In_451);
nor U1302 (N_1302,In_2146,In_2252);
and U1303 (N_1303,In_2909,In_1090);
xnor U1304 (N_1304,In_2988,In_1557);
and U1305 (N_1305,In_2892,In_1577);
and U1306 (N_1306,In_1665,In_1587);
xnor U1307 (N_1307,In_1817,In_1984);
nor U1308 (N_1308,In_613,In_1653);
nand U1309 (N_1309,In_1900,In_883);
xnor U1310 (N_1310,In_1882,In_2740);
or U1311 (N_1311,In_1781,In_1006);
nor U1312 (N_1312,In_707,In_1066);
nor U1313 (N_1313,In_769,In_259);
xnor U1314 (N_1314,In_1150,In_345);
xnor U1315 (N_1315,In_1084,In_1988);
nor U1316 (N_1316,In_1768,In_1160);
xor U1317 (N_1317,In_1479,In_2719);
nor U1318 (N_1318,In_1569,In_70);
xnor U1319 (N_1319,In_2063,In_1838);
xor U1320 (N_1320,In_569,In_2214);
nand U1321 (N_1321,In_723,In_1247);
or U1322 (N_1322,In_2696,In_2191);
xor U1323 (N_1323,In_816,In_2768);
and U1324 (N_1324,In_1322,In_2465);
xnor U1325 (N_1325,In_481,In_1108);
nor U1326 (N_1326,In_2454,In_2278);
and U1327 (N_1327,In_2329,In_1139);
xor U1328 (N_1328,In_340,In_169);
nor U1329 (N_1329,In_2353,In_2120);
xnor U1330 (N_1330,In_1429,In_587);
nand U1331 (N_1331,In_1375,In_1950);
and U1332 (N_1332,In_2948,In_302);
nand U1333 (N_1333,In_2343,In_2520);
nor U1334 (N_1334,In_1659,In_714);
or U1335 (N_1335,In_1849,In_364);
and U1336 (N_1336,In_2763,In_2084);
nor U1337 (N_1337,In_2110,In_2485);
xor U1338 (N_1338,In_99,In_542);
or U1339 (N_1339,In_2356,In_1904);
nand U1340 (N_1340,In_515,In_936);
xor U1341 (N_1341,In_2656,In_286);
and U1342 (N_1342,In_2526,In_2101);
xnor U1343 (N_1343,In_862,In_2835);
nor U1344 (N_1344,In_2539,In_1663);
nor U1345 (N_1345,In_699,In_680);
nand U1346 (N_1346,In_2319,In_1170);
and U1347 (N_1347,In_1656,In_1717);
nor U1348 (N_1348,In_1835,In_1485);
nand U1349 (N_1349,In_59,In_49);
xor U1350 (N_1350,In_2289,In_2946);
and U1351 (N_1351,In_1780,In_37);
and U1352 (N_1352,In_1871,In_2080);
and U1353 (N_1353,In_820,In_2384);
xor U1354 (N_1354,In_815,In_384);
or U1355 (N_1355,In_1074,In_323);
and U1356 (N_1356,In_646,In_848);
and U1357 (N_1357,In_344,In_2256);
nor U1358 (N_1358,In_1338,In_976);
nor U1359 (N_1359,In_1725,In_2660);
xor U1360 (N_1360,In_2856,In_1867);
or U1361 (N_1361,In_817,In_448);
or U1362 (N_1362,In_1816,In_2673);
and U1363 (N_1363,In_1622,In_155);
nor U1364 (N_1364,In_491,In_2680);
nor U1365 (N_1365,In_1328,In_759);
xnor U1366 (N_1366,In_835,In_694);
nand U1367 (N_1367,In_1676,In_93);
or U1368 (N_1368,In_2959,In_1765);
nor U1369 (N_1369,In_2555,In_2075);
nor U1370 (N_1370,In_1151,In_1204);
or U1371 (N_1371,In_1152,In_692);
nor U1372 (N_1372,In_1729,In_899);
nand U1373 (N_1373,In_1007,In_2794);
and U1374 (N_1374,In_2810,In_2153);
xor U1375 (N_1375,In_2481,In_1397);
xnor U1376 (N_1376,In_2784,In_1212);
nor U1377 (N_1377,In_1323,In_1591);
nand U1378 (N_1378,In_2295,In_2625);
and U1379 (N_1379,In_708,In_1180);
and U1380 (N_1380,In_772,In_2529);
or U1381 (N_1381,In_1033,In_706);
or U1382 (N_1382,In_1448,In_2358);
xor U1383 (N_1383,In_2870,In_2583);
xnor U1384 (N_1384,In_2307,In_453);
and U1385 (N_1385,In_1709,In_589);
nand U1386 (N_1386,In_1639,In_2582);
and U1387 (N_1387,In_559,In_598);
xnor U1388 (N_1388,In_1357,In_1544);
or U1389 (N_1389,In_2317,In_1880);
nor U1390 (N_1390,In_2021,In_457);
nor U1391 (N_1391,In_2464,In_1414);
xor U1392 (N_1392,In_1992,In_897);
nand U1393 (N_1393,In_2482,In_2281);
nand U1394 (N_1394,In_1978,In_2440);
or U1395 (N_1395,In_2221,In_2029);
nand U1396 (N_1396,In_1964,In_2799);
and U1397 (N_1397,In_1175,In_2635);
or U1398 (N_1398,In_368,In_2858);
or U1399 (N_1399,In_521,In_508);
or U1400 (N_1400,In_2257,In_479);
xnor U1401 (N_1401,In_1230,In_2468);
xnor U1402 (N_1402,In_2796,In_2293);
nor U1403 (N_1403,In_774,In_938);
or U1404 (N_1404,In_61,In_2500);
nor U1405 (N_1405,In_36,In_610);
or U1406 (N_1406,In_1504,In_489);
and U1407 (N_1407,In_2551,In_307);
and U1408 (N_1408,In_2531,In_1250);
xnor U1409 (N_1409,In_873,In_1145);
or U1410 (N_1410,In_18,In_629);
and U1411 (N_1411,In_212,In_1095);
and U1412 (N_1412,In_2241,In_241);
and U1413 (N_1413,In_1293,In_392);
xor U1414 (N_1414,In_48,In_619);
xor U1415 (N_1415,In_390,In_2126);
nor U1416 (N_1416,In_1013,In_2837);
and U1417 (N_1417,In_228,In_969);
or U1418 (N_1418,In_874,In_455);
and U1419 (N_1419,In_331,In_2027);
xnor U1420 (N_1420,In_1797,In_2425);
nand U1421 (N_1421,In_1354,In_1353);
or U1422 (N_1422,In_1792,In_303);
xnor U1423 (N_1423,In_1636,In_229);
and U1424 (N_1424,In_427,In_2751);
nor U1425 (N_1425,In_2274,In_333);
nand U1426 (N_1426,In_1112,In_133);
xnor U1427 (N_1427,In_2648,In_1233);
xnor U1428 (N_1428,In_2690,In_2134);
or U1429 (N_1429,In_830,In_2222);
and U1430 (N_1430,In_0,In_1001);
nor U1431 (N_1431,In_2783,In_2461);
and U1432 (N_1432,In_2865,In_2336);
and U1433 (N_1433,In_23,In_2702);
nand U1434 (N_1434,In_227,In_2245);
nor U1435 (N_1435,In_1987,In_1563);
xor U1436 (N_1436,In_2199,In_1789);
and U1437 (N_1437,In_2847,In_971);
or U1438 (N_1438,In_525,In_1897);
nor U1439 (N_1439,In_564,In_1844);
xnor U1440 (N_1440,In_956,In_560);
and U1441 (N_1441,In_1800,In_1873);
nand U1442 (N_1442,In_1551,In_2770);
and U1443 (N_1443,In_2767,In_1902);
and U1444 (N_1444,In_2613,In_2248);
nor U1445 (N_1445,In_2006,In_314);
nand U1446 (N_1446,In_1568,In_1794);
and U1447 (N_1447,In_2406,In_379);
xor U1448 (N_1448,In_1512,In_2612);
or U1449 (N_1449,In_1682,In_1881);
nand U1450 (N_1450,In_1660,In_1819);
and U1451 (N_1451,In_1533,In_2125);
and U1452 (N_1452,In_1662,In_803);
xor U1453 (N_1453,In_2341,In_151);
and U1454 (N_1454,In_1454,In_657);
and U1455 (N_1455,In_2630,In_516);
nor U1456 (N_1456,In_2467,In_1814);
or U1457 (N_1457,In_1920,In_330);
or U1458 (N_1458,In_995,In_111);
xor U1459 (N_1459,In_661,In_1617);
nand U1460 (N_1460,In_466,In_130);
and U1461 (N_1461,In_315,In_1511);
and U1462 (N_1462,In_2092,In_1931);
and U1463 (N_1463,In_1421,In_2915);
or U1464 (N_1464,In_2119,In_311);
nor U1465 (N_1465,In_778,In_20);
and U1466 (N_1466,In_2709,In_2792);
nor U1467 (N_1467,In_2372,In_1621);
and U1468 (N_1468,In_1965,In_554);
nor U1469 (N_1469,In_2859,In_1236);
or U1470 (N_1470,In_2573,In_320);
and U1471 (N_1471,In_2432,In_1735);
nor U1472 (N_1472,In_1248,In_1440);
and U1473 (N_1473,In_129,In_675);
nor U1474 (N_1474,In_2145,In_2079);
and U1475 (N_1475,In_1521,In_1302);
and U1476 (N_1476,In_1874,In_1937);
nand U1477 (N_1477,In_1959,In_1144);
nand U1478 (N_1478,In_2538,In_1418);
and U1479 (N_1479,In_1625,In_2587);
xor U1480 (N_1480,In_2149,In_1879);
xnor U1481 (N_1481,In_687,In_254);
xnor U1482 (N_1482,In_570,In_863);
xnor U1483 (N_1483,In_2430,In_2322);
nand U1484 (N_1484,In_2695,In_1887);
and U1485 (N_1485,In_2550,In_1134);
xor U1486 (N_1486,In_295,In_1167);
nor U1487 (N_1487,In_1684,In_207);
xor U1488 (N_1488,In_1522,In_1754);
nand U1489 (N_1489,In_948,In_1314);
xor U1490 (N_1490,In_2804,In_51);
or U1491 (N_1491,In_56,In_643);
or U1492 (N_1492,In_1847,In_2446);
and U1493 (N_1493,In_1501,In_2641);
xor U1494 (N_1494,In_2147,In_464);
or U1495 (N_1495,In_970,In_2945);
or U1496 (N_1496,In_2228,In_2217);
nor U1497 (N_1497,In_2754,In_1229);
nor U1498 (N_1498,In_2717,In_602);
nand U1499 (N_1499,In_1648,In_78);
and U1500 (N_1500,In_336,In_2349);
nand U1501 (N_1501,In_566,In_1830);
xor U1502 (N_1502,In_47,In_2399);
and U1503 (N_1503,In_2835,In_2562);
and U1504 (N_1504,In_1373,In_611);
xor U1505 (N_1505,In_2799,In_493);
or U1506 (N_1506,In_1920,In_941);
and U1507 (N_1507,In_2833,In_1068);
and U1508 (N_1508,In_1825,In_2835);
and U1509 (N_1509,In_682,In_267);
xor U1510 (N_1510,In_2490,In_1330);
xor U1511 (N_1511,In_481,In_2371);
nand U1512 (N_1512,In_2706,In_1538);
nor U1513 (N_1513,In_2070,In_952);
nand U1514 (N_1514,In_980,In_2560);
nor U1515 (N_1515,In_704,In_81);
or U1516 (N_1516,In_109,In_394);
xor U1517 (N_1517,In_1899,In_1274);
or U1518 (N_1518,In_1430,In_2938);
xor U1519 (N_1519,In_482,In_916);
nor U1520 (N_1520,In_558,In_185);
xnor U1521 (N_1521,In_2882,In_2588);
and U1522 (N_1522,In_1259,In_2000);
nor U1523 (N_1523,In_2063,In_2594);
xnor U1524 (N_1524,In_2793,In_2449);
nor U1525 (N_1525,In_1234,In_511);
nand U1526 (N_1526,In_60,In_746);
and U1527 (N_1527,In_1107,In_812);
nand U1528 (N_1528,In_531,In_2528);
and U1529 (N_1529,In_460,In_1858);
xor U1530 (N_1530,In_1083,In_1501);
xor U1531 (N_1531,In_1919,In_2681);
and U1532 (N_1532,In_1900,In_1785);
nor U1533 (N_1533,In_1970,In_717);
nor U1534 (N_1534,In_2768,In_806);
nand U1535 (N_1535,In_622,In_1390);
nand U1536 (N_1536,In_2718,In_2457);
xor U1537 (N_1537,In_2367,In_1236);
nand U1538 (N_1538,In_1291,In_2547);
and U1539 (N_1539,In_2119,In_1414);
xnor U1540 (N_1540,In_633,In_853);
xnor U1541 (N_1541,In_783,In_529);
or U1542 (N_1542,In_2864,In_1696);
and U1543 (N_1543,In_931,In_2087);
nand U1544 (N_1544,In_934,In_2815);
or U1545 (N_1545,In_2499,In_2177);
or U1546 (N_1546,In_2703,In_2009);
nor U1547 (N_1547,In_2648,In_402);
nand U1548 (N_1548,In_434,In_2182);
or U1549 (N_1549,In_2972,In_1442);
and U1550 (N_1550,In_668,In_958);
or U1551 (N_1551,In_1297,In_1745);
xor U1552 (N_1552,In_1346,In_1985);
and U1553 (N_1553,In_852,In_2999);
nand U1554 (N_1554,In_632,In_2319);
and U1555 (N_1555,In_2827,In_1573);
and U1556 (N_1556,In_1836,In_2038);
and U1557 (N_1557,In_812,In_1599);
and U1558 (N_1558,In_1127,In_1746);
nand U1559 (N_1559,In_2390,In_2321);
xor U1560 (N_1560,In_1257,In_2610);
nor U1561 (N_1561,In_2807,In_1199);
nand U1562 (N_1562,In_658,In_229);
nand U1563 (N_1563,In_2843,In_2391);
nor U1564 (N_1564,In_2692,In_2249);
and U1565 (N_1565,In_2275,In_1585);
or U1566 (N_1566,In_2206,In_225);
and U1567 (N_1567,In_2969,In_1064);
xor U1568 (N_1568,In_1324,In_2413);
xnor U1569 (N_1569,In_1312,In_858);
nor U1570 (N_1570,In_228,In_168);
nor U1571 (N_1571,In_587,In_1263);
or U1572 (N_1572,In_1892,In_294);
and U1573 (N_1573,In_1427,In_1488);
and U1574 (N_1574,In_1823,In_2343);
nor U1575 (N_1575,In_934,In_1546);
and U1576 (N_1576,In_2592,In_1639);
nand U1577 (N_1577,In_453,In_2409);
nor U1578 (N_1578,In_1650,In_1660);
or U1579 (N_1579,In_831,In_913);
or U1580 (N_1580,In_1321,In_2819);
and U1581 (N_1581,In_824,In_1512);
and U1582 (N_1582,In_614,In_2676);
and U1583 (N_1583,In_1808,In_1061);
nor U1584 (N_1584,In_2912,In_1512);
nand U1585 (N_1585,In_1167,In_2916);
nand U1586 (N_1586,In_2034,In_2168);
xnor U1587 (N_1587,In_2817,In_2825);
or U1588 (N_1588,In_2632,In_2364);
nor U1589 (N_1589,In_2473,In_722);
xor U1590 (N_1590,In_1481,In_1221);
xnor U1591 (N_1591,In_2681,In_2742);
xnor U1592 (N_1592,In_1984,In_108);
or U1593 (N_1593,In_1376,In_2960);
and U1594 (N_1594,In_1861,In_762);
or U1595 (N_1595,In_2412,In_1853);
nand U1596 (N_1596,In_296,In_1082);
nor U1597 (N_1597,In_2845,In_2713);
or U1598 (N_1598,In_1501,In_711);
or U1599 (N_1599,In_2645,In_458);
nor U1600 (N_1600,In_1213,In_1357);
nand U1601 (N_1601,In_721,In_2987);
or U1602 (N_1602,In_2531,In_1958);
and U1603 (N_1603,In_2949,In_1827);
xnor U1604 (N_1604,In_581,In_2134);
and U1605 (N_1605,In_2178,In_1208);
nand U1606 (N_1606,In_2270,In_202);
nand U1607 (N_1607,In_2966,In_2014);
nand U1608 (N_1608,In_93,In_2585);
or U1609 (N_1609,In_329,In_13);
and U1610 (N_1610,In_1579,In_2954);
xnor U1611 (N_1611,In_1560,In_1996);
nor U1612 (N_1612,In_185,In_886);
xnor U1613 (N_1613,In_1630,In_1261);
nor U1614 (N_1614,In_2623,In_640);
nand U1615 (N_1615,In_27,In_810);
nand U1616 (N_1616,In_1422,In_2641);
and U1617 (N_1617,In_628,In_787);
nand U1618 (N_1618,In_2074,In_2018);
nand U1619 (N_1619,In_2596,In_536);
nand U1620 (N_1620,In_1431,In_1793);
and U1621 (N_1621,In_2199,In_2771);
nor U1622 (N_1622,In_1712,In_405);
or U1623 (N_1623,In_457,In_1009);
and U1624 (N_1624,In_1312,In_950);
xnor U1625 (N_1625,In_2700,In_1541);
nor U1626 (N_1626,In_1110,In_1379);
and U1627 (N_1627,In_2834,In_472);
and U1628 (N_1628,In_1076,In_2110);
or U1629 (N_1629,In_1767,In_932);
or U1630 (N_1630,In_1494,In_1859);
or U1631 (N_1631,In_2645,In_26);
nand U1632 (N_1632,In_1024,In_139);
or U1633 (N_1633,In_716,In_2474);
or U1634 (N_1634,In_2601,In_1914);
nor U1635 (N_1635,In_1002,In_1281);
nand U1636 (N_1636,In_2744,In_1166);
xnor U1637 (N_1637,In_2766,In_1219);
nor U1638 (N_1638,In_321,In_887);
nor U1639 (N_1639,In_2425,In_996);
xor U1640 (N_1640,In_1087,In_2537);
nor U1641 (N_1641,In_1385,In_2015);
nand U1642 (N_1642,In_986,In_2655);
or U1643 (N_1643,In_2618,In_1695);
or U1644 (N_1644,In_2294,In_1983);
and U1645 (N_1645,In_1069,In_166);
or U1646 (N_1646,In_2660,In_2047);
or U1647 (N_1647,In_947,In_1892);
nand U1648 (N_1648,In_1624,In_457);
and U1649 (N_1649,In_2205,In_555);
nand U1650 (N_1650,In_264,In_1531);
nand U1651 (N_1651,In_1559,In_1593);
or U1652 (N_1652,In_2781,In_2130);
nor U1653 (N_1653,In_1968,In_1236);
or U1654 (N_1654,In_1841,In_2711);
and U1655 (N_1655,In_2195,In_2441);
xnor U1656 (N_1656,In_1677,In_1409);
or U1657 (N_1657,In_1364,In_2709);
nor U1658 (N_1658,In_753,In_1537);
and U1659 (N_1659,In_2988,In_1690);
xnor U1660 (N_1660,In_1828,In_154);
and U1661 (N_1661,In_848,In_59);
nor U1662 (N_1662,In_1762,In_2125);
or U1663 (N_1663,In_1562,In_1316);
nor U1664 (N_1664,In_2482,In_394);
nand U1665 (N_1665,In_2818,In_832);
nand U1666 (N_1666,In_2495,In_1389);
xnor U1667 (N_1667,In_1435,In_279);
or U1668 (N_1668,In_448,In_723);
xnor U1669 (N_1669,In_2369,In_198);
xnor U1670 (N_1670,In_893,In_2744);
or U1671 (N_1671,In_2180,In_2959);
nand U1672 (N_1672,In_188,In_530);
and U1673 (N_1673,In_415,In_2019);
and U1674 (N_1674,In_1127,In_2623);
nand U1675 (N_1675,In_1803,In_942);
nor U1676 (N_1676,In_1793,In_624);
nand U1677 (N_1677,In_1353,In_1797);
nand U1678 (N_1678,In_2944,In_2977);
and U1679 (N_1679,In_1513,In_1517);
nor U1680 (N_1680,In_1375,In_1612);
xor U1681 (N_1681,In_894,In_1545);
nand U1682 (N_1682,In_2098,In_1851);
nand U1683 (N_1683,In_1292,In_2203);
xor U1684 (N_1684,In_471,In_962);
or U1685 (N_1685,In_1664,In_1446);
xnor U1686 (N_1686,In_1365,In_2065);
or U1687 (N_1687,In_2066,In_580);
xnor U1688 (N_1688,In_491,In_2934);
or U1689 (N_1689,In_2587,In_731);
xor U1690 (N_1690,In_1145,In_2011);
or U1691 (N_1691,In_1064,In_1918);
or U1692 (N_1692,In_1550,In_1376);
nor U1693 (N_1693,In_534,In_2311);
nand U1694 (N_1694,In_1069,In_1274);
or U1695 (N_1695,In_2674,In_2756);
or U1696 (N_1696,In_2993,In_2376);
nand U1697 (N_1697,In_790,In_1377);
or U1698 (N_1698,In_2577,In_2723);
xnor U1699 (N_1699,In_2433,In_1435);
xnor U1700 (N_1700,In_82,In_2901);
nand U1701 (N_1701,In_1456,In_114);
or U1702 (N_1702,In_1655,In_786);
and U1703 (N_1703,In_355,In_1924);
or U1704 (N_1704,In_2056,In_771);
and U1705 (N_1705,In_2367,In_2987);
nand U1706 (N_1706,In_498,In_1655);
nand U1707 (N_1707,In_852,In_2516);
and U1708 (N_1708,In_1881,In_2090);
and U1709 (N_1709,In_2911,In_2400);
nor U1710 (N_1710,In_1212,In_1531);
and U1711 (N_1711,In_231,In_670);
xnor U1712 (N_1712,In_286,In_2000);
nor U1713 (N_1713,In_2250,In_2667);
xor U1714 (N_1714,In_2797,In_550);
xor U1715 (N_1715,In_436,In_615);
and U1716 (N_1716,In_1380,In_688);
or U1717 (N_1717,In_2971,In_2644);
xnor U1718 (N_1718,In_1284,In_2712);
and U1719 (N_1719,In_973,In_357);
nand U1720 (N_1720,In_1742,In_450);
or U1721 (N_1721,In_1573,In_1522);
xor U1722 (N_1722,In_720,In_871);
and U1723 (N_1723,In_1130,In_2439);
nor U1724 (N_1724,In_1605,In_2689);
nand U1725 (N_1725,In_506,In_354);
nand U1726 (N_1726,In_2224,In_1150);
and U1727 (N_1727,In_2545,In_1022);
and U1728 (N_1728,In_2650,In_443);
nor U1729 (N_1729,In_2430,In_320);
nor U1730 (N_1730,In_1346,In_903);
xnor U1731 (N_1731,In_180,In_2739);
or U1732 (N_1732,In_2209,In_912);
nor U1733 (N_1733,In_2476,In_2423);
xor U1734 (N_1734,In_1343,In_2333);
or U1735 (N_1735,In_2214,In_1122);
nand U1736 (N_1736,In_2462,In_650);
or U1737 (N_1737,In_552,In_1505);
or U1738 (N_1738,In_1369,In_988);
and U1739 (N_1739,In_2252,In_651);
nand U1740 (N_1740,In_442,In_266);
nor U1741 (N_1741,In_1041,In_1604);
or U1742 (N_1742,In_1937,In_905);
nand U1743 (N_1743,In_467,In_1161);
nand U1744 (N_1744,In_199,In_318);
nor U1745 (N_1745,In_848,In_2441);
xor U1746 (N_1746,In_658,In_795);
nor U1747 (N_1747,In_1095,In_1280);
or U1748 (N_1748,In_882,In_2785);
nand U1749 (N_1749,In_1,In_2407);
or U1750 (N_1750,In_2963,In_217);
nor U1751 (N_1751,In_1527,In_2697);
or U1752 (N_1752,In_410,In_1611);
and U1753 (N_1753,In_2507,In_2234);
nor U1754 (N_1754,In_500,In_2220);
and U1755 (N_1755,In_2506,In_770);
nor U1756 (N_1756,In_1641,In_2706);
nor U1757 (N_1757,In_1259,In_487);
and U1758 (N_1758,In_335,In_245);
xor U1759 (N_1759,In_2667,In_2189);
or U1760 (N_1760,In_1618,In_461);
and U1761 (N_1761,In_2532,In_1755);
nand U1762 (N_1762,In_1345,In_612);
or U1763 (N_1763,In_2925,In_2806);
xnor U1764 (N_1764,In_976,In_545);
xnor U1765 (N_1765,In_556,In_677);
nand U1766 (N_1766,In_958,In_1731);
xor U1767 (N_1767,In_1696,In_2056);
nor U1768 (N_1768,In_2973,In_1344);
nor U1769 (N_1769,In_2426,In_255);
xor U1770 (N_1770,In_1818,In_231);
nand U1771 (N_1771,In_341,In_535);
or U1772 (N_1772,In_1680,In_2858);
xnor U1773 (N_1773,In_1168,In_275);
or U1774 (N_1774,In_1614,In_493);
nand U1775 (N_1775,In_1200,In_1278);
xor U1776 (N_1776,In_359,In_700);
nor U1777 (N_1777,In_1846,In_381);
nand U1778 (N_1778,In_166,In_2860);
nor U1779 (N_1779,In_2486,In_2009);
nor U1780 (N_1780,In_1154,In_551);
and U1781 (N_1781,In_131,In_1357);
or U1782 (N_1782,In_1489,In_2189);
and U1783 (N_1783,In_955,In_1469);
and U1784 (N_1784,In_2498,In_672);
nor U1785 (N_1785,In_2582,In_1653);
nor U1786 (N_1786,In_822,In_2516);
nor U1787 (N_1787,In_155,In_294);
and U1788 (N_1788,In_973,In_2036);
nand U1789 (N_1789,In_1055,In_258);
nor U1790 (N_1790,In_1437,In_1273);
nand U1791 (N_1791,In_1915,In_212);
or U1792 (N_1792,In_2628,In_1232);
or U1793 (N_1793,In_1639,In_609);
nor U1794 (N_1794,In_2553,In_1534);
xor U1795 (N_1795,In_1660,In_2454);
nand U1796 (N_1796,In_1302,In_2413);
and U1797 (N_1797,In_1704,In_1716);
and U1798 (N_1798,In_1374,In_1479);
xor U1799 (N_1799,In_230,In_2126);
xor U1800 (N_1800,In_522,In_1219);
xnor U1801 (N_1801,In_1853,In_2098);
or U1802 (N_1802,In_922,In_2092);
xnor U1803 (N_1803,In_1625,In_334);
nand U1804 (N_1804,In_1598,In_838);
and U1805 (N_1805,In_2804,In_2981);
nor U1806 (N_1806,In_650,In_2726);
and U1807 (N_1807,In_25,In_1179);
and U1808 (N_1808,In_2563,In_641);
nand U1809 (N_1809,In_2564,In_1385);
or U1810 (N_1810,In_468,In_249);
xnor U1811 (N_1811,In_2116,In_142);
or U1812 (N_1812,In_1145,In_2996);
xor U1813 (N_1813,In_1391,In_1776);
and U1814 (N_1814,In_1521,In_566);
nor U1815 (N_1815,In_893,In_717);
nor U1816 (N_1816,In_1808,In_2392);
or U1817 (N_1817,In_929,In_1392);
nand U1818 (N_1818,In_2448,In_1365);
nor U1819 (N_1819,In_915,In_267);
and U1820 (N_1820,In_2836,In_2652);
nand U1821 (N_1821,In_2420,In_324);
and U1822 (N_1822,In_2064,In_1020);
and U1823 (N_1823,In_184,In_2087);
nor U1824 (N_1824,In_1306,In_216);
or U1825 (N_1825,In_2164,In_1259);
nand U1826 (N_1826,In_2611,In_2365);
nor U1827 (N_1827,In_1507,In_466);
xnor U1828 (N_1828,In_258,In_1874);
or U1829 (N_1829,In_42,In_1321);
or U1830 (N_1830,In_940,In_136);
xor U1831 (N_1831,In_2557,In_2325);
nand U1832 (N_1832,In_1206,In_2141);
nand U1833 (N_1833,In_2123,In_1360);
nand U1834 (N_1834,In_367,In_1256);
and U1835 (N_1835,In_1679,In_1523);
nand U1836 (N_1836,In_2900,In_1675);
nand U1837 (N_1837,In_2085,In_985);
nor U1838 (N_1838,In_2722,In_1796);
and U1839 (N_1839,In_618,In_1335);
or U1840 (N_1840,In_2856,In_1925);
nand U1841 (N_1841,In_1573,In_2378);
nor U1842 (N_1842,In_2441,In_2989);
nand U1843 (N_1843,In_2709,In_1974);
or U1844 (N_1844,In_1813,In_279);
xor U1845 (N_1845,In_1436,In_1383);
or U1846 (N_1846,In_1830,In_1113);
xnor U1847 (N_1847,In_1628,In_878);
or U1848 (N_1848,In_2927,In_297);
nand U1849 (N_1849,In_2930,In_2593);
or U1850 (N_1850,In_2439,In_2001);
xor U1851 (N_1851,In_2724,In_1685);
xor U1852 (N_1852,In_552,In_1885);
and U1853 (N_1853,In_2873,In_957);
and U1854 (N_1854,In_652,In_2941);
nor U1855 (N_1855,In_996,In_2050);
nor U1856 (N_1856,In_2980,In_2851);
xnor U1857 (N_1857,In_2395,In_1412);
nand U1858 (N_1858,In_2964,In_640);
and U1859 (N_1859,In_1245,In_1079);
nand U1860 (N_1860,In_1144,In_2149);
nor U1861 (N_1861,In_1375,In_468);
nor U1862 (N_1862,In_1117,In_2398);
nor U1863 (N_1863,In_789,In_2884);
and U1864 (N_1864,In_2532,In_59);
or U1865 (N_1865,In_560,In_1857);
nor U1866 (N_1866,In_2262,In_1993);
xnor U1867 (N_1867,In_2930,In_572);
nor U1868 (N_1868,In_326,In_1909);
and U1869 (N_1869,In_1455,In_1669);
and U1870 (N_1870,In_2472,In_1747);
and U1871 (N_1871,In_2001,In_76);
xnor U1872 (N_1872,In_1020,In_2708);
xor U1873 (N_1873,In_981,In_2465);
xnor U1874 (N_1874,In_2989,In_393);
xnor U1875 (N_1875,In_1742,In_2594);
and U1876 (N_1876,In_2660,In_191);
or U1877 (N_1877,In_1583,In_655);
nor U1878 (N_1878,In_376,In_829);
nor U1879 (N_1879,In_2494,In_263);
xnor U1880 (N_1880,In_2023,In_855);
and U1881 (N_1881,In_1817,In_2045);
or U1882 (N_1882,In_1767,In_2760);
xor U1883 (N_1883,In_2032,In_2687);
and U1884 (N_1884,In_111,In_603);
nor U1885 (N_1885,In_1938,In_2043);
or U1886 (N_1886,In_2430,In_1701);
xnor U1887 (N_1887,In_2245,In_570);
xnor U1888 (N_1888,In_2725,In_2072);
xor U1889 (N_1889,In_1324,In_2524);
or U1890 (N_1890,In_1120,In_1735);
nor U1891 (N_1891,In_1436,In_2485);
or U1892 (N_1892,In_2874,In_2308);
and U1893 (N_1893,In_622,In_2208);
or U1894 (N_1894,In_2143,In_374);
or U1895 (N_1895,In_87,In_1260);
nand U1896 (N_1896,In_1763,In_2313);
nand U1897 (N_1897,In_2942,In_400);
and U1898 (N_1898,In_263,In_2613);
xnor U1899 (N_1899,In_2224,In_521);
nand U1900 (N_1900,In_2208,In_810);
nand U1901 (N_1901,In_2742,In_349);
or U1902 (N_1902,In_524,In_2142);
nor U1903 (N_1903,In_1967,In_408);
and U1904 (N_1904,In_1055,In_744);
and U1905 (N_1905,In_2790,In_1641);
nand U1906 (N_1906,In_2692,In_2459);
nor U1907 (N_1907,In_1540,In_362);
xnor U1908 (N_1908,In_1944,In_1116);
and U1909 (N_1909,In_2524,In_902);
nand U1910 (N_1910,In_1813,In_1124);
xnor U1911 (N_1911,In_47,In_777);
and U1912 (N_1912,In_1765,In_257);
nor U1913 (N_1913,In_2064,In_2725);
nor U1914 (N_1914,In_492,In_2682);
nand U1915 (N_1915,In_1098,In_1261);
or U1916 (N_1916,In_322,In_2586);
xor U1917 (N_1917,In_399,In_2857);
nor U1918 (N_1918,In_2074,In_1998);
nand U1919 (N_1919,In_539,In_2391);
and U1920 (N_1920,In_1881,In_785);
nor U1921 (N_1921,In_667,In_116);
nor U1922 (N_1922,In_2956,In_173);
and U1923 (N_1923,In_2645,In_121);
nor U1924 (N_1924,In_2962,In_2504);
xnor U1925 (N_1925,In_1472,In_1145);
xnor U1926 (N_1926,In_932,In_1062);
or U1927 (N_1927,In_1677,In_1888);
xor U1928 (N_1928,In_2196,In_22);
nand U1929 (N_1929,In_1711,In_500);
nor U1930 (N_1930,In_13,In_817);
xnor U1931 (N_1931,In_2903,In_536);
or U1932 (N_1932,In_862,In_231);
xor U1933 (N_1933,In_497,In_1684);
xnor U1934 (N_1934,In_468,In_371);
or U1935 (N_1935,In_660,In_2232);
or U1936 (N_1936,In_1938,In_2418);
or U1937 (N_1937,In_1452,In_2879);
nand U1938 (N_1938,In_216,In_811);
and U1939 (N_1939,In_26,In_1168);
xnor U1940 (N_1940,In_1399,In_17);
nor U1941 (N_1941,In_2793,In_339);
nor U1942 (N_1942,In_294,In_887);
nand U1943 (N_1943,In_2230,In_385);
xor U1944 (N_1944,In_2364,In_1492);
or U1945 (N_1945,In_2253,In_2891);
xor U1946 (N_1946,In_579,In_1014);
nand U1947 (N_1947,In_2621,In_1299);
nor U1948 (N_1948,In_503,In_743);
and U1949 (N_1949,In_383,In_1858);
nand U1950 (N_1950,In_869,In_201);
and U1951 (N_1951,In_2334,In_1246);
nor U1952 (N_1952,In_2382,In_785);
and U1953 (N_1953,In_2898,In_1099);
or U1954 (N_1954,In_2691,In_2145);
and U1955 (N_1955,In_2064,In_1405);
nor U1956 (N_1956,In_2850,In_1939);
nand U1957 (N_1957,In_942,In_933);
or U1958 (N_1958,In_606,In_2267);
nor U1959 (N_1959,In_202,In_442);
or U1960 (N_1960,In_929,In_1966);
nor U1961 (N_1961,In_66,In_734);
or U1962 (N_1962,In_1053,In_2010);
or U1963 (N_1963,In_1756,In_2635);
nor U1964 (N_1964,In_693,In_1995);
nand U1965 (N_1965,In_1014,In_262);
nand U1966 (N_1966,In_1283,In_96);
xnor U1967 (N_1967,In_2050,In_2766);
nor U1968 (N_1968,In_436,In_1278);
nand U1969 (N_1969,In_951,In_2499);
nor U1970 (N_1970,In_1386,In_521);
or U1971 (N_1971,In_242,In_2191);
and U1972 (N_1972,In_2047,In_2455);
xnor U1973 (N_1973,In_99,In_969);
nor U1974 (N_1974,In_1683,In_1900);
or U1975 (N_1975,In_1150,In_2101);
and U1976 (N_1976,In_2698,In_2302);
and U1977 (N_1977,In_515,In_1933);
nor U1978 (N_1978,In_2500,In_1553);
xnor U1979 (N_1979,In_1295,In_217);
or U1980 (N_1980,In_994,In_655);
xor U1981 (N_1981,In_849,In_2411);
xor U1982 (N_1982,In_1786,In_1243);
xor U1983 (N_1983,In_1077,In_2485);
xnor U1984 (N_1984,In_2239,In_1860);
xor U1985 (N_1985,In_1913,In_729);
nand U1986 (N_1986,In_1287,In_1582);
nor U1987 (N_1987,In_495,In_1608);
and U1988 (N_1988,In_1441,In_2018);
nand U1989 (N_1989,In_836,In_2256);
nor U1990 (N_1990,In_589,In_2808);
and U1991 (N_1991,In_374,In_2940);
and U1992 (N_1992,In_807,In_2146);
nand U1993 (N_1993,In_2180,In_2280);
nand U1994 (N_1994,In_2255,In_1493);
or U1995 (N_1995,In_565,In_1454);
nor U1996 (N_1996,In_1203,In_1438);
and U1997 (N_1997,In_1531,In_1508);
nor U1998 (N_1998,In_1524,In_1970);
or U1999 (N_1999,In_1448,In_440);
xor U2000 (N_2000,N_1401,N_1148);
and U2001 (N_2001,N_1963,N_131);
xnor U2002 (N_2002,N_970,N_202);
nand U2003 (N_2003,N_1600,N_723);
nand U2004 (N_2004,N_60,N_1270);
nor U2005 (N_2005,N_956,N_1491);
nand U2006 (N_2006,N_656,N_688);
and U2007 (N_2007,N_941,N_222);
nor U2008 (N_2008,N_7,N_242);
nand U2009 (N_2009,N_1102,N_1828);
xor U2010 (N_2010,N_159,N_1510);
or U2011 (N_2011,N_254,N_573);
nor U2012 (N_2012,N_1895,N_71);
xor U2013 (N_2013,N_862,N_179);
nor U2014 (N_2014,N_973,N_170);
or U2015 (N_2015,N_874,N_1788);
or U2016 (N_2016,N_1745,N_745);
nand U2017 (N_2017,N_1168,N_1883);
nor U2018 (N_2018,N_1040,N_1667);
and U2019 (N_2019,N_1243,N_67);
nand U2020 (N_2020,N_712,N_258);
nand U2021 (N_2021,N_905,N_598);
and U2022 (N_2022,N_1646,N_857);
xor U2023 (N_2023,N_1096,N_334);
nor U2024 (N_2024,N_111,N_284);
nand U2025 (N_2025,N_1022,N_1088);
xor U2026 (N_2026,N_1409,N_31);
xor U2027 (N_2027,N_462,N_1124);
xor U2028 (N_2028,N_1501,N_313);
nor U2029 (N_2029,N_136,N_1271);
and U2030 (N_2030,N_1651,N_1793);
nand U2031 (N_2031,N_383,N_20);
or U2032 (N_2032,N_1568,N_1245);
or U2033 (N_2033,N_609,N_1875);
nand U2034 (N_2034,N_1388,N_1311);
or U2035 (N_2035,N_515,N_901);
xnor U2036 (N_2036,N_1251,N_1371);
nor U2037 (N_2037,N_225,N_110);
or U2038 (N_2038,N_1261,N_25);
nor U2039 (N_2039,N_1320,N_356);
nand U2040 (N_2040,N_483,N_1855);
nand U2041 (N_2041,N_1654,N_747);
nand U2042 (N_2042,N_848,N_363);
or U2043 (N_2043,N_909,N_1464);
nand U2044 (N_2044,N_1601,N_1304);
and U2045 (N_2045,N_387,N_156);
nand U2046 (N_2046,N_154,N_1700);
or U2047 (N_2047,N_1607,N_1581);
or U2048 (N_2048,N_1323,N_58);
and U2049 (N_2049,N_397,N_1871);
nand U2050 (N_2050,N_499,N_1685);
nand U2051 (N_2051,N_1310,N_1649);
nand U2052 (N_2052,N_101,N_1236);
and U2053 (N_2053,N_1241,N_1122);
nor U2054 (N_2054,N_168,N_1321);
or U2055 (N_2055,N_837,N_1385);
xnor U2056 (N_2056,N_793,N_1201);
or U2057 (N_2057,N_748,N_514);
xor U2058 (N_2058,N_288,N_1092);
nor U2059 (N_2059,N_1199,N_1132);
xnor U2060 (N_2060,N_1114,N_1493);
and U2061 (N_2061,N_1127,N_1695);
xnor U2062 (N_2062,N_1852,N_833);
or U2063 (N_2063,N_261,N_41);
or U2064 (N_2064,N_991,N_1711);
and U2065 (N_2065,N_1768,N_1712);
nor U2066 (N_2066,N_923,N_472);
nand U2067 (N_2067,N_791,N_4);
xor U2068 (N_2068,N_1880,N_321);
xnor U2069 (N_2069,N_68,N_1773);
and U2070 (N_2070,N_1566,N_1790);
and U2071 (N_2071,N_1746,N_722);
xnor U2072 (N_2072,N_1334,N_425);
or U2073 (N_2073,N_1373,N_38);
xnor U2074 (N_2074,N_892,N_1670);
nand U2075 (N_2075,N_986,N_177);
nor U2076 (N_2076,N_1424,N_1546);
nor U2077 (N_2077,N_819,N_1597);
xor U2078 (N_2078,N_730,N_593);
nor U2079 (N_2079,N_1561,N_616);
and U2080 (N_2080,N_1846,N_437);
and U2081 (N_2081,N_81,N_1342);
and U2082 (N_2082,N_1503,N_91);
nand U2083 (N_2083,N_689,N_1351);
xnor U2084 (N_2084,N_1544,N_559);
nor U2085 (N_2085,N_1553,N_965);
xnor U2086 (N_2086,N_1337,N_871);
and U2087 (N_2087,N_1387,N_705);
or U2088 (N_2088,N_1262,N_1499);
nor U2089 (N_2089,N_384,N_1489);
xor U2090 (N_2090,N_858,N_600);
and U2091 (N_2091,N_1580,N_660);
nand U2092 (N_2092,N_1984,N_153);
and U2093 (N_2093,N_1346,N_196);
nor U2094 (N_2094,N_714,N_280);
xnor U2095 (N_2095,N_860,N_434);
nor U2096 (N_2096,N_1329,N_1397);
nand U2097 (N_2097,N_999,N_1297);
nand U2098 (N_2098,N_1727,N_1569);
and U2099 (N_2099,N_644,N_916);
or U2100 (N_2100,N_266,N_30);
and U2101 (N_2101,N_324,N_808);
nor U2102 (N_2102,N_33,N_729);
nand U2103 (N_2103,N_1172,N_1827);
nand U2104 (N_2104,N_1956,N_1823);
nor U2105 (N_2105,N_1953,N_1454);
or U2106 (N_2106,N_1490,N_846);
nor U2107 (N_2107,N_1964,N_863);
nor U2108 (N_2108,N_9,N_134);
xor U2109 (N_2109,N_1706,N_255);
nor U2110 (N_2110,N_1624,N_840);
nor U2111 (N_2111,N_35,N_40);
or U2112 (N_2112,N_1997,N_538);
nand U2113 (N_2113,N_1308,N_1998);
nand U2114 (N_2114,N_693,N_1770);
and U2115 (N_2115,N_116,N_560);
xnor U2116 (N_2116,N_140,N_1690);
nand U2117 (N_2117,N_454,N_706);
nand U2118 (N_2118,N_129,N_1925);
nand U2119 (N_2119,N_798,N_1878);
nor U2120 (N_2120,N_763,N_1748);
nand U2121 (N_2121,N_1940,N_1713);
nand U2122 (N_2122,N_1897,N_754);
or U2123 (N_2123,N_1158,N_1989);
and U2124 (N_2124,N_1350,N_1724);
nor U2125 (N_2125,N_1567,N_409);
nand U2126 (N_2126,N_251,N_964);
nand U2127 (N_2127,N_1459,N_1630);
nand U2128 (N_2128,N_1604,N_709);
nand U2129 (N_2129,N_172,N_1742);
xnor U2130 (N_2130,N_954,N_346);
xnor U2131 (N_2131,N_369,N_1888);
nor U2132 (N_2132,N_1405,N_317);
xnor U2133 (N_2133,N_496,N_1287);
nor U2134 (N_2134,N_733,N_199);
nand U2135 (N_2135,N_413,N_420);
and U2136 (N_2136,N_180,N_1286);
or U2137 (N_2137,N_966,N_1634);
nor U2138 (N_2138,N_175,N_1867);
nand U2139 (N_2139,N_539,N_930);
xnor U2140 (N_2140,N_928,N_1596);
nor U2141 (N_2141,N_882,N_1162);
nor U2142 (N_2142,N_1171,N_200);
nand U2143 (N_2143,N_680,N_904);
nor U2144 (N_2144,N_137,N_1256);
nor U2145 (N_2145,N_993,N_1502);
xnor U2146 (N_2146,N_1228,N_711);
or U2147 (N_2147,N_792,N_193);
xor U2148 (N_2148,N_888,N_1259);
nor U2149 (N_2149,N_1368,N_554);
or U2150 (N_2150,N_1315,N_1717);
or U2151 (N_2151,N_1534,N_699);
or U2152 (N_2152,N_16,N_1097);
nand U2153 (N_2153,N_1240,N_1804);
xnor U2154 (N_2154,N_1402,N_341);
nor U2155 (N_2155,N_1660,N_1086);
and U2156 (N_2156,N_1066,N_147);
nand U2157 (N_2157,N_1794,N_1856);
or U2158 (N_2158,N_329,N_1862);
nor U2159 (N_2159,N_152,N_1353);
nand U2160 (N_2160,N_1431,N_374);
nand U2161 (N_2161,N_365,N_290);
xor U2162 (N_2162,N_1492,N_1186);
nor U2163 (N_2163,N_1811,N_273);
xor U2164 (N_2164,N_155,N_239);
nand U2165 (N_2165,N_234,N_957);
xnor U2166 (N_2166,N_1861,N_1539);
nand U2167 (N_2167,N_781,N_415);
nor U2168 (N_2168,N_1520,N_1303);
or U2169 (N_2169,N_1786,N_55);
nand U2170 (N_2170,N_1011,N_885);
nor U2171 (N_2171,N_1797,N_347);
nand U2172 (N_2172,N_1289,N_1521);
or U2173 (N_2173,N_1707,N_1117);
and U2174 (N_2174,N_213,N_1576);
xor U2175 (N_2175,N_488,N_626);
and U2176 (N_2176,N_1235,N_1896);
nand U2177 (N_2177,N_197,N_469);
nor U2178 (N_2178,N_678,N_1758);
nor U2179 (N_2179,N_1523,N_382);
nor U2180 (N_2180,N_676,N_979);
nand U2181 (N_2181,N_1535,N_570);
or U2182 (N_2182,N_1306,N_546);
xnor U2183 (N_2183,N_1087,N_1054);
or U2184 (N_2184,N_1187,N_1574);
or U2185 (N_2185,N_48,N_800);
nor U2186 (N_2186,N_1709,N_96);
or U2187 (N_2187,N_1893,N_204);
and U2188 (N_2188,N_1967,N_1173);
nor U2189 (N_2189,N_1543,N_533);
xnor U2190 (N_2190,N_1126,N_1694);
nor U2191 (N_2191,N_1428,N_674);
and U2192 (N_2192,N_1027,N_1957);
nand U2193 (N_2193,N_1033,N_113);
and U2194 (N_2194,N_734,N_1865);
or U2195 (N_2195,N_174,N_395);
nor U2196 (N_2196,N_1882,N_1549);
xor U2197 (N_2197,N_785,N_1741);
nand U2198 (N_2198,N_80,N_1150);
nand U2199 (N_2199,N_283,N_1747);
and U2200 (N_2200,N_52,N_992);
nor U2201 (N_2201,N_1756,N_1229);
xor U2202 (N_2202,N_919,N_1935);
xnor U2203 (N_2203,N_1265,N_574);
xor U2204 (N_2204,N_1218,N_173);
or U2205 (N_2205,N_740,N_1047);
xor U2206 (N_2206,N_344,N_1141);
or U2207 (N_2207,N_1588,N_400);
nand U2208 (N_2208,N_223,N_1042);
xor U2209 (N_2209,N_1795,N_1250);
nand U2210 (N_2210,N_1932,N_985);
and U2211 (N_2211,N_1010,N_1599);
nand U2212 (N_2212,N_1032,N_638);
and U2213 (N_2213,N_1947,N_1556);
or U2214 (N_2214,N_596,N_1121);
xnor U2215 (N_2215,N_364,N_191);
nand U2216 (N_2216,N_1826,N_1853);
nand U2217 (N_2217,N_1198,N_150);
nor U2218 (N_2218,N_1911,N_278);
or U2219 (N_2219,N_1336,N_1467);
nor U2220 (N_2220,N_1246,N_1441);
and U2221 (N_2221,N_653,N_1035);
or U2222 (N_2222,N_1417,N_1889);
nand U2223 (N_2223,N_476,N_355);
and U2224 (N_2224,N_1468,N_750);
nor U2225 (N_2225,N_1200,N_1698);
xor U2226 (N_2226,N_962,N_1732);
xnor U2227 (N_2227,N_1729,N_1191);
nand U2228 (N_2228,N_1083,N_545);
xor U2229 (N_2229,N_380,N_1194);
or U2230 (N_2230,N_332,N_1550);
or U2231 (N_2231,N_1583,N_1196);
and U2232 (N_2232,N_1374,N_209);
nand U2233 (N_2233,N_29,N_587);
nor U2234 (N_2234,N_349,N_589);
xnor U2235 (N_2235,N_797,N_1723);
nor U2236 (N_2236,N_1045,N_1067);
xor U2237 (N_2237,N_884,N_226);
and U2238 (N_2238,N_583,N_377);
nand U2239 (N_2239,N_92,N_1909);
or U2240 (N_2240,N_298,N_83);
nand U2241 (N_2241,N_1926,N_1918);
or U2242 (N_2242,N_1999,N_1907);
nand U2243 (N_2243,N_1007,N_1681);
and U2244 (N_2244,N_1085,N_19);
nand U2245 (N_2245,N_590,N_807);
or U2246 (N_2246,N_1146,N_731);
or U2247 (N_2247,N_971,N_1605);
nand U2248 (N_2248,N_1781,N_1825);
and U2249 (N_2249,N_362,N_1447);
xnor U2250 (N_2250,N_891,N_504);
and U2251 (N_2251,N_1332,N_491);
and U2252 (N_2252,N_72,N_522);
and U2253 (N_2253,N_235,N_1157);
and U2254 (N_2254,N_783,N_974);
and U2255 (N_2255,N_315,N_1716);
nor U2256 (N_2256,N_1626,N_963);
xor U2257 (N_2257,N_1620,N_1969);
or U2258 (N_2258,N_903,N_1873);
or U2259 (N_2259,N_987,N_1129);
or U2260 (N_2260,N_508,N_1938);
xor U2261 (N_2261,N_74,N_10);
and U2262 (N_2262,N_1061,N_1750);
and U2263 (N_2263,N_1872,N_691);
or U2264 (N_2264,N_259,N_1369);
xnor U2265 (N_2265,N_1398,N_1041);
nand U2266 (N_2266,N_938,N_184);
xnor U2267 (N_2267,N_1153,N_618);
or U2268 (N_2268,N_123,N_900);
nor U2269 (N_2269,N_749,N_1902);
nor U2270 (N_2270,N_562,N_386);
or U2271 (N_2271,N_815,N_1419);
nor U2272 (N_2272,N_1831,N_1328);
nand U2273 (N_2273,N_648,N_677);
or U2274 (N_2274,N_1592,N_1536);
nand U2275 (N_2275,N_1390,N_310);
nor U2276 (N_2276,N_1179,N_490);
or U2277 (N_2277,N_1113,N_1365);
or U2278 (N_2278,N_1736,N_360);
and U2279 (N_2279,N_481,N_838);
nand U2280 (N_2280,N_224,N_569);
nand U2281 (N_2281,N_325,N_553);
xnor U2282 (N_2282,N_351,N_1575);
nor U2283 (N_2283,N_248,N_1589);
and U2284 (N_2284,N_564,N_1710);
xnor U2285 (N_2285,N_1922,N_742);
xnor U2286 (N_2286,N_519,N_980);
nor U2287 (N_2287,N_1635,N_1832);
nand U2288 (N_2288,N_1197,N_458);
and U2289 (N_2289,N_813,N_881);
and U2290 (N_2290,N_1691,N_972);
and U2291 (N_2291,N_1257,N_664);
xnor U2292 (N_2292,N_544,N_1817);
and U2293 (N_2293,N_289,N_1212);
xor U2294 (N_2294,N_338,N_1623);
or U2295 (N_2295,N_1993,N_424);
or U2296 (N_2296,N_1435,N_1813);
nand U2297 (N_2297,N_1248,N_1341);
and U2298 (N_2298,N_1128,N_746);
xor U2299 (N_2299,N_447,N_907);
or U2300 (N_2300,N_1586,N_1578);
and U2301 (N_2301,N_1326,N_592);
xor U2302 (N_2302,N_201,N_484);
nand U2303 (N_2303,N_465,N_643);
or U2304 (N_2304,N_1498,N_1663);
nor U2305 (N_2305,N_1975,N_936);
nor U2306 (N_2306,N_1404,N_527);
xor U2307 (N_2307,N_1319,N_473);
and U2308 (N_2308,N_687,N_127);
xor U2309 (N_2309,N_1174,N_879);
nand U2310 (N_2310,N_169,N_779);
and U2311 (N_2311,N_1481,N_1992);
xnor U2312 (N_2312,N_1704,N_1743);
or U2313 (N_2313,N_636,N_1841);
xor U2314 (N_2314,N_803,N_1609);
nor U2315 (N_2315,N_1119,N_652);
nor U2316 (N_2316,N_468,N_145);
or U2317 (N_2317,N_507,N_109);
nor U2318 (N_2318,N_824,N_1516);
and U2319 (N_2319,N_1343,N_940);
xor U2320 (N_2320,N_487,N_1991);
xor U2321 (N_2321,N_1293,N_893);
and U2322 (N_2322,N_620,N_852);
xnor U2323 (N_2323,N_1427,N_1386);
nor U2324 (N_2324,N_1759,N_878);
and U2325 (N_2325,N_133,N_820);
xor U2326 (N_2326,N_716,N_1622);
and U2327 (N_2327,N_186,N_207);
or U2328 (N_2328,N_1737,N_372);
or U2329 (N_2329,N_612,N_375);
and U2330 (N_2330,N_1043,N_1190);
nor U2331 (N_2331,N_1625,N_926);
nor U2332 (N_2332,N_1970,N_1809);
or U2333 (N_2333,N_417,N_1933);
xnor U2334 (N_2334,N_1439,N_1457);
or U2335 (N_2335,N_21,N_421);
or U2336 (N_2336,N_602,N_802);
nor U2337 (N_2337,N_523,N_739);
nor U2338 (N_2338,N_877,N_1616);
or U2339 (N_2339,N_100,N_1152);
xnor U2340 (N_2340,N_299,N_1411);
nand U2341 (N_2341,N_335,N_410);
nand U2342 (N_2342,N_761,N_287);
or U2343 (N_2343,N_1288,N_1924);
nor U2344 (N_2344,N_1392,N_1784);
nor U2345 (N_2345,N_120,N_700);
nor U2346 (N_2346,N_835,N_1090);
nor U2347 (N_2347,N_122,N_1327);
xor U2348 (N_2348,N_1548,N_208);
and U2349 (N_2349,N_1749,N_138);
or U2350 (N_2350,N_330,N_607);
xor U2351 (N_2351,N_1541,N_17);
xor U2352 (N_2352,N_1791,N_1779);
nor U2353 (N_2353,N_1836,N_1440);
nand U2354 (N_2354,N_274,N_1661);
or U2355 (N_2355,N_880,N_28);
or U2356 (N_2356,N_1894,N_241);
or U2357 (N_2357,N_718,N_516);
or U2358 (N_2358,N_1149,N_671);
and U2359 (N_2359,N_1864,N_1552);
nor U2360 (N_2360,N_751,N_49);
or U2361 (N_2361,N_780,N_702);
nor U2362 (N_2362,N_442,N_1952);
xor U2363 (N_2363,N_552,N_189);
xnor U2364 (N_2364,N_918,N_845);
nor U2365 (N_2365,N_485,N_924);
nor U2366 (N_2366,N_106,N_642);
or U2367 (N_2367,N_43,N_625);
and U2368 (N_2368,N_931,N_623);
xnor U2369 (N_2369,N_316,N_1943);
nand U2370 (N_2370,N_654,N_265);
nand U2371 (N_2371,N_670,N_872);
nor U2372 (N_2372,N_1805,N_1776);
and U2373 (N_2373,N_6,N_1513);
xor U2374 (N_2374,N_1585,N_1664);
xor U2375 (N_2375,N_1966,N_336);
and U2376 (N_2376,N_1961,N_1118);
nor U2377 (N_2377,N_45,N_1094);
or U2378 (N_2378,N_1740,N_1942);
nor U2379 (N_2379,N_912,N_1029);
nand U2380 (N_2380,N_1116,N_1526);
or U2381 (N_2381,N_211,N_890);
nor U2382 (N_2382,N_498,N_1093);
nand U2383 (N_2383,N_163,N_1068);
xor U2384 (N_2384,N_1269,N_238);
xor U2385 (N_2385,N_1820,N_1);
nor U2386 (N_2386,N_640,N_1590);
nor U2387 (N_2387,N_1358,N_439);
nor U2388 (N_2388,N_844,N_1900);
nand U2389 (N_2389,N_989,N_822);
xnor U2390 (N_2390,N_1725,N_396);
xor U2391 (N_2391,N_753,N_1848);
xnor U2392 (N_2392,N_1214,N_836);
or U2393 (N_2393,N_646,N_128);
or U2394 (N_2394,N_1842,N_1211);
nand U2395 (N_2395,N_1612,N_1475);
or U2396 (N_2396,N_404,N_764);
or U2397 (N_2397,N_768,N_1296);
or U2398 (N_2398,N_641,N_1808);
xnor U2399 (N_2399,N_268,N_1514);
nand U2400 (N_2400,N_1486,N_1112);
nor U2401 (N_2401,N_719,N_1920);
or U2402 (N_2402,N_1231,N_406);
xor U2403 (N_2403,N_1379,N_301);
nand U2404 (N_2404,N_1363,N_118);
nand U2405 (N_2405,N_1324,N_1656);
xnor U2406 (N_2406,N_1821,N_1771);
xnor U2407 (N_2407,N_886,N_1432);
or U2408 (N_2408,N_1164,N_1206);
nand U2409 (N_2409,N_1950,N_1854);
xor U2410 (N_2410,N_1163,N_777);
nor U2411 (N_2411,N_1003,N_1079);
nand U2412 (N_2412,N_1608,N_1693);
or U2413 (N_2413,N_98,N_246);
nand U2414 (N_2414,N_1582,N_1115);
nand U2415 (N_2415,N_1430,N_1653);
xnor U2416 (N_2416,N_581,N_1030);
nor U2417 (N_2417,N_512,N_772);
nor U2418 (N_2418,N_657,N_1223);
xnor U2419 (N_2419,N_1533,N_854);
or U2420 (N_2420,N_604,N_1345);
and U2421 (N_2421,N_811,N_818);
nand U2422 (N_2422,N_267,N_1302);
and U2423 (N_2423,N_613,N_1850);
and U2424 (N_2424,N_398,N_1593);
or U2425 (N_2425,N_1264,N_1192);
nor U2426 (N_2426,N_1478,N_90);
or U2427 (N_2427,N_935,N_565);
or U2428 (N_2428,N_1632,N_1718);
and U2429 (N_2429,N_1469,N_260);
nand U2430 (N_2430,N_1139,N_1183);
xnor U2431 (N_2431,N_1182,N_1254);
xnor U2432 (N_2432,N_525,N_1125);
nand U2433 (N_2433,N_1752,N_717);
or U2434 (N_2434,N_855,N_1760);
or U2435 (N_2435,N_506,N_1815);
nand U2436 (N_2436,N_1230,N_2);
or U2437 (N_2437,N_1692,N_1540);
and U2438 (N_2438,N_1249,N_1647);
nor U2439 (N_2439,N_703,N_1565);
or U2440 (N_2440,N_1026,N_1910);
nand U2441 (N_2441,N_187,N_825);
nand U2442 (N_2442,N_896,N_1215);
nor U2443 (N_2443,N_555,N_1666);
xnor U2444 (N_2444,N_1299,N_913);
xor U2445 (N_2445,N_182,N_279);
or U2446 (N_2446,N_1025,N_1189);
or U2447 (N_2447,N_1930,N_579);
xor U2448 (N_2448,N_948,N_1772);
and U2449 (N_2449,N_883,N_114);
or U2450 (N_2450,N_933,N_308);
nand U2451 (N_2451,N_1645,N_39);
nand U2452 (N_2452,N_1280,N_995);
or U2453 (N_2453,N_1673,N_361);
and U2454 (N_2454,N_75,N_1267);
nand U2455 (N_2455,N_1453,N_1237);
nand U2456 (N_2456,N_908,N_1977);
nand U2457 (N_2457,N_1726,N_1835);
or U2458 (N_2458,N_1558,N_551);
nor U2459 (N_2459,N_1506,N_517);
nand U2460 (N_2460,N_176,N_1847);
nand U2461 (N_2461,N_821,N_826);
xnor U2462 (N_2462,N_1073,N_1505);
or U2463 (N_2463,N_390,N_639);
xor U2464 (N_2464,N_358,N_1744);
and U2465 (N_2465,N_1519,N_1721);
xor U2466 (N_2466,N_32,N_1906);
xnor U2467 (N_2467,N_467,N_367);
nand U2468 (N_2468,N_1923,N_1178);
xnor U2469 (N_2469,N_939,N_1104);
and U2470 (N_2470,N_720,N_511);
nand U2471 (N_2471,N_220,N_1266);
and U2472 (N_2472,N_631,N_141);
nor U2473 (N_2473,N_914,N_392);
or U2474 (N_2474,N_401,N_1133);
and U2475 (N_2475,N_64,N_143);
or U2476 (N_2476,N_591,N_1881);
nor U2477 (N_2477,N_1364,N_1822);
and U2478 (N_2478,N_696,N_1408);
or U2479 (N_2479,N_1542,N_381);
or U2480 (N_2480,N_46,N_276);
or U2481 (N_2481,N_1789,N_804);
nand U2482 (N_2482,N_306,N_236);
or U2483 (N_2483,N_1739,N_12);
or U2484 (N_2484,N_769,N_850);
xnor U2485 (N_2485,N_23,N_759);
nand U2486 (N_2486,N_1451,N_927);
or U2487 (N_2487,N_97,N_399);
nor U2488 (N_2488,N_853,N_1354);
and U2489 (N_2489,N_1470,N_1699);
and U2490 (N_2490,N_124,N_1362);
or U2491 (N_2491,N_586,N_1564);
and U2492 (N_2492,N_105,N_823);
and U2493 (N_2493,N_103,N_431);
and U2494 (N_2494,N_1239,N_550);
nand U2495 (N_2495,N_302,N_125);
nor U2496 (N_2496,N_1180,N_1518);
nand U2497 (N_2497,N_1165,N_1980);
xor U2498 (N_2498,N_566,N_1378);
xnor U2499 (N_2499,N_1352,N_524);
and U2500 (N_2500,N_1399,N_601);
nor U2501 (N_2501,N_1509,N_1951);
nor U2502 (N_2502,N_1074,N_951);
xor U2503 (N_2503,N_326,N_1803);
and U2504 (N_2504,N_1049,N_937);
nand U2505 (N_2505,N_432,N_1837);
nor U2506 (N_2506,N_1985,N_252);
or U2507 (N_2507,N_1487,N_1325);
xor U2508 (N_2508,N_1001,N_1017);
xnor U2509 (N_2509,N_181,N_292);
xor U2510 (N_2510,N_388,N_1274);
and U2511 (N_2511,N_1044,N_1678);
nand U2512 (N_2512,N_492,N_1954);
or U2513 (N_2513,N_1140,N_333);
xnor U2514 (N_2514,N_887,N_864);
nand U2515 (N_2515,N_1330,N_448);
nor U2516 (N_2516,N_1863,N_665);
xnor U2517 (N_2517,N_1219,N_146);
nand U2518 (N_2518,N_194,N_983);
xor U2519 (N_2519,N_997,N_1504);
nor U2520 (N_2520,N_1688,N_969);
and U2521 (N_2521,N_1314,N_1446);
or U2522 (N_2522,N_1990,N_1203);
and U2523 (N_2523,N_978,N_1078);
and U2524 (N_2524,N_628,N_1037);
or U2525 (N_2525,N_635,N_1484);
nand U2526 (N_2526,N_542,N_1458);
nand U2527 (N_2527,N_379,N_1367);
or U2528 (N_2528,N_1719,N_1800);
nor U2529 (N_2529,N_1309,N_1123);
nand U2530 (N_2530,N_603,N_300);
xor U2531 (N_2531,N_244,N_1331);
nor U2532 (N_2532,N_1611,N_1410);
nand U2533 (N_2533,N_520,N_1473);
or U2534 (N_2534,N_1960,N_1801);
nor U2535 (N_2535,N_790,N_1994);
or U2536 (N_2536,N_1476,N_1065);
nand U2537 (N_2537,N_1221,N_1301);
or U2538 (N_2538,N_1898,N_672);
nand U2539 (N_2539,N_130,N_744);
xor U2540 (N_2540,N_88,N_827);
nor U2541 (N_2541,N_402,N_166);
nor U2542 (N_2542,N_1829,N_85);
nand U2543 (N_2543,N_405,N_578);
and U2544 (N_2544,N_249,N_1763);
nand U2545 (N_2545,N_1668,N_911);
nand U2546 (N_2546,N_385,N_521);
nor U2547 (N_2547,N_451,N_1291);
xnor U2548 (N_2548,N_724,N_1005);
nand U2549 (N_2549,N_62,N_1782);
nor U2550 (N_2550,N_658,N_243);
xor U2551 (N_2551,N_178,N_1751);
or U2552 (N_2552,N_461,N_171);
nor U2553 (N_2553,N_416,N_1874);
nand U2554 (N_2554,N_662,N_408);
or U2555 (N_2555,N_1675,N_394);
xor U2556 (N_2556,N_1095,N_1006);
nand U2557 (N_2557,N_743,N_1708);
xor U2558 (N_2558,N_414,N_1396);
or U2559 (N_2559,N_206,N_423);
and U2560 (N_2560,N_445,N_1019);
nor U2561 (N_2561,N_1429,N_444);
or U2562 (N_2562,N_869,N_1497);
and U2563 (N_2563,N_942,N_263);
and U2564 (N_2564,N_708,N_1004);
and U2565 (N_2565,N_1009,N_1089);
or U2566 (N_2566,N_205,N_1557);
nor U2567 (N_2567,N_1715,N_1477);
nand U2568 (N_2568,N_1802,N_1677);
nand U2569 (N_2569,N_78,N_757);
nand U2570 (N_2570,N_428,N_1731);
xor U2571 (N_2571,N_1703,N_760);
nor U2572 (N_2572,N_1166,N_1816);
and U2573 (N_2573,N_1886,N_1472);
or U2574 (N_2574,N_54,N_832);
nor U2575 (N_2575,N_1921,N_162);
and U2576 (N_2576,N_650,N_353);
nor U2577 (N_2577,N_1147,N_1234);
nand U2578 (N_2578,N_1335,N_1644);
nor U2579 (N_2579,N_661,N_1834);
nor U2580 (N_2580,N_1738,N_1077);
and U2581 (N_2581,N_944,N_588);
or U2582 (N_2582,N_1525,N_1076);
xnor U2583 (N_2583,N_810,N_411);
xor U2584 (N_2584,N_253,N_786);
nor U2585 (N_2585,N_1071,N_1807);
xnor U2586 (N_2586,N_1627,N_1081);
nor U2587 (N_2587,N_1347,N_932);
or U2588 (N_2588,N_975,N_1305);
xnor U2589 (N_2589,N_801,N_1438);
xnor U2590 (N_2590,N_929,N_1381);
nand U2591 (N_2591,N_1253,N_486);
and U2592 (N_2592,N_575,N_460);
nand U2593 (N_2593,N_264,N_495);
nand U2594 (N_2594,N_1532,N_1818);
nand U2595 (N_2595,N_15,N_1614);
and U2596 (N_2596,N_624,N_307);
nor U2597 (N_2597,N_796,N_1416);
nand U2598 (N_2598,N_1461,N_647);
and U2599 (N_2599,N_1023,N_1948);
nor U2600 (N_2600,N_1722,N_1217);
nand U2601 (N_2601,N_37,N_1244);
or U2602 (N_2602,N_736,N_441);
nand U2603 (N_2603,N_1151,N_679);
and U2604 (N_2604,N_1610,N_323);
nand U2605 (N_2605,N_429,N_1107);
xnor U2606 (N_2606,N_1159,N_1591);
and U2607 (N_2607,N_770,N_1904);
or U2608 (N_2608,N_1339,N_1383);
xor U2609 (N_2609,N_1639,N_861);
xnor U2610 (N_2610,N_1413,N_1425);
or U2611 (N_2611,N_946,N_1819);
and U2612 (N_2612,N_470,N_240);
nor U2613 (N_2613,N_1082,N_167);
or U2614 (N_2614,N_794,N_314);
and U2615 (N_2615,N_286,N_257);
or U2616 (N_2616,N_285,N_1134);
or U2617 (N_2617,N_440,N_1313);
nor U2618 (N_2618,N_1021,N_450);
xor U2619 (N_2619,N_1785,N_952);
nor U2620 (N_2620,N_1437,N_1573);
nand U2621 (N_2621,N_1928,N_1207);
and U2622 (N_2622,N_1176,N_108);
or U2623 (N_2623,N_1903,N_960);
nor U2624 (N_2624,N_1359,N_1444);
nor U2625 (N_2625,N_1016,N_1355);
nor U2626 (N_2626,N_1761,N_1051);
or U2627 (N_2627,N_1720,N_805);
xor U2628 (N_2628,N_477,N_1375);
nor U2629 (N_2629,N_296,N_1662);
or U2630 (N_2630,N_725,N_1884);
xor U2631 (N_2631,N_1474,N_728);
nor U2632 (N_2632,N_686,N_945);
nand U2633 (N_2633,N_959,N_1858);
nor U2634 (N_2634,N_1931,N_1220);
xor U2635 (N_2635,N_1370,N_1272);
or U2636 (N_2636,N_1679,N_1833);
and U2637 (N_2637,N_1238,N_537);
xor U2638 (N_2638,N_112,N_212);
nor U2639 (N_2639,N_73,N_1420);
or U2640 (N_2640,N_667,N_917);
xor U2641 (N_2641,N_304,N_982);
nor U2642 (N_2642,N_328,N_430);
or U2643 (N_2643,N_1316,N_1479);
and U2644 (N_2644,N_1142,N_192);
xor U2645 (N_2645,N_1485,N_1110);
and U2646 (N_2646,N_505,N_11);
nor U2647 (N_2647,N_955,N_1395);
nand U2648 (N_2648,N_1508,N_1048);
nor U2649 (N_2649,N_1885,N_967);
and U2650 (N_2650,N_1137,N_1412);
or U2651 (N_2651,N_921,N_526);
or U2652 (N_2652,N_1184,N_94);
nand U2653 (N_2653,N_876,N_1908);
or U2654 (N_2654,N_1979,N_535);
and U2655 (N_2655,N_1394,N_1615);
xor U2656 (N_2656,N_269,N_1554);
and U2657 (N_2657,N_1891,N_1422);
nand U2658 (N_2658,N_541,N_1774);
nor U2659 (N_2659,N_1450,N_26);
or U2660 (N_2660,N_1946,N_1460);
nand U2661 (N_2661,N_219,N_1055);
nor U2662 (N_2662,N_1344,N_617);
nand U2663 (N_2663,N_1275,N_13);
xor U2664 (N_2664,N_1000,N_1814);
nor U2665 (N_2665,N_1669,N_1547);
xor U2666 (N_2666,N_1755,N_1193);
or U2667 (N_2667,N_418,N_1167);
and U2668 (N_2668,N_331,N_144);
or U2669 (N_2669,N_1511,N_1012);
nor U2670 (N_2670,N_1560,N_1415);
or U2671 (N_2671,N_121,N_619);
xor U2672 (N_2672,N_471,N_1298);
nand U2673 (N_2673,N_457,N_1433);
nor U2674 (N_2674,N_1161,N_1282);
nor U2675 (N_2675,N_765,N_1224);
and U2676 (N_2676,N_327,N_270);
xor U2677 (N_2677,N_422,N_536);
xor U2678 (N_2678,N_1767,N_528);
nand U2679 (N_2679,N_1056,N_1628);
and U2680 (N_2680,N_1631,N_817);
or U2681 (N_2681,N_350,N_1697);
nand U2682 (N_2682,N_57,N_1263);
or U2683 (N_2683,N_1849,N_577);
or U2684 (N_2684,N_1777,N_984);
nor U2685 (N_2685,N_1968,N_1810);
xnor U2686 (N_2686,N_1792,N_732);
xor U2687 (N_2687,N_1366,N_1579);
or U2688 (N_2688,N_633,N_1205);
nor U2689 (N_2689,N_655,N_1949);
nand U2690 (N_2690,N_1945,N_943);
nand U2691 (N_2691,N_5,N_343);
and U2692 (N_2692,N_1637,N_1471);
xnor U2693 (N_2693,N_66,N_1619);
and U2694 (N_2694,N_899,N_1838);
xor U2695 (N_2695,N_1418,N_1659);
nor U2696 (N_2696,N_126,N_572);
or U2697 (N_2697,N_297,N_165);
nor U2698 (N_2698,N_1100,N_897);
xor U2699 (N_2699,N_217,N_1072);
nand U2700 (N_2700,N_1340,N_322);
or U2701 (N_2701,N_1912,N_295);
xnor U2702 (N_2702,N_1941,N_1643);
xnor U2703 (N_2703,N_272,N_685);
nor U2704 (N_2704,N_1887,N_340);
nor U2705 (N_2705,N_464,N_1764);
and U2706 (N_2706,N_1039,N_738);
or U2707 (N_2707,N_210,N_119);
or U2708 (N_2708,N_684,N_449);
xnor U2709 (N_2709,N_1522,N_622);
or U2710 (N_2710,N_1389,N_950);
nand U2711 (N_2711,N_540,N_1105);
xor U2712 (N_2712,N_1080,N_1225);
or U2713 (N_2713,N_1901,N_1273);
nand U2714 (N_2714,N_634,N_1292);
nand U2715 (N_2715,N_1131,N_789);
and U2716 (N_2716,N_681,N_1641);
nand U2717 (N_2717,N_1798,N_1512);
or U2718 (N_2718,N_568,N_216);
nand U2719 (N_2719,N_1276,N_894);
and U2720 (N_2720,N_1642,N_337);
nor U2721 (N_2721,N_161,N_3);
nand U2722 (N_2722,N_1530,N_1799);
and U2723 (N_2723,N_478,N_994);
nand U2724 (N_2724,N_645,N_1917);
xor U2725 (N_2725,N_51,N_889);
or U2726 (N_2726,N_726,N_459);
or U2727 (N_2727,N_489,N_843);
nand U2728 (N_2728,N_1448,N_758);
and U2729 (N_2729,N_502,N_1845);
nor U2730 (N_2730,N_1099,N_1138);
and U2731 (N_2731,N_530,N_503);
or U2732 (N_2732,N_977,N_1689);
and U2733 (N_2733,N_1232,N_1024);
or U2734 (N_2734,N_1445,N_1069);
xnor U2735 (N_2735,N_1015,N_1876);
nand U2736 (N_2736,N_795,N_695);
xor U2737 (N_2737,N_1890,N_1913);
xor U2738 (N_2738,N_203,N_1322);
nand U2739 (N_2739,N_1955,N_1603);
nor U2740 (N_2740,N_1188,N_669);
and U2741 (N_2741,N_376,N_1870);
and U2742 (N_2742,N_1463,N_1442);
nand U2743 (N_2743,N_1062,N_727);
or U2744 (N_2744,N_44,N_368);
or U2745 (N_2745,N_291,N_27);
or U2746 (N_2746,N_76,N_961);
nand U2747 (N_2747,N_1633,N_1260);
and U2748 (N_2748,N_1202,N_814);
nand U2749 (N_2749,N_501,N_1859);
and U2750 (N_2750,N_1529,N_582);
xor U2751 (N_2751,N_1734,N_1064);
and U2752 (N_2752,N_713,N_605);
nand U2753 (N_2753,N_294,N_925);
and U2754 (N_2754,N_875,N_741);
nand U2755 (N_2755,N_104,N_1155);
or U2756 (N_2756,N_1284,N_1500);
nand U2757 (N_2757,N_1929,N_1851);
and U2758 (N_2758,N_1488,N_968);
or U2759 (N_2759,N_93,N_412);
and U2760 (N_2760,N_1840,N_1866);
or U2761 (N_2761,N_370,N_1934);
and U2762 (N_2762,N_1915,N_1587);
nand U2763 (N_2763,N_668,N_1959);
xnor U2764 (N_2764,N_1209,N_1563);
and U2765 (N_2765,N_1844,N_1300);
or U2766 (N_2766,N_1058,N_345);
and U2767 (N_2767,N_531,N_766);
xnor U2768 (N_2768,N_1333,N_1769);
and U2769 (N_2769,N_247,N_303);
xnor U2770 (N_2770,N_1974,N_42);
nor U2771 (N_2771,N_762,N_233);
or U2772 (N_2772,N_148,N_1046);
and U2773 (N_2773,N_497,N_309);
nor U2774 (N_2774,N_1775,N_529);
or U2775 (N_2775,N_1537,N_584);
nor U2776 (N_2776,N_446,N_910);
nor U2777 (N_2777,N_1312,N_856);
nand U2778 (N_2778,N_312,N_755);
xnor U2779 (N_2779,N_1098,N_547);
nor U2780 (N_2780,N_1524,N_629);
or U2781 (N_2781,N_102,N_1730);
xnor U2782 (N_2782,N_737,N_651);
xor U2783 (N_2783,N_463,N_1057);
or U2784 (N_2784,N_1783,N_1407);
nor U2785 (N_2785,N_305,N_915);
or U2786 (N_2786,N_816,N_576);
xor U2787 (N_2787,N_1278,N_1754);
xor U2788 (N_2788,N_1830,N_610);
nor U2789 (N_2789,N_1962,N_1222);
xor U2790 (N_2790,N_117,N_36);
or U2791 (N_2791,N_1507,N_1944);
xor U2792 (N_2792,N_149,N_692);
xnor U2793 (N_2793,N_627,N_787);
nor U2794 (N_2794,N_782,N_867);
nor U2795 (N_2795,N_870,N_453);
xor U2796 (N_2796,N_1145,N_1028);
nor U2797 (N_2797,N_237,N_1135);
xnor U2798 (N_2798,N_683,N_1683);
and U2799 (N_2799,N_953,N_151);
nand U2800 (N_2800,N_1702,N_649);
nand U2801 (N_2801,N_906,N_1986);
nand U2802 (N_2802,N_1059,N_1973);
or U2803 (N_2803,N_1572,N_215);
or U2804 (N_2804,N_895,N_1031);
xor U2805 (N_2805,N_69,N_513);
nor U2806 (N_2806,N_756,N_1682);
or U2807 (N_2807,N_1652,N_812);
nor U2808 (N_2808,N_1384,N_419);
and U2809 (N_2809,N_70,N_615);
nor U2810 (N_2810,N_611,N_1465);
nor U2811 (N_2811,N_1349,N_630);
nand U2812 (N_2812,N_1562,N_65);
or U2813 (N_2813,N_1084,N_50);
nor U2814 (N_2814,N_1671,N_1013);
nand U2815 (N_2815,N_357,N_1839);
xnor U2816 (N_2816,N_475,N_1400);
nor U2817 (N_2817,N_868,N_139);
and U2818 (N_2818,N_1939,N_1216);
nor U2819 (N_2819,N_86,N_698);
xnor U2820 (N_2820,N_666,N_996);
xnor U2821 (N_2821,N_1154,N_34);
xor U2822 (N_2822,N_958,N_1103);
and U2823 (N_2823,N_24,N_1971);
or U2824 (N_2824,N_230,N_510);
nor U2825 (N_2825,N_1595,N_1766);
xnor U2826 (N_2826,N_548,N_1106);
nor U2827 (N_2827,N_1571,N_571);
nand U2828 (N_2828,N_1602,N_1053);
or U2829 (N_2829,N_1348,N_183);
and U2830 (N_2830,N_659,N_1294);
xor U2831 (N_2831,N_1796,N_1618);
or U2832 (N_2832,N_393,N_831);
nor U2833 (N_2833,N_188,N_1290);
or U2834 (N_2834,N_190,N_1528);
nor U2835 (N_2835,N_859,N_1765);
nor U2836 (N_2836,N_1899,N_1606);
or U2837 (N_2837,N_158,N_1101);
or U2838 (N_2838,N_1279,N_1295);
nand U2839 (N_2839,N_1640,N_227);
or U2840 (N_2840,N_1227,N_1714);
nor U2841 (N_2841,N_606,N_1136);
nand U2842 (N_2842,N_1860,N_1995);
xnor U2843 (N_2843,N_673,N_1806);
nor U2844 (N_2844,N_250,N_1735);
nand U2845 (N_2845,N_776,N_1981);
and U2846 (N_2846,N_834,N_1978);
or U2847 (N_2847,N_493,N_1676);
nor U2848 (N_2848,N_556,N_1517);
or U2849 (N_2849,N_1778,N_157);
xor U2850 (N_2850,N_543,N_558);
nor U2851 (N_2851,N_976,N_61);
and U2852 (N_2852,N_371,N_1482);
nor U2853 (N_2853,N_1462,N_1255);
or U2854 (N_2854,N_232,N_988);
and U2855 (N_2855,N_1824,N_1143);
and U2856 (N_2856,N_1002,N_1495);
nand U2857 (N_2857,N_1213,N_752);
xnor U2858 (N_2858,N_1034,N_1494);
nor U2859 (N_2859,N_1382,N_426);
nor U2860 (N_2860,N_998,N_354);
xor U2861 (N_2861,N_1391,N_715);
and U2862 (N_2862,N_319,N_771);
and U2863 (N_2863,N_378,N_1976);
or U2864 (N_2864,N_1144,N_784);
and U2865 (N_2865,N_1594,N_1843);
and U2866 (N_2866,N_231,N_271);
or U2867 (N_2867,N_348,N_342);
xor U2868 (N_2868,N_1545,N_1658);
nand U2869 (N_2869,N_585,N_1414);
nor U2870 (N_2870,N_1988,N_277);
xor U2871 (N_2871,N_922,N_690);
nor U2872 (N_2872,N_1733,N_594);
and U2873 (N_2873,N_1927,N_773);
nand U2874 (N_2874,N_1108,N_466);
and U2875 (N_2875,N_865,N_198);
and U2876 (N_2876,N_1787,N_842);
nand U2877 (N_2877,N_561,N_1050);
nand U2878 (N_2878,N_663,N_164);
nor U2879 (N_2879,N_195,N_898);
and U2880 (N_2880,N_8,N_1456);
nor U2881 (N_2881,N_433,N_1008);
or U2882 (N_2882,N_1996,N_1665);
and U2883 (N_2883,N_775,N_608);
nand U2884 (N_2884,N_1466,N_1443);
xnor U2885 (N_2885,N_1014,N_282);
or U2886 (N_2886,N_275,N_1403);
nor U2887 (N_2887,N_1621,N_1857);
nor U2888 (N_2888,N_682,N_595);
xnor U2889 (N_2889,N_1449,N_427);
and U2890 (N_2890,N_1169,N_403);
nor U2891 (N_2891,N_563,N_707);
or U2892 (N_2892,N_456,N_830);
nor U2893 (N_2893,N_1258,N_95);
nor U2894 (N_2894,N_1655,N_621);
nor U2895 (N_2895,N_1937,N_1177);
xor U2896 (N_2896,N_1185,N_866);
and U2897 (N_2897,N_1052,N_809);
nand U2898 (N_2898,N_214,N_1982);
nor U2899 (N_2899,N_710,N_1120);
or U2900 (N_2900,N_391,N_1252);
or U2901 (N_2901,N_1496,N_1020);
xor U2902 (N_2902,N_281,N_1686);
nand U2903 (N_2903,N_1075,N_339);
and U2904 (N_2904,N_567,N_806);
or U2905 (N_2905,N_828,N_1170);
or U2906 (N_2906,N_59,N_132);
nor U2907 (N_2907,N_1038,N_1983);
or U2908 (N_2908,N_1361,N_82);
and U2909 (N_2909,N_990,N_799);
xnor U2910 (N_2910,N_1538,N_721);
and U2911 (N_2911,N_53,N_1111);
or U2912 (N_2912,N_1317,N_0);
xnor U2913 (N_2913,N_599,N_482);
and U2914 (N_2914,N_1780,N_320);
and U2915 (N_2915,N_1247,N_1919);
nor U2916 (N_2916,N_1063,N_352);
nand U2917 (N_2917,N_500,N_735);
nand U2918 (N_2918,N_1674,N_185);
or U2919 (N_2919,N_1515,N_480);
or U2920 (N_2920,N_774,N_1283);
nor U2921 (N_2921,N_1204,N_107);
nor U2922 (N_2922,N_455,N_518);
nor U2923 (N_2923,N_557,N_1060);
nand U2924 (N_2924,N_1531,N_1434);
nor U2925 (N_2925,N_614,N_839);
or U2926 (N_2926,N_115,N_1613);
xor U2927 (N_2927,N_675,N_142);
and U2928 (N_2928,N_1555,N_79);
nor U2929 (N_2929,N_1936,N_1357);
and U2930 (N_2930,N_1181,N_981);
and U2931 (N_2931,N_1680,N_373);
xnor U2932 (N_2932,N_262,N_873);
and U2933 (N_2933,N_1338,N_1372);
and U2934 (N_2934,N_1701,N_1156);
or U2935 (N_2935,N_99,N_1377);
xor U2936 (N_2936,N_1965,N_218);
nor U2937 (N_2937,N_1877,N_359);
or U2938 (N_2938,N_632,N_597);
nand U2939 (N_2939,N_1480,N_841);
nand U2940 (N_2940,N_1455,N_767);
nand U2941 (N_2941,N_311,N_1753);
nand U2942 (N_2942,N_436,N_89);
and U2943 (N_2943,N_1268,N_1636);
or U2944 (N_2944,N_1307,N_1036);
xor U2945 (N_2945,N_532,N_902);
or U2946 (N_2946,N_1916,N_443);
and U2947 (N_2947,N_221,N_366);
and U2948 (N_2948,N_947,N_452);
or U2949 (N_2949,N_1584,N_229);
xnor U2950 (N_2950,N_1559,N_851);
and U2951 (N_2951,N_1318,N_1577);
nand U2952 (N_2952,N_1527,N_849);
or U2953 (N_2953,N_701,N_1195);
xnor U2954 (N_2954,N_494,N_1421);
nand U2955 (N_2955,N_1705,N_87);
xor U2956 (N_2956,N_1868,N_1762);
xnor U2957 (N_2957,N_1812,N_1208);
or U2958 (N_2958,N_1687,N_56);
nor U2959 (N_2959,N_534,N_1356);
nand U2960 (N_2960,N_1226,N_1657);
nand U2961 (N_2961,N_474,N_934);
nor U2962 (N_2962,N_1696,N_704);
xor U2963 (N_2963,N_160,N_1892);
nand U2964 (N_2964,N_1483,N_22);
nand U2965 (N_2965,N_1598,N_1380);
xor U2966 (N_2966,N_1879,N_1242);
nor U2967 (N_2967,N_920,N_1638);
xor U2968 (N_2968,N_1728,N_949);
xnor U2969 (N_2969,N_1277,N_509);
nand U2970 (N_2970,N_1281,N_1210);
xnor U2971 (N_2971,N_1617,N_1905);
nand U2972 (N_2972,N_1972,N_580);
or U2973 (N_2973,N_435,N_1426);
or U2974 (N_2974,N_1130,N_1650);
and U2975 (N_2975,N_1629,N_1684);
nor U2976 (N_2976,N_847,N_84);
xnor U2977 (N_2977,N_245,N_1376);
and U2978 (N_2978,N_1091,N_389);
xor U2979 (N_2979,N_1869,N_318);
xnor U2980 (N_2980,N_256,N_549);
nand U2981 (N_2981,N_135,N_1551);
nor U2982 (N_2982,N_293,N_829);
nor U2983 (N_2983,N_1452,N_1914);
nand U2984 (N_2984,N_1672,N_77);
and U2985 (N_2985,N_637,N_788);
nand U2986 (N_2986,N_228,N_1070);
or U2987 (N_2987,N_1757,N_1109);
nor U2988 (N_2988,N_1570,N_47);
nand U2989 (N_2989,N_1360,N_1436);
nor U2990 (N_2990,N_1018,N_1160);
and U2991 (N_2991,N_1987,N_1648);
nand U2992 (N_2992,N_407,N_697);
xor U2993 (N_2993,N_63,N_1285);
nand U2994 (N_2994,N_1233,N_1406);
and U2995 (N_2995,N_778,N_1958);
xor U2996 (N_2996,N_1393,N_479);
nand U2997 (N_2997,N_1423,N_694);
and U2998 (N_2998,N_438,N_18);
nor U2999 (N_2999,N_1175,N_14);
or U3000 (N_3000,N_341,N_1467);
nor U3001 (N_3001,N_1172,N_1722);
xnor U3002 (N_3002,N_1547,N_396);
and U3003 (N_3003,N_1923,N_340);
nand U3004 (N_3004,N_248,N_1745);
nor U3005 (N_3005,N_1762,N_1826);
and U3006 (N_3006,N_1891,N_309);
nor U3007 (N_3007,N_98,N_1772);
xnor U3008 (N_3008,N_1942,N_1163);
nand U3009 (N_3009,N_1760,N_1089);
and U3010 (N_3010,N_1820,N_529);
xor U3011 (N_3011,N_599,N_837);
nor U3012 (N_3012,N_199,N_437);
nor U3013 (N_3013,N_620,N_839);
nand U3014 (N_3014,N_867,N_1855);
or U3015 (N_3015,N_1544,N_1363);
nand U3016 (N_3016,N_1776,N_1666);
xnor U3017 (N_3017,N_667,N_1168);
or U3018 (N_3018,N_285,N_454);
xor U3019 (N_3019,N_1900,N_146);
nand U3020 (N_3020,N_354,N_1826);
nor U3021 (N_3021,N_1981,N_1193);
nand U3022 (N_3022,N_779,N_1608);
xnor U3023 (N_3023,N_1078,N_120);
nor U3024 (N_3024,N_1122,N_896);
nand U3025 (N_3025,N_1659,N_1853);
nand U3026 (N_3026,N_855,N_1176);
xor U3027 (N_3027,N_52,N_1869);
nor U3028 (N_3028,N_148,N_1102);
or U3029 (N_3029,N_1106,N_1908);
nand U3030 (N_3030,N_847,N_955);
or U3031 (N_3031,N_1365,N_1988);
xnor U3032 (N_3032,N_661,N_1349);
and U3033 (N_3033,N_495,N_1358);
and U3034 (N_3034,N_154,N_816);
and U3035 (N_3035,N_366,N_775);
and U3036 (N_3036,N_936,N_1461);
nand U3037 (N_3037,N_980,N_207);
xor U3038 (N_3038,N_1336,N_622);
nor U3039 (N_3039,N_1278,N_1568);
xnor U3040 (N_3040,N_1282,N_820);
nand U3041 (N_3041,N_1344,N_605);
nand U3042 (N_3042,N_295,N_1877);
nand U3043 (N_3043,N_11,N_1754);
nand U3044 (N_3044,N_826,N_570);
xnor U3045 (N_3045,N_638,N_296);
and U3046 (N_3046,N_1946,N_401);
nor U3047 (N_3047,N_1981,N_400);
nor U3048 (N_3048,N_1409,N_446);
and U3049 (N_3049,N_370,N_1933);
nor U3050 (N_3050,N_1249,N_1408);
nand U3051 (N_3051,N_1658,N_1308);
and U3052 (N_3052,N_425,N_154);
and U3053 (N_3053,N_1805,N_913);
xor U3054 (N_3054,N_1592,N_825);
nand U3055 (N_3055,N_1672,N_685);
nand U3056 (N_3056,N_471,N_617);
or U3057 (N_3057,N_809,N_1253);
nand U3058 (N_3058,N_985,N_350);
nand U3059 (N_3059,N_90,N_1329);
xnor U3060 (N_3060,N_1025,N_568);
or U3061 (N_3061,N_1306,N_238);
and U3062 (N_3062,N_100,N_1598);
nand U3063 (N_3063,N_1856,N_284);
nand U3064 (N_3064,N_644,N_1750);
nor U3065 (N_3065,N_1565,N_628);
xor U3066 (N_3066,N_512,N_1662);
or U3067 (N_3067,N_8,N_1636);
xnor U3068 (N_3068,N_560,N_562);
and U3069 (N_3069,N_1736,N_1535);
and U3070 (N_3070,N_83,N_55);
and U3071 (N_3071,N_594,N_1674);
or U3072 (N_3072,N_252,N_1382);
nor U3073 (N_3073,N_683,N_1461);
or U3074 (N_3074,N_279,N_492);
and U3075 (N_3075,N_736,N_255);
nand U3076 (N_3076,N_1662,N_1009);
nand U3077 (N_3077,N_1932,N_25);
nand U3078 (N_3078,N_370,N_1768);
xnor U3079 (N_3079,N_1197,N_322);
and U3080 (N_3080,N_1973,N_606);
and U3081 (N_3081,N_1573,N_1841);
and U3082 (N_3082,N_1851,N_1201);
or U3083 (N_3083,N_51,N_1659);
nor U3084 (N_3084,N_327,N_242);
xor U3085 (N_3085,N_1054,N_829);
nor U3086 (N_3086,N_1605,N_5);
or U3087 (N_3087,N_737,N_1587);
and U3088 (N_3088,N_1003,N_246);
nor U3089 (N_3089,N_1830,N_353);
nand U3090 (N_3090,N_635,N_497);
nor U3091 (N_3091,N_1150,N_1057);
xor U3092 (N_3092,N_1571,N_1969);
nor U3093 (N_3093,N_1652,N_1459);
or U3094 (N_3094,N_1077,N_1407);
or U3095 (N_3095,N_1848,N_206);
nor U3096 (N_3096,N_1770,N_736);
xor U3097 (N_3097,N_994,N_1218);
and U3098 (N_3098,N_1288,N_1283);
nand U3099 (N_3099,N_1216,N_1657);
xor U3100 (N_3100,N_1360,N_1409);
or U3101 (N_3101,N_1571,N_1586);
nor U3102 (N_3102,N_869,N_1857);
xnor U3103 (N_3103,N_360,N_1296);
nand U3104 (N_3104,N_804,N_963);
xor U3105 (N_3105,N_1214,N_1204);
nor U3106 (N_3106,N_524,N_724);
and U3107 (N_3107,N_256,N_1591);
and U3108 (N_3108,N_1207,N_540);
xnor U3109 (N_3109,N_1306,N_1239);
xnor U3110 (N_3110,N_1978,N_1552);
xnor U3111 (N_3111,N_950,N_1916);
nor U3112 (N_3112,N_1132,N_147);
xnor U3113 (N_3113,N_1462,N_662);
xnor U3114 (N_3114,N_107,N_116);
nor U3115 (N_3115,N_1011,N_1167);
nor U3116 (N_3116,N_610,N_1295);
xnor U3117 (N_3117,N_110,N_375);
xor U3118 (N_3118,N_1842,N_689);
nor U3119 (N_3119,N_1932,N_330);
xnor U3120 (N_3120,N_1486,N_797);
and U3121 (N_3121,N_1655,N_1314);
nor U3122 (N_3122,N_1847,N_1000);
nor U3123 (N_3123,N_1367,N_91);
nor U3124 (N_3124,N_224,N_763);
nor U3125 (N_3125,N_1521,N_1609);
or U3126 (N_3126,N_580,N_200);
xor U3127 (N_3127,N_944,N_781);
nand U3128 (N_3128,N_1295,N_1031);
nor U3129 (N_3129,N_1172,N_627);
nand U3130 (N_3130,N_539,N_1614);
nand U3131 (N_3131,N_92,N_436);
nand U3132 (N_3132,N_1584,N_1563);
or U3133 (N_3133,N_110,N_490);
xnor U3134 (N_3134,N_1429,N_799);
xnor U3135 (N_3135,N_226,N_563);
or U3136 (N_3136,N_198,N_80);
nor U3137 (N_3137,N_1538,N_767);
xor U3138 (N_3138,N_920,N_1376);
xor U3139 (N_3139,N_781,N_1083);
and U3140 (N_3140,N_417,N_1787);
or U3141 (N_3141,N_132,N_1500);
or U3142 (N_3142,N_179,N_632);
xor U3143 (N_3143,N_1651,N_187);
nor U3144 (N_3144,N_699,N_766);
nand U3145 (N_3145,N_1099,N_680);
or U3146 (N_3146,N_371,N_1730);
and U3147 (N_3147,N_917,N_1493);
nor U3148 (N_3148,N_771,N_1664);
and U3149 (N_3149,N_1639,N_883);
xor U3150 (N_3150,N_1699,N_66);
xnor U3151 (N_3151,N_1194,N_1599);
and U3152 (N_3152,N_330,N_1469);
xnor U3153 (N_3153,N_844,N_127);
or U3154 (N_3154,N_1487,N_1494);
nand U3155 (N_3155,N_526,N_1239);
and U3156 (N_3156,N_448,N_1156);
nor U3157 (N_3157,N_715,N_1963);
nor U3158 (N_3158,N_1171,N_379);
nor U3159 (N_3159,N_902,N_679);
nor U3160 (N_3160,N_623,N_830);
xor U3161 (N_3161,N_1205,N_1831);
xor U3162 (N_3162,N_144,N_1212);
or U3163 (N_3163,N_1205,N_1801);
nor U3164 (N_3164,N_90,N_595);
nand U3165 (N_3165,N_1558,N_1764);
nor U3166 (N_3166,N_383,N_823);
nor U3167 (N_3167,N_1443,N_609);
xnor U3168 (N_3168,N_550,N_1008);
nand U3169 (N_3169,N_229,N_1173);
nor U3170 (N_3170,N_1477,N_19);
nor U3171 (N_3171,N_1556,N_1858);
or U3172 (N_3172,N_1036,N_1333);
nor U3173 (N_3173,N_1104,N_316);
xor U3174 (N_3174,N_555,N_1672);
xor U3175 (N_3175,N_1270,N_352);
nor U3176 (N_3176,N_891,N_1573);
xnor U3177 (N_3177,N_214,N_1734);
nand U3178 (N_3178,N_946,N_941);
nor U3179 (N_3179,N_504,N_726);
or U3180 (N_3180,N_839,N_1991);
xnor U3181 (N_3181,N_1928,N_1504);
nor U3182 (N_3182,N_1208,N_928);
nor U3183 (N_3183,N_1847,N_1999);
or U3184 (N_3184,N_1748,N_198);
and U3185 (N_3185,N_86,N_1760);
and U3186 (N_3186,N_186,N_397);
nand U3187 (N_3187,N_1708,N_940);
nor U3188 (N_3188,N_1708,N_944);
nor U3189 (N_3189,N_385,N_325);
nor U3190 (N_3190,N_361,N_1359);
nand U3191 (N_3191,N_1016,N_221);
nor U3192 (N_3192,N_863,N_669);
nand U3193 (N_3193,N_1246,N_1709);
nand U3194 (N_3194,N_383,N_713);
nand U3195 (N_3195,N_1736,N_1732);
and U3196 (N_3196,N_294,N_911);
xnor U3197 (N_3197,N_250,N_1832);
and U3198 (N_3198,N_714,N_53);
or U3199 (N_3199,N_1192,N_254);
xor U3200 (N_3200,N_456,N_165);
nor U3201 (N_3201,N_731,N_1065);
and U3202 (N_3202,N_1589,N_1403);
nand U3203 (N_3203,N_1967,N_1501);
xor U3204 (N_3204,N_1414,N_52);
nor U3205 (N_3205,N_1022,N_847);
nor U3206 (N_3206,N_133,N_491);
nor U3207 (N_3207,N_992,N_1933);
nand U3208 (N_3208,N_1315,N_1493);
nor U3209 (N_3209,N_1816,N_1503);
and U3210 (N_3210,N_1113,N_1514);
nand U3211 (N_3211,N_1079,N_298);
nor U3212 (N_3212,N_1927,N_663);
nand U3213 (N_3213,N_773,N_1050);
nand U3214 (N_3214,N_552,N_730);
or U3215 (N_3215,N_683,N_1350);
or U3216 (N_3216,N_245,N_1515);
nand U3217 (N_3217,N_1750,N_1045);
xor U3218 (N_3218,N_625,N_677);
or U3219 (N_3219,N_223,N_988);
and U3220 (N_3220,N_1096,N_619);
nand U3221 (N_3221,N_1284,N_1189);
or U3222 (N_3222,N_1875,N_358);
or U3223 (N_3223,N_407,N_986);
xor U3224 (N_3224,N_1846,N_1713);
and U3225 (N_3225,N_189,N_921);
and U3226 (N_3226,N_1997,N_195);
nand U3227 (N_3227,N_342,N_426);
nand U3228 (N_3228,N_518,N_1592);
nor U3229 (N_3229,N_1713,N_369);
xor U3230 (N_3230,N_1576,N_742);
nand U3231 (N_3231,N_958,N_165);
nor U3232 (N_3232,N_483,N_853);
and U3233 (N_3233,N_1460,N_1092);
xnor U3234 (N_3234,N_990,N_1014);
nor U3235 (N_3235,N_1854,N_1324);
nor U3236 (N_3236,N_1285,N_1635);
xor U3237 (N_3237,N_336,N_1119);
nor U3238 (N_3238,N_602,N_1375);
nand U3239 (N_3239,N_404,N_851);
nor U3240 (N_3240,N_718,N_1507);
xnor U3241 (N_3241,N_1533,N_227);
nand U3242 (N_3242,N_575,N_75);
nand U3243 (N_3243,N_772,N_1835);
or U3244 (N_3244,N_1034,N_1054);
xor U3245 (N_3245,N_1951,N_1449);
nand U3246 (N_3246,N_1925,N_1135);
nor U3247 (N_3247,N_594,N_778);
and U3248 (N_3248,N_1008,N_55);
or U3249 (N_3249,N_273,N_733);
xor U3250 (N_3250,N_938,N_1307);
nor U3251 (N_3251,N_378,N_984);
or U3252 (N_3252,N_1364,N_255);
or U3253 (N_3253,N_1370,N_720);
nand U3254 (N_3254,N_1520,N_305);
or U3255 (N_3255,N_272,N_317);
xnor U3256 (N_3256,N_585,N_1897);
nor U3257 (N_3257,N_1703,N_1994);
nand U3258 (N_3258,N_1822,N_1098);
and U3259 (N_3259,N_1205,N_1730);
nand U3260 (N_3260,N_1978,N_764);
xnor U3261 (N_3261,N_1831,N_1034);
and U3262 (N_3262,N_1614,N_1132);
or U3263 (N_3263,N_1598,N_1705);
nand U3264 (N_3264,N_272,N_618);
nand U3265 (N_3265,N_270,N_887);
nor U3266 (N_3266,N_598,N_56);
or U3267 (N_3267,N_46,N_1971);
nor U3268 (N_3268,N_611,N_617);
or U3269 (N_3269,N_1364,N_750);
or U3270 (N_3270,N_1475,N_1088);
or U3271 (N_3271,N_620,N_107);
nand U3272 (N_3272,N_1196,N_864);
xnor U3273 (N_3273,N_984,N_1869);
or U3274 (N_3274,N_491,N_690);
and U3275 (N_3275,N_1739,N_849);
nor U3276 (N_3276,N_1827,N_1321);
and U3277 (N_3277,N_1430,N_661);
nor U3278 (N_3278,N_284,N_713);
or U3279 (N_3279,N_862,N_1505);
nand U3280 (N_3280,N_1759,N_1715);
or U3281 (N_3281,N_1608,N_1311);
nor U3282 (N_3282,N_712,N_1633);
or U3283 (N_3283,N_851,N_994);
nand U3284 (N_3284,N_1168,N_764);
nor U3285 (N_3285,N_1072,N_1316);
or U3286 (N_3286,N_1346,N_1758);
xnor U3287 (N_3287,N_1688,N_840);
nor U3288 (N_3288,N_1283,N_1883);
nand U3289 (N_3289,N_1957,N_1891);
nand U3290 (N_3290,N_1495,N_109);
nand U3291 (N_3291,N_651,N_1756);
nand U3292 (N_3292,N_1150,N_1196);
xor U3293 (N_3293,N_314,N_960);
or U3294 (N_3294,N_1043,N_1136);
xnor U3295 (N_3295,N_370,N_1956);
or U3296 (N_3296,N_989,N_1001);
xor U3297 (N_3297,N_1444,N_964);
or U3298 (N_3298,N_297,N_679);
nor U3299 (N_3299,N_1416,N_860);
nor U3300 (N_3300,N_1777,N_527);
and U3301 (N_3301,N_611,N_422);
nor U3302 (N_3302,N_1743,N_723);
nor U3303 (N_3303,N_1574,N_291);
xor U3304 (N_3304,N_119,N_1153);
and U3305 (N_3305,N_1671,N_1348);
nor U3306 (N_3306,N_1736,N_1563);
and U3307 (N_3307,N_517,N_1504);
nor U3308 (N_3308,N_1422,N_1301);
and U3309 (N_3309,N_446,N_1957);
nor U3310 (N_3310,N_981,N_1000);
nor U3311 (N_3311,N_1809,N_1048);
nor U3312 (N_3312,N_174,N_439);
and U3313 (N_3313,N_98,N_63);
xnor U3314 (N_3314,N_939,N_1766);
nor U3315 (N_3315,N_990,N_1506);
nor U3316 (N_3316,N_1375,N_1236);
xnor U3317 (N_3317,N_1238,N_1308);
nor U3318 (N_3318,N_1518,N_969);
nand U3319 (N_3319,N_776,N_472);
or U3320 (N_3320,N_1624,N_1612);
and U3321 (N_3321,N_408,N_499);
and U3322 (N_3322,N_1649,N_1893);
and U3323 (N_3323,N_738,N_1879);
nand U3324 (N_3324,N_1303,N_1410);
nand U3325 (N_3325,N_1635,N_1646);
nand U3326 (N_3326,N_1096,N_522);
and U3327 (N_3327,N_1993,N_953);
or U3328 (N_3328,N_61,N_628);
xor U3329 (N_3329,N_1020,N_302);
xor U3330 (N_3330,N_951,N_123);
nand U3331 (N_3331,N_852,N_1088);
xor U3332 (N_3332,N_1422,N_1359);
nand U3333 (N_3333,N_743,N_1533);
xor U3334 (N_3334,N_165,N_1429);
or U3335 (N_3335,N_1120,N_1317);
nand U3336 (N_3336,N_610,N_842);
nor U3337 (N_3337,N_1677,N_1835);
or U3338 (N_3338,N_584,N_132);
nand U3339 (N_3339,N_831,N_729);
xnor U3340 (N_3340,N_55,N_1866);
and U3341 (N_3341,N_559,N_227);
and U3342 (N_3342,N_1686,N_929);
or U3343 (N_3343,N_1206,N_1526);
or U3344 (N_3344,N_1071,N_276);
xor U3345 (N_3345,N_1135,N_1222);
or U3346 (N_3346,N_1715,N_1186);
nand U3347 (N_3347,N_161,N_54);
nor U3348 (N_3348,N_1513,N_314);
nand U3349 (N_3349,N_650,N_331);
nor U3350 (N_3350,N_916,N_1576);
xnor U3351 (N_3351,N_1460,N_827);
nand U3352 (N_3352,N_1769,N_278);
xor U3353 (N_3353,N_1880,N_112);
and U3354 (N_3354,N_1385,N_1734);
or U3355 (N_3355,N_333,N_883);
or U3356 (N_3356,N_1520,N_1066);
or U3357 (N_3357,N_1357,N_1316);
xor U3358 (N_3358,N_134,N_195);
xor U3359 (N_3359,N_1239,N_388);
nor U3360 (N_3360,N_973,N_1094);
or U3361 (N_3361,N_1709,N_905);
xnor U3362 (N_3362,N_1926,N_840);
nand U3363 (N_3363,N_1335,N_207);
xnor U3364 (N_3364,N_6,N_880);
and U3365 (N_3365,N_1265,N_945);
or U3366 (N_3366,N_1443,N_1582);
nor U3367 (N_3367,N_634,N_968);
or U3368 (N_3368,N_1903,N_396);
nand U3369 (N_3369,N_1578,N_652);
and U3370 (N_3370,N_1418,N_1173);
xnor U3371 (N_3371,N_183,N_866);
nand U3372 (N_3372,N_532,N_1154);
and U3373 (N_3373,N_838,N_1599);
nor U3374 (N_3374,N_1852,N_469);
and U3375 (N_3375,N_1413,N_440);
nor U3376 (N_3376,N_1744,N_1296);
xor U3377 (N_3377,N_1848,N_1023);
or U3378 (N_3378,N_1089,N_191);
and U3379 (N_3379,N_1315,N_1208);
nor U3380 (N_3380,N_1450,N_1570);
and U3381 (N_3381,N_1603,N_1100);
or U3382 (N_3382,N_1155,N_1895);
and U3383 (N_3383,N_1626,N_1253);
and U3384 (N_3384,N_316,N_259);
or U3385 (N_3385,N_169,N_1008);
nand U3386 (N_3386,N_1355,N_87);
or U3387 (N_3387,N_189,N_967);
or U3388 (N_3388,N_384,N_898);
nor U3389 (N_3389,N_1385,N_289);
or U3390 (N_3390,N_1384,N_1173);
nand U3391 (N_3391,N_482,N_471);
and U3392 (N_3392,N_252,N_837);
nor U3393 (N_3393,N_1900,N_132);
nand U3394 (N_3394,N_686,N_962);
nand U3395 (N_3395,N_83,N_514);
and U3396 (N_3396,N_11,N_1198);
and U3397 (N_3397,N_1549,N_1060);
or U3398 (N_3398,N_1791,N_673);
or U3399 (N_3399,N_1005,N_1137);
or U3400 (N_3400,N_1066,N_1713);
or U3401 (N_3401,N_604,N_638);
xnor U3402 (N_3402,N_1913,N_1908);
nor U3403 (N_3403,N_277,N_399);
xor U3404 (N_3404,N_1043,N_1947);
or U3405 (N_3405,N_779,N_1588);
xnor U3406 (N_3406,N_1980,N_962);
or U3407 (N_3407,N_1590,N_638);
nor U3408 (N_3408,N_1585,N_1148);
xnor U3409 (N_3409,N_629,N_1118);
or U3410 (N_3410,N_1065,N_792);
nor U3411 (N_3411,N_741,N_1412);
and U3412 (N_3412,N_1337,N_535);
nand U3413 (N_3413,N_1346,N_1302);
or U3414 (N_3414,N_1201,N_1677);
and U3415 (N_3415,N_1419,N_747);
nand U3416 (N_3416,N_671,N_1320);
or U3417 (N_3417,N_695,N_259);
and U3418 (N_3418,N_1695,N_1170);
nor U3419 (N_3419,N_562,N_1515);
or U3420 (N_3420,N_493,N_1825);
xnor U3421 (N_3421,N_1827,N_1601);
xnor U3422 (N_3422,N_1525,N_44);
nor U3423 (N_3423,N_1808,N_1588);
and U3424 (N_3424,N_1644,N_1682);
and U3425 (N_3425,N_359,N_1293);
and U3426 (N_3426,N_591,N_265);
xnor U3427 (N_3427,N_1300,N_301);
or U3428 (N_3428,N_1761,N_1664);
or U3429 (N_3429,N_145,N_221);
and U3430 (N_3430,N_1208,N_402);
nand U3431 (N_3431,N_785,N_1624);
or U3432 (N_3432,N_619,N_1727);
and U3433 (N_3433,N_1638,N_244);
xor U3434 (N_3434,N_1288,N_981);
xnor U3435 (N_3435,N_1506,N_619);
and U3436 (N_3436,N_1173,N_826);
nor U3437 (N_3437,N_152,N_229);
xor U3438 (N_3438,N_313,N_889);
and U3439 (N_3439,N_66,N_101);
or U3440 (N_3440,N_477,N_1858);
nand U3441 (N_3441,N_251,N_920);
or U3442 (N_3442,N_786,N_312);
and U3443 (N_3443,N_764,N_70);
nor U3444 (N_3444,N_387,N_497);
or U3445 (N_3445,N_843,N_477);
nand U3446 (N_3446,N_1183,N_1773);
nor U3447 (N_3447,N_764,N_842);
or U3448 (N_3448,N_1235,N_155);
nand U3449 (N_3449,N_1459,N_1354);
nand U3450 (N_3450,N_92,N_1285);
nor U3451 (N_3451,N_310,N_991);
xor U3452 (N_3452,N_847,N_1500);
nor U3453 (N_3453,N_1016,N_938);
nand U3454 (N_3454,N_1383,N_771);
and U3455 (N_3455,N_1732,N_1234);
xor U3456 (N_3456,N_815,N_866);
and U3457 (N_3457,N_1289,N_248);
xnor U3458 (N_3458,N_540,N_1799);
and U3459 (N_3459,N_234,N_402);
or U3460 (N_3460,N_716,N_352);
or U3461 (N_3461,N_286,N_1169);
and U3462 (N_3462,N_1282,N_489);
nand U3463 (N_3463,N_399,N_5);
or U3464 (N_3464,N_1026,N_433);
xnor U3465 (N_3465,N_504,N_1206);
or U3466 (N_3466,N_1692,N_1869);
nor U3467 (N_3467,N_894,N_1173);
or U3468 (N_3468,N_845,N_637);
nand U3469 (N_3469,N_926,N_708);
nand U3470 (N_3470,N_722,N_1621);
nor U3471 (N_3471,N_875,N_1814);
or U3472 (N_3472,N_1215,N_1360);
and U3473 (N_3473,N_496,N_1440);
and U3474 (N_3474,N_1789,N_413);
nand U3475 (N_3475,N_1672,N_1258);
nor U3476 (N_3476,N_1054,N_535);
nand U3477 (N_3477,N_1807,N_1108);
xor U3478 (N_3478,N_1268,N_784);
nand U3479 (N_3479,N_848,N_1198);
nor U3480 (N_3480,N_1971,N_1549);
xnor U3481 (N_3481,N_1832,N_1974);
nor U3482 (N_3482,N_1177,N_143);
or U3483 (N_3483,N_485,N_221);
nand U3484 (N_3484,N_720,N_478);
or U3485 (N_3485,N_735,N_1000);
and U3486 (N_3486,N_1583,N_154);
xnor U3487 (N_3487,N_608,N_1822);
and U3488 (N_3488,N_596,N_924);
and U3489 (N_3489,N_1127,N_101);
and U3490 (N_3490,N_877,N_437);
nand U3491 (N_3491,N_1714,N_617);
nor U3492 (N_3492,N_415,N_540);
nand U3493 (N_3493,N_1362,N_1561);
nor U3494 (N_3494,N_96,N_275);
nor U3495 (N_3495,N_891,N_1937);
and U3496 (N_3496,N_61,N_812);
nand U3497 (N_3497,N_748,N_975);
nor U3498 (N_3498,N_1872,N_901);
nand U3499 (N_3499,N_103,N_1014);
nand U3500 (N_3500,N_370,N_1845);
or U3501 (N_3501,N_1924,N_926);
or U3502 (N_3502,N_1382,N_116);
or U3503 (N_3503,N_1045,N_1475);
xnor U3504 (N_3504,N_176,N_1421);
nor U3505 (N_3505,N_984,N_733);
nor U3506 (N_3506,N_1740,N_1172);
nand U3507 (N_3507,N_1698,N_406);
and U3508 (N_3508,N_1757,N_1798);
and U3509 (N_3509,N_285,N_1765);
and U3510 (N_3510,N_1650,N_310);
and U3511 (N_3511,N_1682,N_1190);
and U3512 (N_3512,N_1429,N_1596);
or U3513 (N_3513,N_1317,N_992);
xor U3514 (N_3514,N_1918,N_691);
nand U3515 (N_3515,N_1664,N_554);
and U3516 (N_3516,N_870,N_443);
and U3517 (N_3517,N_967,N_1134);
xnor U3518 (N_3518,N_1014,N_1365);
or U3519 (N_3519,N_217,N_554);
and U3520 (N_3520,N_1850,N_1332);
nor U3521 (N_3521,N_346,N_217);
nor U3522 (N_3522,N_1789,N_181);
xor U3523 (N_3523,N_1803,N_181);
nand U3524 (N_3524,N_1178,N_843);
xor U3525 (N_3525,N_1546,N_426);
or U3526 (N_3526,N_1148,N_73);
nand U3527 (N_3527,N_926,N_623);
and U3528 (N_3528,N_1244,N_280);
xor U3529 (N_3529,N_1479,N_292);
xnor U3530 (N_3530,N_1918,N_395);
xor U3531 (N_3531,N_923,N_1242);
or U3532 (N_3532,N_1159,N_1916);
or U3533 (N_3533,N_1414,N_600);
nor U3534 (N_3534,N_595,N_1519);
xnor U3535 (N_3535,N_704,N_237);
nand U3536 (N_3536,N_619,N_1663);
nor U3537 (N_3537,N_1774,N_847);
xnor U3538 (N_3538,N_50,N_284);
nor U3539 (N_3539,N_45,N_1611);
nor U3540 (N_3540,N_1336,N_540);
nor U3541 (N_3541,N_1421,N_1333);
or U3542 (N_3542,N_1061,N_1700);
and U3543 (N_3543,N_242,N_1400);
or U3544 (N_3544,N_1164,N_1064);
and U3545 (N_3545,N_1191,N_268);
nand U3546 (N_3546,N_1569,N_369);
nor U3547 (N_3547,N_1324,N_29);
and U3548 (N_3548,N_19,N_1935);
and U3549 (N_3549,N_1921,N_1956);
and U3550 (N_3550,N_627,N_1415);
nor U3551 (N_3551,N_1558,N_1597);
nand U3552 (N_3552,N_209,N_358);
and U3553 (N_3553,N_219,N_1584);
or U3554 (N_3554,N_1853,N_1152);
and U3555 (N_3555,N_1228,N_326);
or U3556 (N_3556,N_761,N_1050);
nand U3557 (N_3557,N_1023,N_149);
or U3558 (N_3558,N_1689,N_1285);
nand U3559 (N_3559,N_1814,N_333);
xor U3560 (N_3560,N_1127,N_1472);
or U3561 (N_3561,N_1955,N_1052);
nor U3562 (N_3562,N_1668,N_405);
or U3563 (N_3563,N_1308,N_1983);
xor U3564 (N_3564,N_591,N_443);
nand U3565 (N_3565,N_772,N_1013);
nor U3566 (N_3566,N_1454,N_1453);
xnor U3567 (N_3567,N_24,N_1162);
nand U3568 (N_3568,N_1229,N_380);
xnor U3569 (N_3569,N_1433,N_1801);
or U3570 (N_3570,N_1983,N_1520);
xnor U3571 (N_3571,N_148,N_706);
xnor U3572 (N_3572,N_1344,N_1642);
or U3573 (N_3573,N_1017,N_1384);
nor U3574 (N_3574,N_1349,N_1730);
xor U3575 (N_3575,N_214,N_662);
nor U3576 (N_3576,N_1774,N_482);
nor U3577 (N_3577,N_1601,N_854);
nor U3578 (N_3578,N_455,N_4);
nor U3579 (N_3579,N_370,N_251);
xnor U3580 (N_3580,N_989,N_81);
nor U3581 (N_3581,N_1482,N_1018);
nor U3582 (N_3582,N_393,N_132);
nand U3583 (N_3583,N_1045,N_307);
nor U3584 (N_3584,N_1903,N_500);
nor U3585 (N_3585,N_324,N_810);
or U3586 (N_3586,N_922,N_645);
nand U3587 (N_3587,N_1428,N_850);
and U3588 (N_3588,N_862,N_1498);
nor U3589 (N_3589,N_1803,N_1475);
and U3590 (N_3590,N_1410,N_35);
or U3591 (N_3591,N_84,N_371);
nor U3592 (N_3592,N_448,N_398);
and U3593 (N_3593,N_1170,N_258);
nor U3594 (N_3594,N_760,N_1458);
xor U3595 (N_3595,N_188,N_1746);
and U3596 (N_3596,N_308,N_554);
nand U3597 (N_3597,N_510,N_1364);
xor U3598 (N_3598,N_788,N_893);
nand U3599 (N_3599,N_821,N_801);
nand U3600 (N_3600,N_1967,N_351);
and U3601 (N_3601,N_655,N_1015);
and U3602 (N_3602,N_511,N_591);
or U3603 (N_3603,N_621,N_1178);
nor U3604 (N_3604,N_60,N_1654);
and U3605 (N_3605,N_395,N_789);
xnor U3606 (N_3606,N_1041,N_1161);
xnor U3607 (N_3607,N_175,N_15);
nand U3608 (N_3608,N_1830,N_916);
nor U3609 (N_3609,N_634,N_963);
and U3610 (N_3610,N_766,N_1031);
xor U3611 (N_3611,N_859,N_541);
nor U3612 (N_3612,N_1822,N_1067);
nor U3613 (N_3613,N_1004,N_1287);
or U3614 (N_3614,N_1655,N_1832);
nand U3615 (N_3615,N_621,N_1080);
nor U3616 (N_3616,N_182,N_499);
or U3617 (N_3617,N_179,N_1681);
nor U3618 (N_3618,N_324,N_870);
nor U3619 (N_3619,N_1039,N_1189);
nand U3620 (N_3620,N_743,N_389);
nor U3621 (N_3621,N_366,N_806);
nand U3622 (N_3622,N_963,N_1296);
and U3623 (N_3623,N_356,N_1698);
and U3624 (N_3624,N_540,N_625);
nand U3625 (N_3625,N_1315,N_1878);
nand U3626 (N_3626,N_357,N_1091);
nand U3627 (N_3627,N_75,N_1771);
or U3628 (N_3628,N_500,N_1121);
nand U3629 (N_3629,N_1685,N_474);
or U3630 (N_3630,N_1730,N_865);
nand U3631 (N_3631,N_1895,N_224);
nor U3632 (N_3632,N_1903,N_330);
nor U3633 (N_3633,N_830,N_946);
and U3634 (N_3634,N_1811,N_1812);
nor U3635 (N_3635,N_135,N_1525);
nor U3636 (N_3636,N_12,N_767);
xor U3637 (N_3637,N_981,N_1476);
or U3638 (N_3638,N_1293,N_632);
and U3639 (N_3639,N_1346,N_422);
nor U3640 (N_3640,N_1581,N_1547);
and U3641 (N_3641,N_1752,N_525);
xor U3642 (N_3642,N_1952,N_621);
xnor U3643 (N_3643,N_1085,N_918);
xor U3644 (N_3644,N_27,N_459);
nor U3645 (N_3645,N_633,N_1875);
nand U3646 (N_3646,N_814,N_1077);
nand U3647 (N_3647,N_1902,N_1006);
or U3648 (N_3648,N_1787,N_475);
xnor U3649 (N_3649,N_1948,N_1990);
or U3650 (N_3650,N_1320,N_784);
nand U3651 (N_3651,N_1655,N_532);
xor U3652 (N_3652,N_788,N_1986);
xnor U3653 (N_3653,N_68,N_218);
nor U3654 (N_3654,N_1796,N_1059);
or U3655 (N_3655,N_191,N_232);
nand U3656 (N_3656,N_1875,N_1473);
or U3657 (N_3657,N_1351,N_192);
nand U3658 (N_3658,N_1572,N_120);
xor U3659 (N_3659,N_513,N_1623);
xnor U3660 (N_3660,N_1481,N_639);
nor U3661 (N_3661,N_1230,N_955);
or U3662 (N_3662,N_248,N_1312);
nor U3663 (N_3663,N_1093,N_834);
or U3664 (N_3664,N_1202,N_986);
nand U3665 (N_3665,N_1847,N_382);
nor U3666 (N_3666,N_1597,N_1162);
or U3667 (N_3667,N_1563,N_611);
and U3668 (N_3668,N_1752,N_497);
and U3669 (N_3669,N_1310,N_1327);
and U3670 (N_3670,N_1713,N_1987);
nand U3671 (N_3671,N_1052,N_1523);
nor U3672 (N_3672,N_562,N_229);
or U3673 (N_3673,N_1108,N_1572);
nor U3674 (N_3674,N_985,N_296);
or U3675 (N_3675,N_882,N_149);
nand U3676 (N_3676,N_366,N_1861);
or U3677 (N_3677,N_1999,N_436);
and U3678 (N_3678,N_1130,N_405);
nor U3679 (N_3679,N_1608,N_811);
or U3680 (N_3680,N_329,N_87);
or U3681 (N_3681,N_755,N_567);
nor U3682 (N_3682,N_1984,N_875);
nand U3683 (N_3683,N_625,N_491);
xnor U3684 (N_3684,N_1173,N_622);
or U3685 (N_3685,N_441,N_596);
or U3686 (N_3686,N_618,N_670);
and U3687 (N_3687,N_1019,N_339);
xnor U3688 (N_3688,N_1246,N_1017);
nor U3689 (N_3689,N_946,N_945);
nand U3690 (N_3690,N_436,N_1739);
and U3691 (N_3691,N_1565,N_1470);
nor U3692 (N_3692,N_879,N_366);
or U3693 (N_3693,N_1188,N_671);
nand U3694 (N_3694,N_1459,N_321);
or U3695 (N_3695,N_799,N_44);
nor U3696 (N_3696,N_1223,N_279);
xnor U3697 (N_3697,N_1029,N_1069);
xnor U3698 (N_3698,N_177,N_1719);
nor U3699 (N_3699,N_1561,N_1435);
nand U3700 (N_3700,N_1459,N_962);
nand U3701 (N_3701,N_1771,N_1237);
nor U3702 (N_3702,N_481,N_1745);
nand U3703 (N_3703,N_424,N_937);
nand U3704 (N_3704,N_1795,N_1642);
nand U3705 (N_3705,N_856,N_995);
xor U3706 (N_3706,N_171,N_1706);
nor U3707 (N_3707,N_693,N_1484);
nand U3708 (N_3708,N_456,N_1456);
and U3709 (N_3709,N_179,N_390);
and U3710 (N_3710,N_1323,N_1343);
nor U3711 (N_3711,N_1482,N_1951);
nor U3712 (N_3712,N_1357,N_75);
nand U3713 (N_3713,N_1508,N_485);
xnor U3714 (N_3714,N_1708,N_482);
nand U3715 (N_3715,N_1592,N_1662);
xor U3716 (N_3716,N_1999,N_475);
xor U3717 (N_3717,N_818,N_1369);
nand U3718 (N_3718,N_1692,N_1065);
nor U3719 (N_3719,N_714,N_1995);
and U3720 (N_3720,N_366,N_1078);
nand U3721 (N_3721,N_1404,N_1524);
or U3722 (N_3722,N_1204,N_65);
and U3723 (N_3723,N_1984,N_97);
nor U3724 (N_3724,N_1210,N_731);
nor U3725 (N_3725,N_485,N_1849);
nand U3726 (N_3726,N_237,N_560);
nand U3727 (N_3727,N_1111,N_1508);
nor U3728 (N_3728,N_716,N_938);
or U3729 (N_3729,N_849,N_552);
nor U3730 (N_3730,N_303,N_1824);
xnor U3731 (N_3731,N_1301,N_1580);
xor U3732 (N_3732,N_848,N_616);
or U3733 (N_3733,N_1693,N_1947);
or U3734 (N_3734,N_436,N_1969);
nor U3735 (N_3735,N_1330,N_1755);
and U3736 (N_3736,N_1110,N_325);
nand U3737 (N_3737,N_1308,N_853);
or U3738 (N_3738,N_1254,N_1812);
nor U3739 (N_3739,N_1602,N_1340);
or U3740 (N_3740,N_1996,N_858);
or U3741 (N_3741,N_1834,N_1122);
or U3742 (N_3742,N_1306,N_828);
nor U3743 (N_3743,N_1826,N_424);
xor U3744 (N_3744,N_1709,N_1895);
xnor U3745 (N_3745,N_294,N_1989);
xor U3746 (N_3746,N_587,N_61);
or U3747 (N_3747,N_880,N_1292);
nand U3748 (N_3748,N_170,N_696);
and U3749 (N_3749,N_1053,N_538);
nand U3750 (N_3750,N_1825,N_841);
and U3751 (N_3751,N_637,N_91);
or U3752 (N_3752,N_431,N_613);
or U3753 (N_3753,N_897,N_922);
or U3754 (N_3754,N_1953,N_330);
nand U3755 (N_3755,N_555,N_139);
and U3756 (N_3756,N_1318,N_1913);
and U3757 (N_3757,N_985,N_1793);
nor U3758 (N_3758,N_180,N_1723);
xnor U3759 (N_3759,N_457,N_839);
nor U3760 (N_3760,N_1965,N_776);
or U3761 (N_3761,N_506,N_473);
and U3762 (N_3762,N_947,N_540);
and U3763 (N_3763,N_1651,N_314);
or U3764 (N_3764,N_988,N_447);
or U3765 (N_3765,N_1256,N_1008);
xnor U3766 (N_3766,N_1288,N_1417);
nor U3767 (N_3767,N_197,N_213);
xnor U3768 (N_3768,N_452,N_432);
nor U3769 (N_3769,N_616,N_492);
nand U3770 (N_3770,N_1026,N_1014);
nor U3771 (N_3771,N_34,N_676);
and U3772 (N_3772,N_1243,N_1526);
xnor U3773 (N_3773,N_1966,N_1638);
and U3774 (N_3774,N_1026,N_309);
or U3775 (N_3775,N_1777,N_1316);
nor U3776 (N_3776,N_1659,N_1733);
and U3777 (N_3777,N_1295,N_898);
xor U3778 (N_3778,N_261,N_896);
or U3779 (N_3779,N_1651,N_1243);
xnor U3780 (N_3780,N_384,N_1746);
and U3781 (N_3781,N_487,N_1241);
and U3782 (N_3782,N_838,N_1132);
xnor U3783 (N_3783,N_363,N_1343);
or U3784 (N_3784,N_1260,N_936);
or U3785 (N_3785,N_88,N_529);
xnor U3786 (N_3786,N_1866,N_537);
nand U3787 (N_3787,N_432,N_564);
nand U3788 (N_3788,N_391,N_265);
nor U3789 (N_3789,N_571,N_1853);
nor U3790 (N_3790,N_321,N_115);
or U3791 (N_3791,N_20,N_1822);
and U3792 (N_3792,N_921,N_151);
or U3793 (N_3793,N_881,N_249);
xor U3794 (N_3794,N_1394,N_1439);
xnor U3795 (N_3795,N_736,N_959);
or U3796 (N_3796,N_150,N_215);
nand U3797 (N_3797,N_739,N_810);
nand U3798 (N_3798,N_368,N_259);
or U3799 (N_3799,N_938,N_956);
xnor U3800 (N_3800,N_995,N_1861);
or U3801 (N_3801,N_763,N_1799);
nor U3802 (N_3802,N_523,N_1547);
xor U3803 (N_3803,N_450,N_1585);
nor U3804 (N_3804,N_1090,N_1453);
xnor U3805 (N_3805,N_1835,N_657);
nand U3806 (N_3806,N_132,N_1326);
or U3807 (N_3807,N_445,N_1839);
xnor U3808 (N_3808,N_63,N_358);
and U3809 (N_3809,N_1305,N_821);
or U3810 (N_3810,N_724,N_181);
xnor U3811 (N_3811,N_1148,N_1430);
nor U3812 (N_3812,N_98,N_622);
or U3813 (N_3813,N_932,N_695);
or U3814 (N_3814,N_790,N_103);
and U3815 (N_3815,N_979,N_279);
and U3816 (N_3816,N_1291,N_1823);
and U3817 (N_3817,N_555,N_1361);
nor U3818 (N_3818,N_1258,N_1416);
nand U3819 (N_3819,N_213,N_381);
and U3820 (N_3820,N_1633,N_23);
or U3821 (N_3821,N_912,N_784);
nand U3822 (N_3822,N_1287,N_731);
and U3823 (N_3823,N_166,N_1483);
and U3824 (N_3824,N_844,N_1465);
or U3825 (N_3825,N_587,N_1215);
or U3826 (N_3826,N_555,N_161);
xnor U3827 (N_3827,N_416,N_285);
and U3828 (N_3828,N_112,N_747);
nor U3829 (N_3829,N_1474,N_166);
nand U3830 (N_3830,N_1845,N_1952);
nor U3831 (N_3831,N_1319,N_1901);
xnor U3832 (N_3832,N_503,N_844);
xnor U3833 (N_3833,N_130,N_1761);
xor U3834 (N_3834,N_420,N_1211);
or U3835 (N_3835,N_1113,N_1675);
or U3836 (N_3836,N_589,N_1354);
xnor U3837 (N_3837,N_1323,N_1340);
xnor U3838 (N_3838,N_1031,N_1602);
nor U3839 (N_3839,N_1544,N_1757);
nor U3840 (N_3840,N_855,N_255);
nand U3841 (N_3841,N_256,N_173);
nor U3842 (N_3842,N_105,N_1477);
and U3843 (N_3843,N_1881,N_1957);
or U3844 (N_3844,N_178,N_354);
and U3845 (N_3845,N_729,N_903);
nor U3846 (N_3846,N_255,N_1222);
nor U3847 (N_3847,N_25,N_1447);
xnor U3848 (N_3848,N_1820,N_1848);
and U3849 (N_3849,N_324,N_1378);
nand U3850 (N_3850,N_1251,N_1305);
and U3851 (N_3851,N_1728,N_1827);
nor U3852 (N_3852,N_1744,N_1785);
xor U3853 (N_3853,N_28,N_1156);
nor U3854 (N_3854,N_46,N_1785);
or U3855 (N_3855,N_1172,N_1168);
nor U3856 (N_3856,N_917,N_185);
xor U3857 (N_3857,N_1110,N_1456);
nand U3858 (N_3858,N_1805,N_1825);
or U3859 (N_3859,N_1025,N_1872);
nand U3860 (N_3860,N_499,N_1636);
nor U3861 (N_3861,N_734,N_161);
and U3862 (N_3862,N_697,N_748);
and U3863 (N_3863,N_667,N_819);
or U3864 (N_3864,N_227,N_349);
or U3865 (N_3865,N_389,N_621);
nand U3866 (N_3866,N_1224,N_237);
or U3867 (N_3867,N_1430,N_1475);
nor U3868 (N_3868,N_1023,N_267);
xnor U3869 (N_3869,N_1490,N_201);
and U3870 (N_3870,N_941,N_1089);
nand U3871 (N_3871,N_1170,N_457);
nor U3872 (N_3872,N_727,N_1027);
nor U3873 (N_3873,N_468,N_1457);
or U3874 (N_3874,N_449,N_59);
nor U3875 (N_3875,N_1089,N_518);
nand U3876 (N_3876,N_543,N_1924);
and U3877 (N_3877,N_1259,N_584);
xnor U3878 (N_3878,N_434,N_169);
nand U3879 (N_3879,N_353,N_254);
or U3880 (N_3880,N_149,N_850);
xnor U3881 (N_3881,N_1298,N_79);
nand U3882 (N_3882,N_1145,N_45);
nor U3883 (N_3883,N_1363,N_1136);
xor U3884 (N_3884,N_1920,N_78);
or U3885 (N_3885,N_295,N_1556);
and U3886 (N_3886,N_334,N_1996);
or U3887 (N_3887,N_479,N_1259);
and U3888 (N_3888,N_1149,N_65);
nor U3889 (N_3889,N_678,N_1753);
xor U3890 (N_3890,N_1173,N_814);
nand U3891 (N_3891,N_476,N_1074);
nor U3892 (N_3892,N_1727,N_534);
xor U3893 (N_3893,N_1261,N_413);
xor U3894 (N_3894,N_1602,N_1692);
nor U3895 (N_3895,N_989,N_719);
xnor U3896 (N_3896,N_1849,N_824);
and U3897 (N_3897,N_755,N_1911);
nand U3898 (N_3898,N_95,N_547);
nor U3899 (N_3899,N_1203,N_1286);
nand U3900 (N_3900,N_1579,N_1818);
nand U3901 (N_3901,N_1470,N_1130);
nor U3902 (N_3902,N_1662,N_1349);
xnor U3903 (N_3903,N_309,N_292);
nand U3904 (N_3904,N_1045,N_427);
and U3905 (N_3905,N_1727,N_894);
xnor U3906 (N_3906,N_1423,N_432);
nor U3907 (N_3907,N_1258,N_599);
nand U3908 (N_3908,N_423,N_607);
and U3909 (N_3909,N_888,N_1741);
or U3910 (N_3910,N_315,N_165);
and U3911 (N_3911,N_342,N_309);
xnor U3912 (N_3912,N_875,N_1620);
or U3913 (N_3913,N_1422,N_1314);
nand U3914 (N_3914,N_1354,N_1964);
and U3915 (N_3915,N_1538,N_1087);
xnor U3916 (N_3916,N_1963,N_1564);
nor U3917 (N_3917,N_1532,N_441);
or U3918 (N_3918,N_708,N_233);
or U3919 (N_3919,N_229,N_538);
xor U3920 (N_3920,N_278,N_661);
or U3921 (N_3921,N_1505,N_1500);
xor U3922 (N_3922,N_1485,N_1186);
nor U3923 (N_3923,N_654,N_524);
and U3924 (N_3924,N_829,N_1614);
and U3925 (N_3925,N_749,N_172);
xnor U3926 (N_3926,N_1740,N_100);
or U3927 (N_3927,N_440,N_1118);
nand U3928 (N_3928,N_1827,N_1428);
nand U3929 (N_3929,N_1529,N_1236);
or U3930 (N_3930,N_835,N_1502);
or U3931 (N_3931,N_826,N_1278);
and U3932 (N_3932,N_815,N_697);
or U3933 (N_3933,N_1730,N_823);
and U3934 (N_3934,N_937,N_185);
nand U3935 (N_3935,N_1759,N_1537);
or U3936 (N_3936,N_1757,N_1735);
nor U3937 (N_3937,N_966,N_1429);
nand U3938 (N_3938,N_1820,N_1054);
xor U3939 (N_3939,N_197,N_384);
nor U3940 (N_3940,N_748,N_1708);
or U3941 (N_3941,N_1104,N_110);
and U3942 (N_3942,N_1137,N_445);
or U3943 (N_3943,N_1837,N_1309);
nor U3944 (N_3944,N_1529,N_1686);
nand U3945 (N_3945,N_1627,N_226);
and U3946 (N_3946,N_1032,N_1357);
and U3947 (N_3947,N_1886,N_609);
nand U3948 (N_3948,N_710,N_967);
nor U3949 (N_3949,N_816,N_272);
xor U3950 (N_3950,N_448,N_1835);
and U3951 (N_3951,N_143,N_529);
or U3952 (N_3952,N_1048,N_1931);
or U3953 (N_3953,N_1413,N_252);
xor U3954 (N_3954,N_1645,N_174);
and U3955 (N_3955,N_126,N_330);
xnor U3956 (N_3956,N_682,N_351);
and U3957 (N_3957,N_1499,N_5);
xnor U3958 (N_3958,N_1736,N_431);
or U3959 (N_3959,N_1550,N_76);
nand U3960 (N_3960,N_408,N_1839);
nand U3961 (N_3961,N_993,N_1878);
nand U3962 (N_3962,N_1953,N_1637);
nand U3963 (N_3963,N_1024,N_1013);
or U3964 (N_3964,N_1080,N_227);
and U3965 (N_3965,N_1551,N_1707);
and U3966 (N_3966,N_270,N_1397);
and U3967 (N_3967,N_1575,N_1144);
nand U3968 (N_3968,N_590,N_1152);
nor U3969 (N_3969,N_1454,N_568);
nand U3970 (N_3970,N_5,N_289);
nand U3971 (N_3971,N_479,N_795);
and U3972 (N_3972,N_1382,N_1752);
nor U3973 (N_3973,N_14,N_1551);
and U3974 (N_3974,N_950,N_564);
and U3975 (N_3975,N_786,N_363);
nand U3976 (N_3976,N_334,N_205);
nand U3977 (N_3977,N_920,N_156);
nor U3978 (N_3978,N_604,N_1885);
or U3979 (N_3979,N_1736,N_1780);
nand U3980 (N_3980,N_1701,N_1930);
nor U3981 (N_3981,N_1609,N_1847);
and U3982 (N_3982,N_1629,N_228);
xor U3983 (N_3983,N_968,N_582);
nand U3984 (N_3984,N_519,N_335);
nand U3985 (N_3985,N_28,N_990);
nor U3986 (N_3986,N_723,N_1178);
xor U3987 (N_3987,N_1158,N_1251);
xor U3988 (N_3988,N_197,N_1442);
nor U3989 (N_3989,N_1526,N_1585);
xor U3990 (N_3990,N_1575,N_184);
nand U3991 (N_3991,N_1981,N_1626);
nand U3992 (N_3992,N_1079,N_1013);
or U3993 (N_3993,N_997,N_1646);
nor U3994 (N_3994,N_1891,N_1797);
nor U3995 (N_3995,N_1112,N_1841);
xnor U3996 (N_3996,N_1776,N_1685);
nand U3997 (N_3997,N_1864,N_563);
nor U3998 (N_3998,N_1679,N_287);
xnor U3999 (N_3999,N_107,N_1565);
nor U4000 (N_4000,N_2441,N_2391);
or U4001 (N_4001,N_3039,N_3250);
or U4002 (N_4002,N_3676,N_2621);
xor U4003 (N_4003,N_3218,N_2640);
xor U4004 (N_4004,N_3681,N_3663);
and U4005 (N_4005,N_3203,N_3683);
xor U4006 (N_4006,N_2458,N_2919);
or U4007 (N_4007,N_3343,N_2720);
or U4008 (N_4008,N_3712,N_3713);
or U4009 (N_4009,N_2547,N_2426);
or U4010 (N_4010,N_2428,N_2718);
nand U4011 (N_4011,N_3269,N_3767);
or U4012 (N_4012,N_3276,N_2339);
xnor U4013 (N_4013,N_2750,N_2662);
nor U4014 (N_4014,N_2132,N_2664);
nor U4015 (N_4015,N_3346,N_2337);
or U4016 (N_4016,N_3848,N_2590);
xor U4017 (N_4017,N_2273,N_3809);
xor U4018 (N_4018,N_3193,N_3520);
nand U4019 (N_4019,N_3065,N_2767);
and U4020 (N_4020,N_2144,N_3449);
xnor U4021 (N_4021,N_2442,N_2446);
or U4022 (N_4022,N_2581,N_3407);
and U4023 (N_4023,N_2372,N_3188);
or U4024 (N_4024,N_2466,N_3644);
and U4025 (N_4025,N_3004,N_2198);
or U4026 (N_4026,N_3647,N_3811);
xor U4027 (N_4027,N_3655,N_3966);
xor U4028 (N_4028,N_3883,N_2934);
nand U4029 (N_4029,N_2418,N_3884);
and U4030 (N_4030,N_2912,N_3476);
xor U4031 (N_4031,N_2052,N_3175);
xor U4032 (N_4032,N_2184,N_3168);
or U4033 (N_4033,N_3961,N_3492);
xnor U4034 (N_4034,N_3500,N_2569);
nor U4035 (N_4035,N_2048,N_3873);
xor U4036 (N_4036,N_3808,N_2849);
nor U4037 (N_4037,N_3324,N_2051);
and U4038 (N_4038,N_2702,N_3301);
xnor U4039 (N_4039,N_2097,N_2141);
xnor U4040 (N_4040,N_2482,N_2510);
nand U4041 (N_4041,N_3064,N_2787);
nor U4042 (N_4042,N_3041,N_3121);
nand U4043 (N_4043,N_2264,N_3765);
nor U4044 (N_4044,N_3026,N_3745);
nand U4045 (N_4045,N_2576,N_3552);
nor U4046 (N_4046,N_3742,N_3442);
nand U4047 (N_4047,N_3003,N_3758);
and U4048 (N_4048,N_3351,N_2743);
or U4049 (N_4049,N_3378,N_2447);
and U4050 (N_4050,N_3825,N_3399);
or U4051 (N_4051,N_2570,N_2354);
nor U4052 (N_4052,N_2082,N_3381);
or U4053 (N_4053,N_3969,N_3697);
nand U4054 (N_4054,N_3423,N_3143);
nand U4055 (N_4055,N_3137,N_3976);
nor U4056 (N_4056,N_2083,N_3487);
nor U4057 (N_4057,N_2881,N_2479);
and U4058 (N_4058,N_3228,N_3802);
and U4059 (N_4059,N_3155,N_3219);
nor U4060 (N_4060,N_3362,N_3229);
nor U4061 (N_4061,N_3521,N_3959);
or U4062 (N_4062,N_3769,N_2660);
xor U4063 (N_4063,N_3634,N_2328);
nor U4064 (N_4064,N_2394,N_2413);
and U4065 (N_4065,N_2712,N_2452);
or U4066 (N_4066,N_2939,N_3861);
nor U4067 (N_4067,N_3158,N_2682);
xnor U4068 (N_4068,N_2115,N_2758);
xnor U4069 (N_4069,N_2281,N_3119);
and U4070 (N_4070,N_3128,N_3135);
or U4071 (N_4071,N_2403,N_3295);
nor U4072 (N_4072,N_2782,N_3877);
xnor U4073 (N_4073,N_2322,N_2665);
xnor U4074 (N_4074,N_2754,N_2131);
and U4075 (N_4075,N_3293,N_2270);
xnor U4076 (N_4076,N_3240,N_2099);
and U4077 (N_4077,N_2521,N_3865);
or U4078 (N_4078,N_2074,N_3149);
or U4079 (N_4079,N_3899,N_2859);
nor U4080 (N_4080,N_3584,N_3093);
xor U4081 (N_4081,N_3666,N_3816);
nand U4082 (N_4082,N_3331,N_3245);
nor U4083 (N_4083,N_2562,N_3148);
xnor U4084 (N_4084,N_2795,N_2398);
xnor U4085 (N_4085,N_3360,N_3614);
nand U4086 (N_4086,N_3429,N_2799);
nor U4087 (N_4087,N_3267,N_2639);
nand U4088 (N_4088,N_3033,N_3220);
nor U4089 (N_4089,N_2777,N_3886);
nor U4090 (N_4090,N_2142,N_3989);
and U4091 (N_4091,N_2381,N_2701);
xor U4092 (N_4092,N_2683,N_3673);
xor U4093 (N_4093,N_2415,N_2488);
nand U4094 (N_4094,N_3537,N_2265);
or U4095 (N_4095,N_3791,N_2648);
nand U4096 (N_4096,N_2967,N_2651);
and U4097 (N_4097,N_3044,N_3479);
nand U4098 (N_4098,N_2686,N_3856);
xnor U4099 (N_4099,N_2745,N_3024);
and U4100 (N_4100,N_2538,N_2386);
nand U4101 (N_4101,N_2926,N_2755);
xor U4102 (N_4102,N_3624,N_2535);
nand U4103 (N_4103,N_2757,N_2587);
nor U4104 (N_4104,N_2916,N_3935);
xnor U4105 (N_4105,N_2788,N_2460);
xnor U4106 (N_4106,N_2243,N_2716);
xnor U4107 (N_4107,N_3785,N_2455);
or U4108 (N_4108,N_3784,N_3023);
nand U4109 (N_4109,N_2242,N_3287);
xor U4110 (N_4110,N_2780,N_3080);
or U4111 (N_4111,N_3129,N_2943);
nand U4112 (N_4112,N_2953,N_3872);
or U4113 (N_4113,N_3179,N_2719);
nor U4114 (N_4114,N_3425,N_2399);
and U4115 (N_4115,N_2707,N_3600);
or U4116 (N_4116,N_2171,N_2039);
xor U4117 (N_4117,N_2042,N_3377);
or U4118 (N_4118,N_3231,N_2540);
and U4119 (N_4119,N_3262,N_3012);
nand U4120 (N_4120,N_2101,N_2526);
nand U4121 (N_4121,N_2993,N_3938);
or U4122 (N_4122,N_3857,N_3268);
nor U4123 (N_4123,N_3067,N_2670);
nand U4124 (N_4124,N_3868,N_3007);
nor U4125 (N_4125,N_2609,N_3541);
xnor U4126 (N_4126,N_3800,N_3704);
nor U4127 (N_4127,N_3355,N_2313);
or U4128 (N_4128,N_2773,N_2607);
and U4129 (N_4129,N_3009,N_2251);
xor U4130 (N_4130,N_2183,N_3201);
nor U4131 (N_4131,N_3958,N_3528);
and U4132 (N_4132,N_3196,N_3592);
and U4133 (N_4133,N_3933,N_3088);
nor U4134 (N_4134,N_2798,N_2964);
or U4135 (N_4135,N_2721,N_2181);
nor U4136 (N_4136,N_2071,N_2697);
nor U4137 (N_4137,N_2524,N_3798);
xor U4138 (N_4138,N_2143,N_3167);
and U4139 (N_4139,N_2899,N_2734);
xnor U4140 (N_4140,N_2962,N_3912);
xor U4141 (N_4141,N_2661,N_3187);
or U4142 (N_4142,N_3512,N_2935);
nor U4143 (N_4143,N_2778,N_3757);
xnor U4144 (N_4144,N_3733,N_3968);
nor U4145 (N_4145,N_2797,N_2692);
nand U4146 (N_4146,N_3599,N_3172);
and U4147 (N_4147,N_3553,N_2204);
and U4148 (N_4148,N_2362,N_3635);
nand U4149 (N_4149,N_3519,N_2401);
nor U4150 (N_4150,N_3475,N_3412);
xnor U4151 (N_4151,N_2383,N_3709);
nand U4152 (N_4152,N_3146,N_3332);
and U4153 (N_4153,N_3527,N_3543);
nor U4154 (N_4154,N_3402,N_3907);
nor U4155 (N_4155,N_3740,N_2998);
xor U4156 (N_4156,N_2388,N_3236);
or U4157 (N_4157,N_3894,N_3507);
xor U4158 (N_4158,N_3762,N_3028);
xnor U4159 (N_4159,N_3214,N_3781);
nor U4160 (N_4160,N_3680,N_2496);
or U4161 (N_4161,N_2477,N_3169);
nand U4162 (N_4162,N_3040,N_3794);
nand U4163 (N_4163,N_3133,N_3288);
nand U4164 (N_4164,N_3893,N_3754);
xnor U4165 (N_4165,N_3498,N_3109);
xnor U4166 (N_4166,N_3855,N_2594);
or U4167 (N_4167,N_2595,N_3387);
xor U4168 (N_4168,N_3439,N_3300);
xnor U4169 (N_4169,N_2948,N_3692);
nor U4170 (N_4170,N_3385,N_2325);
nor U4171 (N_4171,N_3864,N_2667);
or U4172 (N_4172,N_2634,N_3059);
nor U4173 (N_4173,N_2599,N_2542);
nor U4174 (N_4174,N_3951,N_2913);
or U4175 (N_4175,N_2128,N_3918);
or U4176 (N_4176,N_3678,N_3180);
nand U4177 (N_4177,N_2494,N_2221);
nor U4178 (N_4178,N_2098,N_3780);
nor U4179 (N_4179,N_3750,N_3084);
and U4180 (N_4180,N_3474,N_2009);
and U4181 (N_4181,N_2461,N_2223);
xnor U4182 (N_4182,N_3820,N_3730);
nand U4183 (N_4183,N_2073,N_2266);
and U4184 (N_4184,N_2192,N_2803);
and U4185 (N_4185,N_2200,N_2503);
nor U4186 (N_4186,N_2515,N_2825);
or U4187 (N_4187,N_2019,N_2218);
and U4188 (N_4188,N_3403,N_2980);
nor U4189 (N_4189,N_3650,N_3303);
or U4190 (N_4190,N_3424,N_3141);
xnor U4191 (N_4191,N_3207,N_3013);
nand U4192 (N_4192,N_2997,N_2088);
or U4193 (N_4193,N_3693,N_2714);
xor U4194 (N_4194,N_3726,N_3889);
or U4195 (N_4195,N_3689,N_3944);
nand U4196 (N_4196,N_2196,N_3448);
nor U4197 (N_4197,N_2434,N_3055);
xor U4198 (N_4198,N_3092,N_3652);
nand U4199 (N_4199,N_3834,N_2116);
xnor U4200 (N_4200,N_3459,N_3761);
nor U4201 (N_4201,N_2829,N_3797);
nor U4202 (N_4202,N_3255,N_3379);
nand U4203 (N_4203,N_3111,N_2968);
nand U4204 (N_4204,N_2598,N_3783);
nand U4205 (N_4205,N_2213,N_2404);
nand U4206 (N_4206,N_3192,N_2041);
nor U4207 (N_4207,N_3720,N_3263);
xor U4208 (N_4208,N_3395,N_3558);
and U4209 (N_4209,N_2827,N_2933);
and U4210 (N_4210,N_3994,N_3595);
or U4211 (N_4211,N_3075,N_3435);
nor U4212 (N_4212,N_2150,N_2380);
xor U4213 (N_4213,N_2037,N_2378);
xnor U4214 (N_4214,N_2032,N_2427);
xor U4215 (N_4215,N_2024,N_3194);
and U4216 (N_4216,N_3383,N_3923);
and U4217 (N_4217,N_3839,N_2681);
or U4218 (N_4218,N_2384,N_2812);
nand U4219 (N_4219,N_2571,N_3842);
and U4220 (N_4220,N_2591,N_3322);
xnor U4221 (N_4221,N_2696,N_2880);
xor U4222 (N_4222,N_2317,N_2627);
or U4223 (N_4223,N_2152,N_3586);
nand U4224 (N_4224,N_3656,N_3759);
or U4225 (N_4225,N_2272,N_2285);
nand U4226 (N_4226,N_2638,N_3509);
nor U4227 (N_4227,N_2557,N_2624);
xnor U4228 (N_4228,N_3513,N_3392);
and U4229 (N_4229,N_2275,N_2431);
nand U4230 (N_4230,N_2345,N_2653);
nor U4231 (N_4231,N_2261,N_2654);
or U4232 (N_4232,N_2089,N_2256);
and U4233 (N_4233,N_2885,N_3421);
or U4234 (N_4234,N_3570,N_3357);
xnor U4235 (N_4235,N_2616,N_3675);
and U4236 (N_4236,N_3197,N_2257);
nor U4237 (N_4237,N_2911,N_3506);
nor U4238 (N_4238,N_2886,N_3799);
xor U4239 (N_4239,N_3422,N_3627);
xnor U4240 (N_4240,N_2730,N_3460);
and U4241 (N_4241,N_3753,N_3508);
xnor U4242 (N_4242,N_2561,N_2080);
or U4243 (N_4243,N_3514,N_2874);
nor U4244 (N_4244,N_2269,N_3525);
or U4245 (N_4245,N_2018,N_2956);
or U4246 (N_4246,N_2249,N_3190);
nand U4247 (N_4247,N_2991,N_2338);
nand U4248 (N_4248,N_3140,N_2583);
and U4249 (N_4249,N_3481,N_2230);
nand U4250 (N_4250,N_3056,N_2672);
xor U4251 (N_4251,N_3482,N_3913);
nand U4252 (N_4252,N_3568,N_3131);
or U4253 (N_4253,N_2501,N_2689);
xor U4254 (N_4254,N_3625,N_3364);
xor U4255 (N_4255,N_3696,N_2597);
xor U4256 (N_4256,N_3497,N_2532);
nand U4257 (N_4257,N_3574,N_3036);
xor U4258 (N_4258,N_2924,N_2095);
nand U4259 (N_4259,N_2465,N_3555);
nor U4260 (N_4260,N_2695,N_2070);
and U4261 (N_4261,N_2843,N_2333);
and U4262 (N_4262,N_2642,N_2010);
or U4263 (N_4263,N_3311,N_3037);
xor U4264 (N_4264,N_2279,N_2564);
xor U4265 (N_4265,N_3027,N_2835);
and U4266 (N_4266,N_2981,N_2974);
xnor U4267 (N_4267,N_2472,N_2842);
and U4268 (N_4268,N_2582,N_2193);
xor U4269 (N_4269,N_3151,N_3401);
xor U4270 (N_4270,N_2077,N_2484);
or U4271 (N_4271,N_2170,N_3921);
xor U4272 (N_4272,N_3778,N_2172);
xor U4273 (N_4273,N_2055,N_3916);
or U4274 (N_4274,N_3309,N_2687);
or U4275 (N_4275,N_3587,N_2314);
or U4276 (N_4276,N_3937,N_2989);
nand U4277 (N_4277,N_3076,N_2303);
or U4278 (N_4278,N_2444,N_3828);
xnor U4279 (N_4279,N_2584,N_3598);
nand U4280 (N_4280,N_3536,N_3078);
or U4281 (N_4281,N_2226,N_2965);
and U4282 (N_4282,N_3843,N_3363);
xor U4283 (N_4283,N_2347,N_3165);
nand U4284 (N_4284,N_2632,N_2514);
or U4285 (N_4285,N_2861,N_2485);
nor U4286 (N_4286,N_3618,N_3330);
and U4287 (N_4287,N_2868,N_3159);
xnor U4288 (N_4288,N_3620,N_2613);
or U4289 (N_4289,N_3623,N_2112);
or U4290 (N_4290,N_2884,N_3610);
and U4291 (N_4291,N_3885,N_3838);
or U4292 (N_4292,N_3317,N_3290);
nand U4293 (N_4293,N_3217,N_3896);
nor U4294 (N_4294,N_3538,N_2355);
and U4295 (N_4295,N_3182,N_2065);
or U4296 (N_4296,N_3202,N_3621);
xnor U4297 (N_4297,N_2093,N_2704);
and U4298 (N_4298,N_3826,N_3132);
xor U4299 (N_4299,N_2832,N_2847);
or U4300 (N_4300,N_2853,N_3242);
nand U4301 (N_4301,N_2839,N_2500);
nand U4302 (N_4302,N_3665,N_3427);
nand U4303 (N_4303,N_2016,N_3089);
xnor U4304 (N_4304,N_3639,N_2614);
nor U4305 (N_4305,N_2026,N_3394);
or U4306 (N_4306,N_2910,N_3557);
nand U4307 (N_4307,N_2480,N_2909);
nor U4308 (N_4308,N_3996,N_3882);
and U4309 (N_4309,N_3336,N_2940);
and U4310 (N_4310,N_2674,N_2845);
nor U4311 (N_4311,N_2931,N_2129);
and U4312 (N_4312,N_3420,N_3531);
nand U4313 (N_4313,N_3943,N_3768);
nor U4314 (N_4314,N_2499,N_3849);
xnor U4315 (N_4315,N_2768,N_3561);
and U4316 (N_4316,N_3022,N_2457);
or U4317 (N_4317,N_3273,N_2894);
nand U4318 (N_4318,N_2212,N_2293);
xor U4319 (N_4319,N_2146,N_3211);
nand U4320 (N_4320,N_3939,N_3279);
or U4321 (N_4321,N_2781,N_3567);
nor U4322 (N_4322,N_2250,N_3563);
and U4323 (N_4323,N_3284,N_2330);
nand U4324 (N_4324,N_3812,N_2315);
and U4325 (N_4325,N_3747,N_3393);
and U4326 (N_4326,N_3184,N_3609);
and U4327 (N_4327,N_2545,N_2342);
xnor U4328 (N_4328,N_2211,N_2858);
or U4329 (N_4329,N_2100,N_3386);
or U4330 (N_4330,N_2530,N_3619);
nor U4331 (N_4331,N_3501,N_3703);
or U4332 (N_4332,N_3682,N_2182);
nand U4333 (N_4333,N_3806,N_2879);
or U4334 (N_4334,N_3473,N_2700);
and U4335 (N_4335,N_3348,N_3252);
or U4336 (N_4336,N_2691,N_3087);
nor U4337 (N_4337,N_3134,N_2332);
nand U4338 (N_4338,N_3410,N_3283);
and U4339 (N_4339,N_3947,N_3281);
or U4340 (N_4340,N_3455,N_2722);
xor U4341 (N_4341,N_2202,N_2469);
and U4342 (N_4342,N_2240,N_2505);
and U4343 (N_4343,N_2114,N_3591);
nand U4344 (N_4344,N_2895,N_3156);
or U4345 (N_4345,N_3977,N_2451);
nand U4346 (N_4346,N_3396,N_3350);
nor U4347 (N_4347,N_3888,N_2887);
xor U4348 (N_4348,N_2647,N_3462);
nor U4349 (N_4349,N_3851,N_2331);
nand U4350 (N_4350,N_3315,N_3047);
xnor U4351 (N_4351,N_2625,N_2905);
or U4352 (N_4352,N_3206,N_3174);
or U4353 (N_4353,N_3480,N_3391);
xor U4354 (N_4354,N_3814,N_3787);
nand U4355 (N_4355,N_3897,N_3850);
or U4356 (N_4356,N_2102,N_2785);
nor U4357 (N_4357,N_2851,N_3737);
nor U4358 (N_4358,N_3551,N_3296);
or U4359 (N_4359,N_2476,N_3082);
nand U4360 (N_4360,N_2475,N_3565);
and U4361 (N_4361,N_2007,N_2929);
and U4362 (N_4362,N_3967,N_3000);
xor U4363 (N_4363,N_2405,N_2808);
nand U4364 (N_4364,N_3819,N_3370);
or U4365 (N_4365,N_3562,N_2208);
and U4366 (N_4366,N_2326,N_3719);
and U4367 (N_4367,N_2786,N_2869);
nor U4368 (N_4368,N_2214,N_3323);
nor U4369 (N_4369,N_2263,N_2891);
and U4370 (N_4370,N_3583,N_2814);
nand U4371 (N_4371,N_3622,N_3212);
xnor U4372 (N_4372,N_2489,N_2134);
or U4373 (N_4373,N_3588,N_2274);
or U4374 (N_4374,N_2365,N_3199);
nor U4375 (N_4375,N_2680,N_2040);
nand U4376 (N_4376,N_2155,N_2126);
and U4377 (N_4377,N_3216,N_3428);
and U4378 (N_4378,N_3289,N_3575);
and U4379 (N_4379,N_3903,N_3260);
and U4380 (N_4380,N_3988,N_2137);
or U4381 (N_4381,N_3071,N_2066);
or U4382 (N_4382,N_2602,N_3018);
and U4383 (N_4383,N_3698,N_2944);
xnor U4384 (N_4384,N_2603,N_2729);
xnor U4385 (N_4385,N_2081,N_3775);
and U4386 (N_4386,N_2920,N_2059);
xnor U4387 (N_4387,N_2988,N_3069);
or U4388 (N_4388,N_3265,N_3549);
nand U4389 (N_4389,N_3472,N_2844);
or U4390 (N_4390,N_3359,N_2575);
or U4391 (N_4391,N_2927,N_3342);
or U4392 (N_4392,N_2278,N_2225);
nor U4393 (N_4393,N_2950,N_2207);
and U4394 (N_4394,N_2229,N_3942);
xnor U4395 (N_4395,N_2541,N_2973);
nand U4396 (N_4396,N_2318,N_3251);
and U4397 (N_4397,N_3468,N_3915);
nor U4398 (N_4398,N_3960,N_2543);
nand U4399 (N_4399,N_2292,N_2657);
and U4400 (N_4400,N_2731,N_2283);
and U4401 (N_4401,N_3679,N_2246);
or U4402 (N_4402,N_2034,N_2820);
or U4403 (N_4403,N_3408,N_3605);
or U4404 (N_4404,N_3734,N_2806);
nor U4405 (N_4405,N_2149,N_2079);
nor U4406 (N_4406,N_2772,N_2057);
and U4407 (N_4407,N_2685,N_3239);
nor U4408 (N_4408,N_2908,N_2177);
nand U4409 (N_4409,N_3491,N_2320);
nor U4410 (N_4410,N_3971,N_3774);
and U4411 (N_4411,N_2675,N_3547);
xor U4412 (N_4412,N_3796,N_3936);
nand U4413 (N_4413,N_2348,N_2506);
nor U4414 (N_4414,N_3486,N_3478);
nand U4415 (N_4415,N_3743,N_3608);
nor U4416 (N_4416,N_2357,N_3454);
and U4417 (N_4417,N_2713,N_2669);
xor U4418 (N_4418,N_3900,N_3540);
nand U4419 (N_4419,N_2118,N_3259);
xor U4420 (N_4420,N_3560,N_3653);
or U4421 (N_4421,N_2531,N_3006);
or U4422 (N_4422,N_3496,N_3891);
xor U4423 (N_4423,N_3788,N_3594);
or U4424 (N_4424,N_2021,N_2368);
or U4425 (N_4425,N_3702,N_3505);
and U4426 (N_4426,N_2507,N_2893);
nand U4427 (N_4427,N_2421,N_3249);
or U4428 (N_4428,N_2299,N_2197);
nor U4429 (N_4429,N_3795,N_2110);
or U4430 (N_4430,N_2433,N_3672);
nand U4431 (N_4431,N_3782,N_3285);
nand U4432 (N_4432,N_2677,N_2508);
xnor U4433 (N_4433,N_3739,N_2739);
nor U4434 (N_4434,N_3997,N_3941);
or U4435 (N_4435,N_2828,N_3038);
or U4436 (N_4436,N_3398,N_2736);
nand U4437 (N_4437,N_3919,N_3706);
nor U4438 (N_4438,N_2996,N_3548);
xnor U4439 (N_4439,N_3215,N_2986);
nand U4440 (N_4440,N_2572,N_3057);
nor U4441 (N_4441,N_3645,N_3438);
xor U4442 (N_4442,N_3426,N_3471);
or U4443 (N_4443,N_3646,N_3337);
nand U4444 (N_4444,N_3773,N_2219);
and U4445 (N_4445,N_3443,N_2222);
nor U4446 (N_4446,N_3264,N_2140);
or U4447 (N_4447,N_2834,N_3335);
xor U4448 (N_4448,N_3477,N_3320);
xor U4449 (N_4449,N_3107,N_2619);
nor U4450 (N_4450,N_2244,N_3312);
or U4451 (N_4451,N_3444,N_3927);
or U4452 (N_4452,N_3684,N_2179);
nand U4453 (N_4453,N_2726,N_2280);
or U4454 (N_4454,N_3982,N_3792);
nor U4455 (N_4455,N_2789,N_2186);
or U4456 (N_4456,N_3400,N_2429);
or U4457 (N_4457,N_2589,N_3566);
xor U4458 (N_4458,N_3327,N_2113);
and U4459 (N_4459,N_3366,N_2316);
and U4460 (N_4460,N_3887,N_2992);
nand U4461 (N_4461,N_2862,N_3451);
or U4462 (N_4462,N_2025,N_2703);
nor U4463 (N_4463,N_3981,N_2258);
and U4464 (N_4464,N_3998,N_3361);
and U4465 (N_4465,N_3829,N_3338);
xor U4466 (N_4466,N_3494,N_2124);
and U4467 (N_4467,N_3905,N_3633);
nand U4468 (N_4468,N_2206,N_3596);
nor U4469 (N_4469,N_3928,N_3375);
and U4470 (N_4470,N_2872,N_3611);
nand U4471 (N_4471,N_2076,N_2856);
and U4472 (N_4472,N_2706,N_3637);
and U4473 (N_4473,N_2054,N_3083);
or U4474 (N_4474,N_3081,N_2023);
xor U4475 (N_4475,N_3949,N_3911);
nand U4476 (N_4476,N_3685,N_3470);
xor U4477 (N_4477,N_3417,N_2649);
xor U4478 (N_4478,N_2883,N_2063);
or U4479 (N_4479,N_2817,N_3844);
nor U4480 (N_4480,N_2605,N_2645);
nand U4481 (N_4481,N_3751,N_3329);
nand U4482 (N_4482,N_3298,N_3050);
nand U4483 (N_4483,N_3397,N_3931);
and U4484 (N_4484,N_3147,N_2783);
nor U4485 (N_4485,N_3721,N_2617);
or U4486 (N_4486,N_3840,N_2904);
and U4487 (N_4487,N_2031,N_3578);
or U4488 (N_4488,N_3445,N_3741);
xnor U4489 (N_4489,N_3127,N_3356);
or U4490 (N_4490,N_3409,N_3823);
and U4491 (N_4491,N_2903,N_2166);
or U4492 (N_4492,N_3237,N_3643);
xnor U4493 (N_4493,N_2554,N_2191);
nor U4494 (N_4494,N_3021,N_2033);
xor U4495 (N_4495,N_3875,N_3272);
xnor U4496 (N_4496,N_2363,N_3573);
nand U4497 (N_4497,N_2690,N_3863);
and U4498 (N_4498,N_2459,N_3384);
nand U4499 (N_4499,N_2533,N_3546);
nor U4500 (N_4500,N_3554,N_2287);
or U4501 (N_4501,N_3029,N_3510);
or U4502 (N_4502,N_3995,N_3371);
and U4503 (N_4503,N_2498,N_3970);
or U4504 (N_4504,N_2245,N_3764);
nand U4505 (N_4505,N_2741,N_2189);
xnor U4506 (N_4506,N_3483,N_2323);
and U4507 (N_4507,N_2906,N_2568);
nor U4508 (N_4508,N_3198,N_3490);
xor U4509 (N_4509,N_3015,N_3670);
nand U4510 (N_4510,N_2437,N_2050);
nand U4511 (N_4511,N_3962,N_3690);
nor U4512 (N_4512,N_2776,N_2840);
and U4513 (N_4513,N_3660,N_2120);
or U4514 (N_4514,N_3576,N_2865);
and U4515 (N_4515,N_2923,N_3223);
nand U4516 (N_4516,N_2710,N_3389);
or U4517 (N_4517,N_3171,N_3854);
or U4518 (N_4518,N_3051,N_3440);
or U4519 (N_4519,N_3125,N_2976);
nor U4520 (N_4520,N_2864,N_3511);
nand U4521 (N_4521,N_2813,N_2454);
or U4522 (N_4522,N_3178,N_3984);
or U4523 (N_4523,N_2043,N_2949);
xnor U4524 (N_4524,N_3489,N_2738);
nor U4525 (N_4525,N_3777,N_2056);
xnor U4526 (N_4526,N_2014,N_3590);
nand U4527 (N_4527,N_2938,N_2523);
and U4528 (N_4528,N_2321,N_2511);
and U4529 (N_4529,N_3045,N_2830);
or U4530 (N_4530,N_3458,N_2746);
or U4531 (N_4531,N_2492,N_2958);
nand U4532 (N_4532,N_3822,N_3048);
nand U4533 (N_4533,N_3728,N_2539);
and U4534 (N_4534,N_2668,N_3805);
nand U4535 (N_4535,N_2400,N_3948);
xor U4536 (N_4536,N_3085,N_3755);
nand U4537 (N_4537,N_3054,N_3271);
or U4538 (N_4538,N_2195,N_3658);
and U4539 (N_4539,N_2068,N_3817);
nor U4540 (N_4540,N_3581,N_2307);
nand U4541 (N_4541,N_2169,N_3999);
nor U4542 (N_4542,N_2168,N_2260);
or U4543 (N_4543,N_2424,N_2982);
nor U4544 (N_4544,N_2705,N_2450);
nand U4545 (N_4545,N_2860,N_3108);
nand U4546 (N_4546,N_2644,N_2364);
nor U4547 (N_4547,N_3310,N_3373);
nor U4548 (N_4548,N_2611,N_2020);
and U4549 (N_4549,N_2406,N_3105);
xor U4550 (N_4550,N_2359,N_3368);
or U4551 (N_4551,N_3382,N_3908);
or U4552 (N_4552,N_2676,N_2423);
nor U4553 (N_4553,N_3657,N_2493);
xor U4554 (N_4554,N_2267,N_2504);
and U4555 (N_4555,N_3274,N_3859);
nand U4556 (N_4556,N_3688,N_3807);
nor U4557 (N_4557,N_3299,N_2119);
and U4558 (N_4558,N_2977,N_2090);
nand U4559 (N_4559,N_3163,N_2804);
nand U4560 (N_4560,N_2271,N_2029);
nand U4561 (N_4561,N_2392,N_3469);
xnor U4562 (N_4562,N_2878,N_2936);
xnor U4563 (N_4563,N_3112,N_2922);
or U4564 (N_4564,N_3845,N_3020);
or U4565 (N_4565,N_2176,N_2567);
nor U4566 (N_4566,N_2838,N_2495);
nand U4567 (N_4567,N_3965,N_2094);
xor U4568 (N_4568,N_2103,N_2304);
nand U4569 (N_4569,N_2520,N_3801);
nand U4570 (N_4570,N_3846,N_3177);
or U4571 (N_4571,N_2527,N_3333);
nand U4572 (N_4572,N_2154,N_2740);
nand U4573 (N_4573,N_3414,N_3835);
or U4574 (N_4574,N_2136,N_3975);
and U4575 (N_4575,N_2544,N_3302);
nand U4576 (N_4576,N_3963,N_3779);
nor U4577 (N_4577,N_3031,N_2159);
or U4578 (N_4578,N_2153,N_3304);
xor U4579 (N_4579,N_2422,N_2462);
and U4580 (N_4580,N_2216,N_3654);
or U4581 (N_4581,N_2268,N_3195);
or U4582 (N_4582,N_2556,N_3254);
nand U4583 (N_4583,N_3874,N_2174);
nor U4584 (N_4584,N_2559,N_3722);
nor U4585 (N_4585,N_2443,N_3542);
or U4586 (N_4586,N_2369,N_3749);
nand U4587 (N_4587,N_2294,N_2688);
xor U4588 (N_4588,N_2629,N_3871);
and U4589 (N_4589,N_2000,N_2833);
and U4590 (N_4590,N_3222,N_2420);
xor U4591 (N_4591,N_2105,N_2435);
xnor U4592 (N_4592,N_2069,N_2382);
nor U4593 (N_4593,N_2379,N_3956);
nor U4594 (N_4594,N_2866,N_2735);
xor U4595 (N_4595,N_3014,N_2402);
nand U4596 (N_4596,N_2407,N_3433);
and U4597 (N_4597,N_2376,N_3106);
or U4598 (N_4598,N_3736,N_3241);
xor U4599 (N_4599,N_2127,N_2588);
and U4600 (N_4600,N_3144,N_2252);
xnor U4601 (N_4601,N_2167,N_2578);
nor U4602 (N_4602,N_2324,N_3316);
or U4603 (N_4603,N_2774,N_2942);
and U4604 (N_4604,N_3437,N_3945);
nor U4605 (N_4605,N_2641,N_2291);
nand U4606 (N_4606,N_3499,N_2419);
or U4607 (N_4607,N_3522,N_3668);
or U4608 (N_4608,N_2044,N_3793);
nand U4609 (N_4609,N_3307,N_2237);
and U4610 (N_4610,N_3235,N_2478);
or U4611 (N_4611,N_2826,N_2646);
nand U4612 (N_4612,N_3524,N_2658);
xor U4613 (N_4613,N_3636,N_2753);
nand U4614 (N_4614,N_2277,N_3091);
and U4615 (N_4615,N_2852,N_3987);
nor U4616 (N_4616,N_2282,N_3671);
xor U4617 (N_4617,N_3833,N_3390);
or U4618 (N_4618,N_3166,N_3354);
nor U4619 (N_4619,N_3616,N_2724);
nand U4620 (N_4620,N_3374,N_2412);
nand U4621 (N_4621,N_2941,N_3042);
nand U4622 (N_4622,N_2109,N_2305);
or U4623 (N_4623,N_2284,N_2121);
nor U4624 (N_4624,N_2106,N_3341);
nor U4625 (N_4625,N_3752,N_2678);
nand U4626 (N_4626,N_3325,N_2635);
nor U4627 (N_4627,N_2162,N_3597);
nor U4628 (N_4628,N_3488,N_2809);
xor U4629 (N_4629,N_2633,N_2491);
nand U4630 (N_4630,N_3154,N_3104);
xnor U4631 (N_4631,N_2536,N_3365);
and U4632 (N_4632,N_2125,N_2486);
and U4633 (N_4633,N_2464,N_3095);
nor U4634 (N_4634,N_2566,N_2512);
nor U4635 (N_4635,N_2002,N_3858);
nor U4636 (N_4636,N_2350,N_2604);
and U4637 (N_4637,N_2979,N_2053);
nand U4638 (N_4638,N_2550,N_2652);
and U4639 (N_4639,N_3532,N_3130);
or U4640 (N_4640,N_3418,N_3097);
or U4641 (N_4641,N_3946,N_2210);
xor U4642 (N_4642,N_3415,N_3319);
nor U4643 (N_4643,N_2439,N_3630);
or U4644 (N_4644,N_3464,N_2796);
xnor U4645 (N_4645,N_2694,N_2837);
xor U4646 (N_4646,N_2175,N_2917);
nor U4647 (N_4647,N_2580,N_3205);
nor U4648 (N_4648,N_3258,N_2302);
or U4649 (N_4649,N_3818,N_2436);
or U4650 (N_4650,N_3210,N_2311);
or U4651 (N_4651,N_2474,N_2513);
or U4652 (N_4652,N_3550,N_2139);
or U4653 (N_4653,N_2620,N_3725);
nand U4654 (N_4654,N_3631,N_2519);
nor U4655 (N_4655,N_3602,N_3306);
nor U4656 (N_4656,N_2563,N_2855);
or U4657 (N_4657,N_3136,N_2091);
and U4658 (N_4658,N_2387,N_2471);
and U4659 (N_4659,N_3016,N_2698);
nand U4660 (N_4660,N_2699,N_3345);
and U4661 (N_4661,N_3232,N_3227);
xnor U4662 (N_4662,N_2742,N_2728);
nor U4663 (N_4663,N_2289,N_2548);
nand U4664 (N_4664,N_2610,N_2343);
or U4665 (N_4665,N_2078,N_2393);
xor U4666 (N_4666,N_2440,N_3953);
nand U4667 (N_4667,N_2650,N_2356);
xor U4668 (N_4668,N_3841,N_2666);
nor U4669 (N_4669,N_3053,N_3213);
and U4670 (N_4670,N_3649,N_3717);
and U4671 (N_4671,N_3723,N_2715);
nor U4672 (N_4672,N_2373,N_3124);
and U4673 (N_4673,N_2161,N_2027);
and U4674 (N_4674,N_2072,N_3034);
and U4675 (N_4675,N_2453,N_2396);
nand U4676 (N_4676,N_2445,N_2896);
nor U4677 (N_4677,N_3367,N_3406);
or U4678 (N_4678,N_2807,N_2165);
and U4679 (N_4679,N_2971,N_3277);
nor U4680 (N_4680,N_3746,N_3504);
nand U4681 (N_4681,N_3257,N_2483);
xor U4682 (N_4682,N_2235,N_3866);
or U4683 (N_4683,N_2857,N_3162);
nor U4684 (N_4684,N_3909,N_2630);
nand U4685 (N_4685,N_2717,N_3867);
or U4686 (N_4686,N_2295,N_2552);
xor U4687 (N_4687,N_2727,N_2107);
and U4688 (N_4688,N_3786,N_3173);
or U4689 (N_4689,N_3530,N_2353);
nor U4690 (N_4690,N_2038,N_3694);
and U4691 (N_4691,N_3691,N_2408);
and U4692 (N_4692,N_3579,N_2417);
nand U4693 (N_4693,N_3072,N_3572);
nand U4694 (N_4694,N_2209,N_2873);
nor U4695 (N_4695,N_2636,N_3986);
nand U4696 (N_4696,N_3606,N_2233);
or U4697 (N_4697,N_2747,N_2737);
nand U4698 (N_4698,N_3314,N_2117);
or U4699 (N_4699,N_2761,N_3079);
xnor U4700 (N_4700,N_2987,N_2203);
or U4701 (N_4701,N_3804,N_2430);
nand U4702 (N_4702,N_3294,N_3280);
and U4703 (N_4703,N_3208,N_2004);
nor U4704 (N_4704,N_2579,N_2049);
xnor U4705 (N_4705,N_2188,N_2130);
xor U4706 (N_4706,N_2537,N_2810);
nor U4707 (N_4707,N_3744,N_2766);
nor U4708 (N_4708,N_3347,N_3544);
and U4709 (N_4709,N_3074,N_3446);
nor U4710 (N_4710,N_2232,N_2889);
nor U4711 (N_4711,N_2199,N_2087);
nor U4712 (N_4712,N_2955,N_2067);
nand U4713 (N_4713,N_3145,N_3604);
or U4714 (N_4714,N_2205,N_3077);
nand U4715 (N_4715,N_2606,N_3209);
and U4716 (N_4716,N_3275,N_3529);
xor U4717 (N_4717,N_3101,N_3878);
and U4718 (N_4718,N_2148,N_2111);
xor U4719 (N_4719,N_3138,N_2901);
nor U4720 (N_4720,N_3117,N_3710);
xor U4721 (N_4721,N_2358,N_3523);
or U4722 (N_4722,N_3419,N_2631);
xor U4723 (N_4723,N_3950,N_3261);
nand U4724 (N_4724,N_2086,N_3122);
or U4725 (N_4725,N_3589,N_3224);
or U4726 (N_4726,N_2036,N_3929);
and U4727 (N_4727,N_2395,N_3432);
and U4728 (N_4728,N_3465,N_3266);
nor U4729 (N_4729,N_2928,N_3305);
and U4730 (N_4730,N_2301,N_3651);
or U4731 (N_4731,N_2622,N_2925);
xnor U4732 (N_4732,N_3830,N_3103);
nand U4733 (N_4733,N_3043,N_3060);
nor U4734 (N_4734,N_3226,N_2972);
nor U4735 (N_4735,N_2823,N_2995);
xor U4736 (N_4736,N_3230,N_2351);
nor U4737 (N_4737,N_2999,N_2871);
nor U4738 (N_4738,N_3890,N_3910);
nor U4739 (N_4739,N_2349,N_2970);
nand U4740 (N_4740,N_3534,N_3436);
xor U4741 (N_4741,N_2975,N_2771);
and U4742 (N_4742,N_3142,N_2551);
or U4743 (N_4743,N_3629,N_2930);
or U4744 (N_4744,N_2060,N_2882);
nand U4745 (N_4745,N_2663,N_2907);
or U4746 (N_4746,N_3836,N_2762);
and U4747 (N_4747,N_3827,N_2259);
nand U4748 (N_4748,N_3932,N_2811);
xnor U4749 (N_4749,N_3358,N_3687);
and U4750 (N_4750,N_2846,N_2800);
and U4751 (N_4751,N_3126,N_2518);
nand U4752 (N_4752,N_3990,N_3434);
xor U4753 (N_4753,N_3766,N_2978);
or U4754 (N_4754,N_2558,N_3025);
or U4755 (N_4755,N_3526,N_3113);
or U4756 (N_4756,N_3659,N_2824);
or U4757 (N_4757,N_3954,N_3924);
or U4758 (N_4758,N_2375,N_2084);
and U4759 (N_4759,N_3535,N_3847);
or U4760 (N_4760,N_2185,N_2888);
or U4761 (N_4761,N_2104,N_3297);
and U4762 (N_4762,N_2708,N_3161);
xnor U4763 (N_4763,N_3411,N_2759);
and U4764 (N_4764,N_3005,N_3369);
and U4765 (N_4765,N_2410,N_2487);
nor U4766 (N_4766,N_3221,N_2615);
nand U4767 (N_4767,N_3983,N_3447);
or U4768 (N_4768,N_3070,N_2534);
xnor U4769 (N_4769,N_2659,N_3638);
nand U4770 (N_4770,N_3763,N_2802);
and U4771 (N_4771,N_2190,N_2329);
xor U4772 (N_4772,N_3467,N_3934);
nor U4773 (N_4773,N_2985,N_3860);
and U4774 (N_4774,N_2096,N_3789);
and U4775 (N_4775,N_2769,N_3253);
and U4776 (N_4776,N_3869,N_3503);
xnor U4777 (N_4777,N_3270,N_2947);
and U4778 (N_4778,N_2217,N_2612);
xnor U4779 (N_4779,N_3593,N_2957);
nand U4780 (N_4780,N_2238,N_3700);
nor U4781 (N_4781,N_2775,N_2448);
nand U4782 (N_4782,N_3898,N_3516);
xor U4783 (N_4783,N_2565,N_3291);
nand U4784 (N_4784,N_3098,N_3904);
or U4785 (N_4785,N_2028,N_3405);
nand U4786 (N_4786,N_3416,N_2784);
and U4787 (N_4787,N_2585,N_3189);
and U4788 (N_4788,N_2201,N_3248);
or U4789 (N_4789,N_2414,N_2490);
xnor U4790 (N_4790,N_2764,N_3972);
xnor U4791 (N_4791,N_2003,N_3862);
and U4792 (N_4792,N_3515,N_2850);
xnor U4793 (N_4793,N_2628,N_3120);
xnor U4794 (N_4794,N_2236,N_2470);
and U4795 (N_4795,N_2135,N_3181);
xor U4796 (N_4796,N_2180,N_3686);
or U4797 (N_4797,N_3642,N_2733);
nand U4798 (N_4798,N_2310,N_2637);
nand U4799 (N_4799,N_3813,N_3321);
and U4800 (N_4800,N_2456,N_3914);
nand U4801 (N_4801,N_2046,N_3556);
or U4802 (N_4802,N_2234,N_3090);
xnor U4803 (N_4803,N_2085,N_3063);
nor U4804 (N_4804,N_2608,N_2145);
nor U4805 (N_4805,N_2960,N_2801);
and U4806 (N_4806,N_2779,N_2959);
or U4807 (N_4807,N_2819,N_2763);
nand U4808 (N_4808,N_3061,N_3585);
and U4809 (N_4809,N_3282,N_2752);
or U4810 (N_4810,N_3920,N_3339);
nor U4811 (N_4811,N_3735,N_3917);
nand U4812 (N_4812,N_2300,N_3881);
xnor U4813 (N_4813,N_3940,N_2336);
or U4814 (N_4814,N_2528,N_2377);
and U4815 (N_4815,N_2673,N_3344);
or U4816 (N_4816,N_2308,N_3456);
and U4817 (N_4817,N_3170,N_3738);
nor U4818 (N_4818,N_3662,N_2215);
nor U4819 (N_4819,N_3803,N_3313);
and U4820 (N_4820,N_3748,N_2848);
nor U4821 (N_4821,N_3648,N_3716);
nor U4822 (N_4822,N_3466,N_2516);
nand U4823 (N_4823,N_2618,N_2151);
and U4824 (N_4824,N_2952,N_3677);
nand U4825 (N_4825,N_3895,N_3973);
nor U4826 (N_4826,N_2863,N_3925);
xor U4827 (N_4827,N_2312,N_2370);
or U4828 (N_4828,N_3086,N_2164);
and U4829 (N_4829,N_3695,N_3334);
or U4830 (N_4830,N_3278,N_3349);
xor U4831 (N_4831,N_2600,N_2123);
nor U4832 (N_4832,N_3980,N_3626);
and U4833 (N_4833,N_2560,N_2725);
xnor U4834 (N_4834,N_3353,N_3244);
xnor U4835 (N_4835,N_2816,N_2792);
and U4836 (N_4836,N_2138,N_3545);
xnor U4837 (N_4837,N_3729,N_2290);
xor U4838 (N_4838,N_3760,N_2008);
nor U4839 (N_4839,N_3233,N_2821);
nor U4840 (N_4840,N_3617,N_2918);
and U4841 (N_4841,N_2319,N_2723);
and U4842 (N_4842,N_2643,N_2409);
xnor U4843 (N_4843,N_2158,N_2255);
nor U4844 (N_4844,N_2227,N_3430);
nor U4845 (N_4845,N_3978,N_3001);
nor U4846 (N_4846,N_2108,N_2449);
nor U4847 (N_4847,N_3096,N_3225);
and U4848 (N_4848,N_3640,N_3058);
or U4849 (N_4849,N_2467,N_3152);
or U4850 (N_4850,N_3380,N_2744);
nor U4851 (N_4851,N_3580,N_2684);
and U4852 (N_4852,N_3256,N_2990);
nor U4853 (N_4853,N_2553,N_2867);
xnor U4854 (N_4854,N_3853,N_2822);
or U4855 (N_4855,N_3286,N_3441);
and U4856 (N_4856,N_2309,N_3246);
and U4857 (N_4857,N_3669,N_3732);
nand U4858 (N_4858,N_2239,N_2438);
nand U4859 (N_4859,N_2062,N_3957);
nand U4860 (N_4860,N_2914,N_3066);
xor U4861 (N_4861,N_2760,N_3569);
or U4862 (N_4862,N_2693,N_2224);
nand U4863 (N_4863,N_3701,N_2656);
xnor U4864 (N_4864,N_3518,N_3191);
and U4865 (N_4865,N_2709,N_2075);
and U4866 (N_4866,N_2122,N_2231);
xor U4867 (N_4867,N_3008,N_3186);
or U4868 (N_4868,N_2297,N_3340);
and U4869 (N_4869,N_2306,N_3035);
nand U4870 (N_4870,N_3017,N_3837);
or U4871 (N_4871,N_3413,N_2748);
or U4872 (N_4872,N_2932,N_2791);
and U4873 (N_4873,N_3115,N_3238);
nor U4874 (N_4874,N_2951,N_2425);
nor U4875 (N_4875,N_3376,N_2163);
or U4876 (N_4876,N_2984,N_3674);
xor U4877 (N_4877,N_2220,N_3641);
nand U4878 (N_4878,N_2711,N_3308);
xnor U4879 (N_4879,N_3715,N_2341);
or U4880 (N_4880,N_2366,N_3613);
or U4881 (N_4881,N_3118,N_2389);
xor U4882 (N_4882,N_3832,N_3906);
nor U4883 (N_4883,N_3699,N_3533);
and U4884 (N_4884,N_3463,N_3183);
xor U4885 (N_4885,N_2011,N_2679);
xor U4886 (N_4886,N_2574,N_3711);
or U4887 (N_4887,N_3901,N_2432);
or U4888 (N_4888,N_2655,N_2340);
xnor U4889 (N_4889,N_2374,N_3852);
or U4890 (N_4890,N_3068,N_2035);
nand U4891 (N_4891,N_3404,N_2463);
or U4892 (N_4892,N_2870,N_2790);
xor U4893 (N_4893,N_2481,N_3153);
nand U4894 (N_4894,N_3292,N_2509);
and U4895 (N_4895,N_2173,N_2006);
xnor U4896 (N_4896,N_2473,N_2966);
nand U4897 (N_4897,N_2522,N_2921);
or U4898 (N_4898,N_3876,N_2047);
xor U4899 (N_4899,N_2416,N_3539);
and U4900 (N_4900,N_3930,N_2751);
and U4901 (N_4901,N_2497,N_2749);
or U4902 (N_4902,N_2793,N_2854);
and U4903 (N_4903,N_3831,N_3352);
nand U4904 (N_4904,N_2058,N_2937);
or U4905 (N_4905,N_2969,N_2983);
nand U4906 (N_4906,N_3964,N_3603);
and U4907 (N_4907,N_2228,N_2897);
or U4908 (N_4908,N_3157,N_2344);
nand U4909 (N_4909,N_2367,N_2626);
xnor U4910 (N_4910,N_3993,N_2335);
and U4911 (N_4911,N_3724,N_3204);
nor U4912 (N_4912,N_2017,N_3493);
and U4913 (N_4913,N_3049,N_2623);
and U4914 (N_4914,N_2898,N_2092);
and U4915 (N_4915,N_2876,N_2875);
and U4916 (N_4916,N_2327,N_3824);
nand U4917 (N_4917,N_3714,N_3032);
nand U4918 (N_4918,N_2288,N_2818);
xnor U4919 (N_4919,N_3062,N_2468);
and U4920 (N_4920,N_2890,N_3756);
or U4921 (N_4921,N_3564,N_2900);
nand U4922 (N_4922,N_2836,N_3431);
or U4923 (N_4923,N_2549,N_2756);
nor U4924 (N_4924,N_3010,N_2022);
or U4925 (N_4925,N_2298,N_3705);
nor U4926 (N_4926,N_3247,N_2276);
xor U4927 (N_4927,N_2012,N_3116);
xor U4928 (N_4928,N_2015,N_2831);
nand U4929 (N_4929,N_2892,N_3502);
nor U4930 (N_4930,N_2586,N_3243);
xnor U4931 (N_4931,N_2254,N_3707);
nand U4932 (N_4932,N_3559,N_2946);
nand U4933 (N_4933,N_2794,N_3902);
xnor U4934 (N_4934,N_2194,N_2001);
and U4935 (N_4935,N_3718,N_2133);
or U4936 (N_4936,N_2841,N_3484);
xor U4937 (N_4937,N_3582,N_3176);
xnor U4938 (N_4938,N_3776,N_2601);
nor U4939 (N_4939,N_3326,N_3770);
nor U4940 (N_4940,N_3955,N_2390);
and U4941 (N_4941,N_2945,N_2147);
nor U4942 (N_4942,N_2178,N_2253);
nand U4943 (N_4943,N_3667,N_2241);
and U4944 (N_4944,N_3453,N_3234);
and U4945 (N_4945,N_2061,N_3731);
nor U4946 (N_4946,N_3810,N_3985);
nor U4947 (N_4947,N_3892,N_3318);
nand U4948 (N_4948,N_2248,N_2805);
and U4949 (N_4949,N_3664,N_2502);
nand U4950 (N_4950,N_3979,N_3328);
nor U4951 (N_4951,N_3019,N_2157);
nand U4952 (N_4952,N_3815,N_2352);
or U4953 (N_4953,N_2334,N_3601);
or U4954 (N_4954,N_3388,N_2013);
or U4955 (N_4955,N_2877,N_3099);
or U4956 (N_4956,N_2770,N_2815);
or U4957 (N_4957,N_3628,N_3992);
and U4958 (N_4958,N_2385,N_3615);
and U4959 (N_4959,N_3110,N_3461);
or U4960 (N_4960,N_3094,N_3661);
xnor U4961 (N_4961,N_2361,N_2346);
xor U4962 (N_4962,N_3571,N_3164);
nor U4963 (N_4963,N_3200,N_3452);
nor U4964 (N_4964,N_2525,N_2546);
or U4965 (N_4965,N_2961,N_3002);
and U4966 (N_4966,N_2963,N_3046);
or U4967 (N_4967,N_3790,N_2005);
nor U4968 (N_4968,N_2411,N_3612);
and U4969 (N_4969,N_3485,N_3771);
and U4970 (N_4970,N_3991,N_2296);
or U4971 (N_4971,N_3772,N_2593);
nand U4972 (N_4972,N_3139,N_3727);
and U4973 (N_4973,N_3879,N_2915);
and U4974 (N_4974,N_3495,N_3632);
and U4975 (N_4975,N_2517,N_2045);
and U4976 (N_4976,N_2397,N_3821);
xor U4977 (N_4977,N_3102,N_2160);
xor U4978 (N_4978,N_2030,N_2994);
and U4979 (N_4979,N_2555,N_3457);
and U4980 (N_4980,N_2765,N_3114);
or U4981 (N_4981,N_3123,N_2262);
and U4982 (N_4982,N_3150,N_3880);
and U4983 (N_4983,N_3870,N_2286);
xnor U4984 (N_4984,N_3974,N_3922);
and U4985 (N_4985,N_3160,N_3185);
or U4986 (N_4986,N_2187,N_3372);
xor U4987 (N_4987,N_2954,N_2732);
and U4988 (N_4988,N_3708,N_3450);
or U4989 (N_4989,N_2596,N_3052);
xnor U4990 (N_4990,N_3577,N_3926);
nor U4991 (N_4991,N_3100,N_3030);
nor U4992 (N_4992,N_2247,N_2592);
nand U4993 (N_4993,N_3607,N_2573);
or U4994 (N_4994,N_2671,N_2371);
xnor U4995 (N_4995,N_2156,N_3517);
xnor U4996 (N_4996,N_3073,N_3011);
nor U4997 (N_4997,N_3952,N_2529);
xnor U4998 (N_4998,N_2902,N_2360);
nand U4999 (N_4999,N_2577,N_2064);
xor U5000 (N_5000,N_3816,N_3737);
or U5001 (N_5001,N_2667,N_3786);
xor U5002 (N_5002,N_3820,N_3494);
xnor U5003 (N_5003,N_3540,N_3430);
or U5004 (N_5004,N_3175,N_2392);
and U5005 (N_5005,N_3802,N_2856);
xor U5006 (N_5006,N_3909,N_2448);
and U5007 (N_5007,N_3968,N_3524);
nand U5008 (N_5008,N_3672,N_2665);
nor U5009 (N_5009,N_3558,N_2259);
xor U5010 (N_5010,N_3691,N_2761);
or U5011 (N_5011,N_3075,N_3646);
nor U5012 (N_5012,N_2608,N_3470);
or U5013 (N_5013,N_3298,N_2185);
and U5014 (N_5014,N_3163,N_3388);
and U5015 (N_5015,N_3196,N_3476);
xor U5016 (N_5016,N_2717,N_2152);
and U5017 (N_5017,N_3784,N_2629);
nand U5018 (N_5018,N_2436,N_2272);
xor U5019 (N_5019,N_3073,N_3009);
xor U5020 (N_5020,N_2852,N_3091);
nand U5021 (N_5021,N_3141,N_3243);
or U5022 (N_5022,N_3154,N_2997);
nand U5023 (N_5023,N_2727,N_2028);
xnor U5024 (N_5024,N_3340,N_3787);
nand U5025 (N_5025,N_3323,N_3658);
nand U5026 (N_5026,N_3176,N_2141);
and U5027 (N_5027,N_2910,N_2717);
xor U5028 (N_5028,N_2630,N_2146);
and U5029 (N_5029,N_3072,N_2906);
nor U5030 (N_5030,N_3755,N_2077);
or U5031 (N_5031,N_3342,N_3952);
nor U5032 (N_5032,N_3771,N_2955);
nand U5033 (N_5033,N_2517,N_2719);
or U5034 (N_5034,N_2395,N_3188);
nor U5035 (N_5035,N_2888,N_3042);
or U5036 (N_5036,N_3425,N_3544);
xor U5037 (N_5037,N_2226,N_3345);
or U5038 (N_5038,N_2646,N_3766);
nand U5039 (N_5039,N_2166,N_3942);
xnor U5040 (N_5040,N_3733,N_3816);
and U5041 (N_5041,N_3276,N_2845);
xnor U5042 (N_5042,N_3695,N_2913);
xor U5043 (N_5043,N_3078,N_3696);
and U5044 (N_5044,N_3500,N_3367);
and U5045 (N_5045,N_3186,N_2165);
xnor U5046 (N_5046,N_3023,N_2649);
nand U5047 (N_5047,N_3710,N_2521);
or U5048 (N_5048,N_2765,N_3424);
xor U5049 (N_5049,N_3957,N_3636);
xnor U5050 (N_5050,N_3405,N_3633);
nor U5051 (N_5051,N_2923,N_3460);
nor U5052 (N_5052,N_3023,N_3865);
nand U5053 (N_5053,N_2994,N_3543);
or U5054 (N_5054,N_3825,N_3140);
and U5055 (N_5055,N_3431,N_2300);
xnor U5056 (N_5056,N_2732,N_2139);
xnor U5057 (N_5057,N_3173,N_3544);
or U5058 (N_5058,N_2618,N_2227);
nor U5059 (N_5059,N_3276,N_3726);
xor U5060 (N_5060,N_3980,N_3226);
and U5061 (N_5061,N_3037,N_3947);
or U5062 (N_5062,N_2911,N_3034);
or U5063 (N_5063,N_3889,N_3784);
xnor U5064 (N_5064,N_2869,N_2274);
xnor U5065 (N_5065,N_2545,N_2742);
nand U5066 (N_5066,N_3447,N_2936);
nor U5067 (N_5067,N_2041,N_3804);
xor U5068 (N_5068,N_2728,N_2934);
or U5069 (N_5069,N_3914,N_3217);
nand U5070 (N_5070,N_3437,N_3482);
and U5071 (N_5071,N_3295,N_3474);
nand U5072 (N_5072,N_3570,N_3788);
and U5073 (N_5073,N_3252,N_2806);
nand U5074 (N_5074,N_2550,N_3765);
nand U5075 (N_5075,N_3707,N_2977);
and U5076 (N_5076,N_2907,N_3220);
xnor U5077 (N_5077,N_2109,N_3974);
nor U5078 (N_5078,N_3013,N_2965);
and U5079 (N_5079,N_2659,N_2560);
nand U5080 (N_5080,N_2253,N_2859);
and U5081 (N_5081,N_3909,N_3298);
nand U5082 (N_5082,N_3241,N_3985);
or U5083 (N_5083,N_3140,N_3933);
and U5084 (N_5084,N_3825,N_3487);
xor U5085 (N_5085,N_3801,N_2638);
nor U5086 (N_5086,N_3590,N_2559);
xor U5087 (N_5087,N_2895,N_2202);
nand U5088 (N_5088,N_3894,N_3381);
and U5089 (N_5089,N_3847,N_3789);
nand U5090 (N_5090,N_3082,N_3733);
nor U5091 (N_5091,N_2114,N_3132);
xor U5092 (N_5092,N_2509,N_3412);
nor U5093 (N_5093,N_3532,N_3979);
nand U5094 (N_5094,N_3391,N_2031);
nand U5095 (N_5095,N_3760,N_2723);
nor U5096 (N_5096,N_3697,N_2612);
nor U5097 (N_5097,N_2857,N_2498);
nor U5098 (N_5098,N_3257,N_2008);
nand U5099 (N_5099,N_2111,N_2186);
xor U5100 (N_5100,N_2937,N_3351);
and U5101 (N_5101,N_2986,N_3846);
and U5102 (N_5102,N_3466,N_3886);
xnor U5103 (N_5103,N_3297,N_3647);
nor U5104 (N_5104,N_2927,N_2219);
nor U5105 (N_5105,N_3361,N_2718);
and U5106 (N_5106,N_3627,N_3552);
nor U5107 (N_5107,N_3150,N_2223);
and U5108 (N_5108,N_3987,N_2294);
xor U5109 (N_5109,N_3551,N_3168);
or U5110 (N_5110,N_2360,N_3869);
or U5111 (N_5111,N_2287,N_2791);
or U5112 (N_5112,N_3178,N_2957);
or U5113 (N_5113,N_2344,N_3401);
nor U5114 (N_5114,N_2327,N_3609);
nand U5115 (N_5115,N_2437,N_2231);
xor U5116 (N_5116,N_3980,N_3555);
and U5117 (N_5117,N_2794,N_2529);
and U5118 (N_5118,N_3347,N_2806);
and U5119 (N_5119,N_3878,N_2710);
and U5120 (N_5120,N_2990,N_2257);
or U5121 (N_5121,N_3022,N_2689);
and U5122 (N_5122,N_2114,N_2584);
xnor U5123 (N_5123,N_3925,N_2026);
xnor U5124 (N_5124,N_2921,N_3476);
xor U5125 (N_5125,N_3919,N_3273);
and U5126 (N_5126,N_3692,N_3232);
nand U5127 (N_5127,N_3907,N_3126);
or U5128 (N_5128,N_3794,N_2962);
nand U5129 (N_5129,N_3706,N_2905);
nor U5130 (N_5130,N_3829,N_2341);
nor U5131 (N_5131,N_2983,N_2315);
or U5132 (N_5132,N_2645,N_2989);
nand U5133 (N_5133,N_3933,N_2130);
nand U5134 (N_5134,N_3685,N_3978);
nand U5135 (N_5135,N_2280,N_2238);
nor U5136 (N_5136,N_2943,N_3595);
or U5137 (N_5137,N_2569,N_3788);
and U5138 (N_5138,N_3719,N_3778);
nor U5139 (N_5139,N_2746,N_2729);
or U5140 (N_5140,N_3390,N_3227);
nand U5141 (N_5141,N_2770,N_3615);
xnor U5142 (N_5142,N_3096,N_3740);
xnor U5143 (N_5143,N_3704,N_2510);
and U5144 (N_5144,N_2597,N_2387);
nor U5145 (N_5145,N_3620,N_3512);
nor U5146 (N_5146,N_2809,N_2230);
xnor U5147 (N_5147,N_2222,N_3324);
xnor U5148 (N_5148,N_3677,N_2978);
and U5149 (N_5149,N_2768,N_2729);
or U5150 (N_5150,N_2248,N_3113);
or U5151 (N_5151,N_3325,N_2644);
or U5152 (N_5152,N_3153,N_2138);
or U5153 (N_5153,N_3085,N_2352);
nor U5154 (N_5154,N_2455,N_2504);
or U5155 (N_5155,N_2841,N_2507);
nand U5156 (N_5156,N_2517,N_2966);
nor U5157 (N_5157,N_2696,N_3199);
or U5158 (N_5158,N_3545,N_3054);
nor U5159 (N_5159,N_2746,N_3237);
xor U5160 (N_5160,N_3893,N_2732);
or U5161 (N_5161,N_3649,N_2645);
nor U5162 (N_5162,N_3592,N_3787);
and U5163 (N_5163,N_2127,N_3058);
and U5164 (N_5164,N_3290,N_2780);
xnor U5165 (N_5165,N_3236,N_3486);
and U5166 (N_5166,N_3368,N_3208);
nand U5167 (N_5167,N_3805,N_2220);
nand U5168 (N_5168,N_3220,N_2307);
nand U5169 (N_5169,N_3977,N_3766);
nand U5170 (N_5170,N_3187,N_2978);
and U5171 (N_5171,N_2214,N_2028);
xnor U5172 (N_5172,N_3458,N_3105);
nand U5173 (N_5173,N_3386,N_2069);
nor U5174 (N_5174,N_2949,N_2265);
xnor U5175 (N_5175,N_3051,N_3981);
and U5176 (N_5176,N_3056,N_2449);
nand U5177 (N_5177,N_3023,N_2415);
nand U5178 (N_5178,N_3803,N_2229);
nand U5179 (N_5179,N_3079,N_3306);
or U5180 (N_5180,N_2327,N_2399);
nor U5181 (N_5181,N_2597,N_2870);
xor U5182 (N_5182,N_2505,N_2402);
or U5183 (N_5183,N_3295,N_2027);
or U5184 (N_5184,N_3159,N_3921);
nand U5185 (N_5185,N_3458,N_2129);
or U5186 (N_5186,N_3544,N_2105);
and U5187 (N_5187,N_2521,N_3459);
nor U5188 (N_5188,N_2674,N_2991);
nand U5189 (N_5189,N_3145,N_3883);
or U5190 (N_5190,N_2468,N_3942);
xor U5191 (N_5191,N_3033,N_2300);
and U5192 (N_5192,N_2172,N_3596);
nand U5193 (N_5193,N_2103,N_3911);
xor U5194 (N_5194,N_3589,N_2981);
xor U5195 (N_5195,N_2348,N_2737);
nor U5196 (N_5196,N_2970,N_3394);
or U5197 (N_5197,N_3685,N_3303);
nand U5198 (N_5198,N_3115,N_2288);
nand U5199 (N_5199,N_2488,N_2461);
xor U5200 (N_5200,N_2672,N_3017);
nor U5201 (N_5201,N_3770,N_3343);
and U5202 (N_5202,N_3460,N_2469);
xor U5203 (N_5203,N_2114,N_2623);
nor U5204 (N_5204,N_3996,N_2902);
or U5205 (N_5205,N_3609,N_2871);
xnor U5206 (N_5206,N_2088,N_3275);
and U5207 (N_5207,N_2155,N_2381);
xnor U5208 (N_5208,N_2504,N_2186);
nor U5209 (N_5209,N_2787,N_2335);
xnor U5210 (N_5210,N_3367,N_2502);
and U5211 (N_5211,N_3506,N_3659);
and U5212 (N_5212,N_2313,N_3924);
or U5213 (N_5213,N_3971,N_2447);
or U5214 (N_5214,N_3768,N_2118);
nand U5215 (N_5215,N_2261,N_3571);
nand U5216 (N_5216,N_2242,N_2653);
nand U5217 (N_5217,N_2299,N_2677);
and U5218 (N_5218,N_3762,N_3137);
and U5219 (N_5219,N_3690,N_3663);
nand U5220 (N_5220,N_3805,N_2387);
nor U5221 (N_5221,N_2490,N_2089);
nand U5222 (N_5222,N_3616,N_2962);
xor U5223 (N_5223,N_2543,N_2615);
nand U5224 (N_5224,N_2455,N_2683);
nand U5225 (N_5225,N_2582,N_2767);
or U5226 (N_5226,N_2446,N_3072);
and U5227 (N_5227,N_3133,N_2926);
nor U5228 (N_5228,N_3876,N_2085);
nand U5229 (N_5229,N_3108,N_3715);
xnor U5230 (N_5230,N_2279,N_3341);
nand U5231 (N_5231,N_3614,N_3692);
xor U5232 (N_5232,N_2281,N_3628);
nand U5233 (N_5233,N_3549,N_2298);
nor U5234 (N_5234,N_3907,N_3376);
and U5235 (N_5235,N_2526,N_3997);
xor U5236 (N_5236,N_3179,N_2838);
xor U5237 (N_5237,N_3664,N_3150);
and U5238 (N_5238,N_2682,N_3396);
nand U5239 (N_5239,N_2128,N_3088);
or U5240 (N_5240,N_3210,N_2262);
nand U5241 (N_5241,N_2794,N_3107);
or U5242 (N_5242,N_2820,N_2389);
xor U5243 (N_5243,N_2240,N_3678);
and U5244 (N_5244,N_2280,N_3657);
nand U5245 (N_5245,N_3546,N_2815);
or U5246 (N_5246,N_3914,N_2463);
or U5247 (N_5247,N_2124,N_3609);
nand U5248 (N_5248,N_2238,N_3329);
or U5249 (N_5249,N_3825,N_2881);
xnor U5250 (N_5250,N_2631,N_2587);
or U5251 (N_5251,N_3388,N_2855);
or U5252 (N_5252,N_3894,N_2398);
nand U5253 (N_5253,N_3954,N_2537);
and U5254 (N_5254,N_2639,N_3024);
nand U5255 (N_5255,N_2471,N_3243);
nor U5256 (N_5256,N_3404,N_3583);
xor U5257 (N_5257,N_2511,N_3327);
nor U5258 (N_5258,N_3894,N_2547);
nor U5259 (N_5259,N_2783,N_2610);
or U5260 (N_5260,N_2195,N_2323);
or U5261 (N_5261,N_2007,N_2337);
and U5262 (N_5262,N_3239,N_3712);
and U5263 (N_5263,N_2176,N_2593);
nor U5264 (N_5264,N_2546,N_2225);
nor U5265 (N_5265,N_2138,N_3843);
or U5266 (N_5266,N_2983,N_3345);
or U5267 (N_5267,N_2719,N_2344);
nor U5268 (N_5268,N_2785,N_2237);
or U5269 (N_5269,N_3017,N_3423);
and U5270 (N_5270,N_2012,N_2125);
nor U5271 (N_5271,N_2497,N_2571);
xor U5272 (N_5272,N_2675,N_3160);
nor U5273 (N_5273,N_3230,N_2979);
or U5274 (N_5274,N_2086,N_3913);
or U5275 (N_5275,N_2339,N_3688);
nor U5276 (N_5276,N_3716,N_2299);
nand U5277 (N_5277,N_3100,N_2774);
nand U5278 (N_5278,N_2719,N_3687);
nand U5279 (N_5279,N_2121,N_3095);
nand U5280 (N_5280,N_3142,N_2777);
and U5281 (N_5281,N_3271,N_3245);
nor U5282 (N_5282,N_2429,N_3966);
xor U5283 (N_5283,N_2565,N_2761);
nand U5284 (N_5284,N_2871,N_3927);
xnor U5285 (N_5285,N_3043,N_2905);
and U5286 (N_5286,N_3676,N_2308);
or U5287 (N_5287,N_3413,N_2282);
or U5288 (N_5288,N_3848,N_3601);
nand U5289 (N_5289,N_3279,N_3669);
or U5290 (N_5290,N_2203,N_2222);
xor U5291 (N_5291,N_2723,N_3613);
nor U5292 (N_5292,N_3436,N_3553);
nand U5293 (N_5293,N_2090,N_2252);
xnor U5294 (N_5294,N_2216,N_2050);
nor U5295 (N_5295,N_3355,N_2633);
or U5296 (N_5296,N_3243,N_2692);
xnor U5297 (N_5297,N_3124,N_3176);
or U5298 (N_5298,N_2211,N_2234);
or U5299 (N_5299,N_3986,N_3672);
nand U5300 (N_5300,N_3367,N_2653);
and U5301 (N_5301,N_3311,N_2012);
and U5302 (N_5302,N_2918,N_3099);
and U5303 (N_5303,N_3928,N_3740);
nor U5304 (N_5304,N_2534,N_2201);
nand U5305 (N_5305,N_3406,N_2236);
or U5306 (N_5306,N_3277,N_2984);
or U5307 (N_5307,N_2445,N_2060);
nand U5308 (N_5308,N_2360,N_3770);
xnor U5309 (N_5309,N_2909,N_3948);
xnor U5310 (N_5310,N_2655,N_2821);
nor U5311 (N_5311,N_3882,N_3040);
and U5312 (N_5312,N_3751,N_3995);
and U5313 (N_5313,N_2763,N_3345);
xnor U5314 (N_5314,N_3087,N_3135);
xnor U5315 (N_5315,N_2011,N_3371);
xnor U5316 (N_5316,N_3861,N_3766);
or U5317 (N_5317,N_3073,N_2722);
nor U5318 (N_5318,N_2805,N_2860);
and U5319 (N_5319,N_3258,N_3644);
nand U5320 (N_5320,N_2509,N_2492);
xor U5321 (N_5321,N_3130,N_3676);
and U5322 (N_5322,N_3501,N_3072);
and U5323 (N_5323,N_2246,N_3088);
and U5324 (N_5324,N_2767,N_3446);
or U5325 (N_5325,N_3711,N_3147);
nand U5326 (N_5326,N_3460,N_3097);
nor U5327 (N_5327,N_2473,N_2361);
nor U5328 (N_5328,N_3111,N_2926);
nand U5329 (N_5329,N_3022,N_3820);
nand U5330 (N_5330,N_2716,N_2607);
xor U5331 (N_5331,N_3818,N_2345);
xor U5332 (N_5332,N_2500,N_3738);
xor U5333 (N_5333,N_2049,N_3145);
or U5334 (N_5334,N_3184,N_3023);
nor U5335 (N_5335,N_3538,N_3478);
and U5336 (N_5336,N_2982,N_2241);
or U5337 (N_5337,N_3209,N_3812);
nor U5338 (N_5338,N_3466,N_2713);
nand U5339 (N_5339,N_3136,N_3490);
nand U5340 (N_5340,N_3430,N_2869);
or U5341 (N_5341,N_2394,N_2741);
or U5342 (N_5342,N_3443,N_2639);
nor U5343 (N_5343,N_3244,N_3952);
or U5344 (N_5344,N_2238,N_3029);
xnor U5345 (N_5345,N_2473,N_3624);
xnor U5346 (N_5346,N_2430,N_3330);
xnor U5347 (N_5347,N_2778,N_3431);
xnor U5348 (N_5348,N_2251,N_2285);
nand U5349 (N_5349,N_2458,N_2696);
nor U5350 (N_5350,N_2927,N_2616);
and U5351 (N_5351,N_2653,N_2891);
nor U5352 (N_5352,N_3403,N_2206);
or U5353 (N_5353,N_3087,N_3088);
nand U5354 (N_5354,N_3103,N_3628);
xnor U5355 (N_5355,N_2634,N_2939);
nand U5356 (N_5356,N_2944,N_3070);
nor U5357 (N_5357,N_2608,N_2376);
and U5358 (N_5358,N_3857,N_3793);
nor U5359 (N_5359,N_3062,N_3539);
and U5360 (N_5360,N_3276,N_3950);
nor U5361 (N_5361,N_3618,N_2694);
nor U5362 (N_5362,N_3425,N_2552);
xnor U5363 (N_5363,N_3806,N_2684);
nand U5364 (N_5364,N_2200,N_3966);
xor U5365 (N_5365,N_3959,N_3979);
or U5366 (N_5366,N_3235,N_3145);
or U5367 (N_5367,N_2284,N_2379);
xor U5368 (N_5368,N_3732,N_3573);
or U5369 (N_5369,N_2464,N_2934);
nand U5370 (N_5370,N_2965,N_3436);
xnor U5371 (N_5371,N_2773,N_2011);
nor U5372 (N_5372,N_3478,N_2621);
nor U5373 (N_5373,N_3019,N_3972);
and U5374 (N_5374,N_3656,N_2314);
nand U5375 (N_5375,N_2353,N_3762);
nor U5376 (N_5376,N_2665,N_2682);
nor U5377 (N_5377,N_2930,N_2858);
and U5378 (N_5378,N_2544,N_3434);
xnor U5379 (N_5379,N_3999,N_2482);
xor U5380 (N_5380,N_3217,N_3545);
and U5381 (N_5381,N_2559,N_2700);
and U5382 (N_5382,N_2589,N_3350);
and U5383 (N_5383,N_3309,N_3123);
nor U5384 (N_5384,N_3532,N_3445);
or U5385 (N_5385,N_3071,N_3051);
nand U5386 (N_5386,N_2681,N_3953);
and U5387 (N_5387,N_3967,N_3278);
or U5388 (N_5388,N_3908,N_3303);
nand U5389 (N_5389,N_2128,N_3524);
nand U5390 (N_5390,N_3234,N_3887);
or U5391 (N_5391,N_2764,N_3119);
nand U5392 (N_5392,N_3178,N_2776);
or U5393 (N_5393,N_2943,N_3077);
and U5394 (N_5394,N_2940,N_2656);
or U5395 (N_5395,N_3863,N_2237);
nor U5396 (N_5396,N_2626,N_3098);
or U5397 (N_5397,N_2808,N_2516);
and U5398 (N_5398,N_3869,N_2128);
and U5399 (N_5399,N_3213,N_3145);
nand U5400 (N_5400,N_2810,N_2476);
nand U5401 (N_5401,N_2426,N_2659);
or U5402 (N_5402,N_2675,N_3919);
or U5403 (N_5403,N_2949,N_2095);
or U5404 (N_5404,N_2519,N_2378);
or U5405 (N_5405,N_2734,N_3249);
nand U5406 (N_5406,N_3265,N_2829);
xnor U5407 (N_5407,N_3690,N_3238);
nor U5408 (N_5408,N_3639,N_2528);
and U5409 (N_5409,N_3991,N_3137);
or U5410 (N_5410,N_3132,N_3115);
xor U5411 (N_5411,N_3629,N_3887);
xnor U5412 (N_5412,N_3085,N_3895);
nor U5413 (N_5413,N_2332,N_2687);
and U5414 (N_5414,N_2647,N_2756);
xor U5415 (N_5415,N_3714,N_3364);
or U5416 (N_5416,N_3490,N_3157);
and U5417 (N_5417,N_2489,N_3056);
nand U5418 (N_5418,N_2773,N_2754);
xnor U5419 (N_5419,N_2681,N_2510);
and U5420 (N_5420,N_2145,N_2218);
nor U5421 (N_5421,N_3267,N_2669);
and U5422 (N_5422,N_2418,N_2542);
xor U5423 (N_5423,N_2932,N_2289);
nor U5424 (N_5424,N_2806,N_3207);
nand U5425 (N_5425,N_3246,N_2045);
nand U5426 (N_5426,N_3686,N_2704);
xnor U5427 (N_5427,N_2562,N_3877);
nand U5428 (N_5428,N_3229,N_2734);
nor U5429 (N_5429,N_3714,N_2142);
nor U5430 (N_5430,N_3617,N_3187);
nor U5431 (N_5431,N_3373,N_2362);
xnor U5432 (N_5432,N_2940,N_3066);
nor U5433 (N_5433,N_3625,N_2001);
nand U5434 (N_5434,N_2877,N_3200);
nor U5435 (N_5435,N_2929,N_2559);
and U5436 (N_5436,N_2306,N_2291);
or U5437 (N_5437,N_3146,N_2982);
nand U5438 (N_5438,N_3484,N_3660);
nor U5439 (N_5439,N_2977,N_2198);
or U5440 (N_5440,N_2021,N_3668);
or U5441 (N_5441,N_3482,N_2829);
or U5442 (N_5442,N_2320,N_2544);
or U5443 (N_5443,N_3361,N_3817);
and U5444 (N_5444,N_2338,N_2393);
or U5445 (N_5445,N_2708,N_2819);
and U5446 (N_5446,N_2851,N_3481);
nand U5447 (N_5447,N_3518,N_3753);
nor U5448 (N_5448,N_2877,N_3934);
or U5449 (N_5449,N_3898,N_2720);
nor U5450 (N_5450,N_3208,N_3088);
nand U5451 (N_5451,N_3935,N_3705);
nor U5452 (N_5452,N_2937,N_2130);
nor U5453 (N_5453,N_3147,N_2415);
xnor U5454 (N_5454,N_3835,N_2874);
nand U5455 (N_5455,N_2034,N_3949);
nand U5456 (N_5456,N_3486,N_3754);
nand U5457 (N_5457,N_2630,N_2651);
and U5458 (N_5458,N_2516,N_2145);
nand U5459 (N_5459,N_2332,N_2952);
nand U5460 (N_5460,N_2625,N_3142);
nand U5461 (N_5461,N_2790,N_2085);
or U5462 (N_5462,N_2288,N_2555);
and U5463 (N_5463,N_3665,N_2094);
or U5464 (N_5464,N_3067,N_2754);
nand U5465 (N_5465,N_3516,N_2561);
nor U5466 (N_5466,N_3418,N_2404);
or U5467 (N_5467,N_3803,N_3749);
nor U5468 (N_5468,N_3144,N_3947);
nor U5469 (N_5469,N_2688,N_3183);
xor U5470 (N_5470,N_2964,N_2936);
and U5471 (N_5471,N_3192,N_2348);
or U5472 (N_5472,N_2557,N_3231);
xor U5473 (N_5473,N_2699,N_3641);
xnor U5474 (N_5474,N_2226,N_3629);
or U5475 (N_5475,N_3336,N_2324);
nor U5476 (N_5476,N_2487,N_3126);
nand U5477 (N_5477,N_3543,N_2899);
xnor U5478 (N_5478,N_2192,N_2410);
nor U5479 (N_5479,N_2333,N_2014);
or U5480 (N_5480,N_2331,N_2170);
and U5481 (N_5481,N_2621,N_3823);
or U5482 (N_5482,N_3183,N_2928);
or U5483 (N_5483,N_3776,N_3619);
or U5484 (N_5484,N_3496,N_3154);
or U5485 (N_5485,N_2635,N_2155);
or U5486 (N_5486,N_2968,N_2030);
or U5487 (N_5487,N_3179,N_2141);
and U5488 (N_5488,N_2391,N_2890);
and U5489 (N_5489,N_3035,N_3708);
or U5490 (N_5490,N_2918,N_2937);
nor U5491 (N_5491,N_3332,N_3626);
and U5492 (N_5492,N_2430,N_2266);
and U5493 (N_5493,N_2701,N_3100);
xor U5494 (N_5494,N_3683,N_3405);
and U5495 (N_5495,N_2832,N_2627);
nand U5496 (N_5496,N_3168,N_2512);
xor U5497 (N_5497,N_2978,N_2047);
nor U5498 (N_5498,N_3453,N_3154);
nand U5499 (N_5499,N_2175,N_2947);
and U5500 (N_5500,N_3980,N_2263);
xnor U5501 (N_5501,N_2009,N_2197);
nand U5502 (N_5502,N_2041,N_3024);
nor U5503 (N_5503,N_2636,N_2142);
and U5504 (N_5504,N_2825,N_2994);
and U5505 (N_5505,N_2433,N_2796);
nor U5506 (N_5506,N_3851,N_2694);
xor U5507 (N_5507,N_2832,N_3023);
or U5508 (N_5508,N_2785,N_2018);
and U5509 (N_5509,N_3077,N_2630);
and U5510 (N_5510,N_3790,N_3635);
and U5511 (N_5511,N_2254,N_3139);
or U5512 (N_5512,N_2344,N_3671);
nor U5513 (N_5513,N_3618,N_3405);
nor U5514 (N_5514,N_2682,N_2764);
or U5515 (N_5515,N_2822,N_2520);
or U5516 (N_5516,N_3545,N_3645);
nand U5517 (N_5517,N_3235,N_2970);
or U5518 (N_5518,N_2949,N_2434);
and U5519 (N_5519,N_3549,N_2714);
and U5520 (N_5520,N_3961,N_2984);
nand U5521 (N_5521,N_2328,N_2728);
and U5522 (N_5522,N_3341,N_2737);
nor U5523 (N_5523,N_3586,N_3246);
xor U5524 (N_5524,N_2996,N_3994);
nor U5525 (N_5525,N_2774,N_3013);
nand U5526 (N_5526,N_2937,N_3936);
nand U5527 (N_5527,N_2288,N_3448);
xor U5528 (N_5528,N_2183,N_2796);
nor U5529 (N_5529,N_3951,N_2229);
nor U5530 (N_5530,N_3287,N_2168);
xor U5531 (N_5531,N_3763,N_2838);
nor U5532 (N_5532,N_3741,N_2675);
and U5533 (N_5533,N_2822,N_3418);
nand U5534 (N_5534,N_2474,N_2217);
nor U5535 (N_5535,N_2077,N_3878);
or U5536 (N_5536,N_2860,N_2067);
nand U5537 (N_5537,N_2714,N_3942);
nand U5538 (N_5538,N_2603,N_3678);
or U5539 (N_5539,N_3371,N_3775);
nor U5540 (N_5540,N_3791,N_2227);
nor U5541 (N_5541,N_3883,N_3770);
xnor U5542 (N_5542,N_2569,N_2397);
xnor U5543 (N_5543,N_3205,N_2271);
and U5544 (N_5544,N_2807,N_2673);
or U5545 (N_5545,N_3009,N_3978);
nor U5546 (N_5546,N_3927,N_3770);
and U5547 (N_5547,N_2322,N_3736);
xor U5548 (N_5548,N_2880,N_3078);
xnor U5549 (N_5549,N_2156,N_3877);
xor U5550 (N_5550,N_2394,N_2513);
xnor U5551 (N_5551,N_2590,N_2325);
xnor U5552 (N_5552,N_2774,N_2155);
xnor U5553 (N_5553,N_3207,N_2465);
xnor U5554 (N_5554,N_2296,N_2686);
xor U5555 (N_5555,N_2456,N_2151);
nand U5556 (N_5556,N_3268,N_2481);
or U5557 (N_5557,N_3189,N_3332);
nor U5558 (N_5558,N_2847,N_3625);
and U5559 (N_5559,N_3700,N_3211);
xnor U5560 (N_5560,N_2678,N_3302);
and U5561 (N_5561,N_2641,N_2429);
xor U5562 (N_5562,N_2942,N_2196);
nor U5563 (N_5563,N_2775,N_2631);
nand U5564 (N_5564,N_3854,N_3017);
xnor U5565 (N_5565,N_2755,N_3396);
or U5566 (N_5566,N_3682,N_3859);
nand U5567 (N_5567,N_2627,N_2233);
and U5568 (N_5568,N_2666,N_3564);
and U5569 (N_5569,N_2817,N_3174);
xor U5570 (N_5570,N_2029,N_2609);
or U5571 (N_5571,N_2382,N_2580);
nor U5572 (N_5572,N_2876,N_3933);
and U5573 (N_5573,N_2197,N_2417);
nand U5574 (N_5574,N_3400,N_2830);
or U5575 (N_5575,N_2736,N_2606);
xnor U5576 (N_5576,N_3287,N_3251);
or U5577 (N_5577,N_3041,N_2558);
nand U5578 (N_5578,N_3478,N_3445);
nor U5579 (N_5579,N_3400,N_3472);
nor U5580 (N_5580,N_3079,N_3950);
or U5581 (N_5581,N_2622,N_3258);
nand U5582 (N_5582,N_3588,N_2647);
nor U5583 (N_5583,N_2300,N_3651);
nand U5584 (N_5584,N_3314,N_3108);
and U5585 (N_5585,N_3074,N_2830);
and U5586 (N_5586,N_2294,N_2396);
nor U5587 (N_5587,N_2866,N_3834);
nand U5588 (N_5588,N_3579,N_3811);
nand U5589 (N_5589,N_3187,N_3974);
or U5590 (N_5590,N_3960,N_3772);
or U5591 (N_5591,N_2985,N_3885);
or U5592 (N_5592,N_3146,N_3735);
nand U5593 (N_5593,N_3533,N_2656);
or U5594 (N_5594,N_2173,N_3454);
or U5595 (N_5595,N_2014,N_3789);
nand U5596 (N_5596,N_3508,N_3868);
nand U5597 (N_5597,N_2649,N_3837);
nand U5598 (N_5598,N_3362,N_2984);
and U5599 (N_5599,N_2723,N_2376);
or U5600 (N_5600,N_2603,N_3945);
xnor U5601 (N_5601,N_3621,N_3234);
nor U5602 (N_5602,N_3218,N_3984);
xnor U5603 (N_5603,N_2439,N_3485);
nor U5604 (N_5604,N_2946,N_2655);
and U5605 (N_5605,N_2350,N_2840);
nand U5606 (N_5606,N_3091,N_2760);
or U5607 (N_5607,N_2090,N_3231);
nand U5608 (N_5608,N_2366,N_3626);
nand U5609 (N_5609,N_3679,N_3327);
nor U5610 (N_5610,N_2892,N_3941);
or U5611 (N_5611,N_3129,N_3445);
and U5612 (N_5612,N_3060,N_3728);
or U5613 (N_5613,N_3308,N_3128);
xnor U5614 (N_5614,N_2816,N_2118);
and U5615 (N_5615,N_3085,N_3388);
nor U5616 (N_5616,N_3907,N_3453);
and U5617 (N_5617,N_2246,N_3638);
nor U5618 (N_5618,N_3446,N_2486);
and U5619 (N_5619,N_2688,N_3187);
or U5620 (N_5620,N_3572,N_3887);
and U5621 (N_5621,N_3301,N_2157);
xor U5622 (N_5622,N_2921,N_2552);
nand U5623 (N_5623,N_2328,N_3356);
xnor U5624 (N_5624,N_3571,N_3858);
or U5625 (N_5625,N_3025,N_2731);
or U5626 (N_5626,N_3664,N_3529);
or U5627 (N_5627,N_2947,N_2211);
xor U5628 (N_5628,N_3538,N_2795);
and U5629 (N_5629,N_2488,N_3169);
and U5630 (N_5630,N_3083,N_3651);
and U5631 (N_5631,N_2906,N_3969);
and U5632 (N_5632,N_2977,N_2672);
and U5633 (N_5633,N_3397,N_3914);
and U5634 (N_5634,N_3715,N_3718);
nand U5635 (N_5635,N_3258,N_3468);
xor U5636 (N_5636,N_2122,N_2841);
nand U5637 (N_5637,N_3841,N_3790);
and U5638 (N_5638,N_3142,N_3447);
xnor U5639 (N_5639,N_2531,N_2248);
and U5640 (N_5640,N_3725,N_3890);
and U5641 (N_5641,N_3452,N_2670);
nor U5642 (N_5642,N_2722,N_3321);
xor U5643 (N_5643,N_3917,N_3988);
and U5644 (N_5644,N_2832,N_2707);
nor U5645 (N_5645,N_3789,N_3861);
nand U5646 (N_5646,N_3048,N_2028);
or U5647 (N_5647,N_3248,N_3450);
nor U5648 (N_5648,N_3481,N_3111);
and U5649 (N_5649,N_2229,N_3786);
xor U5650 (N_5650,N_3800,N_3360);
xor U5651 (N_5651,N_3427,N_2707);
xnor U5652 (N_5652,N_3449,N_2473);
xor U5653 (N_5653,N_3235,N_2999);
and U5654 (N_5654,N_3835,N_2988);
nor U5655 (N_5655,N_2829,N_3869);
or U5656 (N_5656,N_3553,N_2988);
and U5657 (N_5657,N_3742,N_3193);
and U5658 (N_5658,N_2220,N_3450);
and U5659 (N_5659,N_3646,N_3113);
nand U5660 (N_5660,N_3275,N_3079);
xnor U5661 (N_5661,N_2955,N_3348);
nor U5662 (N_5662,N_2221,N_3032);
nand U5663 (N_5663,N_2127,N_3661);
or U5664 (N_5664,N_3438,N_2658);
xor U5665 (N_5665,N_3358,N_2523);
nand U5666 (N_5666,N_3129,N_2828);
and U5667 (N_5667,N_2454,N_2518);
nor U5668 (N_5668,N_2799,N_2702);
or U5669 (N_5669,N_2437,N_3796);
nor U5670 (N_5670,N_3042,N_2674);
or U5671 (N_5671,N_3339,N_3652);
or U5672 (N_5672,N_3203,N_2621);
nor U5673 (N_5673,N_3264,N_2260);
nor U5674 (N_5674,N_2216,N_3285);
nor U5675 (N_5675,N_3300,N_3249);
xor U5676 (N_5676,N_2086,N_2857);
and U5677 (N_5677,N_2259,N_2012);
nand U5678 (N_5678,N_2254,N_3964);
nor U5679 (N_5679,N_3646,N_3848);
nor U5680 (N_5680,N_3498,N_2467);
or U5681 (N_5681,N_3500,N_2154);
and U5682 (N_5682,N_2454,N_2755);
and U5683 (N_5683,N_2419,N_2180);
nor U5684 (N_5684,N_3579,N_3666);
or U5685 (N_5685,N_2195,N_3615);
nand U5686 (N_5686,N_2540,N_3862);
nand U5687 (N_5687,N_2782,N_2000);
or U5688 (N_5688,N_3950,N_2833);
and U5689 (N_5689,N_3273,N_2680);
nand U5690 (N_5690,N_3105,N_2396);
nand U5691 (N_5691,N_2900,N_3108);
nand U5692 (N_5692,N_2065,N_3993);
or U5693 (N_5693,N_3641,N_2755);
xor U5694 (N_5694,N_2578,N_2005);
nand U5695 (N_5695,N_2272,N_3321);
xnor U5696 (N_5696,N_2909,N_3215);
nor U5697 (N_5697,N_2377,N_2050);
nand U5698 (N_5698,N_3884,N_3045);
nand U5699 (N_5699,N_2606,N_3485);
or U5700 (N_5700,N_2645,N_2026);
or U5701 (N_5701,N_2853,N_2410);
and U5702 (N_5702,N_2566,N_2660);
nor U5703 (N_5703,N_3459,N_3203);
nor U5704 (N_5704,N_3905,N_2548);
nor U5705 (N_5705,N_3501,N_3085);
or U5706 (N_5706,N_3721,N_2574);
and U5707 (N_5707,N_3782,N_2567);
and U5708 (N_5708,N_3204,N_2981);
and U5709 (N_5709,N_2400,N_2403);
and U5710 (N_5710,N_2731,N_3102);
and U5711 (N_5711,N_2599,N_2269);
nor U5712 (N_5712,N_2808,N_3977);
nor U5713 (N_5713,N_3716,N_3265);
xnor U5714 (N_5714,N_3172,N_2219);
nor U5715 (N_5715,N_2860,N_3808);
and U5716 (N_5716,N_2457,N_3895);
and U5717 (N_5717,N_2341,N_3267);
or U5718 (N_5718,N_2096,N_3986);
nor U5719 (N_5719,N_2665,N_3307);
nand U5720 (N_5720,N_3270,N_3693);
nand U5721 (N_5721,N_3713,N_2850);
nand U5722 (N_5722,N_2598,N_3686);
and U5723 (N_5723,N_2555,N_3532);
and U5724 (N_5724,N_3618,N_2283);
xnor U5725 (N_5725,N_2999,N_3054);
xnor U5726 (N_5726,N_3633,N_3065);
and U5727 (N_5727,N_3711,N_2514);
nand U5728 (N_5728,N_3853,N_3961);
xnor U5729 (N_5729,N_2615,N_3365);
xnor U5730 (N_5730,N_2659,N_3644);
nand U5731 (N_5731,N_3995,N_2315);
nor U5732 (N_5732,N_2239,N_3700);
nor U5733 (N_5733,N_3434,N_2985);
nand U5734 (N_5734,N_3974,N_3088);
xnor U5735 (N_5735,N_2099,N_2108);
xnor U5736 (N_5736,N_2151,N_3133);
or U5737 (N_5737,N_2037,N_3628);
or U5738 (N_5738,N_3631,N_2089);
and U5739 (N_5739,N_2974,N_2729);
and U5740 (N_5740,N_2213,N_2918);
xor U5741 (N_5741,N_3091,N_2466);
xnor U5742 (N_5742,N_3066,N_2881);
nand U5743 (N_5743,N_2835,N_3858);
or U5744 (N_5744,N_2500,N_2192);
nand U5745 (N_5745,N_2250,N_3654);
xor U5746 (N_5746,N_2197,N_2133);
xor U5747 (N_5747,N_2891,N_3540);
and U5748 (N_5748,N_3253,N_2026);
or U5749 (N_5749,N_3421,N_2127);
nand U5750 (N_5750,N_2287,N_3499);
xor U5751 (N_5751,N_3896,N_3082);
and U5752 (N_5752,N_2426,N_3440);
nand U5753 (N_5753,N_3981,N_3923);
or U5754 (N_5754,N_3340,N_2929);
or U5755 (N_5755,N_2320,N_3745);
nor U5756 (N_5756,N_3852,N_2419);
nand U5757 (N_5757,N_3477,N_2150);
xor U5758 (N_5758,N_2747,N_3220);
nand U5759 (N_5759,N_2734,N_2032);
xor U5760 (N_5760,N_3002,N_3791);
and U5761 (N_5761,N_3600,N_2723);
or U5762 (N_5762,N_2680,N_2053);
or U5763 (N_5763,N_3399,N_3034);
nor U5764 (N_5764,N_3946,N_3980);
nand U5765 (N_5765,N_3141,N_3875);
nor U5766 (N_5766,N_2691,N_2369);
nand U5767 (N_5767,N_3336,N_3058);
nand U5768 (N_5768,N_2073,N_3238);
nor U5769 (N_5769,N_2922,N_3045);
nand U5770 (N_5770,N_3663,N_2908);
and U5771 (N_5771,N_2288,N_3106);
xnor U5772 (N_5772,N_3822,N_2149);
xor U5773 (N_5773,N_3510,N_2645);
nand U5774 (N_5774,N_2377,N_2898);
or U5775 (N_5775,N_3873,N_2777);
or U5776 (N_5776,N_2270,N_3306);
nand U5777 (N_5777,N_2980,N_3686);
xor U5778 (N_5778,N_2488,N_2964);
xnor U5779 (N_5779,N_3392,N_2325);
and U5780 (N_5780,N_3481,N_3671);
nand U5781 (N_5781,N_2779,N_3545);
or U5782 (N_5782,N_2245,N_2047);
nand U5783 (N_5783,N_2273,N_2777);
xnor U5784 (N_5784,N_3925,N_2414);
and U5785 (N_5785,N_2978,N_2443);
nand U5786 (N_5786,N_2394,N_3310);
nand U5787 (N_5787,N_3135,N_2549);
nand U5788 (N_5788,N_3444,N_2623);
and U5789 (N_5789,N_3031,N_3011);
nand U5790 (N_5790,N_3976,N_3545);
nand U5791 (N_5791,N_3780,N_2936);
and U5792 (N_5792,N_3643,N_2419);
nor U5793 (N_5793,N_3160,N_2749);
or U5794 (N_5794,N_3375,N_2862);
nand U5795 (N_5795,N_3210,N_2270);
and U5796 (N_5796,N_3998,N_2420);
xor U5797 (N_5797,N_2818,N_3287);
xor U5798 (N_5798,N_2770,N_3565);
xor U5799 (N_5799,N_3730,N_2713);
xor U5800 (N_5800,N_3246,N_3716);
nand U5801 (N_5801,N_3352,N_2178);
nand U5802 (N_5802,N_2809,N_2759);
and U5803 (N_5803,N_2094,N_2046);
or U5804 (N_5804,N_3398,N_3961);
nand U5805 (N_5805,N_3710,N_3019);
or U5806 (N_5806,N_2822,N_3112);
or U5807 (N_5807,N_2203,N_3389);
xor U5808 (N_5808,N_3014,N_2561);
or U5809 (N_5809,N_2573,N_3023);
nand U5810 (N_5810,N_2404,N_3927);
nand U5811 (N_5811,N_2961,N_2587);
nand U5812 (N_5812,N_3159,N_3422);
or U5813 (N_5813,N_2569,N_2060);
and U5814 (N_5814,N_2868,N_2430);
xor U5815 (N_5815,N_2493,N_3621);
and U5816 (N_5816,N_2546,N_3500);
nor U5817 (N_5817,N_3307,N_3340);
xor U5818 (N_5818,N_3857,N_2323);
nor U5819 (N_5819,N_3102,N_2982);
nand U5820 (N_5820,N_3139,N_2557);
and U5821 (N_5821,N_3790,N_3468);
nor U5822 (N_5822,N_3083,N_2376);
nor U5823 (N_5823,N_2983,N_3990);
or U5824 (N_5824,N_3402,N_3686);
nor U5825 (N_5825,N_2316,N_3763);
nor U5826 (N_5826,N_3484,N_3597);
and U5827 (N_5827,N_3468,N_2793);
xnor U5828 (N_5828,N_2430,N_2166);
xnor U5829 (N_5829,N_2588,N_2481);
nor U5830 (N_5830,N_3142,N_3170);
nand U5831 (N_5831,N_2137,N_2487);
or U5832 (N_5832,N_2599,N_2535);
nor U5833 (N_5833,N_2468,N_2987);
and U5834 (N_5834,N_2200,N_2961);
xnor U5835 (N_5835,N_3770,N_2821);
nand U5836 (N_5836,N_3659,N_2175);
nor U5837 (N_5837,N_3710,N_3190);
nand U5838 (N_5838,N_2210,N_2172);
and U5839 (N_5839,N_3584,N_2813);
and U5840 (N_5840,N_2512,N_2464);
and U5841 (N_5841,N_2947,N_2909);
or U5842 (N_5842,N_3784,N_2374);
or U5843 (N_5843,N_3203,N_2660);
xor U5844 (N_5844,N_2814,N_3728);
nor U5845 (N_5845,N_2393,N_3619);
nor U5846 (N_5846,N_3615,N_3505);
xor U5847 (N_5847,N_3354,N_2496);
or U5848 (N_5848,N_3244,N_2003);
and U5849 (N_5849,N_3912,N_3546);
or U5850 (N_5850,N_2852,N_2001);
nand U5851 (N_5851,N_3444,N_2890);
nor U5852 (N_5852,N_2367,N_3145);
xor U5853 (N_5853,N_2551,N_2743);
xor U5854 (N_5854,N_2190,N_3659);
nor U5855 (N_5855,N_3887,N_2877);
and U5856 (N_5856,N_2797,N_2431);
and U5857 (N_5857,N_3671,N_2386);
nand U5858 (N_5858,N_3639,N_2740);
nor U5859 (N_5859,N_2422,N_3020);
and U5860 (N_5860,N_2014,N_2629);
nand U5861 (N_5861,N_2078,N_3352);
nand U5862 (N_5862,N_2592,N_2686);
nand U5863 (N_5863,N_2195,N_3927);
or U5864 (N_5864,N_2709,N_2670);
or U5865 (N_5865,N_3045,N_3722);
xor U5866 (N_5866,N_2619,N_3650);
or U5867 (N_5867,N_3254,N_3140);
nand U5868 (N_5868,N_2196,N_3593);
and U5869 (N_5869,N_2822,N_2688);
nor U5870 (N_5870,N_3230,N_2218);
nand U5871 (N_5871,N_2714,N_3711);
xnor U5872 (N_5872,N_3600,N_2910);
xor U5873 (N_5873,N_2949,N_2072);
nor U5874 (N_5874,N_2950,N_3681);
nand U5875 (N_5875,N_2671,N_2461);
or U5876 (N_5876,N_3551,N_2657);
nand U5877 (N_5877,N_2306,N_2410);
xor U5878 (N_5878,N_2369,N_2113);
or U5879 (N_5879,N_2659,N_2073);
and U5880 (N_5880,N_2032,N_3529);
and U5881 (N_5881,N_2108,N_3206);
or U5882 (N_5882,N_3676,N_3524);
and U5883 (N_5883,N_3003,N_2448);
xor U5884 (N_5884,N_2586,N_2246);
nand U5885 (N_5885,N_2837,N_2904);
or U5886 (N_5886,N_3388,N_2632);
and U5887 (N_5887,N_3190,N_3819);
and U5888 (N_5888,N_2334,N_2721);
and U5889 (N_5889,N_3851,N_3849);
nor U5890 (N_5890,N_2241,N_2108);
nand U5891 (N_5891,N_3075,N_2347);
nor U5892 (N_5892,N_2406,N_2765);
xor U5893 (N_5893,N_3656,N_2323);
xnor U5894 (N_5894,N_2374,N_3270);
nand U5895 (N_5895,N_2714,N_3720);
nor U5896 (N_5896,N_2776,N_2635);
nor U5897 (N_5897,N_3630,N_2538);
nor U5898 (N_5898,N_3132,N_2132);
xor U5899 (N_5899,N_2243,N_3603);
nor U5900 (N_5900,N_3891,N_2195);
nor U5901 (N_5901,N_3619,N_3700);
nor U5902 (N_5902,N_3408,N_2172);
and U5903 (N_5903,N_3422,N_3338);
and U5904 (N_5904,N_2781,N_2770);
nand U5905 (N_5905,N_2426,N_2918);
xnor U5906 (N_5906,N_2658,N_2057);
xnor U5907 (N_5907,N_3427,N_3960);
or U5908 (N_5908,N_2426,N_2291);
nand U5909 (N_5909,N_3780,N_2844);
xnor U5910 (N_5910,N_3370,N_2846);
or U5911 (N_5911,N_2120,N_3295);
nor U5912 (N_5912,N_2039,N_2296);
or U5913 (N_5913,N_2491,N_3894);
nor U5914 (N_5914,N_3818,N_3225);
nor U5915 (N_5915,N_2976,N_2205);
nand U5916 (N_5916,N_2166,N_2425);
nor U5917 (N_5917,N_2105,N_2690);
nand U5918 (N_5918,N_3925,N_3579);
and U5919 (N_5919,N_2685,N_3708);
xor U5920 (N_5920,N_2724,N_2219);
nor U5921 (N_5921,N_3049,N_3133);
nand U5922 (N_5922,N_2428,N_2374);
nand U5923 (N_5923,N_3547,N_2255);
nand U5924 (N_5924,N_3420,N_3849);
nor U5925 (N_5925,N_2367,N_2782);
nand U5926 (N_5926,N_3719,N_3121);
xnor U5927 (N_5927,N_2392,N_3220);
nor U5928 (N_5928,N_2753,N_2250);
or U5929 (N_5929,N_3385,N_3457);
nand U5930 (N_5930,N_2876,N_3870);
nand U5931 (N_5931,N_3798,N_3556);
and U5932 (N_5932,N_3460,N_2048);
nor U5933 (N_5933,N_3419,N_3784);
and U5934 (N_5934,N_3148,N_2252);
or U5935 (N_5935,N_2080,N_3896);
nor U5936 (N_5936,N_2923,N_3404);
and U5937 (N_5937,N_2353,N_3257);
xnor U5938 (N_5938,N_2946,N_3144);
nor U5939 (N_5939,N_3417,N_2402);
nor U5940 (N_5940,N_3621,N_2925);
xnor U5941 (N_5941,N_3296,N_3119);
xor U5942 (N_5942,N_2670,N_3240);
nor U5943 (N_5943,N_3380,N_2423);
and U5944 (N_5944,N_3520,N_3555);
and U5945 (N_5945,N_3438,N_2092);
or U5946 (N_5946,N_2962,N_2093);
nand U5947 (N_5947,N_3835,N_2108);
xor U5948 (N_5948,N_2689,N_3556);
and U5949 (N_5949,N_2562,N_2347);
xor U5950 (N_5950,N_3814,N_3707);
xnor U5951 (N_5951,N_2928,N_2693);
nor U5952 (N_5952,N_3366,N_2398);
and U5953 (N_5953,N_3083,N_3100);
nor U5954 (N_5954,N_3361,N_3233);
xnor U5955 (N_5955,N_2343,N_2109);
nand U5956 (N_5956,N_3029,N_2872);
xor U5957 (N_5957,N_3626,N_2269);
nor U5958 (N_5958,N_2905,N_3569);
and U5959 (N_5959,N_3694,N_3839);
or U5960 (N_5960,N_2097,N_2461);
or U5961 (N_5961,N_3942,N_3120);
or U5962 (N_5962,N_3740,N_3641);
or U5963 (N_5963,N_3781,N_2185);
xor U5964 (N_5964,N_3432,N_2239);
xor U5965 (N_5965,N_3121,N_3145);
xor U5966 (N_5966,N_3554,N_2935);
nand U5967 (N_5967,N_2963,N_3817);
nor U5968 (N_5968,N_3577,N_3268);
nand U5969 (N_5969,N_2401,N_2548);
nand U5970 (N_5970,N_2338,N_2054);
and U5971 (N_5971,N_3252,N_2449);
xor U5972 (N_5972,N_3497,N_3825);
nor U5973 (N_5973,N_3889,N_2190);
xor U5974 (N_5974,N_3547,N_3425);
nor U5975 (N_5975,N_2109,N_3649);
xnor U5976 (N_5976,N_2797,N_3124);
nand U5977 (N_5977,N_3185,N_3907);
nor U5978 (N_5978,N_3366,N_2992);
and U5979 (N_5979,N_3464,N_2430);
xor U5980 (N_5980,N_3462,N_2154);
or U5981 (N_5981,N_3842,N_2881);
and U5982 (N_5982,N_2320,N_3802);
or U5983 (N_5983,N_3185,N_3044);
nor U5984 (N_5984,N_2796,N_3522);
nand U5985 (N_5985,N_2603,N_3175);
or U5986 (N_5986,N_3298,N_2791);
xnor U5987 (N_5987,N_2255,N_2870);
and U5988 (N_5988,N_3864,N_2616);
and U5989 (N_5989,N_3288,N_3335);
nor U5990 (N_5990,N_2607,N_2055);
xnor U5991 (N_5991,N_3035,N_2923);
nand U5992 (N_5992,N_2791,N_3591);
and U5993 (N_5993,N_2061,N_3256);
xor U5994 (N_5994,N_3959,N_2649);
or U5995 (N_5995,N_2962,N_3160);
nand U5996 (N_5996,N_2616,N_2391);
or U5997 (N_5997,N_3586,N_3692);
nor U5998 (N_5998,N_2830,N_3670);
and U5999 (N_5999,N_2232,N_3899);
and U6000 (N_6000,N_4267,N_4439);
or U6001 (N_6001,N_5857,N_4612);
xor U6002 (N_6002,N_5100,N_5845);
and U6003 (N_6003,N_4356,N_5583);
and U6004 (N_6004,N_5682,N_4746);
or U6005 (N_6005,N_5210,N_4374);
xor U6006 (N_6006,N_4655,N_4384);
and U6007 (N_6007,N_4838,N_4254);
or U6008 (N_6008,N_5205,N_4240);
nor U6009 (N_6009,N_4306,N_4079);
nor U6010 (N_6010,N_5843,N_5971);
and U6011 (N_6011,N_4493,N_5495);
nand U6012 (N_6012,N_4429,N_4408);
xor U6013 (N_6013,N_4728,N_5946);
and U6014 (N_6014,N_5496,N_5123);
or U6015 (N_6015,N_4435,N_4665);
nand U6016 (N_6016,N_5372,N_5860);
nor U6017 (N_6017,N_4709,N_4901);
and U6018 (N_6018,N_4874,N_5368);
nor U6019 (N_6019,N_5671,N_5085);
nor U6020 (N_6020,N_4363,N_4480);
or U6021 (N_6021,N_5806,N_4636);
nand U6022 (N_6022,N_5624,N_4689);
nor U6023 (N_6023,N_5509,N_5535);
and U6024 (N_6024,N_5244,N_4292);
nand U6025 (N_6025,N_4073,N_4335);
xnor U6026 (N_6026,N_4872,N_4390);
xnor U6027 (N_6027,N_5579,N_5033);
xnor U6028 (N_6028,N_5343,N_5842);
and U6029 (N_6029,N_4725,N_5730);
nor U6030 (N_6030,N_4446,N_4772);
nor U6031 (N_6031,N_5111,N_4692);
xnor U6032 (N_6032,N_5555,N_5022);
xnor U6033 (N_6033,N_5737,N_4150);
nand U6034 (N_6034,N_5596,N_5177);
or U6035 (N_6035,N_5020,N_5136);
nand U6036 (N_6036,N_5521,N_5872);
xnor U6037 (N_6037,N_5018,N_4332);
and U6038 (N_6038,N_5571,N_4940);
nor U6039 (N_6039,N_4337,N_4017);
xor U6040 (N_6040,N_4207,N_5969);
nand U6041 (N_6041,N_4540,N_5537);
nand U6042 (N_6042,N_4633,N_4794);
nand U6043 (N_6043,N_5303,N_5081);
nand U6044 (N_6044,N_4591,N_4600);
or U6045 (N_6045,N_4066,N_4127);
or U6046 (N_6046,N_5246,N_4237);
or U6047 (N_6047,N_5327,N_5601);
xor U6048 (N_6048,N_4737,N_5217);
or U6049 (N_6049,N_4536,N_5121);
nor U6050 (N_6050,N_4625,N_4830);
or U6051 (N_6051,N_4022,N_5153);
nor U6052 (N_6052,N_4667,N_5347);
or U6053 (N_6053,N_4648,N_4382);
or U6054 (N_6054,N_4474,N_4489);
nor U6055 (N_6055,N_4327,N_4690);
xor U6056 (N_6056,N_4112,N_4657);
xor U6057 (N_6057,N_5215,N_4557);
and U6058 (N_6058,N_4727,N_5065);
and U6059 (N_6059,N_4232,N_4302);
xnor U6060 (N_6060,N_4119,N_4915);
nand U6061 (N_6061,N_5344,N_4683);
nor U6062 (N_6062,N_5181,N_4475);
xor U6063 (N_6063,N_5233,N_4851);
nand U6064 (N_6064,N_5900,N_4279);
or U6065 (N_6065,N_5798,N_4551);
nand U6066 (N_6066,N_5300,N_4831);
nand U6067 (N_6067,N_4009,N_5278);
or U6068 (N_6068,N_5649,N_5142);
and U6069 (N_6069,N_5286,N_4021);
and U6070 (N_6070,N_5744,N_4849);
nor U6071 (N_6071,N_4415,N_5106);
nor U6072 (N_6072,N_5049,N_5876);
and U6073 (N_6073,N_5885,N_4740);
nor U6074 (N_6074,N_4959,N_4710);
xnor U6075 (N_6075,N_5625,N_5301);
and U6076 (N_6076,N_5058,N_5166);
or U6077 (N_6077,N_5441,N_5784);
nor U6078 (N_6078,N_5013,N_5680);
nand U6079 (N_6079,N_5720,N_5428);
xor U6080 (N_6080,N_5965,N_5665);
nor U6081 (N_6081,N_5200,N_4804);
nor U6082 (N_6082,N_4873,N_5848);
nor U6083 (N_6083,N_5975,N_4847);
nand U6084 (N_6084,N_4205,N_4993);
nand U6085 (N_6085,N_4140,N_4920);
and U6086 (N_6086,N_5526,N_5283);
xnor U6087 (N_6087,N_4441,N_4258);
nor U6088 (N_6088,N_4266,N_4013);
or U6089 (N_6089,N_4425,N_5588);
nand U6090 (N_6090,N_4360,N_5002);
nor U6091 (N_6091,N_5641,N_4063);
nor U6092 (N_6092,N_5414,N_4183);
or U6093 (N_6093,N_5140,N_5145);
nor U6094 (N_6094,N_4813,N_4691);
xnor U6095 (N_6095,N_4860,N_4752);
nor U6096 (N_6096,N_4743,N_5174);
nor U6097 (N_6097,N_5718,N_5925);
nand U6098 (N_6098,N_4513,N_4229);
nand U6099 (N_6099,N_4914,N_4679);
and U6100 (N_6100,N_5775,N_4913);
or U6101 (N_6101,N_4724,N_4840);
or U6102 (N_6102,N_4147,N_5739);
nand U6103 (N_6103,N_5189,N_4869);
nor U6104 (N_6104,N_5948,N_4133);
or U6105 (N_6105,N_4464,N_4190);
xnor U6106 (N_6106,N_4179,N_4385);
nor U6107 (N_6107,N_4865,N_4260);
and U6108 (N_6108,N_5893,N_5619);
nand U6109 (N_6109,N_5547,N_5817);
or U6110 (N_6110,N_5989,N_4652);
nor U6111 (N_6111,N_5460,N_5960);
nand U6112 (N_6112,N_4589,N_5406);
or U6113 (N_6113,N_4854,N_5201);
nor U6114 (N_6114,N_5991,N_4399);
nor U6115 (N_6115,N_5556,N_5810);
or U6116 (N_6116,N_4421,N_4841);
xnor U6117 (N_6117,N_5685,N_4729);
xor U6118 (N_6118,N_5855,N_5875);
nand U6119 (N_6119,N_5059,N_4387);
nor U6120 (N_6120,N_4388,N_5239);
nor U6121 (N_6121,N_4981,N_4074);
xor U6122 (N_6122,N_5729,N_5191);
nor U6123 (N_6123,N_5563,N_4383);
or U6124 (N_6124,N_5748,N_4918);
nand U6125 (N_6125,N_5019,N_5006);
nand U6126 (N_6126,N_4686,N_5915);
nand U6127 (N_6127,N_5334,N_5150);
xor U6128 (N_6128,N_5773,N_5903);
or U6129 (N_6129,N_4580,N_5771);
nand U6130 (N_6130,N_4814,N_5149);
nor U6131 (N_6131,N_4644,N_5356);
nand U6132 (N_6132,N_4823,N_4701);
or U6133 (N_6133,N_5178,N_5733);
nand U6134 (N_6134,N_5417,N_4058);
or U6135 (N_6135,N_5035,N_4542);
nor U6136 (N_6136,N_4396,N_5467);
or U6137 (N_6137,N_5287,N_4333);
or U6138 (N_6138,N_4836,N_4635);
nand U6139 (N_6139,N_4738,N_5724);
and U6140 (N_6140,N_4601,N_4694);
nor U6141 (N_6141,N_5905,N_5118);
or U6142 (N_6142,N_5726,N_4085);
or U6143 (N_6143,N_5346,N_4817);
and U6144 (N_6144,N_5949,N_4811);
and U6145 (N_6145,N_5310,N_4307);
nand U6146 (N_6146,N_4111,N_4379);
and U6147 (N_6147,N_5216,N_4257);
or U6148 (N_6148,N_5632,N_4026);
or U6149 (N_6149,N_5740,N_5812);
nand U6150 (N_6150,N_5955,N_5886);
xnor U6151 (N_6151,N_4771,N_4929);
nand U6152 (N_6152,N_5398,N_5599);
and U6153 (N_6153,N_4592,N_4708);
or U6154 (N_6154,N_4016,N_5389);
and U6155 (N_6155,N_4883,N_5912);
and U6156 (N_6156,N_4410,N_4569);
or U6157 (N_6157,N_4990,N_4061);
and U6158 (N_6158,N_4001,N_4007);
nor U6159 (N_6159,N_5137,N_4622);
and U6160 (N_6160,N_4336,N_5466);
nor U6161 (N_6161,N_4904,N_4977);
or U6162 (N_6162,N_5034,N_5404);
and U6163 (N_6163,N_4653,N_4141);
nor U6164 (N_6164,N_4104,N_5274);
xor U6165 (N_6165,N_4039,N_4576);
nand U6166 (N_6166,N_5306,N_4145);
or U6167 (N_6167,N_4351,N_5318);
nor U6168 (N_6168,N_5281,N_5182);
xnor U6169 (N_6169,N_4443,N_5209);
nand U6170 (N_6170,N_5071,N_5159);
nand U6171 (N_6171,N_5291,N_4247);
nor U6172 (N_6172,N_5375,N_4884);
or U6173 (N_6173,N_5587,N_4163);
xnor U6174 (N_6174,N_5158,N_4695);
nor U6175 (N_6175,N_5592,N_5208);
nand U6176 (N_6176,N_4843,N_5899);
or U6177 (N_6177,N_5970,N_5319);
xor U6178 (N_6178,N_5669,N_5052);
nor U6179 (N_6179,N_4658,N_5976);
or U6180 (N_6180,N_4659,N_4099);
or U6181 (N_6181,N_4564,N_4437);
and U6182 (N_6182,N_4611,N_4138);
and U6183 (N_6183,N_5175,N_4974);
nand U6184 (N_6184,N_4068,N_5552);
and U6185 (N_6185,N_5042,N_4113);
nand U6186 (N_6186,N_4452,N_5524);
or U6187 (N_6187,N_5869,N_4172);
nor U6188 (N_6188,N_4535,N_4520);
nand U6189 (N_6189,N_4250,N_4666);
or U6190 (N_6190,N_5736,N_5336);
and U6191 (N_6191,N_4559,N_4142);
nand U6192 (N_6192,N_4821,N_5293);
or U6193 (N_6193,N_4548,N_5694);
and U6194 (N_6194,N_5439,N_4093);
and U6195 (N_6195,N_4075,N_5681);
nor U6196 (N_6196,N_4481,N_4420);
nand U6197 (N_6197,N_4642,N_5577);
and U6198 (N_6198,N_4354,N_4646);
or U6199 (N_6199,N_5838,N_4365);
xnor U6200 (N_6200,N_5972,N_4087);
xor U6201 (N_6201,N_5004,N_5546);
or U6202 (N_6202,N_5187,N_5009);
nor U6203 (N_6203,N_4196,N_5358);
or U6204 (N_6204,N_5672,N_4015);
xor U6205 (N_6205,N_5797,N_4858);
xor U6206 (N_6206,N_4985,N_4032);
and U6207 (N_6207,N_5800,N_4832);
nor U6208 (N_6208,N_5364,N_4756);
nor U6209 (N_6209,N_4103,N_4298);
and U6210 (N_6210,N_4370,N_5533);
xor U6211 (N_6211,N_5824,N_5792);
nor U6212 (N_6212,N_4781,N_5361);
and U6213 (N_6213,N_5422,N_4894);
and U6214 (N_6214,N_4597,N_4731);
nand U6215 (N_6215,N_4288,N_4936);
nor U6216 (N_6216,N_5934,N_4467);
nor U6217 (N_6217,N_5513,N_4297);
nand U6218 (N_6218,N_5138,N_5908);
nand U6219 (N_6219,N_5691,N_4230);
nand U6220 (N_6220,N_5407,N_4182);
and U6221 (N_6221,N_4765,N_5594);
nand U6222 (N_6222,N_5440,N_5904);
or U6223 (N_6223,N_5937,N_5820);
nand U6224 (N_6224,N_5001,N_4186);
nand U6225 (N_6225,N_4720,N_4468);
nand U6226 (N_6226,N_5043,N_5270);
and U6227 (N_6227,N_4673,N_4792);
xnor U6228 (N_6228,N_5362,N_5352);
nor U6229 (N_6229,N_4704,N_4194);
xnor U6230 (N_6230,N_5710,N_5854);
and U6231 (N_6231,N_4510,N_5015);
nor U6232 (N_6232,N_4844,N_5804);
xnor U6233 (N_6233,N_5223,N_4466);
or U6234 (N_6234,N_4139,N_4159);
xor U6235 (N_6235,N_5944,N_5234);
nand U6236 (N_6236,N_5853,N_5627);
and U6237 (N_6237,N_5017,N_4151);
nand U6238 (N_6238,N_4960,N_5894);
xnor U6239 (N_6239,N_5927,N_5896);
xnor U6240 (N_6240,N_5054,N_5036);
nand U6241 (N_6241,N_5402,N_4373);
nor U6242 (N_6242,N_4275,N_5534);
or U6243 (N_6243,N_4024,N_4101);
nor U6244 (N_6244,N_4668,N_5692);
nand U6245 (N_6245,N_4639,N_5721);
xnor U6246 (N_6246,N_5092,N_4008);
nand U6247 (N_6247,N_4184,N_4706);
xor U6248 (N_6248,N_4699,N_4958);
or U6249 (N_6249,N_4067,N_4060);
nand U6250 (N_6250,N_5194,N_5039);
xnor U6251 (N_6251,N_4381,N_5117);
or U6252 (N_6252,N_4942,N_4684);
nor U6253 (N_6253,N_5288,N_4460);
nor U6254 (N_6254,N_5105,N_5553);
and U6255 (N_6255,N_4545,N_5664);
and U6256 (N_6256,N_4835,N_4148);
nor U6257 (N_6257,N_4485,N_4806);
and U6258 (N_6258,N_5161,N_5708);
nand U6259 (N_6259,N_4712,N_5427);
xnor U6260 (N_6260,N_5661,N_4216);
xnor U6261 (N_6261,N_4011,N_4871);
or U6262 (N_6262,N_4681,N_4206);
or U6263 (N_6263,N_4610,N_4574);
or U6264 (N_6264,N_4457,N_4054);
xnor U6265 (N_6265,N_5559,N_5990);
xnor U6266 (N_6266,N_5408,N_4780);
nor U6267 (N_6267,N_5119,N_5858);
xor U6268 (N_6268,N_4604,N_4766);
and U6269 (N_6269,N_4560,N_5597);
nor U6270 (N_6270,N_4192,N_4989);
nor U6271 (N_6271,N_5828,N_4939);
nor U6272 (N_6272,N_4896,N_4952);
and U6273 (N_6273,N_5500,N_5846);
nand U6274 (N_6274,N_4006,N_5076);
nand U6275 (N_6275,N_4033,N_5272);
or U6276 (N_6276,N_4189,N_4910);
and U6277 (N_6277,N_5566,N_4476);
nand U6278 (N_6278,N_4294,N_5712);
or U6279 (N_6279,N_4080,N_4144);
or U6280 (N_6280,N_4546,N_4721);
or U6281 (N_6281,N_4329,N_5867);
nor U6282 (N_6282,N_4431,N_5134);
nor U6283 (N_6283,N_4750,N_5508);
or U6284 (N_6284,N_5723,N_5998);
nor U6285 (N_6285,N_4497,N_5608);
nand U6286 (N_6286,N_4870,N_4330);
and U6287 (N_6287,N_4393,N_4051);
xnor U6288 (N_6288,N_5574,N_4912);
or U6289 (N_6289,N_5634,N_4453);
and U6290 (N_6290,N_4524,N_4682);
xor U6291 (N_6291,N_4777,N_4676);
nand U6292 (N_6292,N_5522,N_4059);
nand U6293 (N_6293,N_4590,N_5675);
or U6294 (N_6294,N_4040,N_5844);
nand U6295 (N_6295,N_5888,N_5430);
or U6296 (N_6296,N_4293,N_5751);
nor U6297 (N_6297,N_5295,N_5626);
and U6298 (N_6298,N_5219,N_5863);
and U6299 (N_6299,N_4083,N_4776);
nand U6300 (N_6300,N_5492,N_5808);
xor U6301 (N_6301,N_4095,N_4899);
nor U6302 (N_6302,N_5224,N_5228);
nand U6303 (N_6303,N_5435,N_5767);
nand U6304 (N_6304,N_4309,N_5371);
nor U6305 (N_6305,N_5928,N_4323);
nor U6306 (N_6306,N_5884,N_4369);
or U6307 (N_6307,N_5699,N_4598);
and U6308 (N_6308,N_4881,N_5921);
or U6309 (N_6309,N_5676,N_5097);
nand U6310 (N_6310,N_4494,N_5603);
nand U6311 (N_6311,N_4579,N_5424);
nor U6312 (N_6312,N_5220,N_5069);
nor U6313 (N_6313,N_4403,N_5247);
nor U6314 (N_6314,N_5628,N_5501);
xnor U6315 (N_6315,N_4758,N_4328);
and U6316 (N_6316,N_5419,N_5891);
or U6317 (N_6317,N_5523,N_5110);
nand U6318 (N_6318,N_4164,N_4947);
nor U6319 (N_6319,N_5835,N_4097);
nor U6320 (N_6320,N_5585,N_5135);
and U6321 (N_6321,N_4585,N_4605);
xnor U6322 (N_6322,N_4783,N_5674);
nor U6323 (N_6323,N_5713,N_4500);
or U6324 (N_6324,N_5923,N_4417);
nand U6325 (N_6325,N_4173,N_4617);
xor U6326 (N_6326,N_5539,N_5570);
and U6327 (N_6327,N_5469,N_5515);
nand U6328 (N_6328,N_4359,N_5686);
xnor U6329 (N_6329,N_5707,N_5996);
nand U6330 (N_6330,N_4308,N_4857);
and U6331 (N_6331,N_5330,N_5504);
nand U6332 (N_6332,N_5906,N_4715);
nor U6333 (N_6333,N_5130,N_5662);
xor U6334 (N_6334,N_5133,N_5048);
or U6335 (N_6335,N_4810,N_5431);
and U6336 (N_6336,N_5768,N_5581);
xnor U6337 (N_6337,N_5637,N_5243);
nor U6338 (N_6338,N_5394,N_5816);
xor U6339 (N_6339,N_5517,N_5068);
nor U6340 (N_6340,N_4745,N_5008);
and U6341 (N_6341,N_5892,N_4925);
or U6342 (N_6342,N_4921,N_4943);
or U6343 (N_6343,N_5116,N_5070);
nor U6344 (N_6344,N_4406,N_5266);
nand U6345 (N_6345,N_4711,N_5289);
or U6346 (N_6346,N_5438,N_5734);
and U6347 (N_6347,N_4325,N_5889);
nand U6348 (N_6348,N_5755,N_4326);
nand U6349 (N_6349,N_4038,N_5512);
nand U6350 (N_6350,N_5236,N_5225);
and U6351 (N_6351,N_4558,N_5482);
xor U6352 (N_6352,N_4043,N_5757);
nor U6353 (N_6353,N_5956,N_4512);
and U6354 (N_6354,N_5605,N_5591);
and U6355 (N_6355,N_4770,N_5218);
or U6356 (N_6356,N_4069,N_4447);
nor U6357 (N_6357,N_4241,N_5329);
nand U6358 (N_6358,N_5311,N_5560);
nor U6359 (N_6359,N_5831,N_5421);
and U6360 (N_6360,N_5237,N_5322);
nor U6361 (N_6361,N_4158,N_4933);
and U6362 (N_6362,N_4459,N_5502);
xor U6363 (N_6363,N_5761,N_5871);
and U6364 (N_6364,N_4296,N_5342);
and U6365 (N_6365,N_5355,N_4175);
xnor U6366 (N_6366,N_5543,N_4553);
xnor U6367 (N_6367,N_4168,N_5108);
or U6368 (N_6368,N_4320,N_5683);
nand U6369 (N_6369,N_4850,N_5687);
and U6370 (N_6370,N_4656,N_5055);
nand U6371 (N_6371,N_4623,N_4999);
or U6372 (N_6372,N_4193,N_4228);
or U6373 (N_6373,N_5629,N_4732);
and U6374 (N_6374,N_5379,N_5498);
xnor U6375 (N_6375,N_5992,N_5007);
nand U6376 (N_6376,N_5870,N_5657);
nand U6377 (N_6377,N_4782,N_4048);
or U6378 (N_6378,N_5284,N_4027);
xnor U6379 (N_6379,N_4908,N_5813);
or U6380 (N_6380,N_5829,N_4707);
nand U6381 (N_6381,N_5016,N_4790);
and U6382 (N_6382,N_4848,N_4115);
or U6383 (N_6383,N_5769,N_4321);
and U6384 (N_6384,N_5621,N_5171);
nor U6385 (N_6385,N_5510,N_4143);
and U6386 (N_6386,N_5302,N_4152);
xor U6387 (N_6387,N_4726,N_4803);
nor U6388 (N_6388,N_5112,N_5320);
and U6389 (N_6389,N_4176,N_5143);
nand U6390 (N_6390,N_5264,N_4478);
xnor U6391 (N_6391,N_5984,N_4491);
or U6392 (N_6392,N_4091,N_5256);
xor U6393 (N_6393,N_4313,N_4318);
or U6394 (N_6394,N_4669,N_5101);
and U6395 (N_6395,N_5620,N_4191);
xnor U6396 (N_6396,N_4234,N_5102);
xnor U6397 (N_6397,N_5811,N_4096);
nor U6398 (N_6398,N_5113,N_5477);
nor U6399 (N_6399,N_4253,N_5308);
or U6400 (N_6400,N_4519,N_5511);
nor U6401 (N_6401,N_4347,N_4433);
xnor U6402 (N_6402,N_5207,N_5814);
and U6403 (N_6403,N_5933,N_5061);
xnor U6404 (N_6404,N_4331,N_5981);
and U6405 (N_6405,N_5339,N_4123);
nor U6406 (N_6406,N_5483,N_4675);
xor U6407 (N_6407,N_4317,N_5643);
and U6408 (N_6408,N_5689,N_4809);
and U6409 (N_6409,N_5192,N_5677);
nand U6410 (N_6410,N_4995,N_5663);
nor U6411 (N_6411,N_5668,N_5918);
xor U6412 (N_6412,N_5514,N_4525);
or U6413 (N_6413,N_4131,N_4411);
or U6414 (N_6414,N_5050,N_5850);
or U6415 (N_6415,N_4227,N_5727);
xnor U6416 (N_6416,N_4735,N_4377);
and U6417 (N_6417,N_5146,N_5617);
nor U6418 (N_6418,N_4938,N_5741);
nor U6419 (N_6419,N_5750,N_5554);
or U6420 (N_6420,N_5084,N_5476);
and U6421 (N_6421,N_5943,N_4153);
nand U6422 (N_6422,N_5160,N_5732);
or U6423 (N_6423,N_4537,N_5005);
xnor U6424 (N_6424,N_4764,N_4607);
or U6425 (N_6425,N_5540,N_5666);
nor U6426 (N_6426,N_5091,N_5323);
xnor U6427 (N_6427,N_5114,N_4364);
or U6428 (N_6428,N_5575,N_4816);
or U6429 (N_6429,N_4931,N_4618);
and U6430 (N_6430,N_4825,N_5456);
or U6431 (N_6431,N_5126,N_5772);
nor U6432 (N_6432,N_5080,N_4252);
xnor U6433 (N_6433,N_4730,N_5821);
nor U6434 (N_6434,N_5759,N_5156);
xor U6435 (N_6435,N_4967,N_4584);
nand U6436 (N_6436,N_5693,N_5584);
xnor U6437 (N_6437,N_5589,N_4508);
and U6438 (N_6438,N_5936,N_4878);
or U6439 (N_6439,N_4982,N_4368);
or U6440 (N_6440,N_4670,N_4290);
or U6441 (N_6441,N_5938,N_5979);
xor U6442 (N_6442,N_5258,N_4859);
nor U6443 (N_6443,N_5305,N_4395);
or U6444 (N_6444,N_5204,N_4344);
and U6445 (N_6445,N_4049,N_4755);
and U6446 (N_6446,N_4541,N_4786);
nand U6447 (N_6447,N_4641,N_5382);
xor U6448 (N_6448,N_4409,N_5487);
xor U6449 (N_6449,N_5499,N_4053);
nand U6450 (N_6450,N_4955,N_4672);
xor U6451 (N_6451,N_5941,N_4213);
nor U6452 (N_6452,N_5432,N_4934);
nand U6453 (N_6453,N_4852,N_5077);
or U6454 (N_6454,N_4086,N_5011);
or U6455 (N_6455,N_4877,N_5709);
nor U6456 (N_6456,N_5880,N_4162);
nand U6457 (N_6457,N_4917,N_4451);
and U6458 (N_6458,N_4301,N_4544);
nand U6459 (N_6459,N_4271,N_5095);
nand U6460 (N_6460,N_4802,N_5047);
nand U6461 (N_6461,N_5877,N_4577);
or U6462 (N_6462,N_4092,N_4319);
and U6463 (N_6463,N_5383,N_4282);
and U6464 (N_6464,N_5785,N_4495);
nand U6465 (N_6465,N_5935,N_4349);
nand U6466 (N_6466,N_4400,N_4900);
nor U6467 (N_6467,N_5484,N_4311);
or U6468 (N_6468,N_5072,N_5527);
nand U6469 (N_6469,N_5655,N_4076);
nor U6470 (N_6470,N_5836,N_4490);
xnor U6471 (N_6471,N_4117,N_5451);
nand U6472 (N_6472,N_4304,N_5787);
xnor U6473 (N_6473,N_4041,N_5648);
xnor U6474 (N_6474,N_5259,N_4346);
nor U6475 (N_6475,N_4880,N_5129);
xor U6476 (N_6476,N_5746,N_5473);
and U6477 (N_6477,N_4450,N_5044);
nand U6478 (N_6478,N_5078,N_4487);
nor U6479 (N_6479,N_4445,N_5519);
xor U6480 (N_6480,N_5604,N_4352);
xnor U6481 (N_6481,N_4621,N_4898);
nand U6482 (N_6482,N_5485,N_5849);
or U6483 (N_6483,N_4987,N_5611);
and U6484 (N_6484,N_5144,N_4366);
nor U6485 (N_6485,N_4090,N_4338);
or U6486 (N_6486,N_4029,N_5444);
nand U6487 (N_6487,N_4595,N_4554);
nor U6488 (N_6488,N_4020,N_4640);
nor U6489 (N_6489,N_4444,N_5961);
nand U6490 (N_6490,N_5959,N_5298);
or U6491 (N_6491,N_5195,N_4842);
and U6492 (N_6492,N_4787,N_4563);
and U6493 (N_6493,N_5962,N_5359);
xnor U6494 (N_6494,N_5745,N_4963);
or U6495 (N_6495,N_5098,N_4654);
and U6496 (N_6496,N_4208,N_5185);
xor U6497 (N_6497,N_4507,N_4807);
nor U6498 (N_6498,N_5388,N_4440);
xor U6499 (N_6499,N_4769,N_4469);
or U6500 (N_6500,N_5345,N_5788);
or U6501 (N_6501,N_5999,N_5653);
xor U6502 (N_6502,N_5883,N_4567);
nor U6503 (N_6503,N_4788,N_4998);
and U6504 (N_6504,N_5609,N_5315);
nor U6505 (N_6505,N_5914,N_5249);
nor U6506 (N_6506,N_5380,N_5317);
xor U6507 (N_6507,N_5267,N_5468);
nand U6508 (N_6508,N_4345,N_5725);
nor U6509 (N_6509,N_4923,N_4566);
nand U6510 (N_6510,N_4833,N_5494);
nand U6511 (N_6511,N_5847,N_5839);
nand U6512 (N_6512,N_5988,N_4341);
nand U6513 (N_6513,N_4978,N_5947);
nand U6514 (N_6514,N_5716,N_5425);
nand U6515 (N_6515,N_4853,N_5924);
and U6516 (N_6516,N_4948,N_4118);
xnor U6517 (N_6517,N_5436,N_4935);
or U6518 (N_6518,N_5565,N_4596);
or U6519 (N_6519,N_5569,N_5028);
xor U6520 (N_6520,N_5109,N_4285);
nor U6521 (N_6521,N_4685,N_4233);
or U6522 (N_6522,N_4866,N_4315);
or U6523 (N_6523,N_4789,N_5252);
nand U6524 (N_6524,N_5275,N_5154);
xnor U6525 (N_6525,N_4828,N_5263);
and U6526 (N_6526,N_4578,N_4300);
and U6527 (N_6527,N_4797,N_5333);
xor U6528 (N_6528,N_5087,N_4624);
or U6529 (N_6529,N_4742,N_4218);
and U6530 (N_6530,N_4547,N_4223);
nand U6531 (N_6531,N_4556,N_5434);
and U6532 (N_6532,N_4734,N_5437);
xnor U6533 (N_6533,N_5262,N_4518);
nand U6534 (N_6534,N_4697,N_4187);
or U6535 (N_6535,N_4343,N_5590);
or U6536 (N_6536,N_4757,N_5994);
nand U6537 (N_6537,N_5276,N_4157);
and U6538 (N_6538,N_5268,N_4889);
xnor U6539 (N_6539,N_4517,N_5879);
and U6540 (N_6540,N_4503,N_5312);
nor U6541 (N_6541,N_4523,N_5616);
nand U6542 (N_6542,N_5958,N_5749);
xnor U6543 (N_6543,N_4608,N_4471);
and U6544 (N_6544,N_4107,N_4972);
nand U6545 (N_6545,N_5917,N_5913);
xnor U6546 (N_6546,N_5774,N_5595);
nand U6547 (N_6547,N_5702,N_5612);
nor U6548 (N_6548,N_5572,N_4089);
and U6549 (N_6549,N_5082,N_5909);
xor U6550 (N_6550,N_4005,N_4965);
nand U6551 (N_6551,N_4586,N_4988);
and U6552 (N_6552,N_5488,N_4484);
or U6553 (N_6553,N_4583,N_5815);
nor U6554 (N_6554,N_5640,N_4968);
xor U6555 (N_6555,N_5152,N_4800);
nor U6556 (N_6556,N_5541,N_5202);
and U6557 (N_6557,N_5697,N_5805);
nor U6558 (N_6558,N_5401,N_5309);
or U6559 (N_6559,N_5931,N_5465);
nand U6560 (N_6560,N_5328,N_4573);
nor U6561 (N_6561,N_4378,N_4615);
nor U6562 (N_6562,N_5770,N_4645);
nor U6563 (N_6563,N_5400,N_4845);
or U6564 (N_6564,N_5341,N_4950);
xor U6565 (N_6565,N_5776,N_4180);
xnor U6566 (N_6566,N_5679,N_5809);
and U6567 (N_6567,N_5507,N_4798);
nand U6568 (N_6568,N_5942,N_5297);
nand U6569 (N_6569,N_4239,N_5782);
nand U6570 (N_6570,N_5997,N_4310);
and U6571 (N_6571,N_5193,N_4826);
and U6572 (N_6572,N_5503,N_4128);
nor U6573 (N_6573,N_4827,N_5396);
nor U6574 (N_6574,N_5030,N_4255);
nand U6575 (N_6575,N_4477,N_4470);
or U6576 (N_6576,N_4886,N_5012);
nand U6577 (N_6577,N_4019,N_4238);
nand U6578 (N_6578,N_4287,N_5093);
xor U6579 (N_6579,N_4472,N_4166);
or U6580 (N_6580,N_4932,N_5251);
nor U6581 (N_6581,N_4570,N_4661);
nand U6582 (N_6582,N_4791,N_4174);
nand U6583 (N_6583,N_5409,N_5075);
xnor U6584 (N_6584,N_5794,N_4276);
or U6585 (N_6585,N_5373,N_5586);
nand U6586 (N_6586,N_4012,N_4132);
and U6587 (N_6587,N_4299,N_5658);
nand U6588 (N_6588,N_5157,N_5180);
xor U6589 (N_6589,N_4201,N_4256);
or U6590 (N_6590,N_4538,N_4065);
and U6591 (N_6591,N_5722,N_5285);
and U6592 (N_6592,N_5717,N_4651);
nand U6593 (N_6593,N_4767,N_4116);
or U6594 (N_6594,N_5593,N_5832);
nand U6595 (N_6595,N_5378,N_4242);
or U6596 (N_6596,N_5125,N_5269);
nand U6597 (N_6597,N_5530,N_4696);
nand U6598 (N_6598,N_4716,N_5060);
and U6599 (N_6599,N_4634,N_5922);
and U6600 (N_6600,N_5881,N_5051);
and U6601 (N_6601,N_5292,N_5023);
nand U6602 (N_6602,N_5176,N_5861);
xnor U6603 (N_6603,N_5395,N_5963);
nor U6604 (N_6604,N_5418,N_4084);
or U6605 (N_6605,N_4951,N_5211);
nor U6606 (N_6606,N_5542,N_5939);
and U6607 (N_6607,N_5910,N_5280);
nand U6608 (N_6608,N_5520,N_5410);
nor U6609 (N_6609,N_4779,N_4057);
nor U6610 (N_6610,N_4161,N_5974);
xor U6611 (N_6611,N_5715,N_5376);
and U6612 (N_6612,N_5742,N_5557);
or U6613 (N_6613,N_5830,N_4203);
nor U6614 (N_6614,N_5987,N_4818);
nand U6615 (N_6615,N_4528,N_4571);
and U6616 (N_6616,N_4124,N_5167);
and U6617 (N_6617,N_5325,N_4837);
nand U6618 (N_6618,N_4070,N_5659);
or U6619 (N_6619,N_4202,N_5196);
nor U6620 (N_6620,N_5413,N_5448);
and U6621 (N_6621,N_5929,N_4295);
or U6622 (N_6622,N_4062,N_4550);
nor U6623 (N_6623,N_4045,N_4081);
and U6624 (N_6624,N_4350,N_5562);
or U6625 (N_6625,N_5442,N_4748);
nor U6626 (N_6626,N_4879,N_5706);
and U6627 (N_6627,N_4272,N_4527);
xor U6628 (N_6628,N_4593,N_5551);
and U6629 (N_6629,N_4100,N_5756);
nor U6630 (N_6630,N_5128,N_4273);
and U6631 (N_6631,N_4004,N_4199);
and U6632 (N_6632,N_4195,N_5155);
or U6633 (N_6633,N_4121,N_5426);
nand U6634 (N_6634,N_5529,N_4773);
or U6635 (N_6635,N_4264,N_5841);
or U6636 (N_6636,N_4463,N_5973);
nor U6637 (N_6637,N_5902,N_5827);
xnor U6638 (N_6638,N_5231,N_5954);
xor U6639 (N_6639,N_5753,N_4372);
xnor U6640 (N_6640,N_4862,N_4875);
or U6641 (N_6641,N_5478,N_5010);
or U6642 (N_6642,N_4486,N_5766);
xnor U6643 (N_6643,N_4885,N_4514);
and U6644 (N_6644,N_5528,N_4627);
nor U6645 (N_6645,N_4479,N_4643);
and U6646 (N_6646,N_4109,N_5564);
or U6647 (N_6647,N_5186,N_4867);
nand U6648 (N_6648,N_4398,N_4815);
nor U6649 (N_6649,N_5147,N_5807);
or U6650 (N_6650,N_4515,N_5610);
or U6651 (N_6651,N_4217,N_5067);
nand U6652 (N_6652,N_5622,N_4221);
xnor U6653 (N_6653,N_4055,N_5235);
nand U6654 (N_6654,N_5645,N_4506);
and U6655 (N_6655,N_4839,N_4680);
and U6656 (N_6656,N_4511,N_4994);
or U6657 (N_6657,N_4976,N_5027);
nor U6658 (N_6658,N_5452,N_5462);
xor U6659 (N_6659,N_5728,N_5536);
nand U6660 (N_6660,N_4375,N_4407);
xor U6661 (N_6661,N_5654,N_5678);
nor U6662 (N_6662,N_4246,N_5550);
nand U6663 (N_6663,N_4419,N_5053);
nand U6664 (N_6664,N_4448,N_5719);
nand U6665 (N_6665,N_5040,N_4534);
nor U6666 (N_6666,N_4855,N_4714);
or U6667 (N_6667,N_4718,N_5045);
nand U6668 (N_6668,N_4973,N_4283);
nor U6669 (N_6669,N_5738,N_4502);
xnor U6670 (N_6670,N_5642,N_4970);
xor U6671 (N_6671,N_5472,N_4088);
or U6672 (N_6672,N_5688,N_5120);
nand U6673 (N_6673,N_5470,N_4945);
and U6674 (N_6674,N_4028,N_4749);
nor U6675 (N_6675,N_5711,N_5895);
nor U6676 (N_6676,N_4723,N_4423);
and U6677 (N_6677,N_5169,N_5455);
xnor U6678 (N_6678,N_4361,N_4188);
nor U6679 (N_6679,N_5837,N_5141);
xor U6680 (N_6680,N_4979,N_4997);
and U6681 (N_6681,N_4606,N_5793);
or U6682 (N_6682,N_4268,N_4137);
nand U6683 (N_6683,N_5115,N_4928);
or U6684 (N_6684,N_4037,N_4122);
or U6685 (N_6685,N_4930,N_4170);
and U6686 (N_6686,N_5214,N_4532);
and U6687 (N_6687,N_5652,N_5340);
nand U6688 (N_6688,N_4941,N_4430);
xnor U6689 (N_6689,N_4397,N_5558);
or U6690 (N_6690,N_4863,N_5980);
nor U6691 (N_6691,N_4171,N_5480);
nor U6692 (N_6692,N_4284,N_4768);
and U6693 (N_6693,N_4760,N_4278);
xor U6694 (N_6694,N_4820,N_5802);
nor U6695 (N_6695,N_5104,N_5090);
and U6696 (N_6696,N_4992,N_4244);
xor U6697 (N_6697,N_4222,N_5203);
and U6698 (N_6698,N_5489,N_5094);
nor U6699 (N_6699,N_4418,N_4215);
xor U6700 (N_6700,N_5840,N_4263);
or U6701 (N_6701,N_4154,N_5791);
and U6702 (N_6702,N_4262,N_4984);
or U6703 (N_6703,N_5324,N_4530);
and U6704 (N_6704,N_5463,N_5474);
nor U6705 (N_6705,N_4582,N_5365);
nand U6706 (N_6706,N_4165,N_4160);
and U6707 (N_6707,N_4394,N_4784);
and U6708 (N_6708,N_5277,N_5786);
or U6709 (N_6709,N_4025,N_5764);
and U6710 (N_6710,N_5932,N_5760);
and U6711 (N_6711,N_4616,N_4499);
xor U6712 (N_6712,N_5213,N_4671);
nor U6713 (N_6713,N_5781,N_4663);
and U6714 (N_6714,N_4212,N_5952);
and U6715 (N_6715,N_5580,N_4426);
or U6716 (N_6716,N_4236,N_4861);
nor U6717 (N_6717,N_5148,N_5391);
or U6718 (N_6718,N_4156,N_5164);
or U6719 (N_6719,N_4733,N_4042);
nor U6720 (N_6720,N_5803,N_5253);
nor U6721 (N_6721,N_4353,N_5703);
and U6722 (N_6722,N_5795,N_4376);
and U6723 (N_6723,N_4897,N_5412);
nand U6724 (N_6724,N_5964,N_4599);
and U6725 (N_6725,N_5374,N_4824);
xnor U6726 (N_6726,N_4907,N_4488);
or U6727 (N_6727,N_4717,N_4647);
and U6728 (N_6728,N_5516,N_4581);
or U6729 (N_6729,N_5993,N_5454);
nand U6730 (N_6730,N_4834,N_4401);
or U6731 (N_6731,N_5014,N_4181);
nand U6732 (N_6732,N_5919,N_4371);
or U6733 (N_6733,N_5573,N_4983);
xnor U6734 (N_6734,N_4722,N_4281);
and U6735 (N_6735,N_4922,N_5545);
nor U6736 (N_6736,N_5471,N_5852);
xnor U6737 (N_6737,N_5222,N_4539);
nand U6738 (N_6738,N_4077,N_4626);
xor U6739 (N_6739,N_4455,N_5907);
and U6740 (N_6740,N_4386,N_5183);
nand U6741 (N_6741,N_4102,N_4094);
nor U6742 (N_6742,N_5046,N_4664);
nor U6743 (N_6743,N_5505,N_4868);
nor U6744 (N_6744,N_5967,N_4130);
xor U6745 (N_6745,N_4031,N_4286);
or U6746 (N_6746,N_5833,N_4705);
nor U6747 (N_6747,N_4438,N_5864);
and U6748 (N_6748,N_4316,N_4944);
nand U6749 (N_6749,N_4846,N_5357);
and U6750 (N_6750,N_4614,N_4763);
xnor U6751 (N_6751,N_5254,N_5518);
xor U6752 (N_6752,N_5957,N_5122);
nand U6753 (N_6753,N_5066,N_4693);
nor U6754 (N_6754,N_4903,N_5651);
nor U6755 (N_6755,N_4509,N_5614);
xor U6756 (N_6756,N_5977,N_4198);
nand U6757 (N_6757,N_4245,N_4047);
and U6758 (N_6758,N_5940,N_4110);
or U6759 (N_6759,N_4924,N_4129);
or U6760 (N_6760,N_5667,N_5796);
or U6761 (N_6761,N_5461,N_5083);
nand U6762 (N_6762,N_4106,N_5074);
and U6763 (N_6763,N_5568,N_4314);
or U6764 (N_6764,N_4876,N_4796);
xor U6765 (N_6765,N_5304,N_4249);
and U6766 (N_6766,N_5490,N_4277);
xnor U6767 (N_6767,N_5321,N_4357);
nand U6768 (N_6768,N_5765,N_4754);
or U6769 (N_6769,N_5377,N_5443);
and U6770 (N_6770,N_5021,N_4562);
nor U6771 (N_6771,N_4795,N_4362);
nand U6772 (N_6772,N_5107,N_5475);
and U6773 (N_6773,N_4888,N_5714);
or U6774 (N_6774,N_5025,N_4674);
xnor U6775 (N_6775,N_4587,N_5890);
xnor U6776 (N_6776,N_5636,N_4392);
xnor U6777 (N_6777,N_5411,N_5226);
nand U6778 (N_6778,N_5673,N_4906);
or U6779 (N_6779,N_5901,N_4105);
nand U6780 (N_6780,N_4736,N_5758);
xnor U6781 (N_6781,N_5690,N_4892);
xor U6782 (N_6782,N_5198,N_5834);
xor U6783 (N_6783,N_5926,N_4465);
and U6784 (N_6784,N_4588,N_5405);
or U6785 (N_6785,N_5897,N_4018);
and U6786 (N_6786,N_4751,N_5647);
nand U6787 (N_6787,N_4473,N_5985);
and U6788 (N_6788,N_4902,N_4568);
xor U6789 (N_6789,N_4251,N_5898);
or U6790 (N_6790,N_4402,N_5660);
nor U6791 (N_6791,N_5866,N_5777);
nor U6792 (N_6792,N_5212,N_4204);
nor U6793 (N_6793,N_5790,N_5851);
xor U6794 (N_6794,N_4211,N_4010);
nor U6795 (N_6795,N_4200,N_4630);
xor U6796 (N_6796,N_4637,N_4367);
and U6797 (N_6797,N_5618,N_5103);
xnor U6798 (N_6798,N_5088,N_5024);
nand U6799 (N_6799,N_4521,N_4056);
and U6800 (N_6800,N_5367,N_4046);
nand U6801 (N_6801,N_5331,N_5307);
nand U6802 (N_6802,N_4358,N_5506);
and U6803 (N_6803,N_5403,N_5783);
and U6804 (N_6804,N_5873,N_5294);
nor U6805 (N_6805,N_4214,N_5206);
nand U6806 (N_6806,N_5316,N_4185);
nor U6807 (N_6807,N_5497,N_4322);
xor U6808 (N_6808,N_4887,N_4261);
and U6809 (N_6809,N_5856,N_5695);
or U6810 (N_6810,N_5240,N_4458);
nor U6811 (N_6811,N_5780,N_4996);
nand U6812 (N_6812,N_4572,N_4687);
and U6813 (N_6813,N_4937,N_4000);
xor U6814 (N_6814,N_5433,N_5190);
or U6815 (N_6815,N_4741,N_5747);
and U6816 (N_6816,N_5602,N_4909);
xor U6817 (N_6817,N_4954,N_5644);
xnor U6818 (N_6818,N_5630,N_4072);
nor U6819 (N_6819,N_4543,N_4504);
nand U6820 (N_6820,N_4565,N_4169);
nand U6821 (N_6821,N_4078,N_5392);
nand U6822 (N_6822,N_4340,N_5313);
and U6823 (N_6823,N_5887,N_5623);
nor U6824 (N_6824,N_5995,N_5056);
nor U6825 (N_6825,N_4155,N_4785);
and U6826 (N_6826,N_4660,N_5227);
and U6827 (N_6827,N_4404,N_4482);
and U6828 (N_6828,N_4864,N_5168);
xnor U6829 (N_6829,N_5450,N_5819);
xnor U6830 (N_6830,N_4946,N_5386);
nand U6831 (N_6831,N_5613,N_5062);
nor U6832 (N_6832,N_5387,N_4980);
nand U6833 (N_6833,N_5911,N_4703);
xor U6834 (N_6834,N_4428,N_5464);
xor U6835 (N_6835,N_5701,N_4149);
xnor U6836 (N_6836,N_4324,N_5491);
and U6837 (N_6837,N_5370,N_5032);
and U6838 (N_6838,N_5086,N_5132);
nor U6839 (N_6839,N_5360,N_5242);
nor U6840 (N_6840,N_4146,N_5420);
nand U6841 (N_6841,N_5859,N_5241);
nand U6842 (N_6842,N_5458,N_5656);
nand U6843 (N_6843,N_5531,N_4501);
nor U6844 (N_6844,N_5548,N_4739);
or U6845 (N_6845,N_4135,N_4035);
nor U6846 (N_6846,N_4226,N_5041);
xnor U6847 (N_6847,N_5037,N_5822);
xnor U6848 (N_6848,N_5735,N_5983);
and U6849 (N_6849,N_4555,N_5754);
or U6850 (N_6850,N_5865,N_4529);
or U6851 (N_6851,N_4134,N_4071);
xnor U6852 (N_6852,N_5457,N_5799);
nor U6853 (N_6853,N_5638,N_5257);
nand U6854 (N_6854,N_4422,N_4991);
nor U6855 (N_6855,N_4197,N_5397);
xnor U6856 (N_6856,N_4224,N_4819);
xnor U6857 (N_6857,N_4432,N_5337);
and U6858 (N_6858,N_4126,N_4603);
or U6859 (N_6859,N_4291,N_5029);
and U6860 (N_6860,N_4462,N_5950);
and U6861 (N_6861,N_4964,N_5446);
nand U6862 (N_6862,N_5173,N_4688);
and U6863 (N_6863,N_5162,N_4243);
nor U6864 (N_6864,N_4044,N_4957);
or U6865 (N_6865,N_5124,N_4762);
nand U6866 (N_6866,N_5099,N_4829);
nand U6867 (N_6867,N_5743,N_5423);
nand U6868 (N_6868,N_4650,N_4890);
nand U6869 (N_6869,N_4926,N_4108);
and U6870 (N_6870,N_4380,N_5493);
nand U6871 (N_6871,N_5874,N_5778);
nand U6872 (N_6872,N_4355,N_5248);
xnor U6873 (N_6873,N_4822,N_5953);
or U6874 (N_6874,N_4235,N_4744);
or U6875 (N_6875,N_5459,N_4461);
xor U6876 (N_6876,N_5698,N_5338);
xnor U6877 (N_6877,N_5447,N_5079);
or U6878 (N_6878,N_4927,N_4231);
or U6879 (N_6879,N_4971,N_5567);
xnor U6880 (N_6880,N_5261,N_4334);
and U6881 (N_6881,N_4414,N_5779);
or U6882 (N_6882,N_4209,N_5271);
or U6883 (N_6883,N_5561,N_4891);
xor U6884 (N_6884,N_5429,N_4248);
nand U6885 (N_6885,N_4312,N_4405);
nand U6886 (N_6886,N_5230,N_5481);
or U6887 (N_6887,N_4389,N_5752);
and U6888 (N_6888,N_4034,N_4549);
nand U6889 (N_6889,N_4969,N_5003);
nor U6890 (N_6890,N_4949,N_5250);
and U6891 (N_6891,N_4454,N_4436);
or U6892 (N_6892,N_5600,N_5172);
or U6893 (N_6893,N_5299,N_4619);
and U6894 (N_6894,N_4427,N_5705);
nor U6895 (N_6895,N_4516,N_4775);
or U6896 (N_6896,N_5057,N_4052);
and U6897 (N_6897,N_5273,N_4649);
and U6898 (N_6898,N_4919,N_4531);
xnor U6899 (N_6899,N_4178,N_5350);
and U6900 (N_6900,N_5700,N_5038);
xnor U6901 (N_6901,N_5582,N_5290);
nor U6902 (N_6902,N_4966,N_4629);
nor U6903 (N_6903,N_5314,N_4975);
xor U6904 (N_6904,N_4391,N_4713);
or U6905 (N_6905,N_5260,N_5762);
and U6906 (N_6906,N_5073,N_5139);
and U6907 (N_6907,N_4442,N_4505);
nor U6908 (N_6908,N_4064,N_4893);
and U6909 (N_6909,N_4801,N_5878);
nor U6910 (N_6910,N_5930,N_5598);
or U6911 (N_6911,N_4120,N_5096);
nand U6912 (N_6912,N_4882,N_4449);
nand U6913 (N_6913,N_5385,N_5416);
or U6914 (N_6914,N_4575,N_4434);
or U6915 (N_6915,N_4793,N_5188);
or U6916 (N_6916,N_4023,N_5131);
nor U6917 (N_6917,N_5063,N_4002);
or U6918 (N_6918,N_5199,N_4632);
and U6919 (N_6919,N_5255,N_5825);
nand U6920 (N_6920,N_4594,N_5279);
nor U6921 (N_6921,N_5332,N_5818);
nor U6922 (N_6922,N_4805,N_5982);
or U6923 (N_6923,N_4986,N_5479);
and U6924 (N_6924,N_5449,N_4719);
or U6925 (N_6925,N_5229,N_4274);
or U6926 (N_6926,N_5986,N_4339);
nand U6927 (N_6927,N_5351,N_4424);
or U6928 (N_6928,N_4753,N_4962);
nor U6929 (N_6929,N_5165,N_4259);
nor U6930 (N_6930,N_4561,N_5384);
and U6931 (N_6931,N_4620,N_5968);
nor U6932 (N_6932,N_4533,N_4114);
xor U6933 (N_6933,N_5348,N_5238);
nor U6934 (N_6934,N_5393,N_5184);
nand U6935 (N_6935,N_5245,N_5453);
nor U6936 (N_6936,N_5525,N_4961);
xnor U6937 (N_6937,N_4003,N_5606);
nand U6938 (N_6938,N_5966,N_4677);
and U6939 (N_6939,N_4698,N_4177);
or U6940 (N_6940,N_4289,N_5763);
nor U6941 (N_6941,N_5823,N_4916);
or U6942 (N_6942,N_5696,N_5826);
nand U6943 (N_6943,N_5399,N_4761);
and U6944 (N_6944,N_4305,N_4702);
or U6945 (N_6945,N_5862,N_5232);
nor U6946 (N_6946,N_5163,N_4956);
nand U6947 (N_6947,N_4678,N_5670);
nor U6948 (N_6948,N_4303,N_5920);
xor U6949 (N_6949,N_4413,N_5978);
nand U6950 (N_6950,N_5650,N_5633);
nor U6951 (N_6951,N_5064,N_5000);
xor U6952 (N_6952,N_5031,N_4631);
and U6953 (N_6953,N_5089,N_4050);
and U6954 (N_6954,N_5615,N_5868);
xnor U6955 (N_6955,N_4492,N_5704);
or U6956 (N_6956,N_5282,N_5635);
nand U6957 (N_6957,N_4082,N_5353);
and U6958 (N_6958,N_5127,N_5296);
or U6959 (N_6959,N_4609,N_4270);
xor U6960 (N_6960,N_5576,N_4412);
and U6961 (N_6961,N_5170,N_4483);
nand U6962 (N_6962,N_4856,N_5265);
nor U6963 (N_6963,N_5335,N_4167);
nand U6964 (N_6964,N_4220,N_4342);
nand U6965 (N_6965,N_4613,N_5882);
nand U6966 (N_6966,N_4456,N_4602);
and U6967 (N_6967,N_5578,N_4014);
xnor U6968 (N_6968,N_5349,N_5197);
or U6969 (N_6969,N_5731,N_5631);
xor U6970 (N_6970,N_4812,N_4953);
nor U6971 (N_6971,N_4700,N_4136);
and U6972 (N_6972,N_5801,N_4911);
and U6973 (N_6973,N_5951,N_5538);
and U6974 (N_6974,N_4774,N_5151);
and U6975 (N_6975,N_4526,N_5381);
nor U6976 (N_6976,N_5789,N_5221);
xnor U6977 (N_6977,N_5354,N_4125);
xnor U6978 (N_6978,N_4280,N_4778);
and U6979 (N_6979,N_4759,N_5363);
or U6980 (N_6980,N_5390,N_4905);
nand U6981 (N_6981,N_5369,N_4628);
nor U6982 (N_6982,N_5945,N_4210);
nor U6983 (N_6983,N_5026,N_5179);
nand U6984 (N_6984,N_4638,N_4808);
or U6985 (N_6985,N_5366,N_4895);
nand U6986 (N_6986,N_4225,N_4799);
nor U6987 (N_6987,N_4265,N_5544);
nand U6988 (N_6988,N_4098,N_4552);
xor U6989 (N_6989,N_4522,N_4348);
or U6990 (N_6990,N_5415,N_5607);
xnor U6991 (N_6991,N_5684,N_4498);
nor U6992 (N_6992,N_5486,N_4416);
nor U6993 (N_6993,N_4747,N_4219);
and U6994 (N_6994,N_4269,N_5639);
and U6995 (N_6995,N_5916,N_5445);
nand U6996 (N_6996,N_5549,N_5532);
nor U6997 (N_6997,N_4662,N_4496);
nand U6998 (N_6998,N_4030,N_4036);
and U6999 (N_6999,N_5326,N_5646);
nor U7000 (N_7000,N_5908,N_5167);
nor U7001 (N_7001,N_4974,N_4328);
and U7002 (N_7002,N_5161,N_4939);
nor U7003 (N_7003,N_5820,N_5213);
nand U7004 (N_7004,N_4127,N_4971);
nor U7005 (N_7005,N_4371,N_4516);
nor U7006 (N_7006,N_5845,N_4379);
nand U7007 (N_7007,N_4541,N_5931);
nor U7008 (N_7008,N_4906,N_4134);
or U7009 (N_7009,N_5351,N_4244);
xor U7010 (N_7010,N_4671,N_4198);
nor U7011 (N_7011,N_5643,N_4694);
or U7012 (N_7012,N_4232,N_4270);
xor U7013 (N_7013,N_5055,N_4039);
nand U7014 (N_7014,N_4122,N_4905);
and U7015 (N_7015,N_4960,N_5693);
xor U7016 (N_7016,N_4157,N_5299);
nand U7017 (N_7017,N_4098,N_5084);
nand U7018 (N_7018,N_4385,N_5666);
or U7019 (N_7019,N_4665,N_5318);
xor U7020 (N_7020,N_4561,N_5761);
or U7021 (N_7021,N_4412,N_5827);
nor U7022 (N_7022,N_4039,N_4017);
nand U7023 (N_7023,N_4940,N_5969);
nor U7024 (N_7024,N_4449,N_5892);
xnor U7025 (N_7025,N_4653,N_4917);
or U7026 (N_7026,N_4019,N_4708);
and U7027 (N_7027,N_5131,N_5758);
and U7028 (N_7028,N_5923,N_4291);
and U7029 (N_7029,N_4017,N_5549);
or U7030 (N_7030,N_4621,N_5104);
or U7031 (N_7031,N_4403,N_5674);
xnor U7032 (N_7032,N_5303,N_4073);
xor U7033 (N_7033,N_5961,N_4275);
nor U7034 (N_7034,N_5778,N_4595);
nor U7035 (N_7035,N_4119,N_5497);
nor U7036 (N_7036,N_5345,N_4129);
or U7037 (N_7037,N_5777,N_4915);
nor U7038 (N_7038,N_4694,N_4434);
and U7039 (N_7039,N_5328,N_5113);
nand U7040 (N_7040,N_5368,N_4405);
or U7041 (N_7041,N_4836,N_4390);
nand U7042 (N_7042,N_4255,N_4060);
nor U7043 (N_7043,N_5193,N_4824);
or U7044 (N_7044,N_4561,N_4471);
and U7045 (N_7045,N_5662,N_5994);
nand U7046 (N_7046,N_4338,N_5813);
nand U7047 (N_7047,N_5621,N_4280);
and U7048 (N_7048,N_5497,N_4373);
nor U7049 (N_7049,N_5653,N_4067);
nor U7050 (N_7050,N_5654,N_5446);
and U7051 (N_7051,N_4839,N_4604);
xor U7052 (N_7052,N_5199,N_5266);
or U7053 (N_7053,N_4738,N_5787);
or U7054 (N_7054,N_4137,N_5742);
and U7055 (N_7055,N_5645,N_5163);
nand U7056 (N_7056,N_5006,N_4870);
or U7057 (N_7057,N_5612,N_4243);
nor U7058 (N_7058,N_4333,N_4328);
or U7059 (N_7059,N_5645,N_5046);
nor U7060 (N_7060,N_4863,N_5037);
or U7061 (N_7061,N_4997,N_4181);
nor U7062 (N_7062,N_4914,N_5773);
xor U7063 (N_7063,N_4426,N_5110);
or U7064 (N_7064,N_5549,N_4287);
nor U7065 (N_7065,N_5834,N_4925);
xnor U7066 (N_7066,N_4693,N_5032);
nand U7067 (N_7067,N_4259,N_4103);
nand U7068 (N_7068,N_4634,N_5470);
xor U7069 (N_7069,N_4681,N_5953);
or U7070 (N_7070,N_4354,N_5682);
or U7071 (N_7071,N_4602,N_5040);
nor U7072 (N_7072,N_5571,N_4418);
nor U7073 (N_7073,N_5566,N_5703);
and U7074 (N_7074,N_4049,N_4076);
or U7075 (N_7075,N_5948,N_4039);
xor U7076 (N_7076,N_4791,N_5885);
nor U7077 (N_7077,N_4723,N_4336);
nor U7078 (N_7078,N_5934,N_4387);
or U7079 (N_7079,N_4044,N_5089);
and U7080 (N_7080,N_4462,N_5171);
and U7081 (N_7081,N_4813,N_5732);
or U7082 (N_7082,N_5619,N_4161);
xnor U7083 (N_7083,N_4424,N_4706);
or U7084 (N_7084,N_4574,N_4115);
xnor U7085 (N_7085,N_4999,N_5522);
and U7086 (N_7086,N_5711,N_4401);
nand U7087 (N_7087,N_5341,N_4667);
and U7088 (N_7088,N_5396,N_5512);
and U7089 (N_7089,N_4543,N_4961);
xnor U7090 (N_7090,N_5508,N_5476);
nand U7091 (N_7091,N_5814,N_5526);
xnor U7092 (N_7092,N_5078,N_5351);
xnor U7093 (N_7093,N_5114,N_5687);
and U7094 (N_7094,N_5405,N_5264);
or U7095 (N_7095,N_4390,N_4492);
or U7096 (N_7096,N_5119,N_5787);
or U7097 (N_7097,N_4688,N_5883);
and U7098 (N_7098,N_5405,N_4712);
xnor U7099 (N_7099,N_5478,N_4937);
and U7100 (N_7100,N_5034,N_5965);
nand U7101 (N_7101,N_5665,N_5274);
xnor U7102 (N_7102,N_4239,N_5505);
nor U7103 (N_7103,N_5266,N_4395);
nor U7104 (N_7104,N_5558,N_5357);
and U7105 (N_7105,N_5858,N_4963);
nand U7106 (N_7106,N_5849,N_4217);
nand U7107 (N_7107,N_4613,N_4326);
xnor U7108 (N_7108,N_5782,N_5274);
and U7109 (N_7109,N_4084,N_5441);
nor U7110 (N_7110,N_5450,N_5451);
and U7111 (N_7111,N_4064,N_4440);
nor U7112 (N_7112,N_4037,N_4567);
and U7113 (N_7113,N_4983,N_5578);
nor U7114 (N_7114,N_4491,N_5232);
nor U7115 (N_7115,N_5327,N_5804);
nor U7116 (N_7116,N_4063,N_5956);
or U7117 (N_7117,N_5068,N_4082);
or U7118 (N_7118,N_4521,N_5826);
nor U7119 (N_7119,N_4154,N_4481);
and U7120 (N_7120,N_5611,N_5722);
nand U7121 (N_7121,N_5581,N_5771);
and U7122 (N_7122,N_4289,N_4941);
nand U7123 (N_7123,N_4534,N_4851);
and U7124 (N_7124,N_5863,N_5578);
and U7125 (N_7125,N_5558,N_5551);
or U7126 (N_7126,N_5107,N_4022);
xor U7127 (N_7127,N_4432,N_5530);
or U7128 (N_7128,N_5055,N_5110);
or U7129 (N_7129,N_5600,N_5696);
nand U7130 (N_7130,N_4135,N_5866);
and U7131 (N_7131,N_4791,N_4668);
xnor U7132 (N_7132,N_5083,N_4192);
and U7133 (N_7133,N_4408,N_5450);
and U7134 (N_7134,N_5591,N_4024);
xnor U7135 (N_7135,N_5949,N_4332);
or U7136 (N_7136,N_5715,N_4569);
nand U7137 (N_7137,N_5351,N_5838);
nor U7138 (N_7138,N_4631,N_4980);
and U7139 (N_7139,N_5733,N_5206);
xnor U7140 (N_7140,N_5484,N_5774);
or U7141 (N_7141,N_5159,N_5850);
or U7142 (N_7142,N_5923,N_5913);
xnor U7143 (N_7143,N_4168,N_4841);
and U7144 (N_7144,N_4720,N_4511);
nand U7145 (N_7145,N_5004,N_4218);
xnor U7146 (N_7146,N_4185,N_5060);
xor U7147 (N_7147,N_5758,N_5989);
and U7148 (N_7148,N_4202,N_4743);
and U7149 (N_7149,N_4497,N_5064);
and U7150 (N_7150,N_5282,N_5556);
or U7151 (N_7151,N_4808,N_4030);
or U7152 (N_7152,N_4993,N_4198);
and U7153 (N_7153,N_4570,N_5186);
and U7154 (N_7154,N_5532,N_5793);
xnor U7155 (N_7155,N_5278,N_5077);
or U7156 (N_7156,N_5061,N_4144);
xor U7157 (N_7157,N_5193,N_5128);
or U7158 (N_7158,N_5146,N_4799);
nand U7159 (N_7159,N_4816,N_4175);
xnor U7160 (N_7160,N_4757,N_5735);
and U7161 (N_7161,N_4705,N_4885);
nand U7162 (N_7162,N_5696,N_5114);
nor U7163 (N_7163,N_5342,N_4655);
xnor U7164 (N_7164,N_4497,N_4834);
nand U7165 (N_7165,N_5325,N_4433);
nand U7166 (N_7166,N_4048,N_4967);
xor U7167 (N_7167,N_5718,N_5448);
xnor U7168 (N_7168,N_5544,N_4084);
and U7169 (N_7169,N_4524,N_5121);
nand U7170 (N_7170,N_4909,N_5217);
or U7171 (N_7171,N_4205,N_5675);
or U7172 (N_7172,N_5861,N_5725);
or U7173 (N_7173,N_4828,N_4386);
or U7174 (N_7174,N_5805,N_4611);
nor U7175 (N_7175,N_5353,N_5165);
and U7176 (N_7176,N_5105,N_4264);
nor U7177 (N_7177,N_5689,N_4763);
nand U7178 (N_7178,N_5122,N_4641);
and U7179 (N_7179,N_5628,N_4397);
nor U7180 (N_7180,N_5345,N_5096);
nor U7181 (N_7181,N_4807,N_4603);
or U7182 (N_7182,N_4553,N_5746);
nor U7183 (N_7183,N_5603,N_5663);
nor U7184 (N_7184,N_4061,N_5417);
and U7185 (N_7185,N_5116,N_5030);
and U7186 (N_7186,N_5227,N_5905);
nor U7187 (N_7187,N_4176,N_4161);
and U7188 (N_7188,N_4907,N_4480);
xor U7189 (N_7189,N_5289,N_4999);
and U7190 (N_7190,N_4917,N_5663);
xnor U7191 (N_7191,N_4575,N_5676);
xnor U7192 (N_7192,N_4196,N_4677);
nand U7193 (N_7193,N_5658,N_4793);
nor U7194 (N_7194,N_5457,N_5597);
or U7195 (N_7195,N_4915,N_5207);
nor U7196 (N_7196,N_5219,N_5655);
nand U7197 (N_7197,N_4458,N_4127);
nand U7198 (N_7198,N_5796,N_5351);
or U7199 (N_7199,N_5143,N_5824);
and U7200 (N_7200,N_5822,N_5036);
nand U7201 (N_7201,N_5260,N_4838);
nor U7202 (N_7202,N_4020,N_5115);
nor U7203 (N_7203,N_4470,N_4185);
nor U7204 (N_7204,N_4424,N_5240);
or U7205 (N_7205,N_4422,N_5403);
or U7206 (N_7206,N_4960,N_5646);
nor U7207 (N_7207,N_4188,N_5062);
nand U7208 (N_7208,N_5455,N_4943);
and U7209 (N_7209,N_5272,N_4483);
or U7210 (N_7210,N_4909,N_5697);
nand U7211 (N_7211,N_4387,N_4745);
nand U7212 (N_7212,N_5433,N_4683);
xnor U7213 (N_7213,N_4406,N_4921);
nand U7214 (N_7214,N_4115,N_5102);
nor U7215 (N_7215,N_5829,N_4411);
and U7216 (N_7216,N_5691,N_5854);
or U7217 (N_7217,N_5983,N_5812);
or U7218 (N_7218,N_4255,N_5750);
or U7219 (N_7219,N_4064,N_5458);
nor U7220 (N_7220,N_4459,N_5509);
nand U7221 (N_7221,N_4868,N_4810);
xnor U7222 (N_7222,N_4930,N_4497);
xnor U7223 (N_7223,N_5311,N_5714);
nor U7224 (N_7224,N_4248,N_5235);
xor U7225 (N_7225,N_5164,N_5215);
and U7226 (N_7226,N_4113,N_4323);
and U7227 (N_7227,N_5191,N_4348);
and U7228 (N_7228,N_4450,N_5124);
xnor U7229 (N_7229,N_4615,N_4833);
nor U7230 (N_7230,N_5175,N_5432);
nand U7231 (N_7231,N_4589,N_4970);
and U7232 (N_7232,N_5589,N_4302);
nor U7233 (N_7233,N_5671,N_5686);
nor U7234 (N_7234,N_4521,N_5238);
xnor U7235 (N_7235,N_5128,N_5766);
nor U7236 (N_7236,N_4795,N_4155);
and U7237 (N_7237,N_4554,N_4153);
and U7238 (N_7238,N_4602,N_5071);
or U7239 (N_7239,N_4002,N_5332);
xor U7240 (N_7240,N_4925,N_5077);
and U7241 (N_7241,N_5876,N_4341);
nor U7242 (N_7242,N_4475,N_4286);
or U7243 (N_7243,N_4338,N_4164);
nand U7244 (N_7244,N_5478,N_4413);
nand U7245 (N_7245,N_4169,N_4807);
or U7246 (N_7246,N_5984,N_4428);
nand U7247 (N_7247,N_4537,N_4433);
xor U7248 (N_7248,N_5840,N_5544);
or U7249 (N_7249,N_5452,N_5702);
xor U7250 (N_7250,N_4912,N_5294);
nor U7251 (N_7251,N_5469,N_5254);
nand U7252 (N_7252,N_5782,N_5256);
nand U7253 (N_7253,N_4243,N_5911);
nand U7254 (N_7254,N_5946,N_5058);
or U7255 (N_7255,N_4611,N_4659);
nand U7256 (N_7256,N_5506,N_4126);
or U7257 (N_7257,N_5468,N_5769);
or U7258 (N_7258,N_4029,N_4586);
nand U7259 (N_7259,N_4980,N_4950);
or U7260 (N_7260,N_4768,N_4531);
xnor U7261 (N_7261,N_4487,N_5597);
or U7262 (N_7262,N_4982,N_4719);
nand U7263 (N_7263,N_5619,N_4833);
nor U7264 (N_7264,N_5715,N_4562);
and U7265 (N_7265,N_5341,N_4822);
nor U7266 (N_7266,N_4702,N_5714);
nand U7267 (N_7267,N_5167,N_4426);
nor U7268 (N_7268,N_4553,N_5347);
and U7269 (N_7269,N_5772,N_5978);
or U7270 (N_7270,N_5435,N_5444);
and U7271 (N_7271,N_5021,N_4367);
nor U7272 (N_7272,N_5577,N_4993);
nand U7273 (N_7273,N_5237,N_4392);
and U7274 (N_7274,N_4948,N_5183);
and U7275 (N_7275,N_5806,N_5727);
or U7276 (N_7276,N_5303,N_5418);
and U7277 (N_7277,N_5517,N_5700);
and U7278 (N_7278,N_5351,N_4050);
or U7279 (N_7279,N_4596,N_5109);
nor U7280 (N_7280,N_5581,N_5934);
and U7281 (N_7281,N_4490,N_5938);
xnor U7282 (N_7282,N_4641,N_5290);
nand U7283 (N_7283,N_4490,N_5780);
or U7284 (N_7284,N_5595,N_5042);
or U7285 (N_7285,N_5685,N_5454);
and U7286 (N_7286,N_4519,N_4265);
xor U7287 (N_7287,N_5485,N_5279);
nand U7288 (N_7288,N_5579,N_4384);
xnor U7289 (N_7289,N_5657,N_5767);
nand U7290 (N_7290,N_4492,N_5197);
xnor U7291 (N_7291,N_5735,N_4022);
xnor U7292 (N_7292,N_5567,N_5122);
and U7293 (N_7293,N_5415,N_5127);
nand U7294 (N_7294,N_5801,N_5214);
nand U7295 (N_7295,N_4054,N_4844);
and U7296 (N_7296,N_5590,N_4608);
xor U7297 (N_7297,N_5319,N_5603);
or U7298 (N_7298,N_5564,N_4338);
nand U7299 (N_7299,N_4816,N_5507);
xor U7300 (N_7300,N_4351,N_5227);
or U7301 (N_7301,N_5858,N_4856);
and U7302 (N_7302,N_5114,N_4919);
xnor U7303 (N_7303,N_5893,N_5955);
and U7304 (N_7304,N_5309,N_5481);
nand U7305 (N_7305,N_5360,N_5028);
nand U7306 (N_7306,N_5117,N_4402);
nor U7307 (N_7307,N_4643,N_4336);
nor U7308 (N_7308,N_4519,N_5896);
or U7309 (N_7309,N_5885,N_4873);
xor U7310 (N_7310,N_4198,N_4456);
xor U7311 (N_7311,N_5614,N_5041);
and U7312 (N_7312,N_4820,N_4807);
and U7313 (N_7313,N_5178,N_5699);
and U7314 (N_7314,N_5522,N_4900);
and U7315 (N_7315,N_4243,N_4658);
xor U7316 (N_7316,N_5833,N_4586);
nor U7317 (N_7317,N_4092,N_5597);
nand U7318 (N_7318,N_4683,N_4641);
nor U7319 (N_7319,N_4283,N_5097);
nand U7320 (N_7320,N_4415,N_5757);
and U7321 (N_7321,N_4649,N_5228);
and U7322 (N_7322,N_4370,N_5156);
and U7323 (N_7323,N_5391,N_5624);
or U7324 (N_7324,N_4767,N_4061);
nor U7325 (N_7325,N_5283,N_4295);
or U7326 (N_7326,N_4072,N_5676);
nor U7327 (N_7327,N_4498,N_4989);
or U7328 (N_7328,N_4273,N_4698);
or U7329 (N_7329,N_4441,N_4902);
and U7330 (N_7330,N_5592,N_5307);
nor U7331 (N_7331,N_4370,N_5041);
nor U7332 (N_7332,N_4910,N_5840);
nor U7333 (N_7333,N_4188,N_5837);
nor U7334 (N_7334,N_5241,N_4982);
nand U7335 (N_7335,N_4170,N_5056);
nand U7336 (N_7336,N_5686,N_5097);
or U7337 (N_7337,N_4793,N_5725);
xnor U7338 (N_7338,N_5958,N_4127);
nand U7339 (N_7339,N_5210,N_4142);
nor U7340 (N_7340,N_5620,N_4506);
xor U7341 (N_7341,N_5568,N_4218);
or U7342 (N_7342,N_4060,N_5016);
xor U7343 (N_7343,N_5678,N_5599);
or U7344 (N_7344,N_4193,N_4390);
and U7345 (N_7345,N_4127,N_5078);
nand U7346 (N_7346,N_4002,N_5689);
or U7347 (N_7347,N_5585,N_5565);
nor U7348 (N_7348,N_4669,N_5459);
or U7349 (N_7349,N_5082,N_5410);
nand U7350 (N_7350,N_4611,N_4418);
xnor U7351 (N_7351,N_5876,N_4945);
and U7352 (N_7352,N_5087,N_5406);
nor U7353 (N_7353,N_5227,N_4252);
xnor U7354 (N_7354,N_4749,N_5428);
or U7355 (N_7355,N_4613,N_5082);
nor U7356 (N_7356,N_4921,N_4470);
xor U7357 (N_7357,N_5212,N_5602);
or U7358 (N_7358,N_4343,N_4050);
xor U7359 (N_7359,N_4425,N_4595);
nand U7360 (N_7360,N_4586,N_4519);
and U7361 (N_7361,N_5900,N_5041);
and U7362 (N_7362,N_4698,N_4931);
or U7363 (N_7363,N_5902,N_5324);
nor U7364 (N_7364,N_4021,N_4507);
nor U7365 (N_7365,N_5510,N_5689);
nand U7366 (N_7366,N_5648,N_5619);
or U7367 (N_7367,N_4525,N_5664);
and U7368 (N_7368,N_5997,N_4570);
xor U7369 (N_7369,N_4747,N_4110);
or U7370 (N_7370,N_4148,N_4918);
nor U7371 (N_7371,N_4708,N_5885);
xnor U7372 (N_7372,N_5086,N_5986);
nand U7373 (N_7373,N_5205,N_4938);
xor U7374 (N_7374,N_5259,N_5908);
and U7375 (N_7375,N_5198,N_4115);
xor U7376 (N_7376,N_4895,N_5864);
nand U7377 (N_7377,N_5416,N_5563);
nand U7378 (N_7378,N_4506,N_4735);
nor U7379 (N_7379,N_5782,N_5593);
or U7380 (N_7380,N_4386,N_4937);
and U7381 (N_7381,N_5616,N_4604);
xnor U7382 (N_7382,N_5742,N_4892);
or U7383 (N_7383,N_5908,N_5540);
nor U7384 (N_7384,N_5004,N_5607);
nand U7385 (N_7385,N_5746,N_4944);
or U7386 (N_7386,N_4471,N_4789);
nand U7387 (N_7387,N_4594,N_5397);
nand U7388 (N_7388,N_4430,N_4531);
or U7389 (N_7389,N_5495,N_4753);
and U7390 (N_7390,N_5402,N_5026);
nor U7391 (N_7391,N_5185,N_5961);
and U7392 (N_7392,N_4985,N_5163);
or U7393 (N_7393,N_4441,N_4450);
xor U7394 (N_7394,N_4051,N_4754);
nor U7395 (N_7395,N_5756,N_5102);
nor U7396 (N_7396,N_4267,N_4102);
nor U7397 (N_7397,N_5719,N_5618);
nor U7398 (N_7398,N_5406,N_4077);
nand U7399 (N_7399,N_4240,N_4082);
or U7400 (N_7400,N_4562,N_5288);
xnor U7401 (N_7401,N_4020,N_4834);
xor U7402 (N_7402,N_5663,N_4708);
nand U7403 (N_7403,N_4760,N_5490);
nand U7404 (N_7404,N_5108,N_4248);
xor U7405 (N_7405,N_5666,N_4824);
and U7406 (N_7406,N_5294,N_4791);
xor U7407 (N_7407,N_4219,N_5700);
or U7408 (N_7408,N_4341,N_4679);
xnor U7409 (N_7409,N_4503,N_5958);
nand U7410 (N_7410,N_5420,N_5752);
nand U7411 (N_7411,N_4413,N_4372);
and U7412 (N_7412,N_4329,N_4415);
or U7413 (N_7413,N_5312,N_4339);
or U7414 (N_7414,N_4346,N_5396);
nand U7415 (N_7415,N_4385,N_4390);
xor U7416 (N_7416,N_5701,N_4554);
and U7417 (N_7417,N_4502,N_5623);
and U7418 (N_7418,N_5046,N_5700);
nor U7419 (N_7419,N_5475,N_4618);
and U7420 (N_7420,N_5870,N_4162);
or U7421 (N_7421,N_4768,N_4414);
nor U7422 (N_7422,N_5937,N_4109);
nor U7423 (N_7423,N_4999,N_4610);
xor U7424 (N_7424,N_5766,N_5856);
nor U7425 (N_7425,N_5156,N_4368);
or U7426 (N_7426,N_4066,N_5805);
nor U7427 (N_7427,N_5470,N_5273);
or U7428 (N_7428,N_4727,N_5831);
and U7429 (N_7429,N_5342,N_5234);
or U7430 (N_7430,N_4122,N_4882);
xnor U7431 (N_7431,N_5610,N_4448);
or U7432 (N_7432,N_4466,N_4153);
and U7433 (N_7433,N_5818,N_4600);
nand U7434 (N_7434,N_4241,N_5646);
or U7435 (N_7435,N_5896,N_5361);
and U7436 (N_7436,N_5525,N_5069);
nand U7437 (N_7437,N_4710,N_4416);
nor U7438 (N_7438,N_4717,N_5402);
and U7439 (N_7439,N_5839,N_4446);
xor U7440 (N_7440,N_4099,N_4230);
or U7441 (N_7441,N_4290,N_5099);
or U7442 (N_7442,N_5487,N_5628);
or U7443 (N_7443,N_4288,N_4736);
xor U7444 (N_7444,N_4075,N_4758);
xnor U7445 (N_7445,N_4758,N_5932);
nor U7446 (N_7446,N_5836,N_5125);
or U7447 (N_7447,N_5271,N_4507);
nor U7448 (N_7448,N_4843,N_5111);
nand U7449 (N_7449,N_4361,N_5135);
nor U7450 (N_7450,N_4391,N_4438);
or U7451 (N_7451,N_4528,N_5111);
nand U7452 (N_7452,N_5409,N_5129);
and U7453 (N_7453,N_5180,N_4351);
nor U7454 (N_7454,N_4772,N_4639);
xnor U7455 (N_7455,N_5754,N_5498);
and U7456 (N_7456,N_4044,N_4607);
nand U7457 (N_7457,N_5084,N_5015);
and U7458 (N_7458,N_4020,N_4259);
nor U7459 (N_7459,N_5008,N_5180);
and U7460 (N_7460,N_4770,N_5979);
nor U7461 (N_7461,N_4400,N_4032);
xor U7462 (N_7462,N_5150,N_4537);
nand U7463 (N_7463,N_5686,N_5533);
nand U7464 (N_7464,N_4406,N_4236);
nor U7465 (N_7465,N_4521,N_5764);
nor U7466 (N_7466,N_4428,N_5864);
xor U7467 (N_7467,N_5283,N_5098);
nor U7468 (N_7468,N_4286,N_4673);
nor U7469 (N_7469,N_5311,N_4414);
and U7470 (N_7470,N_4332,N_4800);
and U7471 (N_7471,N_5431,N_5142);
or U7472 (N_7472,N_4972,N_5547);
or U7473 (N_7473,N_5997,N_4726);
nand U7474 (N_7474,N_4322,N_4614);
or U7475 (N_7475,N_5084,N_5525);
xnor U7476 (N_7476,N_5295,N_5702);
nor U7477 (N_7477,N_4733,N_4981);
or U7478 (N_7478,N_4996,N_5269);
nor U7479 (N_7479,N_5897,N_4032);
xor U7480 (N_7480,N_4575,N_4763);
and U7481 (N_7481,N_5643,N_5345);
or U7482 (N_7482,N_5953,N_4253);
or U7483 (N_7483,N_5148,N_4209);
nor U7484 (N_7484,N_4491,N_5090);
xor U7485 (N_7485,N_5912,N_4926);
nand U7486 (N_7486,N_4581,N_4260);
nor U7487 (N_7487,N_4253,N_4317);
xnor U7488 (N_7488,N_5589,N_5840);
and U7489 (N_7489,N_5812,N_5318);
nor U7490 (N_7490,N_4115,N_4026);
or U7491 (N_7491,N_4726,N_5827);
or U7492 (N_7492,N_5202,N_5615);
nand U7493 (N_7493,N_5896,N_5990);
or U7494 (N_7494,N_5811,N_5850);
nand U7495 (N_7495,N_5313,N_5425);
nand U7496 (N_7496,N_5308,N_5737);
nand U7497 (N_7497,N_4117,N_5958);
or U7498 (N_7498,N_4630,N_5070);
nor U7499 (N_7499,N_4874,N_4281);
xnor U7500 (N_7500,N_5037,N_4372);
and U7501 (N_7501,N_4907,N_4375);
and U7502 (N_7502,N_5202,N_4840);
nor U7503 (N_7503,N_5077,N_5073);
or U7504 (N_7504,N_5346,N_5635);
or U7505 (N_7505,N_5035,N_4028);
xnor U7506 (N_7506,N_4611,N_4585);
nor U7507 (N_7507,N_5960,N_4212);
and U7508 (N_7508,N_5297,N_4671);
or U7509 (N_7509,N_5853,N_5691);
nand U7510 (N_7510,N_4131,N_4554);
nor U7511 (N_7511,N_4593,N_5838);
xor U7512 (N_7512,N_4661,N_4810);
xor U7513 (N_7513,N_5340,N_5901);
or U7514 (N_7514,N_4295,N_4719);
nand U7515 (N_7515,N_4140,N_4858);
nand U7516 (N_7516,N_4599,N_4299);
nand U7517 (N_7517,N_4335,N_5591);
xnor U7518 (N_7518,N_5456,N_4743);
xnor U7519 (N_7519,N_4991,N_4327);
or U7520 (N_7520,N_4253,N_5561);
xnor U7521 (N_7521,N_4779,N_5456);
nand U7522 (N_7522,N_4249,N_4346);
nand U7523 (N_7523,N_5415,N_5998);
and U7524 (N_7524,N_5898,N_5705);
and U7525 (N_7525,N_5732,N_4617);
nand U7526 (N_7526,N_5491,N_4787);
and U7527 (N_7527,N_5956,N_4749);
nand U7528 (N_7528,N_4375,N_5779);
or U7529 (N_7529,N_5644,N_4273);
and U7530 (N_7530,N_4020,N_4589);
nand U7531 (N_7531,N_5139,N_4741);
nor U7532 (N_7532,N_4489,N_4567);
nand U7533 (N_7533,N_4798,N_4879);
and U7534 (N_7534,N_4216,N_4585);
xnor U7535 (N_7535,N_5120,N_4250);
and U7536 (N_7536,N_4916,N_5635);
nand U7537 (N_7537,N_5690,N_4645);
nor U7538 (N_7538,N_5984,N_4700);
and U7539 (N_7539,N_4994,N_5984);
xnor U7540 (N_7540,N_4541,N_4330);
xnor U7541 (N_7541,N_4067,N_5623);
nor U7542 (N_7542,N_4736,N_5992);
xnor U7543 (N_7543,N_4860,N_5412);
and U7544 (N_7544,N_4062,N_4597);
nor U7545 (N_7545,N_4070,N_5259);
and U7546 (N_7546,N_4538,N_5095);
nand U7547 (N_7547,N_4850,N_4654);
and U7548 (N_7548,N_4227,N_4268);
nor U7549 (N_7549,N_5282,N_5113);
and U7550 (N_7550,N_5641,N_4694);
or U7551 (N_7551,N_4834,N_4373);
or U7552 (N_7552,N_4747,N_4568);
nor U7553 (N_7553,N_5155,N_4206);
and U7554 (N_7554,N_4994,N_4605);
or U7555 (N_7555,N_4033,N_5989);
xor U7556 (N_7556,N_5391,N_5426);
nand U7557 (N_7557,N_5253,N_5370);
nand U7558 (N_7558,N_5039,N_5164);
nor U7559 (N_7559,N_4570,N_4643);
nor U7560 (N_7560,N_5329,N_5611);
nor U7561 (N_7561,N_5979,N_4402);
xnor U7562 (N_7562,N_5175,N_4117);
nor U7563 (N_7563,N_5070,N_4972);
or U7564 (N_7564,N_5921,N_4211);
and U7565 (N_7565,N_5143,N_4171);
and U7566 (N_7566,N_5778,N_5334);
or U7567 (N_7567,N_5519,N_4114);
nand U7568 (N_7568,N_4095,N_4325);
nand U7569 (N_7569,N_4143,N_4753);
and U7570 (N_7570,N_4659,N_4018);
nand U7571 (N_7571,N_4620,N_5789);
or U7572 (N_7572,N_5822,N_5018);
nor U7573 (N_7573,N_4410,N_5561);
or U7574 (N_7574,N_4242,N_4249);
nand U7575 (N_7575,N_5019,N_4666);
or U7576 (N_7576,N_5636,N_5024);
and U7577 (N_7577,N_4500,N_4021);
or U7578 (N_7578,N_5088,N_5714);
xnor U7579 (N_7579,N_5784,N_5388);
nand U7580 (N_7580,N_4195,N_5142);
nand U7581 (N_7581,N_4339,N_5904);
nor U7582 (N_7582,N_5371,N_4133);
nor U7583 (N_7583,N_4536,N_4969);
or U7584 (N_7584,N_5418,N_4904);
nor U7585 (N_7585,N_4409,N_4993);
and U7586 (N_7586,N_5158,N_4538);
xor U7587 (N_7587,N_4232,N_5339);
xor U7588 (N_7588,N_5944,N_5459);
nor U7589 (N_7589,N_4809,N_5731);
and U7590 (N_7590,N_5442,N_5121);
nor U7591 (N_7591,N_4237,N_5417);
nand U7592 (N_7592,N_4463,N_5326);
nor U7593 (N_7593,N_4291,N_5808);
and U7594 (N_7594,N_5747,N_5696);
nand U7595 (N_7595,N_4601,N_4767);
nor U7596 (N_7596,N_4807,N_4014);
or U7597 (N_7597,N_4215,N_5056);
nor U7598 (N_7598,N_4224,N_4891);
nand U7599 (N_7599,N_5214,N_4674);
and U7600 (N_7600,N_4531,N_4343);
xnor U7601 (N_7601,N_4428,N_5492);
nand U7602 (N_7602,N_4658,N_5550);
and U7603 (N_7603,N_4236,N_5890);
nand U7604 (N_7604,N_4591,N_4833);
and U7605 (N_7605,N_5936,N_4368);
and U7606 (N_7606,N_5079,N_4190);
and U7607 (N_7607,N_4303,N_5265);
nor U7608 (N_7608,N_5806,N_5017);
xor U7609 (N_7609,N_5763,N_5455);
nor U7610 (N_7610,N_4511,N_4183);
and U7611 (N_7611,N_5017,N_4290);
xor U7612 (N_7612,N_4135,N_4585);
or U7613 (N_7613,N_4871,N_5379);
and U7614 (N_7614,N_4716,N_5396);
nand U7615 (N_7615,N_5662,N_4518);
nand U7616 (N_7616,N_4329,N_5911);
nor U7617 (N_7617,N_4634,N_5173);
nor U7618 (N_7618,N_5718,N_4519);
nand U7619 (N_7619,N_5854,N_5300);
or U7620 (N_7620,N_4873,N_5065);
nor U7621 (N_7621,N_4962,N_4462);
xnor U7622 (N_7622,N_4599,N_5720);
nor U7623 (N_7623,N_5656,N_5988);
or U7624 (N_7624,N_4663,N_5455);
nand U7625 (N_7625,N_5820,N_4557);
xnor U7626 (N_7626,N_5607,N_4314);
xnor U7627 (N_7627,N_5152,N_5197);
and U7628 (N_7628,N_4159,N_4365);
xnor U7629 (N_7629,N_5750,N_5583);
nor U7630 (N_7630,N_4153,N_4902);
and U7631 (N_7631,N_5984,N_5694);
and U7632 (N_7632,N_5808,N_4682);
xnor U7633 (N_7633,N_5317,N_4156);
xnor U7634 (N_7634,N_5915,N_5276);
nand U7635 (N_7635,N_4411,N_4716);
xor U7636 (N_7636,N_4257,N_4300);
xor U7637 (N_7637,N_5130,N_4872);
nand U7638 (N_7638,N_5615,N_4184);
nor U7639 (N_7639,N_4531,N_5959);
nand U7640 (N_7640,N_5325,N_5119);
nand U7641 (N_7641,N_4909,N_5159);
or U7642 (N_7642,N_4075,N_5087);
nor U7643 (N_7643,N_5176,N_4669);
and U7644 (N_7644,N_4624,N_5483);
xnor U7645 (N_7645,N_4346,N_5503);
xnor U7646 (N_7646,N_5713,N_5724);
nand U7647 (N_7647,N_5234,N_4554);
nor U7648 (N_7648,N_4037,N_4577);
nor U7649 (N_7649,N_4142,N_5929);
nand U7650 (N_7650,N_4464,N_4739);
nor U7651 (N_7651,N_4301,N_5620);
and U7652 (N_7652,N_5551,N_5139);
and U7653 (N_7653,N_4439,N_4868);
xnor U7654 (N_7654,N_5301,N_4497);
nand U7655 (N_7655,N_5954,N_4574);
or U7656 (N_7656,N_5858,N_5415);
nand U7657 (N_7657,N_5452,N_4687);
nand U7658 (N_7658,N_5311,N_5255);
nor U7659 (N_7659,N_4425,N_5824);
and U7660 (N_7660,N_5868,N_5298);
and U7661 (N_7661,N_5024,N_4186);
xnor U7662 (N_7662,N_4853,N_4269);
and U7663 (N_7663,N_4615,N_5669);
nand U7664 (N_7664,N_4540,N_5644);
and U7665 (N_7665,N_4958,N_4598);
and U7666 (N_7666,N_4759,N_5536);
nor U7667 (N_7667,N_5046,N_4167);
nand U7668 (N_7668,N_5888,N_5367);
nand U7669 (N_7669,N_4586,N_5149);
or U7670 (N_7670,N_5364,N_4063);
xnor U7671 (N_7671,N_4738,N_5502);
and U7672 (N_7672,N_4625,N_4274);
nand U7673 (N_7673,N_4633,N_4210);
nand U7674 (N_7674,N_4494,N_5402);
xor U7675 (N_7675,N_5974,N_5990);
nand U7676 (N_7676,N_5711,N_4332);
nor U7677 (N_7677,N_5827,N_4911);
and U7678 (N_7678,N_4404,N_4178);
xnor U7679 (N_7679,N_4568,N_4053);
or U7680 (N_7680,N_5322,N_5432);
nor U7681 (N_7681,N_5118,N_4419);
nor U7682 (N_7682,N_4557,N_5605);
and U7683 (N_7683,N_4129,N_4955);
xnor U7684 (N_7684,N_5839,N_5457);
nor U7685 (N_7685,N_5993,N_5666);
nand U7686 (N_7686,N_5232,N_5605);
xor U7687 (N_7687,N_4546,N_4513);
and U7688 (N_7688,N_4328,N_5086);
xnor U7689 (N_7689,N_5223,N_4966);
xor U7690 (N_7690,N_5680,N_4296);
or U7691 (N_7691,N_4782,N_4916);
nand U7692 (N_7692,N_4780,N_4979);
nor U7693 (N_7693,N_4400,N_4147);
nor U7694 (N_7694,N_4138,N_4700);
nand U7695 (N_7695,N_4889,N_4882);
and U7696 (N_7696,N_4633,N_5653);
and U7697 (N_7697,N_4526,N_5078);
or U7698 (N_7698,N_5507,N_5516);
nand U7699 (N_7699,N_5586,N_5816);
nand U7700 (N_7700,N_5772,N_4099);
xor U7701 (N_7701,N_4665,N_5819);
or U7702 (N_7702,N_4275,N_4314);
xor U7703 (N_7703,N_5433,N_4823);
nand U7704 (N_7704,N_5575,N_4761);
xnor U7705 (N_7705,N_5219,N_5213);
nor U7706 (N_7706,N_4184,N_5413);
and U7707 (N_7707,N_5299,N_4345);
or U7708 (N_7708,N_5742,N_4805);
and U7709 (N_7709,N_5481,N_4091);
xnor U7710 (N_7710,N_5130,N_4722);
xor U7711 (N_7711,N_4958,N_4629);
or U7712 (N_7712,N_5128,N_5025);
or U7713 (N_7713,N_4189,N_4839);
nand U7714 (N_7714,N_4475,N_5818);
xor U7715 (N_7715,N_5985,N_5483);
nor U7716 (N_7716,N_4129,N_4269);
and U7717 (N_7717,N_4426,N_5569);
and U7718 (N_7718,N_5416,N_4757);
nor U7719 (N_7719,N_5917,N_5989);
or U7720 (N_7720,N_5700,N_4017);
xnor U7721 (N_7721,N_5528,N_5702);
xnor U7722 (N_7722,N_5681,N_5024);
nand U7723 (N_7723,N_4373,N_4061);
xor U7724 (N_7724,N_4128,N_5112);
nand U7725 (N_7725,N_5249,N_4761);
nand U7726 (N_7726,N_5401,N_4143);
or U7727 (N_7727,N_5998,N_5954);
or U7728 (N_7728,N_4176,N_5359);
xnor U7729 (N_7729,N_5721,N_4314);
nand U7730 (N_7730,N_5465,N_4337);
nor U7731 (N_7731,N_4324,N_4329);
and U7732 (N_7732,N_4083,N_5687);
or U7733 (N_7733,N_5254,N_5605);
nor U7734 (N_7734,N_4317,N_4003);
and U7735 (N_7735,N_5452,N_4465);
or U7736 (N_7736,N_5848,N_4216);
nor U7737 (N_7737,N_5944,N_5444);
xor U7738 (N_7738,N_5199,N_4976);
or U7739 (N_7739,N_5259,N_4379);
nand U7740 (N_7740,N_4600,N_4299);
xor U7741 (N_7741,N_5866,N_5163);
or U7742 (N_7742,N_4515,N_5563);
nand U7743 (N_7743,N_4643,N_4827);
and U7744 (N_7744,N_5032,N_5162);
xor U7745 (N_7745,N_5078,N_4274);
nand U7746 (N_7746,N_4522,N_5644);
and U7747 (N_7747,N_5313,N_5885);
nor U7748 (N_7748,N_4673,N_5458);
and U7749 (N_7749,N_5358,N_4575);
nand U7750 (N_7750,N_5818,N_5103);
and U7751 (N_7751,N_4056,N_4805);
nand U7752 (N_7752,N_5472,N_5215);
nand U7753 (N_7753,N_5657,N_4074);
xnor U7754 (N_7754,N_5106,N_5575);
xnor U7755 (N_7755,N_4837,N_5412);
nand U7756 (N_7756,N_5245,N_5978);
nor U7757 (N_7757,N_5129,N_4903);
nor U7758 (N_7758,N_4449,N_5568);
nor U7759 (N_7759,N_4796,N_5823);
and U7760 (N_7760,N_5389,N_4308);
and U7761 (N_7761,N_5535,N_5419);
nand U7762 (N_7762,N_4367,N_4823);
nor U7763 (N_7763,N_4957,N_5324);
nor U7764 (N_7764,N_5460,N_4697);
nor U7765 (N_7765,N_4648,N_5106);
or U7766 (N_7766,N_5855,N_5693);
nor U7767 (N_7767,N_5502,N_4531);
nor U7768 (N_7768,N_5871,N_5601);
nor U7769 (N_7769,N_4067,N_5984);
and U7770 (N_7770,N_4895,N_4125);
nand U7771 (N_7771,N_5358,N_5398);
nor U7772 (N_7772,N_4161,N_5059);
nand U7773 (N_7773,N_5723,N_5930);
or U7774 (N_7774,N_5880,N_5243);
or U7775 (N_7775,N_5841,N_5894);
or U7776 (N_7776,N_4378,N_5586);
xnor U7777 (N_7777,N_4510,N_4438);
and U7778 (N_7778,N_4912,N_5259);
nor U7779 (N_7779,N_4769,N_5673);
or U7780 (N_7780,N_4812,N_4761);
nor U7781 (N_7781,N_4867,N_5774);
or U7782 (N_7782,N_4398,N_5145);
nor U7783 (N_7783,N_5133,N_4669);
and U7784 (N_7784,N_5937,N_5945);
nor U7785 (N_7785,N_4090,N_5827);
xor U7786 (N_7786,N_4566,N_5377);
xor U7787 (N_7787,N_4598,N_5685);
nor U7788 (N_7788,N_4686,N_5133);
or U7789 (N_7789,N_4337,N_4660);
nor U7790 (N_7790,N_5309,N_5621);
nand U7791 (N_7791,N_4985,N_4190);
nor U7792 (N_7792,N_5291,N_5477);
or U7793 (N_7793,N_5668,N_4759);
and U7794 (N_7794,N_4938,N_4910);
xnor U7795 (N_7795,N_4038,N_4869);
xor U7796 (N_7796,N_5326,N_5948);
xor U7797 (N_7797,N_5424,N_4544);
or U7798 (N_7798,N_5822,N_4640);
nand U7799 (N_7799,N_4193,N_4138);
and U7800 (N_7800,N_5659,N_4459);
nand U7801 (N_7801,N_5211,N_4449);
and U7802 (N_7802,N_4378,N_4675);
xnor U7803 (N_7803,N_5444,N_4915);
and U7804 (N_7804,N_5096,N_5277);
xnor U7805 (N_7805,N_4089,N_5403);
nor U7806 (N_7806,N_5563,N_5958);
nand U7807 (N_7807,N_5014,N_5072);
and U7808 (N_7808,N_4712,N_5723);
xnor U7809 (N_7809,N_5752,N_4260);
xor U7810 (N_7810,N_4438,N_5560);
or U7811 (N_7811,N_4728,N_4324);
nand U7812 (N_7812,N_5211,N_5756);
nand U7813 (N_7813,N_4557,N_4333);
and U7814 (N_7814,N_5092,N_5500);
xor U7815 (N_7815,N_4342,N_4150);
or U7816 (N_7816,N_4988,N_4275);
and U7817 (N_7817,N_4092,N_4127);
xor U7818 (N_7818,N_5990,N_4681);
or U7819 (N_7819,N_4264,N_4965);
or U7820 (N_7820,N_4833,N_4414);
or U7821 (N_7821,N_5378,N_5973);
xor U7822 (N_7822,N_4443,N_4243);
nor U7823 (N_7823,N_4244,N_5291);
or U7824 (N_7824,N_5499,N_5966);
or U7825 (N_7825,N_4993,N_4109);
and U7826 (N_7826,N_4489,N_5738);
xor U7827 (N_7827,N_4973,N_5653);
xor U7828 (N_7828,N_5959,N_5113);
nand U7829 (N_7829,N_5737,N_4914);
and U7830 (N_7830,N_5359,N_5902);
or U7831 (N_7831,N_4275,N_4764);
and U7832 (N_7832,N_4169,N_5909);
and U7833 (N_7833,N_5028,N_4161);
nor U7834 (N_7834,N_5467,N_4287);
and U7835 (N_7835,N_5274,N_4643);
nand U7836 (N_7836,N_4436,N_5746);
xnor U7837 (N_7837,N_5210,N_5211);
and U7838 (N_7838,N_4644,N_4979);
nor U7839 (N_7839,N_4142,N_4314);
and U7840 (N_7840,N_5095,N_5627);
nor U7841 (N_7841,N_5880,N_5859);
and U7842 (N_7842,N_5832,N_4419);
xnor U7843 (N_7843,N_5642,N_4187);
xnor U7844 (N_7844,N_5032,N_4382);
and U7845 (N_7845,N_5453,N_4938);
xnor U7846 (N_7846,N_5032,N_5095);
nor U7847 (N_7847,N_5426,N_4603);
xor U7848 (N_7848,N_4177,N_5121);
and U7849 (N_7849,N_4646,N_4677);
nor U7850 (N_7850,N_4737,N_4101);
or U7851 (N_7851,N_4499,N_5107);
and U7852 (N_7852,N_4081,N_5677);
and U7853 (N_7853,N_5716,N_4057);
or U7854 (N_7854,N_5208,N_4137);
nand U7855 (N_7855,N_5621,N_5348);
and U7856 (N_7856,N_5506,N_5852);
nor U7857 (N_7857,N_4848,N_4597);
nor U7858 (N_7858,N_5340,N_4193);
and U7859 (N_7859,N_4411,N_5151);
and U7860 (N_7860,N_5942,N_5904);
nand U7861 (N_7861,N_5534,N_4773);
nor U7862 (N_7862,N_5764,N_4544);
or U7863 (N_7863,N_5155,N_5331);
xnor U7864 (N_7864,N_5835,N_5645);
nor U7865 (N_7865,N_5658,N_4407);
and U7866 (N_7866,N_4263,N_4224);
nor U7867 (N_7867,N_5450,N_5995);
nor U7868 (N_7868,N_4147,N_4621);
or U7869 (N_7869,N_5522,N_5182);
or U7870 (N_7870,N_5284,N_5935);
and U7871 (N_7871,N_5866,N_4839);
xor U7872 (N_7872,N_4946,N_4457);
or U7873 (N_7873,N_4001,N_5600);
nand U7874 (N_7874,N_5728,N_4693);
nor U7875 (N_7875,N_5803,N_4716);
or U7876 (N_7876,N_4883,N_5404);
nor U7877 (N_7877,N_5327,N_4219);
or U7878 (N_7878,N_5873,N_4575);
nor U7879 (N_7879,N_5846,N_5373);
nand U7880 (N_7880,N_5134,N_4589);
and U7881 (N_7881,N_4215,N_5402);
or U7882 (N_7882,N_4182,N_4843);
nand U7883 (N_7883,N_4485,N_4833);
nor U7884 (N_7884,N_4591,N_5769);
and U7885 (N_7885,N_4172,N_5394);
xor U7886 (N_7886,N_4052,N_5606);
nor U7887 (N_7887,N_5536,N_4935);
nand U7888 (N_7888,N_4063,N_4642);
or U7889 (N_7889,N_4353,N_4552);
or U7890 (N_7890,N_5693,N_4551);
nor U7891 (N_7891,N_4301,N_4710);
and U7892 (N_7892,N_4849,N_4438);
xnor U7893 (N_7893,N_5520,N_4953);
or U7894 (N_7894,N_5518,N_5375);
or U7895 (N_7895,N_4375,N_5522);
nand U7896 (N_7896,N_5794,N_5426);
xor U7897 (N_7897,N_5660,N_5857);
nand U7898 (N_7898,N_5312,N_5041);
and U7899 (N_7899,N_5880,N_5038);
and U7900 (N_7900,N_5646,N_4946);
and U7901 (N_7901,N_4358,N_5518);
xnor U7902 (N_7902,N_5416,N_4429);
xor U7903 (N_7903,N_5615,N_4525);
and U7904 (N_7904,N_4173,N_5609);
nand U7905 (N_7905,N_5757,N_4262);
nor U7906 (N_7906,N_4187,N_5484);
nand U7907 (N_7907,N_4684,N_5237);
nand U7908 (N_7908,N_4201,N_4322);
nor U7909 (N_7909,N_4876,N_5322);
or U7910 (N_7910,N_4373,N_5391);
or U7911 (N_7911,N_4702,N_4290);
or U7912 (N_7912,N_4553,N_5501);
xor U7913 (N_7913,N_5405,N_4490);
and U7914 (N_7914,N_4957,N_4437);
and U7915 (N_7915,N_5600,N_5683);
nor U7916 (N_7916,N_5612,N_4653);
xor U7917 (N_7917,N_4481,N_4435);
nor U7918 (N_7918,N_4497,N_5188);
xor U7919 (N_7919,N_4745,N_4763);
nor U7920 (N_7920,N_5089,N_5705);
nor U7921 (N_7921,N_5227,N_4001);
xor U7922 (N_7922,N_5507,N_5926);
nor U7923 (N_7923,N_4220,N_4147);
and U7924 (N_7924,N_4318,N_5445);
nand U7925 (N_7925,N_5133,N_4788);
nand U7926 (N_7926,N_5087,N_4739);
nor U7927 (N_7927,N_5494,N_5262);
nor U7928 (N_7928,N_4665,N_5331);
nor U7929 (N_7929,N_4829,N_5518);
nor U7930 (N_7930,N_4873,N_4132);
nor U7931 (N_7931,N_5479,N_4390);
nor U7932 (N_7932,N_4392,N_4844);
xnor U7933 (N_7933,N_4451,N_5241);
or U7934 (N_7934,N_4949,N_4718);
or U7935 (N_7935,N_4720,N_5513);
nor U7936 (N_7936,N_4022,N_4972);
xnor U7937 (N_7937,N_5135,N_5717);
nor U7938 (N_7938,N_5015,N_4691);
and U7939 (N_7939,N_4176,N_5207);
xor U7940 (N_7940,N_4378,N_5355);
or U7941 (N_7941,N_5906,N_4750);
xor U7942 (N_7942,N_4593,N_5208);
and U7943 (N_7943,N_4979,N_4155);
and U7944 (N_7944,N_4997,N_5981);
xor U7945 (N_7945,N_5858,N_4988);
or U7946 (N_7946,N_4126,N_5705);
or U7947 (N_7947,N_4652,N_4499);
nand U7948 (N_7948,N_5870,N_5974);
xnor U7949 (N_7949,N_4440,N_5535);
and U7950 (N_7950,N_5188,N_5622);
and U7951 (N_7951,N_4492,N_4143);
xor U7952 (N_7952,N_4740,N_5291);
nand U7953 (N_7953,N_4421,N_5602);
xor U7954 (N_7954,N_5220,N_4078);
nor U7955 (N_7955,N_5714,N_4913);
and U7956 (N_7956,N_4165,N_4137);
and U7957 (N_7957,N_4808,N_5447);
and U7958 (N_7958,N_4618,N_4044);
nor U7959 (N_7959,N_4519,N_5043);
nand U7960 (N_7960,N_5481,N_4503);
or U7961 (N_7961,N_4560,N_4248);
or U7962 (N_7962,N_4807,N_4585);
nand U7963 (N_7963,N_5339,N_4422);
xnor U7964 (N_7964,N_5339,N_5236);
or U7965 (N_7965,N_5966,N_4084);
xor U7966 (N_7966,N_5067,N_5218);
and U7967 (N_7967,N_4564,N_4327);
nor U7968 (N_7968,N_5933,N_5049);
nor U7969 (N_7969,N_4853,N_5651);
xnor U7970 (N_7970,N_5240,N_5857);
nor U7971 (N_7971,N_4013,N_5071);
or U7972 (N_7972,N_5518,N_4943);
nand U7973 (N_7973,N_4921,N_4647);
nor U7974 (N_7974,N_4794,N_5051);
or U7975 (N_7975,N_4560,N_5431);
or U7976 (N_7976,N_5847,N_4378);
and U7977 (N_7977,N_4620,N_4234);
nand U7978 (N_7978,N_4826,N_4392);
nor U7979 (N_7979,N_4540,N_5483);
nor U7980 (N_7980,N_5867,N_4201);
or U7981 (N_7981,N_4209,N_5124);
xor U7982 (N_7982,N_4796,N_4130);
nand U7983 (N_7983,N_4682,N_5846);
and U7984 (N_7984,N_4196,N_5497);
xor U7985 (N_7985,N_4866,N_4521);
nand U7986 (N_7986,N_4895,N_5492);
nor U7987 (N_7987,N_4735,N_5434);
and U7988 (N_7988,N_4127,N_4445);
and U7989 (N_7989,N_5970,N_5117);
or U7990 (N_7990,N_5253,N_5792);
nor U7991 (N_7991,N_4880,N_5540);
and U7992 (N_7992,N_5955,N_5040);
nand U7993 (N_7993,N_4851,N_4734);
and U7994 (N_7994,N_5922,N_4414);
nor U7995 (N_7995,N_4759,N_4751);
xor U7996 (N_7996,N_5523,N_5933);
or U7997 (N_7997,N_4344,N_5852);
or U7998 (N_7998,N_5035,N_5347);
nor U7999 (N_7999,N_4906,N_5735);
nand U8000 (N_8000,N_7347,N_6175);
nor U8001 (N_8001,N_6152,N_7410);
xor U8002 (N_8002,N_6696,N_7663);
nand U8003 (N_8003,N_6521,N_6868);
nand U8004 (N_8004,N_6739,N_6370);
xnor U8005 (N_8005,N_7291,N_6892);
and U8006 (N_8006,N_6207,N_7704);
xor U8007 (N_8007,N_6281,N_6598);
nor U8008 (N_8008,N_7137,N_6493);
xnor U8009 (N_8009,N_6985,N_7354);
nor U8010 (N_8010,N_6742,N_7191);
nand U8011 (N_8011,N_7668,N_6421);
and U8012 (N_8012,N_6798,N_6267);
xnor U8013 (N_8013,N_7740,N_7956);
nand U8014 (N_8014,N_7068,N_7805);
xor U8015 (N_8015,N_7705,N_6752);
xnor U8016 (N_8016,N_7263,N_6271);
and U8017 (N_8017,N_6083,N_6825);
xnor U8018 (N_8018,N_6070,N_6209);
nand U8019 (N_8019,N_6645,N_6806);
nor U8020 (N_8020,N_6098,N_6009);
or U8021 (N_8021,N_6389,N_6213);
nand U8022 (N_8022,N_6390,N_6460);
and U8023 (N_8023,N_7276,N_7193);
nor U8024 (N_8024,N_7883,N_6865);
nor U8025 (N_8025,N_6140,N_6080);
or U8026 (N_8026,N_6759,N_7449);
xnor U8027 (N_8027,N_7848,N_6330);
nor U8028 (N_8028,N_6566,N_6807);
and U8029 (N_8029,N_7625,N_7101);
nor U8030 (N_8030,N_7149,N_7031);
or U8031 (N_8031,N_6135,N_7714);
nor U8032 (N_8032,N_7759,N_6294);
nor U8033 (N_8033,N_7837,N_6369);
and U8034 (N_8034,N_6901,N_7262);
xor U8035 (N_8035,N_7116,N_6932);
xor U8036 (N_8036,N_7044,N_6260);
and U8037 (N_8037,N_6804,N_6795);
or U8038 (N_8038,N_6220,N_6619);
and U8039 (N_8039,N_6709,N_7008);
nand U8040 (N_8040,N_6134,N_7758);
xor U8041 (N_8041,N_7074,N_7878);
and U8042 (N_8042,N_6713,N_6764);
nor U8043 (N_8043,N_7158,N_6324);
nor U8044 (N_8044,N_6494,N_7588);
nor U8045 (N_8045,N_6897,N_6719);
nand U8046 (N_8046,N_7518,N_6087);
and U8047 (N_8047,N_6669,N_7983);
and U8048 (N_8048,N_6658,N_6238);
nor U8049 (N_8049,N_7159,N_6997);
nand U8050 (N_8050,N_6419,N_6636);
or U8051 (N_8051,N_6071,N_7160);
nor U8052 (N_8052,N_6151,N_6304);
or U8053 (N_8053,N_7596,N_6986);
xnor U8054 (N_8054,N_7648,N_7163);
nor U8055 (N_8055,N_7363,N_7283);
or U8056 (N_8056,N_7808,N_6477);
or U8057 (N_8057,N_7634,N_6156);
nand U8058 (N_8058,N_7317,N_7818);
nor U8059 (N_8059,N_7644,N_6301);
or U8060 (N_8060,N_7732,N_7122);
nand U8061 (N_8061,N_7350,N_7065);
nor U8062 (N_8062,N_6553,N_6778);
or U8063 (N_8063,N_6474,N_7810);
nor U8064 (N_8064,N_6699,N_7426);
nand U8065 (N_8065,N_7982,N_6172);
and U8066 (N_8066,N_6701,N_7215);
xnor U8067 (N_8067,N_7378,N_7667);
or U8068 (N_8068,N_7735,N_7727);
nand U8069 (N_8069,N_7132,N_6189);
or U8070 (N_8070,N_7840,N_7242);
nand U8071 (N_8071,N_7854,N_7573);
and U8072 (N_8072,N_6791,N_7995);
or U8073 (N_8073,N_7693,N_6674);
nor U8074 (N_8074,N_7866,N_6657);
or U8075 (N_8075,N_6782,N_6184);
and U8076 (N_8076,N_7485,N_7201);
xor U8077 (N_8077,N_6854,N_6642);
nand U8078 (N_8078,N_7330,N_6857);
xnor U8079 (N_8079,N_7429,N_6763);
nor U8080 (N_8080,N_6983,N_7670);
nand U8081 (N_8081,N_7974,N_6864);
nor U8082 (N_8082,N_6462,N_7170);
and U8083 (N_8083,N_7722,N_6218);
or U8084 (N_8084,N_6451,N_6679);
or U8085 (N_8085,N_7367,N_7927);
nand U8086 (N_8086,N_7130,N_6723);
or U8087 (N_8087,N_7638,N_7233);
nand U8088 (N_8088,N_7587,N_7297);
xnor U8089 (N_8089,N_7929,N_6092);
and U8090 (N_8090,N_7917,N_7277);
xor U8091 (N_8091,N_7738,N_6736);
nand U8092 (N_8092,N_7100,N_7084);
nor U8093 (N_8093,N_7308,N_7779);
xor U8094 (N_8094,N_6393,N_6362);
or U8095 (N_8095,N_7076,N_7822);
or U8096 (N_8096,N_7870,N_6771);
nor U8097 (N_8097,N_6289,N_6631);
or U8098 (N_8098,N_6863,N_7846);
xnor U8099 (N_8099,N_7978,N_7522);
nand U8100 (N_8100,N_7821,N_6131);
xor U8101 (N_8101,N_6240,N_7775);
and U8102 (N_8102,N_7348,N_7510);
nor U8103 (N_8103,N_6177,N_6671);
nand U8104 (N_8104,N_7585,N_7462);
and U8105 (N_8105,N_7112,N_7636);
or U8106 (N_8106,N_7285,N_6746);
xnor U8107 (N_8107,N_7453,N_6323);
and U8108 (N_8108,N_6327,N_6517);
and U8109 (N_8109,N_6640,N_7514);
xnor U8110 (N_8110,N_6809,N_7723);
and U8111 (N_8111,N_6457,N_7405);
and U8112 (N_8112,N_6833,N_6757);
and U8113 (N_8113,N_6168,N_6575);
or U8114 (N_8114,N_6380,N_6020);
nand U8115 (N_8115,N_6832,N_7706);
nand U8116 (N_8116,N_7454,N_6336);
nand U8117 (N_8117,N_6247,N_7024);
nand U8118 (N_8118,N_6905,N_6360);
or U8119 (N_8119,N_7914,N_7039);
nor U8120 (N_8120,N_6384,N_7582);
nand U8121 (N_8121,N_6193,N_6399);
or U8122 (N_8122,N_6257,N_6141);
nor U8123 (N_8123,N_6202,N_7411);
nor U8124 (N_8124,N_7835,N_7649);
or U8125 (N_8125,N_7515,N_7994);
and U8126 (N_8126,N_7279,N_7494);
nor U8127 (N_8127,N_6219,N_7780);
or U8128 (N_8128,N_6871,N_6149);
nor U8129 (N_8129,N_6208,N_7507);
nand U8130 (N_8130,N_6483,N_7432);
nor U8131 (N_8131,N_7896,N_7496);
xnor U8132 (N_8132,N_7105,N_7940);
nor U8133 (N_8133,N_6976,N_7859);
nand U8134 (N_8134,N_7402,N_7544);
and U8135 (N_8135,N_7671,N_6758);
nand U8136 (N_8136,N_6712,N_7408);
or U8137 (N_8137,N_6632,N_6125);
nand U8138 (N_8138,N_7369,N_7689);
xnor U8139 (N_8139,N_7501,N_6829);
xor U8140 (N_8140,N_6826,N_7568);
nor U8141 (N_8141,N_6760,N_7679);
and U8142 (N_8142,N_7968,N_7465);
and U8143 (N_8143,N_6443,N_6527);
nand U8144 (N_8144,N_7591,N_7245);
nor U8145 (N_8145,N_6600,N_7628);
or U8146 (N_8146,N_6287,N_6046);
xor U8147 (N_8147,N_6680,N_6879);
nor U8148 (N_8148,N_7003,N_7652);
xnor U8149 (N_8149,N_6793,N_7920);
nand U8150 (N_8150,N_6463,N_7803);
xor U8151 (N_8151,N_7907,N_7720);
and U8152 (N_8152,N_6023,N_7404);
nand U8153 (N_8153,N_6198,N_7483);
nand U8154 (N_8154,N_6303,N_6533);
or U8155 (N_8155,N_7928,N_7502);
nor U8156 (N_8156,N_7087,N_7776);
or U8157 (N_8157,N_6424,N_7179);
xnor U8158 (N_8158,N_7401,N_7653);
xor U8159 (N_8159,N_7126,N_7464);
xnor U8160 (N_8160,N_6053,N_7340);
nand U8161 (N_8161,N_7578,N_7358);
nand U8162 (N_8162,N_7612,N_7973);
or U8163 (N_8163,N_7232,N_7890);
or U8164 (N_8164,N_6111,N_6112);
and U8165 (N_8165,N_7725,N_7615);
nand U8166 (N_8166,N_6993,N_7602);
nand U8167 (N_8167,N_7447,N_6430);
nand U8168 (N_8168,N_6122,N_6041);
and U8169 (N_8169,N_6497,N_6056);
nand U8170 (N_8170,N_6059,N_6559);
and U8171 (N_8171,N_6613,N_7490);
nor U8172 (N_8172,N_7998,N_6848);
nor U8173 (N_8173,N_7082,N_7187);
nand U8174 (N_8174,N_6311,N_7287);
and U8175 (N_8175,N_7230,N_6475);
xnor U8176 (N_8176,N_7858,N_7083);
xnor U8177 (N_8177,N_7841,N_6639);
and U8178 (N_8178,N_7090,N_6312);
or U8179 (N_8179,N_7060,N_6363);
xnor U8180 (N_8180,N_6341,N_7729);
nor U8181 (N_8181,N_6085,N_7417);
xor U8182 (N_8182,N_6565,N_7177);
nand U8183 (N_8183,N_6622,N_7796);
or U8184 (N_8184,N_7924,N_6291);
and U8185 (N_8185,N_6423,N_6138);
nor U8186 (N_8186,N_6322,N_6651);
nor U8187 (N_8187,N_6345,N_6524);
xor U8188 (N_8188,N_7111,N_6919);
or U8189 (N_8189,N_7434,N_6195);
or U8190 (N_8190,N_6552,N_6132);
nand U8191 (N_8191,N_7202,N_7984);
or U8192 (N_8192,N_6979,N_6342);
nor U8193 (N_8193,N_6990,N_7512);
nor U8194 (N_8194,N_6358,N_7477);
nand U8195 (N_8195,N_7004,N_6837);
or U8196 (N_8196,N_6163,N_7220);
xor U8197 (N_8197,N_7071,N_6678);
xor U8198 (N_8198,N_7042,N_6321);
and U8199 (N_8199,N_6922,N_7366);
nor U8200 (N_8200,N_6274,N_7356);
nand U8201 (N_8201,N_6432,N_7343);
nand U8202 (N_8202,N_6373,N_7789);
xnor U8203 (N_8203,N_6957,N_7875);
or U8204 (N_8204,N_6016,N_6144);
xor U8205 (N_8205,N_6718,N_7659);
nand U8206 (N_8206,N_6654,N_7229);
nand U8207 (N_8207,N_6623,N_6661);
xnor U8208 (N_8208,N_6630,N_7150);
or U8209 (N_8209,N_7416,N_6438);
xor U8210 (N_8210,N_6968,N_7696);
and U8211 (N_8211,N_7892,N_7590);
and U8212 (N_8212,N_7894,N_7761);
and U8213 (N_8213,N_7778,N_7771);
and U8214 (N_8214,N_6212,N_7221);
nor U8215 (N_8215,N_7395,N_7254);
and U8216 (N_8216,N_7196,N_6627);
nor U8217 (N_8217,N_7499,N_7344);
nand U8218 (N_8218,N_7383,N_6347);
and U8219 (N_8219,N_6811,N_6297);
and U8220 (N_8220,N_6720,N_6013);
nand U8221 (N_8221,N_6354,N_7301);
xor U8222 (N_8222,N_6405,N_7881);
nor U8223 (N_8223,N_6402,N_7981);
nor U8224 (N_8224,N_6729,N_7373);
nand U8225 (N_8225,N_6526,N_7933);
and U8226 (N_8226,N_6467,N_6861);
xnor U8227 (N_8227,N_6052,N_7852);
xnor U8228 (N_8228,N_7651,N_6387);
nor U8229 (N_8229,N_7533,N_7397);
nand U8230 (N_8230,N_7786,N_7709);
xnor U8231 (N_8231,N_7794,N_7884);
or U8232 (N_8232,N_7699,N_6556);
nand U8233 (N_8233,N_7057,N_6139);
and U8234 (N_8234,N_7966,N_6513);
nor U8235 (N_8235,N_6692,N_7941);
xnor U8236 (N_8236,N_7244,N_7099);
or U8237 (N_8237,N_7156,N_7631);
and U8238 (N_8238,N_6884,N_7799);
and U8239 (N_8239,N_7175,N_6024);
nand U8240 (N_8240,N_7441,N_6256);
or U8241 (N_8241,N_6150,N_7181);
nor U8242 (N_8242,N_6043,N_6855);
or U8243 (N_8243,N_6398,N_7213);
or U8244 (N_8244,N_6368,N_6951);
xnor U8245 (N_8245,N_6844,N_6616);
xor U8246 (N_8246,N_6136,N_6996);
xor U8247 (N_8247,N_7227,N_6755);
and U8248 (N_8248,N_7243,N_7888);
or U8249 (N_8249,N_7406,N_6183);
and U8250 (N_8250,N_6974,N_6359);
nand U8251 (N_8251,N_6120,N_6621);
xnor U8252 (N_8252,N_6000,N_6454);
xor U8253 (N_8253,N_7570,N_6749);
and U8254 (N_8254,N_7467,N_6687);
or U8255 (N_8255,N_7007,N_7571);
and U8256 (N_8256,N_6081,N_6610);
or U8257 (N_8257,N_6102,N_6383);
nand U8258 (N_8258,N_6813,N_7751);
and U8259 (N_8259,N_7937,N_6581);
and U8260 (N_8260,N_7479,N_7932);
nor U8261 (N_8261,N_7601,N_7530);
or U8262 (N_8262,N_6110,N_7463);
or U8263 (N_8263,N_7773,N_7619);
xnor U8264 (N_8264,N_6499,N_7903);
nand U8265 (N_8265,N_6529,N_6515);
or U8266 (N_8266,N_6551,N_7214);
nand U8267 (N_8267,N_6505,N_6061);
nor U8268 (N_8268,N_6594,N_7802);
and U8269 (N_8269,N_6506,N_6532);
or U8270 (N_8270,N_7639,N_6744);
or U8271 (N_8271,N_6166,N_7609);
or U8272 (N_8272,N_6821,N_6548);
or U8273 (N_8273,N_6161,N_7461);
nand U8274 (N_8274,N_7091,N_7136);
nand U8275 (N_8275,N_6950,N_7339);
and U8276 (N_8276,N_6650,N_7577);
xnor U8277 (N_8277,N_6038,N_7938);
nor U8278 (N_8278,N_7868,N_6465);
nor U8279 (N_8279,N_6171,N_6040);
xor U8280 (N_8280,N_7774,N_7707);
and U8281 (N_8281,N_7528,N_6980);
or U8282 (N_8282,N_7346,N_7509);
nand U8283 (N_8283,N_6534,N_7217);
xor U8284 (N_8284,N_6512,N_6253);
nand U8285 (N_8285,N_6285,N_6444);
nand U8286 (N_8286,N_7874,N_6843);
nand U8287 (N_8287,N_6767,N_6459);
or U8288 (N_8288,N_6649,N_6776);
nand U8289 (N_8289,N_7944,N_6747);
nor U8290 (N_8290,N_7660,N_6181);
xor U8291 (N_8291,N_7913,N_6337);
nand U8292 (N_8292,N_7764,N_6113);
nand U8293 (N_8293,N_6574,N_7445);
and U8294 (N_8294,N_7828,N_6891);
or U8295 (N_8295,N_6819,N_7311);
nand U8296 (N_8296,N_7341,N_7152);
nand U8297 (N_8297,N_7986,N_7438);
xor U8298 (N_8298,N_7621,N_7425);
xor U8299 (N_8299,N_7166,N_7716);
xnor U8300 (N_8300,N_6894,N_7294);
nand U8301 (N_8301,N_7873,N_7919);
and U8302 (N_8302,N_7871,N_7752);
nor U8303 (N_8303,N_7123,N_7532);
and U8304 (N_8304,N_6708,N_7926);
and U8305 (N_8305,N_7041,N_6391);
xnor U8306 (N_8306,N_7414,N_7918);
nor U8307 (N_8307,N_7880,N_7320);
or U8308 (N_8308,N_6114,N_6277);
nand U8309 (N_8309,N_6266,N_7993);
and U8310 (N_8310,N_6039,N_6075);
and U8311 (N_8311,N_6774,N_6576);
xnor U8312 (N_8312,N_7807,N_6873);
or U8313 (N_8313,N_6376,N_7203);
nor U8314 (N_8314,N_6780,N_6118);
or U8315 (N_8315,N_7012,N_7174);
and U8316 (N_8316,N_6557,N_7225);
and U8317 (N_8317,N_6935,N_6196);
nand U8318 (N_8318,N_7027,N_6721);
nor U8319 (N_8319,N_7876,N_7762);
nor U8320 (N_8320,N_7692,N_6447);
nand U8321 (N_8321,N_6918,N_6305);
or U8322 (N_8322,N_7861,N_7106);
xor U8323 (N_8323,N_6597,N_7862);
xnor U8324 (N_8324,N_7258,N_7026);
nor U8325 (N_8325,N_6191,N_6546);
and U8326 (N_8326,N_6062,N_7384);
or U8327 (N_8327,N_6890,N_7249);
nor U8328 (N_8328,N_6355,N_6593);
and U8329 (N_8329,N_6072,N_6555);
nor U8330 (N_8330,N_7763,N_6981);
and U8331 (N_8331,N_6801,N_7872);
nor U8332 (N_8332,N_6893,N_6302);
xor U8333 (N_8333,N_7669,N_6488);
nor U8334 (N_8334,N_6315,N_7192);
and U8335 (N_8335,N_6262,N_6353);
and U8336 (N_8336,N_7478,N_7307);
nor U8337 (N_8337,N_7856,N_7228);
and U8338 (N_8338,N_6695,N_7288);
or U8339 (N_8339,N_7772,N_6940);
nor U8340 (N_8340,N_6796,N_6895);
or U8341 (N_8341,N_6814,N_6924);
and U8342 (N_8342,N_7538,N_7980);
nor U8343 (N_8343,N_7857,N_7239);
and U8344 (N_8344,N_7672,N_6216);
nor U8345 (N_8345,N_6926,N_6299);
nand U8346 (N_8346,N_7142,N_7853);
or U8347 (N_8347,N_6944,N_7409);
xnor U8348 (N_8348,N_7766,N_6668);
nand U8349 (N_8349,N_6751,N_6022);
and U8350 (N_8350,N_7224,N_6095);
nor U8351 (N_8351,N_7186,N_6265);
nor U8352 (N_8352,N_6280,N_7198);
nand U8353 (N_8353,N_6605,N_7999);
or U8354 (N_8354,N_6766,N_6603);
or U8355 (N_8355,N_7726,N_6915);
xor U8356 (N_8356,N_7327,N_7690);
xnor U8357 (N_8357,N_6628,N_7143);
xnor U8358 (N_8358,N_7313,N_7593);
and U8359 (N_8359,N_6730,N_7023);
xnor U8360 (N_8360,N_6648,N_7744);
and U8361 (N_8361,N_6361,N_6777);
and U8362 (N_8362,N_6820,N_7559);
nand U8363 (N_8363,N_7172,N_7902);
or U8364 (N_8364,N_6033,N_7627);
and U8365 (N_8365,N_6756,N_6035);
and U8366 (N_8366,N_7178,N_7419);
nor U8367 (N_8367,N_6587,N_7148);
nand U8368 (N_8368,N_6002,N_7792);
or U8369 (N_8369,N_6550,N_7931);
xor U8370 (N_8370,N_7540,N_7812);
and U8371 (N_8371,N_6026,N_6316);
and U8372 (N_8372,N_6097,N_6270);
or U8373 (N_8373,N_6818,N_7289);
xor U8374 (N_8374,N_7210,N_6828);
and U8375 (N_8375,N_7770,N_7829);
nor U8376 (N_8376,N_7377,N_7739);
or U8377 (N_8377,N_6231,N_6292);
and U8378 (N_8378,N_6065,N_7484);
xor U8379 (N_8379,N_7519,N_6914);
xnor U8380 (N_8380,N_7131,N_7686);
nor U8381 (N_8381,N_7736,N_7169);
nand U8382 (N_8382,N_6074,N_6812);
or U8383 (N_8383,N_7022,N_6929);
nand U8384 (N_8384,N_7552,N_6885);
nor U8385 (N_8385,N_7877,N_6842);
and U8386 (N_8386,N_6822,N_6750);
xnor U8387 (N_8387,N_7013,N_7608);
or U8388 (N_8388,N_6706,N_7475);
nor U8389 (N_8389,N_7019,N_6579);
xnor U8390 (N_8390,N_7269,N_6235);
and U8391 (N_8391,N_6063,N_7618);
nor U8392 (N_8392,N_6977,N_6229);
and U8393 (N_8393,N_7115,N_7053);
nand U8394 (N_8394,N_6364,N_7657);
and U8395 (N_8395,N_7960,N_7760);
or U8396 (N_8396,N_7543,N_6006);
or U8397 (N_8397,N_6442,N_6217);
xor U8398 (N_8398,N_7604,N_6954);
nand U8399 (N_8399,N_7094,N_6167);
or U8400 (N_8400,N_7492,N_7581);
xor U8401 (N_8401,N_7466,N_7715);
nand U8402 (N_8402,N_6400,N_7468);
nand U8403 (N_8403,N_7240,N_6934);
nand U8404 (N_8404,N_6561,N_7266);
xnor U8405 (N_8405,N_7379,N_7887);
xnor U8406 (N_8406,N_6704,N_7079);
nor U8407 (N_8407,N_6414,N_6510);
nor U8408 (N_8408,N_6049,N_7531);
nand U8409 (N_8409,N_7038,N_6146);
nand U8410 (N_8410,N_7793,N_6728);
nand U8411 (N_8411,N_7171,N_6458);
xnor U8412 (N_8412,N_6624,N_6965);
nor U8413 (N_8413,N_7403,N_6525);
and U8414 (N_8414,N_7002,N_7700);
and U8415 (N_8415,N_6810,N_7948);
or U8416 (N_8416,N_7626,N_6130);
nor U8417 (N_8417,N_6276,N_6275);
xor U8418 (N_8418,N_7556,N_7867);
xor U8419 (N_8419,N_7635,N_6314);
and U8420 (N_8420,N_6356,N_7879);
and U8421 (N_8421,N_6325,N_6582);
nor U8422 (N_8422,N_6154,N_6121);
nor U8423 (N_8423,N_7072,N_7349);
nor U8424 (N_8424,N_6164,N_6346);
and U8425 (N_8425,N_6137,N_6975);
and U8426 (N_8426,N_7088,N_6123);
and U8427 (N_8427,N_7309,N_7959);
or U8428 (N_8428,N_7503,N_7421);
nor U8429 (N_8429,N_6057,N_6007);
nand U8430 (N_8430,N_7505,N_7458);
xor U8431 (N_8431,N_7691,N_7730);
or U8432 (N_8432,N_6602,N_6158);
or U8433 (N_8433,N_6288,N_7357);
nand U8434 (N_8434,N_6541,N_7655);
or U8435 (N_8435,N_7493,N_6601);
or U8436 (N_8436,N_7371,N_6931);
nor U8437 (N_8437,N_6883,N_6108);
or U8438 (N_8438,N_6169,N_6381);
xnor U8439 (N_8439,N_7062,N_6439);
or U8440 (N_8440,N_7190,N_7260);
nor U8441 (N_8441,N_6044,N_7610);
xor U8442 (N_8442,N_7656,N_6831);
nor U8443 (N_8443,N_7117,N_6745);
nand U8444 (N_8444,N_7476,N_7089);
or U8445 (N_8445,N_6567,N_6994);
or U8446 (N_8446,N_7048,N_6786);
or U8447 (N_8447,N_6662,N_6964);
and U8448 (N_8448,N_6272,N_7860);
nand U8449 (N_8449,N_7145,N_6664);
nand U8450 (N_8450,N_7180,N_6875);
xnor U8451 (N_8451,N_7970,N_6609);
and U8452 (N_8452,N_7574,N_7708);
nor U8453 (N_8453,N_6435,N_7553);
nand U8454 (N_8454,N_7248,N_6107);
nor U8455 (N_8455,N_7303,N_7208);
xnor U8456 (N_8456,N_6549,N_6003);
nand U8457 (N_8457,N_6468,N_6273);
xnor U8458 (N_8458,N_7731,N_6055);
nand U8459 (N_8459,N_6343,N_6104);
nor U8460 (N_8460,N_7790,N_6660);
and U8461 (N_8461,N_6881,N_6449);
nor U8462 (N_8462,N_6332,N_6836);
xnor U8463 (N_8463,N_6320,N_6082);
and U8464 (N_8464,N_7650,N_6481);
nor U8465 (N_8465,N_7755,N_6258);
and U8466 (N_8466,N_6973,N_7939);
and U8467 (N_8467,N_6740,N_6165);
xor U8468 (N_8468,N_7641,N_7622);
nand U8469 (N_8469,N_7508,N_7855);
or U8470 (N_8470,N_6943,N_7495);
nor U8471 (N_8471,N_6656,N_6461);
xnor U8472 (N_8472,N_6377,N_7592);
xnor U8473 (N_8473,N_6450,N_6507);
and U8474 (N_8474,N_6670,N_7678);
xnor U8475 (N_8475,N_7319,N_6911);
or U8476 (N_8476,N_7488,N_7005);
or U8477 (N_8477,N_7662,N_7539);
nand U8478 (N_8478,N_7282,N_6232);
nand U8479 (N_8479,N_6385,N_7010);
nand U8480 (N_8480,N_7067,N_6366);
nand U8481 (N_8481,N_6872,N_7050);
nand U8482 (N_8482,N_7420,N_7199);
or U8483 (N_8483,N_6583,N_7527);
nor U8484 (N_8484,N_6407,N_7745);
nor U8485 (N_8485,N_6953,N_7197);
nor U8486 (N_8486,N_7565,N_6800);
and U8487 (N_8487,N_7184,N_7957);
xnor U8488 (N_8488,N_6735,N_6962);
nand U8489 (N_8489,N_7882,N_7093);
nand U8490 (N_8490,N_6987,N_6489);
xor U8491 (N_8491,N_6094,N_7305);
nor U8492 (N_8492,N_7424,N_7607);
and U8493 (N_8493,N_6519,N_7457);
nor U8494 (N_8494,N_6928,N_6518);
or U8495 (N_8495,N_6697,N_7216);
nand U8496 (N_8496,N_7281,N_6535);
or U8497 (N_8497,N_6495,N_7234);
nand U8498 (N_8498,N_7945,N_7834);
nand U8499 (N_8499,N_7302,N_6959);
xnor U8500 (N_8500,N_6073,N_7949);
xor U8501 (N_8501,N_7721,N_6473);
xor U8502 (N_8502,N_6180,N_6485);
and U8503 (N_8503,N_7661,N_7274);
xnor U8504 (N_8504,N_6963,N_7823);
nand U8505 (N_8505,N_6947,N_6612);
nand U8506 (N_8506,N_6874,N_6734);
and U8507 (N_8507,N_6592,N_7869);
and U8508 (N_8508,N_6328,N_6862);
and U8509 (N_8509,N_6017,N_7525);
nor U8510 (N_8510,N_6418,N_7788);
and U8511 (N_8511,N_6773,N_7257);
or U8512 (N_8512,N_6768,N_6480);
xnor U8513 (N_8513,N_6076,N_6543);
nor U8514 (N_8514,N_6241,N_7561);
or U8515 (N_8515,N_6211,N_7943);
or U8516 (N_8516,N_6214,N_7912);
or U8517 (N_8517,N_7081,N_6923);
and U8518 (N_8518,N_7728,N_7842);
xor U8519 (N_8519,N_7701,N_7753);
and U8520 (N_8520,N_6830,N_6170);
and U8521 (N_8521,N_7200,N_7127);
and U8522 (N_8522,N_6251,N_7025);
and U8523 (N_8523,N_6604,N_7161);
nor U8524 (N_8524,N_7698,N_6775);
nor U8525 (N_8525,N_7703,N_6084);
nor U8526 (N_8526,N_6545,N_7128);
nor U8527 (N_8527,N_7817,N_6961);
or U8528 (N_8528,N_7951,N_7337);
or U8529 (N_8529,N_6227,N_6230);
or U8530 (N_8530,N_7250,N_7645);
and U8531 (N_8531,N_6264,N_6942);
nor U8532 (N_8532,N_6397,N_6127);
and U8533 (N_8533,N_6427,N_6470);
or U8534 (N_8534,N_7576,N_7376);
nor U8535 (N_8535,N_6279,N_7267);
nand U8536 (N_8536,N_6840,N_7750);
or U8537 (N_8537,N_7777,N_7237);
and U8538 (N_8538,N_6412,N_6936);
xor U8539 (N_8539,N_7911,N_6124);
or U8540 (N_8540,N_7767,N_6453);
or U8541 (N_8541,N_7825,N_7833);
or U8542 (N_8542,N_6243,N_7643);
nand U8543 (N_8543,N_6147,N_6991);
or U8544 (N_8544,N_6210,N_6858);
xor U8545 (N_8545,N_6710,N_7365);
nor U8546 (N_8546,N_7063,N_6520);
or U8547 (N_8547,N_7756,N_7815);
xnor U8548 (N_8548,N_6700,N_6909);
nand U8549 (N_8549,N_7387,N_6596);
and U8550 (N_8550,N_6382,N_7222);
nand U8551 (N_8551,N_7733,N_7811);
or U8552 (N_8552,N_6446,N_6464);
or U8553 (N_8553,N_7109,N_7306);
nor U8554 (N_8554,N_7905,N_7442);
or U8555 (N_8555,N_6245,N_6790);
xor U8556 (N_8556,N_6903,N_7889);
nand U8557 (N_8557,N_6927,N_6091);
xor U8558 (N_8558,N_7135,N_6647);
or U8559 (N_8559,N_6500,N_6665);
nor U8560 (N_8560,N_6192,N_6233);
or U8561 (N_8561,N_7697,N_7563);
nand U8562 (N_8562,N_6835,N_7361);
or U8563 (N_8563,N_6205,N_6378);
and U8564 (N_8564,N_7962,N_7595);
nor U8565 (N_8565,N_6783,N_6037);
and U8566 (N_8566,N_7963,N_6106);
nand U8567 (N_8567,N_6036,N_7391);
and U8568 (N_8568,N_7617,N_6185);
nand U8569 (N_8569,N_6589,N_7754);
nor U8570 (N_8570,N_6001,N_6870);
nor U8571 (N_8571,N_7272,N_7235);
or U8572 (N_8572,N_7629,N_6808);
or U8573 (N_8573,N_7151,N_7826);
or U8574 (N_8574,N_7298,N_6025);
xnor U8575 (N_8575,N_7427,N_6225);
nand U8576 (N_8576,N_6867,N_7637);
xor U8577 (N_8577,N_7173,N_6340);
nand U8578 (N_8578,N_7440,N_7801);
or U8579 (N_8579,N_7749,N_6371);
nand U8580 (N_8580,N_6536,N_7992);
and U8581 (N_8581,N_6945,N_7976);
or U8582 (N_8582,N_7047,N_7548);
xnor U8583 (N_8583,N_7584,N_7782);
and U8584 (N_8584,N_6420,N_7677);
nor U8585 (N_8585,N_7300,N_7021);
nor U8586 (N_8586,N_7832,N_7334);
nor U8587 (N_8587,N_7969,N_6876);
or U8588 (N_8588,N_6117,N_7472);
xnor U8589 (N_8589,N_7323,N_7954);
nor U8590 (N_8590,N_6068,N_7040);
nand U8591 (N_8591,N_7557,N_7359);
nand U8592 (N_8592,N_6333,N_7839);
nand U8593 (N_8593,N_6607,N_6242);
nor U8594 (N_8594,N_6921,N_7393);
xor U8595 (N_8595,N_7849,N_7212);
nand U8596 (N_8596,N_6078,N_7315);
nand U8597 (N_8597,N_7114,N_6514);
nor U8598 (N_8598,N_7471,N_7121);
or U8599 (N_8599,N_7147,N_6203);
nor U8600 (N_8600,N_7437,N_7188);
nor U8601 (N_8601,N_7054,N_6530);
nand U8602 (N_8602,N_7746,N_7850);
nor U8603 (N_8603,N_6417,N_6307);
and U8604 (N_8604,N_7140,N_7734);
or U8605 (N_8605,N_7001,N_6298);
nor U8606 (N_8606,N_6173,N_7900);
and U8607 (N_8607,N_7535,N_6999);
and U8608 (N_8608,N_7972,N_6523);
nor U8609 (N_8609,N_6789,N_7489);
nand U8610 (N_8610,N_7431,N_7967);
nor U8611 (N_8611,N_7781,N_6615);
xnor U8612 (N_8612,N_7304,N_6004);
nor U8613 (N_8613,N_7695,N_7864);
xor U8614 (N_8614,N_6365,N_7444);
nor U8615 (N_8615,N_6667,N_6269);
and U8616 (N_8616,N_6045,N_6686);
and U8617 (N_8617,N_6248,N_6988);
xnor U8618 (N_8618,N_6077,N_6350);
or U8619 (N_8619,N_6672,N_7886);
and U8620 (N_8620,N_6608,N_7906);
nor U8621 (N_8621,N_6434,N_6731);
nor U8622 (N_8622,N_7195,N_6109);
xor U8623 (N_8623,N_6946,N_7630);
and U8624 (N_8624,N_7018,N_6741);
and U8625 (N_8625,N_7353,N_7583);
and U8626 (N_8626,N_7086,N_6693);
nor U8627 (N_8627,N_6498,N_6455);
xnor U8628 (N_8628,N_7558,N_7329);
xnor U8629 (N_8629,N_7977,N_7898);
nor U8630 (N_8630,N_7394,N_7506);
nand U8631 (N_8631,N_7095,N_7586);
nand U8632 (N_8632,N_7205,N_7987);
nand U8633 (N_8633,N_6148,N_6584);
and U8634 (N_8634,N_7119,N_7529);
and U8635 (N_8635,N_6522,N_7342);
and U8636 (N_8636,N_6503,N_6012);
and U8637 (N_8637,N_7742,N_7975);
nand U8638 (N_8638,N_7153,N_6433);
and U8639 (N_8639,N_6319,N_7555);
nand U8640 (N_8640,N_7064,N_6509);
nor U8641 (N_8641,N_7513,N_7675);
xor U8642 (N_8642,N_7328,N_6290);
xor U8643 (N_8643,N_6484,N_6743);
or U8644 (N_8644,N_7398,N_7165);
or U8645 (N_8645,N_7606,N_7211);
or U8646 (N_8646,N_7418,N_7748);
and U8647 (N_8647,N_6846,N_6716);
or U8648 (N_8648,N_7255,N_6676);
or U8649 (N_8649,N_6727,N_7654);
xor U8650 (N_8650,N_6222,N_7554);
and U8651 (N_8651,N_6295,N_6197);
or U8652 (N_8652,N_6199,N_7443);
nand U8653 (N_8653,N_7412,N_6411);
nor U8654 (N_8654,N_7487,N_6088);
nor U8655 (N_8655,N_6762,N_7504);
and U8656 (N_8656,N_6847,N_7045);
xor U8657 (N_8657,N_7965,N_6614);
and U8658 (N_8658,N_6153,N_7020);
or U8659 (N_8659,N_7073,N_6765);
nand U8660 (N_8660,N_6595,N_7797);
xor U8661 (N_8661,N_7674,N_6479);
or U8662 (N_8662,N_6313,N_6476);
or U8663 (N_8663,N_7368,N_7390);
xor U8664 (N_8664,N_7719,N_7080);
or U8665 (N_8665,N_6019,N_6617);
nor U8666 (N_8666,N_7958,N_7265);
nand U8667 (N_8667,N_6440,N_7893);
xor U8668 (N_8668,N_6799,N_6586);
xor U8669 (N_8669,N_7542,N_7482);
nor U8670 (N_8670,N_6707,N_6228);
xnor U8671 (N_8671,N_6201,N_7546);
xnor U8672 (N_8672,N_7238,N_7470);
and U8673 (N_8673,N_6788,N_6416);
nand U8674 (N_8674,N_7891,N_6054);
nor U8675 (N_8675,N_7964,N_7800);
or U8676 (N_8676,N_7120,N_6478);
nand U8677 (N_8677,N_7843,N_6956);
xor U8678 (N_8678,N_6492,N_6761);
or U8679 (N_8679,N_6226,N_6571);
or U8680 (N_8680,N_7737,N_6646);
xor U8681 (N_8681,N_6413,N_6972);
xor U8682 (N_8682,N_6851,N_7572);
nor U8683 (N_8683,N_6823,N_7261);
and U8684 (N_8684,N_6794,N_7824);
or U8685 (N_8685,N_7925,N_7061);
nor U8686 (N_8686,N_6174,N_6655);
and U8687 (N_8687,N_6702,N_7077);
xor U8688 (N_8688,N_6375,N_6034);
nor U8689 (N_8689,N_6099,N_6206);
nand U8690 (N_8690,N_7011,N_6599);
xnor U8691 (N_8691,N_7009,N_7428);
nor U8692 (N_8692,N_6572,N_6853);
nor U8693 (N_8693,N_7189,N_6856);
xor U8694 (N_8694,N_7273,N_6011);
and U8695 (N_8695,N_6784,N_6939);
and U8696 (N_8696,N_7321,N_7058);
or U8697 (N_8697,N_7439,N_6803);
and U8698 (N_8698,N_7979,N_7921);
and U8699 (N_8699,N_6200,N_6564);
and U8700 (N_8700,N_7385,N_7168);
nand U8701 (N_8701,N_7757,N_6960);
or U8702 (N_8702,N_6252,N_6090);
nor U8703 (N_8703,N_7827,N_6540);
or U8704 (N_8704,N_6367,N_6190);
and U8705 (N_8705,N_7033,N_7164);
xor U8706 (N_8706,N_7819,N_6816);
nand U8707 (N_8707,N_6969,N_6452);
xor U8708 (N_8708,N_6691,N_6528);
nand U8709 (N_8709,N_7351,N_6029);
nand U8710 (N_8710,N_6103,N_7206);
xor U8711 (N_8711,N_6590,N_7284);
xor U8712 (N_8712,N_7183,N_7989);
xnor U8713 (N_8713,N_7633,N_7511);
nand U8714 (N_8714,N_7813,N_7400);
nand U8715 (N_8715,N_7389,N_6904);
xor U8716 (N_8716,N_6058,N_6129);
xnor U8717 (N_8717,N_6286,N_7451);
nor U8718 (N_8718,N_6221,N_7895);
xnor U8719 (N_8719,N_7688,N_6578);
nand U8720 (N_8720,N_6685,N_6352);
and U8721 (N_8721,N_7108,N_6268);
nand U8722 (N_8722,N_6860,N_6563);
and U8723 (N_8723,N_6998,N_6469);
and U8724 (N_8724,N_7579,N_6724);
xnor U8725 (N_8725,N_6737,N_6705);
xor U8726 (N_8726,N_6781,N_7318);
nor U8727 (N_8727,N_7955,N_6224);
nand U8728 (N_8728,N_6537,N_7316);
and U8729 (N_8729,N_7897,N_6318);
nand U8730 (N_8730,N_6348,N_7916);
nor U8731 (N_8731,N_7381,N_6753);
or U8732 (N_8732,N_7310,N_7241);
xnor U8733 (N_8733,N_6984,N_6042);
xnor U8734 (N_8734,N_6410,N_6644);
nor U8735 (N_8735,N_6558,N_7370);
or U8736 (N_8736,N_6032,N_7640);
and U8737 (N_8737,N_6938,N_7711);
nand U8738 (N_8738,N_7624,N_7847);
nor U8739 (N_8739,N_6133,N_6626);
nor U8740 (N_8740,N_6908,N_7268);
and U8741 (N_8741,N_7364,N_6666);
or U8742 (N_8742,N_6293,N_7333);
nand U8743 (N_8743,N_7611,N_6802);
nand U8744 (N_8744,N_6179,N_6403);
xor U8745 (N_8745,N_7226,N_7806);
nor U8746 (N_8746,N_7322,N_6263);
and U8747 (N_8747,N_7167,N_7392);
or U8748 (N_8748,N_7600,N_6096);
and U8749 (N_8749,N_6143,N_6772);
or U8750 (N_8750,N_7055,N_6620);
or U8751 (N_8751,N_6250,N_6910);
nor U8752 (N_8752,N_6562,N_7107);
nand U8753 (N_8753,N_6357,N_6580);
and U8754 (N_8754,N_6785,N_6283);
or U8755 (N_8755,N_7386,N_7534);
or U8756 (N_8756,N_6069,N_6490);
or U8757 (N_8757,N_7098,N_6683);
and U8758 (N_8758,N_7545,N_7415);
and U8759 (N_8759,N_6282,N_7331);
xnor U8760 (N_8760,N_6028,N_6326);
xor U8761 (N_8761,N_6849,N_6698);
xnor U8762 (N_8762,N_7598,N_7452);
xnor U8763 (N_8763,N_7014,N_7575);
nand U8764 (N_8764,N_6237,N_7293);
nand U8765 (N_8765,N_7336,N_6815);
xnor U8766 (N_8766,N_7613,N_6920);
nor U8767 (N_8767,N_6866,N_6404);
or U8768 (N_8768,N_7207,N_6386);
and U8769 (N_8769,N_6824,N_7605);
xor U8770 (N_8770,N_7104,N_7459);
or U8771 (N_8771,N_7035,N_6018);
nor U8772 (N_8772,N_7747,N_7798);
or U8773 (N_8773,N_6967,N_7899);
nor U8774 (N_8774,N_7520,N_6223);
nor U8775 (N_8775,N_7275,N_6878);
and U8776 (N_8776,N_6344,N_7049);
nand U8777 (N_8777,N_6792,N_6050);
nand U8778 (N_8778,N_6827,N_7138);
nor U8779 (N_8779,N_7718,N_7784);
and U8780 (N_8780,N_6142,N_7204);
and U8781 (N_8781,N_6733,N_6978);
and U8782 (N_8782,N_6955,N_6204);
and U8783 (N_8783,N_6906,N_7270);
nor U8784 (N_8784,N_7809,N_6839);
nand U8785 (N_8785,N_7345,N_6635);
or U8786 (N_8786,N_6437,N_6748);
or U8787 (N_8787,N_7338,N_6845);
xnor U8788 (N_8788,N_7523,N_7795);
or U8789 (N_8789,N_7295,N_7589);
xnor U8790 (N_8790,N_6677,N_6930);
or U8791 (N_8791,N_6544,N_7374);
nand U8792 (N_8792,N_7673,N_6031);
xor U8793 (N_8793,N_7469,N_7562);
xnor U8794 (N_8794,N_6188,N_7251);
and U8795 (N_8795,N_7259,N_6817);
or U8796 (N_8796,N_7830,N_6101);
or U8797 (N_8797,N_7134,N_6538);
nor U8798 (N_8798,N_6877,N_6428);
nor U8799 (N_8799,N_7665,N_6487);
nand U8800 (N_8800,N_6406,N_7658);
nor U8801 (N_8801,N_6841,N_7209);
and U8802 (N_8802,N_7845,N_7851);
nor U8803 (N_8803,N_6255,N_6850);
xnor U8804 (N_8804,N_6888,N_6673);
xnor U8805 (N_8805,N_6379,N_6539);
nor U8806 (N_8806,N_7985,N_7280);
nor U8807 (N_8807,N_6236,N_6300);
xor U8808 (N_8808,N_6436,N_6805);
nor U8809 (N_8809,N_7155,N_7036);
nor U8810 (N_8810,N_6426,N_7059);
xnor U8811 (N_8811,N_6119,N_6941);
nand U8812 (N_8812,N_6725,N_6178);
nand U8813 (N_8813,N_7787,N_7996);
nor U8814 (N_8814,N_6769,N_7299);
nand U8815 (N_8815,N_7516,N_7097);
nand U8816 (N_8816,N_6246,N_7399);
xor U8817 (N_8817,N_7139,N_7144);
or U8818 (N_8818,N_7017,N_7908);
nand U8819 (N_8819,N_6338,N_7564);
or U8820 (N_8820,N_7070,N_6896);
or U8821 (N_8821,N_6899,N_7597);
and U8822 (N_8822,N_6554,N_7743);
or U8823 (N_8823,N_7791,N_6852);
nand U8824 (N_8824,N_7594,N_7075);
nor U8825 (N_8825,N_6472,N_7290);
nand U8826 (N_8826,N_7549,N_7236);
and U8827 (N_8827,N_7278,N_7769);
nor U8828 (N_8828,N_7684,N_6948);
or U8829 (N_8829,N_6339,N_6010);
xor U8830 (N_8830,N_7271,N_6335);
or U8831 (N_8831,N_7526,N_6508);
and U8832 (N_8832,N_7078,N_6496);
or U8833 (N_8833,N_6425,N_6116);
nor U8834 (N_8834,N_6396,N_7685);
and U8835 (N_8835,N_7455,N_7034);
nand U8836 (N_8836,N_6308,N_6834);
and U8837 (N_8837,N_7129,N_6278);
xnor U8838 (N_8838,N_6254,N_6431);
nor U8839 (N_8839,N_7092,N_6573);
and U8840 (N_8840,N_6182,N_7182);
and U8841 (N_8841,N_6787,N_7498);
nor U8842 (N_8842,N_7030,N_7046);
and U8843 (N_8843,N_7296,N_6684);
nor U8844 (N_8844,N_7422,N_7016);
or U8845 (N_8845,N_6570,N_7664);
nand U8846 (N_8846,N_6569,N_7814);
or U8847 (N_8847,N_7264,N_6186);
or U8848 (N_8848,N_6722,N_6162);
nor U8849 (N_8849,N_6714,N_6641);
and U8850 (N_8850,N_7096,N_6907);
nor U8851 (N_8851,N_7551,N_6937);
and U8852 (N_8852,N_7580,N_7517);
nand U8853 (N_8853,N_6047,N_6126);
and U8854 (N_8854,N_6259,N_6115);
xor U8855 (N_8855,N_6060,N_7713);
nor U8856 (N_8856,N_7524,N_6869);
or U8857 (N_8857,N_6157,N_7541);
nor U8858 (N_8858,N_7566,N_7154);
nand U8859 (N_8859,N_6970,N_7536);
or U8860 (N_8860,N_7043,N_7314);
nor U8861 (N_8861,N_6392,N_7647);
xnor U8862 (N_8862,N_6952,N_6694);
xnor U8863 (N_8863,N_7460,N_7162);
nor U8864 (N_8864,N_7500,N_7804);
nand U8865 (N_8865,N_7436,N_7961);
nor U8866 (N_8866,N_6653,N_7360);
xor U8867 (N_8867,N_6606,N_7491);
nand U8868 (N_8868,N_7176,N_6388);
or U8869 (N_8869,N_7683,N_6779);
and U8870 (N_8870,N_6625,N_6880);
and U8871 (N_8871,N_6089,N_6577);
nor U8872 (N_8872,N_7947,N_6971);
nand U8873 (N_8873,N_6501,N_7326);
nor U8874 (N_8874,N_7481,N_6048);
or U8875 (N_8875,N_7741,N_7681);
xnor U8876 (N_8876,N_7219,N_6014);
or U8877 (N_8877,N_7110,N_6898);
or U8878 (N_8878,N_7702,N_6995);
nand U8879 (N_8879,N_6933,N_6471);
and U8880 (N_8880,N_7133,N_6239);
and U8881 (N_8881,N_6234,N_7352);
and U8882 (N_8882,N_7991,N_6585);
or U8883 (N_8883,N_7863,N_6916);
and U8884 (N_8884,N_7380,N_7247);
nor U8885 (N_8885,N_7946,N_6886);
nor U8886 (N_8886,N_7029,N_6194);
and U8887 (N_8887,N_7372,N_7990);
xnor U8888 (N_8888,N_7456,N_6966);
nor U8889 (N_8889,N_6568,N_7146);
nand U8890 (N_8890,N_7118,N_7642);
nor U8891 (N_8891,N_7382,N_6887);
xor U8892 (N_8892,N_6100,N_6331);
and U8893 (N_8893,N_6633,N_7836);
nor U8894 (N_8894,N_7335,N_7831);
and U8895 (N_8895,N_6093,N_7922);
nand U8896 (N_8896,N_7292,N_7015);
nor U8897 (N_8897,N_7423,N_7997);
nand U8898 (N_8898,N_6902,N_6912);
xnor U8899 (N_8899,N_7480,N_7537);
nand U8900 (N_8900,N_6659,N_7844);
nor U8901 (N_8901,N_7362,N_7599);
nor U8902 (N_8902,N_7037,N_6690);
or U8903 (N_8903,N_7632,N_7550);
nor U8904 (N_8904,N_6159,N_7231);
or U8905 (N_8905,N_6917,N_7325);
and U8906 (N_8906,N_6913,N_6638);
xor U8907 (N_8907,N_6021,N_7646);
nor U8908 (N_8908,N_7620,N_7820);
nand U8909 (N_8909,N_7547,N_7185);
nand U8910 (N_8910,N_6187,N_6738);
and U8911 (N_8911,N_6889,N_6317);
nand U8912 (N_8912,N_7051,N_7923);
nand U8913 (N_8913,N_7435,N_7783);
nand U8914 (N_8914,N_6717,N_7355);
or U8915 (N_8915,N_7332,N_7616);
nor U8916 (N_8916,N_7838,N_7971);
and U8917 (N_8917,N_7000,N_7375);
nand U8918 (N_8918,N_7694,N_7473);
xor U8919 (N_8919,N_6711,N_6516);
xnor U8920 (N_8920,N_6334,N_6588);
or U8921 (N_8921,N_6051,N_6859);
nor U8922 (N_8922,N_7569,N_6401);
and U8923 (N_8923,N_7768,N_6296);
xor U8924 (N_8924,N_6542,N_7930);
nand U8925 (N_8925,N_6797,N_7816);
nor U8926 (N_8926,N_7413,N_7623);
and U8927 (N_8927,N_7407,N_6422);
or U8928 (N_8928,N_6491,N_7676);
nand U8929 (N_8929,N_7141,N_6244);
nor U8930 (N_8930,N_6349,N_6663);
or U8931 (N_8931,N_6408,N_6754);
and U8932 (N_8932,N_7430,N_7085);
or U8933 (N_8933,N_6086,N_7904);
and U8934 (N_8934,N_7194,N_6351);
nand U8935 (N_8935,N_7312,N_7450);
xor U8936 (N_8936,N_6456,N_7710);
nand U8937 (N_8937,N_6689,N_7223);
xnor U8938 (N_8938,N_6726,N_7218);
xor U8939 (N_8939,N_7952,N_6949);
and U8940 (N_8940,N_6066,N_6982);
or U8941 (N_8941,N_6989,N_6145);
nor U8942 (N_8942,N_7560,N_7567);
and U8943 (N_8943,N_7056,N_7028);
nor U8944 (N_8944,N_7474,N_6547);
or U8945 (N_8945,N_7901,N_6310);
nand U8946 (N_8946,N_6770,N_6629);
nand U8947 (N_8947,N_7396,N_6688);
xnor U8948 (N_8948,N_6176,N_6652);
nand U8949 (N_8949,N_7910,N_7915);
or U8950 (N_8950,N_6309,N_6618);
nor U8951 (N_8951,N_7113,N_6504);
or U8952 (N_8952,N_6215,N_6306);
and U8953 (N_8953,N_7680,N_7032);
xnor U8954 (N_8954,N_6015,N_6027);
nand U8955 (N_8955,N_6486,N_6249);
and U8956 (N_8956,N_6531,N_7253);
nand U8957 (N_8957,N_6681,N_6284);
nor U8958 (N_8958,N_6445,N_7988);
or U8959 (N_8959,N_7125,N_6105);
and U8960 (N_8960,N_7712,N_6992);
xnor U8961 (N_8961,N_6502,N_6079);
and U8962 (N_8962,N_6448,N_7935);
nor U8963 (N_8963,N_7885,N_6958);
or U8964 (N_8964,N_6415,N_6008);
or U8965 (N_8965,N_7103,N_6372);
or U8966 (N_8966,N_6128,N_7052);
nor U8967 (N_8967,N_7682,N_6637);
and U8968 (N_8968,N_6634,N_7614);
nand U8969 (N_8969,N_7256,N_7246);
xnor U8970 (N_8970,N_6429,N_7942);
xnor U8971 (N_8971,N_6675,N_6882);
nand U8972 (N_8972,N_7066,N_6511);
and U8973 (N_8973,N_6466,N_6329);
and U8974 (N_8974,N_6643,N_7448);
or U8975 (N_8975,N_7724,N_7717);
and U8976 (N_8976,N_7603,N_6160);
and U8977 (N_8977,N_7521,N_7102);
nand U8978 (N_8978,N_7785,N_6409);
nand U8979 (N_8979,N_6441,N_6611);
xnor U8980 (N_8980,N_7765,N_7486);
or U8981 (N_8981,N_6155,N_7687);
and U8982 (N_8982,N_6925,N_7069);
nor U8983 (N_8983,N_7286,N_7124);
and U8984 (N_8984,N_7953,N_7950);
xnor U8985 (N_8985,N_7388,N_6482);
nand U8986 (N_8986,N_6030,N_7497);
and U8987 (N_8987,N_6682,N_6395);
nor U8988 (N_8988,N_7157,N_6374);
and U8989 (N_8989,N_6732,N_6900);
nor U8990 (N_8990,N_6715,N_7252);
and U8991 (N_8991,N_6394,N_6005);
xor U8992 (N_8992,N_7936,N_7934);
and U8993 (N_8993,N_6591,N_6067);
xnor U8994 (N_8994,N_6560,N_7433);
xor U8995 (N_8995,N_6838,N_7006);
xor U8996 (N_8996,N_7909,N_6064);
nand U8997 (N_8997,N_6703,N_7446);
nand U8998 (N_8998,N_7666,N_7865);
or U8999 (N_8999,N_7324,N_6261);
xor U9000 (N_9000,N_6416,N_7985);
xnor U9001 (N_9001,N_7857,N_7322);
nor U9002 (N_9002,N_6129,N_7580);
nand U9003 (N_9003,N_6717,N_6356);
and U9004 (N_9004,N_7993,N_7977);
nand U9005 (N_9005,N_6333,N_7054);
and U9006 (N_9006,N_7592,N_7737);
and U9007 (N_9007,N_7943,N_6503);
nand U9008 (N_9008,N_6550,N_7143);
nand U9009 (N_9009,N_7074,N_7963);
nand U9010 (N_9010,N_6763,N_6700);
xor U9011 (N_9011,N_6100,N_7504);
xor U9012 (N_9012,N_6503,N_7901);
nor U9013 (N_9013,N_6432,N_7342);
xnor U9014 (N_9014,N_7381,N_6718);
xnor U9015 (N_9015,N_7930,N_7961);
xnor U9016 (N_9016,N_6085,N_7833);
or U9017 (N_9017,N_6930,N_6668);
xor U9018 (N_9018,N_7882,N_7767);
xor U9019 (N_9019,N_7580,N_6344);
nor U9020 (N_9020,N_7173,N_6310);
or U9021 (N_9021,N_7081,N_7059);
or U9022 (N_9022,N_7528,N_6345);
or U9023 (N_9023,N_6224,N_7703);
and U9024 (N_9024,N_7821,N_6364);
or U9025 (N_9025,N_6710,N_7069);
nand U9026 (N_9026,N_7612,N_6355);
xnor U9027 (N_9027,N_7256,N_7546);
or U9028 (N_9028,N_7630,N_7322);
nand U9029 (N_9029,N_6743,N_7508);
and U9030 (N_9030,N_7328,N_7808);
nor U9031 (N_9031,N_6527,N_6890);
nor U9032 (N_9032,N_6396,N_7969);
nand U9033 (N_9033,N_7911,N_6055);
and U9034 (N_9034,N_6234,N_7322);
nor U9035 (N_9035,N_6019,N_7984);
nor U9036 (N_9036,N_7505,N_6620);
and U9037 (N_9037,N_6480,N_7978);
xnor U9038 (N_9038,N_6229,N_6497);
xnor U9039 (N_9039,N_7593,N_6269);
xnor U9040 (N_9040,N_6075,N_6214);
or U9041 (N_9041,N_7333,N_7779);
xor U9042 (N_9042,N_7623,N_6591);
nand U9043 (N_9043,N_7161,N_6005);
or U9044 (N_9044,N_7368,N_7708);
nor U9045 (N_9045,N_6168,N_7271);
nand U9046 (N_9046,N_6120,N_6445);
xnor U9047 (N_9047,N_7603,N_7061);
nand U9048 (N_9048,N_6355,N_6077);
nor U9049 (N_9049,N_7799,N_7444);
nor U9050 (N_9050,N_7224,N_7161);
and U9051 (N_9051,N_7041,N_7234);
nand U9052 (N_9052,N_7922,N_7498);
or U9053 (N_9053,N_7866,N_6888);
xor U9054 (N_9054,N_7130,N_7614);
or U9055 (N_9055,N_6554,N_6160);
nand U9056 (N_9056,N_6268,N_7812);
or U9057 (N_9057,N_7787,N_6692);
nand U9058 (N_9058,N_7140,N_6986);
and U9059 (N_9059,N_6169,N_6480);
or U9060 (N_9060,N_6881,N_7625);
xor U9061 (N_9061,N_6079,N_7033);
and U9062 (N_9062,N_7545,N_7617);
nor U9063 (N_9063,N_7241,N_7072);
nor U9064 (N_9064,N_7993,N_6238);
nor U9065 (N_9065,N_7140,N_7520);
and U9066 (N_9066,N_7288,N_7271);
nand U9067 (N_9067,N_7308,N_7948);
xor U9068 (N_9068,N_7784,N_6158);
and U9069 (N_9069,N_7968,N_7046);
or U9070 (N_9070,N_6755,N_6566);
nand U9071 (N_9071,N_6443,N_6598);
or U9072 (N_9072,N_6872,N_6896);
xor U9073 (N_9073,N_7047,N_7231);
xnor U9074 (N_9074,N_6755,N_6651);
or U9075 (N_9075,N_7737,N_6725);
xor U9076 (N_9076,N_7705,N_6324);
nor U9077 (N_9077,N_7986,N_7313);
nor U9078 (N_9078,N_6720,N_7958);
and U9079 (N_9079,N_6353,N_6446);
nor U9080 (N_9080,N_6264,N_6009);
nand U9081 (N_9081,N_7674,N_6310);
or U9082 (N_9082,N_7741,N_6055);
and U9083 (N_9083,N_6014,N_6566);
xnor U9084 (N_9084,N_7987,N_7570);
or U9085 (N_9085,N_6790,N_7703);
nor U9086 (N_9086,N_6875,N_7303);
nand U9087 (N_9087,N_7969,N_7985);
nand U9088 (N_9088,N_6979,N_7409);
or U9089 (N_9089,N_7971,N_7038);
nand U9090 (N_9090,N_6465,N_7475);
nor U9091 (N_9091,N_6652,N_7092);
nand U9092 (N_9092,N_6071,N_6770);
nand U9093 (N_9093,N_6492,N_6611);
and U9094 (N_9094,N_7451,N_6527);
nor U9095 (N_9095,N_6171,N_7547);
or U9096 (N_9096,N_7183,N_6606);
and U9097 (N_9097,N_7483,N_7485);
or U9098 (N_9098,N_6397,N_6937);
xor U9099 (N_9099,N_6193,N_7472);
xor U9100 (N_9100,N_7165,N_6191);
nand U9101 (N_9101,N_7480,N_7026);
or U9102 (N_9102,N_6679,N_6555);
nand U9103 (N_9103,N_6047,N_7089);
xor U9104 (N_9104,N_7435,N_6716);
xor U9105 (N_9105,N_7270,N_7119);
nand U9106 (N_9106,N_6666,N_7615);
nand U9107 (N_9107,N_7187,N_6836);
and U9108 (N_9108,N_7246,N_6996);
xnor U9109 (N_9109,N_7565,N_7646);
xnor U9110 (N_9110,N_6615,N_7510);
and U9111 (N_9111,N_7570,N_6774);
nor U9112 (N_9112,N_6556,N_6780);
or U9113 (N_9113,N_6655,N_7460);
nor U9114 (N_9114,N_7261,N_7809);
or U9115 (N_9115,N_7423,N_6044);
and U9116 (N_9116,N_6888,N_6510);
xnor U9117 (N_9117,N_7502,N_7188);
and U9118 (N_9118,N_6732,N_7641);
nor U9119 (N_9119,N_6252,N_7999);
xor U9120 (N_9120,N_6770,N_6033);
xnor U9121 (N_9121,N_6028,N_7697);
or U9122 (N_9122,N_6254,N_6839);
xnor U9123 (N_9123,N_7929,N_6370);
xor U9124 (N_9124,N_7793,N_6456);
nand U9125 (N_9125,N_7600,N_6856);
and U9126 (N_9126,N_6715,N_6997);
or U9127 (N_9127,N_6136,N_7775);
or U9128 (N_9128,N_7342,N_7979);
nand U9129 (N_9129,N_7417,N_6704);
nor U9130 (N_9130,N_7665,N_7404);
nand U9131 (N_9131,N_7041,N_6396);
or U9132 (N_9132,N_7347,N_6797);
nor U9133 (N_9133,N_6910,N_6899);
or U9134 (N_9134,N_7178,N_7823);
xnor U9135 (N_9135,N_6323,N_6451);
and U9136 (N_9136,N_6990,N_7794);
or U9137 (N_9137,N_7724,N_6400);
and U9138 (N_9138,N_7970,N_6926);
xor U9139 (N_9139,N_7645,N_7145);
xor U9140 (N_9140,N_6701,N_6955);
nor U9141 (N_9141,N_6598,N_6498);
nand U9142 (N_9142,N_6028,N_6439);
xor U9143 (N_9143,N_7438,N_7301);
and U9144 (N_9144,N_7773,N_7384);
or U9145 (N_9145,N_6605,N_7589);
xor U9146 (N_9146,N_7036,N_7051);
or U9147 (N_9147,N_7406,N_6628);
or U9148 (N_9148,N_7044,N_6226);
nor U9149 (N_9149,N_7719,N_7030);
or U9150 (N_9150,N_6721,N_7150);
nand U9151 (N_9151,N_7656,N_6541);
and U9152 (N_9152,N_7868,N_7307);
and U9153 (N_9153,N_7286,N_7864);
xnor U9154 (N_9154,N_7384,N_7047);
nor U9155 (N_9155,N_7964,N_7623);
and U9156 (N_9156,N_6282,N_7743);
nand U9157 (N_9157,N_6985,N_6079);
and U9158 (N_9158,N_6395,N_6524);
or U9159 (N_9159,N_7193,N_7558);
and U9160 (N_9160,N_7166,N_6620);
xor U9161 (N_9161,N_6539,N_7286);
or U9162 (N_9162,N_7869,N_6363);
xnor U9163 (N_9163,N_6901,N_7764);
xnor U9164 (N_9164,N_7466,N_6631);
xnor U9165 (N_9165,N_7371,N_6717);
and U9166 (N_9166,N_6868,N_6968);
nor U9167 (N_9167,N_6968,N_7511);
nand U9168 (N_9168,N_7683,N_6807);
nor U9169 (N_9169,N_7672,N_6251);
xor U9170 (N_9170,N_7200,N_6473);
nor U9171 (N_9171,N_6345,N_6637);
nand U9172 (N_9172,N_6588,N_6345);
and U9173 (N_9173,N_7654,N_6474);
xnor U9174 (N_9174,N_6812,N_7601);
nand U9175 (N_9175,N_6843,N_6533);
nor U9176 (N_9176,N_6695,N_7133);
nand U9177 (N_9177,N_6773,N_7253);
or U9178 (N_9178,N_6207,N_7458);
and U9179 (N_9179,N_7467,N_7968);
or U9180 (N_9180,N_6701,N_6611);
nand U9181 (N_9181,N_7717,N_7045);
nand U9182 (N_9182,N_7760,N_7523);
or U9183 (N_9183,N_7842,N_6718);
nor U9184 (N_9184,N_7202,N_7263);
or U9185 (N_9185,N_7463,N_6952);
nand U9186 (N_9186,N_7735,N_6826);
xnor U9187 (N_9187,N_6527,N_7226);
or U9188 (N_9188,N_7843,N_6369);
xor U9189 (N_9189,N_7418,N_6172);
xor U9190 (N_9190,N_7068,N_6288);
nand U9191 (N_9191,N_6193,N_7756);
xor U9192 (N_9192,N_7322,N_6974);
nor U9193 (N_9193,N_6765,N_7395);
nand U9194 (N_9194,N_7148,N_7998);
nor U9195 (N_9195,N_7108,N_6284);
and U9196 (N_9196,N_6873,N_7741);
or U9197 (N_9197,N_6214,N_7656);
nand U9198 (N_9198,N_6110,N_6211);
and U9199 (N_9199,N_7893,N_7477);
nand U9200 (N_9200,N_6991,N_7512);
nand U9201 (N_9201,N_6850,N_6101);
nor U9202 (N_9202,N_7740,N_7083);
nor U9203 (N_9203,N_6404,N_7262);
nand U9204 (N_9204,N_7750,N_6084);
or U9205 (N_9205,N_6292,N_7646);
xor U9206 (N_9206,N_6906,N_7966);
and U9207 (N_9207,N_6537,N_6356);
or U9208 (N_9208,N_6202,N_6126);
nand U9209 (N_9209,N_7272,N_7059);
xnor U9210 (N_9210,N_6881,N_6909);
or U9211 (N_9211,N_6591,N_7910);
xnor U9212 (N_9212,N_6995,N_7412);
nor U9213 (N_9213,N_6853,N_6622);
nor U9214 (N_9214,N_7349,N_7605);
nor U9215 (N_9215,N_6569,N_6660);
xnor U9216 (N_9216,N_6457,N_6916);
xor U9217 (N_9217,N_7401,N_6819);
nand U9218 (N_9218,N_7170,N_7776);
xnor U9219 (N_9219,N_7444,N_6818);
and U9220 (N_9220,N_6813,N_7486);
and U9221 (N_9221,N_7848,N_6816);
nand U9222 (N_9222,N_7432,N_6531);
nor U9223 (N_9223,N_6123,N_6140);
nand U9224 (N_9224,N_7667,N_6008);
nor U9225 (N_9225,N_7401,N_7627);
nand U9226 (N_9226,N_7987,N_6280);
nor U9227 (N_9227,N_7520,N_7895);
and U9228 (N_9228,N_6736,N_7722);
nand U9229 (N_9229,N_6374,N_7237);
and U9230 (N_9230,N_6955,N_7349);
nor U9231 (N_9231,N_7935,N_6337);
nor U9232 (N_9232,N_6130,N_6801);
or U9233 (N_9233,N_6833,N_7839);
nor U9234 (N_9234,N_7478,N_6356);
xor U9235 (N_9235,N_6750,N_7868);
and U9236 (N_9236,N_7614,N_7415);
or U9237 (N_9237,N_6783,N_7355);
nor U9238 (N_9238,N_7909,N_7734);
nand U9239 (N_9239,N_7715,N_6366);
and U9240 (N_9240,N_6257,N_7535);
nand U9241 (N_9241,N_7620,N_6610);
nor U9242 (N_9242,N_7228,N_6184);
nand U9243 (N_9243,N_6206,N_7751);
and U9244 (N_9244,N_6704,N_6626);
and U9245 (N_9245,N_6308,N_6963);
and U9246 (N_9246,N_6424,N_7132);
nand U9247 (N_9247,N_6677,N_7012);
or U9248 (N_9248,N_6148,N_7028);
xor U9249 (N_9249,N_6901,N_7700);
nand U9250 (N_9250,N_7430,N_6042);
or U9251 (N_9251,N_7612,N_6787);
nand U9252 (N_9252,N_6411,N_7481);
or U9253 (N_9253,N_6975,N_6516);
or U9254 (N_9254,N_7417,N_7329);
and U9255 (N_9255,N_7230,N_6354);
nand U9256 (N_9256,N_6435,N_6450);
xor U9257 (N_9257,N_6272,N_6800);
nor U9258 (N_9258,N_7094,N_7478);
or U9259 (N_9259,N_7459,N_6479);
xor U9260 (N_9260,N_7546,N_6389);
nand U9261 (N_9261,N_7170,N_6258);
nor U9262 (N_9262,N_6333,N_7537);
and U9263 (N_9263,N_6639,N_6983);
xnor U9264 (N_9264,N_7632,N_7717);
or U9265 (N_9265,N_6410,N_7447);
and U9266 (N_9266,N_6969,N_6267);
xor U9267 (N_9267,N_6877,N_6064);
or U9268 (N_9268,N_6725,N_6892);
or U9269 (N_9269,N_7491,N_6828);
or U9270 (N_9270,N_6394,N_7972);
xnor U9271 (N_9271,N_6519,N_6465);
nor U9272 (N_9272,N_7869,N_7086);
or U9273 (N_9273,N_7409,N_7924);
nand U9274 (N_9274,N_6997,N_6207);
nor U9275 (N_9275,N_7866,N_7376);
or U9276 (N_9276,N_7581,N_6175);
xor U9277 (N_9277,N_6432,N_7199);
xnor U9278 (N_9278,N_6198,N_7189);
and U9279 (N_9279,N_6105,N_7427);
nand U9280 (N_9280,N_6295,N_7637);
and U9281 (N_9281,N_7969,N_7895);
nand U9282 (N_9282,N_6608,N_7429);
xor U9283 (N_9283,N_7350,N_7267);
or U9284 (N_9284,N_6672,N_7918);
or U9285 (N_9285,N_7901,N_7421);
xor U9286 (N_9286,N_6832,N_6589);
nor U9287 (N_9287,N_6040,N_6334);
or U9288 (N_9288,N_7771,N_7685);
xor U9289 (N_9289,N_6381,N_7241);
xnor U9290 (N_9290,N_6769,N_7062);
or U9291 (N_9291,N_7771,N_7991);
nand U9292 (N_9292,N_6467,N_6223);
nand U9293 (N_9293,N_6850,N_7549);
and U9294 (N_9294,N_7326,N_7711);
nand U9295 (N_9295,N_7437,N_7021);
nor U9296 (N_9296,N_7814,N_7759);
xnor U9297 (N_9297,N_6485,N_6800);
xnor U9298 (N_9298,N_6541,N_6673);
nand U9299 (N_9299,N_7427,N_7135);
xor U9300 (N_9300,N_7848,N_7762);
nand U9301 (N_9301,N_7703,N_7742);
nor U9302 (N_9302,N_6641,N_6978);
or U9303 (N_9303,N_7679,N_6504);
or U9304 (N_9304,N_6919,N_6333);
xnor U9305 (N_9305,N_7805,N_6673);
or U9306 (N_9306,N_7861,N_7209);
or U9307 (N_9307,N_6766,N_7278);
nor U9308 (N_9308,N_7033,N_6639);
or U9309 (N_9309,N_6461,N_7640);
or U9310 (N_9310,N_6352,N_7705);
or U9311 (N_9311,N_7183,N_7074);
xor U9312 (N_9312,N_6881,N_7910);
nor U9313 (N_9313,N_7166,N_7685);
nor U9314 (N_9314,N_6004,N_6528);
or U9315 (N_9315,N_7377,N_6583);
and U9316 (N_9316,N_7481,N_7758);
nor U9317 (N_9317,N_6516,N_6031);
nand U9318 (N_9318,N_6088,N_7746);
nand U9319 (N_9319,N_6507,N_6425);
and U9320 (N_9320,N_7894,N_6773);
nand U9321 (N_9321,N_7199,N_7521);
nor U9322 (N_9322,N_6200,N_7534);
nand U9323 (N_9323,N_7891,N_7185);
xnor U9324 (N_9324,N_7773,N_7103);
nand U9325 (N_9325,N_6797,N_6862);
nand U9326 (N_9326,N_7198,N_6721);
nor U9327 (N_9327,N_7119,N_7859);
nor U9328 (N_9328,N_6045,N_6044);
and U9329 (N_9329,N_7482,N_7784);
and U9330 (N_9330,N_7142,N_7888);
nand U9331 (N_9331,N_7260,N_6194);
and U9332 (N_9332,N_6319,N_7538);
nor U9333 (N_9333,N_6690,N_6285);
nor U9334 (N_9334,N_6447,N_6182);
nor U9335 (N_9335,N_6827,N_7459);
or U9336 (N_9336,N_7014,N_6473);
nor U9337 (N_9337,N_6973,N_7707);
nor U9338 (N_9338,N_6224,N_7732);
nand U9339 (N_9339,N_7921,N_6560);
nand U9340 (N_9340,N_7821,N_6900);
or U9341 (N_9341,N_7677,N_7098);
or U9342 (N_9342,N_7890,N_6643);
and U9343 (N_9343,N_7718,N_7284);
or U9344 (N_9344,N_7112,N_6335);
nand U9345 (N_9345,N_6603,N_6055);
and U9346 (N_9346,N_6614,N_6508);
or U9347 (N_9347,N_6635,N_7689);
and U9348 (N_9348,N_6207,N_6363);
or U9349 (N_9349,N_6827,N_6285);
nor U9350 (N_9350,N_6162,N_7086);
and U9351 (N_9351,N_6582,N_7825);
xor U9352 (N_9352,N_7462,N_6111);
and U9353 (N_9353,N_7312,N_6195);
or U9354 (N_9354,N_7310,N_7464);
nand U9355 (N_9355,N_7740,N_7940);
nor U9356 (N_9356,N_6554,N_6985);
xnor U9357 (N_9357,N_6227,N_6908);
nor U9358 (N_9358,N_7277,N_6361);
nor U9359 (N_9359,N_6481,N_6674);
nand U9360 (N_9360,N_6512,N_7807);
xor U9361 (N_9361,N_6528,N_6593);
xor U9362 (N_9362,N_7064,N_6883);
or U9363 (N_9363,N_6526,N_7942);
nand U9364 (N_9364,N_6285,N_6281);
nand U9365 (N_9365,N_7836,N_7859);
nand U9366 (N_9366,N_6120,N_7240);
xor U9367 (N_9367,N_7959,N_6317);
nand U9368 (N_9368,N_6133,N_6004);
or U9369 (N_9369,N_7665,N_6958);
and U9370 (N_9370,N_7204,N_6395);
nand U9371 (N_9371,N_6254,N_7252);
or U9372 (N_9372,N_6740,N_7900);
and U9373 (N_9373,N_7101,N_7355);
xor U9374 (N_9374,N_6861,N_7334);
nor U9375 (N_9375,N_7025,N_7109);
nand U9376 (N_9376,N_7477,N_6914);
and U9377 (N_9377,N_6207,N_7782);
nand U9378 (N_9378,N_6629,N_6582);
nor U9379 (N_9379,N_6388,N_7161);
nor U9380 (N_9380,N_7350,N_6074);
nor U9381 (N_9381,N_6371,N_7674);
nand U9382 (N_9382,N_7368,N_7071);
or U9383 (N_9383,N_7705,N_6376);
nand U9384 (N_9384,N_6019,N_7287);
xnor U9385 (N_9385,N_7940,N_6610);
nand U9386 (N_9386,N_6529,N_6676);
or U9387 (N_9387,N_6040,N_6736);
nand U9388 (N_9388,N_7211,N_6254);
nor U9389 (N_9389,N_7530,N_7471);
xor U9390 (N_9390,N_6421,N_6841);
or U9391 (N_9391,N_7413,N_7783);
nor U9392 (N_9392,N_7770,N_6369);
and U9393 (N_9393,N_7496,N_6995);
or U9394 (N_9394,N_7583,N_7417);
xor U9395 (N_9395,N_6383,N_7939);
and U9396 (N_9396,N_7676,N_6182);
nand U9397 (N_9397,N_6238,N_6624);
nor U9398 (N_9398,N_6358,N_7721);
and U9399 (N_9399,N_6363,N_6508);
nand U9400 (N_9400,N_7492,N_7920);
or U9401 (N_9401,N_7700,N_7359);
and U9402 (N_9402,N_7569,N_7870);
nor U9403 (N_9403,N_7772,N_6726);
or U9404 (N_9404,N_7203,N_6829);
and U9405 (N_9405,N_7938,N_6151);
and U9406 (N_9406,N_7579,N_6663);
and U9407 (N_9407,N_7316,N_6617);
nor U9408 (N_9408,N_7046,N_6235);
xnor U9409 (N_9409,N_6345,N_6496);
and U9410 (N_9410,N_7709,N_6148);
nor U9411 (N_9411,N_7535,N_7574);
or U9412 (N_9412,N_7834,N_6841);
xnor U9413 (N_9413,N_6895,N_6694);
and U9414 (N_9414,N_7870,N_6729);
and U9415 (N_9415,N_6970,N_6610);
and U9416 (N_9416,N_6741,N_7385);
nor U9417 (N_9417,N_6923,N_7437);
nand U9418 (N_9418,N_6077,N_6931);
and U9419 (N_9419,N_7298,N_7571);
nand U9420 (N_9420,N_7325,N_6014);
and U9421 (N_9421,N_6648,N_7024);
nand U9422 (N_9422,N_6717,N_6108);
and U9423 (N_9423,N_6832,N_6229);
nand U9424 (N_9424,N_7352,N_6987);
nand U9425 (N_9425,N_6389,N_6280);
xor U9426 (N_9426,N_7948,N_6869);
or U9427 (N_9427,N_6235,N_6034);
and U9428 (N_9428,N_6578,N_7520);
xnor U9429 (N_9429,N_6202,N_6736);
and U9430 (N_9430,N_7115,N_6948);
nand U9431 (N_9431,N_7762,N_6168);
xor U9432 (N_9432,N_6399,N_7483);
nor U9433 (N_9433,N_6131,N_6463);
and U9434 (N_9434,N_6274,N_7272);
or U9435 (N_9435,N_6697,N_7773);
nand U9436 (N_9436,N_7911,N_6809);
nand U9437 (N_9437,N_6601,N_7291);
and U9438 (N_9438,N_7676,N_6870);
and U9439 (N_9439,N_7246,N_7688);
nand U9440 (N_9440,N_7693,N_6801);
nor U9441 (N_9441,N_6725,N_7877);
nor U9442 (N_9442,N_7003,N_7009);
or U9443 (N_9443,N_7964,N_6066);
and U9444 (N_9444,N_6262,N_6047);
and U9445 (N_9445,N_7534,N_7123);
or U9446 (N_9446,N_7898,N_6957);
xnor U9447 (N_9447,N_7514,N_7968);
nand U9448 (N_9448,N_7418,N_6004);
nor U9449 (N_9449,N_7201,N_7781);
nor U9450 (N_9450,N_7355,N_7089);
or U9451 (N_9451,N_7481,N_7747);
nand U9452 (N_9452,N_6373,N_7366);
xnor U9453 (N_9453,N_6698,N_7949);
nand U9454 (N_9454,N_7366,N_7899);
and U9455 (N_9455,N_7257,N_7488);
nand U9456 (N_9456,N_6970,N_6020);
nand U9457 (N_9457,N_7451,N_6300);
nand U9458 (N_9458,N_6670,N_7472);
nand U9459 (N_9459,N_7670,N_7736);
or U9460 (N_9460,N_7312,N_7552);
nor U9461 (N_9461,N_7863,N_7291);
and U9462 (N_9462,N_7504,N_6860);
or U9463 (N_9463,N_6784,N_7839);
or U9464 (N_9464,N_7954,N_6764);
and U9465 (N_9465,N_7930,N_6201);
or U9466 (N_9466,N_7161,N_6876);
xor U9467 (N_9467,N_7737,N_6708);
nor U9468 (N_9468,N_6923,N_7993);
xor U9469 (N_9469,N_7137,N_6574);
and U9470 (N_9470,N_7890,N_6713);
nand U9471 (N_9471,N_7367,N_6919);
and U9472 (N_9472,N_6227,N_6829);
or U9473 (N_9473,N_6610,N_7847);
nor U9474 (N_9474,N_6535,N_6943);
xnor U9475 (N_9475,N_7155,N_6558);
or U9476 (N_9476,N_6251,N_7592);
nor U9477 (N_9477,N_6241,N_7117);
and U9478 (N_9478,N_7273,N_6823);
xnor U9479 (N_9479,N_6111,N_6371);
nor U9480 (N_9480,N_6854,N_6586);
nor U9481 (N_9481,N_7481,N_7376);
nor U9482 (N_9482,N_7186,N_7457);
nand U9483 (N_9483,N_6542,N_6373);
nand U9484 (N_9484,N_7977,N_6698);
xor U9485 (N_9485,N_6849,N_7310);
xnor U9486 (N_9486,N_6189,N_7176);
or U9487 (N_9487,N_6646,N_7234);
xnor U9488 (N_9488,N_7286,N_6754);
xor U9489 (N_9489,N_7145,N_6174);
or U9490 (N_9490,N_6943,N_6920);
and U9491 (N_9491,N_7237,N_7447);
or U9492 (N_9492,N_6933,N_6160);
xnor U9493 (N_9493,N_7272,N_6523);
or U9494 (N_9494,N_6971,N_7158);
and U9495 (N_9495,N_6142,N_7665);
and U9496 (N_9496,N_6959,N_7030);
or U9497 (N_9497,N_6011,N_6353);
nor U9498 (N_9498,N_6222,N_7248);
nor U9499 (N_9499,N_6720,N_7918);
xnor U9500 (N_9500,N_7170,N_6902);
nand U9501 (N_9501,N_7936,N_6940);
nor U9502 (N_9502,N_6818,N_7112);
and U9503 (N_9503,N_6733,N_6970);
or U9504 (N_9504,N_7578,N_7305);
and U9505 (N_9505,N_7260,N_6283);
nand U9506 (N_9506,N_7120,N_7794);
and U9507 (N_9507,N_7375,N_7305);
and U9508 (N_9508,N_7213,N_6448);
nand U9509 (N_9509,N_6590,N_7694);
nand U9510 (N_9510,N_6729,N_7463);
nand U9511 (N_9511,N_7512,N_7639);
xor U9512 (N_9512,N_7237,N_7441);
and U9513 (N_9513,N_6480,N_6628);
and U9514 (N_9514,N_6219,N_6665);
and U9515 (N_9515,N_6391,N_7230);
and U9516 (N_9516,N_7602,N_6272);
and U9517 (N_9517,N_7524,N_7313);
nand U9518 (N_9518,N_6165,N_6489);
and U9519 (N_9519,N_7638,N_7199);
xor U9520 (N_9520,N_6811,N_6880);
and U9521 (N_9521,N_7056,N_7978);
or U9522 (N_9522,N_7077,N_6783);
xnor U9523 (N_9523,N_6926,N_6159);
nor U9524 (N_9524,N_6145,N_7472);
xor U9525 (N_9525,N_6010,N_6303);
xnor U9526 (N_9526,N_7756,N_7343);
or U9527 (N_9527,N_6325,N_6907);
nand U9528 (N_9528,N_6238,N_6430);
nor U9529 (N_9529,N_6692,N_6975);
nor U9530 (N_9530,N_6005,N_6955);
nor U9531 (N_9531,N_7520,N_6108);
or U9532 (N_9532,N_6897,N_6159);
xnor U9533 (N_9533,N_6475,N_6719);
or U9534 (N_9534,N_6775,N_6155);
and U9535 (N_9535,N_7112,N_6734);
nand U9536 (N_9536,N_6013,N_7516);
or U9537 (N_9537,N_6280,N_7410);
or U9538 (N_9538,N_6847,N_7300);
or U9539 (N_9539,N_6355,N_6646);
or U9540 (N_9540,N_6402,N_7814);
nor U9541 (N_9541,N_7249,N_7778);
xnor U9542 (N_9542,N_7139,N_7168);
xor U9543 (N_9543,N_6672,N_6799);
or U9544 (N_9544,N_6403,N_7474);
nor U9545 (N_9545,N_7017,N_6587);
nand U9546 (N_9546,N_7260,N_6895);
or U9547 (N_9547,N_6936,N_6067);
or U9548 (N_9548,N_7956,N_6243);
xnor U9549 (N_9549,N_6352,N_7550);
or U9550 (N_9550,N_6986,N_7200);
nor U9551 (N_9551,N_7695,N_6768);
nor U9552 (N_9552,N_7413,N_6859);
xor U9553 (N_9553,N_6627,N_7379);
nand U9554 (N_9554,N_7975,N_7837);
nor U9555 (N_9555,N_6369,N_7923);
or U9556 (N_9556,N_6723,N_6655);
nor U9557 (N_9557,N_6111,N_7416);
nor U9558 (N_9558,N_7430,N_6737);
and U9559 (N_9559,N_7424,N_6841);
or U9560 (N_9560,N_7228,N_7545);
nand U9561 (N_9561,N_7750,N_6221);
xor U9562 (N_9562,N_7023,N_7806);
or U9563 (N_9563,N_6945,N_7909);
or U9564 (N_9564,N_6834,N_6858);
nand U9565 (N_9565,N_6069,N_6886);
xor U9566 (N_9566,N_6399,N_7262);
nand U9567 (N_9567,N_7568,N_6983);
or U9568 (N_9568,N_6572,N_6807);
nand U9569 (N_9569,N_7654,N_7980);
xnor U9570 (N_9570,N_6379,N_7264);
nor U9571 (N_9571,N_7016,N_7866);
or U9572 (N_9572,N_7814,N_7741);
xor U9573 (N_9573,N_6131,N_6748);
xor U9574 (N_9574,N_6228,N_6765);
nor U9575 (N_9575,N_7620,N_7034);
and U9576 (N_9576,N_6862,N_6702);
xnor U9577 (N_9577,N_7598,N_6814);
and U9578 (N_9578,N_7307,N_7520);
xnor U9579 (N_9579,N_6073,N_6172);
nor U9580 (N_9580,N_7675,N_7219);
and U9581 (N_9581,N_7264,N_7712);
nor U9582 (N_9582,N_7282,N_6784);
and U9583 (N_9583,N_7904,N_7734);
and U9584 (N_9584,N_6890,N_7446);
or U9585 (N_9585,N_7048,N_7698);
and U9586 (N_9586,N_7335,N_7365);
or U9587 (N_9587,N_6516,N_7276);
or U9588 (N_9588,N_7420,N_6298);
nand U9589 (N_9589,N_7871,N_7653);
or U9590 (N_9590,N_6003,N_6423);
and U9591 (N_9591,N_7719,N_6637);
or U9592 (N_9592,N_6359,N_7305);
nor U9593 (N_9593,N_7828,N_6193);
xnor U9594 (N_9594,N_7897,N_7744);
nor U9595 (N_9595,N_7676,N_6657);
nand U9596 (N_9596,N_6944,N_7496);
nor U9597 (N_9597,N_6260,N_6859);
nand U9598 (N_9598,N_7321,N_7952);
nor U9599 (N_9599,N_6147,N_6568);
nor U9600 (N_9600,N_6757,N_7325);
nand U9601 (N_9601,N_7406,N_6571);
xnor U9602 (N_9602,N_7101,N_7333);
nor U9603 (N_9603,N_7318,N_7677);
or U9604 (N_9604,N_6099,N_7967);
nor U9605 (N_9605,N_7206,N_7566);
or U9606 (N_9606,N_7526,N_7433);
xor U9607 (N_9607,N_6207,N_7727);
xor U9608 (N_9608,N_7998,N_7783);
xor U9609 (N_9609,N_7625,N_7028);
and U9610 (N_9610,N_6853,N_6337);
xor U9611 (N_9611,N_6466,N_7071);
nand U9612 (N_9612,N_7147,N_6608);
and U9613 (N_9613,N_6930,N_7491);
or U9614 (N_9614,N_6964,N_6726);
nand U9615 (N_9615,N_6377,N_6022);
and U9616 (N_9616,N_6874,N_6146);
and U9617 (N_9617,N_6249,N_7673);
or U9618 (N_9618,N_7920,N_6689);
and U9619 (N_9619,N_7538,N_6673);
and U9620 (N_9620,N_6479,N_7871);
nor U9621 (N_9621,N_6682,N_6691);
nand U9622 (N_9622,N_7126,N_6522);
nor U9623 (N_9623,N_6305,N_7147);
and U9624 (N_9624,N_6970,N_7912);
nor U9625 (N_9625,N_7855,N_7003);
xor U9626 (N_9626,N_6071,N_6157);
nor U9627 (N_9627,N_7077,N_7232);
or U9628 (N_9628,N_7289,N_7391);
xnor U9629 (N_9629,N_7073,N_7569);
nand U9630 (N_9630,N_6495,N_6241);
nand U9631 (N_9631,N_6868,N_6755);
or U9632 (N_9632,N_7872,N_6338);
or U9633 (N_9633,N_7817,N_7929);
or U9634 (N_9634,N_6985,N_7359);
nand U9635 (N_9635,N_6668,N_7461);
or U9636 (N_9636,N_6430,N_7773);
nand U9637 (N_9637,N_6144,N_6875);
or U9638 (N_9638,N_6055,N_6217);
and U9639 (N_9639,N_7256,N_6950);
xnor U9640 (N_9640,N_6298,N_7241);
nor U9641 (N_9641,N_7166,N_7212);
nor U9642 (N_9642,N_7733,N_6683);
and U9643 (N_9643,N_6286,N_6771);
xnor U9644 (N_9644,N_6465,N_7254);
xor U9645 (N_9645,N_6526,N_6763);
nand U9646 (N_9646,N_6102,N_6965);
or U9647 (N_9647,N_7256,N_6227);
xnor U9648 (N_9648,N_7696,N_6571);
nand U9649 (N_9649,N_6330,N_6176);
nor U9650 (N_9650,N_7878,N_7236);
and U9651 (N_9651,N_6263,N_6331);
or U9652 (N_9652,N_7442,N_6934);
or U9653 (N_9653,N_6682,N_6741);
xor U9654 (N_9654,N_7401,N_6213);
or U9655 (N_9655,N_6636,N_6401);
nand U9656 (N_9656,N_6911,N_6190);
nor U9657 (N_9657,N_6055,N_7124);
xor U9658 (N_9658,N_6665,N_7361);
nand U9659 (N_9659,N_7740,N_7338);
nor U9660 (N_9660,N_6587,N_6139);
and U9661 (N_9661,N_6365,N_6236);
or U9662 (N_9662,N_7070,N_7776);
or U9663 (N_9663,N_6911,N_6703);
and U9664 (N_9664,N_7660,N_7560);
or U9665 (N_9665,N_7230,N_6637);
or U9666 (N_9666,N_7158,N_6400);
or U9667 (N_9667,N_6277,N_7504);
nor U9668 (N_9668,N_7724,N_7046);
or U9669 (N_9669,N_7968,N_6948);
and U9670 (N_9670,N_7525,N_6601);
nor U9671 (N_9671,N_6078,N_6060);
nand U9672 (N_9672,N_6776,N_7870);
nand U9673 (N_9673,N_7680,N_6132);
nand U9674 (N_9674,N_7424,N_7492);
xnor U9675 (N_9675,N_7778,N_7070);
and U9676 (N_9676,N_6442,N_6256);
nor U9677 (N_9677,N_6015,N_7717);
and U9678 (N_9678,N_7394,N_6827);
and U9679 (N_9679,N_6610,N_7989);
or U9680 (N_9680,N_7886,N_6275);
xnor U9681 (N_9681,N_7354,N_7326);
or U9682 (N_9682,N_7433,N_7670);
nand U9683 (N_9683,N_6086,N_6340);
nor U9684 (N_9684,N_6495,N_6568);
nor U9685 (N_9685,N_7892,N_6070);
nor U9686 (N_9686,N_7508,N_6801);
nor U9687 (N_9687,N_7820,N_7092);
nand U9688 (N_9688,N_6677,N_6620);
nor U9689 (N_9689,N_7111,N_7833);
nand U9690 (N_9690,N_6551,N_6694);
xor U9691 (N_9691,N_6290,N_7530);
and U9692 (N_9692,N_7025,N_6943);
and U9693 (N_9693,N_7763,N_7478);
nor U9694 (N_9694,N_7305,N_6460);
nand U9695 (N_9695,N_7471,N_7993);
or U9696 (N_9696,N_7264,N_7705);
or U9697 (N_9697,N_6400,N_6473);
xor U9698 (N_9698,N_6150,N_6649);
and U9699 (N_9699,N_6971,N_7503);
and U9700 (N_9700,N_7410,N_7946);
xnor U9701 (N_9701,N_6359,N_7873);
nand U9702 (N_9702,N_7155,N_7487);
or U9703 (N_9703,N_6083,N_7181);
xor U9704 (N_9704,N_6222,N_6023);
and U9705 (N_9705,N_7730,N_7953);
and U9706 (N_9706,N_6082,N_6211);
or U9707 (N_9707,N_7220,N_6261);
nand U9708 (N_9708,N_7677,N_7459);
nor U9709 (N_9709,N_7114,N_6221);
or U9710 (N_9710,N_7201,N_6674);
and U9711 (N_9711,N_6931,N_6779);
and U9712 (N_9712,N_6688,N_6306);
or U9713 (N_9713,N_7642,N_7516);
or U9714 (N_9714,N_6256,N_6081);
xor U9715 (N_9715,N_6308,N_7936);
xnor U9716 (N_9716,N_7263,N_7560);
xor U9717 (N_9717,N_6235,N_6038);
nand U9718 (N_9718,N_7291,N_6147);
and U9719 (N_9719,N_7723,N_7182);
xor U9720 (N_9720,N_6838,N_7965);
nor U9721 (N_9721,N_7758,N_6735);
nand U9722 (N_9722,N_6710,N_6281);
xor U9723 (N_9723,N_7257,N_7712);
nor U9724 (N_9724,N_6278,N_6833);
nand U9725 (N_9725,N_6525,N_7730);
nand U9726 (N_9726,N_7555,N_6339);
xnor U9727 (N_9727,N_7222,N_7384);
or U9728 (N_9728,N_6765,N_6075);
and U9729 (N_9729,N_7852,N_6067);
xor U9730 (N_9730,N_6608,N_6417);
and U9731 (N_9731,N_7991,N_6033);
and U9732 (N_9732,N_6671,N_7242);
nor U9733 (N_9733,N_6961,N_7566);
nand U9734 (N_9734,N_6631,N_6903);
or U9735 (N_9735,N_7405,N_7914);
nor U9736 (N_9736,N_6494,N_6741);
nor U9737 (N_9737,N_6773,N_7666);
xor U9738 (N_9738,N_7638,N_6945);
and U9739 (N_9739,N_6905,N_6640);
nand U9740 (N_9740,N_6160,N_6118);
xnor U9741 (N_9741,N_7823,N_6236);
and U9742 (N_9742,N_7824,N_7778);
and U9743 (N_9743,N_6529,N_6282);
and U9744 (N_9744,N_7808,N_7931);
xor U9745 (N_9745,N_7845,N_7646);
or U9746 (N_9746,N_6839,N_6043);
and U9747 (N_9747,N_7998,N_7795);
or U9748 (N_9748,N_7379,N_7841);
or U9749 (N_9749,N_7176,N_7984);
nand U9750 (N_9750,N_7090,N_6160);
or U9751 (N_9751,N_7115,N_6195);
xnor U9752 (N_9752,N_6036,N_7189);
nor U9753 (N_9753,N_7551,N_7502);
and U9754 (N_9754,N_7744,N_7851);
nand U9755 (N_9755,N_6017,N_6818);
xor U9756 (N_9756,N_6718,N_6429);
and U9757 (N_9757,N_7989,N_7998);
or U9758 (N_9758,N_6085,N_7057);
xor U9759 (N_9759,N_6233,N_7064);
xor U9760 (N_9760,N_7219,N_7365);
nand U9761 (N_9761,N_6639,N_7872);
or U9762 (N_9762,N_6522,N_6231);
or U9763 (N_9763,N_6695,N_6740);
xor U9764 (N_9764,N_7108,N_6110);
nor U9765 (N_9765,N_6929,N_7696);
nor U9766 (N_9766,N_6585,N_6560);
nor U9767 (N_9767,N_6981,N_7203);
or U9768 (N_9768,N_7447,N_7706);
or U9769 (N_9769,N_6347,N_7485);
nand U9770 (N_9770,N_7269,N_7659);
or U9771 (N_9771,N_7088,N_6781);
nand U9772 (N_9772,N_6332,N_7824);
xor U9773 (N_9773,N_6548,N_6993);
nor U9774 (N_9774,N_7996,N_7647);
and U9775 (N_9775,N_7798,N_6882);
nor U9776 (N_9776,N_7229,N_6046);
nand U9777 (N_9777,N_7579,N_6683);
xor U9778 (N_9778,N_6377,N_6781);
nor U9779 (N_9779,N_6933,N_7213);
and U9780 (N_9780,N_6135,N_6196);
nor U9781 (N_9781,N_7093,N_6412);
xor U9782 (N_9782,N_6334,N_6933);
and U9783 (N_9783,N_7754,N_6097);
or U9784 (N_9784,N_7138,N_7569);
and U9785 (N_9785,N_6523,N_6212);
nor U9786 (N_9786,N_6268,N_7702);
and U9787 (N_9787,N_6358,N_7402);
nor U9788 (N_9788,N_7125,N_6595);
nand U9789 (N_9789,N_7970,N_6249);
xnor U9790 (N_9790,N_6285,N_7974);
or U9791 (N_9791,N_7190,N_7446);
or U9792 (N_9792,N_7417,N_6955);
nand U9793 (N_9793,N_7319,N_6113);
or U9794 (N_9794,N_7543,N_6062);
nor U9795 (N_9795,N_7812,N_6582);
nand U9796 (N_9796,N_6317,N_6343);
xor U9797 (N_9797,N_7351,N_6242);
and U9798 (N_9798,N_6968,N_6698);
or U9799 (N_9799,N_6865,N_6928);
or U9800 (N_9800,N_7057,N_6042);
xor U9801 (N_9801,N_6450,N_6023);
or U9802 (N_9802,N_7094,N_6608);
nand U9803 (N_9803,N_6748,N_6962);
or U9804 (N_9804,N_7666,N_6481);
and U9805 (N_9805,N_6984,N_7079);
nor U9806 (N_9806,N_7651,N_6686);
xnor U9807 (N_9807,N_6465,N_7161);
nor U9808 (N_9808,N_6322,N_6235);
xor U9809 (N_9809,N_6531,N_6103);
and U9810 (N_9810,N_7719,N_7999);
nor U9811 (N_9811,N_7477,N_7564);
nor U9812 (N_9812,N_6741,N_7520);
xnor U9813 (N_9813,N_6810,N_7196);
nor U9814 (N_9814,N_6737,N_7297);
xor U9815 (N_9815,N_7203,N_7598);
or U9816 (N_9816,N_7118,N_6166);
nand U9817 (N_9817,N_7508,N_7698);
and U9818 (N_9818,N_7010,N_6701);
nor U9819 (N_9819,N_6836,N_6110);
nand U9820 (N_9820,N_7733,N_7211);
nor U9821 (N_9821,N_6069,N_6047);
nand U9822 (N_9822,N_7268,N_6683);
nand U9823 (N_9823,N_7272,N_6915);
nand U9824 (N_9824,N_6645,N_7700);
and U9825 (N_9825,N_7818,N_6524);
and U9826 (N_9826,N_6067,N_7401);
and U9827 (N_9827,N_6211,N_6216);
xor U9828 (N_9828,N_7819,N_6066);
xnor U9829 (N_9829,N_6374,N_6160);
or U9830 (N_9830,N_7642,N_6109);
xor U9831 (N_9831,N_7784,N_6510);
nand U9832 (N_9832,N_7960,N_7477);
xor U9833 (N_9833,N_6030,N_7289);
nor U9834 (N_9834,N_7793,N_6149);
xor U9835 (N_9835,N_7421,N_6472);
or U9836 (N_9836,N_7114,N_7942);
or U9837 (N_9837,N_6239,N_6245);
nand U9838 (N_9838,N_6071,N_7065);
and U9839 (N_9839,N_6027,N_7481);
nand U9840 (N_9840,N_6231,N_6384);
or U9841 (N_9841,N_7003,N_6626);
nor U9842 (N_9842,N_7009,N_7609);
nor U9843 (N_9843,N_7270,N_6815);
and U9844 (N_9844,N_6649,N_6910);
xnor U9845 (N_9845,N_6777,N_7397);
nor U9846 (N_9846,N_7584,N_7327);
and U9847 (N_9847,N_6539,N_6544);
or U9848 (N_9848,N_6499,N_7310);
xor U9849 (N_9849,N_6979,N_6470);
nor U9850 (N_9850,N_7037,N_6440);
xnor U9851 (N_9851,N_6581,N_6975);
or U9852 (N_9852,N_6294,N_7476);
or U9853 (N_9853,N_6480,N_6244);
and U9854 (N_9854,N_6635,N_7372);
xnor U9855 (N_9855,N_6815,N_7660);
xor U9856 (N_9856,N_7053,N_6958);
xnor U9857 (N_9857,N_7027,N_6844);
xor U9858 (N_9858,N_6628,N_6546);
or U9859 (N_9859,N_7768,N_7432);
or U9860 (N_9860,N_7425,N_7950);
nand U9861 (N_9861,N_7402,N_6176);
xor U9862 (N_9862,N_6969,N_7783);
nor U9863 (N_9863,N_6306,N_6478);
nand U9864 (N_9864,N_7572,N_6241);
nand U9865 (N_9865,N_7371,N_7508);
xor U9866 (N_9866,N_7841,N_7709);
xnor U9867 (N_9867,N_6453,N_6064);
nor U9868 (N_9868,N_7791,N_6830);
nand U9869 (N_9869,N_7222,N_7438);
nand U9870 (N_9870,N_7628,N_7861);
nand U9871 (N_9871,N_7476,N_7536);
nand U9872 (N_9872,N_7068,N_7646);
xor U9873 (N_9873,N_6328,N_7070);
or U9874 (N_9874,N_7472,N_6969);
nand U9875 (N_9875,N_7224,N_7555);
or U9876 (N_9876,N_6627,N_6082);
nor U9877 (N_9877,N_6347,N_6395);
and U9878 (N_9878,N_6291,N_7761);
nor U9879 (N_9879,N_6104,N_6569);
nand U9880 (N_9880,N_7040,N_6382);
xnor U9881 (N_9881,N_7598,N_7509);
xor U9882 (N_9882,N_7107,N_7455);
nand U9883 (N_9883,N_7516,N_7961);
nand U9884 (N_9884,N_7302,N_7044);
xor U9885 (N_9885,N_7728,N_7122);
and U9886 (N_9886,N_6199,N_7831);
nand U9887 (N_9887,N_6614,N_7555);
nand U9888 (N_9888,N_7769,N_6797);
and U9889 (N_9889,N_7418,N_6477);
xnor U9890 (N_9890,N_7074,N_6003);
nand U9891 (N_9891,N_7628,N_7587);
or U9892 (N_9892,N_7867,N_6945);
nand U9893 (N_9893,N_6924,N_7042);
or U9894 (N_9894,N_6579,N_6269);
or U9895 (N_9895,N_7222,N_7591);
nor U9896 (N_9896,N_7762,N_6653);
nor U9897 (N_9897,N_7111,N_6158);
nor U9898 (N_9898,N_6362,N_6566);
and U9899 (N_9899,N_6989,N_6831);
nand U9900 (N_9900,N_7318,N_6731);
nand U9901 (N_9901,N_7812,N_7953);
or U9902 (N_9902,N_6537,N_6501);
xor U9903 (N_9903,N_7091,N_6942);
and U9904 (N_9904,N_7400,N_7295);
xnor U9905 (N_9905,N_6135,N_6030);
and U9906 (N_9906,N_7885,N_6524);
nand U9907 (N_9907,N_7102,N_6622);
nand U9908 (N_9908,N_7973,N_6039);
xor U9909 (N_9909,N_7344,N_6293);
and U9910 (N_9910,N_7145,N_6491);
or U9911 (N_9911,N_7820,N_6600);
nand U9912 (N_9912,N_6650,N_7124);
nor U9913 (N_9913,N_6039,N_6511);
nand U9914 (N_9914,N_6006,N_7634);
nand U9915 (N_9915,N_6947,N_6627);
and U9916 (N_9916,N_6064,N_6297);
nor U9917 (N_9917,N_7617,N_7309);
or U9918 (N_9918,N_6782,N_6594);
nand U9919 (N_9919,N_6281,N_6887);
nor U9920 (N_9920,N_6809,N_6186);
and U9921 (N_9921,N_6586,N_6379);
or U9922 (N_9922,N_7662,N_7791);
nor U9923 (N_9923,N_6690,N_7462);
nor U9924 (N_9924,N_6465,N_6228);
and U9925 (N_9925,N_6803,N_7722);
or U9926 (N_9926,N_7965,N_6319);
and U9927 (N_9927,N_6040,N_7192);
or U9928 (N_9928,N_6727,N_7041);
nor U9929 (N_9929,N_6347,N_6255);
nor U9930 (N_9930,N_6498,N_6055);
or U9931 (N_9931,N_7937,N_7842);
nor U9932 (N_9932,N_6201,N_7731);
nor U9933 (N_9933,N_7688,N_6963);
and U9934 (N_9934,N_6993,N_7630);
nand U9935 (N_9935,N_6425,N_6560);
or U9936 (N_9936,N_7514,N_7157);
and U9937 (N_9937,N_7206,N_7195);
or U9938 (N_9938,N_7014,N_6928);
or U9939 (N_9939,N_7991,N_6799);
or U9940 (N_9940,N_7112,N_7200);
or U9941 (N_9941,N_6646,N_7464);
and U9942 (N_9942,N_6653,N_7154);
nand U9943 (N_9943,N_7535,N_7105);
and U9944 (N_9944,N_6755,N_6025);
and U9945 (N_9945,N_6740,N_7353);
nand U9946 (N_9946,N_6098,N_6535);
nor U9947 (N_9947,N_6277,N_7150);
or U9948 (N_9948,N_6045,N_7334);
or U9949 (N_9949,N_6379,N_6038);
nor U9950 (N_9950,N_7428,N_6928);
nand U9951 (N_9951,N_7274,N_6579);
nor U9952 (N_9952,N_7364,N_6261);
or U9953 (N_9953,N_7043,N_6344);
nand U9954 (N_9954,N_7324,N_6503);
nor U9955 (N_9955,N_6545,N_7312);
and U9956 (N_9956,N_7577,N_7535);
or U9957 (N_9957,N_7385,N_7683);
nor U9958 (N_9958,N_7550,N_7102);
and U9959 (N_9959,N_7930,N_6847);
xor U9960 (N_9960,N_7145,N_6639);
or U9961 (N_9961,N_7916,N_7866);
or U9962 (N_9962,N_6110,N_7603);
nor U9963 (N_9963,N_7611,N_7357);
xnor U9964 (N_9964,N_6631,N_6832);
nand U9965 (N_9965,N_7398,N_6563);
nand U9966 (N_9966,N_6760,N_7596);
nand U9967 (N_9967,N_7521,N_6395);
or U9968 (N_9968,N_6723,N_6986);
xor U9969 (N_9969,N_7251,N_7895);
xor U9970 (N_9970,N_7074,N_7524);
and U9971 (N_9971,N_6203,N_7648);
xnor U9972 (N_9972,N_7184,N_6593);
nor U9973 (N_9973,N_7872,N_7262);
or U9974 (N_9974,N_7071,N_7502);
nand U9975 (N_9975,N_6683,N_7044);
or U9976 (N_9976,N_7842,N_7316);
and U9977 (N_9977,N_7860,N_6534);
xor U9978 (N_9978,N_7798,N_6979);
and U9979 (N_9979,N_7463,N_7227);
xnor U9980 (N_9980,N_6862,N_6664);
and U9981 (N_9981,N_6764,N_6251);
and U9982 (N_9982,N_7039,N_7978);
or U9983 (N_9983,N_7883,N_6107);
xor U9984 (N_9984,N_6162,N_7393);
nand U9985 (N_9985,N_7242,N_6100);
or U9986 (N_9986,N_6250,N_7512);
nor U9987 (N_9987,N_7925,N_6899);
nand U9988 (N_9988,N_6341,N_6994);
xor U9989 (N_9989,N_7085,N_7277);
nor U9990 (N_9990,N_7375,N_6236);
and U9991 (N_9991,N_7059,N_7011);
and U9992 (N_9992,N_6409,N_7099);
nor U9993 (N_9993,N_7415,N_6928);
xnor U9994 (N_9994,N_6665,N_6097);
and U9995 (N_9995,N_7402,N_7079);
xnor U9996 (N_9996,N_6068,N_7598);
and U9997 (N_9997,N_6795,N_6093);
and U9998 (N_9998,N_6771,N_7597);
nand U9999 (N_9999,N_6000,N_6290);
xor U10000 (N_10000,N_8057,N_9017);
or U10001 (N_10001,N_8082,N_9124);
nand U10002 (N_10002,N_8758,N_9871);
nand U10003 (N_10003,N_8982,N_8967);
and U10004 (N_10004,N_8553,N_8478);
xnor U10005 (N_10005,N_9183,N_8364);
and U10006 (N_10006,N_8606,N_8937);
nand U10007 (N_10007,N_8083,N_9331);
xnor U10008 (N_10008,N_9199,N_9329);
or U10009 (N_10009,N_8262,N_8915);
xnor U10010 (N_10010,N_8298,N_9317);
and U10011 (N_10011,N_9729,N_8064);
or U10012 (N_10012,N_9578,N_8702);
and U10013 (N_10013,N_8344,N_9401);
or U10014 (N_10014,N_9351,N_9007);
and U10015 (N_10015,N_8030,N_9090);
and U10016 (N_10016,N_9024,N_8407);
nor U10017 (N_10017,N_9405,N_9256);
xor U10018 (N_10018,N_8384,N_8871);
nand U10019 (N_10019,N_8315,N_8366);
nand U10020 (N_10020,N_9078,N_9043);
or U10021 (N_10021,N_9733,N_9192);
or U10022 (N_10022,N_9867,N_9113);
or U10023 (N_10023,N_9369,N_8657);
nand U10024 (N_10024,N_9925,N_8971);
or U10025 (N_10025,N_8374,N_9986);
and U10026 (N_10026,N_9518,N_9559);
and U10027 (N_10027,N_8746,N_9533);
or U10028 (N_10028,N_8129,N_8730);
nor U10029 (N_10029,N_9220,N_9773);
and U10030 (N_10030,N_9900,N_8261);
and U10031 (N_10031,N_9165,N_8097);
nor U10032 (N_10032,N_8290,N_9276);
or U10033 (N_10033,N_8334,N_8470);
xor U10034 (N_10034,N_8667,N_8922);
and U10035 (N_10035,N_8940,N_8049);
nand U10036 (N_10036,N_9501,N_8965);
xnor U10037 (N_10037,N_9715,N_8080);
and U10038 (N_10038,N_9621,N_9308);
and U10039 (N_10039,N_9380,N_8009);
nand U10040 (N_10040,N_8681,N_9130);
nor U10041 (N_10041,N_9322,N_9747);
and U10042 (N_10042,N_8095,N_9321);
and U10043 (N_10043,N_9262,N_9623);
nor U10044 (N_10044,N_8687,N_8398);
xor U10045 (N_10045,N_8283,N_9544);
or U10046 (N_10046,N_8905,N_8427);
and U10047 (N_10047,N_8012,N_9525);
and U10048 (N_10048,N_9253,N_8775);
xnor U10049 (N_10049,N_9575,N_8980);
nor U10050 (N_10050,N_9981,N_9516);
nor U10051 (N_10051,N_8647,N_8753);
xor U10052 (N_10052,N_9683,N_8409);
nand U10053 (N_10053,N_8093,N_9497);
nor U10054 (N_10054,N_8473,N_8482);
or U10055 (N_10055,N_9645,N_9954);
or U10056 (N_10056,N_9615,N_9837);
xor U10057 (N_10057,N_8695,N_8063);
and U10058 (N_10058,N_8259,N_8472);
xor U10059 (N_10059,N_8287,N_9073);
xor U10060 (N_10060,N_9144,N_8679);
or U10061 (N_10061,N_8782,N_9147);
xnor U10062 (N_10062,N_8300,N_8458);
or U10063 (N_10063,N_9161,N_9422);
nor U10064 (N_10064,N_8068,N_8737);
xnor U10065 (N_10065,N_9781,N_9899);
xnor U10066 (N_10066,N_9096,N_8588);
and U10067 (N_10067,N_8425,N_8579);
xor U10068 (N_10068,N_9806,N_8763);
or U10069 (N_10069,N_9601,N_8524);
and U10070 (N_10070,N_9242,N_9085);
nor U10071 (N_10071,N_8581,N_8600);
or U10072 (N_10072,N_9767,N_9949);
nand U10073 (N_10073,N_8826,N_9528);
nand U10074 (N_10074,N_9968,N_9931);
xor U10075 (N_10075,N_9841,N_9857);
xor U10076 (N_10076,N_9226,N_8860);
or U10077 (N_10077,N_8304,N_8712);
nor U10078 (N_10078,N_8123,N_8224);
xnor U10079 (N_10079,N_9038,N_9500);
or U10080 (N_10080,N_9221,N_8680);
and U10081 (N_10081,N_9983,N_9285);
and U10082 (N_10082,N_9917,N_9785);
nand U10083 (N_10083,N_8421,N_9919);
and U10084 (N_10084,N_9157,N_8430);
nand U10085 (N_10085,N_9873,N_9265);
nor U10086 (N_10086,N_9803,N_9102);
xor U10087 (N_10087,N_9774,N_8833);
xor U10088 (N_10088,N_9959,N_8279);
or U10089 (N_10089,N_9456,N_9576);
and U10090 (N_10090,N_9622,N_8174);
xnor U10091 (N_10091,N_9977,N_8343);
nor U10092 (N_10092,N_8997,N_9200);
and U10093 (N_10093,N_8120,N_8518);
nand U10094 (N_10094,N_9674,N_9882);
and U10095 (N_10095,N_9318,N_8335);
nor U10096 (N_10096,N_8992,N_8620);
xnor U10097 (N_10097,N_9418,N_9269);
nand U10098 (N_10098,N_8011,N_8875);
nor U10099 (N_10099,N_8501,N_8928);
or U10100 (N_10100,N_9975,N_8526);
nand U10101 (N_10101,N_8358,N_9398);
nand U10102 (N_10102,N_9914,N_8655);
nand U10103 (N_10103,N_8154,N_8053);
nor U10104 (N_10104,N_9039,N_8769);
nand U10105 (N_10105,N_8329,N_9897);
or U10106 (N_10106,N_8172,N_8943);
or U10107 (N_10107,N_9514,N_8295);
nand U10108 (N_10108,N_9783,N_8449);
and U10109 (N_10109,N_9376,N_8536);
nand U10110 (N_10110,N_9540,N_8079);
nor U10111 (N_10111,N_8622,N_9379);
nor U10112 (N_10112,N_9435,N_8502);
and U10113 (N_10113,N_8133,N_9554);
nand U10114 (N_10114,N_8336,N_8217);
nor U10115 (N_10115,N_8519,N_8312);
and U10116 (N_10116,N_9423,N_9598);
xnor U10117 (N_10117,N_9313,N_9104);
xnor U10118 (N_10118,N_9833,N_8525);
nand U10119 (N_10119,N_8929,N_8834);
or U10120 (N_10120,N_8515,N_9595);
nand U10121 (N_10121,N_9128,N_9698);
nor U10122 (N_10122,N_9574,N_8453);
or U10123 (N_10123,N_9413,N_8465);
nand U10124 (N_10124,N_8031,N_8350);
nor U10125 (N_10125,N_9805,N_9976);
and U10126 (N_10126,N_8050,N_8894);
nand U10127 (N_10127,N_9924,N_8020);
nand U10128 (N_10128,N_9932,N_9241);
nor U10129 (N_10129,N_9270,N_8991);
and U10130 (N_10130,N_8459,N_8561);
or U10131 (N_10131,N_8511,N_9403);
xor U10132 (N_10132,N_9772,N_8745);
nand U10133 (N_10133,N_8109,N_9510);
and U10134 (N_10134,N_8665,N_9751);
nand U10135 (N_10135,N_9964,N_9667);
nor U10136 (N_10136,N_9929,N_9235);
xor U10137 (N_10137,N_9439,N_8069);
xor U10138 (N_10138,N_8917,N_8925);
nor U10139 (N_10139,N_9709,N_9569);
nor U10140 (N_10140,N_9126,N_8740);
nand U10141 (N_10141,N_8062,N_9912);
and U10142 (N_10142,N_8564,N_9196);
xor U10143 (N_10143,N_9030,N_9763);
nor U10144 (N_10144,N_8151,N_9652);
and U10145 (N_10145,N_8642,N_8978);
nor U10146 (N_10146,N_8110,N_8509);
and U10147 (N_10147,N_9362,N_8999);
or U10148 (N_10148,N_9400,N_8376);
xor U10149 (N_10149,N_8193,N_9182);
or U10150 (N_10150,N_8149,N_8682);
nand U10151 (N_10151,N_9207,N_9489);
or U10152 (N_10152,N_8005,N_9287);
and U10153 (N_10153,N_9014,N_8504);
nor U10154 (N_10154,N_8206,N_9381);
or U10155 (N_10155,N_9771,N_9260);
or U10156 (N_10156,N_8963,N_9672);
xnor U10157 (N_10157,N_9033,N_9546);
nand U10158 (N_10158,N_8241,N_8571);
and U10159 (N_10159,N_8400,N_8696);
xnor U10160 (N_10160,N_9795,N_8408);
nand U10161 (N_10161,N_8480,N_9465);
nor U10162 (N_10162,N_8061,N_8533);
and U10163 (N_10163,N_8264,N_8896);
nand U10164 (N_10164,N_9719,N_9116);
nor U10165 (N_10165,N_9635,N_8071);
and U10166 (N_10166,N_8729,N_8497);
nand U10167 (N_10167,N_8603,N_9300);
nand U10168 (N_10168,N_8495,N_9708);
xnor U10169 (N_10169,N_9835,N_9630);
nand U10170 (N_10170,N_9868,N_8773);
xnor U10171 (N_10171,N_8195,N_9099);
nand U10172 (N_10172,N_9086,N_9206);
or U10173 (N_10173,N_8327,N_8945);
and U10174 (N_10174,N_8878,N_8332);
nor U10175 (N_10175,N_8556,N_9442);
nand U10176 (N_10176,N_9408,N_9399);
nor U10177 (N_10177,N_8722,N_8422);
and U10178 (N_10178,N_8897,N_8245);
and U10179 (N_10179,N_8612,N_9586);
or U10180 (N_10180,N_8212,N_8662);
nand U10181 (N_10181,N_8218,N_8546);
xnor U10182 (N_10182,N_8469,N_8727);
nor U10183 (N_10183,N_8522,N_8903);
nor U10184 (N_10184,N_9738,N_8957);
nand U10185 (N_10185,N_9666,N_9108);
xnor U10186 (N_10186,N_9892,N_9168);
nand U10187 (N_10187,N_9962,N_9686);
xnor U10188 (N_10188,N_9943,N_8951);
or U10189 (N_10189,N_8067,N_8391);
nor U10190 (N_10190,N_9972,N_8652);
xnor U10191 (N_10191,N_8454,N_9676);
nand U10192 (N_10192,N_8705,N_9987);
xor U10193 (N_10193,N_9561,N_9343);
and U10194 (N_10194,N_9885,N_8370);
nand U10195 (N_10195,N_8508,N_9046);
xor U10196 (N_10196,N_8537,N_9764);
or U10197 (N_10197,N_9958,N_9813);
nand U10198 (N_10198,N_8013,N_9591);
nand U10199 (N_10199,N_8186,N_9011);
nand U10200 (N_10200,N_8242,N_8165);
nor U10201 (N_10201,N_9947,N_9498);
nand U10202 (N_10202,N_8790,N_8555);
nor U10203 (N_10203,N_9349,N_8293);
xnor U10204 (N_10204,N_9816,N_8969);
xor U10205 (N_10205,N_8395,N_8260);
xnor U10206 (N_10206,N_9850,N_8314);
nor U10207 (N_10207,N_8565,N_8285);
nand U10208 (N_10208,N_8200,N_9117);
nand U10209 (N_10209,N_9750,N_9992);
nor U10210 (N_10210,N_9861,N_9782);
or U10211 (N_10211,N_8590,N_8568);
xnor U10212 (N_10212,N_8498,N_8551);
nor U10213 (N_10213,N_8631,N_9565);
nor U10214 (N_10214,N_8448,N_9524);
nor U10215 (N_10215,N_9072,N_9583);
xor U10216 (N_10216,N_9197,N_9682);
xnor U10217 (N_10217,N_9848,N_9870);
and U10218 (N_10218,N_8379,N_8308);
nand U10219 (N_10219,N_8204,N_8791);
xor U10220 (N_10220,N_9452,N_9557);
nor U10221 (N_10221,N_8911,N_9809);
nand U10222 (N_10222,N_9890,N_8996);
nand U10223 (N_10223,N_8108,N_8091);
or U10224 (N_10224,N_9286,N_9801);
and U10225 (N_10225,N_8514,N_9991);
nand U10226 (N_10226,N_8443,N_9617);
or U10227 (N_10227,N_9780,N_8641);
or U10228 (N_10228,N_8632,N_9891);
nor U10229 (N_10229,N_9082,N_8716);
nor U10230 (N_10230,N_9984,N_8222);
or U10231 (N_10231,N_9603,N_9307);
xnor U10232 (N_10232,N_8356,N_9315);
and U10233 (N_10233,N_9215,N_8294);
and U10234 (N_10234,N_9471,N_9744);
nand U10235 (N_10235,N_8816,N_9697);
nand U10236 (N_10236,N_8948,N_8263);
nor U10237 (N_10237,N_8693,N_9228);
xor U10238 (N_10238,N_8118,N_9732);
xnor U10239 (N_10239,N_9211,N_8254);
and U10240 (N_10240,N_8277,N_9702);
nor U10241 (N_10241,N_9083,N_9613);
and U10242 (N_10242,N_8764,N_9787);
xnor U10243 (N_10243,N_9414,N_9704);
nand U10244 (N_10244,N_8196,N_9999);
nor U10245 (N_10245,N_8756,N_8543);
or U10246 (N_10246,N_8851,N_8780);
or U10247 (N_10247,N_9974,N_9110);
nor U10248 (N_10248,N_9677,N_9012);
and U10249 (N_10249,N_8732,N_8209);
xor U10250 (N_10250,N_8574,N_9409);
nand U10251 (N_10251,N_9004,N_8248);
or U10252 (N_10252,N_8309,N_8220);
nand U10253 (N_10253,N_9469,N_8070);
or U10254 (N_10254,N_8893,N_9556);
nor U10255 (N_10255,N_9365,N_9188);
and U10256 (N_10256,N_9626,N_8055);
nand U10257 (N_10257,N_8906,N_9736);
and U10258 (N_10258,N_8168,N_9716);
or U10259 (N_10259,N_8651,N_8862);
nor U10260 (N_10260,N_8086,N_8988);
or U10261 (N_10261,N_9955,N_8231);
nand U10262 (N_10262,N_8914,N_8866);
nand U10263 (N_10263,N_8783,N_8723);
nand U10264 (N_10264,N_9155,N_9386);
or U10265 (N_10265,N_9830,N_9768);
and U10266 (N_10266,N_8022,N_8836);
xor U10267 (N_10267,N_8240,N_8252);
or U10268 (N_10268,N_9597,N_9132);
xnor U10269 (N_10269,N_8964,N_9378);
nand U10270 (N_10270,N_8461,N_9258);
nand U10271 (N_10271,N_8197,N_8023);
or U10272 (N_10272,N_8827,N_8138);
nand U10273 (N_10273,N_9415,N_8008);
xor U10274 (N_10274,N_9874,N_9859);
nand U10275 (N_10275,N_9562,N_8406);
nor U10276 (N_10276,N_8349,N_8238);
and U10277 (N_10277,N_8132,N_8604);
xnor U10278 (N_10278,N_9411,N_8800);
or U10279 (N_10279,N_9190,N_9163);
and U10280 (N_10280,N_8365,N_8128);
nor U10281 (N_10281,N_9948,N_8595);
or U10282 (N_10282,N_8090,N_8778);
nor U10283 (N_10283,N_8001,N_8414);
nor U10284 (N_10284,N_8301,N_9552);
xor U10285 (N_10285,N_8829,N_9394);
xor U10286 (N_10286,N_8249,N_9358);
xnor U10287 (N_10287,N_8542,N_8513);
nand U10288 (N_10288,N_8962,N_8239);
nor U10289 (N_10289,N_8396,N_8664);
or U10290 (N_10290,N_8328,N_9057);
nor U10291 (N_10291,N_8188,N_9926);
and U10292 (N_10292,N_9000,N_8203);
and U10293 (N_10293,N_8105,N_8500);
or U10294 (N_10294,N_9884,N_8506);
and U10295 (N_10295,N_8496,N_8340);
or U10296 (N_10296,N_8942,N_8464);
or U10297 (N_10297,N_8767,N_9081);
nor U10298 (N_10298,N_8706,N_8171);
nand U10299 (N_10299,N_9808,N_9407);
or U10300 (N_10300,N_9105,N_9657);
nand U10301 (N_10301,N_8228,N_8257);
nor U10302 (N_10302,N_9055,N_9725);
and U10303 (N_10303,N_8912,N_9311);
nand U10304 (N_10304,N_8699,N_8968);
nand U10305 (N_10305,N_8768,N_9205);
or U10306 (N_10306,N_8970,N_8939);
xnor U10307 (N_10307,N_8910,N_9222);
nand U10308 (N_10308,N_9723,N_9034);
nand U10309 (N_10309,N_9076,N_9208);
or U10310 (N_10310,N_8688,N_8845);
nor U10311 (N_10311,N_8490,N_9445);
nor U10312 (N_10312,N_8191,N_8347);
or U10313 (N_10313,N_8813,N_8385);
or U10314 (N_10314,N_9154,N_9338);
xor U10315 (N_10315,N_9600,N_8724);
xor U10316 (N_10316,N_8798,N_9015);
or U10317 (N_10317,N_8831,N_9555);
or U10318 (N_10318,N_9450,N_8666);
and U10319 (N_10319,N_8380,N_8796);
or U10320 (N_10320,N_8236,N_9960);
nor U10321 (N_10321,N_8100,N_8265);
nor U10322 (N_10322,N_9075,N_8394);
xnor U10323 (N_10323,N_8182,N_8742);
xnor U10324 (N_10324,N_9864,N_9171);
and U10325 (N_10325,N_8362,N_8529);
xor U10326 (N_10326,N_9920,N_9519);
nor U10327 (N_10327,N_9520,N_8886);
nand U10328 (N_10328,N_8021,N_8268);
nand U10329 (N_10329,N_9137,N_8754);
xor U10330 (N_10330,N_9934,N_9969);
xor U10331 (N_10331,N_9181,N_8690);
and U10332 (N_10332,N_8145,N_9189);
xor U10333 (N_10333,N_8296,N_9582);
and U10334 (N_10334,N_9037,N_8368);
or U10335 (N_10335,N_8802,N_9599);
xor U10336 (N_10336,N_8572,N_9843);
xor U10337 (N_10337,N_8272,N_9614);
xor U10338 (N_10338,N_9941,N_8479);
nand U10339 (N_10339,N_9254,N_9443);
nor U10340 (N_10340,N_8985,N_8616);
nor U10341 (N_10341,N_9695,N_8330);
xor U10342 (N_10342,N_9511,N_8507);
and U10343 (N_10343,N_8981,N_8383);
and U10344 (N_10344,N_8435,N_9397);
xnor U10345 (N_10345,N_8270,N_9508);
nand U10346 (N_10346,N_9333,N_8441);
or U10347 (N_10347,N_9690,N_8460);
xor U10348 (N_10348,N_9204,N_8934);
nand U10349 (N_10349,N_8805,N_9323);
and U10350 (N_10350,N_8892,N_8960);
nand U10351 (N_10351,N_9939,N_9566);
nand U10352 (N_10352,N_9010,N_8205);
xor U10353 (N_10353,N_8772,N_8499);
or U10354 (N_10354,N_9143,N_9389);
and U10355 (N_10355,N_8865,N_9392);
nor U10356 (N_10356,N_8671,N_9093);
or U10357 (N_10357,N_9122,N_9480);
nor U10358 (N_10358,N_8351,N_8403);
xnor U10359 (N_10359,N_9526,N_9357);
or U10360 (N_10360,N_9827,N_9769);
nor U10361 (N_10361,N_8078,N_8438);
or U10362 (N_10362,N_8809,N_9250);
and U10363 (N_10363,N_9361,N_9754);
nand U10364 (N_10364,N_9743,N_9167);
nor U10365 (N_10365,N_8202,N_8444);
and U10366 (N_10366,N_9304,N_9506);
nor U10367 (N_10367,N_8413,N_8255);
and U10368 (N_10368,N_8879,N_8434);
nor U10369 (N_10369,N_9956,N_9921);
nand U10370 (N_10370,N_9457,N_8440);
xor U10371 (N_10371,N_9354,N_9573);
or U10372 (N_10372,N_9374,N_8361);
nor U10373 (N_10373,N_9066,N_8986);
xnor U10374 (N_10374,N_9098,N_8776);
or U10375 (N_10375,N_9340,N_9728);
xor U10376 (N_10376,N_8375,N_9474);
nor U10377 (N_10377,N_8872,N_8602);
nor U10378 (N_10378,N_8748,N_9918);
nor U10379 (N_10379,N_9838,N_8321);
nor U10380 (N_10380,N_9640,N_9044);
nand U10381 (N_10381,N_9326,N_9458);
xor U10382 (N_10382,N_9114,N_8787);
nor U10383 (N_10383,N_8784,N_9159);
or U10384 (N_10384,N_9359,N_8855);
nor U10385 (N_10385,N_9701,N_8562);
xnor U10386 (N_10386,N_8142,N_8420);
or U10387 (N_10387,N_8058,N_9534);
or U10388 (N_10388,N_8491,N_8567);
xor U10389 (N_10389,N_9644,N_8119);
nor U10390 (N_10390,N_8586,N_8794);
or U10391 (N_10391,N_9330,N_9663);
and U10392 (N_10392,N_8274,N_8307);
nand U10393 (N_10393,N_9819,N_9699);
xnor U10394 (N_10394,N_9650,N_9029);
xnor U10395 (N_10395,N_9146,N_9395);
nand U10396 (N_10396,N_8393,N_8734);
and U10397 (N_10397,N_8966,N_8932);
nand U10398 (N_10398,N_9825,N_9097);
nor U10399 (N_10399,N_8369,N_8094);
and U10400 (N_10400,N_9001,N_9735);
xor U10401 (N_10401,N_8346,N_8818);
nand U10402 (N_10402,N_8028,N_9616);
xnor U10403 (N_10403,N_8814,N_9823);
nor U10404 (N_10404,N_8663,N_9971);
nand U10405 (N_10405,N_9472,N_9022);
nor U10406 (N_10406,N_9101,N_8373);
xor U10407 (N_10407,N_8592,N_9404);
or U10408 (N_10408,N_8806,N_8289);
nor U10409 (N_10409,N_9047,N_9995);
nand U10410 (N_10410,N_8000,N_9495);
and U10411 (N_10411,N_8244,N_8733);
nor U10412 (N_10412,N_9726,N_8779);
xnor U10413 (N_10413,N_9305,N_8885);
and U10414 (N_10414,N_9927,N_8042);
nand U10415 (N_10415,N_8534,N_8147);
nand U10416 (N_10416,N_8569,N_9367);
and U10417 (N_10417,N_8326,N_8704);
or U10418 (N_10418,N_9123,N_9145);
or U10419 (N_10419,N_8014,N_8125);
or U10420 (N_10420,N_9278,N_8150);
xnor U10421 (N_10421,N_9517,N_8575);
xnor U10422 (N_10422,N_9180,N_9631);
nand U10423 (N_10423,N_9681,N_9612);
nor U10424 (N_10424,N_8096,N_9063);
nand U10425 (N_10425,N_9289,N_9431);
xor U10426 (N_10426,N_9074,N_8412);
nand U10427 (N_10427,N_8804,N_8505);
nand U10428 (N_10428,N_9910,N_9051);
nor U10429 (N_10429,N_8085,N_8825);
and U10430 (N_10430,N_8956,N_9788);
nor U10431 (N_10431,N_8628,N_8954);
nor U10432 (N_10432,N_9084,N_8726);
xnor U10433 (N_10433,N_9447,N_9855);
nor U10434 (N_10434,N_9527,N_9722);
nand U10435 (N_10435,N_9664,N_8907);
and U10436 (N_10436,N_8528,N_8751);
nor U10437 (N_10437,N_8276,N_8591);
xnor U10438 (N_10438,N_9303,N_8617);
xnor U10439 (N_10439,N_9348,N_9653);
nand U10440 (N_10440,N_9173,N_8003);
or U10441 (N_10441,N_9247,N_8765);
nor U10442 (N_10442,N_9989,N_8757);
and U10443 (N_10443,N_8952,N_9705);
nand U10444 (N_10444,N_9632,N_8432);
xnor U10445 (N_10445,N_8883,N_9179);
or U10446 (N_10446,N_9696,N_9779);
or U10447 (N_10447,N_8402,N_9493);
xor U10448 (N_10448,N_9641,N_8477);
nand U10449 (N_10449,N_9793,N_9761);
or U10450 (N_10450,N_8835,N_8483);
nor U10451 (N_10451,N_9370,N_9261);
and U10452 (N_10452,N_8635,N_8549);
and U10453 (N_10453,N_9230,N_9125);
xor U10454 (N_10454,N_9296,N_8429);
xor U10455 (N_10455,N_9068,N_8913);
or U10456 (N_10456,N_9290,N_9095);
nand U10457 (N_10457,N_9930,N_8801);
nor U10458 (N_10458,N_9255,N_8025);
or U10459 (N_10459,N_9547,N_8760);
or U10460 (N_10460,N_8823,N_8399);
nand U10461 (N_10461,N_8576,N_9945);
nor U10462 (N_10462,N_9814,N_9065);
or U10463 (N_10463,N_8799,N_9027);
nand U10464 (N_10464,N_9319,N_8961);
and U10465 (N_10465,N_8452,N_8707);
nor U10466 (N_10466,N_9755,N_8474);
or U10467 (N_10467,N_8056,N_8051);
xor U10468 (N_10468,N_8207,N_8322);
and U10469 (N_10469,N_9893,N_9268);
or U10470 (N_10470,N_9127,N_9172);
and U10471 (N_10471,N_8153,N_8887);
nand U10472 (N_10472,N_9138,N_9913);
and U10473 (N_10473,N_9152,N_9071);
xnor U10474 (N_10474,N_9203,N_8341);
xnor U10475 (N_10475,N_9002,N_8048);
or U10476 (N_10476,N_9839,N_9866);
or U10477 (N_10477,N_9089,N_9217);
and U10478 (N_10478,N_9703,N_9201);
xor U10479 (N_10479,N_9023,N_8250);
xor U10480 (N_10480,N_8156,N_9312);
xor U10481 (N_10481,N_9025,N_9396);
xnor U10482 (N_10482,N_9572,N_8807);
nor U10483 (N_10483,N_9467,N_8392);
and U10484 (N_10484,N_9232,N_9903);
nand U10485 (N_10485,N_8060,N_8266);
xnor U10486 (N_10486,N_9119,N_9951);
nand U10487 (N_10487,N_9935,N_9713);
xor U10488 (N_10488,N_9462,N_9282);
or U10489 (N_10489,N_8401,N_8035);
nor U10490 (N_10490,N_8233,N_8367);
xnor U10491 (N_10491,N_9150,N_8485);
nand U10492 (N_10492,N_8607,N_9325);
nand U10493 (N_10493,N_9717,N_8348);
xor U10494 (N_10494,N_8319,N_9234);
or U10495 (N_10495,N_8931,N_8708);
xor U10496 (N_10496,N_8643,N_9727);
and U10497 (N_10497,N_8439,N_9342);
or U10498 (N_10498,N_8891,N_8424);
and U10499 (N_10499,N_9088,N_9639);
and U10500 (N_10500,N_8979,N_8541);
xnor U10501 (N_10501,N_8725,N_9902);
nor U10502 (N_10502,N_9106,N_9229);
xnor U10503 (N_10503,N_8691,N_9542);
nand U10504 (N_10504,N_8215,N_8715);
and U10505 (N_10505,N_8089,N_9100);
xor U10506 (N_10506,N_9094,N_9352);
xor U10507 (N_10507,N_9382,N_9994);
and U10508 (N_10508,N_8927,N_8700);
and U10509 (N_10509,N_8098,N_8557);
or U10510 (N_10510,N_8530,N_9053);
nor U10511 (N_10511,N_8735,N_9477);
nand U10512 (N_10512,N_8626,N_9259);
and U10513 (N_10513,N_9654,N_9753);
or U10514 (N_10514,N_8492,N_8987);
and U10515 (N_10515,N_8750,N_9360);
nor U10516 (N_10516,N_8489,N_8993);
or U10517 (N_10517,N_9706,N_9888);
and U10518 (N_10518,N_8868,N_8977);
or U10519 (N_10519,N_8629,N_9822);
nor U10520 (N_10520,N_9901,N_9393);
and U10521 (N_10521,N_8711,N_9804);
and U10522 (N_10522,N_9016,N_9383);
or U10523 (N_10523,N_9406,N_8674);
nor U10524 (N_10524,N_8933,N_9852);
xnor U10525 (N_10525,N_9794,N_9463);
or U10526 (N_10526,N_9069,N_8117);
or U10527 (N_10527,N_8837,N_9120);
or U10528 (N_10528,N_9549,N_8410);
xnor U10529 (N_10529,N_9950,N_8689);
nor U10530 (N_10530,N_8084,N_9740);
and U10531 (N_10531,N_8856,N_9335);
xnor U10532 (N_10532,N_8785,N_8175);
xor U10533 (N_10533,N_8318,N_9385);
xor U10534 (N_10534,N_8299,N_8088);
nor U10535 (N_10535,N_9602,N_8577);
or U10536 (N_10536,N_9784,N_9679);
nand U10537 (N_10537,N_8843,N_8625);
nand U10538 (N_10538,N_9579,N_9210);
xor U10539 (N_10539,N_8797,N_8447);
nor U10540 (N_10540,N_8223,N_9149);
or U10541 (N_10541,N_8701,N_9610);
nand U10542 (N_10542,N_9907,N_8795);
or U10543 (N_10543,N_8324,N_8653);
nor U10544 (N_10544,N_9481,N_8857);
xor U10545 (N_10545,N_8026,N_8678);
nor U10546 (N_10546,N_9236,N_9944);
and U10547 (N_10547,N_9739,N_8848);
or U10548 (N_10548,N_9680,N_9938);
xor U10549 (N_10549,N_8467,N_8623);
xnor U10550 (N_10550,N_9824,N_8876);
or U10551 (N_10551,N_9842,N_8173);
xor U10552 (N_10552,N_9252,N_8558);
and U10553 (N_10553,N_8738,N_8808);
and U10554 (N_10554,N_9731,N_8390);
xor U10555 (N_10555,N_9223,N_8476);
or U10556 (N_10556,N_9845,N_8323);
or U10557 (N_10557,N_8821,N_8728);
or U10558 (N_10558,N_9344,N_9832);
xor U10559 (N_10559,N_9856,N_9064);
or U10560 (N_10560,N_8849,N_9563);
and U10561 (N_10561,N_9077,N_9898);
and U10562 (N_10562,N_9227,N_8357);
and U10563 (N_10563,N_8130,N_9240);
or U10564 (N_10564,N_8455,N_9844);
nand U10565 (N_10565,N_9766,N_8881);
or U10566 (N_10566,N_8882,N_8388);
nor U10567 (N_10567,N_9271,N_9797);
nand U10568 (N_10568,N_9668,N_9453);
nand U10569 (N_10569,N_8924,N_9166);
nor U10570 (N_10570,N_9417,N_8038);
or U10571 (N_10571,N_9812,N_8180);
nor U10572 (N_10572,N_9860,N_9567);
xnor U10573 (N_10573,N_9478,N_8437);
nor U10574 (N_10574,N_9940,N_8076);
xor U10575 (N_10575,N_8972,N_8634);
or U10576 (N_10576,N_9693,N_9185);
and U10577 (N_10577,N_9473,N_9170);
xnor U10578 (N_10578,N_8548,N_8297);
nor U10579 (N_10579,N_9334,N_9537);
xor U10580 (N_10580,N_9800,N_9491);
nor U10581 (N_10581,N_8955,N_9560);
nand U10582 (N_10582,N_8015,N_9432);
or U10583 (N_10583,N_9273,N_9353);
or U10584 (N_10584,N_8077,N_9134);
or U10585 (N_10585,N_9748,N_8633);
and U10586 (N_10586,N_8864,N_8194);
nand U10587 (N_10587,N_9345,N_8320);
xor U10588 (N_10588,N_8761,N_8126);
or U10589 (N_10589,N_9451,N_9248);
nand U10590 (N_10590,N_8890,N_9799);
xnor U10591 (N_10591,N_8815,N_9026);
and U10592 (N_10592,N_9571,N_8850);
or U10593 (N_10593,N_9062,N_8019);
nand U10594 (N_10594,N_9297,N_9153);
or U10595 (N_10595,N_8106,N_8024);
and U10596 (N_10596,N_9483,N_8810);
or U10597 (N_10597,N_9618,N_8941);
xnor U10598 (N_10598,N_8593,N_8908);
nand U10599 (N_10599,N_9018,N_8619);
nor U10600 (N_10600,N_8503,N_8316);
xnor U10601 (N_10601,N_8853,N_8516);
and U10602 (N_10602,N_8423,N_9933);
and U10603 (N_10603,N_9658,N_9515);
nor U10604 (N_10604,N_8610,N_9817);
and U10605 (N_10605,N_8990,N_8353);
nor U10606 (N_10606,N_9757,N_9056);
and U10607 (N_10607,N_8115,N_9908);
nor U10608 (N_10608,N_9426,N_9080);
nand U10609 (N_10609,N_9828,N_9551);
nand U10610 (N_10610,N_8135,N_9742);
or U10611 (N_10611,N_8377,N_8983);
xnor U10612 (N_10612,N_8280,N_9543);
nor U10613 (N_10613,N_8547,N_8136);
nand U10614 (N_10614,N_8898,N_9851);
nor U10615 (N_10615,N_9459,N_9484);
nor U10616 (N_10616,N_8037,N_9589);
nor U10617 (N_10617,N_8159,N_9267);
or U10618 (N_10618,N_8762,N_9320);
nand U10619 (N_10619,N_9020,N_8339);
nand U10620 (N_10620,N_9390,N_8994);
and U10621 (N_10621,N_9580,N_8844);
nor U10622 (N_10622,N_9584,N_8043);
nand U10623 (N_10623,N_9880,N_9636);
or U10624 (N_10624,N_8185,N_9765);
or U10625 (N_10625,N_9624,N_8976);
nand U10626 (N_10626,N_8004,N_9156);
or U10627 (N_10627,N_9887,N_8462);
nor U10628 (N_10628,N_8958,N_9671);
and U10629 (N_10629,N_9662,N_9410);
xor U10630 (N_10630,N_8731,N_8935);
or U10631 (N_10631,N_9107,N_8075);
nor U10632 (N_10632,N_8002,N_9219);
nand U10633 (N_10633,N_8658,N_9169);
nor U10634 (N_10634,N_8419,N_9337);
xor U10635 (N_10635,N_8131,N_8599);
and U10636 (N_10636,N_8397,N_8611);
nor U10637 (N_10637,N_9476,N_8721);
and U10638 (N_10638,N_9049,N_8870);
or U10639 (N_10639,N_9040,N_8709);
and U10640 (N_10640,N_8921,N_9231);
or U10641 (N_10641,N_9499,N_9264);
xnor U10642 (N_10642,N_9590,N_9041);
xnor U10643 (N_10643,N_9876,N_8580);
xor U10644 (N_10644,N_8271,N_8155);
xnor U10645 (N_10645,N_9802,N_8512);
nor U10646 (N_10646,N_9504,N_9328);
xor U10647 (N_10647,N_8141,N_8660);
nor U10648 (N_10648,N_9301,N_9470);
and U10649 (N_10649,N_9627,N_8317);
xor U10650 (N_10650,N_8792,N_9140);
xnor U10651 (N_10651,N_8036,N_9553);
nand U10652 (N_10652,N_9878,N_8124);
and U10653 (N_10653,N_9758,N_8584);
nor U10654 (N_10654,N_9911,N_9283);
nand U10655 (N_10655,N_9996,N_9148);
xor U10656 (N_10656,N_8627,N_9239);
nand U10657 (N_10657,N_8659,N_8686);
and U10658 (N_10658,N_9734,N_9896);
xor U10659 (N_10659,N_9523,N_8523);
and U10660 (N_10660,N_9225,N_9512);
nor U10661 (N_10661,N_9294,N_8121);
nand U10662 (N_10662,N_9836,N_9928);
xor U10663 (N_10663,N_8824,N_9494);
and U10664 (N_10664,N_9036,N_8139);
xnor U10665 (N_10665,N_9388,N_9142);
or U10666 (N_10666,N_9060,N_8984);
and U10667 (N_10667,N_8668,N_9214);
and U10668 (N_10668,N_8847,N_8854);
nand U10669 (N_10669,N_8938,N_9013);
nor U10670 (N_10670,N_9997,N_9529);
nor U10671 (N_10671,N_9121,N_8644);
xor U10672 (N_10672,N_9310,N_9760);
and U10673 (N_10673,N_8127,N_9466);
xnor U10674 (N_10674,N_9087,N_9692);
and U10675 (N_10675,N_8052,N_9059);
xor U10676 (N_10676,N_9558,N_8788);
and U10677 (N_10677,N_8583,N_9741);
or U10678 (N_10678,N_8661,N_9350);
xnor U10679 (N_10679,N_8899,N_8900);
and U10680 (N_10680,N_9141,N_9642);
xnor U10681 (N_10681,N_8111,N_8284);
nand U10682 (N_10682,N_8457,N_8039);
nand U10683 (N_10683,N_8382,N_8947);
xnor U10684 (N_10684,N_8428,N_9243);
nor U10685 (N_10685,N_9973,N_8007);
nand U10686 (N_10686,N_8446,N_8275);
nor U10687 (N_10687,N_9050,N_8415);
nand U10688 (N_10688,N_9826,N_8615);
xnor U10689 (N_10689,N_8072,N_9923);
or U10690 (N_10690,N_8291,N_8920);
xor U10691 (N_10691,N_8614,N_9058);
nand U10692 (N_10692,N_9455,N_9881);
and U10693 (N_10693,N_9299,N_8486);
xnor U10694 (N_10694,N_8578,N_9831);
nor U10695 (N_10695,N_8869,N_8181);
and U10696 (N_10696,N_8527,N_9637);
or U10697 (N_10697,N_9605,N_8841);
nor U10698 (N_10698,N_9048,N_9638);
or U10699 (N_10699,N_9678,N_8672);
nor U10700 (N_10700,N_9606,N_9440);
and U10701 (N_10701,N_8770,N_8027);
nor U10702 (N_10702,N_8717,N_8989);
and U10703 (N_10703,N_8718,N_8047);
and U10704 (N_10704,N_9594,N_8192);
xor U10705 (N_10705,N_8640,N_9212);
or U10706 (N_10706,N_9377,N_8563);
or U10707 (N_10707,N_9346,N_8975);
nor U10708 (N_10708,N_9685,N_8859);
nor U10709 (N_10709,N_9965,N_8311);
or U10710 (N_10710,N_9535,N_9879);
or U10711 (N_10711,N_9790,N_8338);
or U10712 (N_10712,N_8302,N_8998);
nand U10713 (N_10713,N_8179,N_8573);
xnor U10714 (N_10714,N_8286,N_8213);
nand U10715 (N_10715,N_9427,N_8585);
or U10716 (N_10716,N_9186,N_9776);
and U10717 (N_10717,N_9280,N_8995);
nand U10718 (N_10718,N_9752,N_8786);
nor U10719 (N_10719,N_9191,N_8251);
or U10720 (N_10720,N_8433,N_9536);
nand U10721 (N_10721,N_9079,N_8253);
or U10722 (N_10722,N_9649,N_8143);
or U10723 (N_10723,N_8137,N_9587);
xnor U10724 (N_10724,N_9218,N_8842);
or U10725 (N_10725,N_8601,N_8587);
xor U10726 (N_10726,N_8305,N_9436);
xor U10727 (N_10727,N_9889,N_8540);
xnor U10728 (N_10728,N_9460,N_9438);
or U10729 (N_10729,N_9238,N_9193);
and U10730 (N_10730,N_9670,N_8538);
or U10731 (N_10731,N_8822,N_8065);
xor U10732 (N_10732,N_8953,N_8450);
and U10733 (N_10733,N_8074,N_8256);
or U10734 (N_10734,N_8624,N_9607);
or U10735 (N_10735,N_9988,N_8582);
or U10736 (N_10736,N_8487,N_9858);
and U10737 (N_10737,N_9257,N_9877);
or U10738 (N_10738,N_9846,N_9363);
nand U10739 (N_10739,N_8113,N_9957);
and U10740 (N_10740,N_9875,N_9990);
nand U10741 (N_10741,N_9786,N_8066);
or U10742 (N_10742,N_8685,N_9118);
nand U10743 (N_10743,N_8959,N_9777);
nor U10744 (N_10744,N_8861,N_8648);
and U10745 (N_10745,N_8517,N_9922);
or U10746 (N_10746,N_9906,N_9293);
nor U10747 (N_10747,N_9479,N_9112);
xnor U10748 (N_10748,N_8888,N_9611);
nand U10749 (N_10749,N_9316,N_8714);
nand U10750 (N_10750,N_9651,N_9869);
nor U10751 (N_10751,N_9647,N_8521);
nor U10752 (N_10752,N_9496,N_8531);
or U10753 (N_10753,N_8442,N_9746);
and U10754 (N_10754,N_8719,N_8759);
and U10755 (N_10755,N_9009,N_8973);
and U10756 (N_10756,N_8677,N_8589);
nand U10757 (N_10757,N_9673,N_9656);
nand U10758 (N_10758,N_9233,N_9375);
nand U10759 (N_10759,N_9284,N_9045);
xnor U10760 (N_10760,N_8744,N_9619);
and U10761 (N_10761,N_8736,N_9756);
or U10762 (N_10762,N_9021,N_8163);
nand U10763 (N_10763,N_8646,N_8654);
nand U10764 (N_10764,N_9620,N_8858);
xor U10765 (N_10765,N_8184,N_8281);
nor U10766 (N_10766,N_8134,N_8880);
xor U10767 (N_10767,N_8313,N_8475);
xnor U10768 (N_10768,N_8466,N_8103);
nand U10769 (N_10769,N_9532,N_8227);
nor U10770 (N_10770,N_9272,N_8713);
and U10771 (N_10771,N_9811,N_8550);
nor U10772 (N_10772,N_9135,N_8010);
and U10773 (N_10773,N_9894,N_9249);
and U10774 (N_10774,N_8532,N_8481);
nor U10775 (N_10775,N_8418,N_8649);
nand U10776 (N_10776,N_9834,N_8451);
and U10777 (N_10777,N_9263,N_8636);
nand U10778 (N_10778,N_9430,N_8645);
nor U10779 (N_10779,N_8747,N_8046);
and U10780 (N_10780,N_8445,N_9031);
and U10781 (N_10781,N_9291,N_8189);
nand U10782 (N_10782,N_8176,N_8670);
xor U10783 (N_10783,N_8554,N_8029);
or U10784 (N_10784,N_9298,N_9505);
nor U10785 (N_10785,N_9054,N_8793);
xnor U10786 (N_10786,N_9905,N_8918);
and U10787 (N_10787,N_8278,N_9292);
or U10788 (N_10788,N_9548,N_9070);
and U10789 (N_10789,N_9454,N_9688);
nor U10790 (N_10790,N_8178,N_9849);
and U10791 (N_10791,N_9032,N_9129);
nand U10792 (N_10792,N_8216,N_9433);
and U10793 (N_10793,N_9336,N_8471);
xor U10794 (N_10794,N_8006,N_9245);
xnor U10795 (N_10795,N_9865,N_8411);
or U10796 (N_10796,N_9862,N_8597);
nand U10797 (N_10797,N_9295,N_9464);
xnor U10798 (N_10798,N_9530,N_9364);
nor U10799 (N_10799,N_9448,N_9368);
nand U10800 (N_10800,N_8081,N_9371);
xor U10801 (N_10801,N_9821,N_9904);
nand U10802 (N_10802,N_8535,N_9687);
and U10803 (N_10803,N_9509,N_9246);
nor U10804 (N_10804,N_9998,N_8819);
and U10805 (N_10805,N_9655,N_8463);
or U10806 (N_10806,N_9485,N_9721);
or U10807 (N_10807,N_8177,N_9646);
xor U10808 (N_10808,N_8812,N_8288);
and U10809 (N_10809,N_9005,N_8811);
or U10810 (N_10810,N_9840,N_8596);
and U10811 (N_10811,N_9052,N_9347);
nor U10812 (N_10812,N_8638,N_9691);
or U10813 (N_10813,N_8743,N_8749);
xor U10814 (N_10814,N_9720,N_9006);
xor U10815 (N_10815,N_8162,N_8684);
xnor U10816 (N_10816,N_8692,N_8867);
or U10817 (N_10817,N_8034,N_9792);
or U10818 (N_10818,N_8045,N_9184);
xor U10819 (N_10819,N_8214,N_8114);
xor U10820 (N_10820,N_9416,N_8637);
or U10821 (N_10821,N_8230,N_9661);
nand U10822 (N_10822,N_8187,N_8613);
xor U10823 (N_10823,N_9985,N_8656);
xnor U10824 (N_10824,N_8650,N_9391);
or U10825 (N_10825,N_8669,N_8303);
nor U10826 (N_10826,N_9468,N_9942);
nor U10827 (N_10827,N_8386,N_8909);
nor U10828 (N_10828,N_9982,N_9158);
nor U10829 (N_10829,N_8608,N_9251);
xor U10830 (N_10830,N_8234,N_8741);
or U10831 (N_10831,N_9568,N_8360);
nand U10832 (N_10832,N_8710,N_9461);
xnor U10833 (N_10833,N_9541,N_9402);
or U10834 (N_10834,N_9115,N_9490);
or U10835 (N_10835,N_8387,N_9384);
xnor U10836 (N_10836,N_9711,N_8354);
nor U10837 (N_10837,N_8325,N_8889);
xnor U10838 (N_10838,N_9538,N_9895);
and U10839 (N_10839,N_8148,N_9366);
or U10840 (N_10840,N_9872,N_9091);
xnor U10841 (N_10841,N_9550,N_9213);
and U10842 (N_10842,N_9244,N_9428);
xnor U10843 (N_10843,N_9604,N_9502);
or U10844 (N_10844,N_9820,N_8292);
nor U10845 (N_10845,N_8273,N_8488);
or U10846 (N_10846,N_8152,N_8161);
nor U10847 (N_10847,N_9503,N_8246);
nor U10848 (N_10848,N_9324,N_8017);
nor U10849 (N_10849,N_8916,N_8389);
or U10850 (N_10850,N_9111,N_8493);
xnor U10851 (N_10851,N_8164,N_8258);
xnor U10852 (N_10852,N_9028,N_9332);
or U10853 (N_10853,N_9449,N_8372);
and U10854 (N_10854,N_8552,N_8839);
xor U10855 (N_10855,N_8771,N_8950);
xor U10856 (N_10856,N_9570,N_9314);
or U10857 (N_10857,N_8211,N_9202);
and U10858 (N_10858,N_9434,N_8494);
xnor U10859 (N_10859,N_9327,N_9710);
or U10860 (N_10860,N_9486,N_9980);
nand U10861 (N_10861,N_8877,N_9588);
or U10862 (N_10862,N_8902,N_9937);
nand U10863 (N_10863,N_8371,N_8974);
and U10864 (N_10864,N_9545,N_9778);
and U10865 (N_10865,N_8144,N_9209);
xnor U10866 (N_10866,N_8235,N_8884);
nor U10867 (N_10867,N_9978,N_9675);
xnor U10868 (N_10868,N_9531,N_9648);
or U10869 (N_10869,N_9724,N_9737);
and U10870 (N_10870,N_8381,N_8016);
or U10871 (N_10871,N_8237,N_8752);
and U10872 (N_10872,N_9224,N_9577);
nor U10873 (N_10873,N_9198,N_9288);
nand U10874 (N_10874,N_8104,N_9694);
or U10875 (N_10875,N_8781,N_9419);
and U10876 (N_10876,N_9131,N_9669);
nand U10877 (N_10877,N_9356,N_8863);
xnor U10878 (N_10878,N_8766,N_9444);
nand U10879 (N_10879,N_9482,N_9970);
xnor U10880 (N_10880,N_8566,N_9492);
nor U10881 (N_10881,N_8210,N_8116);
nand U10882 (N_10882,N_9507,N_8901);
xor U10883 (N_10883,N_8949,N_9689);
xor U10884 (N_10884,N_9810,N_9585);
xnor U10885 (N_10885,N_8405,N_8404);
nand U10886 (N_10886,N_9372,N_9581);
nand U10887 (N_10887,N_8158,N_9634);
nand U10888 (N_10888,N_8033,N_8140);
xor U10889 (N_10889,N_9936,N_8673);
or U10890 (N_10890,N_9909,N_9665);
and U10891 (N_10891,N_9596,N_9700);
and U10892 (N_10892,N_9160,N_9425);
nor U10893 (N_10893,N_9707,N_9151);
nand U10894 (N_10894,N_8018,N_8777);
nand U10895 (N_10895,N_9625,N_8160);
and U10896 (N_10896,N_9176,N_9593);
nor U10897 (N_10897,N_9643,N_9718);
or U10898 (N_10898,N_8510,N_8694);
and U10899 (N_10899,N_9373,N_8087);
or U10900 (N_10900,N_9035,N_8789);
nor U10901 (N_10901,N_9067,N_8208);
and U10902 (N_10902,N_8229,N_9791);
or U10903 (N_10903,N_9475,N_9863);
or U10904 (N_10904,N_9139,N_9659);
xnor U10905 (N_10905,N_9749,N_9109);
nor U10906 (N_10906,N_8431,N_9592);
nor U10907 (N_10907,N_9775,N_8895);
or U10908 (N_10908,N_8363,N_8840);
or U10909 (N_10909,N_9886,N_8355);
xor U10910 (N_10910,N_9770,N_8426);
or U10911 (N_10911,N_9966,N_9277);
and U10912 (N_10912,N_8904,N_8167);
or U10913 (N_10913,N_8226,N_9420);
nor U10914 (N_10914,N_8944,N_9302);
xor U10915 (N_10915,N_8874,N_8102);
xor U10916 (N_10916,N_8310,N_9387);
xnor U10917 (N_10917,N_8817,N_9424);
or U10918 (N_10918,N_9175,N_8946);
and U10919 (N_10919,N_9847,N_8040);
xor U10920 (N_10920,N_8594,N_9174);
xnor U10921 (N_10921,N_8539,N_9762);
xnor U10922 (N_10922,N_8219,N_9633);
and U10923 (N_10923,N_9341,N_8852);
nand U10924 (N_10924,N_8170,N_9103);
nor U10925 (N_10925,N_8183,N_8436);
xor U10926 (N_10926,N_9355,N_8267);
xor U10927 (N_10927,N_8598,N_9194);
or U10928 (N_10928,N_8232,N_9339);
nor U10929 (N_10929,N_9712,N_8269);
or U10930 (N_10930,N_8820,N_8609);
nand U10931 (N_10931,N_9162,N_9759);
nand U10932 (N_10932,N_8306,N_8675);
nand U10933 (N_10933,N_8378,N_9829);
and U10934 (N_10934,N_8621,N_9946);
or U10935 (N_10935,N_9883,N_9608);
nor U10936 (N_10936,N_8484,N_9967);
nand U10937 (N_10937,N_8054,N_8359);
nand U10938 (N_10938,N_8345,N_9854);
or U10939 (N_10939,N_8559,N_8468);
or U10940 (N_10940,N_9953,N_9745);
nor U10941 (N_10941,N_8342,N_8846);
or U10942 (N_10942,N_8828,N_8605);
or U10943 (N_10943,N_8774,N_8560);
and U10944 (N_10944,N_8416,N_8169);
nor U10945 (N_10945,N_8683,N_8099);
or U10946 (N_10946,N_9275,N_8739);
xnor U10947 (N_10947,N_8417,N_8190);
nand U10948 (N_10948,N_8873,N_9092);
xor U10949 (N_10949,N_8618,N_9684);
and U10950 (N_10950,N_8199,N_8112);
or U10951 (N_10951,N_8225,N_8697);
and U10952 (N_10952,N_8570,N_9714);
and U10953 (N_10953,N_8073,N_9019);
xnor U10954 (N_10954,N_9916,N_9730);
xor U10955 (N_10955,N_9008,N_9003);
nand U10956 (N_10956,N_9853,N_8703);
and U10957 (N_10957,N_8630,N_9963);
or U10958 (N_10958,N_9429,N_8243);
nand U10959 (N_10959,N_8122,N_9628);
xor U10960 (N_10960,N_8032,N_9195);
nor U10961 (N_10961,N_8838,N_8923);
nand U10962 (N_10962,N_9807,N_9177);
xor U10963 (N_10963,N_9216,N_9281);
nand U10964 (N_10964,N_8059,N_9279);
xor U10965 (N_10965,N_8698,N_9513);
nand U10966 (N_10966,N_9961,N_8041);
nor U10967 (N_10967,N_8676,N_8919);
nor U10968 (N_10968,N_8936,N_9915);
or U10969 (N_10969,N_8331,N_9993);
xor U10970 (N_10970,N_9522,N_9488);
nor U10971 (N_10971,N_9609,N_8044);
nor U10972 (N_10972,N_9042,N_9274);
or U10973 (N_10973,N_8101,N_8930);
nor U10974 (N_10974,N_8720,N_9818);
or U10975 (N_10975,N_9187,N_9164);
nand U10976 (N_10976,N_9446,N_8146);
nor U10977 (N_10977,N_8520,N_8107);
and U10978 (N_10978,N_9266,N_8803);
and U10979 (N_10979,N_9979,N_9815);
and U10980 (N_10980,N_9421,N_9309);
or U10981 (N_10981,N_8337,N_8456);
nor U10982 (N_10982,N_9061,N_9237);
nand U10983 (N_10983,N_8198,N_9629);
nor U10984 (N_10984,N_9306,N_9521);
xor U10985 (N_10985,N_9789,N_9660);
nor U10986 (N_10986,N_8545,N_8333);
xor U10987 (N_10987,N_8282,N_8755);
or U10988 (N_10988,N_9133,N_8639);
nand U10989 (N_10989,N_8201,N_9539);
nand U10990 (N_10990,N_8832,N_8926);
xnor U10991 (N_10991,N_9487,N_8166);
nand U10992 (N_10992,N_8352,N_9796);
or U10993 (N_10993,N_8830,N_9564);
nor U10994 (N_10994,N_9441,N_8247);
nor U10995 (N_10995,N_9178,N_9437);
nor U10996 (N_10996,N_8092,N_9798);
nand U10997 (N_10997,N_9136,N_8544);
xor U10998 (N_10998,N_9412,N_8157);
nand U10999 (N_10999,N_9952,N_8221);
or U11000 (N_11000,N_8033,N_9918);
xor U11001 (N_11001,N_9171,N_9957);
nand U11002 (N_11002,N_8799,N_8025);
and U11003 (N_11003,N_9191,N_8318);
xor U11004 (N_11004,N_9110,N_8253);
or U11005 (N_11005,N_8083,N_8429);
or U11006 (N_11006,N_9322,N_8264);
or U11007 (N_11007,N_9093,N_8500);
nor U11008 (N_11008,N_9723,N_9666);
xor U11009 (N_11009,N_9187,N_9783);
xor U11010 (N_11010,N_9971,N_8420);
or U11011 (N_11011,N_9603,N_8566);
nor U11012 (N_11012,N_8092,N_9810);
xnor U11013 (N_11013,N_9056,N_8578);
or U11014 (N_11014,N_9210,N_8444);
nor U11015 (N_11015,N_8312,N_8746);
or U11016 (N_11016,N_9139,N_8884);
and U11017 (N_11017,N_8197,N_8852);
and U11018 (N_11018,N_9548,N_8343);
nor U11019 (N_11019,N_8891,N_8739);
xnor U11020 (N_11020,N_9881,N_9619);
xor U11021 (N_11021,N_9037,N_8301);
and U11022 (N_11022,N_8189,N_9037);
nor U11023 (N_11023,N_8561,N_9230);
nor U11024 (N_11024,N_9829,N_9519);
or U11025 (N_11025,N_9117,N_9679);
xnor U11026 (N_11026,N_8341,N_9365);
xnor U11027 (N_11027,N_9835,N_9927);
xor U11028 (N_11028,N_9289,N_8508);
nor U11029 (N_11029,N_8752,N_8894);
or U11030 (N_11030,N_9194,N_9439);
and U11031 (N_11031,N_9948,N_8685);
or U11032 (N_11032,N_9023,N_9642);
xor U11033 (N_11033,N_8032,N_9697);
nor U11034 (N_11034,N_8275,N_8666);
xnor U11035 (N_11035,N_8259,N_8948);
xor U11036 (N_11036,N_9859,N_9364);
nand U11037 (N_11037,N_9663,N_9624);
and U11038 (N_11038,N_8207,N_8348);
nand U11039 (N_11039,N_9492,N_9169);
and U11040 (N_11040,N_9187,N_9365);
nand U11041 (N_11041,N_8074,N_9376);
and U11042 (N_11042,N_8785,N_8744);
and U11043 (N_11043,N_9115,N_8534);
nand U11044 (N_11044,N_8445,N_8034);
nand U11045 (N_11045,N_9648,N_8061);
or U11046 (N_11046,N_8583,N_8822);
and U11047 (N_11047,N_8995,N_9927);
nand U11048 (N_11048,N_8137,N_9282);
or U11049 (N_11049,N_9674,N_9579);
or U11050 (N_11050,N_9162,N_9217);
nor U11051 (N_11051,N_9387,N_9648);
or U11052 (N_11052,N_9987,N_9405);
or U11053 (N_11053,N_9631,N_8016);
nor U11054 (N_11054,N_9767,N_8151);
or U11055 (N_11055,N_8928,N_8380);
nor U11056 (N_11056,N_8665,N_9535);
or U11057 (N_11057,N_8353,N_9395);
nand U11058 (N_11058,N_9850,N_8657);
or U11059 (N_11059,N_8309,N_8601);
or U11060 (N_11060,N_9833,N_9965);
nor U11061 (N_11061,N_8394,N_9479);
nor U11062 (N_11062,N_8904,N_8991);
or U11063 (N_11063,N_8842,N_8959);
nor U11064 (N_11064,N_8314,N_9957);
nor U11065 (N_11065,N_9366,N_9850);
nand U11066 (N_11066,N_8501,N_8801);
and U11067 (N_11067,N_9015,N_9793);
nor U11068 (N_11068,N_8176,N_8812);
or U11069 (N_11069,N_8471,N_9100);
nand U11070 (N_11070,N_8007,N_8062);
or U11071 (N_11071,N_9500,N_8156);
or U11072 (N_11072,N_8837,N_9047);
nand U11073 (N_11073,N_8595,N_8908);
and U11074 (N_11074,N_9588,N_9566);
nor U11075 (N_11075,N_9916,N_9347);
nor U11076 (N_11076,N_8433,N_9969);
or U11077 (N_11077,N_8439,N_8028);
nor U11078 (N_11078,N_8682,N_8635);
or U11079 (N_11079,N_8990,N_8185);
xor U11080 (N_11080,N_9753,N_9295);
and U11081 (N_11081,N_9523,N_8325);
or U11082 (N_11082,N_9635,N_9781);
and U11083 (N_11083,N_8154,N_9476);
or U11084 (N_11084,N_8217,N_8676);
and U11085 (N_11085,N_8173,N_8197);
or U11086 (N_11086,N_8831,N_9267);
nand U11087 (N_11087,N_9822,N_9871);
xnor U11088 (N_11088,N_9147,N_9158);
and U11089 (N_11089,N_8075,N_9160);
and U11090 (N_11090,N_9066,N_8210);
nor U11091 (N_11091,N_9903,N_9452);
and U11092 (N_11092,N_8376,N_8739);
or U11093 (N_11093,N_8283,N_9127);
nand U11094 (N_11094,N_9659,N_8102);
nand U11095 (N_11095,N_8598,N_9051);
nor U11096 (N_11096,N_8870,N_8192);
nor U11097 (N_11097,N_8380,N_9584);
nand U11098 (N_11098,N_8331,N_8502);
xnor U11099 (N_11099,N_8075,N_9579);
xor U11100 (N_11100,N_9717,N_9157);
xnor U11101 (N_11101,N_9937,N_9510);
or U11102 (N_11102,N_8910,N_9245);
nand U11103 (N_11103,N_8155,N_9378);
nor U11104 (N_11104,N_9650,N_8871);
nand U11105 (N_11105,N_9625,N_9463);
xnor U11106 (N_11106,N_9942,N_8020);
xnor U11107 (N_11107,N_9923,N_8309);
nor U11108 (N_11108,N_9234,N_9103);
nand U11109 (N_11109,N_8443,N_9264);
xnor U11110 (N_11110,N_9853,N_8325);
and U11111 (N_11111,N_9790,N_9863);
and U11112 (N_11112,N_9704,N_9146);
and U11113 (N_11113,N_8869,N_9323);
or U11114 (N_11114,N_8431,N_9615);
nand U11115 (N_11115,N_8470,N_8872);
xor U11116 (N_11116,N_9278,N_9488);
and U11117 (N_11117,N_8670,N_9464);
and U11118 (N_11118,N_8382,N_8757);
or U11119 (N_11119,N_8633,N_8264);
or U11120 (N_11120,N_8877,N_9021);
and U11121 (N_11121,N_8111,N_8296);
or U11122 (N_11122,N_8790,N_9417);
xnor U11123 (N_11123,N_8608,N_8000);
and U11124 (N_11124,N_8796,N_9824);
xnor U11125 (N_11125,N_8745,N_8381);
nor U11126 (N_11126,N_8508,N_9452);
xor U11127 (N_11127,N_8424,N_9194);
or U11128 (N_11128,N_9432,N_9935);
nor U11129 (N_11129,N_8604,N_8925);
or U11130 (N_11130,N_8016,N_9364);
nor U11131 (N_11131,N_8158,N_8281);
xnor U11132 (N_11132,N_9025,N_9637);
nand U11133 (N_11133,N_8374,N_8817);
and U11134 (N_11134,N_8915,N_8385);
xnor U11135 (N_11135,N_9163,N_9376);
nand U11136 (N_11136,N_8091,N_9066);
or U11137 (N_11137,N_8391,N_8856);
nand U11138 (N_11138,N_9033,N_8913);
or U11139 (N_11139,N_9110,N_9964);
and U11140 (N_11140,N_8336,N_9688);
xnor U11141 (N_11141,N_8406,N_9618);
xor U11142 (N_11142,N_8150,N_8645);
nor U11143 (N_11143,N_9613,N_9989);
and U11144 (N_11144,N_8509,N_8865);
and U11145 (N_11145,N_9175,N_8573);
nor U11146 (N_11146,N_8860,N_8267);
or U11147 (N_11147,N_9760,N_9330);
nor U11148 (N_11148,N_9973,N_8414);
nand U11149 (N_11149,N_9790,N_8716);
xnor U11150 (N_11150,N_8556,N_9288);
and U11151 (N_11151,N_8745,N_8478);
or U11152 (N_11152,N_8750,N_9527);
or U11153 (N_11153,N_8910,N_9924);
nor U11154 (N_11154,N_8913,N_9812);
nor U11155 (N_11155,N_9921,N_8709);
nor U11156 (N_11156,N_8936,N_9096);
xnor U11157 (N_11157,N_8214,N_8714);
and U11158 (N_11158,N_8959,N_8888);
nor U11159 (N_11159,N_8268,N_8351);
or U11160 (N_11160,N_8269,N_8597);
nor U11161 (N_11161,N_8624,N_8756);
nand U11162 (N_11162,N_8181,N_9646);
xor U11163 (N_11163,N_9088,N_8331);
nand U11164 (N_11164,N_9047,N_8178);
or U11165 (N_11165,N_8972,N_8654);
and U11166 (N_11166,N_9537,N_9853);
nand U11167 (N_11167,N_8067,N_8102);
xnor U11168 (N_11168,N_8545,N_9988);
nor U11169 (N_11169,N_9715,N_9131);
and U11170 (N_11170,N_8260,N_9773);
xnor U11171 (N_11171,N_8388,N_9450);
and U11172 (N_11172,N_8498,N_9497);
nand U11173 (N_11173,N_8101,N_9978);
xnor U11174 (N_11174,N_8980,N_9029);
or U11175 (N_11175,N_9239,N_8543);
nor U11176 (N_11176,N_8148,N_8220);
nand U11177 (N_11177,N_8617,N_8155);
xor U11178 (N_11178,N_9214,N_8960);
xor U11179 (N_11179,N_8946,N_9398);
nor U11180 (N_11180,N_8276,N_8072);
nor U11181 (N_11181,N_8211,N_8874);
nor U11182 (N_11182,N_8379,N_9286);
and U11183 (N_11183,N_9000,N_9586);
nor U11184 (N_11184,N_8461,N_9581);
or U11185 (N_11185,N_9740,N_8486);
nor U11186 (N_11186,N_8525,N_9482);
xnor U11187 (N_11187,N_9064,N_8216);
xnor U11188 (N_11188,N_8737,N_8554);
xnor U11189 (N_11189,N_8773,N_8905);
xor U11190 (N_11190,N_8607,N_8947);
nand U11191 (N_11191,N_8437,N_8708);
and U11192 (N_11192,N_9842,N_9423);
nand U11193 (N_11193,N_9786,N_8348);
nor U11194 (N_11194,N_8490,N_9177);
nor U11195 (N_11195,N_9768,N_8724);
or U11196 (N_11196,N_8239,N_9286);
nand U11197 (N_11197,N_8341,N_8862);
or U11198 (N_11198,N_8038,N_8446);
xor U11199 (N_11199,N_8074,N_9579);
xnor U11200 (N_11200,N_9403,N_9757);
nand U11201 (N_11201,N_8646,N_8796);
nor U11202 (N_11202,N_9227,N_8163);
or U11203 (N_11203,N_9928,N_9006);
and U11204 (N_11204,N_8027,N_8858);
nor U11205 (N_11205,N_9886,N_9454);
nand U11206 (N_11206,N_9901,N_9754);
or U11207 (N_11207,N_8497,N_9605);
nor U11208 (N_11208,N_8740,N_9350);
xor U11209 (N_11209,N_8719,N_8393);
or U11210 (N_11210,N_9600,N_9834);
and U11211 (N_11211,N_9627,N_8713);
xnor U11212 (N_11212,N_8550,N_9632);
or U11213 (N_11213,N_9987,N_9393);
and U11214 (N_11214,N_8785,N_9590);
xnor U11215 (N_11215,N_9256,N_8056);
xnor U11216 (N_11216,N_9991,N_8234);
nor U11217 (N_11217,N_8537,N_9593);
nand U11218 (N_11218,N_8266,N_9974);
xnor U11219 (N_11219,N_9073,N_9832);
nor U11220 (N_11220,N_9739,N_9392);
xor U11221 (N_11221,N_8258,N_8808);
and U11222 (N_11222,N_9536,N_8715);
xor U11223 (N_11223,N_8107,N_9889);
and U11224 (N_11224,N_9377,N_8998);
nor U11225 (N_11225,N_8165,N_8332);
nand U11226 (N_11226,N_9916,N_8997);
nor U11227 (N_11227,N_8186,N_8942);
nor U11228 (N_11228,N_8473,N_9964);
and U11229 (N_11229,N_9810,N_8254);
nand U11230 (N_11230,N_8779,N_9968);
or U11231 (N_11231,N_9591,N_8839);
and U11232 (N_11232,N_8055,N_9168);
nor U11233 (N_11233,N_9732,N_9499);
nand U11234 (N_11234,N_9746,N_9674);
nand U11235 (N_11235,N_8807,N_9395);
and U11236 (N_11236,N_9849,N_9002);
and U11237 (N_11237,N_8306,N_8659);
nor U11238 (N_11238,N_9530,N_8454);
nor U11239 (N_11239,N_8482,N_8530);
and U11240 (N_11240,N_8719,N_9135);
nor U11241 (N_11241,N_8001,N_8218);
nor U11242 (N_11242,N_8004,N_8317);
and U11243 (N_11243,N_9848,N_9819);
or U11244 (N_11244,N_9341,N_8094);
xnor U11245 (N_11245,N_9324,N_9823);
nand U11246 (N_11246,N_8532,N_8804);
nand U11247 (N_11247,N_9066,N_9033);
nand U11248 (N_11248,N_8812,N_8781);
and U11249 (N_11249,N_9591,N_8231);
xnor U11250 (N_11250,N_8342,N_9499);
nor U11251 (N_11251,N_9624,N_9105);
and U11252 (N_11252,N_9096,N_9147);
xor U11253 (N_11253,N_8844,N_9418);
and U11254 (N_11254,N_8368,N_9755);
nor U11255 (N_11255,N_8147,N_8386);
nor U11256 (N_11256,N_8741,N_9894);
nand U11257 (N_11257,N_9703,N_8356);
xnor U11258 (N_11258,N_8960,N_8339);
and U11259 (N_11259,N_9268,N_9875);
nor U11260 (N_11260,N_8680,N_8634);
and U11261 (N_11261,N_8504,N_8971);
or U11262 (N_11262,N_9827,N_9358);
and U11263 (N_11263,N_8757,N_9750);
or U11264 (N_11264,N_8963,N_9811);
xor U11265 (N_11265,N_8776,N_8612);
or U11266 (N_11266,N_8539,N_9882);
nand U11267 (N_11267,N_8427,N_9803);
nor U11268 (N_11268,N_9284,N_8447);
nor U11269 (N_11269,N_9370,N_9663);
or U11270 (N_11270,N_9484,N_8185);
or U11271 (N_11271,N_8096,N_9256);
nor U11272 (N_11272,N_9602,N_8919);
and U11273 (N_11273,N_8802,N_9465);
and U11274 (N_11274,N_8776,N_9520);
nor U11275 (N_11275,N_9838,N_9942);
or U11276 (N_11276,N_8817,N_9282);
nor U11277 (N_11277,N_8225,N_9083);
nand U11278 (N_11278,N_9150,N_8009);
and U11279 (N_11279,N_9633,N_8204);
or U11280 (N_11280,N_9572,N_9654);
nor U11281 (N_11281,N_9984,N_8919);
xor U11282 (N_11282,N_8312,N_8595);
nor U11283 (N_11283,N_8837,N_9099);
or U11284 (N_11284,N_9458,N_8647);
nand U11285 (N_11285,N_8821,N_8637);
nand U11286 (N_11286,N_8043,N_8547);
nand U11287 (N_11287,N_8019,N_9869);
or U11288 (N_11288,N_9051,N_9886);
or U11289 (N_11289,N_9482,N_9048);
nand U11290 (N_11290,N_9559,N_8211);
nor U11291 (N_11291,N_9540,N_9380);
or U11292 (N_11292,N_9302,N_8371);
xnor U11293 (N_11293,N_8697,N_9151);
xnor U11294 (N_11294,N_9428,N_8064);
nor U11295 (N_11295,N_8127,N_8481);
xnor U11296 (N_11296,N_9609,N_8102);
xor U11297 (N_11297,N_9775,N_9317);
xnor U11298 (N_11298,N_8185,N_8162);
or U11299 (N_11299,N_8906,N_9493);
xnor U11300 (N_11300,N_9425,N_9613);
or U11301 (N_11301,N_8019,N_9645);
nor U11302 (N_11302,N_8659,N_9330);
or U11303 (N_11303,N_8265,N_9535);
xor U11304 (N_11304,N_8797,N_9137);
and U11305 (N_11305,N_9379,N_8569);
and U11306 (N_11306,N_8939,N_8051);
nand U11307 (N_11307,N_8203,N_8227);
nand U11308 (N_11308,N_8390,N_9229);
nand U11309 (N_11309,N_8554,N_8641);
xor U11310 (N_11310,N_9766,N_9931);
or U11311 (N_11311,N_9789,N_8889);
nor U11312 (N_11312,N_9191,N_8888);
and U11313 (N_11313,N_8676,N_8823);
or U11314 (N_11314,N_8201,N_9430);
and U11315 (N_11315,N_9388,N_8662);
nand U11316 (N_11316,N_8108,N_9750);
xor U11317 (N_11317,N_9496,N_8681);
xor U11318 (N_11318,N_8333,N_8757);
and U11319 (N_11319,N_8264,N_9317);
and U11320 (N_11320,N_9627,N_8427);
and U11321 (N_11321,N_9014,N_8077);
or U11322 (N_11322,N_8703,N_9896);
xor U11323 (N_11323,N_9768,N_9660);
and U11324 (N_11324,N_8019,N_9329);
nor U11325 (N_11325,N_8636,N_9384);
and U11326 (N_11326,N_9839,N_9768);
xor U11327 (N_11327,N_8520,N_8422);
nand U11328 (N_11328,N_8896,N_8713);
nand U11329 (N_11329,N_9135,N_8883);
nand U11330 (N_11330,N_9055,N_9728);
or U11331 (N_11331,N_8700,N_9229);
nand U11332 (N_11332,N_8076,N_9170);
or U11333 (N_11333,N_8071,N_9181);
and U11334 (N_11334,N_8770,N_8249);
nor U11335 (N_11335,N_9850,N_9478);
nand U11336 (N_11336,N_9696,N_8922);
nand U11337 (N_11337,N_8738,N_8488);
xor U11338 (N_11338,N_9576,N_9073);
xnor U11339 (N_11339,N_9431,N_9195);
and U11340 (N_11340,N_9031,N_8925);
xnor U11341 (N_11341,N_8460,N_9878);
nor U11342 (N_11342,N_8290,N_9676);
xnor U11343 (N_11343,N_8560,N_8497);
or U11344 (N_11344,N_9616,N_9366);
and U11345 (N_11345,N_8926,N_9365);
xnor U11346 (N_11346,N_9707,N_9489);
or U11347 (N_11347,N_9309,N_9282);
nor U11348 (N_11348,N_9183,N_8297);
or U11349 (N_11349,N_8782,N_9839);
or U11350 (N_11350,N_9511,N_9684);
xor U11351 (N_11351,N_9389,N_9608);
nand U11352 (N_11352,N_8347,N_9136);
nor U11353 (N_11353,N_9483,N_9758);
nand U11354 (N_11354,N_9518,N_9614);
nor U11355 (N_11355,N_8311,N_9295);
and U11356 (N_11356,N_8749,N_8477);
or U11357 (N_11357,N_9295,N_8973);
or U11358 (N_11358,N_8319,N_9902);
nand U11359 (N_11359,N_8217,N_8532);
nand U11360 (N_11360,N_9318,N_9757);
and U11361 (N_11361,N_9861,N_9885);
nand U11362 (N_11362,N_9394,N_8562);
nand U11363 (N_11363,N_9564,N_9207);
nand U11364 (N_11364,N_9297,N_8868);
nor U11365 (N_11365,N_8185,N_9232);
xnor U11366 (N_11366,N_8936,N_8725);
nand U11367 (N_11367,N_8180,N_8561);
nor U11368 (N_11368,N_9667,N_8226);
or U11369 (N_11369,N_8772,N_9588);
nor U11370 (N_11370,N_8379,N_9354);
and U11371 (N_11371,N_9113,N_9444);
xor U11372 (N_11372,N_8386,N_9949);
nand U11373 (N_11373,N_9566,N_9775);
or U11374 (N_11374,N_9515,N_9392);
and U11375 (N_11375,N_8260,N_9178);
and U11376 (N_11376,N_8848,N_8360);
nand U11377 (N_11377,N_9198,N_8270);
and U11378 (N_11378,N_8756,N_8109);
and U11379 (N_11379,N_8463,N_9276);
xnor U11380 (N_11380,N_9447,N_8033);
xnor U11381 (N_11381,N_9570,N_9917);
nand U11382 (N_11382,N_8274,N_8734);
nand U11383 (N_11383,N_8534,N_8193);
xnor U11384 (N_11384,N_9726,N_9761);
nand U11385 (N_11385,N_8017,N_9183);
xnor U11386 (N_11386,N_9415,N_8849);
and U11387 (N_11387,N_9111,N_9160);
nand U11388 (N_11388,N_8492,N_8125);
xor U11389 (N_11389,N_9496,N_9931);
nor U11390 (N_11390,N_9993,N_8653);
or U11391 (N_11391,N_8150,N_9768);
nand U11392 (N_11392,N_9156,N_8573);
nand U11393 (N_11393,N_8734,N_9266);
and U11394 (N_11394,N_8292,N_8046);
or U11395 (N_11395,N_8622,N_8895);
or U11396 (N_11396,N_9144,N_9489);
xor U11397 (N_11397,N_8163,N_9112);
nor U11398 (N_11398,N_8280,N_9631);
or U11399 (N_11399,N_8465,N_8850);
nand U11400 (N_11400,N_8705,N_8426);
and U11401 (N_11401,N_9000,N_9560);
and U11402 (N_11402,N_9837,N_8338);
or U11403 (N_11403,N_9162,N_8391);
and U11404 (N_11404,N_8158,N_9010);
xnor U11405 (N_11405,N_8546,N_9466);
xor U11406 (N_11406,N_8635,N_8870);
nand U11407 (N_11407,N_8882,N_9292);
nor U11408 (N_11408,N_9522,N_9797);
nand U11409 (N_11409,N_8344,N_9297);
or U11410 (N_11410,N_8916,N_8690);
or U11411 (N_11411,N_8474,N_8528);
and U11412 (N_11412,N_9166,N_9237);
or U11413 (N_11413,N_8396,N_8023);
and U11414 (N_11414,N_8309,N_9377);
and U11415 (N_11415,N_8308,N_8330);
xnor U11416 (N_11416,N_8400,N_9474);
xor U11417 (N_11417,N_9472,N_8659);
or U11418 (N_11418,N_9585,N_9118);
xor U11419 (N_11419,N_9036,N_9212);
and U11420 (N_11420,N_9849,N_9036);
xor U11421 (N_11421,N_9912,N_9002);
xnor U11422 (N_11422,N_8050,N_9480);
xor U11423 (N_11423,N_8759,N_8877);
nor U11424 (N_11424,N_9930,N_9351);
xor U11425 (N_11425,N_8239,N_9615);
nor U11426 (N_11426,N_9587,N_8032);
nor U11427 (N_11427,N_9610,N_9909);
and U11428 (N_11428,N_8005,N_8510);
or U11429 (N_11429,N_9576,N_8546);
xor U11430 (N_11430,N_8745,N_8477);
xnor U11431 (N_11431,N_9390,N_8385);
nand U11432 (N_11432,N_8242,N_8745);
or U11433 (N_11433,N_9396,N_9480);
nor U11434 (N_11434,N_8817,N_9076);
or U11435 (N_11435,N_8024,N_9093);
or U11436 (N_11436,N_9650,N_9553);
or U11437 (N_11437,N_8836,N_9105);
xor U11438 (N_11438,N_8162,N_8520);
nand U11439 (N_11439,N_9117,N_8632);
and U11440 (N_11440,N_8137,N_8800);
and U11441 (N_11441,N_8748,N_8166);
xor U11442 (N_11442,N_9465,N_8263);
nand U11443 (N_11443,N_8552,N_8010);
nor U11444 (N_11444,N_8519,N_9035);
xor U11445 (N_11445,N_9946,N_9253);
nor U11446 (N_11446,N_9149,N_9069);
nand U11447 (N_11447,N_9080,N_8445);
nor U11448 (N_11448,N_8436,N_9690);
xor U11449 (N_11449,N_8101,N_8931);
and U11450 (N_11450,N_8335,N_9015);
and U11451 (N_11451,N_9786,N_8524);
or U11452 (N_11452,N_9442,N_9422);
and U11453 (N_11453,N_8870,N_9130);
xnor U11454 (N_11454,N_9797,N_8412);
and U11455 (N_11455,N_9008,N_9828);
or U11456 (N_11456,N_8862,N_8602);
and U11457 (N_11457,N_9106,N_9128);
xor U11458 (N_11458,N_8980,N_8341);
and U11459 (N_11459,N_9107,N_8013);
xor U11460 (N_11460,N_8255,N_9501);
nand U11461 (N_11461,N_9956,N_9027);
and U11462 (N_11462,N_8997,N_9103);
and U11463 (N_11463,N_8067,N_8533);
nor U11464 (N_11464,N_9722,N_8668);
nand U11465 (N_11465,N_8824,N_9235);
xnor U11466 (N_11466,N_9456,N_9406);
xnor U11467 (N_11467,N_8435,N_9613);
nor U11468 (N_11468,N_8914,N_8803);
and U11469 (N_11469,N_9237,N_8963);
nor U11470 (N_11470,N_8363,N_8219);
and U11471 (N_11471,N_8093,N_8828);
nor U11472 (N_11472,N_8497,N_8185);
and U11473 (N_11473,N_8888,N_9385);
nor U11474 (N_11474,N_8964,N_8382);
nand U11475 (N_11475,N_8540,N_9473);
xor U11476 (N_11476,N_9265,N_9040);
nor U11477 (N_11477,N_9054,N_9708);
or U11478 (N_11478,N_8235,N_8337);
nand U11479 (N_11479,N_8664,N_8669);
or U11480 (N_11480,N_8596,N_9564);
or U11481 (N_11481,N_9847,N_8924);
xor U11482 (N_11482,N_8433,N_9314);
or U11483 (N_11483,N_8867,N_9598);
and U11484 (N_11484,N_9054,N_9567);
nor U11485 (N_11485,N_9768,N_9451);
nor U11486 (N_11486,N_9611,N_8773);
xor U11487 (N_11487,N_9280,N_9766);
nand U11488 (N_11488,N_9938,N_9359);
or U11489 (N_11489,N_8900,N_8542);
nor U11490 (N_11490,N_9821,N_8736);
or U11491 (N_11491,N_8497,N_8595);
nand U11492 (N_11492,N_8798,N_8870);
nor U11493 (N_11493,N_9895,N_8129);
nor U11494 (N_11494,N_8331,N_8728);
and U11495 (N_11495,N_8674,N_9651);
xnor U11496 (N_11496,N_9076,N_9059);
nor U11497 (N_11497,N_8640,N_8212);
nand U11498 (N_11498,N_8075,N_8496);
or U11499 (N_11499,N_9795,N_9222);
and U11500 (N_11500,N_8985,N_9905);
and U11501 (N_11501,N_9407,N_8576);
and U11502 (N_11502,N_9756,N_9139);
xor U11503 (N_11503,N_9173,N_9476);
and U11504 (N_11504,N_9412,N_8311);
nor U11505 (N_11505,N_9873,N_9009);
nor U11506 (N_11506,N_8371,N_8790);
nand U11507 (N_11507,N_8787,N_8547);
xor U11508 (N_11508,N_8921,N_9730);
and U11509 (N_11509,N_8725,N_8089);
or U11510 (N_11510,N_8480,N_9863);
xor U11511 (N_11511,N_8359,N_9055);
nor U11512 (N_11512,N_8973,N_9078);
and U11513 (N_11513,N_8829,N_9336);
or U11514 (N_11514,N_9603,N_8831);
nor U11515 (N_11515,N_8400,N_9904);
or U11516 (N_11516,N_9299,N_8373);
nor U11517 (N_11517,N_8985,N_9755);
nand U11518 (N_11518,N_8283,N_9671);
or U11519 (N_11519,N_8350,N_9041);
and U11520 (N_11520,N_8817,N_9524);
nand U11521 (N_11521,N_8847,N_8494);
and U11522 (N_11522,N_8645,N_8920);
and U11523 (N_11523,N_9035,N_9584);
nor U11524 (N_11524,N_8714,N_9189);
and U11525 (N_11525,N_8430,N_8570);
xnor U11526 (N_11526,N_8906,N_8288);
and U11527 (N_11527,N_8290,N_9388);
nor U11528 (N_11528,N_8608,N_9013);
nor U11529 (N_11529,N_9629,N_8582);
xnor U11530 (N_11530,N_8384,N_9632);
nand U11531 (N_11531,N_9264,N_9159);
xnor U11532 (N_11532,N_9667,N_9540);
and U11533 (N_11533,N_9844,N_8320);
or U11534 (N_11534,N_8263,N_9428);
and U11535 (N_11535,N_9896,N_9452);
xnor U11536 (N_11536,N_8909,N_8693);
nand U11537 (N_11537,N_9082,N_9747);
nand U11538 (N_11538,N_8751,N_9498);
and U11539 (N_11539,N_8438,N_9290);
nor U11540 (N_11540,N_9281,N_9114);
nor U11541 (N_11541,N_8622,N_9042);
or U11542 (N_11542,N_8106,N_9408);
and U11543 (N_11543,N_9337,N_9196);
xor U11544 (N_11544,N_8948,N_8230);
and U11545 (N_11545,N_9549,N_8827);
or U11546 (N_11546,N_9418,N_9475);
and U11547 (N_11547,N_8008,N_8847);
nand U11548 (N_11548,N_9174,N_9407);
or U11549 (N_11549,N_9360,N_9564);
xnor U11550 (N_11550,N_8407,N_8595);
xor U11551 (N_11551,N_9640,N_8314);
or U11552 (N_11552,N_9596,N_8938);
nand U11553 (N_11553,N_9084,N_8560);
or U11554 (N_11554,N_9540,N_9386);
nand U11555 (N_11555,N_9566,N_8532);
or U11556 (N_11556,N_9098,N_9082);
xor U11557 (N_11557,N_9582,N_8280);
xnor U11558 (N_11558,N_8529,N_9486);
xnor U11559 (N_11559,N_8210,N_9790);
nor U11560 (N_11560,N_8670,N_9123);
nor U11561 (N_11561,N_8061,N_9311);
or U11562 (N_11562,N_9691,N_8219);
and U11563 (N_11563,N_9141,N_9187);
nand U11564 (N_11564,N_9677,N_8934);
xor U11565 (N_11565,N_8773,N_9113);
nand U11566 (N_11566,N_8508,N_8492);
or U11567 (N_11567,N_8599,N_9946);
nand U11568 (N_11568,N_9589,N_9771);
xnor U11569 (N_11569,N_8745,N_9479);
nor U11570 (N_11570,N_8135,N_9431);
xor U11571 (N_11571,N_9926,N_9466);
nand U11572 (N_11572,N_9234,N_8131);
nor U11573 (N_11573,N_8159,N_8338);
xor U11574 (N_11574,N_8073,N_9553);
and U11575 (N_11575,N_9527,N_9090);
xor U11576 (N_11576,N_9302,N_9861);
and U11577 (N_11577,N_8490,N_9340);
or U11578 (N_11578,N_8889,N_9751);
or U11579 (N_11579,N_8598,N_9363);
nand U11580 (N_11580,N_8176,N_8964);
nor U11581 (N_11581,N_8008,N_8639);
and U11582 (N_11582,N_8807,N_8512);
nand U11583 (N_11583,N_9509,N_9220);
nor U11584 (N_11584,N_9784,N_8163);
xnor U11585 (N_11585,N_9268,N_9521);
and U11586 (N_11586,N_9651,N_9391);
nor U11587 (N_11587,N_9645,N_8858);
or U11588 (N_11588,N_9367,N_8400);
xor U11589 (N_11589,N_9939,N_9518);
xnor U11590 (N_11590,N_9340,N_8910);
or U11591 (N_11591,N_9948,N_8770);
nand U11592 (N_11592,N_8860,N_8733);
nor U11593 (N_11593,N_9877,N_8611);
and U11594 (N_11594,N_8433,N_9413);
xnor U11595 (N_11595,N_8203,N_8507);
nor U11596 (N_11596,N_9374,N_8541);
and U11597 (N_11597,N_9663,N_8686);
or U11598 (N_11598,N_8853,N_8753);
and U11599 (N_11599,N_9718,N_8797);
nor U11600 (N_11600,N_9395,N_9362);
nand U11601 (N_11601,N_8913,N_8370);
xor U11602 (N_11602,N_9405,N_9786);
nand U11603 (N_11603,N_9899,N_8165);
or U11604 (N_11604,N_9516,N_8216);
nand U11605 (N_11605,N_9832,N_8397);
nand U11606 (N_11606,N_8903,N_8437);
nand U11607 (N_11607,N_9229,N_9468);
nand U11608 (N_11608,N_8188,N_9394);
nor U11609 (N_11609,N_8594,N_8903);
and U11610 (N_11610,N_9880,N_8217);
and U11611 (N_11611,N_9590,N_8575);
nand U11612 (N_11612,N_8607,N_9690);
xnor U11613 (N_11613,N_9512,N_9184);
nor U11614 (N_11614,N_8100,N_9388);
and U11615 (N_11615,N_8719,N_9287);
and U11616 (N_11616,N_8404,N_8359);
or U11617 (N_11617,N_9939,N_9669);
xnor U11618 (N_11618,N_9622,N_9925);
and U11619 (N_11619,N_9598,N_8527);
nand U11620 (N_11620,N_9754,N_9566);
and U11621 (N_11621,N_9177,N_8977);
and U11622 (N_11622,N_9737,N_8895);
xor U11623 (N_11623,N_8679,N_9017);
nor U11624 (N_11624,N_8341,N_9053);
nor U11625 (N_11625,N_8688,N_8482);
nand U11626 (N_11626,N_9235,N_8815);
nor U11627 (N_11627,N_9885,N_9848);
or U11628 (N_11628,N_8300,N_9848);
nand U11629 (N_11629,N_8975,N_9128);
nand U11630 (N_11630,N_8064,N_8165);
or U11631 (N_11631,N_9221,N_9865);
nor U11632 (N_11632,N_8241,N_8230);
xor U11633 (N_11633,N_9371,N_9795);
and U11634 (N_11634,N_8933,N_9441);
and U11635 (N_11635,N_9252,N_9276);
nor U11636 (N_11636,N_8716,N_8096);
nand U11637 (N_11637,N_8535,N_9279);
nand U11638 (N_11638,N_9427,N_9405);
and U11639 (N_11639,N_9508,N_8513);
nand U11640 (N_11640,N_9746,N_8315);
nor U11641 (N_11641,N_9437,N_8909);
or U11642 (N_11642,N_8055,N_9649);
and U11643 (N_11643,N_8411,N_8512);
nand U11644 (N_11644,N_9337,N_8758);
or U11645 (N_11645,N_8691,N_9344);
xor U11646 (N_11646,N_8696,N_8083);
nand U11647 (N_11647,N_9324,N_9798);
nand U11648 (N_11648,N_9314,N_9077);
nor U11649 (N_11649,N_9574,N_9184);
nor U11650 (N_11650,N_8659,N_9405);
and U11651 (N_11651,N_8199,N_8791);
or U11652 (N_11652,N_9326,N_8077);
nor U11653 (N_11653,N_8285,N_9004);
nand U11654 (N_11654,N_9482,N_8050);
or U11655 (N_11655,N_8006,N_9772);
xnor U11656 (N_11656,N_8551,N_9633);
or U11657 (N_11657,N_8894,N_8287);
nor U11658 (N_11658,N_9175,N_9725);
or U11659 (N_11659,N_8466,N_9451);
and U11660 (N_11660,N_8503,N_8979);
or U11661 (N_11661,N_9714,N_8914);
nand U11662 (N_11662,N_8170,N_8372);
or U11663 (N_11663,N_9208,N_8519);
and U11664 (N_11664,N_9145,N_9174);
and U11665 (N_11665,N_9934,N_8799);
nor U11666 (N_11666,N_9385,N_8795);
and U11667 (N_11667,N_8524,N_8427);
nor U11668 (N_11668,N_8453,N_8469);
nand U11669 (N_11669,N_9401,N_8243);
nor U11670 (N_11670,N_8602,N_8782);
and U11671 (N_11671,N_8322,N_9409);
and U11672 (N_11672,N_8149,N_8953);
and U11673 (N_11673,N_9653,N_8754);
nor U11674 (N_11674,N_8856,N_9736);
or U11675 (N_11675,N_9545,N_9843);
nand U11676 (N_11676,N_9776,N_9992);
or U11677 (N_11677,N_8007,N_9031);
nor U11678 (N_11678,N_9901,N_9206);
xor U11679 (N_11679,N_8586,N_8715);
nor U11680 (N_11680,N_8812,N_9589);
nand U11681 (N_11681,N_8911,N_9043);
and U11682 (N_11682,N_9385,N_8823);
and U11683 (N_11683,N_9838,N_9172);
xnor U11684 (N_11684,N_9523,N_8608);
nor U11685 (N_11685,N_8676,N_8439);
and U11686 (N_11686,N_9052,N_8241);
nand U11687 (N_11687,N_9378,N_9412);
and U11688 (N_11688,N_9287,N_9908);
xor U11689 (N_11689,N_8168,N_9699);
or U11690 (N_11690,N_8083,N_9102);
and U11691 (N_11691,N_8274,N_8247);
or U11692 (N_11692,N_8643,N_8374);
nor U11693 (N_11693,N_9539,N_8281);
or U11694 (N_11694,N_9847,N_9891);
nor U11695 (N_11695,N_8112,N_8215);
or U11696 (N_11696,N_8112,N_9323);
and U11697 (N_11697,N_8849,N_8898);
xnor U11698 (N_11698,N_8412,N_8400);
nand U11699 (N_11699,N_9266,N_8326);
or U11700 (N_11700,N_8810,N_9449);
or U11701 (N_11701,N_8520,N_8085);
nand U11702 (N_11702,N_8729,N_9978);
nand U11703 (N_11703,N_8281,N_9597);
nor U11704 (N_11704,N_8069,N_8318);
or U11705 (N_11705,N_8171,N_8489);
xor U11706 (N_11706,N_8398,N_8341);
nor U11707 (N_11707,N_8460,N_9322);
or U11708 (N_11708,N_9076,N_8040);
nand U11709 (N_11709,N_8736,N_9357);
xnor U11710 (N_11710,N_8215,N_9996);
nand U11711 (N_11711,N_9299,N_9685);
and U11712 (N_11712,N_8201,N_9109);
nand U11713 (N_11713,N_9067,N_9036);
nor U11714 (N_11714,N_9057,N_9960);
and U11715 (N_11715,N_9537,N_9270);
or U11716 (N_11716,N_8637,N_8581);
nor U11717 (N_11717,N_9360,N_8751);
nor U11718 (N_11718,N_9606,N_9614);
and U11719 (N_11719,N_9443,N_8973);
and U11720 (N_11720,N_8515,N_8234);
nor U11721 (N_11721,N_9355,N_8993);
nor U11722 (N_11722,N_9612,N_8416);
xnor U11723 (N_11723,N_8921,N_8294);
nor U11724 (N_11724,N_9674,N_8995);
or U11725 (N_11725,N_8395,N_9330);
nor U11726 (N_11726,N_9266,N_9319);
nand U11727 (N_11727,N_9532,N_9239);
and U11728 (N_11728,N_9473,N_8327);
nor U11729 (N_11729,N_8110,N_8243);
xnor U11730 (N_11730,N_9920,N_9657);
nand U11731 (N_11731,N_9195,N_8454);
xnor U11732 (N_11732,N_8876,N_9574);
nand U11733 (N_11733,N_8474,N_8071);
and U11734 (N_11734,N_8880,N_9504);
xnor U11735 (N_11735,N_8621,N_9225);
nor U11736 (N_11736,N_9963,N_8158);
or U11737 (N_11737,N_9723,N_9038);
and U11738 (N_11738,N_8137,N_8967);
nand U11739 (N_11739,N_8036,N_8003);
xor U11740 (N_11740,N_8699,N_8170);
xor U11741 (N_11741,N_9008,N_8871);
nand U11742 (N_11742,N_9832,N_8335);
and U11743 (N_11743,N_9064,N_9135);
xor U11744 (N_11744,N_8310,N_9255);
xnor U11745 (N_11745,N_9470,N_9516);
and U11746 (N_11746,N_9212,N_9691);
nor U11747 (N_11747,N_9017,N_9955);
and U11748 (N_11748,N_8570,N_9505);
xnor U11749 (N_11749,N_8801,N_8877);
nor U11750 (N_11750,N_8374,N_8934);
or U11751 (N_11751,N_8848,N_9635);
nand U11752 (N_11752,N_8051,N_9513);
nand U11753 (N_11753,N_8753,N_8099);
or U11754 (N_11754,N_9661,N_9389);
or U11755 (N_11755,N_8921,N_8828);
and U11756 (N_11756,N_8816,N_8826);
nor U11757 (N_11757,N_9015,N_8044);
and U11758 (N_11758,N_8430,N_9370);
or U11759 (N_11759,N_8933,N_8163);
nor U11760 (N_11760,N_9740,N_9283);
xnor U11761 (N_11761,N_9780,N_9179);
or U11762 (N_11762,N_9259,N_8620);
or U11763 (N_11763,N_9499,N_9898);
or U11764 (N_11764,N_8056,N_8104);
or U11765 (N_11765,N_8896,N_9633);
or U11766 (N_11766,N_8617,N_8104);
or U11767 (N_11767,N_8596,N_8264);
xnor U11768 (N_11768,N_9548,N_9140);
and U11769 (N_11769,N_9592,N_9480);
nand U11770 (N_11770,N_8477,N_9332);
or U11771 (N_11771,N_9014,N_8460);
and U11772 (N_11772,N_9685,N_9777);
or U11773 (N_11773,N_8470,N_8917);
and U11774 (N_11774,N_8948,N_8590);
xnor U11775 (N_11775,N_9936,N_9987);
and U11776 (N_11776,N_9255,N_9881);
or U11777 (N_11777,N_8663,N_8246);
xnor U11778 (N_11778,N_8228,N_8299);
nand U11779 (N_11779,N_8937,N_8760);
or U11780 (N_11780,N_8417,N_9240);
nor U11781 (N_11781,N_9703,N_9221);
nand U11782 (N_11782,N_9379,N_8064);
or U11783 (N_11783,N_9203,N_8598);
or U11784 (N_11784,N_9834,N_9197);
and U11785 (N_11785,N_9551,N_9341);
and U11786 (N_11786,N_8485,N_9982);
or U11787 (N_11787,N_9780,N_8585);
xor U11788 (N_11788,N_8912,N_9814);
or U11789 (N_11789,N_9022,N_8179);
nor U11790 (N_11790,N_9754,N_9921);
nor U11791 (N_11791,N_9092,N_9923);
nand U11792 (N_11792,N_8751,N_9321);
and U11793 (N_11793,N_9680,N_8400);
or U11794 (N_11794,N_9545,N_9824);
nor U11795 (N_11795,N_9929,N_9831);
or U11796 (N_11796,N_9681,N_9978);
or U11797 (N_11797,N_9352,N_8759);
nand U11798 (N_11798,N_8799,N_9488);
and U11799 (N_11799,N_8390,N_8379);
nand U11800 (N_11800,N_8070,N_9691);
or U11801 (N_11801,N_9030,N_9421);
xor U11802 (N_11802,N_9467,N_8455);
or U11803 (N_11803,N_9815,N_8657);
nor U11804 (N_11804,N_8364,N_9159);
nor U11805 (N_11805,N_8463,N_9501);
xor U11806 (N_11806,N_8542,N_9440);
and U11807 (N_11807,N_8222,N_8081);
and U11808 (N_11808,N_9758,N_9357);
or U11809 (N_11809,N_9376,N_8129);
or U11810 (N_11810,N_9944,N_8739);
or U11811 (N_11811,N_8164,N_8866);
xnor U11812 (N_11812,N_9013,N_8455);
or U11813 (N_11813,N_8063,N_9000);
nor U11814 (N_11814,N_8422,N_8089);
nand U11815 (N_11815,N_8173,N_9839);
nand U11816 (N_11816,N_9602,N_9913);
xnor U11817 (N_11817,N_8415,N_9336);
or U11818 (N_11818,N_8481,N_8058);
or U11819 (N_11819,N_9366,N_9333);
nand U11820 (N_11820,N_9176,N_9453);
nand U11821 (N_11821,N_8431,N_9642);
xor U11822 (N_11822,N_9321,N_8177);
nor U11823 (N_11823,N_9498,N_8957);
and U11824 (N_11824,N_8416,N_9198);
or U11825 (N_11825,N_9110,N_9323);
xnor U11826 (N_11826,N_8113,N_9385);
nor U11827 (N_11827,N_8908,N_8738);
or U11828 (N_11828,N_9156,N_8278);
nand U11829 (N_11829,N_9436,N_8970);
nand U11830 (N_11830,N_9624,N_9967);
and U11831 (N_11831,N_8175,N_9341);
or U11832 (N_11832,N_9750,N_9775);
and U11833 (N_11833,N_8529,N_8031);
xor U11834 (N_11834,N_8448,N_8782);
xnor U11835 (N_11835,N_9550,N_9320);
and U11836 (N_11836,N_9145,N_8174);
or U11837 (N_11837,N_8601,N_8037);
nand U11838 (N_11838,N_8035,N_9402);
nand U11839 (N_11839,N_9179,N_8734);
and U11840 (N_11840,N_8371,N_9161);
xor U11841 (N_11841,N_8044,N_8377);
nor U11842 (N_11842,N_9707,N_9840);
xor U11843 (N_11843,N_9996,N_9272);
and U11844 (N_11844,N_8299,N_9916);
and U11845 (N_11845,N_8198,N_8637);
or U11846 (N_11846,N_9456,N_9964);
and U11847 (N_11847,N_9291,N_8660);
xnor U11848 (N_11848,N_8724,N_9387);
or U11849 (N_11849,N_9532,N_8420);
or U11850 (N_11850,N_8114,N_9380);
nor U11851 (N_11851,N_8678,N_8888);
nor U11852 (N_11852,N_8341,N_9372);
and U11853 (N_11853,N_9030,N_8275);
or U11854 (N_11854,N_9478,N_9569);
xnor U11855 (N_11855,N_9620,N_9189);
nor U11856 (N_11856,N_9755,N_8163);
nor U11857 (N_11857,N_9598,N_9593);
nor U11858 (N_11858,N_9289,N_9007);
nor U11859 (N_11859,N_9071,N_9189);
nor U11860 (N_11860,N_8574,N_8591);
or U11861 (N_11861,N_8405,N_8324);
or U11862 (N_11862,N_8621,N_8644);
xnor U11863 (N_11863,N_9297,N_9242);
nand U11864 (N_11864,N_8302,N_8211);
or U11865 (N_11865,N_9530,N_8691);
and U11866 (N_11866,N_9293,N_8857);
or U11867 (N_11867,N_9579,N_9202);
nand U11868 (N_11868,N_8222,N_9350);
and U11869 (N_11869,N_8836,N_9620);
nor U11870 (N_11870,N_9905,N_9530);
nor U11871 (N_11871,N_8375,N_9440);
or U11872 (N_11872,N_9146,N_8415);
nor U11873 (N_11873,N_8415,N_8132);
and U11874 (N_11874,N_8721,N_9417);
or U11875 (N_11875,N_8318,N_8386);
or U11876 (N_11876,N_8519,N_9237);
and U11877 (N_11877,N_8111,N_8395);
xnor U11878 (N_11878,N_9194,N_8371);
nor U11879 (N_11879,N_9334,N_8229);
nor U11880 (N_11880,N_8452,N_9100);
xor U11881 (N_11881,N_9749,N_8812);
or U11882 (N_11882,N_8926,N_8803);
or U11883 (N_11883,N_9757,N_9597);
nor U11884 (N_11884,N_8249,N_9486);
and U11885 (N_11885,N_9418,N_8796);
xor U11886 (N_11886,N_8416,N_8826);
and U11887 (N_11887,N_8199,N_9177);
and U11888 (N_11888,N_8299,N_9271);
or U11889 (N_11889,N_9702,N_8401);
nand U11890 (N_11890,N_9809,N_8428);
and U11891 (N_11891,N_8467,N_8083);
xor U11892 (N_11892,N_8673,N_9207);
xor U11893 (N_11893,N_8074,N_8380);
and U11894 (N_11894,N_9215,N_8072);
nor U11895 (N_11895,N_9533,N_8061);
nor U11896 (N_11896,N_8549,N_9434);
xnor U11897 (N_11897,N_9329,N_8582);
xor U11898 (N_11898,N_8198,N_9721);
or U11899 (N_11899,N_8207,N_8858);
xnor U11900 (N_11900,N_8824,N_8778);
xnor U11901 (N_11901,N_9527,N_8311);
nand U11902 (N_11902,N_9192,N_9417);
and U11903 (N_11903,N_9928,N_8671);
nand U11904 (N_11904,N_9820,N_9251);
xnor U11905 (N_11905,N_9776,N_8824);
nor U11906 (N_11906,N_8266,N_9249);
or U11907 (N_11907,N_8403,N_8215);
and U11908 (N_11908,N_9593,N_9040);
nand U11909 (N_11909,N_9700,N_8441);
xor U11910 (N_11910,N_8807,N_8292);
nor U11911 (N_11911,N_9481,N_8509);
and U11912 (N_11912,N_8744,N_8508);
and U11913 (N_11913,N_9726,N_9365);
nor U11914 (N_11914,N_9031,N_9210);
nor U11915 (N_11915,N_8729,N_9629);
nor U11916 (N_11916,N_9002,N_8010);
xor U11917 (N_11917,N_9942,N_9713);
and U11918 (N_11918,N_8586,N_8504);
xor U11919 (N_11919,N_8916,N_8634);
or U11920 (N_11920,N_9796,N_9257);
xnor U11921 (N_11921,N_9916,N_9424);
nor U11922 (N_11922,N_8116,N_9562);
xnor U11923 (N_11923,N_8613,N_9545);
nand U11924 (N_11924,N_8674,N_9006);
nand U11925 (N_11925,N_9898,N_8184);
nand U11926 (N_11926,N_9274,N_8958);
nor U11927 (N_11927,N_8847,N_9170);
xor U11928 (N_11928,N_9981,N_9451);
nand U11929 (N_11929,N_9658,N_9753);
or U11930 (N_11930,N_9761,N_9532);
nand U11931 (N_11931,N_9468,N_9542);
xor U11932 (N_11932,N_8759,N_9556);
or U11933 (N_11933,N_9081,N_8726);
or U11934 (N_11934,N_9323,N_8177);
nand U11935 (N_11935,N_9569,N_8965);
nor U11936 (N_11936,N_8214,N_9040);
nor U11937 (N_11937,N_8744,N_9192);
xnor U11938 (N_11938,N_9341,N_8962);
and U11939 (N_11939,N_8956,N_8131);
xor U11940 (N_11940,N_9559,N_9755);
xor U11941 (N_11941,N_9912,N_8185);
nor U11942 (N_11942,N_8104,N_8005);
xor U11943 (N_11943,N_8179,N_8506);
and U11944 (N_11944,N_9408,N_8571);
xor U11945 (N_11945,N_9056,N_9292);
nor U11946 (N_11946,N_9582,N_9350);
nand U11947 (N_11947,N_8935,N_9462);
nand U11948 (N_11948,N_8453,N_8243);
nand U11949 (N_11949,N_8898,N_9772);
nor U11950 (N_11950,N_9177,N_9505);
and U11951 (N_11951,N_9122,N_9638);
xnor U11952 (N_11952,N_8778,N_8191);
nor U11953 (N_11953,N_8198,N_9746);
nand U11954 (N_11954,N_8451,N_9522);
xnor U11955 (N_11955,N_9487,N_8310);
and U11956 (N_11956,N_9310,N_9456);
nor U11957 (N_11957,N_8495,N_8887);
and U11958 (N_11958,N_8202,N_8935);
and U11959 (N_11959,N_9268,N_9541);
nand U11960 (N_11960,N_9831,N_9600);
nand U11961 (N_11961,N_9857,N_9623);
and U11962 (N_11962,N_9188,N_9652);
and U11963 (N_11963,N_9263,N_8256);
nand U11964 (N_11964,N_9362,N_8881);
and U11965 (N_11965,N_8756,N_9043);
nand U11966 (N_11966,N_8191,N_8368);
or U11967 (N_11967,N_8583,N_8663);
xor U11968 (N_11968,N_8604,N_9562);
or U11969 (N_11969,N_9186,N_8698);
nor U11970 (N_11970,N_8471,N_8138);
or U11971 (N_11971,N_9720,N_9546);
and U11972 (N_11972,N_9474,N_8590);
and U11973 (N_11973,N_8265,N_8176);
xnor U11974 (N_11974,N_9351,N_8356);
nand U11975 (N_11975,N_8738,N_8728);
xor U11976 (N_11976,N_9636,N_9039);
nor U11977 (N_11977,N_8540,N_8326);
nand U11978 (N_11978,N_8695,N_8015);
and U11979 (N_11979,N_9497,N_8148);
xor U11980 (N_11980,N_8464,N_9812);
or U11981 (N_11981,N_9095,N_9416);
and U11982 (N_11982,N_9592,N_9607);
and U11983 (N_11983,N_9202,N_8735);
nor U11984 (N_11984,N_8107,N_8075);
xor U11985 (N_11985,N_9184,N_9035);
nor U11986 (N_11986,N_8992,N_9846);
or U11987 (N_11987,N_9689,N_9164);
nor U11988 (N_11988,N_8235,N_8257);
and U11989 (N_11989,N_8707,N_8425);
xnor U11990 (N_11990,N_8516,N_9246);
xor U11991 (N_11991,N_8520,N_9244);
nand U11992 (N_11992,N_8769,N_9746);
nor U11993 (N_11993,N_8071,N_8743);
and U11994 (N_11994,N_8737,N_8545);
nor U11995 (N_11995,N_8683,N_9286);
or U11996 (N_11996,N_8075,N_8959);
nor U11997 (N_11997,N_9495,N_9468);
nand U11998 (N_11998,N_8676,N_9366);
nor U11999 (N_11999,N_9811,N_9204);
xnor U12000 (N_12000,N_11444,N_11045);
and U12001 (N_12001,N_10222,N_10957);
or U12002 (N_12002,N_10435,N_11244);
and U12003 (N_12003,N_11415,N_10448);
xor U12004 (N_12004,N_11395,N_11913);
nor U12005 (N_12005,N_11915,N_11471);
and U12006 (N_12006,N_11731,N_11636);
xnor U12007 (N_12007,N_11130,N_11073);
nand U12008 (N_12008,N_10889,N_10795);
nor U12009 (N_12009,N_10644,N_11393);
xnor U12010 (N_12010,N_11786,N_11339);
nand U12011 (N_12011,N_10445,N_11310);
xor U12012 (N_12012,N_11533,N_11246);
or U12013 (N_12013,N_10293,N_10755);
nor U12014 (N_12014,N_11142,N_10354);
nor U12015 (N_12015,N_10211,N_11753);
xnor U12016 (N_12016,N_10618,N_10616);
xor U12017 (N_12017,N_10074,N_11080);
or U12018 (N_12018,N_11576,N_11314);
nand U12019 (N_12019,N_10463,N_10377);
and U12020 (N_12020,N_10600,N_11494);
xnor U12021 (N_12021,N_10011,N_11043);
nor U12022 (N_12022,N_10469,N_10754);
or U12023 (N_12023,N_10573,N_11564);
or U12024 (N_12024,N_10908,N_11265);
nor U12025 (N_12025,N_11202,N_11209);
nor U12026 (N_12026,N_11441,N_11146);
and U12027 (N_12027,N_11428,N_11040);
and U12028 (N_12028,N_10916,N_10749);
xnor U12029 (N_12029,N_10457,N_10997);
nor U12030 (N_12030,N_11143,N_11994);
nand U12031 (N_12031,N_10582,N_11907);
or U12032 (N_12032,N_10349,N_10675);
or U12033 (N_12033,N_10687,N_11610);
and U12034 (N_12034,N_10715,N_10841);
or U12035 (N_12035,N_11443,N_11463);
xor U12036 (N_12036,N_10289,N_10932);
nand U12037 (N_12037,N_10054,N_11817);
nor U12038 (N_12038,N_10096,N_10766);
or U12039 (N_12039,N_11460,N_10652);
nand U12040 (N_12040,N_11848,N_11057);
nand U12041 (N_12041,N_10962,N_11120);
xnor U12042 (N_12042,N_11792,N_11135);
xnor U12043 (N_12043,N_11717,N_10295);
or U12044 (N_12044,N_11740,N_10802);
nand U12045 (N_12045,N_11276,N_10403);
or U12046 (N_12046,N_11149,N_10956);
and U12047 (N_12047,N_10868,N_11237);
xor U12048 (N_12048,N_11331,N_10839);
nand U12049 (N_12049,N_10106,N_11936);
or U12050 (N_12050,N_10746,N_10093);
nor U12051 (N_12051,N_11614,N_11499);
xnor U12052 (N_12052,N_11843,N_10659);
and U12053 (N_12053,N_11264,N_10676);
or U12054 (N_12054,N_10039,N_11802);
nor U12055 (N_12055,N_11206,N_10725);
and U12056 (N_12056,N_11529,N_11230);
or U12057 (N_12057,N_10982,N_10660);
or U12058 (N_12058,N_10171,N_10152);
and U12059 (N_12059,N_11249,N_10420);
nand U12060 (N_12060,N_11097,N_11170);
or U12061 (N_12061,N_10155,N_10735);
nor U12062 (N_12062,N_11302,N_10869);
and U12063 (N_12063,N_11183,N_10258);
xor U12064 (N_12064,N_11855,N_10200);
and U12065 (N_12065,N_10433,N_10645);
or U12066 (N_12066,N_11739,N_11211);
xor U12067 (N_12067,N_10043,N_11758);
and U12068 (N_12068,N_11814,N_10127);
xnor U12069 (N_12069,N_10845,N_10415);
nor U12070 (N_12070,N_10462,N_10977);
and U12071 (N_12071,N_10847,N_10124);
nand U12072 (N_12072,N_11121,N_11323);
xnor U12073 (N_12073,N_10928,N_11841);
nand U12074 (N_12074,N_11436,N_10713);
xnor U12075 (N_12075,N_11354,N_10452);
nand U12076 (N_12076,N_11970,N_11932);
nand U12077 (N_12077,N_11307,N_10584);
xnor U12078 (N_12078,N_11705,N_11100);
or U12079 (N_12079,N_11019,N_10595);
nand U12080 (N_12080,N_11693,N_10721);
or U12081 (N_12081,N_11110,N_11447);
xor U12082 (N_12082,N_10282,N_10743);
nor U12083 (N_12083,N_10995,N_11222);
nor U12084 (N_12084,N_10070,N_11001);
nor U12085 (N_12085,N_11488,N_11173);
nor U12086 (N_12086,N_10164,N_10303);
xor U12087 (N_12087,N_11596,N_10590);
nand U12088 (N_12088,N_10213,N_11965);
and U12089 (N_12089,N_10261,N_10064);
or U12090 (N_12090,N_10234,N_10712);
and U12091 (N_12091,N_10207,N_11945);
xnor U12092 (N_12092,N_10091,N_10084);
nor U12093 (N_12093,N_11652,N_11710);
and U12094 (N_12094,N_11526,N_11150);
nor U12095 (N_12095,N_10035,N_11939);
nand U12096 (N_12096,N_10414,N_10820);
and U12097 (N_12097,N_10188,N_11383);
xnor U12098 (N_12098,N_10671,N_10292);
xnor U12099 (N_12099,N_11165,N_10972);
nand U12100 (N_12100,N_11303,N_11096);
and U12101 (N_12101,N_10505,N_10895);
xor U12102 (N_12102,N_10009,N_10203);
nand U12103 (N_12103,N_11726,N_11585);
xnor U12104 (N_12104,N_11182,N_11122);
xnor U12105 (N_12105,N_11766,N_10422);
nand U12106 (N_12106,N_11133,N_11708);
and U12107 (N_12107,N_10384,N_11741);
xor U12108 (N_12108,N_10513,N_10340);
xnor U12109 (N_12109,N_10430,N_11508);
or U12110 (N_12110,N_11951,N_10148);
or U12111 (N_12111,N_10413,N_11257);
or U12112 (N_12112,N_11933,N_11995);
and U12113 (N_12113,N_10287,N_10739);
or U12114 (N_12114,N_11125,N_11049);
or U12115 (N_12115,N_11525,N_11520);
nand U12116 (N_12116,N_10036,N_10242);
or U12117 (N_12117,N_10767,N_11860);
xnor U12118 (N_12118,N_11634,N_11485);
nor U12119 (N_12119,N_11558,N_11159);
or U12120 (N_12120,N_11947,N_11465);
or U12121 (N_12121,N_11335,N_11926);
nor U12122 (N_12122,N_10611,N_10664);
nand U12123 (N_12123,N_11899,N_10855);
or U12124 (N_12124,N_10619,N_11824);
or U12125 (N_12125,N_10232,N_10756);
nor U12126 (N_12126,N_11891,N_10110);
and U12127 (N_12127,N_10197,N_11002);
nor U12128 (N_12128,N_10807,N_11780);
nor U12129 (N_12129,N_11200,N_11538);
and U12130 (N_12130,N_11176,N_10734);
nand U12131 (N_12131,N_10459,N_11114);
xor U12132 (N_12132,N_11836,N_11338);
nand U12133 (N_12133,N_10753,N_11623);
xor U12134 (N_12134,N_10166,N_11111);
and U12135 (N_12135,N_10192,N_11190);
and U12136 (N_12136,N_10466,N_11104);
or U12137 (N_12137,N_11233,N_11458);
or U12138 (N_12138,N_11232,N_10798);
xor U12139 (N_12139,N_11999,N_11702);
nor U12140 (N_12140,N_11734,N_11448);
nor U12141 (N_12141,N_11388,N_10714);
xor U12142 (N_12142,N_10313,N_11643);
or U12143 (N_12143,N_11470,N_10708);
nor U12144 (N_12144,N_10720,N_10129);
and U12145 (N_12145,N_11506,N_11501);
xnor U12146 (N_12146,N_11827,N_11664);
nor U12147 (N_12147,N_11369,N_11409);
and U12148 (N_12148,N_10131,N_10477);
nand U12149 (N_12149,N_11069,N_10539);
or U12150 (N_12150,N_11648,N_10780);
nor U12151 (N_12151,N_10220,N_10794);
and U12152 (N_12152,N_10602,N_11703);
xnor U12153 (N_12153,N_11723,N_11489);
or U12154 (N_12154,N_10711,N_10160);
xnor U12155 (N_12155,N_10575,N_11810);
and U12156 (N_12156,N_10126,N_10971);
and U12157 (N_12157,N_11832,N_11955);
or U12158 (N_12158,N_11351,N_11280);
nand U12159 (N_12159,N_10964,N_11322);
nor U12160 (N_12160,N_10389,N_10812);
xnor U12161 (N_12161,N_11025,N_11577);
xor U12162 (N_12162,N_10813,N_11737);
and U12163 (N_12163,N_10394,N_11086);
nand U12164 (N_12164,N_10731,N_11895);
and U12165 (N_12165,N_11884,N_10880);
and U12166 (N_12166,N_10874,N_11451);
or U12167 (N_12167,N_11980,N_11414);
and U12168 (N_12168,N_10598,N_11851);
nor U12169 (N_12169,N_11886,N_11628);
nand U12170 (N_12170,N_11006,N_11433);
nor U12171 (N_12171,N_11658,N_11132);
nor U12172 (N_12172,N_11145,N_11361);
or U12173 (N_12173,N_10509,N_11192);
nand U12174 (N_12174,N_10046,N_11888);
nor U12175 (N_12175,N_10680,N_10073);
nor U12176 (N_12176,N_10159,N_11603);
nor U12177 (N_12177,N_11271,N_10861);
xnor U12178 (N_12178,N_11712,N_11781);
xnor U12179 (N_12179,N_11897,N_10274);
or U12180 (N_12180,N_10216,N_11517);
nor U12181 (N_12181,N_10305,N_11290);
nand U12182 (N_12182,N_11730,N_11553);
nand U12183 (N_12183,N_10272,N_10085);
nand U12184 (N_12184,N_10507,N_10641);
and U12185 (N_12185,N_10117,N_10737);
nor U12186 (N_12186,N_10773,N_11337);
or U12187 (N_12187,N_10467,N_11055);
nand U12188 (N_12188,N_10386,N_11608);
or U12189 (N_12189,N_11692,N_11277);
nor U12190 (N_12190,N_11226,N_11287);
nor U12191 (N_12191,N_10699,N_10759);
nor U12192 (N_12192,N_11358,N_11735);
nand U12193 (N_12193,N_11949,N_10239);
and U12194 (N_12194,N_10760,N_11665);
nand U12195 (N_12195,N_10314,N_10399);
xnor U12196 (N_12196,N_10730,N_10989);
nand U12197 (N_12197,N_11456,N_11992);
and U12198 (N_12198,N_11185,N_10361);
or U12199 (N_12199,N_10194,N_11340);
nor U12200 (N_12200,N_11243,N_10633);
and U12201 (N_12201,N_11124,N_11597);
nor U12202 (N_12202,N_11467,N_11738);
xor U12203 (N_12203,N_10105,N_10825);
nor U12204 (N_12204,N_10331,N_10439);
or U12205 (N_12205,N_10661,N_10534);
nand U12206 (N_12206,N_11203,N_11207);
and U12207 (N_12207,N_11656,N_11591);
and U12208 (N_12208,N_11342,N_11716);
nor U12209 (N_12209,N_11026,N_10357);
xnor U12210 (N_12210,N_10072,N_11675);
xnor U12211 (N_12211,N_10873,N_11707);
and U12212 (N_12212,N_11912,N_11650);
and U12213 (N_12213,N_10960,N_10592);
or U12214 (N_12214,N_11077,N_10623);
nand U12215 (N_12215,N_10373,N_11733);
and U12216 (N_12216,N_11474,N_11695);
nor U12217 (N_12217,N_11399,N_10921);
nand U12218 (N_12218,N_11906,N_11773);
nand U12219 (N_12219,N_11959,N_11497);
nor U12220 (N_12220,N_10900,N_10481);
xnor U12221 (N_12221,N_10089,N_11205);
xor U12222 (N_12222,N_11437,N_11898);
nor U12223 (N_12223,N_11362,N_10934);
nor U12224 (N_12224,N_10887,N_10020);
nand U12225 (N_12225,N_10913,N_11350);
or U12226 (N_12226,N_10284,N_10175);
and U12227 (N_12227,N_11957,N_10271);
or U12228 (N_12228,N_11106,N_10180);
xor U12229 (N_12229,N_11262,N_11224);
xnor U12230 (N_12230,N_10961,N_10102);
xnor U12231 (N_12231,N_11548,N_10770);
nor U12232 (N_12232,N_10267,N_10352);
and U12233 (N_12233,N_10973,N_10029);
or U12234 (N_12234,N_11820,N_11327);
and U12235 (N_12235,N_11540,N_10917);
xnor U12236 (N_12236,N_10844,N_11425);
xor U12237 (N_12237,N_10436,N_10034);
xor U12238 (N_12238,N_10526,N_10547);
or U12239 (N_12239,N_11927,N_11727);
nor U12240 (N_12240,N_11438,N_11498);
xor U12241 (N_12241,N_11682,N_10483);
nor U12242 (N_12242,N_10495,N_10364);
or U12243 (N_12243,N_11245,N_10134);
nor U12244 (N_12244,N_11154,N_11946);
or U12245 (N_12245,N_11059,N_10083);
nor U12246 (N_12246,N_11539,N_10473);
xor U12247 (N_12247,N_11248,N_10028);
nand U12248 (N_12248,N_11390,N_11366);
and U12249 (N_12249,N_10974,N_10543);
nor U12250 (N_12250,N_10022,N_11023);
nor U12251 (N_12251,N_11070,N_11584);
nor U12252 (N_12252,N_10503,N_11619);
and U12253 (N_12253,N_11866,N_10922);
or U12254 (N_12254,N_10051,N_11819);
or U12255 (N_12255,N_10980,N_10589);
or U12256 (N_12256,N_10338,N_10886);
and U12257 (N_12257,N_10324,N_11213);
or U12258 (N_12258,N_10008,N_10062);
nor U12259 (N_12259,N_10706,N_11536);
nor U12260 (N_12260,N_10943,N_11177);
and U12261 (N_12261,N_11089,N_11424);
nor U12262 (N_12262,N_10252,N_10648);
or U12263 (N_12263,N_11904,N_11223);
nor U12264 (N_12264,N_10401,N_11285);
or U12265 (N_12265,N_11775,N_11621);
xnor U12266 (N_12266,N_11732,N_11071);
nor U12267 (N_12267,N_10821,N_11941);
nor U12268 (N_12268,N_11381,N_10642);
or U12269 (N_12269,N_11861,N_10410);
or U12270 (N_12270,N_11782,N_10094);
nand U12271 (N_12271,N_10210,N_10061);
xnor U12272 (N_12272,N_10967,N_10925);
or U12273 (N_12273,N_10907,N_11627);
xnor U12274 (N_12274,N_11326,N_11403);
nand U12275 (N_12275,N_11446,N_10638);
xor U12276 (N_12276,N_11432,N_10214);
nand U12277 (N_12277,N_10285,N_10854);
nor U12278 (N_12278,N_10275,N_10850);
nor U12279 (N_12279,N_11996,N_11178);
xor U12280 (N_12280,N_10787,N_11127);
nand U12281 (N_12281,N_11639,N_11058);
nand U12282 (N_12282,N_10681,N_11027);
or U12283 (N_12283,N_11098,N_11968);
nand U12284 (N_12284,N_11943,N_10360);
nor U12285 (N_12285,N_11147,N_10601);
and U12286 (N_12286,N_10692,N_11197);
nor U12287 (N_12287,N_11210,N_10992);
and U12288 (N_12288,N_11477,N_11806);
or U12289 (N_12289,N_10793,N_11763);
nor U12290 (N_12290,N_10947,N_11850);
and U12291 (N_12291,N_10451,N_11566);
and U12292 (N_12292,N_11598,N_11760);
or U12293 (N_12293,N_11751,N_10443);
and U12294 (N_12294,N_11632,N_10751);
or U12295 (N_12295,N_11099,N_11954);
or U12296 (N_12296,N_11373,N_10255);
or U12297 (N_12297,N_11622,N_10783);
and U12298 (N_12298,N_10550,N_10882);
or U12299 (N_12299,N_10668,N_11768);
nor U12300 (N_12300,N_10165,N_11484);
nand U12301 (N_12301,N_11048,N_10672);
nand U12302 (N_12302,N_11486,N_11605);
and U12303 (N_12303,N_11604,N_11989);
and U12304 (N_12304,N_10649,N_11807);
nand U12305 (N_12305,N_10017,N_10914);
nand U12306 (N_12306,N_10178,N_11718);
nor U12307 (N_12307,N_11567,N_10639);
or U12308 (N_12308,N_11667,N_10518);
nand U12309 (N_12309,N_10883,N_10111);
xnor U12310 (N_12310,N_10000,N_11826);
or U12311 (N_12311,N_11266,N_11595);
nor U12312 (N_12312,N_10390,N_10496);
nand U12313 (N_12313,N_10350,N_10704);
nor U12314 (N_12314,N_10149,N_10497);
nor U12315 (N_12315,N_11549,N_10741);
and U12316 (N_12316,N_10270,N_11053);
or U12317 (N_12317,N_10524,N_10818);
xnor U12318 (N_12318,N_11215,N_11016);
xor U12319 (N_12319,N_11160,N_11208);
xnor U12320 (N_12320,N_11316,N_11199);
nor U12321 (N_12321,N_10673,N_11301);
or U12322 (N_12322,N_11583,N_10190);
nand U12323 (N_12323,N_11082,N_11005);
nor U12324 (N_12324,N_10571,N_11075);
nor U12325 (N_12325,N_11227,N_10201);
and U12326 (N_12326,N_11445,N_11812);
xor U12327 (N_12327,N_10878,N_11187);
nor U12328 (N_12328,N_11831,N_10315);
and U12329 (N_12329,N_11606,N_10612);
xor U12330 (N_12330,N_10183,N_11638);
nor U12331 (N_12331,N_10815,N_10221);
and U12332 (N_12332,N_10341,N_10750);
and U12333 (N_12333,N_10263,N_11123);
and U12334 (N_12334,N_10247,N_11309);
and U12335 (N_12335,N_11914,N_10556);
nor U12336 (N_12336,N_11618,N_10304);
nor U12337 (N_12337,N_10891,N_10736);
nand U12338 (N_12338,N_11166,N_11808);
and U12339 (N_12339,N_10437,N_11715);
nand U12340 (N_12340,N_10309,N_10257);
nand U12341 (N_12341,N_11570,N_10139);
xnor U12342 (N_12342,N_11278,N_10256);
nor U12343 (N_12343,N_10470,N_10187);
xor U12344 (N_12344,N_10005,N_10343);
and U12345 (N_12345,N_11803,N_10808);
or U12346 (N_12346,N_10748,N_11565);
and U12347 (N_12347,N_11672,N_11364);
and U12348 (N_12348,N_11126,N_11937);
nand U12349 (N_12349,N_11527,N_11789);
and U12350 (N_12350,N_10297,N_10196);
xor U12351 (N_12351,N_11261,N_11236);
nand U12352 (N_12352,N_11204,N_10366);
or U12353 (N_12353,N_11919,N_11341);
nor U12354 (N_12354,N_10635,N_11218);
nand U12355 (N_12355,N_11683,N_11374);
nor U12356 (N_12356,N_11318,N_11902);
or U12357 (N_12357,N_11985,N_10594);
or U12358 (N_12358,N_11181,N_11518);
and U12359 (N_12359,N_10141,N_11516);
nand U12360 (N_12360,N_11599,N_11167);
nand U12361 (N_12361,N_10682,N_11776);
nor U12362 (N_12362,N_10732,N_11095);
nand U12363 (N_12363,N_10041,N_10336);
or U12364 (N_12364,N_10065,N_11252);
nand U12365 (N_12365,N_10788,N_11201);
nand U12366 (N_12366,N_10701,N_10519);
and U12367 (N_12367,N_10156,N_11896);
and U12368 (N_12368,N_11876,N_10049);
and U12369 (N_12369,N_11010,N_11018);
and U12370 (N_12370,N_11713,N_10674);
nor U12371 (N_12371,N_10689,N_11091);
nor U12372 (N_12372,N_11637,N_10050);
xnor U12373 (N_12373,N_11856,N_10015);
and U12374 (N_12374,N_10945,N_11039);
or U12375 (N_12375,N_11616,N_10525);
or U12376 (N_12376,N_11511,N_10488);
nor U12377 (N_12377,N_10060,N_10176);
xor U12378 (N_12378,N_10599,N_10407);
nand U12379 (N_12379,N_10940,N_11816);
nand U12380 (N_12380,N_10132,N_10351);
or U12381 (N_12381,N_10378,N_10605);
and U12382 (N_12382,N_11028,N_10078);
nand U12383 (N_12383,N_11908,N_11171);
nor U12384 (N_12384,N_10388,N_10245);
or U12385 (N_12385,N_11847,N_10108);
xor U12386 (N_12386,N_10076,N_10241);
xnor U12387 (N_12387,N_11311,N_11649);
nor U12388 (N_12388,N_11429,N_10764);
nand U12389 (N_12389,N_11701,N_11960);
xor U12390 (N_12390,N_10137,N_11778);
nor U12391 (N_12391,N_11587,N_11944);
and U12392 (N_12392,N_11845,N_10658);
nand U12393 (N_12393,N_11988,N_10321);
nor U12394 (N_12394,N_11483,N_11743);
xnor U12395 (N_12395,N_10333,N_10266);
nand U12396 (N_12396,N_10607,N_11535);
or U12397 (N_12397,N_11544,N_11853);
nor U12398 (N_12398,N_10702,N_11887);
nor U12399 (N_12399,N_11813,N_10935);
or U12400 (N_12400,N_11214,N_10740);
nor U12401 (N_12401,N_11893,N_11042);
nor U12402 (N_12402,N_10686,N_11212);
nor U12403 (N_12403,N_10248,N_11983);
and U12404 (N_12404,N_10849,N_11569);
xor U12405 (N_12405,N_10100,N_11690);
nand U12406 (N_12406,N_10233,N_11973);
nand U12407 (N_12407,N_10586,N_11882);
and U12408 (N_12408,N_10071,N_11552);
and U12409 (N_12409,N_11993,N_10244);
nor U12410 (N_12410,N_10797,N_11346);
or U12411 (N_12411,N_11537,N_10606);
and U12412 (N_12412,N_11347,N_11607);
and U12413 (N_12413,N_11825,N_11797);
and U12414 (N_12414,N_10508,N_10262);
xor U12415 (N_12415,N_11481,N_11515);
or U12416 (N_12416,N_10742,N_10717);
nor U12417 (N_12417,N_10792,N_11653);
xnor U12418 (N_12418,N_11950,N_11297);
nand U12419 (N_12419,N_11334,N_10032);
nand U12420 (N_12420,N_10195,N_10569);
nor U12421 (N_12421,N_10938,N_10450);
and U12422 (N_12422,N_11295,N_11925);
nand U12423 (N_12423,N_10796,N_10016);
or U12424 (N_12424,N_10814,N_10727);
and U12425 (N_12425,N_10225,N_11367);
and U12426 (N_12426,N_10565,N_11263);
xnor U12427 (N_12427,N_11629,N_11063);
and U12428 (N_12428,N_11240,N_10118);
nand U12429 (N_12429,N_11066,N_11052);
nor U12430 (N_12430,N_11380,N_11298);
and U12431 (N_12431,N_11811,N_10707);
xor U12432 (N_12432,N_11697,N_10561);
or U12433 (N_12433,N_10958,N_11699);
or U12434 (N_12434,N_10970,N_11356);
and U12435 (N_12435,N_10030,N_11034);
nand U12436 (N_12436,N_11956,N_10208);
and U12437 (N_12437,N_11044,N_11714);
or U12438 (N_12438,N_11355,N_10951);
nand U12439 (N_12439,N_10905,N_10955);
and U12440 (N_12440,N_11777,N_10291);
nor U12441 (N_12441,N_11920,N_11416);
nand U12442 (N_12442,N_10294,N_10426);
nand U12443 (N_12443,N_10944,N_10622);
nor U12444 (N_12444,N_10987,N_10809);
nand U12445 (N_12445,N_11435,N_10722);
or U12446 (N_12446,N_11102,N_10348);
nor U12447 (N_12447,N_10710,N_10237);
and U12448 (N_12448,N_10901,N_11910);
xnor U12449 (N_12449,N_10185,N_10493);
nand U12450 (N_12450,N_11241,N_10299);
nand U12451 (N_12451,N_10002,N_10918);
nand U12452 (N_12452,N_11296,N_11007);
and U12453 (N_12453,N_10230,N_10816);
nor U12454 (N_12454,N_11952,N_11784);
nand U12455 (N_12455,N_10238,N_11804);
and U12456 (N_12456,N_10359,N_11449);
nor U12457 (N_12457,N_11575,N_11461);
or U12458 (N_12458,N_10608,N_11559);
xnor U12459 (N_12459,N_11796,N_10651);
and U12460 (N_12460,N_11343,N_10738);
xor U12461 (N_12461,N_11455,N_11854);
xnor U12462 (N_12462,N_11427,N_10830);
or U12463 (N_12463,N_11004,N_11491);
or U12464 (N_12464,N_11815,N_11017);
or U12465 (N_12465,N_11094,N_11514);
and U12466 (N_12466,N_11074,N_11958);
nand U12467 (N_12467,N_10438,N_11869);
and U12468 (N_12468,N_10993,N_11376);
nor U12469 (N_12469,N_10217,N_10963);
or U12470 (N_12470,N_10975,N_10548);
or U12471 (N_12471,N_11586,N_10829);
or U12472 (N_12472,N_10425,N_11858);
nor U12473 (N_12473,N_10828,N_10824);
nand U12474 (N_12474,N_11163,N_11156);
xor U12475 (N_12475,N_10075,N_10574);
nor U12476 (N_12476,N_10991,N_11384);
nor U12477 (N_12477,N_10647,N_11875);
nand U12478 (N_12478,N_10339,N_10719);
xnor U12479 (N_12479,N_10231,N_10610);
xor U12480 (N_12480,N_10578,N_11431);
xnor U12481 (N_12481,N_11169,N_10236);
xnor U12482 (N_12482,N_11523,N_11408);
and U12483 (N_12483,N_11589,N_10475);
nor U12484 (N_12484,N_11308,N_11375);
or U12485 (N_12485,N_11279,N_11188);
nor U12486 (N_12486,N_11291,N_11195);
nor U12487 (N_12487,N_10894,N_11709);
xor U12488 (N_12488,N_11021,N_11267);
or U12489 (N_12489,N_10931,N_10976);
and U12490 (N_12490,N_10052,N_11545);
xor U12491 (N_12491,N_10374,N_11251);
nor U12492 (N_12492,N_11986,N_10662);
or U12493 (N_12493,N_10498,N_11054);
or U12494 (N_12494,N_10540,N_10512);
nor U12495 (N_12495,N_11088,N_10862);
nor U12496 (N_12496,N_11631,N_11273);
xnor U12497 (N_12497,N_11711,N_11987);
or U12498 (N_12498,N_10206,N_10580);
and U12499 (N_12499,N_10223,N_11754);
or U12500 (N_12500,N_10409,N_10936);
and U12501 (N_12501,N_11056,N_10521);
nand U12502 (N_12502,N_10881,N_10915);
nor U12503 (N_12503,N_10650,N_10801);
or U12504 (N_12504,N_11401,N_10308);
xnor U12505 (N_12505,N_11398,N_10082);
and U12506 (N_12506,N_11761,N_11592);
nor U12507 (N_12507,N_11736,N_11547);
xor U12508 (N_12508,N_11818,N_11676);
and U12509 (N_12509,N_10228,N_10460);
nand U12510 (N_12510,N_11368,N_11180);
or U12511 (N_12511,N_10246,N_10968);
nand U12512 (N_12512,N_10986,N_10226);
or U12513 (N_12513,N_10520,N_10202);
or U12514 (N_12514,N_11971,N_11281);
and U12515 (N_12515,N_11020,N_11269);
and U12516 (N_12516,N_11141,N_11293);
nor U12517 (N_12517,N_10781,N_10107);
and U12518 (N_12518,N_10122,N_11581);
and U12519 (N_12519,N_11228,N_11392);
or U12520 (N_12520,N_11008,N_10380);
nor U12521 (N_12521,N_11928,N_11640);
and U12522 (N_12522,N_11153,N_11967);
xnor U12523 (N_12523,N_10570,N_10001);
or U12524 (N_12524,N_11883,N_11571);
or U12525 (N_12525,N_10310,N_11242);
xor U12526 (N_12526,N_11885,N_10040);
and U12527 (N_12527,N_10479,N_10038);
nor U12528 (N_12528,N_10670,N_11642);
and U12529 (N_12529,N_10444,N_10066);
or U12530 (N_12530,N_11344,N_10365);
nand U12531 (N_12531,N_10836,N_11580);
nand U12532 (N_12532,N_11462,N_10863);
and U12533 (N_12533,N_10092,N_11868);
nand U12534 (N_12534,N_11659,N_10342);
and U12535 (N_12535,N_10597,N_10551);
or U12536 (N_12536,N_10157,N_11493);
and U12537 (N_12537,N_10006,N_11609);
or U12538 (N_12538,N_11757,N_11829);
nand U12539 (N_12539,N_10871,N_10179);
nor U12540 (N_12540,N_11990,N_11573);
nand U12541 (N_12541,N_10902,N_10103);
nand U12542 (N_12542,N_11454,N_11247);
nand U12543 (N_12543,N_10803,N_10301);
nand U12544 (N_12544,N_10269,N_11822);
nand U12545 (N_12545,N_10018,N_10240);
nand U12546 (N_12546,N_11630,N_10279);
or U12547 (N_12547,N_11466,N_11030);
nand U12548 (N_12548,N_11352,N_11360);
and U12549 (N_12549,N_11684,N_10398);
nand U12550 (N_12550,N_10130,N_10627);
nor U12551 (N_12551,N_11478,N_11411);
nand U12552 (N_12552,N_10209,N_10577);
and U12553 (N_12553,N_11231,N_11953);
and U12554 (N_12554,N_11336,N_11917);
or U12555 (N_12555,N_10805,N_10625);
and U12556 (N_12556,N_11617,N_10033);
or U12557 (N_12557,N_11889,N_10966);
or U12558 (N_12558,N_10581,N_10278);
and U12559 (N_12559,N_11671,N_10499);
and U12560 (N_12560,N_11528,N_11909);
nor U12561 (N_12561,N_10564,N_11563);
nand U12562 (N_12562,N_11931,N_11250);
xnor U12563 (N_12563,N_10919,N_11905);
nor U12564 (N_12564,N_11357,N_11116);
nor U12565 (N_12565,N_10544,N_11107);
nand U12566 (N_12566,N_10392,N_11108);
and U12567 (N_12567,N_11767,N_11748);
nand U12568 (N_12568,N_11239,N_11216);
and U12569 (N_12569,N_11426,N_10516);
or U12570 (N_12570,N_10227,N_11918);
or U12571 (N_12571,N_10058,N_10777);
or U12572 (N_12572,N_11601,N_11772);
nor U12573 (N_12573,N_10596,N_11502);
xor U12574 (N_12574,N_11700,N_10640);
nand U12575 (N_12575,N_10328,N_11655);
xor U12576 (N_12576,N_10381,N_10927);
nor U12577 (N_12577,N_10954,N_10624);
and U12578 (N_12578,N_11292,N_10853);
nand U12579 (N_12579,N_10037,N_10429);
nand U12580 (N_12580,N_11085,N_10529);
nor U12581 (N_12581,N_10003,N_10265);
nor U12582 (N_12582,N_10044,N_10910);
xor U12583 (N_12583,N_10705,N_11469);
or U12584 (N_12584,N_10572,N_11272);
and U12585 (N_12585,N_10666,N_10504);
or U12586 (N_12586,N_10557,N_11979);
nor U12587 (N_12587,N_10172,N_10875);
nand U12588 (N_12588,N_11865,N_11258);
and U12589 (N_12589,N_11260,N_11072);
and U12590 (N_12590,N_10298,N_10283);
nor U12591 (N_12591,N_11742,N_10694);
nand U12592 (N_12592,N_10988,N_10023);
nor U12593 (N_12593,N_10568,N_11128);
and U12594 (N_12594,N_10109,N_10879);
nand U12595 (N_12595,N_10690,N_10800);
xnor U12596 (N_12596,N_10567,N_11119);
and U12597 (N_12597,N_11036,N_11378);
or U12598 (N_12598,N_11982,N_10810);
or U12599 (N_12599,N_11530,N_11720);
nand U12600 (N_12600,N_11546,N_10097);
xor U12601 (N_12601,N_11668,N_11359);
nand U12602 (N_12602,N_11064,N_10335);
and U12603 (N_12603,N_10191,N_10133);
or U12604 (N_12604,N_10542,N_11787);
or U12605 (N_12605,N_11756,N_10631);
nand U12606 (N_12606,N_11259,N_11911);
nor U12607 (N_12607,N_10142,N_11134);
nand U12608 (N_12608,N_11235,N_10440);
nand U12609 (N_12609,N_11363,N_11835);
or U12610 (N_12610,N_10170,N_11964);
xnor U12611 (N_12611,N_10454,N_11706);
nand U12612 (N_12612,N_10726,N_11903);
nand U12613 (N_12613,N_10456,N_11003);
nand U12614 (N_12614,N_10929,N_10260);
nor U12615 (N_12615,N_10150,N_11900);
or U12616 (N_12616,N_10045,N_11268);
and U12617 (N_12617,N_11852,N_11833);
nor U12618 (N_12618,N_10418,N_10337);
or U12619 (N_12619,N_11473,N_10502);
nor U12620 (N_12620,N_11476,N_10629);
or U12621 (N_12621,N_11076,N_10146);
and U12622 (N_12622,N_11976,N_10969);
nand U12623 (N_12623,N_11220,N_11299);
or U12624 (N_12624,N_10786,N_10491);
or U12625 (N_12625,N_11839,N_11771);
or U12626 (N_12626,N_11809,N_10449);
xnor U12627 (N_12627,N_10177,N_10541);
nand U12628 (N_12628,N_11513,N_11140);
xor U12629 (N_12629,N_11661,N_11783);
or U12630 (N_12630,N_11698,N_10696);
nor U12631 (N_12631,N_11997,N_11752);
nand U12632 (N_12632,N_11844,N_11749);
and U12633 (N_12633,N_10121,N_10613);
xnor U12634 (N_12634,N_10555,N_10636);
or U12635 (N_12635,N_10432,N_11219);
nor U12636 (N_12636,N_11112,N_11155);
nor U12637 (N_12637,N_11413,N_11068);
nor U12638 (N_12638,N_11924,N_11798);
xnor U12639 (N_12639,N_10286,N_10937);
nor U12640 (N_12640,N_11500,N_11521);
and U12641 (N_12641,N_10933,N_10585);
xnor U12642 (N_12642,N_11332,N_11793);
xor U12643 (N_12643,N_10428,N_11651);
or U12644 (N_12644,N_10723,N_10375);
nor U12645 (N_12645,N_10474,N_11440);
nand U12646 (N_12646,N_11613,N_11090);
nor U12647 (N_12647,N_11084,N_10080);
xnor U12648 (N_12648,N_11198,N_10920);
xor U12649 (N_12649,N_10522,N_10884);
or U12650 (N_12650,N_10535,N_10229);
nand U12651 (N_12651,N_10042,N_10909);
and U12652 (N_12652,N_11840,N_10684);
or U12653 (N_12653,N_11404,N_10757);
and U12654 (N_12654,N_11079,N_10877);
and U12655 (N_12655,N_11503,N_11300);
nand U12656 (N_12656,N_11161,N_10698);
xor U12657 (N_12657,N_11118,N_10465);
and U12658 (N_12658,N_11152,N_10326);
xnor U12659 (N_12659,N_10531,N_10930);
or U12660 (N_12660,N_11410,N_10779);
nand U12661 (N_12661,N_10999,N_11385);
or U12662 (N_12662,N_10811,N_11894);
and U12663 (N_12663,N_10173,N_10709);
xnor U12664 (N_12664,N_11625,N_10776);
nand U12665 (N_12665,N_10487,N_10514);
nand U12666 (N_12666,N_11305,N_10846);
xor U12667 (N_12667,N_10199,N_10576);
and U12668 (N_12668,N_10840,N_11870);
nand U12669 (N_12669,N_10771,N_11184);
and U12670 (N_12670,N_11938,N_11193);
nand U12671 (N_12671,N_10031,N_10243);
or U12672 (N_12672,N_11061,N_11313);
xor U12673 (N_12673,N_11452,N_11038);
nand U12674 (N_12674,N_11328,N_10860);
nor U12675 (N_12675,N_11009,N_10558);
nor U12676 (N_12676,N_10385,N_10656);
or U12677 (N_12677,N_10296,N_10325);
nand U12678 (N_12678,N_10205,N_11421);
xnor U12679 (N_12679,N_11050,N_11590);
and U12680 (N_12680,N_11168,N_10476);
or U12681 (N_12681,N_10344,N_11602);
nor U12682 (N_12682,N_11289,N_11418);
nor U12683 (N_12683,N_11221,N_11174);
nand U12684 (N_12684,N_10620,N_11333);
or U12685 (N_12685,N_10458,N_11386);
nand U12686 (N_12686,N_10182,N_11144);
and U12687 (N_12687,N_10087,N_10353);
or U12688 (N_12688,N_11093,N_11031);
or U12689 (N_12689,N_10626,N_10387);
and U12690 (N_12690,N_10446,N_10994);
and U12691 (N_12691,N_11389,N_11560);
xor U12692 (N_12692,N_11475,N_11472);
xnor U12693 (N_12693,N_10424,N_11834);
and U12694 (N_12694,N_11283,N_10789);
and U12695 (N_12695,N_10804,N_10758);
xnor U12696 (N_12696,N_11179,N_10941);
xor U12697 (N_12697,N_11729,N_11823);
or U12698 (N_12698,N_10685,N_10747);
nand U12699 (N_12699,N_10579,N_10614);
or U12700 (N_12700,N_11871,N_11750);
xor U12701 (N_12701,N_11015,N_10026);
nor U12702 (N_12702,N_10663,N_10530);
or U12703 (N_12703,N_11382,N_11755);
xor U12704 (N_12704,N_10370,N_11148);
or U12705 (N_12705,N_10899,N_10857);
or U12706 (N_12706,N_10290,N_11255);
nor U12707 (N_12707,N_11724,N_11966);
or U12708 (N_12708,N_11083,N_11412);
nand U12709 (N_12709,N_10515,N_10025);
and U12710 (N_12710,N_10566,N_10332);
nor U12711 (N_12711,N_10383,N_11704);
and U12712 (N_12712,N_11722,N_11788);
nor U12713 (N_12713,N_11620,N_11129);
and U12714 (N_12714,N_10055,N_10774);
xnor U12715 (N_12715,N_11867,N_10125);
nor U12716 (N_12716,N_10397,N_10402);
xor U12717 (N_12717,N_10480,N_10892);
nor U12718 (N_12718,N_11510,N_10204);
nand U12719 (N_12719,N_11325,N_11948);
xnor U12720 (N_12720,N_11880,N_10396);
nand U12721 (N_12721,N_10604,N_10224);
nor U12722 (N_12722,N_11492,N_10472);
and U12723 (N_12723,N_10021,N_10677);
or U12724 (N_12724,N_10168,N_10464);
or U12725 (N_12725,N_10588,N_10653);
xnor U12726 (N_12726,N_11694,N_10912);
and U12727 (N_12727,N_11689,N_10300);
nor U12728 (N_12728,N_10665,N_11000);
nor U12729 (N_12729,N_11379,N_10198);
or U12730 (N_12730,N_11105,N_10630);
nor U12731 (N_12731,N_10318,N_10553);
and U12732 (N_12732,N_10949,N_10838);
or U12733 (N_12733,N_11315,N_11849);
nor U12734 (N_12734,N_10250,N_10048);
nand U12735 (N_12735,N_10896,N_10193);
nand U12736 (N_12736,N_10081,N_11136);
nand U12737 (N_12737,N_10145,N_11654);
xnor U12738 (N_12738,N_11117,N_11794);
xor U12739 (N_12739,N_11194,N_11624);
xnor U12740 (N_12740,N_11974,N_11372);
nand U12741 (N_12741,N_10996,N_10984);
and U12742 (N_12742,N_10431,N_10688);
or U12743 (N_12743,N_10634,N_10135);
nor U12744 (N_12744,N_11345,N_10559);
or U12745 (N_12745,N_11138,N_10101);
nand U12746 (N_12746,N_11464,N_10924);
nor U12747 (N_12747,N_10468,N_11669);
or U12748 (N_12748,N_10890,N_10140);
nor U12749 (N_12749,N_10865,N_11507);
nand U12750 (N_12750,N_11770,N_11837);
or U12751 (N_12751,N_10859,N_10019);
or U12752 (N_12752,N_10434,N_10056);
and U12753 (N_12753,N_11678,N_10189);
or U12754 (N_12754,N_10885,N_11578);
nor U12755 (N_12755,N_11842,N_10784);
and U12756 (N_12756,N_11430,N_10842);
and U12757 (N_12757,N_11131,N_11977);
and U12758 (N_12758,N_10316,N_10835);
nand U12759 (N_12759,N_10186,N_10485);
and U12760 (N_12760,N_11657,N_11644);
and U12761 (N_12761,N_10151,N_10471);
or U12762 (N_12762,N_11881,N_11482);
nor U12763 (N_12763,N_10536,N_11568);
xnor U12764 (N_12764,N_11329,N_11531);
nand U12765 (N_12765,N_11863,N_11646);
or U12766 (N_12766,N_11696,N_11645);
or U12767 (N_12767,N_11541,N_11037);
nand U12768 (N_12768,N_11312,N_10591);
nand U12769 (N_12769,N_10416,N_11306);
xor U12770 (N_12770,N_10288,N_10254);
xnor U12771 (N_12771,N_11400,N_10953);
xnor U12772 (N_12772,N_10482,N_11524);
or U12773 (N_12773,N_11162,N_11975);
and U12774 (N_12774,N_10897,N_10158);
nor U12775 (N_12775,N_10823,N_11402);
nand U12776 (N_12776,N_11065,N_11680);
and U12777 (N_12777,N_11929,N_10716);
or U12778 (N_12778,N_11542,N_10492);
nor U12779 (N_12779,N_11961,N_11821);
or U12780 (N_12780,N_10632,N_11113);
xnor U12781 (N_12781,N_10047,N_11725);
nand U12782 (N_12782,N_11157,N_11353);
xor U12783 (N_12783,N_11468,N_10837);
nand U12784 (N_12784,N_10114,N_11728);
xnor U12785 (N_12785,N_10998,N_11582);
and U12786 (N_12786,N_11480,N_10400);
or U12787 (N_12787,N_10791,N_11765);
and U12788 (N_12788,N_10086,N_11838);
and U12789 (N_12789,N_10212,N_11158);
nand U12790 (N_12790,N_11320,N_11670);
and U12791 (N_12791,N_11663,N_10527);
nand U12792 (N_12792,N_10785,N_10501);
xor U12793 (N_12793,N_11588,N_10643);
nand U12794 (N_12794,N_11719,N_10406);
xor U12795 (N_12795,N_10729,N_10024);
and U12796 (N_12796,N_11419,N_10752);
nor U12797 (N_12797,N_11101,N_11319);
and U12798 (N_12798,N_10762,N_10484);
nor U12799 (N_12799,N_10990,N_11791);
or U12800 (N_12800,N_10163,N_11626);
or U12801 (N_12801,N_11921,N_10560);
nand U12802 (N_12802,N_10965,N_10251);
xor U12803 (N_12803,N_11012,N_11991);
or U12804 (N_12804,N_10154,N_11972);
nor U12805 (N_12805,N_11666,N_10533);
xnor U12806 (N_12806,N_11963,N_10382);
xor U12807 (N_12807,N_10184,N_11304);
or U12808 (N_12808,N_11046,N_10302);
nor U12809 (N_12809,N_10852,N_11901);
xor U12810 (N_12810,N_10562,N_10112);
or U12811 (N_12811,N_10679,N_10678);
or U12812 (N_12812,N_11164,N_10782);
nor U12813 (N_12813,N_11828,N_10563);
or U12814 (N_12814,N_10799,N_10546);
xor U12815 (N_12815,N_11229,N_11137);
or U12816 (N_12816,N_10904,N_10517);
nand U12817 (N_12817,N_10369,N_11922);
xor U12818 (N_12818,N_10362,N_10356);
and U12819 (N_12819,N_11024,N_11762);
nor U12820 (N_12820,N_11420,N_10549);
nor U12821 (N_12821,N_10427,N_10703);
and U12822 (N_12822,N_10162,N_11394);
nor U12823 (N_12823,N_10952,N_11284);
xnor U12824 (N_12824,N_11857,N_11764);
and U12825 (N_12825,N_10831,N_10393);
or U12826 (N_12826,N_11878,N_11348);
and U12827 (N_12827,N_10490,N_10317);
nand U12828 (N_12828,N_11864,N_10778);
or U12829 (N_12829,N_11172,N_10007);
nor U12830 (N_12830,N_11600,N_10983);
nor U12831 (N_12831,N_10806,N_10979);
xor U12832 (N_12832,N_11189,N_11317);
or U12833 (N_12833,N_11790,N_11035);
xnor U12834 (N_12834,N_10167,N_10330);
xnor U12835 (N_12835,N_10946,N_10405);
nor U12836 (N_12836,N_11321,N_11998);
and U12837 (N_12837,N_11087,N_10371);
nor U12838 (N_12838,N_11397,N_10978);
and U12839 (N_12839,N_11686,N_11612);
or U12840 (N_12840,N_10523,N_11562);
nor U12841 (N_12841,N_10942,N_10637);
nor U12842 (N_12842,N_10099,N_11442);
nor U12843 (N_12843,N_10115,N_11846);
and U12844 (N_12844,N_11225,N_11032);
nand U12845 (N_12845,N_11641,N_10421);
or U12846 (N_12846,N_11370,N_11270);
xor U12847 (N_12847,N_10113,N_10215);
xnor U12848 (N_12848,N_11962,N_10306);
nand U12849 (N_12849,N_11572,N_10010);
xnor U12850 (N_12850,N_11377,N_11505);
and U12851 (N_12851,N_10068,N_11434);
or U12852 (N_12852,N_10320,N_10367);
or U12853 (N_12853,N_11274,N_10368);
and U12854 (N_12854,N_10528,N_11969);
xnor U12855 (N_12855,N_10856,N_10411);
nand U12856 (N_12856,N_10700,N_10069);
xor U12857 (N_12857,N_10138,N_11551);
nand U12858 (N_12858,N_10537,N_11417);
or U12859 (N_12859,N_10981,N_11872);
and U12860 (N_12860,N_11555,N_11579);
nor U12861 (N_12861,N_11014,N_11439);
nor U12862 (N_12862,N_10669,N_11349);
or U12863 (N_12863,N_11635,N_11406);
nor U12864 (N_12864,N_10822,N_11479);
or U12865 (N_12865,N_11873,N_11151);
nor U12866 (N_12866,N_10098,N_10259);
or U12867 (N_12867,N_10552,N_11013);
nor U12868 (N_12868,N_10120,N_11254);
nand U12869 (N_12869,N_10079,N_11175);
xor U12870 (N_12870,N_10453,N_10834);
or U12871 (N_12871,N_10412,N_10765);
xor U12872 (N_12872,N_11371,N_11745);
xor U12873 (N_12873,N_10334,N_10583);
xnor U12874 (N_12874,N_11490,N_10423);
nand U12875 (N_12875,N_10218,N_11109);
nor U12876 (N_12876,N_10408,N_11022);
or U12877 (N_12877,N_10511,N_10872);
nand U12878 (N_12878,N_11923,N_10587);
xnor U12879 (N_12879,N_11594,N_10264);
xnor U12880 (N_12880,N_10617,N_11688);
and U12881 (N_12881,N_10851,N_10104);
or U12882 (N_12882,N_10143,N_10355);
nor U12883 (N_12883,N_10280,N_10817);
and U12884 (N_12884,N_11092,N_11674);
or U12885 (N_12885,N_10923,N_11282);
xnor U12886 (N_12886,N_11532,N_11611);
and U12887 (N_12887,N_11687,N_11554);
or U12888 (N_12888,N_10404,N_10911);
nand U12889 (N_12889,N_10898,N_10181);
xor U12890 (N_12890,N_10832,N_11759);
and U12891 (N_12891,N_10312,N_10346);
and U12892 (N_12892,N_10858,N_11795);
or U12893 (N_12893,N_11522,N_11288);
or U12894 (N_12894,N_10281,N_10876);
nor U12895 (N_12895,N_10379,N_10628);
and U12896 (N_12896,N_11859,N_11387);
nand U12897 (N_12897,N_10027,N_10603);
xnor U12898 (N_12898,N_10123,N_10667);
nor U12899 (N_12899,N_11275,N_10268);
nand U12900 (N_12900,N_10733,N_11405);
nor U12901 (N_12901,N_10948,N_11935);
nand U12902 (N_12902,N_11801,N_10621);
and U12903 (N_12903,N_10745,N_11365);
nor U12904 (N_12904,N_11450,N_10090);
xor U12905 (N_12905,N_11391,N_11747);
xor U12906 (N_12906,N_11940,N_11294);
nor U12907 (N_12907,N_10311,N_10013);
nand U12908 (N_12908,N_11930,N_10724);
xnor U12909 (N_12909,N_10095,N_10615);
nand U12910 (N_12910,N_10461,N_10827);
nor U12911 (N_12911,N_10277,N_10538);
and U12912 (N_12912,N_11457,N_10693);
and U12913 (N_12913,N_11984,N_11081);
or U12914 (N_12914,N_10772,N_11519);
xnor U12915 (N_12915,N_11744,N_10323);
nor U12916 (N_12916,N_11561,N_11234);
nand U12917 (N_12917,N_10088,N_11673);
and U12918 (N_12918,N_11534,N_10276);
and U12919 (N_12919,N_10077,N_10657);
nand U12920 (N_12920,N_10153,N_10506);
or U12921 (N_12921,N_10864,N_10775);
nand U12922 (N_12922,N_10695,N_11029);
and U12923 (N_12923,N_10870,N_11679);
and U12924 (N_12924,N_11504,N_11721);
and U12925 (N_12925,N_10345,N_10116);
nand U12926 (N_12926,N_10790,N_10819);
nor U12927 (N_12927,N_10494,N_11509);
nor U12928 (N_12928,N_11256,N_11396);
xnor U12929 (N_12929,N_10395,N_10593);
nor U12930 (N_12930,N_11041,N_10545);
xor U12931 (N_12931,N_11238,N_11191);
nand U12932 (N_12932,N_10906,N_11805);
or U12933 (N_12933,N_10866,N_10728);
nand U12934 (N_12934,N_10419,N_10489);
nand U12935 (N_12935,N_10478,N_10417);
nor U12936 (N_12936,N_10128,N_10486);
and U12937 (N_12937,N_10893,N_11512);
and U12938 (N_12938,N_11647,N_10161);
xnor U12939 (N_12939,N_11785,N_10510);
or U12940 (N_12940,N_11691,N_11286);
nor U12941 (N_12941,N_10319,N_10327);
nand U12942 (N_12942,N_11916,N_10768);
nor U12943 (N_12943,N_11186,N_11253);
or U12944 (N_12944,N_10174,N_10053);
nand U12945 (N_12945,N_11890,N_11779);
and U12946 (N_12946,N_11942,N_10761);
nor U12947 (N_12947,N_10826,N_10147);
nor U12948 (N_12948,N_10144,N_10926);
nor U12949 (N_12949,N_10442,N_11978);
or U12950 (N_12950,N_11033,N_10655);
or U12951 (N_12951,N_11550,N_11422);
and U12952 (N_12952,N_10063,N_11407);
xor U12953 (N_12953,N_11060,N_10903);
or U12954 (N_12954,N_11799,N_11556);
or U12955 (N_12955,N_10833,N_10447);
or U12956 (N_12956,N_11800,N_10744);
nand U12957 (N_12957,N_11487,N_10848);
xnor U12958 (N_12958,N_11051,N_10329);
nand U12959 (N_12959,N_10867,N_10136);
or U12960 (N_12960,N_11496,N_11423);
nand U12961 (N_12961,N_11593,N_10372);
or U12962 (N_12962,N_10532,N_11495);
xnor U12963 (N_12963,N_10985,N_10697);
nand U12964 (N_12964,N_10376,N_11862);
and U12965 (N_12965,N_10253,N_10646);
or U12966 (N_12966,N_11078,N_10067);
and U12967 (N_12967,N_11067,N_11217);
nor U12968 (N_12968,N_11662,N_10391);
and U12969 (N_12969,N_11660,N_11681);
or U12970 (N_12970,N_10500,N_11103);
nand U12971 (N_12971,N_10691,N_11892);
nor U12972 (N_12972,N_10888,N_10769);
xor U12973 (N_12973,N_10014,N_10235);
xor U12974 (N_12974,N_10609,N_10654);
nand U12975 (N_12975,N_10363,N_10219);
nor U12976 (N_12976,N_11330,N_10249);
xor U12977 (N_12977,N_11543,N_11324);
and U12978 (N_12978,N_11196,N_11139);
nand U12979 (N_12979,N_11685,N_11557);
nand U12980 (N_12980,N_11453,N_10059);
or U12981 (N_12981,N_11830,N_10273);
nor U12982 (N_12982,N_10358,N_11879);
nand U12983 (N_12983,N_11047,N_10455);
xnor U12984 (N_12984,N_11769,N_11062);
nor U12985 (N_12985,N_11459,N_10939);
nor U12986 (N_12986,N_10307,N_10057);
or U12987 (N_12987,N_10683,N_10718);
xor U12988 (N_12988,N_10012,N_11633);
nand U12989 (N_12989,N_10959,N_11981);
nand U12990 (N_12990,N_10843,N_11934);
xnor U12991 (N_12991,N_11115,N_10119);
nor U12992 (N_12992,N_10004,N_11677);
nor U12993 (N_12993,N_11615,N_10169);
and U12994 (N_12994,N_10347,N_10554);
nand U12995 (N_12995,N_11746,N_11774);
xnor U12996 (N_12996,N_11874,N_11011);
or U12997 (N_12997,N_11574,N_10322);
and U12998 (N_12998,N_11877,N_10441);
or U12999 (N_12999,N_10950,N_10763);
nor U13000 (N_13000,N_11660,N_11328);
or U13001 (N_13001,N_10252,N_11352);
xor U13002 (N_13002,N_10800,N_10598);
nor U13003 (N_13003,N_10670,N_10495);
xor U13004 (N_13004,N_11953,N_11275);
xnor U13005 (N_13005,N_11825,N_11119);
xor U13006 (N_13006,N_10534,N_11655);
and U13007 (N_13007,N_10201,N_11239);
and U13008 (N_13008,N_10819,N_11329);
or U13009 (N_13009,N_11293,N_11473);
nor U13010 (N_13010,N_10479,N_11540);
xnor U13011 (N_13011,N_11660,N_11004);
nor U13012 (N_13012,N_10048,N_10751);
and U13013 (N_13013,N_10272,N_10150);
nor U13014 (N_13014,N_10410,N_10689);
nand U13015 (N_13015,N_11320,N_11548);
or U13016 (N_13016,N_10709,N_10058);
nand U13017 (N_13017,N_11397,N_11447);
or U13018 (N_13018,N_10079,N_11766);
and U13019 (N_13019,N_10999,N_11755);
or U13020 (N_13020,N_10443,N_11819);
or U13021 (N_13021,N_10238,N_10247);
xor U13022 (N_13022,N_10111,N_11910);
nor U13023 (N_13023,N_10591,N_10508);
nor U13024 (N_13024,N_11221,N_10371);
nand U13025 (N_13025,N_10946,N_11348);
or U13026 (N_13026,N_10334,N_11454);
xor U13027 (N_13027,N_10023,N_11256);
xnor U13028 (N_13028,N_10772,N_10099);
nor U13029 (N_13029,N_10209,N_11761);
xor U13030 (N_13030,N_11340,N_10831);
xnor U13031 (N_13031,N_10078,N_10562);
and U13032 (N_13032,N_10023,N_11991);
nor U13033 (N_13033,N_10261,N_10232);
and U13034 (N_13034,N_11997,N_10541);
and U13035 (N_13035,N_10162,N_10303);
xor U13036 (N_13036,N_11958,N_10062);
and U13037 (N_13037,N_10473,N_11755);
or U13038 (N_13038,N_10402,N_10772);
nor U13039 (N_13039,N_10103,N_11415);
nor U13040 (N_13040,N_11896,N_11447);
nand U13041 (N_13041,N_11247,N_11294);
nand U13042 (N_13042,N_10813,N_10877);
or U13043 (N_13043,N_11551,N_11719);
or U13044 (N_13044,N_10364,N_10857);
and U13045 (N_13045,N_10628,N_10873);
or U13046 (N_13046,N_11143,N_11303);
nand U13047 (N_13047,N_11880,N_11727);
and U13048 (N_13048,N_10502,N_11938);
nand U13049 (N_13049,N_11397,N_11355);
and U13050 (N_13050,N_10591,N_11941);
or U13051 (N_13051,N_10031,N_10801);
or U13052 (N_13052,N_11133,N_11330);
nor U13053 (N_13053,N_10051,N_11661);
nand U13054 (N_13054,N_10672,N_11380);
xnor U13055 (N_13055,N_11380,N_10700);
nor U13056 (N_13056,N_10876,N_11602);
nor U13057 (N_13057,N_11933,N_11986);
nor U13058 (N_13058,N_11799,N_10924);
or U13059 (N_13059,N_10914,N_10310);
and U13060 (N_13060,N_10015,N_11725);
nor U13061 (N_13061,N_11570,N_11753);
xor U13062 (N_13062,N_11746,N_11373);
or U13063 (N_13063,N_10381,N_10101);
xor U13064 (N_13064,N_11973,N_10228);
nor U13065 (N_13065,N_10710,N_11221);
nand U13066 (N_13066,N_11952,N_11792);
and U13067 (N_13067,N_10113,N_11879);
and U13068 (N_13068,N_10060,N_11107);
nor U13069 (N_13069,N_11155,N_11608);
nor U13070 (N_13070,N_10364,N_10765);
nand U13071 (N_13071,N_10334,N_11467);
nor U13072 (N_13072,N_10461,N_11679);
and U13073 (N_13073,N_11498,N_10652);
nor U13074 (N_13074,N_11892,N_10009);
or U13075 (N_13075,N_11881,N_10158);
and U13076 (N_13076,N_10953,N_11340);
and U13077 (N_13077,N_11386,N_10328);
nand U13078 (N_13078,N_10594,N_11247);
and U13079 (N_13079,N_11507,N_10497);
xnor U13080 (N_13080,N_11142,N_11724);
nor U13081 (N_13081,N_11854,N_11017);
and U13082 (N_13082,N_11294,N_10024);
nor U13083 (N_13083,N_11574,N_10920);
or U13084 (N_13084,N_10701,N_10554);
xor U13085 (N_13085,N_11839,N_10073);
and U13086 (N_13086,N_10816,N_11127);
xor U13087 (N_13087,N_10629,N_10035);
xnor U13088 (N_13088,N_11020,N_10303);
and U13089 (N_13089,N_11778,N_10792);
or U13090 (N_13090,N_10094,N_11077);
nand U13091 (N_13091,N_11796,N_11657);
or U13092 (N_13092,N_11517,N_11380);
nor U13093 (N_13093,N_11912,N_10259);
nor U13094 (N_13094,N_10884,N_10477);
or U13095 (N_13095,N_11177,N_11818);
nor U13096 (N_13096,N_10611,N_11002);
or U13097 (N_13097,N_10829,N_10216);
xnor U13098 (N_13098,N_11870,N_10804);
and U13099 (N_13099,N_10586,N_10583);
nand U13100 (N_13100,N_11663,N_10580);
nor U13101 (N_13101,N_10974,N_10577);
nand U13102 (N_13102,N_11516,N_11230);
nor U13103 (N_13103,N_11133,N_11885);
nand U13104 (N_13104,N_11936,N_11939);
xor U13105 (N_13105,N_11463,N_11282);
or U13106 (N_13106,N_11999,N_10533);
xor U13107 (N_13107,N_11970,N_10750);
and U13108 (N_13108,N_11389,N_11310);
nand U13109 (N_13109,N_11388,N_11530);
nor U13110 (N_13110,N_11195,N_11002);
xor U13111 (N_13111,N_11115,N_11524);
or U13112 (N_13112,N_11323,N_10548);
or U13113 (N_13113,N_10194,N_11744);
nor U13114 (N_13114,N_10608,N_10744);
xor U13115 (N_13115,N_11966,N_10297);
nand U13116 (N_13116,N_10582,N_10786);
nand U13117 (N_13117,N_11365,N_10361);
xor U13118 (N_13118,N_10842,N_10183);
nor U13119 (N_13119,N_11374,N_10794);
nand U13120 (N_13120,N_10403,N_11325);
or U13121 (N_13121,N_10646,N_11251);
or U13122 (N_13122,N_10381,N_11142);
nand U13123 (N_13123,N_10826,N_10422);
or U13124 (N_13124,N_11252,N_11476);
nor U13125 (N_13125,N_11787,N_10091);
nand U13126 (N_13126,N_10882,N_11999);
xnor U13127 (N_13127,N_10411,N_10521);
or U13128 (N_13128,N_11108,N_11382);
xnor U13129 (N_13129,N_10452,N_10295);
nand U13130 (N_13130,N_10201,N_10430);
nor U13131 (N_13131,N_11892,N_11643);
or U13132 (N_13132,N_11562,N_11405);
nand U13133 (N_13133,N_10226,N_10267);
or U13134 (N_13134,N_10662,N_10078);
and U13135 (N_13135,N_11869,N_11587);
xnor U13136 (N_13136,N_11240,N_11744);
or U13137 (N_13137,N_10243,N_10355);
and U13138 (N_13138,N_11840,N_10486);
or U13139 (N_13139,N_11810,N_11797);
xnor U13140 (N_13140,N_11944,N_11257);
xnor U13141 (N_13141,N_10611,N_10928);
and U13142 (N_13142,N_10937,N_10139);
and U13143 (N_13143,N_11699,N_11082);
nand U13144 (N_13144,N_11334,N_10628);
xnor U13145 (N_13145,N_10271,N_11825);
nor U13146 (N_13146,N_10472,N_11720);
or U13147 (N_13147,N_11288,N_11421);
or U13148 (N_13148,N_11820,N_11606);
nand U13149 (N_13149,N_10535,N_11109);
and U13150 (N_13150,N_11187,N_10423);
nor U13151 (N_13151,N_11901,N_10454);
xor U13152 (N_13152,N_10324,N_11044);
or U13153 (N_13153,N_11731,N_11837);
nor U13154 (N_13154,N_10548,N_10260);
or U13155 (N_13155,N_11790,N_10647);
nor U13156 (N_13156,N_11630,N_10450);
nand U13157 (N_13157,N_10667,N_11021);
nor U13158 (N_13158,N_10587,N_11823);
and U13159 (N_13159,N_10823,N_10035);
or U13160 (N_13160,N_10240,N_10110);
nor U13161 (N_13161,N_11271,N_10733);
and U13162 (N_13162,N_11031,N_10457);
xor U13163 (N_13163,N_11008,N_11103);
xnor U13164 (N_13164,N_10217,N_10103);
and U13165 (N_13165,N_10355,N_11575);
nor U13166 (N_13166,N_11799,N_11421);
and U13167 (N_13167,N_11622,N_10032);
or U13168 (N_13168,N_10705,N_10839);
nand U13169 (N_13169,N_11317,N_10458);
nor U13170 (N_13170,N_10881,N_11010);
nand U13171 (N_13171,N_11340,N_10822);
and U13172 (N_13172,N_10875,N_11493);
and U13173 (N_13173,N_10587,N_11933);
xor U13174 (N_13174,N_11720,N_10521);
and U13175 (N_13175,N_11185,N_11078);
or U13176 (N_13176,N_10500,N_11762);
nor U13177 (N_13177,N_11025,N_10099);
or U13178 (N_13178,N_10034,N_11750);
and U13179 (N_13179,N_11427,N_10920);
and U13180 (N_13180,N_10035,N_10086);
nand U13181 (N_13181,N_11520,N_10609);
nand U13182 (N_13182,N_10562,N_11439);
xor U13183 (N_13183,N_11847,N_11777);
nor U13184 (N_13184,N_11082,N_11544);
and U13185 (N_13185,N_10435,N_11362);
nand U13186 (N_13186,N_10365,N_11821);
xnor U13187 (N_13187,N_11741,N_11067);
xnor U13188 (N_13188,N_11596,N_10797);
nand U13189 (N_13189,N_11400,N_11386);
or U13190 (N_13190,N_10143,N_10670);
and U13191 (N_13191,N_10844,N_11868);
or U13192 (N_13192,N_10848,N_11875);
or U13193 (N_13193,N_10482,N_11449);
or U13194 (N_13194,N_10310,N_10281);
xor U13195 (N_13195,N_11291,N_11720);
nand U13196 (N_13196,N_11221,N_11242);
and U13197 (N_13197,N_11273,N_10768);
or U13198 (N_13198,N_11063,N_10367);
nor U13199 (N_13199,N_10836,N_10187);
nor U13200 (N_13200,N_10708,N_11860);
or U13201 (N_13201,N_11689,N_10412);
and U13202 (N_13202,N_10517,N_11780);
nand U13203 (N_13203,N_11554,N_10776);
and U13204 (N_13204,N_10608,N_10189);
and U13205 (N_13205,N_11831,N_11718);
xor U13206 (N_13206,N_10365,N_10072);
nand U13207 (N_13207,N_10049,N_10773);
nor U13208 (N_13208,N_10652,N_10752);
or U13209 (N_13209,N_11771,N_10939);
or U13210 (N_13210,N_10710,N_11249);
xor U13211 (N_13211,N_11516,N_10158);
xor U13212 (N_13212,N_11912,N_10942);
and U13213 (N_13213,N_11681,N_11609);
xnor U13214 (N_13214,N_11375,N_10268);
xor U13215 (N_13215,N_11559,N_11371);
and U13216 (N_13216,N_11775,N_11042);
or U13217 (N_13217,N_10617,N_10211);
or U13218 (N_13218,N_11970,N_10019);
and U13219 (N_13219,N_10978,N_10326);
nand U13220 (N_13220,N_10589,N_11410);
and U13221 (N_13221,N_11702,N_11824);
nor U13222 (N_13222,N_10599,N_11567);
xnor U13223 (N_13223,N_10711,N_11072);
nor U13224 (N_13224,N_10269,N_10313);
nor U13225 (N_13225,N_11503,N_11273);
and U13226 (N_13226,N_10195,N_11241);
nor U13227 (N_13227,N_10154,N_10854);
and U13228 (N_13228,N_10255,N_10677);
and U13229 (N_13229,N_10211,N_11392);
nand U13230 (N_13230,N_10956,N_11752);
xnor U13231 (N_13231,N_10539,N_10448);
xor U13232 (N_13232,N_10496,N_10487);
xnor U13233 (N_13233,N_11030,N_10881);
or U13234 (N_13234,N_10100,N_11168);
xnor U13235 (N_13235,N_11152,N_10772);
nor U13236 (N_13236,N_11888,N_11949);
xor U13237 (N_13237,N_10319,N_10259);
nand U13238 (N_13238,N_10902,N_11598);
xnor U13239 (N_13239,N_11974,N_11279);
or U13240 (N_13240,N_10563,N_10133);
nor U13241 (N_13241,N_10651,N_11872);
xor U13242 (N_13242,N_11122,N_10437);
or U13243 (N_13243,N_11731,N_11496);
nand U13244 (N_13244,N_11939,N_11879);
nor U13245 (N_13245,N_11815,N_10132);
xor U13246 (N_13246,N_11663,N_10960);
xor U13247 (N_13247,N_10642,N_10866);
and U13248 (N_13248,N_11667,N_10396);
nor U13249 (N_13249,N_11721,N_11164);
nand U13250 (N_13250,N_10940,N_11175);
and U13251 (N_13251,N_11950,N_11198);
nor U13252 (N_13252,N_10141,N_11955);
or U13253 (N_13253,N_10671,N_11246);
nand U13254 (N_13254,N_10763,N_10819);
xnor U13255 (N_13255,N_10706,N_11589);
and U13256 (N_13256,N_10618,N_11914);
nand U13257 (N_13257,N_10688,N_10928);
nand U13258 (N_13258,N_11254,N_10522);
nor U13259 (N_13259,N_11168,N_10025);
nand U13260 (N_13260,N_10315,N_10946);
and U13261 (N_13261,N_10103,N_10433);
nand U13262 (N_13262,N_10574,N_11817);
xnor U13263 (N_13263,N_11477,N_10728);
nor U13264 (N_13264,N_10230,N_11237);
nand U13265 (N_13265,N_10302,N_10562);
xor U13266 (N_13266,N_10232,N_11155);
and U13267 (N_13267,N_10269,N_10308);
or U13268 (N_13268,N_10944,N_10695);
xor U13269 (N_13269,N_11902,N_11486);
or U13270 (N_13270,N_11361,N_10072);
or U13271 (N_13271,N_11332,N_10029);
nor U13272 (N_13272,N_11047,N_11803);
nor U13273 (N_13273,N_10661,N_10890);
xor U13274 (N_13274,N_10037,N_11837);
or U13275 (N_13275,N_11302,N_10749);
or U13276 (N_13276,N_10277,N_10401);
xor U13277 (N_13277,N_10968,N_10035);
nand U13278 (N_13278,N_11690,N_10432);
nand U13279 (N_13279,N_10568,N_11248);
or U13280 (N_13280,N_11488,N_11217);
nand U13281 (N_13281,N_10639,N_11687);
xor U13282 (N_13282,N_10599,N_10684);
xnor U13283 (N_13283,N_11986,N_11369);
or U13284 (N_13284,N_11702,N_10833);
nor U13285 (N_13285,N_11586,N_10593);
or U13286 (N_13286,N_11762,N_10020);
nor U13287 (N_13287,N_11175,N_10267);
nor U13288 (N_13288,N_11944,N_10757);
xor U13289 (N_13289,N_11511,N_10468);
nand U13290 (N_13290,N_11447,N_11993);
nor U13291 (N_13291,N_11352,N_11340);
xnor U13292 (N_13292,N_10908,N_11591);
xnor U13293 (N_13293,N_10513,N_10912);
xnor U13294 (N_13294,N_11973,N_10568);
and U13295 (N_13295,N_10816,N_10335);
xnor U13296 (N_13296,N_10763,N_11872);
nor U13297 (N_13297,N_11091,N_10099);
nor U13298 (N_13298,N_11683,N_10045);
or U13299 (N_13299,N_11963,N_11877);
or U13300 (N_13300,N_11332,N_11071);
nor U13301 (N_13301,N_10696,N_11015);
nand U13302 (N_13302,N_10850,N_10517);
nor U13303 (N_13303,N_11669,N_11117);
or U13304 (N_13304,N_10639,N_10273);
nand U13305 (N_13305,N_11954,N_11236);
xnor U13306 (N_13306,N_11032,N_10043);
or U13307 (N_13307,N_10059,N_10096);
or U13308 (N_13308,N_11875,N_11215);
nand U13309 (N_13309,N_10298,N_10252);
nand U13310 (N_13310,N_10673,N_10819);
and U13311 (N_13311,N_11735,N_11281);
xnor U13312 (N_13312,N_10816,N_11356);
xor U13313 (N_13313,N_10411,N_10725);
nor U13314 (N_13314,N_10244,N_11623);
or U13315 (N_13315,N_10861,N_10557);
or U13316 (N_13316,N_10369,N_10484);
nand U13317 (N_13317,N_10304,N_11925);
xor U13318 (N_13318,N_11756,N_11369);
nand U13319 (N_13319,N_11039,N_11336);
or U13320 (N_13320,N_11037,N_10974);
or U13321 (N_13321,N_10181,N_10054);
and U13322 (N_13322,N_10486,N_10617);
and U13323 (N_13323,N_10075,N_10180);
nand U13324 (N_13324,N_11767,N_10404);
nand U13325 (N_13325,N_11009,N_10349);
nand U13326 (N_13326,N_10362,N_11279);
nand U13327 (N_13327,N_10082,N_10801);
or U13328 (N_13328,N_10802,N_11338);
nor U13329 (N_13329,N_11716,N_10758);
nand U13330 (N_13330,N_11965,N_10413);
and U13331 (N_13331,N_10094,N_11184);
xnor U13332 (N_13332,N_11845,N_11887);
nor U13333 (N_13333,N_11362,N_11377);
nand U13334 (N_13334,N_11212,N_11570);
nand U13335 (N_13335,N_10571,N_10163);
xor U13336 (N_13336,N_11490,N_10983);
xor U13337 (N_13337,N_10788,N_11401);
and U13338 (N_13338,N_11253,N_10526);
or U13339 (N_13339,N_10694,N_11179);
or U13340 (N_13340,N_10197,N_11090);
and U13341 (N_13341,N_10740,N_11077);
xor U13342 (N_13342,N_10162,N_11665);
nor U13343 (N_13343,N_10930,N_10662);
nor U13344 (N_13344,N_11284,N_11068);
nor U13345 (N_13345,N_11014,N_11812);
and U13346 (N_13346,N_11375,N_10615);
xor U13347 (N_13347,N_11333,N_11857);
nand U13348 (N_13348,N_10589,N_10870);
xor U13349 (N_13349,N_10599,N_10997);
xnor U13350 (N_13350,N_10060,N_11578);
or U13351 (N_13351,N_11419,N_11984);
xnor U13352 (N_13352,N_11415,N_11613);
nor U13353 (N_13353,N_11158,N_11285);
xor U13354 (N_13354,N_11517,N_10704);
nand U13355 (N_13355,N_11994,N_11656);
nor U13356 (N_13356,N_11427,N_10996);
and U13357 (N_13357,N_10823,N_10694);
nand U13358 (N_13358,N_10886,N_10014);
xnor U13359 (N_13359,N_10108,N_11865);
nand U13360 (N_13360,N_11157,N_10148);
or U13361 (N_13361,N_11295,N_10270);
nor U13362 (N_13362,N_10708,N_11956);
and U13363 (N_13363,N_10388,N_11829);
xor U13364 (N_13364,N_11692,N_10804);
nor U13365 (N_13365,N_11317,N_10708);
xor U13366 (N_13366,N_10405,N_11485);
xnor U13367 (N_13367,N_10393,N_10330);
xor U13368 (N_13368,N_10766,N_10298);
and U13369 (N_13369,N_11612,N_10167);
nand U13370 (N_13370,N_11061,N_10434);
xnor U13371 (N_13371,N_11297,N_11416);
nand U13372 (N_13372,N_10801,N_11827);
xor U13373 (N_13373,N_11231,N_11285);
or U13374 (N_13374,N_10555,N_11547);
or U13375 (N_13375,N_10388,N_10369);
and U13376 (N_13376,N_10352,N_11157);
nand U13377 (N_13377,N_10397,N_10513);
and U13378 (N_13378,N_11197,N_11346);
xor U13379 (N_13379,N_11189,N_10803);
nand U13380 (N_13380,N_11493,N_10410);
and U13381 (N_13381,N_11246,N_11633);
and U13382 (N_13382,N_10121,N_10592);
or U13383 (N_13383,N_11637,N_10836);
xnor U13384 (N_13384,N_11170,N_10013);
nand U13385 (N_13385,N_10353,N_10229);
or U13386 (N_13386,N_11185,N_11334);
and U13387 (N_13387,N_11488,N_11120);
nand U13388 (N_13388,N_11360,N_11251);
nor U13389 (N_13389,N_11039,N_10343);
nand U13390 (N_13390,N_11208,N_11962);
or U13391 (N_13391,N_10803,N_10779);
nand U13392 (N_13392,N_10384,N_10636);
nor U13393 (N_13393,N_10164,N_11107);
xnor U13394 (N_13394,N_10964,N_10144);
xnor U13395 (N_13395,N_11297,N_10731);
nand U13396 (N_13396,N_10100,N_11994);
or U13397 (N_13397,N_11200,N_10849);
or U13398 (N_13398,N_11209,N_10356);
nor U13399 (N_13399,N_11138,N_11542);
and U13400 (N_13400,N_11163,N_11653);
nor U13401 (N_13401,N_10605,N_10594);
xor U13402 (N_13402,N_11008,N_10349);
nand U13403 (N_13403,N_11696,N_11430);
or U13404 (N_13404,N_10509,N_10453);
and U13405 (N_13405,N_11181,N_11072);
or U13406 (N_13406,N_11730,N_11196);
and U13407 (N_13407,N_10334,N_11597);
and U13408 (N_13408,N_11259,N_10206);
or U13409 (N_13409,N_11235,N_10274);
and U13410 (N_13410,N_10413,N_10298);
xnor U13411 (N_13411,N_10057,N_10357);
nor U13412 (N_13412,N_10310,N_11500);
xor U13413 (N_13413,N_10033,N_11766);
xor U13414 (N_13414,N_10230,N_11564);
xnor U13415 (N_13415,N_10103,N_10266);
xnor U13416 (N_13416,N_11940,N_10147);
xnor U13417 (N_13417,N_11334,N_10023);
xnor U13418 (N_13418,N_10313,N_10806);
and U13419 (N_13419,N_11701,N_10755);
nand U13420 (N_13420,N_10336,N_10419);
nand U13421 (N_13421,N_10900,N_10974);
xor U13422 (N_13422,N_11336,N_11773);
xnor U13423 (N_13423,N_11556,N_10888);
nand U13424 (N_13424,N_10626,N_11286);
nor U13425 (N_13425,N_11049,N_10236);
xor U13426 (N_13426,N_11003,N_10062);
nor U13427 (N_13427,N_10667,N_11086);
nand U13428 (N_13428,N_11007,N_10699);
nand U13429 (N_13429,N_11162,N_11312);
and U13430 (N_13430,N_10790,N_10671);
nor U13431 (N_13431,N_10971,N_11919);
and U13432 (N_13432,N_10101,N_11651);
xor U13433 (N_13433,N_10114,N_11252);
xnor U13434 (N_13434,N_10994,N_10862);
nand U13435 (N_13435,N_10434,N_11903);
xnor U13436 (N_13436,N_11046,N_11476);
nand U13437 (N_13437,N_10714,N_11640);
nand U13438 (N_13438,N_10365,N_10684);
nand U13439 (N_13439,N_11846,N_11062);
nand U13440 (N_13440,N_11659,N_11068);
or U13441 (N_13441,N_11016,N_10182);
nand U13442 (N_13442,N_11373,N_10279);
and U13443 (N_13443,N_11387,N_11965);
xnor U13444 (N_13444,N_10136,N_11132);
and U13445 (N_13445,N_10017,N_11998);
nand U13446 (N_13446,N_11183,N_11629);
or U13447 (N_13447,N_11932,N_11250);
or U13448 (N_13448,N_10112,N_11487);
nand U13449 (N_13449,N_11463,N_11910);
nand U13450 (N_13450,N_10865,N_11053);
and U13451 (N_13451,N_10521,N_11598);
nor U13452 (N_13452,N_10122,N_10743);
nand U13453 (N_13453,N_11966,N_10301);
nor U13454 (N_13454,N_10394,N_11475);
xnor U13455 (N_13455,N_10314,N_11601);
xnor U13456 (N_13456,N_11386,N_10757);
or U13457 (N_13457,N_11985,N_10975);
nand U13458 (N_13458,N_10306,N_10421);
and U13459 (N_13459,N_11787,N_11050);
nor U13460 (N_13460,N_10012,N_11441);
nor U13461 (N_13461,N_10879,N_11845);
nor U13462 (N_13462,N_10509,N_10304);
nor U13463 (N_13463,N_11679,N_10201);
or U13464 (N_13464,N_11650,N_10955);
or U13465 (N_13465,N_10048,N_11292);
nor U13466 (N_13466,N_11289,N_10290);
nand U13467 (N_13467,N_11709,N_10966);
xnor U13468 (N_13468,N_10588,N_10331);
xnor U13469 (N_13469,N_10684,N_10296);
nor U13470 (N_13470,N_10510,N_10438);
or U13471 (N_13471,N_10006,N_11980);
xnor U13472 (N_13472,N_11070,N_10935);
and U13473 (N_13473,N_11253,N_11460);
nor U13474 (N_13474,N_11421,N_11080);
nor U13475 (N_13475,N_11916,N_11764);
or U13476 (N_13476,N_11934,N_10565);
and U13477 (N_13477,N_11963,N_10676);
xnor U13478 (N_13478,N_11057,N_10948);
and U13479 (N_13479,N_11727,N_11215);
or U13480 (N_13480,N_10449,N_11895);
and U13481 (N_13481,N_10592,N_11010);
and U13482 (N_13482,N_10977,N_10580);
nor U13483 (N_13483,N_10643,N_10937);
xor U13484 (N_13484,N_10658,N_11093);
nand U13485 (N_13485,N_10436,N_11726);
nand U13486 (N_13486,N_10819,N_11232);
xnor U13487 (N_13487,N_10103,N_11731);
or U13488 (N_13488,N_10867,N_11777);
nand U13489 (N_13489,N_10332,N_10842);
xnor U13490 (N_13490,N_10828,N_11286);
xor U13491 (N_13491,N_11760,N_11162);
or U13492 (N_13492,N_11879,N_11554);
nand U13493 (N_13493,N_10979,N_11532);
xnor U13494 (N_13494,N_11633,N_11992);
xnor U13495 (N_13495,N_11138,N_10758);
xor U13496 (N_13496,N_11144,N_10557);
or U13497 (N_13497,N_10197,N_10783);
xnor U13498 (N_13498,N_11349,N_11786);
or U13499 (N_13499,N_10647,N_11444);
nor U13500 (N_13500,N_11181,N_10496);
nor U13501 (N_13501,N_10489,N_11874);
nand U13502 (N_13502,N_10519,N_10987);
and U13503 (N_13503,N_11204,N_11065);
and U13504 (N_13504,N_10126,N_10333);
and U13505 (N_13505,N_11934,N_11680);
nor U13506 (N_13506,N_11503,N_10001);
and U13507 (N_13507,N_11465,N_11265);
and U13508 (N_13508,N_11274,N_10795);
and U13509 (N_13509,N_10367,N_11886);
nor U13510 (N_13510,N_10581,N_10008);
or U13511 (N_13511,N_10544,N_11544);
nor U13512 (N_13512,N_11813,N_11608);
xor U13513 (N_13513,N_10043,N_11841);
nor U13514 (N_13514,N_10916,N_11056);
xnor U13515 (N_13515,N_10626,N_11092);
and U13516 (N_13516,N_11324,N_10632);
nor U13517 (N_13517,N_10472,N_10640);
or U13518 (N_13518,N_11753,N_11448);
and U13519 (N_13519,N_11002,N_11775);
nand U13520 (N_13520,N_11548,N_10715);
xnor U13521 (N_13521,N_10397,N_11774);
or U13522 (N_13522,N_11633,N_10240);
nor U13523 (N_13523,N_11220,N_10196);
and U13524 (N_13524,N_10987,N_11617);
nand U13525 (N_13525,N_11010,N_10045);
xnor U13526 (N_13526,N_11073,N_10581);
and U13527 (N_13527,N_10524,N_10398);
xor U13528 (N_13528,N_11758,N_11157);
xor U13529 (N_13529,N_11195,N_10633);
xnor U13530 (N_13530,N_11238,N_10916);
nand U13531 (N_13531,N_11112,N_10051);
xor U13532 (N_13532,N_11468,N_11424);
nor U13533 (N_13533,N_10808,N_11661);
xor U13534 (N_13534,N_11611,N_10314);
or U13535 (N_13535,N_10467,N_10671);
nand U13536 (N_13536,N_11557,N_11978);
and U13537 (N_13537,N_10455,N_10414);
nand U13538 (N_13538,N_10745,N_11867);
nor U13539 (N_13539,N_10706,N_11523);
nor U13540 (N_13540,N_11806,N_11459);
and U13541 (N_13541,N_11679,N_11856);
and U13542 (N_13542,N_10752,N_10501);
xnor U13543 (N_13543,N_11749,N_11065);
or U13544 (N_13544,N_11050,N_10792);
or U13545 (N_13545,N_11113,N_10341);
nor U13546 (N_13546,N_10070,N_10351);
and U13547 (N_13547,N_10607,N_10735);
or U13548 (N_13548,N_10404,N_10951);
or U13549 (N_13549,N_11143,N_10125);
or U13550 (N_13550,N_11440,N_11457);
nor U13551 (N_13551,N_10979,N_10657);
or U13552 (N_13552,N_10423,N_11682);
or U13553 (N_13553,N_11739,N_10238);
xor U13554 (N_13554,N_11157,N_10471);
nand U13555 (N_13555,N_11717,N_11113);
or U13556 (N_13556,N_11390,N_10989);
nor U13557 (N_13557,N_11742,N_11168);
xor U13558 (N_13558,N_11401,N_11528);
or U13559 (N_13559,N_11438,N_10324);
and U13560 (N_13560,N_11724,N_11084);
and U13561 (N_13561,N_10116,N_10337);
nor U13562 (N_13562,N_10324,N_10393);
nand U13563 (N_13563,N_11804,N_10970);
nand U13564 (N_13564,N_11449,N_11981);
nand U13565 (N_13565,N_10052,N_10642);
and U13566 (N_13566,N_11010,N_10820);
or U13567 (N_13567,N_10541,N_11775);
and U13568 (N_13568,N_10966,N_11516);
nand U13569 (N_13569,N_11989,N_11314);
nand U13570 (N_13570,N_11298,N_10996);
xnor U13571 (N_13571,N_10722,N_11319);
and U13572 (N_13572,N_11135,N_11382);
xnor U13573 (N_13573,N_10081,N_11351);
or U13574 (N_13574,N_10550,N_10460);
xnor U13575 (N_13575,N_11371,N_11076);
and U13576 (N_13576,N_10519,N_11986);
nand U13577 (N_13577,N_11482,N_10345);
nor U13578 (N_13578,N_10557,N_11653);
or U13579 (N_13579,N_11656,N_11451);
or U13580 (N_13580,N_11145,N_10456);
nand U13581 (N_13581,N_10934,N_11412);
nand U13582 (N_13582,N_11469,N_11880);
nor U13583 (N_13583,N_10621,N_10873);
nand U13584 (N_13584,N_10503,N_10898);
nand U13585 (N_13585,N_11256,N_11413);
xor U13586 (N_13586,N_11057,N_11652);
and U13587 (N_13587,N_10063,N_11293);
nor U13588 (N_13588,N_10316,N_11137);
nand U13589 (N_13589,N_10850,N_10183);
and U13590 (N_13590,N_10189,N_10590);
nand U13591 (N_13591,N_11576,N_10353);
nand U13592 (N_13592,N_10583,N_11037);
nand U13593 (N_13593,N_11862,N_10047);
xnor U13594 (N_13594,N_11087,N_10259);
xnor U13595 (N_13595,N_11963,N_10608);
or U13596 (N_13596,N_11473,N_10520);
nor U13597 (N_13597,N_11340,N_10711);
xor U13598 (N_13598,N_11629,N_10902);
nor U13599 (N_13599,N_11401,N_10537);
and U13600 (N_13600,N_10949,N_11128);
and U13601 (N_13601,N_10417,N_11761);
and U13602 (N_13602,N_10885,N_10667);
xor U13603 (N_13603,N_11605,N_11036);
or U13604 (N_13604,N_10016,N_10256);
nor U13605 (N_13605,N_10033,N_10160);
nand U13606 (N_13606,N_10672,N_11765);
nand U13607 (N_13607,N_10746,N_10944);
or U13608 (N_13608,N_10558,N_11690);
and U13609 (N_13609,N_11248,N_10197);
and U13610 (N_13610,N_10893,N_11343);
or U13611 (N_13611,N_10407,N_11476);
nand U13612 (N_13612,N_10139,N_11713);
xor U13613 (N_13613,N_10101,N_10747);
or U13614 (N_13614,N_11203,N_10596);
or U13615 (N_13615,N_11798,N_11840);
nor U13616 (N_13616,N_10841,N_11502);
or U13617 (N_13617,N_10277,N_10795);
or U13618 (N_13618,N_10368,N_10887);
or U13619 (N_13619,N_11097,N_10840);
and U13620 (N_13620,N_10408,N_10465);
or U13621 (N_13621,N_11861,N_11094);
or U13622 (N_13622,N_10779,N_10730);
xor U13623 (N_13623,N_10488,N_10992);
nor U13624 (N_13624,N_10307,N_11299);
and U13625 (N_13625,N_11399,N_11673);
and U13626 (N_13626,N_11668,N_10109);
or U13627 (N_13627,N_11076,N_10177);
or U13628 (N_13628,N_11074,N_10635);
or U13629 (N_13629,N_10427,N_11784);
xnor U13630 (N_13630,N_10229,N_10114);
nand U13631 (N_13631,N_11099,N_11740);
nor U13632 (N_13632,N_10360,N_10523);
nand U13633 (N_13633,N_11434,N_11633);
xor U13634 (N_13634,N_11311,N_11107);
xnor U13635 (N_13635,N_11898,N_11372);
or U13636 (N_13636,N_11913,N_10886);
nand U13637 (N_13637,N_11964,N_10281);
or U13638 (N_13638,N_11245,N_10674);
and U13639 (N_13639,N_10334,N_11828);
nor U13640 (N_13640,N_11755,N_11975);
or U13641 (N_13641,N_10062,N_11036);
xor U13642 (N_13642,N_11329,N_10960);
xor U13643 (N_13643,N_11209,N_11637);
and U13644 (N_13644,N_10799,N_10234);
nor U13645 (N_13645,N_10449,N_10712);
and U13646 (N_13646,N_10453,N_10271);
or U13647 (N_13647,N_10603,N_11411);
nand U13648 (N_13648,N_10463,N_10367);
nor U13649 (N_13649,N_10270,N_10206);
and U13650 (N_13650,N_11580,N_10316);
xnor U13651 (N_13651,N_10824,N_11059);
or U13652 (N_13652,N_11529,N_10558);
and U13653 (N_13653,N_11626,N_10791);
or U13654 (N_13654,N_10869,N_11445);
nor U13655 (N_13655,N_10302,N_10037);
xnor U13656 (N_13656,N_10257,N_10603);
nor U13657 (N_13657,N_10805,N_10834);
or U13658 (N_13658,N_11196,N_11281);
nand U13659 (N_13659,N_11085,N_11672);
or U13660 (N_13660,N_11901,N_10513);
nand U13661 (N_13661,N_11701,N_11060);
nand U13662 (N_13662,N_11172,N_10189);
xnor U13663 (N_13663,N_10513,N_11563);
nand U13664 (N_13664,N_10802,N_10155);
or U13665 (N_13665,N_11515,N_10461);
nand U13666 (N_13666,N_10094,N_10990);
xor U13667 (N_13667,N_10548,N_10212);
nor U13668 (N_13668,N_10509,N_10584);
nor U13669 (N_13669,N_10621,N_10788);
xor U13670 (N_13670,N_11590,N_10064);
and U13671 (N_13671,N_10249,N_10529);
xor U13672 (N_13672,N_10508,N_11271);
or U13673 (N_13673,N_11000,N_10628);
nor U13674 (N_13674,N_11301,N_10578);
and U13675 (N_13675,N_10640,N_11580);
or U13676 (N_13676,N_11489,N_11425);
nand U13677 (N_13677,N_11678,N_10583);
and U13678 (N_13678,N_10773,N_10131);
xnor U13679 (N_13679,N_11270,N_10872);
or U13680 (N_13680,N_10314,N_11925);
nand U13681 (N_13681,N_10343,N_10625);
xnor U13682 (N_13682,N_11069,N_10558);
or U13683 (N_13683,N_11232,N_10781);
xnor U13684 (N_13684,N_11479,N_10450);
nand U13685 (N_13685,N_11228,N_10539);
and U13686 (N_13686,N_11948,N_10782);
nand U13687 (N_13687,N_11538,N_10132);
nand U13688 (N_13688,N_11264,N_11920);
or U13689 (N_13689,N_10506,N_10255);
nand U13690 (N_13690,N_11223,N_11013);
or U13691 (N_13691,N_11601,N_11989);
nor U13692 (N_13692,N_10025,N_10252);
and U13693 (N_13693,N_10766,N_11013);
and U13694 (N_13694,N_11741,N_11036);
nand U13695 (N_13695,N_10661,N_10517);
nand U13696 (N_13696,N_11233,N_10523);
and U13697 (N_13697,N_10455,N_10561);
nor U13698 (N_13698,N_10984,N_10200);
nor U13699 (N_13699,N_10462,N_10672);
xor U13700 (N_13700,N_11037,N_11743);
and U13701 (N_13701,N_10394,N_10525);
nand U13702 (N_13702,N_11825,N_10515);
xnor U13703 (N_13703,N_10760,N_10361);
nand U13704 (N_13704,N_10694,N_10452);
nor U13705 (N_13705,N_11419,N_11525);
nand U13706 (N_13706,N_11184,N_10122);
nor U13707 (N_13707,N_10604,N_10481);
and U13708 (N_13708,N_11515,N_10658);
nor U13709 (N_13709,N_11088,N_11866);
or U13710 (N_13710,N_10447,N_11177);
or U13711 (N_13711,N_10457,N_11718);
nor U13712 (N_13712,N_10638,N_10040);
nand U13713 (N_13713,N_10771,N_10063);
nand U13714 (N_13714,N_11220,N_11369);
xor U13715 (N_13715,N_10517,N_11374);
nand U13716 (N_13716,N_10524,N_10764);
nand U13717 (N_13717,N_11267,N_10633);
xor U13718 (N_13718,N_11995,N_11842);
or U13719 (N_13719,N_10500,N_10594);
nand U13720 (N_13720,N_11881,N_10858);
and U13721 (N_13721,N_10675,N_11792);
xor U13722 (N_13722,N_11741,N_11680);
nand U13723 (N_13723,N_11289,N_11910);
or U13724 (N_13724,N_11239,N_11884);
and U13725 (N_13725,N_10811,N_11321);
xnor U13726 (N_13726,N_10891,N_11217);
nor U13727 (N_13727,N_10179,N_10356);
nand U13728 (N_13728,N_11174,N_10928);
nor U13729 (N_13729,N_10213,N_11465);
or U13730 (N_13730,N_10208,N_11279);
xnor U13731 (N_13731,N_11054,N_11856);
and U13732 (N_13732,N_11521,N_10359);
xnor U13733 (N_13733,N_11456,N_11885);
and U13734 (N_13734,N_11907,N_11030);
or U13735 (N_13735,N_10014,N_11004);
nor U13736 (N_13736,N_10407,N_10147);
xor U13737 (N_13737,N_11173,N_11475);
nor U13738 (N_13738,N_11161,N_10902);
or U13739 (N_13739,N_10118,N_10134);
and U13740 (N_13740,N_11672,N_11025);
nor U13741 (N_13741,N_11282,N_10257);
or U13742 (N_13742,N_10244,N_10557);
and U13743 (N_13743,N_10191,N_11141);
or U13744 (N_13744,N_10354,N_10103);
nand U13745 (N_13745,N_11495,N_11953);
xor U13746 (N_13746,N_10570,N_11751);
nor U13747 (N_13747,N_11978,N_11603);
or U13748 (N_13748,N_10533,N_10466);
nor U13749 (N_13749,N_11831,N_10463);
and U13750 (N_13750,N_11307,N_11354);
and U13751 (N_13751,N_10013,N_10901);
xor U13752 (N_13752,N_11690,N_11539);
nand U13753 (N_13753,N_11283,N_10066);
xor U13754 (N_13754,N_11137,N_11126);
or U13755 (N_13755,N_10423,N_11719);
xor U13756 (N_13756,N_11658,N_10052);
xor U13757 (N_13757,N_10162,N_11485);
nand U13758 (N_13758,N_10313,N_11946);
and U13759 (N_13759,N_11383,N_10473);
nand U13760 (N_13760,N_11005,N_11116);
nand U13761 (N_13761,N_10428,N_10987);
nand U13762 (N_13762,N_11112,N_11399);
and U13763 (N_13763,N_11965,N_10404);
nor U13764 (N_13764,N_11760,N_10599);
xor U13765 (N_13765,N_10622,N_10446);
and U13766 (N_13766,N_10660,N_11214);
nand U13767 (N_13767,N_11260,N_10887);
or U13768 (N_13768,N_10877,N_10000);
and U13769 (N_13769,N_10886,N_11230);
nor U13770 (N_13770,N_11607,N_11256);
nor U13771 (N_13771,N_10095,N_11249);
xnor U13772 (N_13772,N_10381,N_10249);
nor U13773 (N_13773,N_11133,N_11683);
and U13774 (N_13774,N_11448,N_10226);
nor U13775 (N_13775,N_10300,N_10817);
nor U13776 (N_13776,N_10060,N_10434);
or U13777 (N_13777,N_11589,N_10357);
xnor U13778 (N_13778,N_10621,N_11746);
nand U13779 (N_13779,N_11535,N_11884);
nor U13780 (N_13780,N_10309,N_10691);
and U13781 (N_13781,N_11061,N_10322);
and U13782 (N_13782,N_10671,N_11544);
nor U13783 (N_13783,N_10270,N_11474);
or U13784 (N_13784,N_10998,N_11404);
and U13785 (N_13785,N_11557,N_10400);
nor U13786 (N_13786,N_11663,N_11254);
or U13787 (N_13787,N_10547,N_11882);
nand U13788 (N_13788,N_11957,N_10842);
or U13789 (N_13789,N_10805,N_11709);
or U13790 (N_13790,N_10587,N_10238);
nor U13791 (N_13791,N_10174,N_10825);
nand U13792 (N_13792,N_11611,N_10436);
and U13793 (N_13793,N_10620,N_10014);
nand U13794 (N_13794,N_11661,N_11027);
nor U13795 (N_13795,N_11033,N_11966);
xor U13796 (N_13796,N_10089,N_11703);
nor U13797 (N_13797,N_10377,N_10158);
xnor U13798 (N_13798,N_11905,N_11360);
xnor U13799 (N_13799,N_10554,N_10961);
nor U13800 (N_13800,N_10866,N_10732);
or U13801 (N_13801,N_11142,N_10245);
nand U13802 (N_13802,N_10983,N_10449);
nor U13803 (N_13803,N_10995,N_11939);
or U13804 (N_13804,N_10672,N_11353);
or U13805 (N_13805,N_11337,N_10638);
xor U13806 (N_13806,N_10000,N_10975);
and U13807 (N_13807,N_11286,N_10287);
xnor U13808 (N_13808,N_11332,N_11722);
and U13809 (N_13809,N_10742,N_10400);
and U13810 (N_13810,N_10902,N_10070);
nor U13811 (N_13811,N_10109,N_10852);
and U13812 (N_13812,N_10253,N_11895);
and U13813 (N_13813,N_10002,N_10792);
xor U13814 (N_13814,N_11673,N_11142);
xnor U13815 (N_13815,N_10028,N_11827);
xor U13816 (N_13816,N_11223,N_11682);
nand U13817 (N_13817,N_10514,N_10320);
xor U13818 (N_13818,N_10989,N_10018);
xnor U13819 (N_13819,N_11000,N_10265);
and U13820 (N_13820,N_11285,N_10957);
nand U13821 (N_13821,N_11027,N_11301);
or U13822 (N_13822,N_11535,N_10513);
nand U13823 (N_13823,N_11362,N_10919);
nand U13824 (N_13824,N_10107,N_10557);
nand U13825 (N_13825,N_10581,N_11803);
nand U13826 (N_13826,N_10153,N_10923);
nand U13827 (N_13827,N_10172,N_11991);
nand U13828 (N_13828,N_10108,N_10560);
xor U13829 (N_13829,N_11003,N_10000);
and U13830 (N_13830,N_10671,N_10695);
or U13831 (N_13831,N_11129,N_10071);
nor U13832 (N_13832,N_10136,N_11359);
nand U13833 (N_13833,N_10995,N_10259);
and U13834 (N_13834,N_11065,N_11176);
nor U13835 (N_13835,N_11524,N_11094);
or U13836 (N_13836,N_10998,N_11337);
nor U13837 (N_13837,N_11653,N_10090);
nor U13838 (N_13838,N_11731,N_11713);
nand U13839 (N_13839,N_11704,N_11030);
or U13840 (N_13840,N_11791,N_10054);
nor U13841 (N_13841,N_10817,N_10573);
or U13842 (N_13842,N_10818,N_11565);
nor U13843 (N_13843,N_10221,N_10428);
or U13844 (N_13844,N_10533,N_11942);
nand U13845 (N_13845,N_11080,N_11880);
nand U13846 (N_13846,N_10298,N_11124);
and U13847 (N_13847,N_11725,N_10625);
nand U13848 (N_13848,N_11041,N_10223);
nand U13849 (N_13849,N_11267,N_10271);
nand U13850 (N_13850,N_10687,N_11147);
xnor U13851 (N_13851,N_10368,N_10534);
or U13852 (N_13852,N_11025,N_11347);
or U13853 (N_13853,N_10515,N_10186);
nand U13854 (N_13854,N_11363,N_10464);
or U13855 (N_13855,N_11071,N_10043);
and U13856 (N_13856,N_11267,N_10169);
nand U13857 (N_13857,N_11060,N_11002);
and U13858 (N_13858,N_10633,N_11053);
xnor U13859 (N_13859,N_10830,N_11700);
and U13860 (N_13860,N_11321,N_11904);
nor U13861 (N_13861,N_10389,N_10186);
nand U13862 (N_13862,N_11348,N_11520);
nor U13863 (N_13863,N_10237,N_10202);
and U13864 (N_13864,N_10568,N_10587);
nand U13865 (N_13865,N_10402,N_11691);
xnor U13866 (N_13866,N_10799,N_11235);
and U13867 (N_13867,N_11274,N_11664);
and U13868 (N_13868,N_11383,N_10820);
and U13869 (N_13869,N_10384,N_11549);
nand U13870 (N_13870,N_11591,N_10690);
xnor U13871 (N_13871,N_11683,N_11626);
xor U13872 (N_13872,N_11107,N_11880);
nand U13873 (N_13873,N_11967,N_11352);
and U13874 (N_13874,N_11327,N_10326);
nor U13875 (N_13875,N_10751,N_11384);
nor U13876 (N_13876,N_10828,N_11495);
and U13877 (N_13877,N_10903,N_11544);
and U13878 (N_13878,N_10427,N_10913);
xor U13879 (N_13879,N_10462,N_11552);
and U13880 (N_13880,N_10585,N_10049);
and U13881 (N_13881,N_11042,N_11531);
and U13882 (N_13882,N_11686,N_11682);
and U13883 (N_13883,N_10443,N_10690);
xnor U13884 (N_13884,N_11769,N_10664);
nand U13885 (N_13885,N_10209,N_10070);
and U13886 (N_13886,N_10355,N_11626);
xnor U13887 (N_13887,N_11697,N_11228);
nor U13888 (N_13888,N_11518,N_10646);
or U13889 (N_13889,N_10188,N_10055);
and U13890 (N_13890,N_10062,N_11600);
or U13891 (N_13891,N_11021,N_11984);
or U13892 (N_13892,N_10392,N_10135);
and U13893 (N_13893,N_11702,N_11334);
xor U13894 (N_13894,N_10572,N_11846);
xnor U13895 (N_13895,N_11262,N_10215);
or U13896 (N_13896,N_10986,N_11419);
and U13897 (N_13897,N_10162,N_10449);
xnor U13898 (N_13898,N_10413,N_11293);
nor U13899 (N_13899,N_10227,N_11807);
nand U13900 (N_13900,N_10699,N_10120);
and U13901 (N_13901,N_11756,N_11430);
nand U13902 (N_13902,N_11024,N_11408);
nand U13903 (N_13903,N_10742,N_10846);
and U13904 (N_13904,N_10279,N_11254);
or U13905 (N_13905,N_11625,N_11781);
or U13906 (N_13906,N_11983,N_11259);
xnor U13907 (N_13907,N_10889,N_10574);
xor U13908 (N_13908,N_10514,N_11438);
xnor U13909 (N_13909,N_11027,N_10809);
xnor U13910 (N_13910,N_11159,N_10740);
and U13911 (N_13911,N_11281,N_11625);
or U13912 (N_13912,N_11472,N_10681);
and U13913 (N_13913,N_11959,N_10880);
and U13914 (N_13914,N_11958,N_11483);
xnor U13915 (N_13915,N_10937,N_11212);
xor U13916 (N_13916,N_11385,N_11253);
nand U13917 (N_13917,N_10119,N_10073);
xnor U13918 (N_13918,N_11989,N_11874);
xor U13919 (N_13919,N_10400,N_10851);
nor U13920 (N_13920,N_10015,N_11912);
and U13921 (N_13921,N_10639,N_10865);
and U13922 (N_13922,N_11400,N_11645);
nor U13923 (N_13923,N_10223,N_11452);
nor U13924 (N_13924,N_10810,N_10394);
nand U13925 (N_13925,N_11872,N_10538);
nand U13926 (N_13926,N_11570,N_11729);
nand U13927 (N_13927,N_11423,N_11272);
and U13928 (N_13928,N_11135,N_11096);
or U13929 (N_13929,N_10774,N_11679);
and U13930 (N_13930,N_10301,N_10922);
nand U13931 (N_13931,N_10910,N_11415);
and U13932 (N_13932,N_11181,N_10879);
or U13933 (N_13933,N_10588,N_10930);
xor U13934 (N_13934,N_10561,N_10921);
or U13935 (N_13935,N_10876,N_11545);
and U13936 (N_13936,N_11466,N_10554);
and U13937 (N_13937,N_10540,N_10876);
xor U13938 (N_13938,N_10324,N_11459);
nor U13939 (N_13939,N_10152,N_11245);
nor U13940 (N_13940,N_10622,N_11927);
and U13941 (N_13941,N_11073,N_11730);
xor U13942 (N_13942,N_10794,N_11316);
nand U13943 (N_13943,N_10603,N_10625);
xnor U13944 (N_13944,N_11455,N_11742);
xnor U13945 (N_13945,N_11872,N_11405);
or U13946 (N_13946,N_10614,N_11111);
or U13947 (N_13947,N_10696,N_10901);
and U13948 (N_13948,N_10168,N_11197);
and U13949 (N_13949,N_10662,N_10570);
nor U13950 (N_13950,N_11436,N_11811);
nor U13951 (N_13951,N_10619,N_10266);
xnor U13952 (N_13952,N_10026,N_11762);
or U13953 (N_13953,N_10801,N_11690);
nand U13954 (N_13954,N_11551,N_10710);
and U13955 (N_13955,N_10879,N_11116);
xnor U13956 (N_13956,N_10819,N_11008);
and U13957 (N_13957,N_10139,N_11404);
nor U13958 (N_13958,N_10178,N_10657);
or U13959 (N_13959,N_11526,N_11630);
and U13960 (N_13960,N_11336,N_10366);
nor U13961 (N_13961,N_10972,N_11957);
nand U13962 (N_13962,N_11345,N_10666);
or U13963 (N_13963,N_10048,N_11172);
and U13964 (N_13964,N_10201,N_11258);
and U13965 (N_13965,N_10608,N_11286);
or U13966 (N_13966,N_11039,N_11998);
and U13967 (N_13967,N_11796,N_11435);
or U13968 (N_13968,N_10222,N_11027);
and U13969 (N_13969,N_11669,N_11718);
nor U13970 (N_13970,N_11084,N_10265);
and U13971 (N_13971,N_10635,N_10682);
xnor U13972 (N_13972,N_10712,N_10388);
or U13973 (N_13973,N_11341,N_11810);
xor U13974 (N_13974,N_11413,N_11626);
nor U13975 (N_13975,N_11702,N_11919);
xor U13976 (N_13976,N_11653,N_10511);
nand U13977 (N_13977,N_10248,N_10497);
nand U13978 (N_13978,N_11008,N_10081);
nand U13979 (N_13979,N_10818,N_11159);
xnor U13980 (N_13980,N_11402,N_11725);
xor U13981 (N_13981,N_11245,N_10622);
or U13982 (N_13982,N_10272,N_10808);
nor U13983 (N_13983,N_10820,N_10274);
nand U13984 (N_13984,N_10282,N_10028);
nor U13985 (N_13985,N_10960,N_11135);
or U13986 (N_13986,N_10847,N_11530);
or U13987 (N_13987,N_11434,N_10183);
and U13988 (N_13988,N_11742,N_10510);
nor U13989 (N_13989,N_11870,N_11666);
or U13990 (N_13990,N_10074,N_11632);
xnor U13991 (N_13991,N_10287,N_10725);
and U13992 (N_13992,N_11808,N_11836);
and U13993 (N_13993,N_11735,N_10388);
nand U13994 (N_13994,N_11596,N_10217);
nor U13995 (N_13995,N_11774,N_10941);
nand U13996 (N_13996,N_11281,N_10068);
nor U13997 (N_13997,N_10349,N_10039);
nand U13998 (N_13998,N_10345,N_10537);
xor U13999 (N_13999,N_10554,N_11333);
xnor U14000 (N_14000,N_13914,N_12867);
and U14001 (N_14001,N_12648,N_12481);
or U14002 (N_14002,N_12830,N_13849);
nor U14003 (N_14003,N_12617,N_12152);
and U14004 (N_14004,N_12088,N_13236);
or U14005 (N_14005,N_13628,N_12026);
nor U14006 (N_14006,N_12076,N_12126);
or U14007 (N_14007,N_12091,N_13964);
nor U14008 (N_14008,N_13650,N_12354);
or U14009 (N_14009,N_13103,N_12628);
xnor U14010 (N_14010,N_12285,N_12164);
or U14011 (N_14011,N_12491,N_13657);
nor U14012 (N_14012,N_13741,N_12658);
and U14013 (N_14013,N_13416,N_13181);
nand U14014 (N_14014,N_12644,N_13438);
and U14015 (N_14015,N_13187,N_12567);
nand U14016 (N_14016,N_12016,N_13107);
and U14017 (N_14017,N_12103,N_13868);
nor U14018 (N_14018,N_12868,N_13592);
xor U14019 (N_14019,N_13493,N_12142);
nand U14020 (N_14020,N_12504,N_12849);
nand U14021 (N_14021,N_12257,N_13535);
nor U14022 (N_14022,N_12028,N_12559);
nand U14023 (N_14023,N_13118,N_12121);
and U14024 (N_14024,N_13803,N_12515);
nand U14025 (N_14025,N_13699,N_13003);
nor U14026 (N_14026,N_12966,N_13182);
xor U14027 (N_14027,N_13071,N_12826);
nand U14028 (N_14028,N_13109,N_12011);
nand U14029 (N_14029,N_13262,N_13464);
or U14030 (N_14030,N_12926,N_13128);
or U14031 (N_14031,N_12978,N_13058);
xnor U14032 (N_14032,N_13888,N_13225);
and U14033 (N_14033,N_13990,N_12937);
nor U14034 (N_14034,N_12700,N_12078);
xnor U14035 (N_14035,N_12056,N_13057);
nor U14036 (N_14036,N_13363,N_12842);
nand U14037 (N_14037,N_12097,N_13802);
nand U14038 (N_14038,N_13922,N_12009);
xnor U14039 (N_14039,N_12706,N_13101);
or U14040 (N_14040,N_13756,N_13596);
xor U14041 (N_14041,N_12450,N_13320);
nor U14042 (N_14042,N_12785,N_13916);
nand U14043 (N_14043,N_12642,N_13144);
and U14044 (N_14044,N_12203,N_12145);
nor U14045 (N_14045,N_13481,N_12513);
xor U14046 (N_14046,N_13085,N_12659);
nand U14047 (N_14047,N_12122,N_13510);
or U14048 (N_14048,N_13082,N_13078);
and U14049 (N_14049,N_13471,N_13897);
and U14050 (N_14050,N_12235,N_13745);
or U14051 (N_14051,N_12878,N_12095);
nand U14052 (N_14052,N_13069,N_12541);
nor U14053 (N_14053,N_12821,N_12034);
nor U14054 (N_14054,N_13525,N_13346);
and U14055 (N_14055,N_12753,N_12461);
xor U14056 (N_14056,N_12948,N_12347);
and U14057 (N_14057,N_12162,N_13534);
xor U14058 (N_14058,N_13726,N_12792);
and U14059 (N_14059,N_13976,N_13074);
or U14060 (N_14060,N_12917,N_12955);
nand U14061 (N_14061,N_13957,N_13517);
xor U14062 (N_14062,N_13893,N_13958);
and U14063 (N_14063,N_12805,N_13938);
nor U14064 (N_14064,N_13064,N_13806);
or U14065 (N_14065,N_12958,N_13828);
xnor U14066 (N_14066,N_13361,N_12265);
nor U14067 (N_14067,N_12176,N_13981);
and U14068 (N_14068,N_12580,N_13417);
xnor U14069 (N_14069,N_12277,N_12775);
nor U14070 (N_14070,N_13325,N_13436);
and U14071 (N_14071,N_13117,N_12987);
or U14072 (N_14072,N_12779,N_13560);
and U14073 (N_14073,N_13638,N_12673);
and U14074 (N_14074,N_12360,N_12272);
and U14075 (N_14075,N_13646,N_13848);
or U14076 (N_14076,N_12804,N_12199);
xor U14077 (N_14077,N_12799,N_12790);
or U14078 (N_14078,N_13676,N_12731);
xnor U14079 (N_14079,N_13904,N_13659);
xnor U14080 (N_14080,N_13331,N_12367);
or U14081 (N_14081,N_13029,N_12260);
nor U14082 (N_14082,N_12953,N_12287);
or U14083 (N_14083,N_13420,N_12940);
nand U14084 (N_14084,N_12189,N_12465);
or U14085 (N_14085,N_13739,N_13090);
and U14086 (N_14086,N_13165,N_13094);
nand U14087 (N_14087,N_12857,N_13096);
nor U14088 (N_14088,N_12601,N_12668);
or U14089 (N_14089,N_13915,N_13430);
or U14090 (N_14090,N_12426,N_12378);
or U14091 (N_14091,N_12242,N_12568);
nor U14092 (N_14092,N_13686,N_13546);
nand U14093 (N_14093,N_13454,N_12197);
or U14094 (N_14094,N_13286,N_13448);
nand U14095 (N_14095,N_13087,N_12661);
xor U14096 (N_14096,N_13786,N_12518);
nand U14097 (N_14097,N_13251,N_13402);
xor U14098 (N_14098,N_12240,N_12968);
and U14099 (N_14099,N_13813,N_12425);
and U14100 (N_14100,N_13776,N_12362);
or U14101 (N_14101,N_12839,N_12664);
nor U14102 (N_14102,N_13293,N_12050);
or U14103 (N_14103,N_13511,N_12971);
and U14104 (N_14104,N_13671,N_13642);
nor U14105 (N_14105,N_13937,N_12886);
nand U14106 (N_14106,N_13805,N_13954);
nor U14107 (N_14107,N_13788,N_12906);
nand U14108 (N_14108,N_12818,N_13495);
xnor U14109 (N_14109,N_12527,N_12024);
nor U14110 (N_14110,N_12557,N_12042);
or U14111 (N_14111,N_12333,N_13449);
xnor U14112 (N_14112,N_13912,N_13791);
xnor U14113 (N_14113,N_13451,N_12087);
xor U14114 (N_14114,N_12787,N_12548);
or U14115 (N_14115,N_13799,N_12092);
nor U14116 (N_14116,N_13220,N_12634);
nor U14117 (N_14117,N_12292,N_13947);
nand U14118 (N_14118,N_13162,N_13705);
or U14119 (N_14119,N_13193,N_13426);
or U14120 (N_14120,N_13617,N_13163);
or U14121 (N_14121,N_13291,N_12519);
or U14122 (N_14122,N_13539,N_12690);
xor U14123 (N_14123,N_12094,N_13861);
nand U14124 (N_14124,N_13266,N_13605);
and U14125 (N_14125,N_13401,N_12813);
and U14126 (N_14126,N_12411,N_12326);
xor U14127 (N_14127,N_13939,N_13250);
xor U14128 (N_14128,N_13318,N_13298);
xor U14129 (N_14129,N_13512,N_13649);
nor U14130 (N_14130,N_12707,N_13825);
xnor U14131 (N_14131,N_13407,N_13431);
and U14132 (N_14132,N_13886,N_13554);
nor U14133 (N_14133,N_13682,N_12616);
nor U14134 (N_14134,N_12119,N_12205);
nand U14135 (N_14135,N_12531,N_12536);
nor U14136 (N_14136,N_12043,N_13081);
xnor U14137 (N_14137,N_12381,N_13950);
and U14138 (N_14138,N_13382,N_12049);
nor U14139 (N_14139,N_12751,N_13767);
nor U14140 (N_14140,N_12832,N_12669);
xnor U14141 (N_14141,N_12068,N_12851);
and U14142 (N_14142,N_12607,N_13288);
nor U14143 (N_14143,N_13159,N_12363);
or U14144 (N_14144,N_13940,N_12371);
nor U14145 (N_14145,N_12517,N_13877);
nor U14146 (N_14146,N_13555,N_13782);
nand U14147 (N_14147,N_12848,N_13004);
or U14148 (N_14148,N_12942,N_13818);
and U14149 (N_14149,N_12105,N_12772);
or U14150 (N_14150,N_12035,N_12633);
nand U14151 (N_14151,N_13365,N_12179);
or U14152 (N_14152,N_12113,N_12332);
nand U14153 (N_14153,N_13487,N_12214);
nor U14154 (N_14154,N_12258,N_13235);
nand U14155 (N_14155,N_13344,N_13845);
or U14156 (N_14156,N_13866,N_12671);
and U14157 (N_14157,N_13993,N_12727);
xor U14158 (N_14158,N_13651,N_12720);
nand U14159 (N_14159,N_13390,N_13373);
nor U14160 (N_14160,N_13059,N_12928);
nor U14161 (N_14161,N_13906,N_12337);
or U14162 (N_14162,N_13932,N_12489);
nor U14163 (N_14163,N_12086,N_13450);
xnor U14164 (N_14164,N_12823,N_13027);
xor U14165 (N_14165,N_12865,N_13244);
nand U14166 (N_14166,N_12036,N_12138);
nand U14167 (N_14167,N_12484,N_13854);
nand U14168 (N_14168,N_13793,N_12710);
and U14169 (N_14169,N_13785,N_12981);
nor U14170 (N_14170,N_12793,N_12570);
xor U14171 (N_14171,N_13795,N_13614);
xnor U14172 (N_14172,N_12532,N_12336);
or U14173 (N_14173,N_13777,N_12526);
and U14174 (N_14174,N_13789,N_13328);
xnor U14175 (N_14175,N_12623,N_12665);
xnor U14176 (N_14176,N_13062,N_12918);
or U14177 (N_14177,N_12353,N_13393);
nand U14178 (N_14178,N_12863,N_12758);
nand U14179 (N_14179,N_12212,N_13704);
xor U14180 (N_14180,N_13290,N_12188);
or U14181 (N_14181,N_13160,N_12451);
or U14182 (N_14182,N_12789,N_12930);
nand U14183 (N_14183,N_12629,N_13584);
xor U14184 (N_14184,N_13025,N_12810);
nand U14185 (N_14185,N_12679,N_13405);
and U14186 (N_14186,N_12657,N_12296);
nor U14187 (N_14187,N_13282,N_13891);
or U14188 (N_14188,N_12429,N_13558);
xor U14189 (N_14189,N_13043,N_13122);
or U14190 (N_14190,N_13368,N_13017);
xor U14191 (N_14191,N_13229,N_12428);
xnor U14192 (N_14192,N_13590,N_12158);
nor U14193 (N_14193,N_13237,N_13701);
and U14194 (N_14194,N_13689,N_12038);
or U14195 (N_14195,N_12972,N_12402);
nand U14196 (N_14196,N_12936,N_12494);
nand U14197 (N_14197,N_13885,N_13427);
or U14198 (N_14198,N_13456,N_12973);
nor U14199 (N_14199,N_12870,N_12058);
xnor U14200 (N_14200,N_12074,N_13720);
and U14201 (N_14201,N_13624,N_12374);
nor U14202 (N_14202,N_13292,N_13052);
nand U14203 (N_14203,N_13284,N_12469);
nor U14204 (N_14204,N_12675,N_13223);
nand U14205 (N_14205,N_13227,N_12912);
xor U14206 (N_14206,N_12651,N_13551);
nand U14207 (N_14207,N_13507,N_13790);
and U14208 (N_14208,N_13724,N_12027);
nand U14209 (N_14209,N_12811,N_13158);
and U14210 (N_14210,N_12396,N_12072);
nor U14211 (N_14211,N_12008,N_12010);
nand U14212 (N_14212,N_13597,N_13717);
xnor U14213 (N_14213,N_13413,N_12649);
nand U14214 (N_14214,N_13092,N_12443);
nand U14215 (N_14215,N_13210,N_13145);
nand U14216 (N_14216,N_13760,N_12471);
and U14217 (N_14217,N_13870,N_13364);
xor U14218 (N_14218,N_12051,N_13688);
nand U14219 (N_14219,N_12488,N_12406);
and U14220 (N_14220,N_13046,N_13600);
or U14221 (N_14221,N_13484,N_13569);
and U14222 (N_14222,N_12713,N_12639);
and U14223 (N_14223,N_13977,N_12167);
and U14224 (N_14224,N_13809,N_13821);
nor U14225 (N_14225,N_13974,N_13421);
nor U14226 (N_14226,N_13312,N_12773);
nor U14227 (N_14227,N_13541,N_12029);
nand U14228 (N_14228,N_12756,N_13956);
and U14229 (N_14229,N_13224,N_12304);
nor U14230 (N_14230,N_12259,N_13833);
nand U14231 (N_14231,N_13611,N_12213);
nand U14232 (N_14232,N_13553,N_12183);
and U14233 (N_14233,N_13710,N_12542);
nand U14234 (N_14234,N_12275,N_13556);
or U14235 (N_14235,N_13826,N_12284);
and U14236 (N_14236,N_12646,N_13972);
nand U14237 (N_14237,N_13690,N_12874);
and U14238 (N_14238,N_13911,N_12514);
xnor U14239 (N_14239,N_12047,N_12195);
nor U14240 (N_14240,N_13437,N_13340);
xor U14241 (N_14241,N_12576,N_12127);
or U14242 (N_14242,N_12916,N_12654);
nand U14243 (N_14243,N_13441,N_13567);
nand U14244 (N_14244,N_13696,N_13549);
or U14245 (N_14245,N_13547,N_12533);
and U14246 (N_14246,N_13585,N_13028);
nor U14247 (N_14247,N_13858,N_12635);
nand U14248 (N_14248,N_13113,N_12650);
nor U14249 (N_14249,N_12237,N_12090);
or U14250 (N_14250,N_12390,N_13816);
xor U14251 (N_14251,N_13189,N_13254);
nand U14252 (N_14252,N_13422,N_13734);
and U14253 (N_14253,N_12717,N_12460);
or U14254 (N_14254,N_12175,N_12636);
nor U14255 (N_14255,N_13719,N_12967);
and U14256 (N_14256,N_13377,N_12512);
and U14257 (N_14257,N_12828,N_13475);
xor U14258 (N_14258,N_12156,N_13662);
and U14259 (N_14259,N_13761,N_13149);
xor U14260 (N_14260,N_12831,N_12077);
xnor U14261 (N_14261,N_12022,N_13385);
or U14262 (N_14262,N_13079,N_13751);
nand U14263 (N_14263,N_12031,N_13141);
xor U14264 (N_14264,N_13342,N_12932);
nand U14265 (N_14265,N_12132,N_12563);
or U14266 (N_14266,N_13499,N_12455);
and U14267 (N_14267,N_12941,N_13006);
xnor U14268 (N_14268,N_13823,N_13133);
nor U14269 (N_14269,N_12314,N_12505);
nor U14270 (N_14270,N_12934,N_12392);
nor U14271 (N_14271,N_13496,N_13781);
nor U14272 (N_14272,N_12282,N_13321);
or U14273 (N_14273,N_13907,N_12018);
nor U14274 (N_14274,N_12879,N_13249);
xnor U14275 (N_14275,N_13852,N_13860);
xnor U14276 (N_14276,N_13980,N_12280);
and U14277 (N_14277,N_12129,N_13458);
nand U14278 (N_14278,N_13768,N_12692);
xor U14279 (N_14279,N_12909,N_12246);
xnor U14280 (N_14280,N_13049,N_13900);
and U14281 (N_14281,N_13301,N_12432);
nand U14282 (N_14282,N_12317,N_12929);
or U14283 (N_14283,N_13953,N_13995);
and U14284 (N_14284,N_13665,N_13440);
nand U14285 (N_14285,N_12446,N_12062);
nand U14286 (N_14286,N_13272,N_13934);
and U14287 (N_14287,N_13930,N_12418);
nand U14288 (N_14288,N_12437,N_13263);
nor U14289 (N_14289,N_12738,N_13199);
or U14290 (N_14290,N_13376,N_13519);
xnor U14291 (N_14291,N_12680,N_12174);
xnor U14292 (N_14292,N_12391,N_13216);
nor U14293 (N_14293,N_13242,N_12053);
or U14294 (N_14294,N_12577,N_12331);
xnor U14295 (N_14295,N_12001,N_13654);
or U14296 (N_14296,N_12903,N_13260);
nor U14297 (N_14297,N_12814,N_13335);
or U14298 (N_14298,N_13479,N_13847);
nor U14299 (N_14299,N_12573,N_13645);
xnor U14300 (N_14300,N_12575,N_13022);
and U14301 (N_14301,N_13687,N_13388);
nand U14302 (N_14302,N_13743,N_12816);
or U14303 (N_14303,N_12670,N_12797);
nand U14304 (N_14304,N_12609,N_12595);
xor U14305 (N_14305,N_13629,N_13559);
nor U14306 (N_14306,N_12073,N_12989);
nor U14307 (N_14307,N_13247,N_12403);
xor U14308 (N_14308,N_12744,N_13276);
xor U14309 (N_14309,N_13123,N_13946);
nor U14310 (N_14310,N_13380,N_12747);
and U14311 (N_14311,N_12896,N_13865);
or U14312 (N_14312,N_12992,N_12422);
nor U14313 (N_14313,N_13086,N_12591);
and U14314 (N_14314,N_12862,N_12012);
or U14315 (N_14315,N_13238,N_12725);
nor U14316 (N_14316,N_13195,N_13391);
xor U14317 (N_14317,N_12254,N_12225);
nand U14318 (N_14318,N_12919,N_13142);
and U14319 (N_14319,N_12477,N_12439);
xnor U14320 (N_14320,N_13604,N_12069);
nand U14321 (N_14321,N_13644,N_12970);
nand U14322 (N_14322,N_12625,N_12410);
nand U14323 (N_14323,N_13051,N_13641);
nor U14324 (N_14324,N_13537,N_13168);
xor U14325 (N_14325,N_12487,N_12998);
nand U14326 (N_14326,N_12757,N_13680);
or U14327 (N_14327,N_13121,N_13208);
xnor U14328 (N_14328,N_12291,N_13194);
nand U14329 (N_14329,N_12441,N_13982);
nand U14330 (N_14330,N_13639,N_13444);
and U14331 (N_14331,N_12734,N_12444);
xnor U14332 (N_14332,N_12276,N_13709);
or U14333 (N_14333,N_13008,N_13672);
or U14334 (N_14334,N_12698,N_12436);
or U14335 (N_14335,N_13652,N_12769);
nand U14336 (N_14336,N_12215,N_13386);
or U14337 (N_14337,N_13742,N_13372);
or U14338 (N_14338,N_12351,N_12478);
nor U14339 (N_14339,N_13289,N_13703);
and U14340 (N_14340,N_13452,N_13829);
or U14341 (N_14341,N_13478,N_13418);
and U14342 (N_14342,N_13787,N_12844);
and U14343 (N_14343,N_12566,N_13613);
xor U14344 (N_14344,N_13524,N_13913);
xnor U14345 (N_14345,N_13898,N_12453);
and U14346 (N_14346,N_13582,N_13513);
nor U14347 (N_14347,N_12185,N_12977);
or U14348 (N_14348,N_12082,N_13076);
nor U14349 (N_14349,N_12303,N_12569);
and U14350 (N_14350,N_12388,N_12550);
or U14351 (N_14351,N_13920,N_12767);
nor U14352 (N_14352,N_13814,N_13986);
xnor U14353 (N_14353,N_12893,N_12462);
and U14354 (N_14354,N_12687,N_12549);
nor U14355 (N_14355,N_12956,N_13764);
and U14356 (N_14356,N_12547,N_12180);
nor U14357 (N_14357,N_13044,N_12125);
and U14358 (N_14358,N_13476,N_12344);
and U14359 (N_14359,N_12606,N_13443);
and U14360 (N_14360,N_13447,N_12829);
or U14361 (N_14361,N_13747,N_12096);
nand U14362 (N_14362,N_12057,N_13231);
or U14363 (N_14363,N_13300,N_13580);
or U14364 (N_14364,N_13504,N_12869);
and U14365 (N_14365,N_13902,N_12715);
nand U14366 (N_14366,N_13856,N_12579);
and U14367 (N_14367,N_13925,N_13397);
and U14368 (N_14368,N_12825,N_12102);
xnor U14369 (N_14369,N_13362,N_12562);
and U14370 (N_14370,N_12216,N_12807);
nor U14371 (N_14371,N_13975,N_13518);
nand U14372 (N_14372,N_12054,N_13152);
nor U14373 (N_14373,N_13942,N_13640);
nor U14374 (N_14374,N_12365,N_12316);
and U14375 (N_14375,N_13396,N_12033);
nor U14376 (N_14376,N_12501,N_12357);
and U14377 (N_14377,N_12473,N_12066);
or U14378 (N_14378,N_13945,N_13048);
nor U14379 (N_14379,N_13486,N_12366);
xnor U14380 (N_14380,N_13246,N_13267);
xnor U14381 (N_14381,N_13574,N_12055);
or U14382 (N_14382,N_13038,N_13089);
nor U14383 (N_14383,N_12630,N_13804);
nor U14384 (N_14384,N_13329,N_12140);
and U14385 (N_14385,N_12976,N_12427);
nor U14386 (N_14386,N_13749,N_13055);
nor U14387 (N_14387,N_12286,N_13603);
or U14388 (N_14388,N_13429,N_13354);
or U14389 (N_14389,N_12424,N_13024);
or U14390 (N_14390,N_13269,N_13068);
xor U14391 (N_14391,N_12841,N_13116);
nand U14392 (N_14392,N_12343,N_12529);
or U14393 (N_14393,N_12298,N_12760);
xnor U14394 (N_14394,N_13273,N_13483);
xnor U14395 (N_14395,N_13005,N_13515);
or U14396 (N_14396,N_13631,N_13998);
nand U14397 (N_14397,N_12433,N_13664);
or U14398 (N_14398,N_12382,N_13350);
or U14399 (N_14399,N_13498,N_13610);
and U14400 (N_14400,N_12834,N_13253);
nor U14401 (N_14401,N_13240,N_12241);
nor U14402 (N_14402,N_13271,N_13632);
xor U14403 (N_14403,N_13457,N_13164);
or U14404 (N_14404,N_12624,N_13763);
xnor U14405 (N_14405,N_13730,N_12666);
nor U14406 (N_14406,N_12017,N_12726);
and U14407 (N_14407,N_13404,N_13936);
xor U14408 (N_14408,N_12369,N_13264);
xor U14409 (N_14409,N_13378,N_12597);
and U14410 (N_14410,N_12622,N_13206);
or U14411 (N_14411,N_13218,N_13581);
xor U14412 (N_14412,N_13316,N_12783);
nor U14413 (N_14413,N_12604,N_13083);
xnor U14414 (N_14414,N_12160,N_13037);
nor U14415 (N_14415,N_13010,N_12190);
nand U14416 (N_14416,N_12641,N_13732);
nand U14417 (N_14417,N_13406,N_13943);
and U14418 (N_14418,N_12342,N_12752);
and U14419 (N_14419,N_12358,N_12921);
xnor U14420 (N_14420,N_13929,N_12880);
and U14421 (N_14421,N_13212,N_12485);
xor U14422 (N_14422,N_13711,N_12268);
and U14423 (N_14423,N_13673,N_13001);
and U14424 (N_14424,N_13084,N_12980);
and U14425 (N_14425,N_13729,N_12269);
and U14426 (N_14426,N_13921,N_12045);
and U14427 (N_14427,N_12249,N_13615);
nand U14428 (N_14428,N_12041,N_12279);
nor U14429 (N_14429,N_12655,N_13572);
xnor U14430 (N_14430,N_12081,N_13473);
and U14431 (N_14431,N_12621,N_12385);
nor U14432 (N_14432,N_12110,N_13215);
xnor U14433 (N_14433,N_13973,N_13878);
nand U14434 (N_14434,N_13105,N_12840);
xnor U14435 (N_14435,N_12809,N_13841);
and U14436 (N_14436,N_13488,N_12196);
nand U14437 (N_14437,N_12328,N_12938);
nor U14438 (N_14438,N_12730,N_13718);
and U14439 (N_14439,N_13634,N_12163);
or U14440 (N_14440,N_12516,N_12270);
and U14441 (N_14441,N_12590,N_13778);
or U14442 (N_14442,N_13691,N_12611);
and U14443 (N_14443,N_13169,N_13623);
or U14444 (N_14444,N_12109,N_12791);
xor U14445 (N_14445,N_13136,N_12721);
or U14446 (N_14446,N_12640,N_12594);
nor U14447 (N_14447,N_13706,N_12714);
xor U14448 (N_14448,N_13735,N_13191);
and U14449 (N_14449,N_13371,N_12614);
xor U14450 (N_14450,N_13815,N_13796);
or U14451 (N_14451,N_13683,N_12794);
and U14452 (N_14452,N_12155,N_12210);
and U14453 (N_14453,N_13233,N_13552);
and U14454 (N_14454,N_12728,N_13991);
and U14455 (N_14455,N_12309,N_12153);
and U14456 (N_14456,N_12892,N_13723);
and U14457 (N_14457,N_12962,N_12891);
or U14458 (N_14458,N_12020,N_13104);
nor U14459 (N_14459,N_12560,N_12368);
nor U14460 (N_14460,N_12776,N_12500);
xor U14461 (N_14461,N_12996,N_13970);
nor U14462 (N_14462,N_13466,N_13800);
nand U14463 (N_14463,N_12434,N_13666);
nor U14464 (N_14464,N_12979,N_12961);
nand U14465 (N_14465,N_12193,N_13207);
nor U14466 (N_14466,N_13924,N_12677);
xnor U14467 (N_14467,N_12871,N_13180);
xor U14468 (N_14468,N_12733,N_13586);
nand U14469 (N_14469,N_12283,N_12534);
nand U14470 (N_14470,N_12339,N_13542);
nor U14471 (N_14471,N_13832,N_12944);
nor U14472 (N_14472,N_13563,N_13589);
xnor U14473 (N_14473,N_12310,N_13339);
nand U14474 (N_14474,N_12697,N_13480);
nand U14475 (N_14475,N_13032,N_13108);
nor U14476 (N_14476,N_13722,N_12850);
and U14477 (N_14477,N_13419,N_12171);
and U14478 (N_14478,N_13453,N_12627);
nor U14479 (N_14479,N_13733,N_13469);
nor U14480 (N_14480,N_12387,N_12846);
nand U14481 (N_14481,N_12290,N_12983);
nor U14482 (N_14482,N_12837,N_12067);
nor U14483 (N_14483,N_13961,N_13151);
nor U14484 (N_14484,N_13154,N_13575);
and U14485 (N_14485,N_13304,N_13923);
and U14486 (N_14486,N_12380,N_12002);
and U14487 (N_14487,N_13583,N_13752);
nor U14488 (N_14488,N_12186,N_13232);
nor U14489 (N_14489,N_12620,N_13358);
and U14490 (N_14490,N_12522,N_13296);
and U14491 (N_14491,N_13277,N_13500);
nand U14492 (N_14492,N_12466,N_13147);
xor U14493 (N_14493,N_12736,N_12191);
xnor U14494 (N_14494,N_13073,N_13088);
or U14495 (N_14495,N_13594,N_12048);
and U14496 (N_14496,N_12603,N_13334);
xnor U14497 (N_14497,N_12384,N_12588);
and U14498 (N_14498,N_13485,N_13348);
and U14499 (N_14499,N_12770,N_13626);
xor U14500 (N_14500,N_13919,N_13762);
and U14501 (N_14501,N_12800,N_12833);
and U14502 (N_14502,N_13261,N_13134);
nor U14503 (N_14503,N_12495,N_13844);
or U14504 (N_14504,N_13978,N_13540);
or U14505 (N_14505,N_13054,N_12632);
nor U14506 (N_14506,N_13810,N_13432);
and U14507 (N_14507,N_13681,N_13315);
nor U14508 (N_14508,N_13302,N_12511);
xor U14509 (N_14509,N_13317,N_13056);
nand U14510 (N_14510,N_13561,N_12100);
or U14511 (N_14511,N_12120,N_12858);
nand U14512 (N_14512,N_12781,N_12046);
nand U14513 (N_14513,N_12373,N_13843);
xor U14514 (N_14514,N_13616,N_12589);
and U14515 (N_14515,N_12691,N_12499);
or U14516 (N_14516,N_12395,N_13864);
xor U14517 (N_14517,N_13562,N_12144);
or U14518 (N_14518,N_12719,N_13492);
xor U14519 (N_14519,N_12302,N_12447);
or U14520 (N_14520,N_12684,N_13532);
nand U14521 (N_14521,N_13067,N_12327);
or U14522 (N_14522,N_13166,N_12168);
nand U14523 (N_14523,N_12990,N_12013);
xnor U14524 (N_14524,N_13409,N_12448);
xnor U14525 (N_14525,N_12995,N_13489);
xnor U14526 (N_14526,N_12605,N_13351);
xor U14527 (N_14527,N_13647,N_13533);
nor U14528 (N_14528,N_13278,N_13908);
nand U14529 (N_14529,N_13817,N_13602);
nand U14530 (N_14530,N_12965,N_12223);
xor U14531 (N_14531,N_13015,N_12490);
and U14532 (N_14532,N_12883,N_12682);
or U14533 (N_14533,N_13307,N_12908);
and U14534 (N_14534,N_13968,N_12946);
xnor U14535 (N_14535,N_12897,N_13869);
and U14536 (N_14536,N_13177,N_13612);
nor U14537 (N_14537,N_13299,N_13305);
or U14538 (N_14538,N_13461,N_13521);
and U14539 (N_14539,N_13347,N_13112);
nor U14540 (N_14540,N_13040,N_13769);
or U14541 (N_14541,N_13538,N_13837);
or U14542 (N_14542,N_13100,N_12025);
nand U14543 (N_14543,N_13176,N_13880);
or U14544 (N_14544,N_13780,N_13337);
nor U14545 (N_14545,N_13987,N_13731);
and U14546 (N_14546,N_12349,N_12116);
nor U14547 (N_14547,N_13294,N_13721);
xor U14548 (N_14548,N_13370,N_12015);
nand U14549 (N_14549,N_13633,N_12716);
or U14550 (N_14550,N_13971,N_12737);
and U14551 (N_14551,N_13910,N_13357);
and U14552 (N_14552,N_12289,N_12209);
xnor U14553 (N_14553,N_13514,N_12412);
nand U14554 (N_14554,N_13999,N_13753);
and U14555 (N_14555,N_12104,N_12106);
or U14556 (N_14556,N_13543,N_13824);
nor U14557 (N_14557,N_12118,N_13526);
and U14558 (N_14558,N_12910,N_12075);
and U14559 (N_14559,N_13445,N_12295);
xor U14560 (N_14560,N_12319,N_12866);
or U14561 (N_14561,N_12699,N_12556);
nand U14562 (N_14562,N_13918,N_12755);
nand U14563 (N_14563,N_13303,N_12474);
nor U14564 (N_14564,N_12943,N_13491);
or U14565 (N_14565,N_12618,N_12743);
nor U14566 (N_14566,N_13280,N_13598);
and U14567 (N_14567,N_12663,N_12653);
and U14568 (N_14568,N_13905,N_12123);
xnor U14569 (N_14569,N_12656,N_12521);
nor U14570 (N_14570,N_12492,N_13192);
xor U14571 (N_14571,N_12935,N_13327);
xor U14572 (N_14572,N_13757,N_13713);
or U14573 (N_14573,N_12986,N_13564);
nor U14574 (N_14574,N_13941,N_12774);
xnor U14575 (N_14575,N_12475,N_12761);
nand U14576 (N_14576,N_13838,N_12889);
xnor U14577 (N_14577,N_12318,N_13606);
nor U14578 (N_14578,N_13297,N_13030);
or U14579 (N_14579,N_13179,N_12457);
and U14580 (N_14580,N_12117,N_13245);
nand U14581 (N_14581,N_12111,N_12574);
and U14582 (N_14582,N_13411,N_13306);
nand U14583 (N_14583,N_12226,N_13111);
xor U14584 (N_14584,N_12293,N_13648);
xnor U14585 (N_14585,N_13228,N_13890);
nand U14586 (N_14586,N_13183,N_12023);
or U14587 (N_14587,N_13595,N_13367);
or U14588 (N_14588,N_12098,N_13031);
xor U14589 (N_14589,N_13736,N_13835);
or U14590 (N_14590,N_13579,N_12211);
xor U14591 (N_14591,N_12112,N_12479);
xnor U14592 (N_14592,N_12581,N_12480);
xor U14593 (N_14593,N_13963,N_13811);
and U14594 (N_14594,N_13002,N_12101);
and U14595 (N_14595,N_12503,N_12399);
nand U14596 (N_14596,N_12525,N_13019);
and U14597 (N_14597,N_13801,N_12749);
or U14598 (N_14598,N_13279,N_12431);
nand U14599 (N_14599,N_13156,N_12824);
or U14600 (N_14600,N_12904,N_13599);
nand U14601 (N_14601,N_12598,N_13313);
and U14602 (N_14602,N_12281,N_12602);
nand U14603 (N_14603,N_13173,N_13523);
and U14604 (N_14604,N_12134,N_13909);
nor U14605 (N_14605,N_13836,N_13379);
xor U14606 (N_14606,N_13871,N_12902);
nor U14607 (N_14607,N_13066,N_12251);
xnor U14608 (N_14608,N_13983,N_13663);
and U14609 (N_14609,N_12524,N_13446);
nor U14610 (N_14610,N_13754,N_13465);
nor U14611 (N_14611,N_12359,N_13150);
xor U14612 (N_14612,N_12459,N_12414);
or U14613 (N_14613,N_13326,N_13063);
or U14614 (N_14614,N_12311,N_13171);
xnor U14615 (N_14615,N_12400,N_13571);
nand U14616 (N_14616,N_13341,N_12389);
or U14617 (N_14617,N_12089,N_13748);
xor U14618 (N_14618,N_12263,N_13497);
xor U14619 (N_14619,N_13901,N_13653);
nor U14620 (N_14620,N_12723,N_13819);
xor U14621 (N_14621,N_13072,N_13677);
xor U14622 (N_14622,N_13792,N_12472);
or U14623 (N_14623,N_13467,N_13050);
nor U14624 (N_14624,N_13374,N_13178);
nor U14625 (N_14625,N_12420,N_12264);
xor U14626 (N_14626,N_13822,N_13423);
or U14627 (N_14627,N_12764,N_13265);
and U14628 (N_14628,N_12416,N_12178);
nand U14629 (N_14629,N_13895,N_12224);
nor U14630 (N_14630,N_12984,N_12877);
nor U14631 (N_14631,N_13275,N_12949);
and U14632 (N_14632,N_13274,N_13333);
nor U14633 (N_14633,N_13258,N_12308);
nand U14634 (N_14634,N_13857,N_12572);
and U14635 (N_14635,N_12364,N_12722);
xnor U14636 (N_14636,N_13153,N_12356);
and U14637 (N_14637,N_13387,N_12482);
and U14638 (N_14638,N_12571,N_12271);
and U14639 (N_14639,N_12021,N_12754);
nand U14640 (N_14640,N_12243,N_12361);
or U14641 (N_14641,N_13463,N_12739);
nand U14642 (N_14642,N_13989,N_12615);
and U14643 (N_14643,N_12039,N_12587);
and U14644 (N_14644,N_12732,N_13130);
xnor U14645 (N_14645,N_12905,N_12796);
nand U14646 (N_14646,N_13366,N_13013);
xnor U14647 (N_14647,N_13544,N_13239);
xor U14648 (N_14648,N_12718,N_12182);
nand U14649 (N_14649,N_12252,N_12626);
nand U14650 (N_14650,N_13834,N_12585);
nor U14651 (N_14651,N_13771,N_13234);
or U14652 (N_14652,N_12004,N_13295);
nand U14653 (N_14653,N_13170,N_12300);
and U14654 (N_14654,N_13707,N_13506);
and U14655 (N_14655,N_13520,N_12564);
nor U14656 (N_14656,N_13203,N_12864);
or U14657 (N_14657,N_13712,N_13281);
nor U14658 (N_14658,N_13636,N_12913);
or U14659 (N_14659,N_13414,N_12920);
or U14660 (N_14660,N_13509,N_12586);
nor U14661 (N_14661,N_13872,N_12198);
or U14662 (N_14662,N_12232,N_12207);
and U14663 (N_14663,N_12079,N_12206);
xnor U14664 (N_14664,N_13755,N_12994);
and U14665 (N_14665,N_12114,N_13960);
and U14666 (N_14666,N_12355,N_13812);
or U14667 (N_14667,N_13969,N_12528);
xnor U14668 (N_14668,N_12593,N_12330);
or U14669 (N_14669,N_13470,N_12063);
nand U14670 (N_14670,N_12662,N_12881);
nand U14671 (N_14671,N_13740,N_12394);
nand U14672 (N_14672,N_12847,N_12667);
nor U14673 (N_14673,N_12900,N_13093);
nor U14674 (N_14674,N_12964,N_12887);
nor U14675 (N_14675,N_12766,N_12685);
xor U14676 (N_14676,N_13021,N_12445);
nand U14677 (N_14677,N_12398,N_13097);
nor U14678 (N_14678,N_12070,N_12146);
nand U14679 (N_14679,N_13794,N_12218);
nor U14680 (N_14680,N_13016,N_12545);
xor U14681 (N_14681,N_13675,N_12712);
xor U14682 (N_14682,N_12404,N_13842);
and U14683 (N_14683,N_12952,N_12037);
nor U14684 (N_14684,N_12817,N_12014);
and U14685 (N_14685,N_12925,N_13927);
nor U14686 (N_14686,N_13360,N_12172);
or U14687 (N_14687,N_13394,N_12150);
or U14688 (N_14688,N_13146,N_13979);
xnor U14689 (N_14689,N_13222,N_13287);
nand U14690 (N_14690,N_12255,N_13172);
and U14691 (N_14691,N_12234,N_13840);
nand U14692 (N_14692,N_12159,N_13161);
nor U14693 (N_14693,N_13186,N_12301);
xnor U14694 (N_14694,N_12227,N_12306);
nor U14695 (N_14695,N_13635,N_12470);
nand U14696 (N_14696,N_13996,N_13308);
or U14697 (N_14697,N_12239,N_12748);
nor U14698 (N_14698,N_13892,N_13007);
nor U14699 (N_14699,N_13332,N_13935);
nand U14700 (N_14700,N_13395,N_12261);
xnor U14701 (N_14701,N_12750,N_12780);
or U14702 (N_14702,N_12376,N_12582);
xnor U14703 (N_14703,N_12873,N_13685);
and U14704 (N_14704,N_12065,N_12544);
nand U14705 (N_14705,N_13529,N_13219);
or U14706 (N_14706,N_12220,N_12975);
and U14707 (N_14707,N_13894,N_12325);
nor U14708 (N_14708,N_13966,N_12405);
nor U14709 (N_14709,N_12421,N_12808);
or U14710 (N_14710,N_13679,N_12044);
xor U14711 (N_14711,N_13850,N_13643);
nand U14712 (N_14712,N_12128,N_13656);
or U14713 (N_14713,N_13899,N_12502);
or U14714 (N_14714,N_12689,N_13928);
nor U14715 (N_14715,N_13126,N_12762);
or U14716 (N_14716,N_12901,N_12982);
and U14717 (N_14717,N_13202,N_13505);
and U14718 (N_14718,N_13243,N_13119);
nor U14719 (N_14719,N_13879,N_13770);
nor U14720 (N_14720,N_12997,N_13214);
nor U14721 (N_14721,N_13873,N_12324);
nand U14722 (N_14722,N_12520,N_12778);
or U14723 (N_14723,N_12763,N_12099);
and U14724 (N_14724,N_13867,N_12133);
or U14725 (N_14725,N_12555,N_13985);
and U14726 (N_14726,N_13204,N_12686);
xnor U14727 (N_14727,N_12338,N_12836);
or U14728 (N_14728,N_12693,N_12933);
nor U14729 (N_14729,N_12085,N_13863);
xnor U14730 (N_14730,N_12888,N_13962);
xor U14731 (N_14731,N_13702,N_13965);
xor U14732 (N_14732,N_12007,N_12139);
nand U14733 (N_14733,N_12985,N_13369);
xnor U14734 (N_14734,N_12812,N_12135);
and U14735 (N_14735,N_12771,N_12509);
xnor U14736 (N_14736,N_13516,N_12184);
and U14737 (N_14737,N_12856,N_12493);
and U14738 (N_14738,N_12885,N_12806);
or U14739 (N_14739,N_13859,N_12498);
or U14740 (N_14740,N_12064,N_13797);
nand U14741 (N_14741,N_13205,N_13917);
or U14742 (N_14742,N_13700,N_12643);
nand U14743 (N_14743,N_12294,N_12137);
or U14744 (N_14744,N_13459,N_12321);
nand U14745 (N_14745,N_12247,N_13188);
nor U14746 (N_14746,N_12245,N_12652);
xor U14747 (N_14747,N_13715,N_12827);
and U14748 (N_14748,N_13355,N_12600);
nor U14749 (N_14749,N_12890,N_12452);
xor U14750 (N_14750,N_12061,N_13255);
xnor U14751 (N_14751,N_13637,N_12273);
xor U14752 (N_14752,N_13992,N_12676);
or U14753 (N_14753,N_12221,N_13550);
and U14754 (N_14754,N_13127,N_12397);
nand U14755 (N_14755,N_13967,N_12678);
xor U14756 (N_14756,N_13399,N_13830);
nor U14757 (N_14757,N_13425,N_13257);
or U14758 (N_14758,N_12147,N_12759);
and U14759 (N_14759,N_12845,N_13591);
nor U14760 (N_14760,N_13060,N_13896);
nor U14761 (N_14761,N_12899,N_12894);
xor U14762 (N_14762,N_12483,N_12177);
nor U14763 (N_14763,N_12988,N_12496);
nor U14764 (N_14764,N_13324,N_13322);
and U14765 (N_14765,N_13660,N_12115);
or U14766 (N_14766,N_12244,N_12401);
and U14767 (N_14767,N_12947,N_13070);
or U14768 (N_14768,N_13674,N_12497);
and U14769 (N_14769,N_13217,N_12884);
or U14770 (N_14770,N_12741,N_12543);
xnor U14771 (N_14771,N_13820,N_13725);
or U14772 (N_14772,N_12423,N_13375);
xnor U14773 (N_14773,N_13047,N_13775);
or U14774 (N_14774,N_13132,N_13750);
or U14775 (N_14775,N_13211,N_12551);
nor U14776 (N_14776,N_12430,N_13197);
nor U14777 (N_14777,N_12329,N_12708);
or U14778 (N_14778,N_12740,N_13323);
xnor U14779 (N_14779,N_12299,N_13174);
or U14780 (N_14780,N_12619,N_12458);
and U14781 (N_14781,N_12711,N_12231);
and U14782 (N_14782,N_12322,N_12413);
and U14783 (N_14783,N_12672,N_13501);
or U14784 (N_14784,N_12578,N_12924);
and U14785 (N_14785,N_12637,N_12202);
and U14786 (N_14786,N_12974,N_13881);
nand U14787 (N_14787,N_13625,N_13381);
nand U14788 (N_14788,N_12546,N_13213);
xor U14789 (N_14789,N_12768,N_13887);
nand U14790 (N_14790,N_13536,N_12742);
and U14791 (N_14791,N_13948,N_12782);
xnor U14792 (N_14792,N_13827,N_12701);
nand U14793 (N_14793,N_12165,N_12005);
nor U14794 (N_14794,N_12843,N_13759);
nand U14795 (N_14795,N_13694,N_13655);
and U14796 (N_14796,N_12688,N_12248);
xor U14797 (N_14797,N_12370,N_13472);
nor U14798 (N_14798,N_13384,N_13014);
nand U14799 (N_14799,N_13115,N_13607);
nor U14800 (N_14800,N_13065,N_12407);
xor U14801 (N_14801,N_13053,N_12233);
nor U14802 (N_14802,N_12194,N_13952);
and U14803 (N_14803,N_13135,N_12596);
nor U14804 (N_14804,N_13695,N_12442);
nor U14805 (N_14805,N_12084,N_12951);
and U14806 (N_14806,N_13774,N_13984);
and U14807 (N_14807,N_12266,N_12638);
or U14808 (N_14808,N_13670,N_13310);
and U14809 (N_14809,N_12993,N_13698);
xnor U14810 (N_14810,N_12735,N_12166);
nor U14811 (N_14811,N_13330,N_13460);
nor U14812 (N_14812,N_12746,N_12003);
nand U14813 (N_14813,N_12914,N_12136);
or U14814 (N_14814,N_12415,N_13110);
nand U14815 (N_14815,N_13667,N_12786);
nor U14816 (N_14816,N_13658,N_13503);
nor U14817 (N_14817,N_13148,N_13508);
or U14818 (N_14818,N_12346,N_12882);
nor U14819 (N_14819,N_13035,N_12032);
or U14820 (N_14820,N_12795,N_13669);
nand U14821 (N_14821,N_12467,N_12435);
and U14822 (N_14822,N_13392,N_12408);
xnor U14823 (N_14823,N_12476,N_12599);
nor U14824 (N_14824,N_13124,N_12463);
or U14825 (N_14825,N_13738,N_12510);
xnor U14826 (N_14826,N_13684,N_13994);
xnor U14827 (N_14827,N_12253,N_12612);
xnor U14828 (N_14828,N_12683,N_12530);
and U14829 (N_14829,N_13190,N_13955);
nor U14830 (N_14830,N_12313,N_13167);
xor U14831 (N_14831,N_13125,N_13621);
nor U14832 (N_14832,N_13959,N_12124);
or U14833 (N_14833,N_12040,N_13314);
nand U14834 (N_14834,N_12181,N_12610);
nor U14835 (N_14835,N_12108,N_13338);
and U14836 (N_14836,N_13442,N_12312);
or U14837 (N_14837,N_13221,N_13576);
nor U14838 (N_14838,N_13727,N_13343);
or U14839 (N_14839,N_13226,N_12861);
xor U14840 (N_14840,N_13023,N_12323);
and U14841 (N_14841,N_12647,N_13692);
nor U14842 (N_14842,N_12141,N_12006);
nand U14843 (N_14843,N_12288,N_13531);
and U14844 (N_14844,N_12554,N_12000);
or U14845 (N_14845,N_13746,N_12704);
xor U14846 (N_14846,N_12815,N_13200);
nand U14847 (N_14847,N_12506,N_13256);
xnor U14848 (N_14848,N_12454,N_13949);
nand U14849 (N_14849,N_12583,N_12348);
nor U14850 (N_14850,N_13129,N_12030);
nor U14851 (N_14851,N_12449,N_13175);
and U14852 (N_14852,N_13528,N_12922);
nand U14853 (N_14853,N_13926,N_12393);
and U14854 (N_14854,N_12340,N_12345);
nor U14855 (N_14855,N_12262,N_12409);
and U14856 (N_14856,N_13846,N_12915);
or U14857 (N_14857,N_13095,N_13045);
or U14858 (N_14858,N_12784,N_12130);
and U14859 (N_14859,N_13435,N_13779);
nand U14860 (N_14860,N_13565,N_12229);
and U14861 (N_14861,N_13241,N_13091);
nand U14862 (N_14862,N_13765,N_12565);
and U14863 (N_14863,N_13353,N_12561);
or U14864 (N_14864,N_13020,N_12315);
nand U14865 (N_14865,N_12876,N_12173);
or U14866 (N_14866,N_13198,N_13566);
and U14867 (N_14867,N_12963,N_13588);
and U14868 (N_14868,N_13882,N_13012);
nor U14869 (N_14869,N_12341,N_12419);
nand U14870 (N_14870,N_12274,N_12278);
and U14871 (N_14871,N_12927,N_12071);
and U14872 (N_14872,N_13889,N_13410);
nor U14873 (N_14873,N_12645,N_12228);
xnor U14874 (N_14874,N_13080,N_13587);
nor U14875 (N_14875,N_12853,N_12080);
nor U14876 (N_14876,N_13627,N_13862);
nand U14877 (N_14877,N_12703,N_12838);
nor U14878 (N_14878,N_13490,N_13268);
or U14879 (N_14879,N_13185,N_13408);
nor U14880 (N_14880,N_12019,N_13494);
xor U14881 (N_14881,N_13714,N_12819);
or U14882 (N_14882,N_12464,N_13568);
or U14883 (N_14883,N_12154,N_12852);
nand U14884 (N_14884,N_13773,N_13831);
and U14885 (N_14885,N_13545,N_13557);
or U14886 (N_14886,N_13601,N_13608);
nor U14887 (N_14887,N_12201,N_13209);
nor U14888 (N_14888,N_13468,N_12681);
and U14889 (N_14889,N_12954,N_12379);
and U14890 (N_14890,N_13041,N_12161);
nor U14891 (N_14891,N_13808,N_13716);
nor U14892 (N_14892,N_13527,N_12939);
xor U14893 (N_14893,N_12959,N_12143);
or U14894 (N_14894,N_13201,N_13138);
nand U14895 (N_14895,N_13157,N_12456);
or U14896 (N_14896,N_12999,N_13798);
nand U14897 (N_14897,N_13577,N_12250);
xor U14898 (N_14898,N_12107,N_13502);
nor U14899 (N_14899,N_12553,N_13270);
nor U14900 (N_14900,N_13630,N_13131);
and U14901 (N_14901,N_12334,N_12950);
xnor U14902 (N_14902,N_13230,N_12540);
or U14903 (N_14903,N_12694,N_13903);
or U14904 (N_14904,N_12724,N_12695);
nand U14905 (N_14905,N_12674,N_13482);
xor U14906 (N_14906,N_13876,N_13345);
nand U14907 (N_14907,N_13783,N_13697);
nand U14908 (N_14908,N_13839,N_12552);
and U14909 (N_14909,N_12059,N_13102);
or U14910 (N_14910,N_13424,N_12417);
nor U14911 (N_14911,N_12631,N_13997);
or U14912 (N_14912,N_13349,N_13099);
and U14913 (N_14913,N_12438,N_12386);
nor U14914 (N_14914,N_12157,N_13728);
xnor U14915 (N_14915,N_12745,N_13155);
xnor U14916 (N_14916,N_12486,N_12957);
or U14917 (N_14917,N_12320,N_13120);
or U14918 (N_14918,N_12535,N_12859);
xor U14919 (N_14919,N_13474,N_12860);
xor U14920 (N_14920,N_12820,N_13137);
and U14921 (N_14921,N_12822,N_12705);
or U14922 (N_14922,N_13114,N_13018);
nor U14923 (N_14923,N_13252,N_13311);
or U14924 (N_14924,N_12131,N_12052);
nor U14925 (N_14925,N_13619,N_13530);
nor U14926 (N_14926,N_13415,N_12895);
or U14927 (N_14927,N_12192,N_13434);
xor U14928 (N_14928,N_13283,N_13522);
nand U14929 (N_14929,N_13356,N_12788);
nor U14930 (N_14930,N_13851,N_13807);
nor U14931 (N_14931,N_12803,N_13036);
xor U14932 (N_14932,N_12083,N_12267);
nand U14933 (N_14933,N_12222,N_13184);
and U14934 (N_14934,N_13106,N_13196);
or U14935 (N_14935,N_13398,N_12801);
nand U14936 (N_14936,N_12350,N_13772);
nor U14937 (N_14937,N_12537,N_13439);
nor U14938 (N_14938,N_13033,N_13383);
nand U14939 (N_14939,N_13693,N_12613);
nand U14940 (N_14940,N_12352,N_12660);
nor U14941 (N_14941,N_13011,N_12372);
nand U14942 (N_14942,N_13570,N_12297);
nor U14943 (N_14943,N_13618,N_13578);
nor U14944 (N_14944,N_13548,N_12709);
or U14945 (N_14945,N_12538,N_12608);
nor U14946 (N_14946,N_12187,N_13477);
and U14947 (N_14947,N_12765,N_13319);
or U14948 (N_14948,N_13609,N_13098);
nand U14949 (N_14949,N_12911,N_12584);
nor U14950 (N_14950,N_12923,N_13884);
and U14951 (N_14951,N_12875,N_12468);
and U14952 (N_14952,N_13853,N_13139);
and U14953 (N_14953,N_12307,N_13400);
nor U14954 (N_14954,N_12093,N_13661);
nand U14955 (N_14955,N_13352,N_12696);
nor U14956 (N_14956,N_12508,N_12729);
and U14957 (N_14957,N_12149,N_13668);
or U14958 (N_14958,N_12872,N_12219);
and U14959 (N_14959,N_12960,N_12969);
xnor U14960 (N_14960,N_13412,N_12305);
and U14961 (N_14961,N_13143,N_13077);
and U14962 (N_14962,N_13593,N_13874);
or U14963 (N_14963,N_13620,N_13708);
nor U14964 (N_14964,N_13737,N_13389);
xnor U14965 (N_14965,N_13034,N_13883);
xnor U14966 (N_14966,N_12440,N_13933);
and U14967 (N_14967,N_12907,N_12256);
nand U14968 (N_14968,N_13784,N_13042);
and U14969 (N_14969,N_12151,N_13359);
or U14970 (N_14970,N_12798,N_12204);
xnor U14971 (N_14971,N_13455,N_12539);
xnor U14972 (N_14972,N_13140,N_13988);
xnor U14973 (N_14973,N_12702,N_13433);
and U14974 (N_14974,N_12931,N_13758);
nor U14975 (N_14975,N_12835,N_12802);
nor U14976 (N_14976,N_13744,N_13766);
nor U14977 (N_14977,N_13309,N_13285);
or U14978 (N_14978,N_12170,N_13248);
xor U14979 (N_14979,N_12991,N_13061);
and U14980 (N_14980,N_12383,N_12945);
nor U14981 (N_14981,N_12238,N_12148);
xor U14982 (N_14982,N_12377,N_12200);
or U14983 (N_14983,N_12217,N_13000);
xor U14984 (N_14984,N_12507,N_13026);
nand U14985 (N_14985,N_12592,N_13573);
xnor U14986 (N_14986,N_13951,N_12060);
nand U14987 (N_14987,N_13075,N_12558);
nand U14988 (N_14988,N_13336,N_13855);
xnor U14989 (N_14989,N_12169,N_13259);
and U14990 (N_14990,N_12777,N_12375);
nor U14991 (N_14991,N_12854,N_13403);
or U14992 (N_14992,N_13931,N_13622);
nand U14993 (N_14993,N_12236,N_13875);
nand U14994 (N_14994,N_12335,N_13678);
and U14995 (N_14995,N_12855,N_12523);
nor U14996 (N_14996,N_13462,N_13428);
or U14997 (N_14997,N_13009,N_12898);
or U14998 (N_14998,N_12208,N_12230);
nor U14999 (N_14999,N_13944,N_13039);
nor U15000 (N_15000,N_12137,N_12405);
xor U15001 (N_15001,N_13219,N_13839);
xor U15002 (N_15002,N_13043,N_12862);
nand U15003 (N_15003,N_12429,N_12920);
or U15004 (N_15004,N_13988,N_12878);
and U15005 (N_15005,N_12767,N_12715);
or U15006 (N_15006,N_13685,N_12025);
nand U15007 (N_15007,N_13990,N_13128);
nor U15008 (N_15008,N_13654,N_12766);
or U15009 (N_15009,N_13096,N_13789);
xnor U15010 (N_15010,N_12593,N_13452);
or U15011 (N_15011,N_13208,N_13618);
nor U15012 (N_15012,N_12702,N_13185);
nor U15013 (N_15013,N_13785,N_12627);
or U15014 (N_15014,N_13934,N_12180);
xor U15015 (N_15015,N_12403,N_13929);
nand U15016 (N_15016,N_12524,N_12646);
nand U15017 (N_15017,N_12271,N_13448);
nand U15018 (N_15018,N_12084,N_13072);
or U15019 (N_15019,N_12264,N_12209);
nand U15020 (N_15020,N_13872,N_12321);
or U15021 (N_15021,N_13485,N_13731);
and U15022 (N_15022,N_13965,N_12211);
nor U15023 (N_15023,N_13433,N_12402);
and U15024 (N_15024,N_12664,N_12675);
or U15025 (N_15025,N_12248,N_13710);
nand U15026 (N_15026,N_13892,N_12589);
xnor U15027 (N_15027,N_13220,N_12975);
nor U15028 (N_15028,N_12417,N_13415);
xor U15029 (N_15029,N_12682,N_13047);
nand U15030 (N_15030,N_12720,N_12191);
xor U15031 (N_15031,N_12113,N_12007);
and U15032 (N_15032,N_12527,N_13560);
and U15033 (N_15033,N_13363,N_13335);
or U15034 (N_15034,N_12672,N_13368);
nor U15035 (N_15035,N_12504,N_13793);
or U15036 (N_15036,N_13570,N_12497);
nor U15037 (N_15037,N_13009,N_12566);
and U15038 (N_15038,N_13250,N_13293);
nor U15039 (N_15039,N_13521,N_13870);
nor U15040 (N_15040,N_12714,N_12793);
nor U15041 (N_15041,N_12042,N_12654);
and U15042 (N_15042,N_12043,N_12977);
xor U15043 (N_15043,N_12223,N_12529);
nor U15044 (N_15044,N_13793,N_13175);
nand U15045 (N_15045,N_12096,N_13788);
nand U15046 (N_15046,N_12328,N_13762);
and U15047 (N_15047,N_12000,N_12488);
and U15048 (N_15048,N_13633,N_13043);
nor U15049 (N_15049,N_12532,N_12737);
nand U15050 (N_15050,N_13968,N_12260);
or U15051 (N_15051,N_12510,N_12589);
nand U15052 (N_15052,N_12795,N_13106);
and U15053 (N_15053,N_13249,N_12511);
nor U15054 (N_15054,N_12257,N_12282);
and U15055 (N_15055,N_12127,N_12303);
nand U15056 (N_15056,N_12465,N_12091);
xor U15057 (N_15057,N_13629,N_12707);
nand U15058 (N_15058,N_13394,N_12158);
and U15059 (N_15059,N_13965,N_13437);
xnor U15060 (N_15060,N_13726,N_12314);
nand U15061 (N_15061,N_13660,N_13097);
or U15062 (N_15062,N_12856,N_12344);
nor U15063 (N_15063,N_12707,N_13315);
xnor U15064 (N_15064,N_13871,N_12052);
and U15065 (N_15065,N_12635,N_12964);
and U15066 (N_15066,N_12555,N_12648);
and U15067 (N_15067,N_13569,N_13969);
or U15068 (N_15068,N_12260,N_13004);
nand U15069 (N_15069,N_13385,N_13821);
nand U15070 (N_15070,N_12124,N_12988);
or U15071 (N_15071,N_12595,N_12587);
or U15072 (N_15072,N_12058,N_13869);
or U15073 (N_15073,N_12428,N_12271);
nand U15074 (N_15074,N_12915,N_13278);
xnor U15075 (N_15075,N_13984,N_12137);
or U15076 (N_15076,N_12114,N_12261);
nand U15077 (N_15077,N_12031,N_12091);
nand U15078 (N_15078,N_12240,N_13728);
or U15079 (N_15079,N_12510,N_12846);
and U15080 (N_15080,N_12742,N_12519);
and U15081 (N_15081,N_13983,N_13795);
or U15082 (N_15082,N_13421,N_13627);
or U15083 (N_15083,N_13818,N_12731);
nand U15084 (N_15084,N_12270,N_13677);
nor U15085 (N_15085,N_12544,N_13252);
nor U15086 (N_15086,N_13457,N_12917);
xor U15087 (N_15087,N_12522,N_13999);
xnor U15088 (N_15088,N_13468,N_13679);
and U15089 (N_15089,N_12920,N_12922);
and U15090 (N_15090,N_13649,N_12876);
xnor U15091 (N_15091,N_13304,N_12078);
or U15092 (N_15092,N_13482,N_13417);
nor U15093 (N_15093,N_13979,N_12951);
nand U15094 (N_15094,N_12768,N_13525);
and U15095 (N_15095,N_13632,N_13330);
nor U15096 (N_15096,N_12644,N_12970);
xnor U15097 (N_15097,N_13684,N_13117);
nand U15098 (N_15098,N_13710,N_12091);
nand U15099 (N_15099,N_13731,N_13803);
nor U15100 (N_15100,N_13530,N_13634);
and U15101 (N_15101,N_13902,N_12180);
xor U15102 (N_15102,N_13272,N_12200);
nand U15103 (N_15103,N_12686,N_13659);
and U15104 (N_15104,N_12183,N_12347);
xor U15105 (N_15105,N_12145,N_12163);
or U15106 (N_15106,N_13336,N_13988);
xnor U15107 (N_15107,N_12664,N_12358);
and U15108 (N_15108,N_13072,N_13544);
nor U15109 (N_15109,N_13070,N_12506);
nor U15110 (N_15110,N_13788,N_12358);
nor U15111 (N_15111,N_12938,N_12735);
or U15112 (N_15112,N_12157,N_13878);
nand U15113 (N_15113,N_12915,N_13903);
nand U15114 (N_15114,N_13981,N_12073);
nor U15115 (N_15115,N_13557,N_12512);
or U15116 (N_15116,N_12911,N_12356);
or U15117 (N_15117,N_12664,N_13107);
nor U15118 (N_15118,N_12290,N_12782);
and U15119 (N_15119,N_13764,N_13646);
nand U15120 (N_15120,N_12026,N_13102);
nand U15121 (N_15121,N_12615,N_13686);
nand U15122 (N_15122,N_13785,N_12670);
or U15123 (N_15123,N_13161,N_13408);
and U15124 (N_15124,N_12493,N_13886);
nor U15125 (N_15125,N_13665,N_13353);
or U15126 (N_15126,N_13134,N_13856);
and U15127 (N_15127,N_13435,N_12332);
or U15128 (N_15128,N_13556,N_12010);
nand U15129 (N_15129,N_12057,N_12134);
xnor U15130 (N_15130,N_12794,N_12485);
nand U15131 (N_15131,N_13261,N_13628);
nor U15132 (N_15132,N_13132,N_12877);
nand U15133 (N_15133,N_12444,N_13197);
and U15134 (N_15134,N_13740,N_12057);
and U15135 (N_15135,N_13711,N_13292);
xor U15136 (N_15136,N_12685,N_12879);
or U15137 (N_15137,N_12837,N_12017);
nand U15138 (N_15138,N_13574,N_13947);
or U15139 (N_15139,N_13531,N_12514);
and U15140 (N_15140,N_12378,N_12880);
nand U15141 (N_15141,N_13562,N_13049);
or U15142 (N_15142,N_13352,N_12224);
and U15143 (N_15143,N_12298,N_13357);
nand U15144 (N_15144,N_12197,N_13741);
nand U15145 (N_15145,N_12996,N_12437);
nand U15146 (N_15146,N_13778,N_13274);
xor U15147 (N_15147,N_13404,N_13300);
or U15148 (N_15148,N_12717,N_12027);
or U15149 (N_15149,N_12395,N_12178);
nand U15150 (N_15150,N_13925,N_12312);
xor U15151 (N_15151,N_13814,N_12643);
nand U15152 (N_15152,N_13200,N_12068);
or U15153 (N_15153,N_13032,N_13216);
xnor U15154 (N_15154,N_12134,N_12418);
nor U15155 (N_15155,N_13172,N_13159);
nand U15156 (N_15156,N_13859,N_13221);
nand U15157 (N_15157,N_12539,N_13917);
nor U15158 (N_15158,N_12688,N_12559);
and U15159 (N_15159,N_13980,N_12772);
and U15160 (N_15160,N_12919,N_13504);
nand U15161 (N_15161,N_12320,N_12930);
and U15162 (N_15162,N_13726,N_13011);
and U15163 (N_15163,N_13036,N_13049);
or U15164 (N_15164,N_13525,N_13211);
or U15165 (N_15165,N_12994,N_12387);
nor U15166 (N_15166,N_13317,N_12999);
and U15167 (N_15167,N_12973,N_13035);
nand U15168 (N_15168,N_13347,N_13291);
xor U15169 (N_15169,N_12156,N_12550);
nand U15170 (N_15170,N_12236,N_12668);
and U15171 (N_15171,N_12432,N_12166);
or U15172 (N_15172,N_12091,N_13803);
nand U15173 (N_15173,N_12828,N_12086);
or U15174 (N_15174,N_13280,N_12166);
nor U15175 (N_15175,N_13112,N_12718);
xor U15176 (N_15176,N_13692,N_12796);
nand U15177 (N_15177,N_12043,N_12497);
nor U15178 (N_15178,N_12695,N_13163);
or U15179 (N_15179,N_13552,N_13971);
and U15180 (N_15180,N_12354,N_12106);
xor U15181 (N_15181,N_12861,N_13648);
xnor U15182 (N_15182,N_13323,N_13597);
xor U15183 (N_15183,N_13322,N_12602);
xor U15184 (N_15184,N_12963,N_12507);
nand U15185 (N_15185,N_13483,N_12400);
or U15186 (N_15186,N_13444,N_13351);
xor U15187 (N_15187,N_13331,N_13002);
nand U15188 (N_15188,N_13147,N_13380);
xnor U15189 (N_15189,N_12591,N_13873);
or U15190 (N_15190,N_12506,N_13935);
nand U15191 (N_15191,N_13506,N_12763);
nand U15192 (N_15192,N_13449,N_13290);
nand U15193 (N_15193,N_13180,N_12670);
and U15194 (N_15194,N_12406,N_13928);
xor U15195 (N_15195,N_12422,N_12031);
nor U15196 (N_15196,N_12271,N_12024);
or U15197 (N_15197,N_13631,N_12628);
or U15198 (N_15198,N_12775,N_13669);
and U15199 (N_15199,N_13926,N_13235);
nand U15200 (N_15200,N_12716,N_13663);
or U15201 (N_15201,N_12816,N_13353);
or U15202 (N_15202,N_13967,N_12043);
xnor U15203 (N_15203,N_13590,N_12100);
nand U15204 (N_15204,N_12722,N_13277);
nor U15205 (N_15205,N_12826,N_12028);
and U15206 (N_15206,N_13363,N_12888);
xnor U15207 (N_15207,N_13151,N_13505);
or U15208 (N_15208,N_13181,N_13425);
nand U15209 (N_15209,N_12814,N_12957);
nor U15210 (N_15210,N_13105,N_12986);
nand U15211 (N_15211,N_12820,N_13859);
nor U15212 (N_15212,N_13302,N_12469);
nand U15213 (N_15213,N_13189,N_12977);
nand U15214 (N_15214,N_13678,N_13465);
xor U15215 (N_15215,N_13393,N_12504);
nand U15216 (N_15216,N_13982,N_13746);
nand U15217 (N_15217,N_12996,N_13475);
xor U15218 (N_15218,N_12682,N_12311);
and U15219 (N_15219,N_13622,N_12415);
nor U15220 (N_15220,N_12822,N_12977);
or U15221 (N_15221,N_13320,N_13390);
or U15222 (N_15222,N_13175,N_13895);
nand U15223 (N_15223,N_13167,N_12903);
or U15224 (N_15224,N_12011,N_12713);
xnor U15225 (N_15225,N_12186,N_13456);
xnor U15226 (N_15226,N_12703,N_13262);
or U15227 (N_15227,N_12467,N_13378);
nor U15228 (N_15228,N_13392,N_12353);
and U15229 (N_15229,N_12438,N_12341);
xor U15230 (N_15230,N_12430,N_13834);
or U15231 (N_15231,N_13361,N_12806);
nand U15232 (N_15232,N_13333,N_12101);
and U15233 (N_15233,N_12796,N_13162);
nand U15234 (N_15234,N_12300,N_12540);
xor U15235 (N_15235,N_12568,N_12829);
nor U15236 (N_15236,N_13829,N_13994);
nand U15237 (N_15237,N_13882,N_12017);
or U15238 (N_15238,N_12018,N_13058);
xor U15239 (N_15239,N_12628,N_12252);
xor U15240 (N_15240,N_13144,N_12427);
and U15241 (N_15241,N_13236,N_13679);
nand U15242 (N_15242,N_12146,N_13064);
nor U15243 (N_15243,N_13787,N_12991);
nand U15244 (N_15244,N_13615,N_13899);
xnor U15245 (N_15245,N_13568,N_13702);
and U15246 (N_15246,N_12319,N_12364);
and U15247 (N_15247,N_12403,N_13422);
and U15248 (N_15248,N_13272,N_12187);
nand U15249 (N_15249,N_12168,N_13941);
xnor U15250 (N_15250,N_12107,N_12938);
nand U15251 (N_15251,N_13417,N_13748);
xnor U15252 (N_15252,N_12315,N_12544);
xnor U15253 (N_15253,N_12396,N_12709);
or U15254 (N_15254,N_12116,N_12030);
nand U15255 (N_15255,N_12938,N_13609);
nor U15256 (N_15256,N_12154,N_13714);
xnor U15257 (N_15257,N_12710,N_13009);
nor U15258 (N_15258,N_13745,N_12267);
nand U15259 (N_15259,N_13815,N_13097);
and U15260 (N_15260,N_13193,N_13526);
and U15261 (N_15261,N_12765,N_13973);
nor U15262 (N_15262,N_13529,N_12319);
nor U15263 (N_15263,N_12264,N_13985);
nor U15264 (N_15264,N_13550,N_13549);
and U15265 (N_15265,N_12224,N_12260);
nor U15266 (N_15266,N_13565,N_13628);
xor U15267 (N_15267,N_12108,N_12716);
and U15268 (N_15268,N_13736,N_13365);
and U15269 (N_15269,N_12862,N_13912);
or U15270 (N_15270,N_12937,N_12590);
nand U15271 (N_15271,N_12896,N_13392);
nand U15272 (N_15272,N_13898,N_12123);
or U15273 (N_15273,N_12614,N_13458);
or U15274 (N_15274,N_12848,N_12480);
or U15275 (N_15275,N_13851,N_12391);
and U15276 (N_15276,N_12514,N_12852);
xor U15277 (N_15277,N_13932,N_13232);
and U15278 (N_15278,N_13748,N_13328);
or U15279 (N_15279,N_13299,N_13785);
nor U15280 (N_15280,N_13158,N_12123);
and U15281 (N_15281,N_13866,N_13710);
nand U15282 (N_15282,N_12285,N_12899);
and U15283 (N_15283,N_12727,N_12968);
nand U15284 (N_15284,N_13591,N_13562);
and U15285 (N_15285,N_12885,N_12782);
or U15286 (N_15286,N_13949,N_12600);
nand U15287 (N_15287,N_12347,N_12083);
nand U15288 (N_15288,N_13526,N_13756);
and U15289 (N_15289,N_13974,N_12182);
nor U15290 (N_15290,N_12062,N_12893);
and U15291 (N_15291,N_12874,N_13488);
or U15292 (N_15292,N_12892,N_12171);
nor U15293 (N_15293,N_12680,N_13676);
xnor U15294 (N_15294,N_13889,N_13130);
or U15295 (N_15295,N_12261,N_12388);
or U15296 (N_15296,N_13146,N_12005);
xor U15297 (N_15297,N_13331,N_13122);
xnor U15298 (N_15298,N_13412,N_12410);
nand U15299 (N_15299,N_13100,N_12174);
nor U15300 (N_15300,N_12355,N_13698);
xor U15301 (N_15301,N_13970,N_12708);
nor U15302 (N_15302,N_12127,N_13010);
nand U15303 (N_15303,N_12571,N_13872);
nor U15304 (N_15304,N_12473,N_12806);
nor U15305 (N_15305,N_12304,N_13071);
nor U15306 (N_15306,N_13923,N_13856);
nor U15307 (N_15307,N_12218,N_13919);
xnor U15308 (N_15308,N_12983,N_13248);
nand U15309 (N_15309,N_12107,N_13192);
nor U15310 (N_15310,N_13676,N_12378);
and U15311 (N_15311,N_12031,N_12625);
and U15312 (N_15312,N_12953,N_12304);
nand U15313 (N_15313,N_12004,N_12319);
nand U15314 (N_15314,N_12220,N_12779);
and U15315 (N_15315,N_13039,N_12507);
or U15316 (N_15316,N_13094,N_12445);
or U15317 (N_15317,N_12258,N_12123);
nor U15318 (N_15318,N_13943,N_13850);
nor U15319 (N_15319,N_12536,N_13900);
nor U15320 (N_15320,N_13917,N_12203);
nor U15321 (N_15321,N_13343,N_12881);
and U15322 (N_15322,N_13592,N_13594);
nand U15323 (N_15323,N_12936,N_13821);
xnor U15324 (N_15324,N_12240,N_12415);
nor U15325 (N_15325,N_12304,N_12862);
nor U15326 (N_15326,N_12139,N_13230);
nand U15327 (N_15327,N_12165,N_12778);
xor U15328 (N_15328,N_12603,N_12009);
and U15329 (N_15329,N_13729,N_13714);
or U15330 (N_15330,N_12400,N_13853);
nor U15331 (N_15331,N_13327,N_12717);
xor U15332 (N_15332,N_13276,N_13476);
nor U15333 (N_15333,N_12496,N_13368);
xor U15334 (N_15334,N_13236,N_13271);
nand U15335 (N_15335,N_12174,N_12514);
nand U15336 (N_15336,N_13146,N_12951);
and U15337 (N_15337,N_13809,N_13432);
xnor U15338 (N_15338,N_13878,N_13439);
nand U15339 (N_15339,N_13039,N_13018);
and U15340 (N_15340,N_12336,N_12399);
xnor U15341 (N_15341,N_12261,N_13048);
nor U15342 (N_15342,N_12138,N_12788);
nor U15343 (N_15343,N_13565,N_12126);
nand U15344 (N_15344,N_13541,N_12059);
nor U15345 (N_15345,N_12061,N_13848);
and U15346 (N_15346,N_12258,N_13338);
nand U15347 (N_15347,N_12629,N_13009);
xnor U15348 (N_15348,N_12517,N_13704);
nor U15349 (N_15349,N_13477,N_12884);
and U15350 (N_15350,N_13222,N_12292);
or U15351 (N_15351,N_13894,N_12435);
and U15352 (N_15352,N_13180,N_12434);
or U15353 (N_15353,N_13662,N_12232);
or U15354 (N_15354,N_12533,N_12014);
or U15355 (N_15355,N_12138,N_13445);
and U15356 (N_15356,N_13762,N_12990);
nor U15357 (N_15357,N_13160,N_12682);
and U15358 (N_15358,N_13228,N_13143);
or U15359 (N_15359,N_13853,N_12230);
or U15360 (N_15360,N_12478,N_12995);
or U15361 (N_15361,N_12357,N_13539);
nand U15362 (N_15362,N_12035,N_12758);
or U15363 (N_15363,N_13220,N_12843);
and U15364 (N_15364,N_13765,N_13850);
and U15365 (N_15365,N_13536,N_13812);
or U15366 (N_15366,N_13016,N_12588);
nor U15367 (N_15367,N_13317,N_13915);
nand U15368 (N_15368,N_13757,N_13243);
and U15369 (N_15369,N_13605,N_12624);
or U15370 (N_15370,N_13975,N_12474);
and U15371 (N_15371,N_13545,N_13588);
nand U15372 (N_15372,N_13243,N_13911);
and U15373 (N_15373,N_12903,N_13809);
nand U15374 (N_15374,N_13104,N_13026);
or U15375 (N_15375,N_12581,N_13664);
and U15376 (N_15376,N_13559,N_12106);
nand U15377 (N_15377,N_12346,N_12289);
xor U15378 (N_15378,N_13935,N_13334);
nand U15379 (N_15379,N_12455,N_12745);
xor U15380 (N_15380,N_13982,N_13147);
nand U15381 (N_15381,N_12490,N_12847);
nor U15382 (N_15382,N_13595,N_13807);
xnor U15383 (N_15383,N_13726,N_13189);
nor U15384 (N_15384,N_13456,N_13038);
nand U15385 (N_15385,N_13551,N_12473);
xor U15386 (N_15386,N_13624,N_12264);
nor U15387 (N_15387,N_12627,N_13662);
nor U15388 (N_15388,N_13303,N_13567);
or U15389 (N_15389,N_12193,N_13644);
nor U15390 (N_15390,N_12640,N_13083);
xnor U15391 (N_15391,N_12200,N_13070);
xnor U15392 (N_15392,N_13943,N_13077);
nand U15393 (N_15393,N_12141,N_13001);
xnor U15394 (N_15394,N_12877,N_12516);
xor U15395 (N_15395,N_13020,N_12396);
or U15396 (N_15396,N_12941,N_13663);
or U15397 (N_15397,N_13998,N_13604);
xnor U15398 (N_15398,N_13332,N_12835);
nand U15399 (N_15399,N_12233,N_13862);
or U15400 (N_15400,N_12339,N_12718);
nand U15401 (N_15401,N_12855,N_12865);
nor U15402 (N_15402,N_12476,N_13552);
or U15403 (N_15403,N_12879,N_13714);
nand U15404 (N_15404,N_12372,N_13368);
and U15405 (N_15405,N_12704,N_12941);
nand U15406 (N_15406,N_13481,N_13819);
or U15407 (N_15407,N_12048,N_12642);
or U15408 (N_15408,N_12948,N_12156);
and U15409 (N_15409,N_13175,N_12433);
xnor U15410 (N_15410,N_12178,N_12385);
nor U15411 (N_15411,N_13103,N_12173);
nand U15412 (N_15412,N_13837,N_13067);
or U15413 (N_15413,N_13698,N_12901);
or U15414 (N_15414,N_12524,N_13760);
or U15415 (N_15415,N_12534,N_13758);
or U15416 (N_15416,N_12086,N_12807);
or U15417 (N_15417,N_13838,N_12049);
xnor U15418 (N_15418,N_13511,N_13205);
and U15419 (N_15419,N_12121,N_12218);
nor U15420 (N_15420,N_13668,N_13745);
and U15421 (N_15421,N_12294,N_12497);
or U15422 (N_15422,N_13253,N_13782);
nand U15423 (N_15423,N_12233,N_13939);
nand U15424 (N_15424,N_13744,N_12195);
nor U15425 (N_15425,N_13032,N_12317);
xor U15426 (N_15426,N_13559,N_12185);
and U15427 (N_15427,N_12179,N_13392);
or U15428 (N_15428,N_13584,N_13761);
nor U15429 (N_15429,N_13231,N_12890);
or U15430 (N_15430,N_12765,N_13096);
nor U15431 (N_15431,N_13503,N_12082);
xor U15432 (N_15432,N_13487,N_13723);
and U15433 (N_15433,N_12751,N_13249);
nor U15434 (N_15434,N_12971,N_12075);
nor U15435 (N_15435,N_13427,N_12752);
or U15436 (N_15436,N_13464,N_12515);
xnor U15437 (N_15437,N_13728,N_13811);
or U15438 (N_15438,N_13023,N_13045);
or U15439 (N_15439,N_12659,N_13865);
xor U15440 (N_15440,N_12478,N_12262);
nor U15441 (N_15441,N_12665,N_12458);
xnor U15442 (N_15442,N_13734,N_12146);
nor U15443 (N_15443,N_12199,N_12528);
xnor U15444 (N_15444,N_13079,N_13993);
xor U15445 (N_15445,N_12093,N_13770);
nand U15446 (N_15446,N_13900,N_12067);
and U15447 (N_15447,N_12760,N_12246);
xnor U15448 (N_15448,N_13840,N_13411);
nor U15449 (N_15449,N_12172,N_12470);
nand U15450 (N_15450,N_12161,N_12854);
nand U15451 (N_15451,N_13191,N_12748);
nor U15452 (N_15452,N_13848,N_12142);
and U15453 (N_15453,N_12092,N_13682);
and U15454 (N_15454,N_12169,N_12254);
or U15455 (N_15455,N_13858,N_13736);
nand U15456 (N_15456,N_13040,N_12130);
nand U15457 (N_15457,N_12326,N_12928);
xor U15458 (N_15458,N_12021,N_13386);
or U15459 (N_15459,N_12626,N_12088);
and U15460 (N_15460,N_12321,N_12628);
nor U15461 (N_15461,N_12190,N_12706);
or U15462 (N_15462,N_12998,N_13444);
and U15463 (N_15463,N_13704,N_13972);
or U15464 (N_15464,N_12855,N_13476);
or U15465 (N_15465,N_13500,N_12322);
xor U15466 (N_15466,N_13366,N_12759);
or U15467 (N_15467,N_12103,N_12560);
nand U15468 (N_15468,N_13648,N_12162);
nor U15469 (N_15469,N_13031,N_13745);
nor U15470 (N_15470,N_13703,N_13751);
nor U15471 (N_15471,N_12790,N_12900);
nor U15472 (N_15472,N_13905,N_13239);
or U15473 (N_15473,N_13515,N_12972);
and U15474 (N_15474,N_12678,N_13924);
nand U15475 (N_15475,N_12922,N_13304);
nand U15476 (N_15476,N_12964,N_13492);
xnor U15477 (N_15477,N_13357,N_12607);
xnor U15478 (N_15478,N_13659,N_12668);
nor U15479 (N_15479,N_12662,N_12296);
nand U15480 (N_15480,N_13373,N_13519);
nand U15481 (N_15481,N_13719,N_13616);
nor U15482 (N_15482,N_13498,N_13668);
nor U15483 (N_15483,N_12572,N_13160);
xnor U15484 (N_15484,N_13392,N_13054);
nor U15485 (N_15485,N_12242,N_13326);
and U15486 (N_15486,N_13575,N_12793);
xor U15487 (N_15487,N_12302,N_12143);
nand U15488 (N_15488,N_12946,N_12817);
xnor U15489 (N_15489,N_13073,N_12179);
xnor U15490 (N_15490,N_12454,N_12140);
or U15491 (N_15491,N_12605,N_13341);
and U15492 (N_15492,N_13626,N_12327);
or U15493 (N_15493,N_13740,N_12893);
or U15494 (N_15494,N_12536,N_13845);
and U15495 (N_15495,N_12633,N_13757);
or U15496 (N_15496,N_12013,N_12531);
nand U15497 (N_15497,N_13163,N_12341);
xnor U15498 (N_15498,N_12242,N_13693);
and U15499 (N_15499,N_12880,N_12153);
nor U15500 (N_15500,N_12589,N_13046);
nand U15501 (N_15501,N_13389,N_12151);
nand U15502 (N_15502,N_12058,N_13723);
nand U15503 (N_15503,N_13656,N_12204);
xor U15504 (N_15504,N_13208,N_12432);
or U15505 (N_15505,N_12582,N_13927);
and U15506 (N_15506,N_13606,N_13498);
xor U15507 (N_15507,N_13180,N_13423);
or U15508 (N_15508,N_13911,N_13880);
nor U15509 (N_15509,N_13665,N_12035);
and U15510 (N_15510,N_13033,N_13275);
or U15511 (N_15511,N_13267,N_13692);
xnor U15512 (N_15512,N_13610,N_13715);
nor U15513 (N_15513,N_12218,N_12558);
and U15514 (N_15514,N_13066,N_13992);
nor U15515 (N_15515,N_13745,N_12636);
or U15516 (N_15516,N_12501,N_12248);
nor U15517 (N_15517,N_13654,N_13403);
nand U15518 (N_15518,N_13045,N_12570);
and U15519 (N_15519,N_12893,N_13751);
nor U15520 (N_15520,N_12547,N_13676);
or U15521 (N_15521,N_12246,N_13351);
nand U15522 (N_15522,N_12267,N_13675);
nand U15523 (N_15523,N_12695,N_12987);
nor U15524 (N_15524,N_13144,N_13474);
xor U15525 (N_15525,N_13722,N_13372);
xor U15526 (N_15526,N_13347,N_12927);
nor U15527 (N_15527,N_13310,N_13348);
and U15528 (N_15528,N_13619,N_12079);
nor U15529 (N_15529,N_13863,N_12933);
nor U15530 (N_15530,N_13397,N_12962);
xor U15531 (N_15531,N_12713,N_12561);
nor U15532 (N_15532,N_12644,N_12609);
or U15533 (N_15533,N_12754,N_13149);
and U15534 (N_15534,N_12617,N_12660);
and U15535 (N_15535,N_12826,N_12784);
nor U15536 (N_15536,N_12076,N_12267);
nor U15537 (N_15537,N_12887,N_12073);
nand U15538 (N_15538,N_12375,N_13008);
or U15539 (N_15539,N_12452,N_12698);
nor U15540 (N_15540,N_12661,N_12423);
or U15541 (N_15541,N_12901,N_13059);
xor U15542 (N_15542,N_13642,N_13539);
nor U15543 (N_15543,N_12283,N_13538);
xnor U15544 (N_15544,N_13041,N_13509);
xnor U15545 (N_15545,N_12339,N_13678);
nor U15546 (N_15546,N_12520,N_13288);
nand U15547 (N_15547,N_12954,N_13299);
nor U15548 (N_15548,N_13839,N_12488);
and U15549 (N_15549,N_13407,N_13482);
nand U15550 (N_15550,N_13396,N_12647);
and U15551 (N_15551,N_12478,N_13124);
and U15552 (N_15552,N_12526,N_13882);
xor U15553 (N_15553,N_13348,N_13401);
xnor U15554 (N_15554,N_13143,N_12533);
nand U15555 (N_15555,N_13552,N_12315);
nand U15556 (N_15556,N_12937,N_12192);
nor U15557 (N_15557,N_13945,N_12690);
or U15558 (N_15558,N_12046,N_13726);
nand U15559 (N_15559,N_12196,N_12779);
nor U15560 (N_15560,N_12975,N_13335);
xor U15561 (N_15561,N_12747,N_12530);
or U15562 (N_15562,N_12926,N_12970);
and U15563 (N_15563,N_12449,N_12830);
nand U15564 (N_15564,N_12028,N_13217);
and U15565 (N_15565,N_12640,N_13874);
and U15566 (N_15566,N_13761,N_12954);
and U15567 (N_15567,N_13708,N_13007);
xnor U15568 (N_15568,N_13701,N_13672);
xnor U15569 (N_15569,N_13680,N_13729);
nand U15570 (N_15570,N_12145,N_12429);
xor U15571 (N_15571,N_12503,N_13864);
or U15572 (N_15572,N_13105,N_12072);
nand U15573 (N_15573,N_13073,N_13442);
nor U15574 (N_15574,N_13819,N_13242);
or U15575 (N_15575,N_13243,N_13668);
xor U15576 (N_15576,N_13888,N_13290);
nor U15577 (N_15577,N_13300,N_13866);
xnor U15578 (N_15578,N_12205,N_13882);
nand U15579 (N_15579,N_13241,N_12765);
nand U15580 (N_15580,N_13233,N_12702);
nand U15581 (N_15581,N_12495,N_13998);
or U15582 (N_15582,N_13286,N_13039);
or U15583 (N_15583,N_12264,N_13117);
nor U15584 (N_15584,N_12014,N_12147);
or U15585 (N_15585,N_12050,N_12595);
and U15586 (N_15586,N_12932,N_13594);
xor U15587 (N_15587,N_13438,N_12875);
nand U15588 (N_15588,N_13107,N_13985);
and U15589 (N_15589,N_13348,N_13426);
xor U15590 (N_15590,N_13986,N_12363);
and U15591 (N_15591,N_12154,N_13034);
nand U15592 (N_15592,N_13109,N_13492);
or U15593 (N_15593,N_12067,N_13870);
nand U15594 (N_15594,N_12960,N_13876);
xnor U15595 (N_15595,N_12488,N_12494);
nor U15596 (N_15596,N_13043,N_13091);
xor U15597 (N_15597,N_13489,N_13436);
nor U15598 (N_15598,N_12875,N_12156);
nand U15599 (N_15599,N_13341,N_12936);
nand U15600 (N_15600,N_13091,N_13030);
nand U15601 (N_15601,N_12074,N_13449);
and U15602 (N_15602,N_12151,N_13844);
nor U15603 (N_15603,N_13514,N_13436);
and U15604 (N_15604,N_12916,N_12513);
nand U15605 (N_15605,N_13952,N_13136);
or U15606 (N_15606,N_12482,N_12658);
xor U15607 (N_15607,N_13445,N_13364);
or U15608 (N_15608,N_12551,N_12428);
or U15609 (N_15609,N_12709,N_12086);
nor U15610 (N_15610,N_13003,N_12709);
xor U15611 (N_15611,N_13585,N_12065);
or U15612 (N_15612,N_12118,N_13035);
nand U15613 (N_15613,N_12884,N_13556);
nor U15614 (N_15614,N_12038,N_13333);
xnor U15615 (N_15615,N_13997,N_12990);
or U15616 (N_15616,N_12318,N_12718);
nand U15617 (N_15617,N_13109,N_13230);
xor U15618 (N_15618,N_12184,N_13557);
xor U15619 (N_15619,N_12494,N_13132);
and U15620 (N_15620,N_12978,N_13404);
nor U15621 (N_15621,N_13039,N_12591);
xor U15622 (N_15622,N_13397,N_12098);
and U15623 (N_15623,N_12208,N_13880);
and U15624 (N_15624,N_12650,N_12694);
nor U15625 (N_15625,N_13181,N_13800);
and U15626 (N_15626,N_12090,N_13961);
nand U15627 (N_15627,N_13863,N_13602);
xor U15628 (N_15628,N_12925,N_12418);
and U15629 (N_15629,N_13202,N_13179);
nor U15630 (N_15630,N_12823,N_13537);
and U15631 (N_15631,N_13472,N_12008);
and U15632 (N_15632,N_13872,N_12759);
nand U15633 (N_15633,N_13206,N_12442);
xnor U15634 (N_15634,N_13458,N_13363);
nand U15635 (N_15635,N_12646,N_12828);
or U15636 (N_15636,N_12923,N_13977);
and U15637 (N_15637,N_13059,N_12504);
or U15638 (N_15638,N_12805,N_13599);
nor U15639 (N_15639,N_12042,N_13364);
nand U15640 (N_15640,N_13760,N_13174);
or U15641 (N_15641,N_12452,N_13933);
xor U15642 (N_15642,N_12768,N_12784);
nand U15643 (N_15643,N_13436,N_13870);
xor U15644 (N_15644,N_13736,N_12869);
or U15645 (N_15645,N_13393,N_13117);
nor U15646 (N_15646,N_13571,N_13595);
or U15647 (N_15647,N_13139,N_12292);
or U15648 (N_15648,N_13297,N_12139);
or U15649 (N_15649,N_13109,N_13584);
xnor U15650 (N_15650,N_13907,N_12270);
nand U15651 (N_15651,N_12482,N_13701);
xor U15652 (N_15652,N_13180,N_12466);
and U15653 (N_15653,N_12694,N_12699);
xor U15654 (N_15654,N_13253,N_12135);
or U15655 (N_15655,N_12188,N_12683);
xor U15656 (N_15656,N_12655,N_13968);
and U15657 (N_15657,N_13724,N_13880);
and U15658 (N_15658,N_12699,N_13741);
and U15659 (N_15659,N_12937,N_13286);
or U15660 (N_15660,N_13650,N_12217);
or U15661 (N_15661,N_13747,N_12388);
xor U15662 (N_15662,N_12964,N_12739);
or U15663 (N_15663,N_12584,N_13342);
nand U15664 (N_15664,N_13312,N_13003);
and U15665 (N_15665,N_12231,N_13982);
or U15666 (N_15666,N_13904,N_12561);
xnor U15667 (N_15667,N_13664,N_12544);
nor U15668 (N_15668,N_13610,N_13103);
and U15669 (N_15669,N_12085,N_13559);
xnor U15670 (N_15670,N_12530,N_12035);
nand U15671 (N_15671,N_12980,N_12215);
nand U15672 (N_15672,N_12739,N_13168);
nor U15673 (N_15673,N_12025,N_13543);
nand U15674 (N_15674,N_12748,N_13541);
nor U15675 (N_15675,N_13435,N_13142);
nand U15676 (N_15676,N_13303,N_13846);
and U15677 (N_15677,N_12983,N_12542);
or U15678 (N_15678,N_13885,N_12684);
and U15679 (N_15679,N_13117,N_13617);
and U15680 (N_15680,N_12637,N_13140);
or U15681 (N_15681,N_12628,N_12934);
nand U15682 (N_15682,N_13854,N_12582);
xnor U15683 (N_15683,N_12015,N_13511);
nand U15684 (N_15684,N_13351,N_12871);
xnor U15685 (N_15685,N_13140,N_12837);
or U15686 (N_15686,N_12956,N_13154);
nand U15687 (N_15687,N_12164,N_13933);
xor U15688 (N_15688,N_13795,N_12969);
and U15689 (N_15689,N_12171,N_12103);
xnor U15690 (N_15690,N_12682,N_13277);
nor U15691 (N_15691,N_13334,N_13291);
nor U15692 (N_15692,N_12738,N_13694);
or U15693 (N_15693,N_12401,N_12211);
or U15694 (N_15694,N_12631,N_13055);
xor U15695 (N_15695,N_12002,N_13924);
nor U15696 (N_15696,N_13508,N_13596);
nand U15697 (N_15697,N_12509,N_12041);
nand U15698 (N_15698,N_12598,N_12804);
and U15699 (N_15699,N_12333,N_13375);
or U15700 (N_15700,N_13599,N_12118);
xnor U15701 (N_15701,N_13148,N_12068);
xor U15702 (N_15702,N_12902,N_12409);
xor U15703 (N_15703,N_13124,N_12574);
nand U15704 (N_15704,N_12482,N_12237);
and U15705 (N_15705,N_12468,N_12325);
or U15706 (N_15706,N_12790,N_12100);
nor U15707 (N_15707,N_13545,N_12296);
nor U15708 (N_15708,N_13685,N_13299);
or U15709 (N_15709,N_12174,N_12345);
or U15710 (N_15710,N_12217,N_13319);
nor U15711 (N_15711,N_13596,N_12710);
nand U15712 (N_15712,N_13520,N_13845);
xor U15713 (N_15713,N_13594,N_13149);
nand U15714 (N_15714,N_12304,N_12880);
nor U15715 (N_15715,N_12107,N_13191);
nor U15716 (N_15716,N_13407,N_13188);
nor U15717 (N_15717,N_12482,N_13310);
nor U15718 (N_15718,N_12630,N_12293);
nor U15719 (N_15719,N_13940,N_12640);
and U15720 (N_15720,N_12422,N_13466);
xnor U15721 (N_15721,N_12494,N_13482);
or U15722 (N_15722,N_12710,N_13351);
nand U15723 (N_15723,N_13889,N_12942);
nor U15724 (N_15724,N_12223,N_13864);
and U15725 (N_15725,N_12581,N_13792);
nand U15726 (N_15726,N_12766,N_12592);
or U15727 (N_15727,N_12338,N_12832);
and U15728 (N_15728,N_13808,N_12837);
or U15729 (N_15729,N_13947,N_12144);
and U15730 (N_15730,N_13111,N_12640);
nand U15731 (N_15731,N_12296,N_12032);
nand U15732 (N_15732,N_12431,N_13393);
nor U15733 (N_15733,N_13517,N_13396);
or U15734 (N_15734,N_13178,N_13796);
nor U15735 (N_15735,N_12595,N_13137);
nor U15736 (N_15736,N_12674,N_12914);
or U15737 (N_15737,N_13482,N_12188);
xor U15738 (N_15738,N_12253,N_13018);
xnor U15739 (N_15739,N_13179,N_12449);
nor U15740 (N_15740,N_13359,N_13724);
nand U15741 (N_15741,N_13925,N_12358);
nand U15742 (N_15742,N_13638,N_12279);
or U15743 (N_15743,N_13225,N_12198);
and U15744 (N_15744,N_12048,N_13511);
nand U15745 (N_15745,N_13336,N_12873);
xor U15746 (N_15746,N_12356,N_12593);
and U15747 (N_15747,N_13643,N_13901);
xor U15748 (N_15748,N_13528,N_13693);
and U15749 (N_15749,N_12395,N_13680);
nand U15750 (N_15750,N_12555,N_13110);
nor U15751 (N_15751,N_12586,N_13344);
nand U15752 (N_15752,N_13619,N_12654);
and U15753 (N_15753,N_13666,N_12911);
nand U15754 (N_15754,N_12585,N_12332);
or U15755 (N_15755,N_12318,N_13216);
and U15756 (N_15756,N_12610,N_12883);
nand U15757 (N_15757,N_13549,N_12052);
nand U15758 (N_15758,N_12431,N_13157);
or U15759 (N_15759,N_12436,N_13203);
or U15760 (N_15760,N_12348,N_12871);
or U15761 (N_15761,N_12549,N_12146);
nor U15762 (N_15762,N_12113,N_12155);
nor U15763 (N_15763,N_12783,N_13672);
and U15764 (N_15764,N_13298,N_12814);
nor U15765 (N_15765,N_13007,N_13406);
and U15766 (N_15766,N_12998,N_12087);
xnor U15767 (N_15767,N_12446,N_13819);
or U15768 (N_15768,N_13478,N_12281);
and U15769 (N_15769,N_13345,N_13529);
xor U15770 (N_15770,N_12515,N_12600);
or U15771 (N_15771,N_13775,N_12092);
nand U15772 (N_15772,N_12461,N_13653);
xnor U15773 (N_15773,N_12150,N_13604);
nand U15774 (N_15774,N_12616,N_12004);
or U15775 (N_15775,N_12574,N_12531);
and U15776 (N_15776,N_13549,N_12964);
xor U15777 (N_15777,N_12361,N_13442);
nor U15778 (N_15778,N_12499,N_13854);
and U15779 (N_15779,N_13071,N_12134);
nor U15780 (N_15780,N_13885,N_12522);
nor U15781 (N_15781,N_13571,N_12190);
and U15782 (N_15782,N_12740,N_13254);
xnor U15783 (N_15783,N_13232,N_12467);
and U15784 (N_15784,N_12186,N_12710);
xnor U15785 (N_15785,N_13647,N_12373);
and U15786 (N_15786,N_13758,N_12257);
and U15787 (N_15787,N_12710,N_13486);
and U15788 (N_15788,N_12904,N_12266);
xor U15789 (N_15789,N_12411,N_12284);
and U15790 (N_15790,N_12268,N_13935);
nor U15791 (N_15791,N_13584,N_13256);
or U15792 (N_15792,N_13482,N_12342);
nor U15793 (N_15793,N_12394,N_12053);
and U15794 (N_15794,N_13687,N_12700);
xnor U15795 (N_15795,N_13300,N_12419);
xnor U15796 (N_15796,N_12853,N_13006);
and U15797 (N_15797,N_12449,N_12795);
or U15798 (N_15798,N_12910,N_13729);
xor U15799 (N_15799,N_13004,N_12962);
nand U15800 (N_15800,N_13067,N_12657);
nand U15801 (N_15801,N_12636,N_13249);
or U15802 (N_15802,N_12099,N_13785);
and U15803 (N_15803,N_12923,N_13174);
and U15804 (N_15804,N_13000,N_13463);
xnor U15805 (N_15805,N_12390,N_13894);
xor U15806 (N_15806,N_12402,N_13744);
and U15807 (N_15807,N_12064,N_12817);
and U15808 (N_15808,N_13018,N_12885);
or U15809 (N_15809,N_12977,N_12771);
nor U15810 (N_15810,N_12777,N_13293);
or U15811 (N_15811,N_12024,N_13025);
or U15812 (N_15812,N_12161,N_13635);
xnor U15813 (N_15813,N_13037,N_12238);
and U15814 (N_15814,N_13780,N_12694);
or U15815 (N_15815,N_13155,N_13453);
and U15816 (N_15816,N_12657,N_13745);
xnor U15817 (N_15817,N_13388,N_12621);
and U15818 (N_15818,N_13976,N_12312);
xor U15819 (N_15819,N_13511,N_13284);
xnor U15820 (N_15820,N_13425,N_12823);
nor U15821 (N_15821,N_13766,N_13032);
nand U15822 (N_15822,N_12141,N_13861);
nor U15823 (N_15823,N_12354,N_12869);
or U15824 (N_15824,N_12075,N_13730);
and U15825 (N_15825,N_12039,N_13091);
xor U15826 (N_15826,N_13617,N_13116);
or U15827 (N_15827,N_12569,N_13107);
nor U15828 (N_15828,N_12808,N_13781);
or U15829 (N_15829,N_12121,N_12860);
or U15830 (N_15830,N_12891,N_13301);
and U15831 (N_15831,N_13023,N_12868);
nand U15832 (N_15832,N_13341,N_13956);
and U15833 (N_15833,N_12494,N_13807);
nand U15834 (N_15834,N_12308,N_12535);
and U15835 (N_15835,N_13068,N_12918);
and U15836 (N_15836,N_13814,N_12233);
or U15837 (N_15837,N_13339,N_13559);
nor U15838 (N_15838,N_12243,N_13600);
xor U15839 (N_15839,N_13479,N_13462);
xnor U15840 (N_15840,N_12531,N_12840);
nor U15841 (N_15841,N_12839,N_12021);
and U15842 (N_15842,N_12477,N_12383);
and U15843 (N_15843,N_12938,N_12284);
or U15844 (N_15844,N_13894,N_13820);
or U15845 (N_15845,N_13144,N_12652);
xor U15846 (N_15846,N_13114,N_13767);
xor U15847 (N_15847,N_12178,N_12760);
or U15848 (N_15848,N_13045,N_13157);
or U15849 (N_15849,N_13451,N_12792);
or U15850 (N_15850,N_12917,N_13307);
xnor U15851 (N_15851,N_13182,N_12297);
or U15852 (N_15852,N_13940,N_12351);
and U15853 (N_15853,N_12511,N_12206);
or U15854 (N_15854,N_13296,N_13808);
and U15855 (N_15855,N_13036,N_13310);
or U15856 (N_15856,N_12283,N_13976);
or U15857 (N_15857,N_13652,N_12956);
or U15858 (N_15858,N_13210,N_12882);
nand U15859 (N_15859,N_12436,N_12888);
xor U15860 (N_15860,N_13559,N_12422);
and U15861 (N_15861,N_12337,N_12962);
nor U15862 (N_15862,N_12439,N_13845);
nor U15863 (N_15863,N_13030,N_13767);
and U15864 (N_15864,N_13312,N_12300);
or U15865 (N_15865,N_12861,N_12670);
nor U15866 (N_15866,N_12640,N_12146);
xor U15867 (N_15867,N_12951,N_12062);
and U15868 (N_15868,N_13970,N_13498);
or U15869 (N_15869,N_13473,N_12755);
or U15870 (N_15870,N_12101,N_13901);
and U15871 (N_15871,N_13797,N_12666);
nand U15872 (N_15872,N_12655,N_13947);
xor U15873 (N_15873,N_12891,N_13614);
or U15874 (N_15874,N_12545,N_12380);
nor U15875 (N_15875,N_12067,N_13297);
nand U15876 (N_15876,N_12501,N_12851);
and U15877 (N_15877,N_12707,N_12745);
and U15878 (N_15878,N_13018,N_13902);
nor U15879 (N_15879,N_13966,N_12436);
or U15880 (N_15880,N_13128,N_13794);
nand U15881 (N_15881,N_13778,N_13636);
nor U15882 (N_15882,N_13659,N_13670);
xor U15883 (N_15883,N_12897,N_12573);
nand U15884 (N_15884,N_12326,N_12514);
and U15885 (N_15885,N_13322,N_13291);
nor U15886 (N_15886,N_12947,N_13424);
and U15887 (N_15887,N_13716,N_13357);
and U15888 (N_15888,N_13628,N_12266);
xnor U15889 (N_15889,N_12917,N_12578);
or U15890 (N_15890,N_13858,N_12181);
nor U15891 (N_15891,N_13851,N_12117);
xnor U15892 (N_15892,N_13874,N_12006);
and U15893 (N_15893,N_13147,N_12935);
or U15894 (N_15894,N_12217,N_13452);
or U15895 (N_15895,N_12455,N_13208);
and U15896 (N_15896,N_13302,N_12861);
or U15897 (N_15897,N_13395,N_13574);
xnor U15898 (N_15898,N_12499,N_12445);
xnor U15899 (N_15899,N_12105,N_13212);
nor U15900 (N_15900,N_13460,N_13918);
xor U15901 (N_15901,N_13492,N_13037);
and U15902 (N_15902,N_12663,N_13760);
nor U15903 (N_15903,N_12755,N_13840);
or U15904 (N_15904,N_12113,N_13345);
and U15905 (N_15905,N_12823,N_12501);
or U15906 (N_15906,N_12062,N_12081);
and U15907 (N_15907,N_12385,N_12205);
or U15908 (N_15908,N_12276,N_13325);
xor U15909 (N_15909,N_13661,N_12702);
xnor U15910 (N_15910,N_12701,N_13536);
and U15911 (N_15911,N_13903,N_12155);
nand U15912 (N_15912,N_12678,N_12103);
nand U15913 (N_15913,N_13926,N_12901);
and U15914 (N_15914,N_13293,N_13487);
nand U15915 (N_15915,N_13441,N_12693);
nor U15916 (N_15916,N_12685,N_12583);
nand U15917 (N_15917,N_13858,N_12458);
and U15918 (N_15918,N_12299,N_12348);
nor U15919 (N_15919,N_13351,N_12396);
or U15920 (N_15920,N_13745,N_12486);
xor U15921 (N_15921,N_13127,N_12989);
xnor U15922 (N_15922,N_13916,N_13152);
and U15923 (N_15923,N_13945,N_12037);
and U15924 (N_15924,N_12128,N_13857);
nand U15925 (N_15925,N_13464,N_13733);
nor U15926 (N_15926,N_12567,N_12675);
nor U15927 (N_15927,N_12761,N_13388);
or U15928 (N_15928,N_13900,N_13448);
nand U15929 (N_15929,N_13969,N_12277);
and U15930 (N_15930,N_12800,N_13129);
or U15931 (N_15931,N_13013,N_13294);
nor U15932 (N_15932,N_12677,N_12640);
nand U15933 (N_15933,N_13866,N_12630);
and U15934 (N_15934,N_13847,N_13749);
or U15935 (N_15935,N_12883,N_12557);
nor U15936 (N_15936,N_13163,N_12909);
and U15937 (N_15937,N_13300,N_13069);
and U15938 (N_15938,N_12635,N_12492);
or U15939 (N_15939,N_13759,N_13044);
nand U15940 (N_15940,N_12369,N_13970);
nor U15941 (N_15941,N_12095,N_12922);
or U15942 (N_15942,N_12200,N_13700);
and U15943 (N_15943,N_12371,N_12915);
and U15944 (N_15944,N_13060,N_13155);
nand U15945 (N_15945,N_12657,N_13184);
and U15946 (N_15946,N_12337,N_12803);
nor U15947 (N_15947,N_13491,N_13404);
nand U15948 (N_15948,N_12051,N_12774);
nor U15949 (N_15949,N_13786,N_13180);
xor U15950 (N_15950,N_12204,N_12343);
nand U15951 (N_15951,N_13108,N_12056);
nor U15952 (N_15952,N_12294,N_13165);
xor U15953 (N_15953,N_13156,N_13287);
and U15954 (N_15954,N_13406,N_13893);
nor U15955 (N_15955,N_12755,N_13966);
nand U15956 (N_15956,N_12184,N_12251);
nand U15957 (N_15957,N_13552,N_12147);
or U15958 (N_15958,N_12665,N_13292);
or U15959 (N_15959,N_13108,N_13946);
xor U15960 (N_15960,N_13678,N_12999);
nor U15961 (N_15961,N_13778,N_12916);
and U15962 (N_15962,N_13799,N_12320);
or U15963 (N_15963,N_12662,N_12805);
xor U15964 (N_15964,N_12534,N_13902);
or U15965 (N_15965,N_12920,N_12935);
nand U15966 (N_15966,N_13803,N_12077);
nand U15967 (N_15967,N_13578,N_13165);
nor U15968 (N_15968,N_13177,N_12477);
and U15969 (N_15969,N_13486,N_13449);
and U15970 (N_15970,N_13638,N_13075);
or U15971 (N_15971,N_12542,N_12043);
or U15972 (N_15972,N_13053,N_13445);
or U15973 (N_15973,N_13437,N_13308);
nand U15974 (N_15974,N_12576,N_13714);
nand U15975 (N_15975,N_13061,N_12057);
nor U15976 (N_15976,N_12105,N_12612);
nand U15977 (N_15977,N_13909,N_12371);
nor U15978 (N_15978,N_13434,N_12343);
or U15979 (N_15979,N_13112,N_12322);
and U15980 (N_15980,N_13779,N_13161);
nor U15981 (N_15981,N_12368,N_13368);
or U15982 (N_15982,N_12495,N_12588);
and U15983 (N_15983,N_12800,N_13206);
nand U15984 (N_15984,N_12706,N_13964);
and U15985 (N_15985,N_12870,N_13386);
nor U15986 (N_15986,N_13213,N_12171);
nand U15987 (N_15987,N_12857,N_12557);
nand U15988 (N_15988,N_13369,N_13600);
xnor U15989 (N_15989,N_13960,N_12615);
or U15990 (N_15990,N_13975,N_12798);
or U15991 (N_15991,N_13787,N_13951);
xor U15992 (N_15992,N_13723,N_12954);
or U15993 (N_15993,N_12836,N_12569);
nor U15994 (N_15994,N_13808,N_12218);
and U15995 (N_15995,N_13893,N_12903);
xnor U15996 (N_15996,N_13195,N_12142);
or U15997 (N_15997,N_12306,N_12821);
or U15998 (N_15998,N_12554,N_12428);
or U15999 (N_15999,N_12251,N_12095);
nand U16000 (N_16000,N_14473,N_15608);
nand U16001 (N_16001,N_14648,N_14950);
xor U16002 (N_16002,N_15208,N_14792);
or U16003 (N_16003,N_14355,N_15124);
xnor U16004 (N_16004,N_14071,N_15479);
nor U16005 (N_16005,N_15559,N_15785);
nor U16006 (N_16006,N_14456,N_14921);
xor U16007 (N_16007,N_15537,N_15623);
and U16008 (N_16008,N_15950,N_14598);
xor U16009 (N_16009,N_15845,N_14870);
nor U16010 (N_16010,N_14748,N_15418);
or U16011 (N_16011,N_14934,N_14961);
or U16012 (N_16012,N_14133,N_14948);
nand U16013 (N_16013,N_14156,N_15987);
xor U16014 (N_16014,N_15597,N_15546);
and U16015 (N_16015,N_15240,N_15259);
nor U16016 (N_16016,N_15017,N_15340);
nor U16017 (N_16017,N_14005,N_14716);
and U16018 (N_16018,N_15134,N_14387);
or U16019 (N_16019,N_15793,N_15449);
xor U16020 (N_16020,N_14059,N_14567);
nor U16021 (N_16021,N_14054,N_15094);
nand U16022 (N_16022,N_15233,N_15994);
nor U16023 (N_16023,N_15056,N_14395);
nor U16024 (N_16024,N_15458,N_15344);
and U16025 (N_16025,N_14370,N_14615);
and U16026 (N_16026,N_14068,N_14541);
xor U16027 (N_16027,N_15780,N_15657);
nand U16028 (N_16028,N_14254,N_14721);
xor U16029 (N_16029,N_14487,N_14882);
and U16030 (N_16030,N_15752,N_14682);
and U16031 (N_16031,N_15505,N_15722);
xor U16032 (N_16032,N_14700,N_15542);
and U16033 (N_16033,N_15273,N_14907);
or U16034 (N_16034,N_14182,N_15452);
and U16035 (N_16035,N_15236,N_15164);
and U16036 (N_16036,N_14694,N_15003);
nand U16037 (N_16037,N_14877,N_15828);
and U16038 (N_16038,N_14462,N_14665);
and U16039 (N_16039,N_15797,N_14287);
and U16040 (N_16040,N_14045,N_14659);
and U16041 (N_16041,N_14526,N_14299);
and U16042 (N_16042,N_15408,N_15843);
nor U16043 (N_16043,N_14952,N_14637);
nand U16044 (N_16044,N_15839,N_15533);
nand U16045 (N_16045,N_14565,N_14266);
or U16046 (N_16046,N_14463,N_15866);
or U16047 (N_16047,N_14431,N_14233);
or U16048 (N_16048,N_14786,N_14649);
and U16049 (N_16049,N_14618,N_14026);
nor U16050 (N_16050,N_15063,N_15123);
and U16051 (N_16051,N_14129,N_15256);
nand U16052 (N_16052,N_14698,N_15510);
xor U16053 (N_16053,N_14739,N_14738);
nand U16054 (N_16054,N_14607,N_14813);
or U16055 (N_16055,N_15761,N_14664);
and U16056 (N_16056,N_14190,N_14602);
and U16057 (N_16057,N_15195,N_15963);
and U16058 (N_16058,N_14745,N_14707);
nor U16059 (N_16059,N_15379,N_14154);
xnor U16060 (N_16060,N_15411,N_14413);
and U16061 (N_16061,N_15946,N_14397);
nor U16062 (N_16062,N_14338,N_14589);
xnor U16063 (N_16063,N_15178,N_14094);
or U16064 (N_16064,N_15052,N_14434);
or U16065 (N_16065,N_15136,N_15663);
or U16066 (N_16066,N_14278,N_14440);
xnor U16067 (N_16067,N_15241,N_15137);
nand U16068 (N_16068,N_15291,N_14920);
and U16069 (N_16069,N_14157,N_14159);
nor U16070 (N_16070,N_14225,N_14232);
or U16071 (N_16071,N_15119,N_15333);
nand U16072 (N_16072,N_15262,N_15374);
or U16073 (N_16073,N_15093,N_14186);
and U16074 (N_16074,N_14075,N_15757);
nor U16075 (N_16075,N_15162,N_14111);
xor U16076 (N_16076,N_15177,N_15816);
nor U16077 (N_16077,N_15806,N_15368);
or U16078 (N_16078,N_14860,N_15530);
and U16079 (N_16079,N_14984,N_14571);
nand U16080 (N_16080,N_15257,N_14679);
and U16081 (N_16081,N_14353,N_15928);
nor U16082 (N_16082,N_15480,N_14422);
xor U16083 (N_16083,N_14687,N_14817);
nor U16084 (N_16084,N_15332,N_15749);
and U16085 (N_16085,N_15297,N_14863);
or U16086 (N_16086,N_15674,N_14873);
nor U16087 (N_16087,N_14505,N_15989);
nand U16088 (N_16088,N_15067,N_14942);
or U16089 (N_16089,N_14670,N_15967);
nor U16090 (N_16090,N_15005,N_14247);
or U16091 (N_16091,N_15978,N_14557);
and U16092 (N_16092,N_14742,N_14409);
nand U16093 (N_16093,N_15009,N_15016);
nor U16094 (N_16094,N_15279,N_15900);
nand U16095 (N_16095,N_14916,N_15500);
xor U16096 (N_16096,N_14173,N_14398);
nand U16097 (N_16097,N_14134,N_14788);
and U16098 (N_16098,N_14241,N_15156);
nor U16099 (N_16099,N_14854,N_14537);
and U16100 (N_16100,N_15531,N_15952);
nor U16101 (N_16101,N_15742,N_15201);
or U16102 (N_16102,N_15721,N_14931);
nand U16103 (N_16103,N_14550,N_15436);
or U16104 (N_16104,N_15842,N_14922);
nand U16105 (N_16105,N_14269,N_14548);
nor U16106 (N_16106,N_14688,N_15941);
xor U16107 (N_16107,N_14556,N_14221);
nand U16108 (N_16108,N_14477,N_14454);
and U16109 (N_16109,N_15281,N_15883);
nor U16110 (N_16110,N_15130,N_14695);
or U16111 (N_16111,N_15909,N_15562);
or U16112 (N_16112,N_15455,N_15388);
nand U16113 (N_16113,N_15927,N_15624);
nor U16114 (N_16114,N_14717,N_14521);
and U16115 (N_16115,N_15868,N_15580);
or U16116 (N_16116,N_15585,N_14351);
nor U16117 (N_16117,N_14193,N_14275);
nand U16118 (N_16118,N_14588,N_14118);
and U16119 (N_16119,N_14296,N_15497);
xnor U16120 (N_16120,N_14329,N_14298);
nand U16121 (N_16121,N_14144,N_15024);
and U16122 (N_16122,N_15518,N_14480);
nand U16123 (N_16123,N_14402,N_15278);
xor U16124 (N_16124,N_14706,N_15371);
nor U16125 (N_16125,N_14751,N_14723);
nor U16126 (N_16126,N_15653,N_15127);
or U16127 (N_16127,N_15028,N_15701);
and U16128 (N_16128,N_14478,N_15292);
nor U16129 (N_16129,N_14325,N_14972);
nand U16130 (N_16130,N_15917,N_14833);
or U16131 (N_16131,N_14077,N_15085);
xor U16132 (N_16132,N_15980,N_15403);
nand U16133 (N_16133,N_14977,N_15747);
xnor U16134 (N_16134,N_15263,N_14966);
nor U16135 (N_16135,N_15008,N_14868);
nor U16136 (N_16136,N_15715,N_14332);
xnor U16137 (N_16137,N_15765,N_14335);
nand U16138 (N_16138,N_14994,N_15414);
or U16139 (N_16139,N_15031,N_14576);
and U16140 (N_16140,N_15534,N_14999);
nor U16141 (N_16141,N_15066,N_15921);
nor U16142 (N_16142,N_14371,N_15694);
nand U16143 (N_16143,N_14640,N_14774);
nand U16144 (N_16144,N_14666,N_15802);
xor U16145 (N_16145,N_15384,N_15831);
nor U16146 (N_16146,N_14773,N_15213);
nor U16147 (N_16147,N_15443,N_15931);
nand U16148 (N_16148,N_15159,N_14196);
or U16149 (N_16149,N_15779,N_15547);
nand U16150 (N_16150,N_15590,N_14262);
nor U16151 (N_16151,N_15687,N_15731);
or U16152 (N_16152,N_14416,N_14746);
or U16153 (N_16153,N_14344,N_14625);
nor U16154 (N_16154,N_14448,N_14291);
nand U16155 (N_16155,N_14601,N_15737);
or U16156 (N_16156,N_15432,N_14284);
nand U16157 (N_16157,N_15270,N_14103);
nor U16158 (N_16158,N_14171,N_14988);
nand U16159 (N_16159,N_14845,N_15935);
nand U16160 (N_16160,N_14904,N_14516);
nand U16161 (N_16161,N_15758,N_15027);
nor U16162 (N_16162,N_15768,N_15914);
xnor U16163 (N_16163,N_15700,N_14295);
xnor U16164 (N_16164,N_15044,N_15956);
and U16165 (N_16165,N_15158,N_14177);
nand U16166 (N_16166,N_14958,N_14437);
nor U16167 (N_16167,N_14840,N_15448);
or U16168 (N_16168,N_14849,N_15954);
nand U16169 (N_16169,N_15026,N_15991);
and U16170 (N_16170,N_14940,N_14658);
nand U16171 (N_16171,N_15431,N_15583);
nand U16172 (N_16172,N_14470,N_15450);
or U16173 (N_16173,N_14689,N_14803);
or U16174 (N_16174,N_15476,N_14092);
nor U16175 (N_16175,N_14013,N_15098);
nor U16176 (N_16176,N_15096,N_14957);
nand U16177 (N_16177,N_14630,N_15284);
nor U16178 (N_16178,N_15668,N_15955);
and U16179 (N_16179,N_14238,N_14307);
nor U16180 (N_16180,N_14878,N_14603);
nand U16181 (N_16181,N_14128,N_15370);
and U16182 (N_16182,N_15901,N_14489);
nand U16183 (N_16183,N_15294,N_15495);
nand U16184 (N_16184,N_14954,N_15633);
xor U16185 (N_16185,N_15968,N_15876);
or U16186 (N_16186,N_15206,N_14216);
or U16187 (N_16187,N_14644,N_15656);
nor U16188 (N_16188,N_14674,N_14753);
xor U16189 (N_16189,N_14458,N_14102);
or U16190 (N_16190,N_14520,N_15413);
xnor U16191 (N_16191,N_15154,N_15364);
and U16192 (N_16192,N_15501,N_15690);
nor U16193 (N_16193,N_15922,N_15526);
nand U16194 (N_16194,N_14158,N_14760);
nor U16195 (N_16195,N_15515,N_15601);
nand U16196 (N_16196,N_14407,N_15251);
xnor U16197 (N_16197,N_15491,N_14794);
nor U16198 (N_16198,N_14302,N_15838);
or U16199 (N_16199,N_15199,N_14919);
nor U16200 (N_16200,N_15059,N_15354);
or U16201 (N_16201,N_14684,N_15361);
nor U16202 (N_16202,N_15880,N_15416);
nor U16203 (N_16203,N_14735,N_14943);
nor U16204 (N_16204,N_14285,N_14729);
and U16205 (N_16205,N_15685,N_15977);
nand U16206 (N_16206,N_14248,N_14373);
and U16207 (N_16207,N_14965,N_15540);
and U16208 (N_16208,N_15675,N_14927);
nand U16209 (N_16209,N_15082,N_14072);
nand U16210 (N_16210,N_15106,N_14428);
and U16211 (N_16211,N_14252,N_14832);
nand U16212 (N_16212,N_15383,N_15695);
and U16213 (N_16213,N_15759,N_14000);
xnor U16214 (N_16214,N_14443,N_15300);
nand U16215 (N_16215,N_15485,N_14595);
or U16216 (N_16216,N_15494,N_15829);
or U16217 (N_16217,N_15184,N_14384);
and U16218 (N_16218,N_15855,N_15025);
or U16219 (N_16219,N_15069,N_14914);
nor U16220 (N_16220,N_15138,N_14982);
and U16221 (N_16221,N_15220,N_14730);
and U16222 (N_16222,N_15397,N_15065);
xor U16223 (N_16223,N_15072,N_15915);
or U16224 (N_16224,N_14875,N_14577);
xnor U16225 (N_16225,N_15556,N_14974);
or U16226 (N_16226,N_14917,N_14787);
xnor U16227 (N_16227,N_15578,N_14476);
nor U16228 (N_16228,N_15645,N_15462);
or U16229 (N_16229,N_15869,N_14217);
and U16230 (N_16230,N_15271,N_15635);
and U16231 (N_16231,N_14949,N_14051);
or U16232 (N_16232,N_15187,N_15867);
nor U16233 (N_16233,N_15525,N_14218);
xor U16234 (N_16234,N_15328,N_15227);
or U16235 (N_16235,N_15461,N_14865);
or U16236 (N_16236,N_15095,N_14529);
and U16237 (N_16237,N_15619,N_14702);
or U16238 (N_16238,N_15075,N_15207);
nor U16239 (N_16239,N_15702,N_14108);
and U16240 (N_16240,N_14354,N_15298);
and U16241 (N_16241,N_15439,N_15899);
or U16242 (N_16242,N_15803,N_15290);
nor U16243 (N_16243,N_15508,N_15125);
nand U16244 (N_16244,N_14810,N_15171);
or U16245 (N_16245,N_15247,N_15372);
nand U16246 (N_16246,N_15216,N_14147);
nand U16247 (N_16247,N_14886,N_14410);
xnor U16248 (N_16248,N_14841,N_14442);
or U16249 (N_16249,N_14078,N_15058);
nor U16250 (N_16250,N_14236,N_15250);
nor U16251 (N_16251,N_15030,N_14992);
xor U16252 (N_16252,N_14194,N_14104);
xor U16253 (N_16253,N_14749,N_14019);
and U16254 (N_16254,N_15173,N_14846);
xor U16255 (N_16255,N_15099,N_15265);
xnor U16256 (N_16256,N_14806,N_14403);
nand U16257 (N_16257,N_15228,N_15873);
or U16258 (N_16258,N_15050,N_14491);
and U16259 (N_16259,N_14479,N_14242);
nand U16260 (N_16260,N_14681,N_15642);
xor U16261 (N_16261,N_15577,N_15239);
nand U16262 (N_16262,N_15183,N_14112);
or U16263 (N_16263,N_15032,N_14925);
nor U16264 (N_16264,N_14547,N_14151);
nand U16265 (N_16265,N_15490,N_14009);
nor U16266 (N_16266,N_15421,N_14752);
or U16267 (N_16267,N_15661,N_14271);
nor U16268 (N_16268,N_15045,N_14264);
xnor U16269 (N_16269,N_15712,N_15640);
or U16270 (N_16270,N_14311,N_14690);
nor U16271 (N_16271,N_14758,N_15975);
nor U16272 (N_16272,N_14754,N_15755);
nor U16273 (N_16273,N_14192,N_14465);
and U16274 (N_16274,N_15548,N_14152);
nor U16275 (N_16275,N_15516,N_14555);
xnor U16276 (N_16276,N_14662,N_14858);
xor U16277 (N_16277,N_15161,N_14861);
nand U16278 (N_16278,N_14148,N_14251);
or U16279 (N_16279,N_15283,N_15079);
nor U16280 (N_16280,N_14951,N_14498);
nor U16281 (N_16281,N_15850,N_14692);
nor U16282 (N_16282,N_15887,N_14174);
and U16283 (N_16283,N_15482,N_15157);
xnor U16284 (N_16284,N_14652,N_14930);
nand U16285 (N_16285,N_15120,N_14484);
nor U16286 (N_16286,N_15316,N_15103);
nor U16287 (N_16287,N_15410,N_15609);
nand U16288 (N_16288,N_14286,N_14481);
or U16289 (N_16289,N_15807,N_15389);
nor U16290 (N_16290,N_14785,N_14627);
nand U16291 (N_16291,N_15871,N_14967);
nand U16292 (N_16292,N_14346,N_15198);
nor U16293 (N_16293,N_14239,N_14256);
and U16294 (N_16294,N_15180,N_15519);
nor U16295 (N_16295,N_15615,N_14944);
nand U16296 (N_16296,N_14691,N_15697);
and U16297 (N_16297,N_15688,N_14895);
nor U16298 (N_16298,N_15276,N_15289);
xor U16299 (N_16299,N_14733,N_15456);
nor U16300 (N_16300,N_15539,N_15684);
or U16301 (N_16301,N_14558,N_15057);
nand U16302 (N_16302,N_15588,N_15463);
xor U16303 (N_16303,N_14046,N_14375);
or U16304 (N_16304,N_15714,N_14114);
nand U16305 (N_16305,N_14839,N_15438);
or U16306 (N_16306,N_14308,N_15840);
nor U16307 (N_16307,N_14215,N_14683);
nor U16308 (N_16308,N_14531,N_15986);
nor U16309 (N_16309,N_14317,N_15762);
nor U16310 (N_16310,N_15948,N_15314);
nor U16311 (N_16311,N_14117,N_15730);
or U16312 (N_16312,N_15068,N_15985);
and U16313 (N_16313,N_14227,N_15434);
nand U16314 (N_16314,N_15390,N_15719);
nand U16315 (N_16315,N_14029,N_14983);
or U16316 (N_16316,N_15744,N_14504);
and U16317 (N_16317,N_15823,N_14765);
nand U16318 (N_16318,N_15859,N_14153);
or U16319 (N_16319,N_15053,N_14208);
nand U16320 (N_16320,N_14620,N_15926);
and U16321 (N_16321,N_15393,N_14561);
nor U16322 (N_16322,N_14512,N_14010);
or U16323 (N_16323,N_14450,N_14997);
nand U16324 (N_16324,N_14824,N_14359);
nor U16325 (N_16325,N_15996,N_14331);
nand U16326 (N_16326,N_15524,N_14012);
nor U16327 (N_16327,N_14605,N_15606);
nand U16328 (N_16328,N_14517,N_14962);
nand U16329 (N_16329,N_14850,N_14036);
nand U16330 (N_16330,N_15426,N_14120);
nor U16331 (N_16331,N_15625,N_14705);
nand U16332 (N_16332,N_14935,N_14418);
and U16333 (N_16333,N_14290,N_15148);
nand U16334 (N_16334,N_15212,N_15732);
xnor U16335 (N_16335,N_14970,N_14769);
xnor U16336 (N_16336,N_15111,N_14015);
xnor U16337 (N_16337,N_14155,N_15232);
nand U16338 (N_16338,N_15629,N_15430);
or U16339 (N_16339,N_15949,N_15155);
xnor U16340 (N_16340,N_15834,N_15570);
xor U16341 (N_16341,N_14380,N_14883);
nor U16342 (N_16342,N_15381,N_14621);
nand U16343 (N_16343,N_14973,N_14368);
xnor U16344 (N_16344,N_14678,N_15725);
nor U16345 (N_16345,N_14096,N_15153);
nor U16346 (N_16346,N_14197,N_15884);
nor U16347 (N_16347,N_14135,N_15160);
nand U16348 (N_16348,N_14341,N_15377);
nor U16349 (N_16349,N_14105,N_15221);
nor U16350 (N_16350,N_14362,N_15821);
and U16351 (N_16351,N_14214,N_14023);
nor U16352 (N_16352,N_15402,N_15784);
or U16353 (N_16353,N_14802,N_14641);
nor U16354 (N_16354,N_15822,N_14900);
nand U16355 (N_16355,N_15550,N_15594);
and U16356 (N_16356,N_15541,N_14088);
nor U16357 (N_16357,N_14539,N_14819);
or U16358 (N_16358,N_14496,N_14634);
or U16359 (N_16359,N_15401,N_14998);
nor U16360 (N_16360,N_14224,N_14888);
and U16361 (N_16361,N_15551,N_14002);
and U16362 (N_16362,N_15614,N_15132);
xnor U16363 (N_16363,N_14844,N_14435);
nor U16364 (N_16364,N_15282,N_15860);
xor U16365 (N_16365,N_15654,N_15766);
and U16366 (N_16366,N_15483,N_14656);
or U16367 (N_16367,N_15444,N_15958);
nand U16368 (N_16368,N_15795,N_15165);
and U16369 (N_16369,N_15943,N_14617);
xnor U16370 (N_16370,N_14899,N_14993);
nor U16371 (N_16371,N_15293,N_15669);
xnor U16372 (N_16372,N_15637,N_15983);
and U16373 (N_16373,N_15567,N_15704);
or U16374 (N_16374,N_15713,N_14055);
nor U16375 (N_16375,N_15424,N_14908);
or U16376 (N_16376,N_14959,N_14645);
nand U16377 (N_16377,N_15708,N_15767);
and U16378 (N_16378,N_15734,N_14777);
nand U16379 (N_16379,N_14048,N_14697);
nor U16380 (N_16380,N_14981,N_15969);
and U16381 (N_16381,N_14772,N_14265);
xor U16382 (N_16382,N_14540,N_15726);
xor U16383 (N_16383,N_14657,N_14425);
nor U16384 (N_16384,N_14654,N_15957);
or U16385 (N_16385,N_14318,N_14074);
nor U16386 (N_16386,N_15367,N_14747);
xor U16387 (N_16387,N_15122,N_14414);
xor U16388 (N_16388,N_14024,N_14898);
or U16389 (N_16389,N_14671,N_14320);
xnor U16390 (N_16390,N_14811,N_15427);
nand U16391 (N_16391,N_14708,N_15587);
or U16392 (N_16392,N_14433,N_14272);
or U16393 (N_16393,N_15077,N_14424);
nand U16394 (N_16394,N_15878,N_14165);
xor U16395 (N_16395,N_14313,N_15959);
or U16396 (N_16396,N_15315,N_15035);
xor U16397 (N_16397,N_15751,N_14590);
nand U16398 (N_16398,N_15617,N_14137);
nor U16399 (N_16399,N_14528,N_15447);
and U16400 (N_16400,N_15607,N_14892);
nand U16401 (N_16401,N_14722,N_14805);
xnor U16402 (N_16402,N_15409,N_14404);
nand U16403 (N_16403,N_14820,N_14101);
xnor U16404 (N_16404,N_15819,N_15353);
xor U16405 (N_16405,N_15611,N_15280);
xor U16406 (N_16406,N_15144,N_14606);
and U16407 (N_16407,N_14490,N_14255);
nor U16408 (N_16408,N_14542,N_14043);
or U16409 (N_16409,N_15561,N_15405);
nor U16410 (N_16410,N_15357,N_14989);
nand U16411 (N_16411,N_14062,N_15960);
nand U16412 (N_16412,N_14807,N_15110);
and U16413 (N_16413,N_15814,N_15193);
or U16414 (N_16414,N_15406,N_15893);
nand U16415 (N_16415,N_14737,N_14881);
nand U16416 (N_16416,N_14168,N_14203);
and U16417 (N_16417,N_15705,N_14783);
nand U16418 (N_16418,N_14179,N_15889);
nor U16419 (N_16419,N_15235,N_15327);
nor U16420 (N_16420,N_14987,N_14070);
nand U16421 (N_16421,N_15788,N_15787);
xor U16422 (N_16422,N_14379,N_15681);
or U16423 (N_16423,N_15083,N_14358);
and U16424 (N_16424,N_15238,N_14638);
nand U16425 (N_16425,N_14231,N_15781);
nand U16426 (N_16426,N_14750,N_15337);
xnor U16427 (N_16427,N_14474,N_15805);
nand U16428 (N_16428,N_15740,N_14503);
and U16429 (N_16429,N_15176,N_14008);
nor U16430 (N_16430,N_15043,N_14816);
and U16431 (N_16431,N_15659,N_15892);
nor U16432 (N_16432,N_15380,N_14025);
nand U16433 (N_16433,N_15496,N_14928);
xor U16434 (N_16434,N_15185,N_14902);
nor U16435 (N_16435,N_14360,N_15832);
nand U16436 (N_16436,N_14432,N_14267);
nand U16437 (N_16437,N_15189,N_14514);
and U16438 (N_16438,N_15792,N_14582);
nor U16439 (N_16439,N_14763,N_15529);
nor U16440 (N_16440,N_15825,N_14623);
nand U16441 (N_16441,N_14200,N_15569);
or U16442 (N_16442,N_14759,N_14412);
and U16443 (N_16443,N_15939,N_14040);
xnor U16444 (N_16444,N_14035,N_15984);
and U16445 (N_16445,N_15150,N_14543);
nand U16446 (N_16446,N_15062,N_14052);
nor U16447 (N_16447,N_14650,N_15387);
xor U16448 (N_16448,N_14609,N_15311);
and U16449 (N_16449,N_14725,N_15924);
xnor U16450 (N_16450,N_14429,N_15299);
xor U16451 (N_16451,N_14534,N_15835);
xor U16452 (N_16452,N_15683,N_14065);
nand U16453 (N_16453,N_14507,N_15029);
nor U16454 (N_16454,N_14471,N_15188);
nor U16455 (N_16455,N_14388,N_15359);
nand U16456 (N_16456,N_15809,N_15244);
nand U16457 (N_16457,N_14085,N_14619);
and U16458 (N_16458,N_14731,N_14890);
nor U16459 (N_16459,N_15269,N_15741);
or U16460 (N_16460,N_15142,N_14007);
or U16461 (N_16461,N_15517,N_15979);
or U16462 (N_16462,N_15798,N_14995);
and U16463 (N_16463,N_15783,N_15890);
and U16464 (N_16464,N_15665,N_14365);
and U16465 (N_16465,N_14639,N_15001);
nor U16466 (N_16466,N_15362,N_15022);
and U16467 (N_16467,N_14109,N_15004);
nor U16468 (N_16468,N_14701,N_14508);
or U16469 (N_16469,N_14668,N_14202);
and U16470 (N_16470,N_14323,N_15114);
or U16471 (N_16471,N_14210,N_14081);
nand U16472 (N_16472,N_14703,N_14969);
xnor U16473 (N_16473,N_14564,N_15776);
nand U16474 (N_16474,N_14439,N_15673);
nor U16475 (N_16475,N_14933,N_14205);
xnor U16476 (N_16476,N_14268,N_14466);
xnor U16477 (N_16477,N_14756,N_15699);
and U16478 (N_16478,N_14600,N_15319);
or U16479 (N_16479,N_15874,N_15895);
nor U16480 (N_16480,N_14084,N_15896);
and U16481 (N_16481,N_14509,N_14243);
nand U16482 (N_16482,N_15507,N_14326);
nor U16483 (N_16483,N_15260,N_15310);
nor U16484 (N_16484,N_15827,N_15571);
xor U16485 (N_16485,N_14506,N_14377);
nand U16486 (N_16486,N_14926,N_14486);
and U16487 (N_16487,N_15287,N_14107);
nor U16488 (N_16488,N_14452,N_15317);
xor U16489 (N_16489,N_14337,N_15771);
xnor U16490 (N_16490,N_15071,N_14884);
or U16491 (N_16491,N_14306,N_15179);
xnor U16492 (N_16492,N_14342,N_14867);
nor U16493 (N_16493,N_14647,N_14667);
nand U16494 (N_16494,N_15801,N_15385);
xor U16495 (N_16495,N_15863,N_14673);
nor U16496 (N_16496,N_14319,N_14406);
nor U16497 (N_16497,N_14677,N_14441);
xor U16498 (N_16498,N_15521,N_15209);
and U16499 (N_16499,N_14176,N_15942);
nand U16500 (N_16500,N_14169,N_15277);
xnor U16501 (N_16501,N_15603,N_15107);
nand U16502 (N_16502,N_15226,N_14814);
or U16503 (N_16503,N_14823,N_14812);
nand U16504 (N_16504,N_14383,N_14929);
nor U16505 (N_16505,N_15033,N_14593);
nor U16506 (N_16506,N_14732,N_14495);
nand U16507 (N_16507,N_14166,N_14309);
or U16508 (N_16508,N_14911,N_15054);
and U16509 (N_16509,N_14339,N_15296);
or U16510 (N_16510,N_14419,N_14206);
nor U16511 (N_16511,N_15729,N_15049);
xnor U16512 (N_16512,N_14488,N_14294);
xor U16513 (N_16513,N_14041,N_14279);
xor U16514 (N_16514,N_15064,N_14340);
or U16515 (N_16515,N_15457,N_14766);
xor U16516 (N_16516,N_15999,N_15808);
nand U16517 (N_16517,N_14838,N_15428);
nand U16518 (N_16518,N_15903,N_14633);
xor U16519 (N_16519,N_15682,N_15976);
nand U16520 (N_16520,N_15538,N_14001);
or U16521 (N_16521,N_14187,N_14562);
or U16522 (N_16522,N_14315,N_15080);
or U16523 (N_16523,N_15486,N_15817);
nand U16524 (N_16524,N_14960,N_14063);
xor U16525 (N_16525,N_15343,N_15313);
or U16526 (N_16526,N_15854,N_14330);
nand U16527 (N_16527,N_14978,N_15910);
xnor U16528 (N_16528,N_15974,N_15170);
xnor U16529 (N_16529,N_15973,N_15618);
or U16530 (N_16530,N_14523,N_14872);
and U16531 (N_16531,N_15568,N_14946);
nand U16532 (N_16532,N_14597,N_15329);
and U16533 (N_16533,N_15990,N_15522);
xor U16534 (N_16534,N_14314,N_14563);
and U16535 (N_16535,N_14511,N_15511);
xnor U16536 (N_16536,N_15630,N_14198);
xor U16537 (N_16537,N_14519,N_15021);
nor U16538 (N_16538,N_14086,N_14420);
nor U16539 (N_16539,N_15811,N_14535);
nor U16540 (N_16540,N_14585,N_15846);
or U16541 (N_16541,N_15325,N_14566);
or U16542 (N_16542,N_14724,N_15575);
or U16543 (N_16543,N_15196,N_15906);
or U16544 (N_16544,N_15477,N_15453);
xnor U16545 (N_16545,N_15902,N_15870);
and U16546 (N_16546,N_14396,N_15940);
xnor U16547 (N_16547,N_14032,N_15543);
nand U16548 (N_16548,N_15350,N_15131);
nor U16549 (N_16549,N_15667,N_15423);
nand U16550 (N_16550,N_14226,N_14906);
xor U16551 (N_16551,N_15373,N_14575);
nor U16552 (N_16552,N_15446,N_15552);
and U16553 (N_16553,N_14310,N_14986);
xor U16554 (N_16554,N_14778,N_15394);
nand U16555 (N_16555,N_14853,N_14903);
xnor U16556 (N_16556,N_15558,N_14188);
nor U16557 (N_16557,N_15579,N_15169);
nand U16558 (N_16558,N_14893,N_14113);
and U16559 (N_16559,N_14980,N_14990);
nand U16560 (N_16560,N_15919,N_14207);
xor U16561 (N_16561,N_14376,N_14494);
nor U16562 (N_16562,N_14282,N_15865);
nand U16563 (N_16563,N_15230,N_14149);
or U16564 (N_16564,N_14530,N_15091);
nor U16565 (N_16565,N_15849,N_15060);
nand U16566 (N_16566,N_14175,N_15356);
xor U16567 (N_16567,N_15881,N_15420);
xnor U16568 (N_16568,N_14276,N_14624);
xor U16569 (N_16569,N_15650,N_14061);
and U16570 (N_16570,N_14991,N_15168);
xor U16571 (N_16571,N_14776,N_15399);
or U16572 (N_16572,N_15475,N_14685);
nor U16573 (N_16573,N_15753,N_14030);
nand U16574 (N_16574,N_15012,N_14400);
or U16575 (N_16575,N_14822,N_15791);
and U16576 (N_16576,N_15506,N_14552);
xnor U16577 (N_16577,N_14363,N_14178);
xnor U16578 (N_16578,N_15215,N_14080);
xnor U16579 (N_16579,N_14324,N_14343);
nor U16580 (N_16580,N_14082,N_14180);
and U16581 (N_16581,N_14364,N_15936);
and U16582 (N_16582,N_15113,N_14831);
nand U16583 (N_16583,N_15717,N_14791);
nand U16584 (N_16584,N_15549,N_15929);
and U16585 (N_16585,N_15912,N_15092);
nand U16586 (N_16586,N_14586,N_14544);
nand U16587 (N_16587,N_14089,N_15487);
xnor U16588 (N_16588,N_14461,N_14246);
xor U16589 (N_16589,N_15591,N_14515);
nand U16590 (N_16590,N_15626,N_15988);
nand U16591 (N_16591,N_14044,N_14297);
xnor U16592 (N_16592,N_14796,N_15152);
or U16593 (N_16593,N_14438,N_15203);
nand U16594 (N_16594,N_15833,N_15369);
and U16595 (N_16595,N_15572,N_14714);
nand U16596 (N_16596,N_14223,N_14316);
nor U16597 (N_16597,N_14580,N_15304);
and U16598 (N_16598,N_14871,N_15565);
or U16599 (N_16599,N_14936,N_15019);
nand U16600 (N_16600,N_14522,N_14592);
nor U16601 (N_16601,N_14181,N_14327);
xnor U16602 (N_16602,N_15581,N_14393);
and U16603 (N_16603,N_15376,N_15466);
and U16604 (N_16604,N_14119,N_14855);
nand U16605 (N_16605,N_15470,N_15225);
nand U16606 (N_16606,N_14613,N_15345);
nor U16607 (N_16607,N_14003,N_15670);
and U16608 (N_16608,N_14956,N_14115);
and U16609 (N_16609,N_14123,N_15288);
and U16610 (N_16610,N_15404,N_14399);
and U16611 (N_16611,N_15078,N_14150);
nor U16612 (N_16612,N_15782,N_14538);
nor U16613 (N_16613,N_14790,N_15326);
nand U16614 (N_16614,N_14126,N_14661);
and U16615 (N_16615,N_15378,N_14423);
or U16616 (N_16616,N_14616,N_15321);
nand U16617 (N_16617,N_15346,N_14367);
nor U16618 (N_16618,N_15644,N_15662);
nand U16619 (N_16619,N_15433,N_14230);
and U16620 (N_16620,N_15141,N_14028);
and U16621 (N_16621,N_14779,N_15386);
nand U16622 (N_16622,N_14764,N_14136);
xnor U16623 (N_16623,N_15716,N_15465);
or U16624 (N_16624,N_15648,N_15677);
xnor U16625 (N_16625,N_15864,N_15918);
or U16626 (N_16626,N_15023,N_14321);
nand U16627 (N_16627,N_14229,N_15348);
or U16628 (N_16628,N_15074,N_15097);
or U16629 (N_16629,N_15813,N_14333);
or U16630 (N_16630,N_15102,N_15925);
or U16631 (N_16631,N_14301,N_15488);
and U16632 (N_16632,N_15613,N_14847);
nor U16633 (N_16633,N_14095,N_15841);
nand U16634 (N_16634,N_15651,N_14006);
and U16635 (N_16635,N_15301,N_14444);
or U16636 (N_16636,N_14880,N_14795);
nand U16637 (N_16637,N_14170,N_15643);
xnor U16638 (N_16638,N_14642,N_15255);
nor U16639 (N_16639,N_15858,N_14655);
or U16640 (N_16640,N_15582,N_15498);
and U16641 (N_16641,N_15815,N_15934);
and U16642 (N_16642,N_14937,N_14430);
xnor U16643 (N_16643,N_15953,N_15395);
or U16644 (N_16644,N_14622,N_14955);
nor U16645 (N_16645,N_14793,N_14583);
nand U16646 (N_16646,N_14713,N_14913);
xnor U16647 (N_16647,N_14305,N_15219);
nand U16648 (N_16648,N_15718,N_15907);
nand U16649 (N_16649,N_15573,N_14047);
or U16650 (N_16650,N_15459,N_15738);
nand U16651 (N_16651,N_14300,N_15339);
nor U16652 (N_16652,N_15763,N_15217);
nand U16653 (N_16653,N_14579,N_15084);
or U16654 (N_16654,N_15360,N_15493);
xnor U16655 (N_16655,N_14525,N_15962);
and U16656 (N_16656,N_15856,N_14021);
nand U16657 (N_16657,N_14381,N_15341);
or U16658 (N_16658,N_15200,N_15720);
and U16659 (N_16659,N_15596,N_15267);
nand U16660 (N_16660,N_15502,N_14069);
nor U16661 (N_16661,N_15324,N_15191);
nor U16662 (N_16662,N_14626,N_14034);
xor U16663 (N_16663,N_14415,N_15503);
nand U16664 (N_16664,N_15998,N_14887);
xor U16665 (N_16665,N_14038,N_14804);
or U16666 (N_16666,N_14411,N_15920);
and U16667 (N_16667,N_14891,N_14056);
nand U16668 (N_16668,N_14941,N_15192);
nor U16669 (N_16669,N_14385,N_14234);
nand U16670 (N_16670,N_15013,N_15037);
xor U16671 (N_16671,N_15818,N_14510);
or U16672 (N_16672,N_14042,N_14211);
nor U16673 (N_16673,N_14222,N_15789);
xor U16674 (N_16674,N_15723,N_14142);
and U16675 (N_16675,N_15852,N_14923);
and U16676 (N_16676,N_15055,N_15070);
nor U16677 (N_16677,N_15599,N_14897);
nor U16678 (N_16678,N_14386,N_14277);
and U16679 (N_16679,N_14289,N_15544);
nand U16680 (N_16680,N_15143,N_14445);
nor U16681 (N_16681,N_14918,N_15115);
and U16682 (N_16682,N_14453,N_15039);
nor U16683 (N_16683,N_14964,N_15557);
xnor U16684 (N_16684,N_15647,N_14258);
nand U16685 (N_16685,N_14636,N_15163);
nor U16686 (N_16686,N_14553,N_14212);
and U16687 (N_16687,N_14532,N_15081);
or U16688 (N_16688,N_14546,N_15897);
nand U16689 (N_16689,N_15145,N_14932);
xor U16690 (N_16690,N_15610,N_15139);
nor U16691 (N_16691,N_15305,N_15109);
xor U16692 (N_16692,N_15652,N_15923);
nor U16693 (N_16693,N_14249,N_15272);
and U16694 (N_16694,N_15347,N_15703);
nor U16695 (N_16695,N_15237,N_15038);
xnor U16696 (N_16696,N_14734,N_14696);
xor U16697 (N_16697,N_15756,N_15666);
or U16698 (N_16698,N_14718,N_14356);
xor U16699 (N_16699,N_14334,N_15087);
or U16700 (N_16700,N_14060,N_15844);
and U16701 (N_16701,N_14401,N_14213);
xor U16702 (N_16702,N_14780,N_14915);
and U16703 (N_16703,N_15853,N_15415);
nand U16704 (N_16704,N_15440,N_15422);
nand U16705 (N_16705,N_15660,N_15499);
xor U16706 (N_16706,N_15309,N_15036);
or U16707 (N_16707,N_14160,N_15743);
nor U16708 (N_16708,N_15484,N_15112);
or U16709 (N_16709,N_15913,N_14093);
nor U16710 (N_16710,N_15698,N_15520);
xnor U16711 (N_16711,N_14132,N_14468);
nor U16712 (N_16712,N_14771,N_14253);
and U16713 (N_16713,N_15437,N_15351);
nand U16714 (N_16714,N_15133,N_15166);
nor U16715 (N_16715,N_14161,N_15847);
or U16716 (N_16716,N_14283,N_15848);
xor U16717 (N_16717,N_14016,N_15535);
nor U16718 (N_16718,N_15391,N_14184);
nand U16719 (N_16719,N_15467,N_14322);
and U16720 (N_16720,N_15862,N_15553);
xnor U16721 (N_16721,N_14349,N_15997);
or U16722 (N_16722,N_15275,N_15307);
or U16723 (N_16723,N_14834,N_14357);
nand U16724 (N_16724,N_14896,N_15658);
and U16725 (N_16725,N_14394,N_15040);
nor U16726 (N_16726,N_15214,N_15750);
nor U16727 (N_16727,N_15891,N_14131);
or U16728 (N_16728,N_14976,N_14457);
or U16729 (N_16729,N_15664,N_15471);
nor U16730 (N_16730,N_15671,N_14185);
or U16731 (N_16731,N_14145,N_14083);
xnor U16732 (N_16732,N_15696,N_14821);
nor U16733 (N_16733,N_14066,N_14825);
nor U16734 (N_16734,N_15268,N_14312);
nor U16735 (N_16735,N_14653,N_15007);
or U16736 (N_16736,N_14139,N_14167);
xor U16737 (N_16737,N_15875,N_15210);
xnor U16738 (N_16738,N_15140,N_15266);
and U16739 (N_16739,N_14874,N_15128);
and U16740 (N_16740,N_15342,N_15489);
xor U16741 (N_16741,N_14460,N_15632);
nor U16742 (N_16742,N_15211,N_14280);
nand U16743 (N_16743,N_15468,N_15894);
nand U16744 (N_16744,N_15937,N_15602);
nand U16745 (N_16745,N_15249,N_14799);
or U16746 (N_16746,N_14843,N_15460);
and U16747 (N_16747,N_14374,N_15800);
or U16748 (N_16748,N_14743,N_14830);
xnor U16749 (N_16749,N_14545,N_15911);
nor U16750 (N_16750,N_15331,N_14632);
xor U16751 (N_16751,N_14612,N_15047);
or U16752 (N_16752,N_14455,N_14859);
nand U16753 (N_16753,N_15382,N_14568);
xnor U16754 (N_16754,N_14391,N_15739);
and U16755 (N_16755,N_14560,N_14502);
nor U16756 (N_16756,N_15190,N_15312);
nor U16757 (N_16757,N_14098,N_15441);
or U16758 (N_16758,N_15646,N_14587);
xor U16759 (N_16759,N_14828,N_14106);
xor U16760 (N_16760,N_14672,N_14121);
xor U16761 (N_16761,N_14975,N_15686);
xor U16762 (N_16762,N_14501,N_14781);
or U16763 (N_16763,N_15754,N_14770);
nand U16764 (N_16764,N_14049,N_15966);
nor U16765 (N_16765,N_14594,N_14492);
or U16766 (N_16766,N_15252,N_14449);
and U16767 (N_16767,N_14837,N_15253);
nor U16768 (N_16768,N_15679,N_15323);
and U16769 (N_16769,N_15736,N_15146);
xor U16770 (N_16770,N_15812,N_14201);
nand U16771 (N_16771,N_14499,N_14274);
nor U16772 (N_16772,N_15745,N_14447);
nand U16773 (N_16773,N_15830,N_14784);
nor U16774 (N_16774,N_15222,N_15820);
nor U16775 (N_16775,N_14050,N_15355);
or U16776 (N_16776,N_15711,N_15970);
nand U16777 (N_16777,N_15264,N_14798);
or U16778 (N_16778,N_14797,N_14693);
or U16779 (N_16779,N_15777,N_15088);
or U16780 (N_16780,N_15116,N_14347);
or U16781 (N_16781,N_14191,N_14704);
xor U16782 (N_16782,N_15308,N_14631);
nand U16783 (N_16783,N_15627,N_14527);
and U16784 (N_16784,N_15469,N_14570);
nand U16785 (N_16785,N_15286,N_14451);
and U16786 (N_16786,N_15612,N_15481);
nand U16787 (N_16787,N_14183,N_14366);
nor U16788 (N_16788,N_14011,N_14680);
and U16789 (N_16789,N_15400,N_15982);
xnor U16790 (N_16790,N_15218,N_15042);
xor U16791 (N_16791,N_14328,N_15243);
and U16792 (N_16792,N_14464,N_15261);
nor U16793 (N_16793,N_15773,N_14894);
nor U16794 (N_16794,N_14740,N_14436);
and U16795 (N_16795,N_15932,N_14110);
xnor U16796 (N_16796,N_15947,N_15051);
nor U16797 (N_16797,N_15972,N_15678);
xnor U16798 (N_16798,N_14757,N_15992);
xor U16799 (N_16799,N_15186,N_14809);
nand U16800 (N_16800,N_15728,N_14996);
nand U16801 (N_16801,N_15474,N_15041);
nor U16802 (N_16802,N_14100,N_15592);
nand U16803 (N_16803,N_14116,N_14826);
and U16804 (N_16804,N_14775,N_15352);
nor U16805 (N_16805,N_14369,N_15981);
xor U16806 (N_16806,N_14204,N_15175);
nor U16807 (N_16807,N_14842,N_14027);
nand U16808 (N_16808,N_15576,N_15204);
or U16809 (N_16809,N_15090,N_14058);
xor U16810 (N_16810,N_15254,N_15930);
nand U16811 (N_16811,N_15320,N_15231);
xor U16812 (N_16812,N_14138,N_15229);
nand U16813 (N_16813,N_14459,N_14130);
nor U16814 (N_16814,N_14715,N_15882);
or U16815 (N_16815,N_14348,N_15365);
nand U16816 (N_16816,N_14905,N_14591);
or U16817 (N_16817,N_14004,N_15532);
xnor U16818 (N_16818,N_14869,N_14303);
and U16819 (N_16819,N_15604,N_14726);
nand U16820 (N_16820,N_15472,N_15879);
xor U16821 (N_16821,N_15514,N_14789);
and U16822 (N_16822,N_14257,N_15554);
xnor U16823 (N_16823,N_15295,N_14020);
nor U16824 (N_16824,N_15407,N_14405);
or U16825 (N_16825,N_15492,N_15772);
xor U16826 (N_16826,N_14712,N_14945);
nor U16827 (N_16827,N_15018,N_15566);
or U16828 (N_16828,N_15086,N_14281);
nor U16829 (N_16829,N_14608,N_14261);
and U16830 (N_16830,N_14018,N_15995);
or U16831 (N_16831,N_15117,N_15454);
nand U16832 (N_16832,N_14014,N_15574);
nor U16833 (N_16833,N_15837,N_15790);
nor U16834 (N_16834,N_14767,N_15451);
or U16835 (N_16835,N_15951,N_14288);
nor U16836 (N_16836,N_15358,N_15689);
or U16837 (N_16837,N_15010,N_15151);
xnor U16838 (N_16838,N_14699,N_15888);
or U16839 (N_16839,N_14876,N_15908);
nor U16840 (N_16840,N_15375,N_14372);
nand U16841 (N_16841,N_14581,N_14475);
or U16842 (N_16842,N_14270,N_14610);
xor U16843 (N_16843,N_15804,N_14596);
or U16844 (N_16844,N_15101,N_15916);
nand U16845 (N_16845,N_14336,N_15174);
or U16846 (N_16846,N_15015,N_14660);
or U16847 (N_16847,N_14635,N_14736);
xor U16848 (N_16848,N_14141,N_14686);
xor U16849 (N_16849,N_15000,N_15877);
xor U16850 (N_16850,N_14574,N_15523);
nor U16851 (N_16851,N_15584,N_14408);
nor U16852 (N_16852,N_14800,N_15692);
and U16853 (N_16853,N_15796,N_14604);
and U16854 (N_16854,N_14885,N_15335);
and U16855 (N_16855,N_15598,N_14901);
nor U16856 (N_16856,N_14304,N_14924);
and U16857 (N_16857,N_14879,N_14971);
or U16858 (N_16858,N_15770,N_14352);
nand U16859 (N_16859,N_14244,N_15760);
and U16860 (N_16860,N_14263,N_14910);
or U16861 (N_16861,N_14866,N_14611);
or U16862 (N_16862,N_14067,N_15746);
xnor U16863 (N_16863,N_14240,N_14675);
and U16864 (N_16864,N_15799,N_15129);
or U16865 (N_16865,N_15563,N_15014);
nand U16866 (N_16866,N_14467,N_15774);
and U16867 (N_16867,N_14651,N_14939);
nor U16868 (N_16868,N_15733,N_14037);
and U16869 (N_16869,N_15223,N_14090);
or U16870 (N_16870,N_14614,N_15135);
or U16871 (N_16871,N_14162,N_15435);
nand U16872 (N_16872,N_14146,N_15061);
or U16873 (N_16873,N_15224,N_14857);
nand U16874 (N_16874,N_14762,N_15769);
and U16875 (N_16875,N_14801,N_15707);
xnor U16876 (N_16876,N_15076,N_15964);
xor U16877 (N_16877,N_15628,N_14578);
or U16878 (N_16878,N_14053,N_14852);
nand U16879 (N_16879,N_15392,N_14985);
nand U16880 (N_16880,N_14127,N_15147);
nor U16881 (N_16881,N_14382,N_14143);
nor U16882 (N_16882,N_15412,N_14827);
nor U16883 (N_16883,N_14856,N_14073);
or U16884 (N_16884,N_14125,N_14209);
xnor U16885 (N_16885,N_15872,N_14076);
nor U16886 (N_16886,N_14584,N_15182);
and U16887 (N_16887,N_14087,N_15639);
nand U16888 (N_16888,N_14864,N_15655);
and U16889 (N_16889,N_14663,N_14755);
nand U16890 (N_16890,N_15242,N_14482);
nor U16891 (N_16891,N_15631,N_14079);
or U16892 (N_16892,N_14245,N_15349);
and U16893 (N_16893,N_15419,N_15398);
xnor U16894 (N_16894,N_15710,N_14862);
nor U16895 (N_16895,N_14235,N_15504);
and U16896 (N_16896,N_15322,N_15089);
xor U16897 (N_16897,N_15234,N_14189);
or U16898 (N_16898,N_15680,N_15104);
xor U16899 (N_16899,N_15616,N_14292);
xnor U16900 (N_16900,N_14195,N_14533);
or U16901 (N_16901,N_14953,N_14835);
or U16902 (N_16902,N_14513,N_15258);
or U16903 (N_16903,N_14815,N_14646);
and U16904 (N_16904,N_14099,N_15478);
nand U16905 (N_16905,N_15898,N_15672);
and U16906 (N_16906,N_15330,N_15417);
or U16907 (N_16907,N_15836,N_14599);
nand U16908 (N_16908,N_14427,N_14719);
nand U16909 (N_16909,N_15429,N_15336);
or U16910 (N_16910,N_15861,N_14744);
nand U16911 (N_16911,N_15993,N_15509);
nor U16912 (N_16912,N_14293,N_15851);
and U16913 (N_16913,N_15810,N_15046);
or U16914 (N_16914,N_14022,N_14559);
or U16915 (N_16915,N_15512,N_14039);
nand U16916 (N_16916,N_14836,N_15205);
nand U16917 (N_16917,N_15634,N_14421);
or U16918 (N_16918,N_15528,N_14549);
or U16919 (N_16919,N_14711,N_14938);
xnor U16920 (N_16920,N_15971,N_14979);
nand U16921 (N_16921,N_15197,N_15302);
xor U16922 (N_16922,N_14033,N_15593);
nor U16923 (N_16923,N_15105,N_15724);
and U16924 (N_16924,N_15020,N_14017);
nand U16925 (N_16925,N_15857,N_15886);
nor U16926 (N_16926,N_15786,N_15118);
nand U16927 (N_16927,N_15938,N_15363);
or U16928 (N_16928,N_15338,N_15775);
or U16929 (N_16929,N_15318,N_15181);
nand U16930 (N_16930,N_14064,N_14140);
nor U16931 (N_16931,N_14741,N_14500);
nor U16932 (N_16932,N_14573,N_15586);
and U16933 (N_16933,N_15034,N_14912);
nor U16934 (N_16934,N_14947,N_15513);
nor U16935 (N_16935,N_15442,N_15595);
nand U16936 (N_16936,N_14361,N_15555);
nor U16937 (N_16937,N_14172,N_15194);
nand U16938 (N_16938,N_15425,N_15167);
and U16939 (N_16939,N_15011,N_15709);
or U16940 (N_16940,N_14676,N_14968);
or U16941 (N_16941,N_15620,N_15564);
and U16942 (N_16942,N_14889,N_15748);
xnor U16943 (N_16943,N_14031,N_14273);
and U16944 (N_16944,N_14199,N_15149);
xnor U16945 (N_16945,N_15464,N_15605);
nor U16946 (N_16946,N_15764,N_14260);
nand U16947 (N_16947,N_15334,N_14250);
nor U16948 (N_16948,N_15108,N_15006);
xnor U16949 (N_16949,N_14097,N_14164);
xnor U16950 (N_16950,N_15638,N_15676);
nand U16951 (N_16951,N_15905,N_15621);
or U16952 (N_16952,N_15826,N_15396);
nor U16953 (N_16953,N_15824,N_15245);
nor U16954 (N_16954,N_14720,N_14469);
nor U16955 (N_16955,N_14446,N_15366);
and U16956 (N_16956,N_14350,N_14091);
or U16957 (N_16957,N_14536,N_14963);
nor U16958 (N_16958,N_14483,N_14237);
nand U16959 (N_16959,N_15649,N_15944);
nand U16960 (N_16960,N_15641,N_15693);
and U16961 (N_16961,N_15126,N_15636);
xnor U16962 (N_16962,N_14728,N_14848);
or U16963 (N_16963,N_14709,N_14808);
nand U16964 (N_16964,N_14524,N_15794);
and U16965 (N_16965,N_14518,N_14710);
and U16966 (N_16966,N_14259,N_15527);
nand U16967 (N_16967,N_14768,N_14572);
and U16968 (N_16968,N_14727,N_14829);
nand U16969 (N_16969,N_15885,N_15246);
xnor U16970 (N_16970,N_15274,N_15589);
and U16971 (N_16971,N_14493,N_14643);
nor U16972 (N_16972,N_15545,N_14228);
and U16973 (N_16973,N_14220,N_15945);
and U16974 (N_16974,N_15048,N_14551);
nor U16975 (N_16975,N_14628,N_15778);
nor U16976 (N_16976,N_15600,N_14782);
or U16977 (N_16977,N_14472,N_14497);
and U16978 (N_16978,N_14390,N_15100);
or U16979 (N_16979,N_14057,N_14392);
nor U16980 (N_16980,N_14554,N_15727);
nand U16981 (N_16981,N_14909,N_14417);
and U16982 (N_16982,N_15202,N_14669);
or U16983 (N_16983,N_15121,N_14761);
nand U16984 (N_16984,N_15904,N_15622);
and U16985 (N_16985,N_15965,N_15691);
and U16986 (N_16986,N_14124,N_14485);
nor U16987 (N_16987,N_14569,N_14219);
nand U16988 (N_16988,N_14818,N_15248);
nor U16989 (N_16989,N_15285,N_15473);
xor U16990 (N_16990,N_14629,N_14345);
nor U16991 (N_16991,N_15536,N_15735);
nand U16992 (N_16992,N_15961,N_15303);
and U16993 (N_16993,N_15560,N_15073);
nor U16994 (N_16994,N_14426,N_15445);
nand U16995 (N_16995,N_15933,N_15706);
and U16996 (N_16996,N_15172,N_15306);
nor U16997 (N_16997,N_14378,N_14122);
nand U16998 (N_16998,N_15002,N_14851);
or U16999 (N_16999,N_14163,N_14389);
nand U17000 (N_17000,N_15755,N_14397);
and U17001 (N_17001,N_14135,N_14607);
nor U17002 (N_17002,N_15128,N_14907);
or U17003 (N_17003,N_15832,N_15658);
nor U17004 (N_17004,N_14292,N_15403);
and U17005 (N_17005,N_14802,N_15595);
nor U17006 (N_17006,N_15814,N_14072);
or U17007 (N_17007,N_15255,N_14088);
xnor U17008 (N_17008,N_14596,N_15560);
xor U17009 (N_17009,N_15365,N_14183);
nand U17010 (N_17010,N_15188,N_15558);
or U17011 (N_17011,N_15441,N_15244);
xor U17012 (N_17012,N_15490,N_14907);
and U17013 (N_17013,N_14033,N_14009);
or U17014 (N_17014,N_15352,N_15940);
and U17015 (N_17015,N_15046,N_14782);
and U17016 (N_17016,N_15679,N_14406);
nand U17017 (N_17017,N_15050,N_14291);
nor U17018 (N_17018,N_15777,N_14957);
or U17019 (N_17019,N_14613,N_14849);
nand U17020 (N_17020,N_14145,N_15786);
nand U17021 (N_17021,N_14187,N_14968);
and U17022 (N_17022,N_14576,N_15972);
nand U17023 (N_17023,N_15229,N_14752);
nor U17024 (N_17024,N_14946,N_15619);
nand U17025 (N_17025,N_14513,N_14052);
or U17026 (N_17026,N_15398,N_14964);
and U17027 (N_17027,N_14700,N_14835);
nand U17028 (N_17028,N_14038,N_15946);
nand U17029 (N_17029,N_14848,N_15656);
or U17030 (N_17030,N_15488,N_14171);
and U17031 (N_17031,N_14180,N_14035);
nor U17032 (N_17032,N_15481,N_14525);
and U17033 (N_17033,N_14324,N_15464);
and U17034 (N_17034,N_14940,N_14397);
nor U17035 (N_17035,N_15330,N_14643);
nand U17036 (N_17036,N_15966,N_14793);
or U17037 (N_17037,N_15819,N_14012);
xnor U17038 (N_17038,N_15552,N_14595);
nor U17039 (N_17039,N_15555,N_14466);
nand U17040 (N_17040,N_15483,N_14764);
nand U17041 (N_17041,N_14494,N_15966);
nand U17042 (N_17042,N_15393,N_15375);
nand U17043 (N_17043,N_14445,N_14295);
nand U17044 (N_17044,N_15040,N_14726);
nor U17045 (N_17045,N_14284,N_14040);
and U17046 (N_17046,N_15579,N_14305);
nor U17047 (N_17047,N_14454,N_15514);
nand U17048 (N_17048,N_14681,N_15308);
or U17049 (N_17049,N_14268,N_14026);
xnor U17050 (N_17050,N_14910,N_14926);
and U17051 (N_17051,N_14624,N_15604);
nand U17052 (N_17052,N_14827,N_14026);
or U17053 (N_17053,N_14315,N_14053);
nand U17054 (N_17054,N_14021,N_14906);
nor U17055 (N_17055,N_14900,N_15393);
nand U17056 (N_17056,N_15311,N_14137);
nor U17057 (N_17057,N_14915,N_14846);
or U17058 (N_17058,N_15661,N_15981);
or U17059 (N_17059,N_15214,N_15065);
xor U17060 (N_17060,N_15444,N_14767);
xor U17061 (N_17061,N_14623,N_15866);
or U17062 (N_17062,N_15252,N_14753);
nand U17063 (N_17063,N_15023,N_14711);
and U17064 (N_17064,N_15610,N_14472);
xor U17065 (N_17065,N_15472,N_15936);
nand U17066 (N_17066,N_15969,N_14983);
nand U17067 (N_17067,N_14535,N_14962);
and U17068 (N_17068,N_14303,N_14970);
or U17069 (N_17069,N_15257,N_15983);
and U17070 (N_17070,N_15340,N_14901);
nor U17071 (N_17071,N_14571,N_15899);
nand U17072 (N_17072,N_14781,N_14428);
nand U17073 (N_17073,N_15644,N_15342);
or U17074 (N_17074,N_14379,N_15487);
nor U17075 (N_17075,N_15726,N_14515);
nor U17076 (N_17076,N_14929,N_15492);
nor U17077 (N_17077,N_14569,N_15867);
nand U17078 (N_17078,N_15941,N_14433);
or U17079 (N_17079,N_15086,N_14555);
and U17080 (N_17080,N_14080,N_15267);
nor U17081 (N_17081,N_15994,N_15272);
and U17082 (N_17082,N_15052,N_15896);
or U17083 (N_17083,N_14964,N_15731);
or U17084 (N_17084,N_14954,N_14595);
or U17085 (N_17085,N_14494,N_15349);
and U17086 (N_17086,N_14243,N_14300);
nand U17087 (N_17087,N_15400,N_15697);
nand U17088 (N_17088,N_15237,N_14843);
nor U17089 (N_17089,N_15901,N_15817);
and U17090 (N_17090,N_14519,N_15204);
xor U17091 (N_17091,N_14385,N_15045);
and U17092 (N_17092,N_15372,N_15730);
or U17093 (N_17093,N_14733,N_15040);
and U17094 (N_17094,N_15141,N_15231);
xor U17095 (N_17095,N_14651,N_14702);
nor U17096 (N_17096,N_15714,N_15303);
nand U17097 (N_17097,N_14997,N_15400);
or U17098 (N_17098,N_14415,N_15583);
and U17099 (N_17099,N_14527,N_14534);
or U17100 (N_17100,N_14625,N_14976);
xor U17101 (N_17101,N_15101,N_15755);
nand U17102 (N_17102,N_15523,N_15529);
nor U17103 (N_17103,N_14372,N_15374);
or U17104 (N_17104,N_14601,N_14268);
or U17105 (N_17105,N_14756,N_14618);
and U17106 (N_17106,N_15421,N_14539);
nand U17107 (N_17107,N_15325,N_14482);
nand U17108 (N_17108,N_15882,N_14659);
and U17109 (N_17109,N_14654,N_15617);
or U17110 (N_17110,N_14912,N_14289);
nor U17111 (N_17111,N_14559,N_15305);
nand U17112 (N_17112,N_14560,N_14330);
nor U17113 (N_17113,N_14067,N_15606);
and U17114 (N_17114,N_14513,N_14528);
or U17115 (N_17115,N_14373,N_14999);
xor U17116 (N_17116,N_14021,N_14726);
nand U17117 (N_17117,N_14074,N_15050);
xor U17118 (N_17118,N_14368,N_14728);
or U17119 (N_17119,N_14014,N_15690);
xor U17120 (N_17120,N_14112,N_14391);
and U17121 (N_17121,N_14543,N_14021);
xor U17122 (N_17122,N_15386,N_15453);
and U17123 (N_17123,N_15043,N_15595);
nor U17124 (N_17124,N_15733,N_15553);
xor U17125 (N_17125,N_15632,N_14222);
and U17126 (N_17126,N_14383,N_15302);
nand U17127 (N_17127,N_15470,N_15762);
xor U17128 (N_17128,N_15885,N_15031);
nand U17129 (N_17129,N_15541,N_14653);
and U17130 (N_17130,N_15268,N_15687);
nand U17131 (N_17131,N_15770,N_15395);
xnor U17132 (N_17132,N_15816,N_15638);
nor U17133 (N_17133,N_14374,N_14219);
and U17134 (N_17134,N_14452,N_14050);
xor U17135 (N_17135,N_15673,N_14748);
nor U17136 (N_17136,N_14443,N_14491);
xor U17137 (N_17137,N_14898,N_15165);
xnor U17138 (N_17138,N_14145,N_15388);
or U17139 (N_17139,N_15238,N_14769);
nor U17140 (N_17140,N_14473,N_14927);
or U17141 (N_17141,N_14415,N_14281);
or U17142 (N_17142,N_15572,N_14586);
nand U17143 (N_17143,N_15899,N_14107);
or U17144 (N_17144,N_14528,N_15535);
and U17145 (N_17145,N_14715,N_14379);
or U17146 (N_17146,N_14655,N_14702);
nand U17147 (N_17147,N_14410,N_14371);
nor U17148 (N_17148,N_15775,N_14758);
nor U17149 (N_17149,N_14131,N_15724);
and U17150 (N_17150,N_14656,N_15674);
nor U17151 (N_17151,N_14124,N_15180);
xnor U17152 (N_17152,N_15987,N_15067);
nor U17153 (N_17153,N_14589,N_14408);
and U17154 (N_17154,N_14330,N_15507);
or U17155 (N_17155,N_14373,N_15450);
nand U17156 (N_17156,N_14691,N_15491);
nor U17157 (N_17157,N_14496,N_15481);
nand U17158 (N_17158,N_15128,N_14279);
or U17159 (N_17159,N_15792,N_14567);
or U17160 (N_17160,N_15783,N_15332);
xor U17161 (N_17161,N_15502,N_14422);
or U17162 (N_17162,N_15341,N_14133);
or U17163 (N_17163,N_14447,N_14278);
or U17164 (N_17164,N_14647,N_15180);
or U17165 (N_17165,N_15582,N_15652);
xnor U17166 (N_17166,N_15603,N_14328);
xor U17167 (N_17167,N_14918,N_15386);
or U17168 (N_17168,N_15764,N_14446);
nor U17169 (N_17169,N_15134,N_14427);
and U17170 (N_17170,N_14150,N_15132);
xnor U17171 (N_17171,N_15920,N_15987);
xnor U17172 (N_17172,N_14808,N_14235);
and U17173 (N_17173,N_15483,N_14822);
or U17174 (N_17174,N_14133,N_14633);
and U17175 (N_17175,N_15942,N_14246);
nor U17176 (N_17176,N_14612,N_15058);
or U17177 (N_17177,N_15862,N_14438);
nor U17178 (N_17178,N_15697,N_15722);
nor U17179 (N_17179,N_15885,N_15138);
xor U17180 (N_17180,N_15991,N_15087);
nor U17181 (N_17181,N_14116,N_15240);
or U17182 (N_17182,N_14612,N_15461);
nand U17183 (N_17183,N_15275,N_15003);
nand U17184 (N_17184,N_14504,N_14129);
nor U17185 (N_17185,N_14835,N_15024);
nor U17186 (N_17186,N_14505,N_14726);
xor U17187 (N_17187,N_14227,N_14794);
or U17188 (N_17188,N_14216,N_15550);
and U17189 (N_17189,N_15092,N_14407);
nor U17190 (N_17190,N_15411,N_15184);
or U17191 (N_17191,N_14957,N_15565);
nand U17192 (N_17192,N_14281,N_15892);
xnor U17193 (N_17193,N_15199,N_14745);
nand U17194 (N_17194,N_15462,N_14574);
nor U17195 (N_17195,N_14735,N_14645);
nor U17196 (N_17196,N_14784,N_14359);
nand U17197 (N_17197,N_14494,N_14903);
and U17198 (N_17198,N_14303,N_15519);
nand U17199 (N_17199,N_14434,N_15570);
and U17200 (N_17200,N_14778,N_14155);
or U17201 (N_17201,N_15066,N_14226);
nor U17202 (N_17202,N_15178,N_15842);
xor U17203 (N_17203,N_15693,N_14419);
or U17204 (N_17204,N_14430,N_14907);
or U17205 (N_17205,N_15278,N_15973);
or U17206 (N_17206,N_15985,N_14820);
and U17207 (N_17207,N_14556,N_14187);
nand U17208 (N_17208,N_15520,N_15052);
nor U17209 (N_17209,N_15803,N_14756);
nand U17210 (N_17210,N_15970,N_15901);
or U17211 (N_17211,N_14885,N_15467);
or U17212 (N_17212,N_15736,N_15518);
and U17213 (N_17213,N_14326,N_15587);
and U17214 (N_17214,N_15056,N_15772);
nor U17215 (N_17215,N_15850,N_15302);
nor U17216 (N_17216,N_14183,N_15106);
xor U17217 (N_17217,N_15675,N_14928);
or U17218 (N_17218,N_14263,N_14708);
or U17219 (N_17219,N_14647,N_14549);
nor U17220 (N_17220,N_14333,N_14816);
xnor U17221 (N_17221,N_14164,N_15445);
or U17222 (N_17222,N_15276,N_15785);
nand U17223 (N_17223,N_14444,N_14012);
or U17224 (N_17224,N_14583,N_14990);
xor U17225 (N_17225,N_15815,N_14539);
or U17226 (N_17226,N_14418,N_14145);
or U17227 (N_17227,N_14176,N_14833);
and U17228 (N_17228,N_14265,N_14893);
nor U17229 (N_17229,N_14592,N_14187);
or U17230 (N_17230,N_14038,N_14041);
nor U17231 (N_17231,N_14876,N_14007);
or U17232 (N_17232,N_14495,N_15703);
or U17233 (N_17233,N_14639,N_14599);
or U17234 (N_17234,N_15178,N_14464);
xnor U17235 (N_17235,N_15567,N_15915);
and U17236 (N_17236,N_14617,N_15292);
and U17237 (N_17237,N_14213,N_15315);
nor U17238 (N_17238,N_15382,N_15954);
nor U17239 (N_17239,N_15621,N_15328);
nand U17240 (N_17240,N_14662,N_14463);
and U17241 (N_17241,N_14204,N_15889);
nand U17242 (N_17242,N_15650,N_14605);
xor U17243 (N_17243,N_14622,N_14821);
or U17244 (N_17244,N_15091,N_15065);
nor U17245 (N_17245,N_14988,N_14206);
xor U17246 (N_17246,N_14960,N_14291);
and U17247 (N_17247,N_15456,N_14761);
nor U17248 (N_17248,N_14827,N_15931);
or U17249 (N_17249,N_15518,N_14597);
or U17250 (N_17250,N_14243,N_15076);
nor U17251 (N_17251,N_14261,N_14011);
nor U17252 (N_17252,N_14043,N_14997);
nor U17253 (N_17253,N_15435,N_15064);
and U17254 (N_17254,N_15235,N_14906);
or U17255 (N_17255,N_15242,N_15900);
and U17256 (N_17256,N_15611,N_15838);
and U17257 (N_17257,N_15708,N_14612);
nor U17258 (N_17258,N_15736,N_15640);
nor U17259 (N_17259,N_14902,N_14805);
xnor U17260 (N_17260,N_14146,N_15999);
nand U17261 (N_17261,N_14741,N_14202);
nor U17262 (N_17262,N_14483,N_15083);
nor U17263 (N_17263,N_14486,N_14223);
or U17264 (N_17264,N_14479,N_14613);
nor U17265 (N_17265,N_15143,N_15480);
xor U17266 (N_17266,N_14173,N_14267);
and U17267 (N_17267,N_14292,N_14385);
nand U17268 (N_17268,N_14379,N_14603);
or U17269 (N_17269,N_14135,N_14114);
nor U17270 (N_17270,N_14547,N_15954);
nand U17271 (N_17271,N_14725,N_15984);
and U17272 (N_17272,N_14320,N_15115);
nor U17273 (N_17273,N_15669,N_15917);
or U17274 (N_17274,N_15166,N_14332);
and U17275 (N_17275,N_14181,N_15751);
nand U17276 (N_17276,N_14414,N_14671);
nor U17277 (N_17277,N_15872,N_14326);
nand U17278 (N_17278,N_14520,N_15390);
and U17279 (N_17279,N_14119,N_14358);
nor U17280 (N_17280,N_15309,N_15731);
xnor U17281 (N_17281,N_15574,N_14402);
and U17282 (N_17282,N_14551,N_15766);
and U17283 (N_17283,N_15961,N_14303);
and U17284 (N_17284,N_14148,N_14419);
nor U17285 (N_17285,N_15772,N_14426);
and U17286 (N_17286,N_14898,N_14353);
and U17287 (N_17287,N_14735,N_14939);
xnor U17288 (N_17288,N_14085,N_15790);
and U17289 (N_17289,N_14019,N_15488);
and U17290 (N_17290,N_15871,N_14111);
nor U17291 (N_17291,N_14208,N_15899);
or U17292 (N_17292,N_14821,N_14222);
nor U17293 (N_17293,N_14122,N_15641);
and U17294 (N_17294,N_15712,N_14220);
and U17295 (N_17295,N_14848,N_14182);
or U17296 (N_17296,N_14568,N_14279);
nor U17297 (N_17297,N_14019,N_15662);
xnor U17298 (N_17298,N_15406,N_14359);
nor U17299 (N_17299,N_15779,N_14810);
nor U17300 (N_17300,N_15388,N_15530);
nor U17301 (N_17301,N_15974,N_15012);
and U17302 (N_17302,N_15739,N_14761);
or U17303 (N_17303,N_15001,N_15148);
nor U17304 (N_17304,N_15529,N_14769);
and U17305 (N_17305,N_15807,N_14346);
xor U17306 (N_17306,N_14808,N_15808);
xnor U17307 (N_17307,N_15681,N_14465);
nor U17308 (N_17308,N_15937,N_14450);
xor U17309 (N_17309,N_15057,N_14981);
and U17310 (N_17310,N_14405,N_15812);
nor U17311 (N_17311,N_15296,N_15500);
nor U17312 (N_17312,N_15689,N_15403);
and U17313 (N_17313,N_14579,N_14798);
or U17314 (N_17314,N_14769,N_15010);
and U17315 (N_17315,N_15577,N_15532);
nor U17316 (N_17316,N_15776,N_14296);
xor U17317 (N_17317,N_14096,N_14996);
and U17318 (N_17318,N_15797,N_14084);
nand U17319 (N_17319,N_15621,N_14104);
nand U17320 (N_17320,N_15017,N_14810);
nor U17321 (N_17321,N_14686,N_15379);
nand U17322 (N_17322,N_14908,N_15477);
nor U17323 (N_17323,N_15069,N_15236);
nand U17324 (N_17324,N_14222,N_15333);
and U17325 (N_17325,N_15377,N_14575);
or U17326 (N_17326,N_15381,N_15642);
xnor U17327 (N_17327,N_14443,N_14848);
nor U17328 (N_17328,N_15014,N_15982);
xor U17329 (N_17329,N_15398,N_15258);
xnor U17330 (N_17330,N_15416,N_14396);
nand U17331 (N_17331,N_15703,N_15662);
and U17332 (N_17332,N_14742,N_14417);
xnor U17333 (N_17333,N_15004,N_15027);
xnor U17334 (N_17334,N_15619,N_14765);
or U17335 (N_17335,N_14028,N_14154);
nor U17336 (N_17336,N_14899,N_14802);
nor U17337 (N_17337,N_15991,N_14911);
nor U17338 (N_17338,N_15052,N_14396);
xor U17339 (N_17339,N_15641,N_15438);
or U17340 (N_17340,N_15896,N_14676);
or U17341 (N_17341,N_14855,N_15575);
or U17342 (N_17342,N_14623,N_15293);
or U17343 (N_17343,N_15253,N_15919);
nor U17344 (N_17344,N_14439,N_14284);
or U17345 (N_17345,N_15828,N_15891);
xnor U17346 (N_17346,N_15402,N_15123);
nor U17347 (N_17347,N_15765,N_14354);
nor U17348 (N_17348,N_15447,N_15497);
or U17349 (N_17349,N_14807,N_14532);
nand U17350 (N_17350,N_14908,N_14508);
nand U17351 (N_17351,N_14484,N_15821);
xnor U17352 (N_17352,N_14863,N_14895);
nor U17353 (N_17353,N_14806,N_15753);
and U17354 (N_17354,N_14299,N_14115);
and U17355 (N_17355,N_14429,N_14887);
nor U17356 (N_17356,N_15576,N_15936);
xnor U17357 (N_17357,N_15939,N_15569);
and U17358 (N_17358,N_15970,N_15529);
nor U17359 (N_17359,N_14332,N_14720);
nor U17360 (N_17360,N_15803,N_15096);
xor U17361 (N_17361,N_15051,N_14365);
nand U17362 (N_17362,N_15722,N_15211);
and U17363 (N_17363,N_14496,N_14471);
nor U17364 (N_17364,N_14474,N_15510);
nand U17365 (N_17365,N_15174,N_15857);
nor U17366 (N_17366,N_14115,N_15023);
nand U17367 (N_17367,N_14436,N_15363);
nor U17368 (N_17368,N_14932,N_15785);
and U17369 (N_17369,N_15684,N_14877);
and U17370 (N_17370,N_15132,N_15615);
nand U17371 (N_17371,N_14743,N_15277);
nor U17372 (N_17372,N_14713,N_15276);
or U17373 (N_17373,N_15301,N_14554);
xor U17374 (N_17374,N_15773,N_15420);
and U17375 (N_17375,N_14766,N_15846);
nor U17376 (N_17376,N_14056,N_14294);
nor U17377 (N_17377,N_14486,N_14502);
or U17378 (N_17378,N_14401,N_14023);
and U17379 (N_17379,N_15026,N_14793);
and U17380 (N_17380,N_15524,N_15243);
or U17381 (N_17381,N_14884,N_14123);
nand U17382 (N_17382,N_15261,N_15324);
nand U17383 (N_17383,N_14777,N_15090);
xnor U17384 (N_17384,N_15009,N_15511);
nor U17385 (N_17385,N_14432,N_15717);
xnor U17386 (N_17386,N_15072,N_14360);
or U17387 (N_17387,N_15858,N_14258);
xnor U17388 (N_17388,N_15385,N_14555);
nand U17389 (N_17389,N_15215,N_15222);
or U17390 (N_17390,N_14876,N_14850);
and U17391 (N_17391,N_15830,N_14839);
nor U17392 (N_17392,N_15451,N_14430);
nor U17393 (N_17393,N_15690,N_15323);
nand U17394 (N_17394,N_15003,N_14315);
nand U17395 (N_17395,N_14166,N_14316);
xnor U17396 (N_17396,N_14094,N_15281);
or U17397 (N_17397,N_14446,N_14557);
nor U17398 (N_17398,N_15276,N_15923);
nand U17399 (N_17399,N_15180,N_14272);
xnor U17400 (N_17400,N_14930,N_14444);
or U17401 (N_17401,N_14609,N_14631);
and U17402 (N_17402,N_15475,N_14469);
or U17403 (N_17403,N_15450,N_14832);
or U17404 (N_17404,N_14352,N_15078);
nand U17405 (N_17405,N_14065,N_15838);
nor U17406 (N_17406,N_15557,N_15068);
xnor U17407 (N_17407,N_14877,N_14834);
nor U17408 (N_17408,N_14541,N_14096);
nor U17409 (N_17409,N_15316,N_14012);
nor U17410 (N_17410,N_14432,N_14545);
or U17411 (N_17411,N_15865,N_14728);
and U17412 (N_17412,N_15774,N_15985);
nor U17413 (N_17413,N_15995,N_15460);
xnor U17414 (N_17414,N_15380,N_14755);
xor U17415 (N_17415,N_14985,N_14884);
or U17416 (N_17416,N_15394,N_15858);
and U17417 (N_17417,N_14300,N_14552);
and U17418 (N_17418,N_14479,N_15175);
nand U17419 (N_17419,N_14608,N_15881);
and U17420 (N_17420,N_15565,N_15641);
xnor U17421 (N_17421,N_14972,N_14789);
xnor U17422 (N_17422,N_14372,N_15096);
or U17423 (N_17423,N_14831,N_15894);
or U17424 (N_17424,N_14910,N_15133);
xor U17425 (N_17425,N_15842,N_14417);
xnor U17426 (N_17426,N_14255,N_15157);
xor U17427 (N_17427,N_14801,N_15845);
nor U17428 (N_17428,N_15275,N_14608);
nand U17429 (N_17429,N_15874,N_15663);
xor U17430 (N_17430,N_15331,N_14399);
nor U17431 (N_17431,N_15243,N_15133);
xor U17432 (N_17432,N_14280,N_14011);
and U17433 (N_17433,N_14015,N_14334);
nand U17434 (N_17434,N_15786,N_14613);
xor U17435 (N_17435,N_14554,N_14348);
and U17436 (N_17436,N_15806,N_15653);
nor U17437 (N_17437,N_14044,N_15033);
xnor U17438 (N_17438,N_14519,N_15563);
or U17439 (N_17439,N_14536,N_14925);
nand U17440 (N_17440,N_15157,N_14619);
xor U17441 (N_17441,N_14105,N_15402);
xor U17442 (N_17442,N_15530,N_14664);
nand U17443 (N_17443,N_14492,N_15288);
nor U17444 (N_17444,N_15351,N_14365);
nand U17445 (N_17445,N_14599,N_15678);
nor U17446 (N_17446,N_14654,N_15930);
nand U17447 (N_17447,N_15249,N_14393);
and U17448 (N_17448,N_14778,N_14168);
or U17449 (N_17449,N_14456,N_14277);
xor U17450 (N_17450,N_14508,N_15685);
xnor U17451 (N_17451,N_15591,N_14538);
and U17452 (N_17452,N_14740,N_15914);
nand U17453 (N_17453,N_15972,N_15742);
nor U17454 (N_17454,N_15808,N_14668);
nand U17455 (N_17455,N_15063,N_15410);
or U17456 (N_17456,N_15465,N_15187);
nand U17457 (N_17457,N_15831,N_14356);
and U17458 (N_17458,N_15059,N_14794);
or U17459 (N_17459,N_15776,N_14084);
or U17460 (N_17460,N_15292,N_15843);
nor U17461 (N_17461,N_14388,N_15442);
xor U17462 (N_17462,N_15190,N_15275);
xor U17463 (N_17463,N_14579,N_15925);
nor U17464 (N_17464,N_15930,N_15892);
nand U17465 (N_17465,N_14536,N_14451);
and U17466 (N_17466,N_14348,N_15651);
or U17467 (N_17467,N_15672,N_15073);
or U17468 (N_17468,N_15652,N_14569);
xnor U17469 (N_17469,N_15461,N_15876);
nand U17470 (N_17470,N_15656,N_15907);
nor U17471 (N_17471,N_15660,N_14299);
nand U17472 (N_17472,N_14551,N_15318);
or U17473 (N_17473,N_15061,N_15475);
or U17474 (N_17474,N_14072,N_15777);
or U17475 (N_17475,N_14798,N_14402);
xnor U17476 (N_17476,N_15933,N_14978);
nor U17477 (N_17477,N_14876,N_14128);
or U17478 (N_17478,N_14775,N_14631);
or U17479 (N_17479,N_15344,N_15414);
xor U17480 (N_17480,N_15983,N_14688);
or U17481 (N_17481,N_14670,N_14122);
or U17482 (N_17482,N_14414,N_14136);
nor U17483 (N_17483,N_14098,N_14790);
and U17484 (N_17484,N_14294,N_14369);
or U17485 (N_17485,N_15670,N_14408);
xnor U17486 (N_17486,N_14561,N_15679);
nand U17487 (N_17487,N_14332,N_14127);
and U17488 (N_17488,N_14185,N_14558);
or U17489 (N_17489,N_14143,N_14110);
nor U17490 (N_17490,N_15214,N_15386);
nand U17491 (N_17491,N_15025,N_14638);
or U17492 (N_17492,N_14399,N_14591);
nand U17493 (N_17493,N_15340,N_15415);
or U17494 (N_17494,N_15990,N_15022);
nand U17495 (N_17495,N_15448,N_14045);
xnor U17496 (N_17496,N_15348,N_14341);
and U17497 (N_17497,N_14919,N_14713);
and U17498 (N_17498,N_14363,N_15786);
xnor U17499 (N_17499,N_14269,N_15230);
nand U17500 (N_17500,N_15604,N_15100);
nor U17501 (N_17501,N_14216,N_15755);
or U17502 (N_17502,N_14122,N_15929);
nor U17503 (N_17503,N_14954,N_14468);
and U17504 (N_17504,N_15432,N_15756);
or U17505 (N_17505,N_14632,N_14421);
and U17506 (N_17506,N_14362,N_14056);
and U17507 (N_17507,N_15453,N_15342);
nand U17508 (N_17508,N_15985,N_15619);
xor U17509 (N_17509,N_14132,N_14241);
or U17510 (N_17510,N_15277,N_15128);
xnor U17511 (N_17511,N_15558,N_14968);
xnor U17512 (N_17512,N_15318,N_15421);
xnor U17513 (N_17513,N_14780,N_14437);
and U17514 (N_17514,N_14578,N_15255);
nor U17515 (N_17515,N_14251,N_14085);
nand U17516 (N_17516,N_15330,N_15678);
xnor U17517 (N_17517,N_14593,N_15682);
nand U17518 (N_17518,N_14251,N_14747);
and U17519 (N_17519,N_15090,N_15879);
or U17520 (N_17520,N_14324,N_15434);
and U17521 (N_17521,N_14705,N_15941);
and U17522 (N_17522,N_15979,N_14967);
nor U17523 (N_17523,N_15226,N_14461);
and U17524 (N_17524,N_14829,N_14231);
or U17525 (N_17525,N_15947,N_15359);
xnor U17526 (N_17526,N_14117,N_14490);
xor U17527 (N_17527,N_15696,N_14011);
or U17528 (N_17528,N_15174,N_15186);
nand U17529 (N_17529,N_14273,N_15181);
and U17530 (N_17530,N_15476,N_15024);
xnor U17531 (N_17531,N_14987,N_14127);
nand U17532 (N_17532,N_15728,N_15692);
nor U17533 (N_17533,N_15443,N_14914);
xnor U17534 (N_17534,N_14575,N_14824);
xnor U17535 (N_17535,N_15045,N_15846);
and U17536 (N_17536,N_14835,N_14850);
or U17537 (N_17537,N_14861,N_14630);
nor U17538 (N_17538,N_15316,N_14370);
or U17539 (N_17539,N_14653,N_15044);
nand U17540 (N_17540,N_15837,N_15481);
xor U17541 (N_17541,N_14874,N_15688);
nor U17542 (N_17542,N_15381,N_15324);
nor U17543 (N_17543,N_15519,N_15021);
nand U17544 (N_17544,N_14013,N_14141);
or U17545 (N_17545,N_14233,N_14572);
or U17546 (N_17546,N_15265,N_14805);
nor U17547 (N_17547,N_15810,N_15826);
or U17548 (N_17548,N_14597,N_14434);
and U17549 (N_17549,N_15682,N_14421);
and U17550 (N_17550,N_14556,N_14600);
or U17551 (N_17551,N_15961,N_14848);
nand U17552 (N_17552,N_14086,N_14296);
or U17553 (N_17553,N_15130,N_15529);
or U17554 (N_17554,N_14223,N_14999);
nand U17555 (N_17555,N_14655,N_14470);
xnor U17556 (N_17556,N_15731,N_15184);
or U17557 (N_17557,N_14673,N_15194);
xor U17558 (N_17558,N_15809,N_14877);
nor U17559 (N_17559,N_15905,N_15671);
and U17560 (N_17560,N_14151,N_15820);
and U17561 (N_17561,N_15677,N_14450);
xor U17562 (N_17562,N_14892,N_15990);
nor U17563 (N_17563,N_15156,N_15916);
and U17564 (N_17564,N_15023,N_14375);
and U17565 (N_17565,N_15045,N_15983);
nand U17566 (N_17566,N_14887,N_15488);
nor U17567 (N_17567,N_14786,N_14008);
nor U17568 (N_17568,N_14178,N_15553);
xnor U17569 (N_17569,N_14850,N_15391);
and U17570 (N_17570,N_15615,N_15254);
nand U17571 (N_17571,N_15923,N_15006);
nor U17572 (N_17572,N_15978,N_15958);
and U17573 (N_17573,N_14169,N_15824);
nor U17574 (N_17574,N_14002,N_15901);
or U17575 (N_17575,N_14819,N_14024);
or U17576 (N_17576,N_14787,N_14898);
nor U17577 (N_17577,N_15760,N_15113);
nand U17578 (N_17578,N_15316,N_15757);
nand U17579 (N_17579,N_15340,N_15226);
nor U17580 (N_17580,N_14590,N_14685);
or U17581 (N_17581,N_15530,N_15938);
or U17582 (N_17582,N_14687,N_15011);
and U17583 (N_17583,N_14627,N_15585);
nand U17584 (N_17584,N_15262,N_14174);
nand U17585 (N_17585,N_14238,N_14581);
or U17586 (N_17586,N_15048,N_14195);
nor U17587 (N_17587,N_15874,N_14300);
nand U17588 (N_17588,N_15428,N_15217);
and U17589 (N_17589,N_15581,N_14675);
nand U17590 (N_17590,N_14220,N_14948);
xnor U17591 (N_17591,N_14202,N_14696);
and U17592 (N_17592,N_15078,N_14468);
nor U17593 (N_17593,N_15309,N_14096);
xor U17594 (N_17594,N_15262,N_15779);
xnor U17595 (N_17595,N_14236,N_15798);
or U17596 (N_17596,N_14600,N_14804);
or U17597 (N_17597,N_15087,N_14088);
nand U17598 (N_17598,N_14069,N_15618);
and U17599 (N_17599,N_15936,N_14200);
xnor U17600 (N_17600,N_14315,N_15352);
nand U17601 (N_17601,N_14260,N_14196);
xnor U17602 (N_17602,N_14798,N_15115);
and U17603 (N_17603,N_14206,N_14942);
xor U17604 (N_17604,N_14451,N_14495);
and U17605 (N_17605,N_14767,N_14505);
nand U17606 (N_17606,N_15683,N_15610);
and U17607 (N_17607,N_14482,N_15938);
and U17608 (N_17608,N_14061,N_14634);
xor U17609 (N_17609,N_14069,N_14495);
or U17610 (N_17610,N_15678,N_14403);
nor U17611 (N_17611,N_14547,N_14712);
nor U17612 (N_17612,N_15138,N_14788);
xnor U17613 (N_17613,N_14442,N_15685);
nand U17614 (N_17614,N_14718,N_14424);
xnor U17615 (N_17615,N_15496,N_15769);
or U17616 (N_17616,N_15919,N_15244);
or U17617 (N_17617,N_15118,N_14550);
and U17618 (N_17618,N_14929,N_15859);
nand U17619 (N_17619,N_15422,N_14961);
nor U17620 (N_17620,N_15286,N_15672);
nand U17621 (N_17621,N_14217,N_15540);
and U17622 (N_17622,N_15663,N_15591);
nor U17623 (N_17623,N_14215,N_14231);
or U17624 (N_17624,N_14376,N_14286);
nor U17625 (N_17625,N_15624,N_14621);
and U17626 (N_17626,N_14023,N_15950);
nand U17627 (N_17627,N_14369,N_15721);
nand U17628 (N_17628,N_14871,N_14720);
nor U17629 (N_17629,N_15605,N_15560);
xnor U17630 (N_17630,N_15472,N_15817);
nand U17631 (N_17631,N_15215,N_14440);
or U17632 (N_17632,N_14315,N_14917);
or U17633 (N_17633,N_14975,N_14741);
nand U17634 (N_17634,N_14642,N_14643);
or U17635 (N_17635,N_15416,N_15478);
or U17636 (N_17636,N_14460,N_15591);
xnor U17637 (N_17637,N_15580,N_15159);
nor U17638 (N_17638,N_14768,N_15554);
and U17639 (N_17639,N_15893,N_15045);
and U17640 (N_17640,N_14066,N_14728);
nor U17641 (N_17641,N_15014,N_14038);
nor U17642 (N_17642,N_15285,N_15531);
nand U17643 (N_17643,N_15861,N_14942);
nand U17644 (N_17644,N_15471,N_14935);
and U17645 (N_17645,N_15500,N_15557);
xor U17646 (N_17646,N_15201,N_14562);
nor U17647 (N_17647,N_15713,N_15183);
or U17648 (N_17648,N_14412,N_15485);
nand U17649 (N_17649,N_14298,N_15080);
and U17650 (N_17650,N_14046,N_14262);
or U17651 (N_17651,N_14516,N_15457);
xor U17652 (N_17652,N_14746,N_14871);
and U17653 (N_17653,N_14682,N_15568);
nand U17654 (N_17654,N_15177,N_15368);
or U17655 (N_17655,N_14316,N_15536);
or U17656 (N_17656,N_15871,N_14373);
nand U17657 (N_17657,N_15134,N_15512);
and U17658 (N_17658,N_15151,N_15898);
nor U17659 (N_17659,N_14430,N_14666);
and U17660 (N_17660,N_14232,N_15508);
nor U17661 (N_17661,N_14454,N_14282);
nor U17662 (N_17662,N_15066,N_14264);
or U17663 (N_17663,N_15409,N_14043);
xnor U17664 (N_17664,N_14781,N_14329);
xor U17665 (N_17665,N_15513,N_14139);
or U17666 (N_17666,N_14250,N_14720);
nor U17667 (N_17667,N_15312,N_14295);
xnor U17668 (N_17668,N_15098,N_14173);
or U17669 (N_17669,N_14962,N_15859);
nor U17670 (N_17670,N_15168,N_14082);
and U17671 (N_17671,N_14878,N_14309);
or U17672 (N_17672,N_14015,N_14711);
xor U17673 (N_17673,N_14635,N_14147);
nand U17674 (N_17674,N_14851,N_15029);
or U17675 (N_17675,N_14862,N_14536);
or U17676 (N_17676,N_15285,N_15079);
and U17677 (N_17677,N_14016,N_14576);
or U17678 (N_17678,N_14983,N_14219);
xnor U17679 (N_17679,N_15714,N_14309);
or U17680 (N_17680,N_15632,N_15918);
xor U17681 (N_17681,N_14658,N_14269);
nor U17682 (N_17682,N_15167,N_15137);
or U17683 (N_17683,N_15321,N_15266);
and U17684 (N_17684,N_14608,N_14080);
and U17685 (N_17685,N_14309,N_14694);
nor U17686 (N_17686,N_14029,N_15059);
nand U17687 (N_17687,N_14291,N_15789);
or U17688 (N_17688,N_15479,N_15835);
and U17689 (N_17689,N_14298,N_14488);
nor U17690 (N_17690,N_14837,N_14513);
and U17691 (N_17691,N_14022,N_15770);
nand U17692 (N_17692,N_15967,N_15189);
and U17693 (N_17693,N_15292,N_15166);
nand U17694 (N_17694,N_14563,N_15142);
xor U17695 (N_17695,N_15389,N_14392);
xor U17696 (N_17696,N_15291,N_14987);
xnor U17697 (N_17697,N_14137,N_15205);
or U17698 (N_17698,N_15179,N_14778);
nand U17699 (N_17699,N_14745,N_15017);
xor U17700 (N_17700,N_14650,N_15880);
and U17701 (N_17701,N_15609,N_15135);
nand U17702 (N_17702,N_15049,N_14347);
nand U17703 (N_17703,N_14906,N_14048);
xnor U17704 (N_17704,N_15588,N_15356);
xnor U17705 (N_17705,N_14315,N_15983);
nand U17706 (N_17706,N_15080,N_15633);
and U17707 (N_17707,N_15795,N_14581);
and U17708 (N_17708,N_15845,N_14864);
xnor U17709 (N_17709,N_14243,N_14891);
xor U17710 (N_17710,N_15473,N_15756);
nand U17711 (N_17711,N_15727,N_14119);
nor U17712 (N_17712,N_15137,N_14309);
nor U17713 (N_17713,N_14578,N_15295);
and U17714 (N_17714,N_15293,N_15740);
nand U17715 (N_17715,N_14205,N_14626);
nor U17716 (N_17716,N_15457,N_15370);
or U17717 (N_17717,N_14859,N_15050);
nor U17718 (N_17718,N_15636,N_15315);
nand U17719 (N_17719,N_14772,N_15973);
xnor U17720 (N_17720,N_15393,N_15022);
and U17721 (N_17721,N_14827,N_15664);
or U17722 (N_17722,N_14447,N_15746);
nand U17723 (N_17723,N_14649,N_14895);
or U17724 (N_17724,N_14653,N_15939);
and U17725 (N_17725,N_14659,N_14446);
and U17726 (N_17726,N_15952,N_14051);
and U17727 (N_17727,N_15648,N_15471);
or U17728 (N_17728,N_15393,N_14091);
or U17729 (N_17729,N_15338,N_15175);
nand U17730 (N_17730,N_14494,N_14462);
or U17731 (N_17731,N_14570,N_14567);
xnor U17732 (N_17732,N_14270,N_15083);
nor U17733 (N_17733,N_14373,N_14816);
nor U17734 (N_17734,N_14927,N_15860);
and U17735 (N_17735,N_15121,N_14588);
nor U17736 (N_17736,N_15230,N_15585);
nand U17737 (N_17737,N_14552,N_15466);
and U17738 (N_17738,N_14326,N_14865);
and U17739 (N_17739,N_14563,N_14564);
and U17740 (N_17740,N_15985,N_15450);
and U17741 (N_17741,N_14688,N_14238);
or U17742 (N_17742,N_15505,N_14324);
nand U17743 (N_17743,N_14736,N_15821);
or U17744 (N_17744,N_14383,N_15689);
nand U17745 (N_17745,N_15125,N_14692);
nand U17746 (N_17746,N_14102,N_14304);
xor U17747 (N_17747,N_15172,N_15068);
or U17748 (N_17748,N_14563,N_14294);
and U17749 (N_17749,N_15062,N_14545);
and U17750 (N_17750,N_14886,N_14180);
and U17751 (N_17751,N_14307,N_14110);
nand U17752 (N_17752,N_14230,N_15883);
or U17753 (N_17753,N_15542,N_14186);
nor U17754 (N_17754,N_15950,N_14918);
nand U17755 (N_17755,N_14494,N_15516);
nand U17756 (N_17756,N_14834,N_14684);
nand U17757 (N_17757,N_14931,N_14199);
or U17758 (N_17758,N_15721,N_14163);
nand U17759 (N_17759,N_15918,N_14515);
or U17760 (N_17760,N_15408,N_15710);
or U17761 (N_17761,N_15855,N_15457);
nor U17762 (N_17762,N_15695,N_14305);
nor U17763 (N_17763,N_14401,N_15223);
nor U17764 (N_17764,N_14598,N_15467);
nor U17765 (N_17765,N_15384,N_15490);
and U17766 (N_17766,N_14384,N_15877);
xor U17767 (N_17767,N_15242,N_15544);
and U17768 (N_17768,N_15691,N_15522);
nor U17769 (N_17769,N_14780,N_14961);
or U17770 (N_17770,N_14915,N_14132);
xor U17771 (N_17771,N_14711,N_14870);
nand U17772 (N_17772,N_14001,N_15548);
and U17773 (N_17773,N_15968,N_14986);
nor U17774 (N_17774,N_15201,N_14473);
or U17775 (N_17775,N_15787,N_14030);
nor U17776 (N_17776,N_15277,N_15889);
xnor U17777 (N_17777,N_14843,N_15394);
nand U17778 (N_17778,N_15654,N_15254);
nand U17779 (N_17779,N_14437,N_14078);
nor U17780 (N_17780,N_14511,N_14235);
and U17781 (N_17781,N_15794,N_14760);
or U17782 (N_17782,N_15463,N_15609);
nor U17783 (N_17783,N_14717,N_14548);
nor U17784 (N_17784,N_14173,N_14739);
nand U17785 (N_17785,N_15478,N_15729);
nor U17786 (N_17786,N_14132,N_14420);
or U17787 (N_17787,N_14017,N_15221);
nand U17788 (N_17788,N_14652,N_14473);
nand U17789 (N_17789,N_14452,N_14924);
or U17790 (N_17790,N_14805,N_15052);
or U17791 (N_17791,N_15450,N_15574);
and U17792 (N_17792,N_15707,N_15756);
or U17793 (N_17793,N_15505,N_15416);
nor U17794 (N_17794,N_14377,N_15393);
or U17795 (N_17795,N_14779,N_15384);
or U17796 (N_17796,N_14343,N_14647);
nand U17797 (N_17797,N_14567,N_15498);
or U17798 (N_17798,N_15822,N_15560);
or U17799 (N_17799,N_14816,N_14330);
xnor U17800 (N_17800,N_15244,N_14195);
and U17801 (N_17801,N_15067,N_15689);
and U17802 (N_17802,N_15021,N_14839);
xor U17803 (N_17803,N_15910,N_14938);
and U17804 (N_17804,N_15284,N_14245);
or U17805 (N_17805,N_14319,N_14143);
or U17806 (N_17806,N_14969,N_15434);
xnor U17807 (N_17807,N_14550,N_14468);
or U17808 (N_17808,N_14854,N_15548);
xnor U17809 (N_17809,N_15077,N_15750);
nand U17810 (N_17810,N_15629,N_15425);
and U17811 (N_17811,N_15940,N_14105);
nor U17812 (N_17812,N_14490,N_15026);
or U17813 (N_17813,N_15751,N_15069);
nor U17814 (N_17814,N_15810,N_14404);
and U17815 (N_17815,N_14835,N_14792);
xor U17816 (N_17816,N_14524,N_14638);
and U17817 (N_17817,N_14707,N_15114);
nor U17818 (N_17818,N_15566,N_15654);
and U17819 (N_17819,N_15476,N_15153);
and U17820 (N_17820,N_15699,N_14481);
and U17821 (N_17821,N_14018,N_15277);
and U17822 (N_17822,N_14485,N_15451);
nor U17823 (N_17823,N_14476,N_15460);
or U17824 (N_17824,N_15631,N_14952);
xor U17825 (N_17825,N_14274,N_15914);
or U17826 (N_17826,N_15921,N_14596);
or U17827 (N_17827,N_14822,N_14378);
nor U17828 (N_17828,N_14438,N_15037);
nand U17829 (N_17829,N_15076,N_15526);
nand U17830 (N_17830,N_14146,N_15869);
nor U17831 (N_17831,N_14157,N_15676);
nand U17832 (N_17832,N_15761,N_15969);
nor U17833 (N_17833,N_15333,N_14312);
nand U17834 (N_17834,N_15818,N_14294);
or U17835 (N_17835,N_15611,N_14722);
and U17836 (N_17836,N_15943,N_15696);
or U17837 (N_17837,N_14404,N_15076);
or U17838 (N_17838,N_14169,N_15349);
and U17839 (N_17839,N_15218,N_15795);
xor U17840 (N_17840,N_14639,N_14984);
nand U17841 (N_17841,N_14776,N_14629);
and U17842 (N_17842,N_14479,N_15506);
nor U17843 (N_17843,N_15186,N_14103);
xor U17844 (N_17844,N_15708,N_15047);
and U17845 (N_17845,N_15513,N_15136);
or U17846 (N_17846,N_14253,N_15619);
xor U17847 (N_17847,N_15032,N_14424);
and U17848 (N_17848,N_15402,N_14700);
nand U17849 (N_17849,N_14088,N_14948);
nor U17850 (N_17850,N_14539,N_14216);
nor U17851 (N_17851,N_15237,N_15431);
xnor U17852 (N_17852,N_15793,N_15252);
nor U17853 (N_17853,N_15921,N_14768);
and U17854 (N_17854,N_15741,N_15765);
or U17855 (N_17855,N_15898,N_15630);
nor U17856 (N_17856,N_14678,N_15946);
nor U17857 (N_17857,N_14377,N_15718);
xor U17858 (N_17858,N_14474,N_15886);
and U17859 (N_17859,N_14433,N_14840);
or U17860 (N_17860,N_14589,N_14403);
and U17861 (N_17861,N_14428,N_14208);
and U17862 (N_17862,N_14590,N_14588);
and U17863 (N_17863,N_14328,N_15414);
xor U17864 (N_17864,N_15323,N_14566);
and U17865 (N_17865,N_14985,N_14987);
and U17866 (N_17866,N_14427,N_15332);
and U17867 (N_17867,N_14660,N_14054);
and U17868 (N_17868,N_15503,N_15682);
and U17869 (N_17869,N_15421,N_15935);
and U17870 (N_17870,N_15128,N_14139);
or U17871 (N_17871,N_15278,N_15047);
and U17872 (N_17872,N_15756,N_15484);
and U17873 (N_17873,N_14792,N_15230);
nand U17874 (N_17874,N_15057,N_15282);
nor U17875 (N_17875,N_15910,N_15343);
or U17876 (N_17876,N_15403,N_14826);
or U17877 (N_17877,N_15190,N_15309);
and U17878 (N_17878,N_14633,N_15931);
or U17879 (N_17879,N_15964,N_15435);
nor U17880 (N_17880,N_15650,N_14842);
and U17881 (N_17881,N_14781,N_15870);
nor U17882 (N_17882,N_14361,N_15995);
nand U17883 (N_17883,N_14320,N_14821);
nand U17884 (N_17884,N_15397,N_14909);
nand U17885 (N_17885,N_14110,N_15670);
and U17886 (N_17886,N_14108,N_14832);
and U17887 (N_17887,N_14049,N_14610);
and U17888 (N_17888,N_15478,N_14383);
and U17889 (N_17889,N_15879,N_14801);
and U17890 (N_17890,N_14860,N_14788);
or U17891 (N_17891,N_14020,N_15304);
nand U17892 (N_17892,N_15841,N_14372);
nand U17893 (N_17893,N_15422,N_15334);
or U17894 (N_17894,N_14702,N_14411);
and U17895 (N_17895,N_15124,N_14232);
or U17896 (N_17896,N_14241,N_14929);
nor U17897 (N_17897,N_15269,N_14196);
nand U17898 (N_17898,N_15467,N_14992);
or U17899 (N_17899,N_14173,N_14889);
or U17900 (N_17900,N_14652,N_15007);
nand U17901 (N_17901,N_15534,N_14513);
nor U17902 (N_17902,N_15903,N_15490);
xnor U17903 (N_17903,N_14696,N_14738);
or U17904 (N_17904,N_14455,N_15982);
and U17905 (N_17905,N_15414,N_14332);
nand U17906 (N_17906,N_15663,N_14342);
or U17907 (N_17907,N_15689,N_14972);
nand U17908 (N_17908,N_15431,N_14975);
xor U17909 (N_17909,N_15107,N_14864);
xnor U17910 (N_17910,N_14258,N_15172);
and U17911 (N_17911,N_14157,N_15048);
or U17912 (N_17912,N_15330,N_15066);
xor U17913 (N_17913,N_15262,N_14078);
xor U17914 (N_17914,N_14702,N_14065);
nor U17915 (N_17915,N_15759,N_14381);
nand U17916 (N_17916,N_15574,N_14761);
nand U17917 (N_17917,N_14351,N_15352);
nor U17918 (N_17918,N_14047,N_14630);
nand U17919 (N_17919,N_15633,N_15386);
nand U17920 (N_17920,N_15907,N_14234);
nand U17921 (N_17921,N_15090,N_14362);
xnor U17922 (N_17922,N_15045,N_14268);
and U17923 (N_17923,N_14057,N_15815);
nand U17924 (N_17924,N_15482,N_14869);
nand U17925 (N_17925,N_14230,N_15071);
nand U17926 (N_17926,N_14431,N_15020);
nand U17927 (N_17927,N_14720,N_15269);
or U17928 (N_17928,N_14836,N_14206);
and U17929 (N_17929,N_14911,N_15234);
or U17930 (N_17930,N_15682,N_14728);
nor U17931 (N_17931,N_15982,N_14181);
or U17932 (N_17932,N_15516,N_15721);
and U17933 (N_17933,N_15818,N_14402);
or U17934 (N_17934,N_15369,N_14618);
or U17935 (N_17935,N_15075,N_14728);
xnor U17936 (N_17936,N_15606,N_15173);
xor U17937 (N_17937,N_15574,N_15776);
and U17938 (N_17938,N_15682,N_14829);
xnor U17939 (N_17939,N_15930,N_15216);
or U17940 (N_17940,N_14842,N_15305);
and U17941 (N_17941,N_14141,N_14417);
or U17942 (N_17942,N_15738,N_15669);
or U17943 (N_17943,N_15549,N_15052);
nor U17944 (N_17944,N_15824,N_14306);
nor U17945 (N_17945,N_14065,N_14024);
nor U17946 (N_17946,N_15613,N_15791);
xor U17947 (N_17947,N_15201,N_15514);
xnor U17948 (N_17948,N_14145,N_15278);
nor U17949 (N_17949,N_15630,N_14562);
nand U17950 (N_17950,N_15466,N_15620);
nand U17951 (N_17951,N_14054,N_15660);
or U17952 (N_17952,N_14896,N_15186);
and U17953 (N_17953,N_15640,N_14141);
xor U17954 (N_17954,N_14934,N_15496);
or U17955 (N_17955,N_14481,N_14402);
or U17956 (N_17956,N_15833,N_14662);
nand U17957 (N_17957,N_14813,N_15135);
xor U17958 (N_17958,N_14610,N_15602);
and U17959 (N_17959,N_14114,N_15458);
xor U17960 (N_17960,N_15830,N_15784);
and U17961 (N_17961,N_14949,N_15883);
and U17962 (N_17962,N_15161,N_14551);
and U17963 (N_17963,N_14551,N_15706);
nand U17964 (N_17964,N_14463,N_14842);
xor U17965 (N_17965,N_14061,N_14870);
xor U17966 (N_17966,N_14839,N_14642);
and U17967 (N_17967,N_15730,N_15471);
and U17968 (N_17968,N_15986,N_14620);
nand U17969 (N_17969,N_14475,N_14314);
xnor U17970 (N_17970,N_15785,N_14639);
nor U17971 (N_17971,N_14222,N_15120);
nor U17972 (N_17972,N_15922,N_14670);
or U17973 (N_17973,N_15628,N_14639);
xor U17974 (N_17974,N_14353,N_15946);
or U17975 (N_17975,N_15734,N_14801);
or U17976 (N_17976,N_14374,N_14630);
nor U17977 (N_17977,N_14977,N_14049);
and U17978 (N_17978,N_15196,N_15634);
nor U17979 (N_17979,N_14062,N_15182);
and U17980 (N_17980,N_15979,N_15155);
xor U17981 (N_17981,N_15798,N_15941);
xor U17982 (N_17982,N_14222,N_15305);
or U17983 (N_17983,N_14466,N_14749);
nand U17984 (N_17984,N_14865,N_15763);
xor U17985 (N_17985,N_14592,N_15629);
nor U17986 (N_17986,N_14288,N_14666);
and U17987 (N_17987,N_14975,N_14152);
nor U17988 (N_17988,N_14328,N_15848);
or U17989 (N_17989,N_15647,N_15034);
nor U17990 (N_17990,N_15327,N_15912);
xnor U17991 (N_17991,N_15657,N_14836);
xnor U17992 (N_17992,N_14867,N_14485);
and U17993 (N_17993,N_14222,N_15078);
nand U17994 (N_17994,N_15578,N_15657);
nand U17995 (N_17995,N_15437,N_15719);
xor U17996 (N_17996,N_14221,N_15853);
nor U17997 (N_17997,N_14389,N_14303);
xnor U17998 (N_17998,N_15640,N_14322);
xor U17999 (N_17999,N_14529,N_15742);
nand U18000 (N_18000,N_16945,N_17267);
or U18001 (N_18001,N_17493,N_16320);
and U18002 (N_18002,N_16365,N_16037);
xnor U18003 (N_18003,N_16327,N_17837);
xor U18004 (N_18004,N_16455,N_16617);
or U18005 (N_18005,N_17399,N_16470);
or U18006 (N_18006,N_17830,N_17858);
or U18007 (N_18007,N_17347,N_17857);
nor U18008 (N_18008,N_17868,N_17632);
nand U18009 (N_18009,N_16414,N_17400);
and U18010 (N_18010,N_17738,N_16423);
xnor U18011 (N_18011,N_17426,N_17051);
nor U18012 (N_18012,N_17379,N_17249);
xnor U18013 (N_18013,N_16877,N_16433);
xor U18014 (N_18014,N_16927,N_17986);
and U18015 (N_18015,N_16534,N_17316);
or U18016 (N_18016,N_17431,N_16641);
nand U18017 (N_18017,N_17303,N_17617);
nor U18018 (N_18018,N_16102,N_17983);
nor U18019 (N_18019,N_16647,N_17045);
and U18020 (N_18020,N_16055,N_16336);
or U18021 (N_18021,N_17147,N_17787);
and U18022 (N_18022,N_17896,N_17615);
and U18023 (N_18023,N_16438,N_17409);
nor U18024 (N_18024,N_16799,N_17958);
xnor U18025 (N_18025,N_17470,N_17319);
xnor U18026 (N_18026,N_17800,N_16409);
nor U18027 (N_18027,N_17245,N_17670);
xnor U18028 (N_18028,N_17818,N_16712);
or U18029 (N_18029,N_17263,N_16563);
nand U18030 (N_18030,N_17481,N_17397);
nor U18031 (N_18031,N_17349,N_17386);
xor U18032 (N_18032,N_16658,N_17534);
nor U18033 (N_18033,N_17772,N_16598);
or U18034 (N_18034,N_17852,N_16407);
xor U18035 (N_18035,N_16491,N_16541);
xnor U18036 (N_18036,N_16187,N_16761);
xnor U18037 (N_18037,N_17079,N_16502);
or U18038 (N_18038,N_17124,N_17658);
xnor U18039 (N_18039,N_16432,N_17626);
xnor U18040 (N_18040,N_17246,N_17304);
or U18041 (N_18041,N_16305,N_16169);
nor U18042 (N_18042,N_16479,N_16946);
nand U18043 (N_18043,N_17086,N_16894);
xnor U18044 (N_18044,N_16477,N_17418);
xnor U18045 (N_18045,N_16752,N_16175);
and U18046 (N_18046,N_17341,N_16258);
nand U18047 (N_18047,N_17491,N_17854);
or U18048 (N_18048,N_16482,N_16329);
or U18049 (N_18049,N_17904,N_17849);
nor U18050 (N_18050,N_17378,N_17111);
and U18051 (N_18051,N_16796,N_16679);
nand U18052 (N_18052,N_17413,N_16643);
xor U18053 (N_18053,N_17106,N_16704);
nor U18054 (N_18054,N_16434,N_17607);
nor U18055 (N_18055,N_17680,N_16552);
and U18056 (N_18056,N_17826,N_17814);
and U18057 (N_18057,N_16772,N_17974);
or U18058 (N_18058,N_16484,N_17699);
xnor U18059 (N_18059,N_17042,N_17411);
and U18060 (N_18060,N_17057,N_16852);
nand U18061 (N_18061,N_16442,N_16039);
and U18062 (N_18062,N_16095,N_16741);
nor U18063 (N_18063,N_17237,N_16141);
nand U18064 (N_18064,N_17564,N_16022);
xnor U18065 (N_18065,N_17601,N_17385);
or U18066 (N_18066,N_17761,N_16122);
and U18067 (N_18067,N_17944,N_17038);
or U18068 (N_18068,N_17192,N_16726);
nand U18069 (N_18069,N_17420,N_17158);
xor U18070 (N_18070,N_16332,N_17355);
or U18071 (N_18071,N_17825,N_16463);
xor U18072 (N_18072,N_17331,N_16357);
nand U18073 (N_18073,N_17724,N_16996);
or U18074 (N_18074,N_16253,N_16871);
and U18075 (N_18075,N_17504,N_17408);
and U18076 (N_18076,N_16801,N_16536);
or U18077 (N_18077,N_17044,N_16924);
nor U18078 (N_18078,N_16225,N_16939);
or U18079 (N_18079,N_16417,N_17628);
xor U18080 (N_18080,N_17438,N_17707);
or U18081 (N_18081,N_16845,N_16166);
nor U18082 (N_18082,N_17821,N_16553);
nand U18083 (N_18083,N_16354,N_16628);
xnor U18084 (N_18084,N_17477,N_17603);
and U18085 (N_18085,N_16256,N_17170);
and U18086 (N_18086,N_16723,N_16908);
nor U18087 (N_18087,N_17040,N_17517);
xnor U18088 (N_18088,N_16465,N_16870);
xnor U18089 (N_18089,N_17643,N_16431);
and U18090 (N_18090,N_17653,N_17667);
and U18091 (N_18091,N_17600,N_16016);
nand U18092 (N_18092,N_16749,N_17046);
nand U18093 (N_18093,N_17965,N_16076);
nor U18094 (N_18094,N_17035,N_16952);
xor U18095 (N_18095,N_17661,N_16065);
nand U18096 (N_18096,N_17563,N_17336);
or U18097 (N_18097,N_16060,N_16675);
nand U18098 (N_18098,N_17613,N_17995);
or U18099 (N_18099,N_16289,N_16367);
xnor U18100 (N_18100,N_17977,N_17796);
xor U18101 (N_18101,N_17509,N_17294);
and U18102 (N_18102,N_16506,N_17082);
nand U18103 (N_18103,N_16212,N_16094);
nor U18104 (N_18104,N_17704,N_17196);
or U18105 (N_18105,N_17165,N_17570);
xnor U18106 (N_18106,N_16974,N_16815);
and U18107 (N_18107,N_17520,N_16269);
xor U18108 (N_18108,N_16021,N_17396);
nor U18109 (N_18109,N_17608,N_17711);
xor U18110 (N_18110,N_17545,N_17903);
or U18111 (N_18111,N_17616,N_17952);
nand U18112 (N_18112,N_17181,N_17898);
or U18113 (N_18113,N_17480,N_16035);
xor U18114 (N_18114,N_16317,N_17195);
nor U18115 (N_18115,N_17930,N_17815);
xnor U18116 (N_18116,N_17332,N_16003);
nor U18117 (N_18117,N_16259,N_17989);
nand U18118 (N_18118,N_17078,N_17164);
nand U18119 (N_18119,N_16048,N_16621);
nand U18120 (N_18120,N_17407,N_16719);
and U18121 (N_18121,N_17033,N_17059);
nor U18122 (N_18122,N_17286,N_16316);
and U18123 (N_18123,N_17573,N_16378);
and U18124 (N_18124,N_16400,N_16958);
nand U18125 (N_18125,N_16152,N_17853);
or U18126 (N_18126,N_16476,N_17424);
nor U18127 (N_18127,N_16464,N_16159);
or U18128 (N_18128,N_17657,N_17173);
or U18129 (N_18129,N_16979,N_16837);
xor U18130 (N_18130,N_17744,N_17076);
xor U18131 (N_18131,N_16177,N_16987);
or U18132 (N_18132,N_16825,N_17439);
nand U18133 (N_18133,N_16383,N_17112);
nand U18134 (N_18134,N_17373,N_16229);
xnor U18135 (N_18135,N_17169,N_16277);
nor U18136 (N_18136,N_16665,N_17143);
xor U18137 (N_18137,N_16827,N_17004);
xnor U18138 (N_18138,N_17968,N_17136);
nor U18139 (N_18139,N_17646,N_16066);
or U18140 (N_18140,N_17978,N_17333);
nor U18141 (N_18141,N_17101,N_17579);
xnor U18142 (N_18142,N_17864,N_17037);
nor U18143 (N_18143,N_16889,N_17931);
nand U18144 (N_18144,N_16089,N_16004);
nand U18145 (N_18145,N_17861,N_17999);
and U18146 (N_18146,N_16707,N_16554);
nand U18147 (N_18147,N_16828,N_17956);
and U18148 (N_18148,N_17257,N_16855);
nor U18149 (N_18149,N_17302,N_17519);
nor U18150 (N_18150,N_16086,N_16309);
or U18151 (N_18151,N_16950,N_17322);
nor U18152 (N_18152,N_16514,N_16411);
or U18153 (N_18153,N_16488,N_17758);
xor U18154 (N_18154,N_17639,N_17532);
xor U18155 (N_18155,N_16054,N_17511);
xnor U18156 (N_18156,N_17911,N_16948);
xor U18157 (N_18157,N_16669,N_16728);
nor U18158 (N_18158,N_17248,N_17940);
xnor U18159 (N_18159,N_17024,N_17406);
and U18160 (N_18160,N_17705,N_17605);
xor U18161 (N_18161,N_17323,N_17924);
nor U18162 (N_18162,N_16914,N_17805);
or U18163 (N_18163,N_16616,N_17116);
xor U18164 (N_18164,N_16452,N_16027);
xnor U18165 (N_18165,N_17630,N_17466);
xnor U18166 (N_18166,N_16623,N_16100);
and U18167 (N_18167,N_16489,N_16765);
xnor U18168 (N_18168,N_17660,N_17404);
nand U18169 (N_18169,N_16687,N_16912);
xor U18170 (N_18170,N_16971,N_17132);
and U18171 (N_18171,N_16597,N_17859);
xnor U18172 (N_18172,N_17186,N_16814);
xnor U18173 (N_18173,N_16018,N_17296);
and U18174 (N_18174,N_16026,N_17812);
xnor U18175 (N_18175,N_17879,N_17395);
nand U18176 (N_18176,N_16267,N_16626);
and U18177 (N_18177,N_16300,N_17951);
xnor U18178 (N_18178,N_16983,N_17593);
xnor U18179 (N_18179,N_16634,N_17065);
xnor U18180 (N_18180,N_17539,N_16943);
xnor U18181 (N_18181,N_17561,N_17054);
and U18182 (N_18182,N_16933,N_17454);
or U18183 (N_18183,N_17401,N_16347);
or U18184 (N_18184,N_17039,N_17732);
or U18185 (N_18185,N_16091,N_17932);
nor U18186 (N_18186,N_17916,N_16053);
nand U18187 (N_18187,N_17206,N_16809);
or U18188 (N_18188,N_16333,N_16802);
or U18189 (N_18189,N_17277,N_16394);
or U18190 (N_18190,N_16330,N_16388);
and U18191 (N_18191,N_16693,N_16263);
nor U18192 (N_18192,N_17364,N_16445);
or U18193 (N_18193,N_17550,N_17856);
xnor U18194 (N_18194,N_16956,N_17394);
xnor U18195 (N_18195,N_17633,N_17252);
nor U18196 (N_18196,N_16603,N_16389);
nand U18197 (N_18197,N_17947,N_16627);
or U18198 (N_18198,N_16072,N_16197);
nor U18199 (N_18199,N_17216,N_17448);
xor U18200 (N_18200,N_16991,N_17749);
and U18201 (N_18201,N_17972,N_17266);
nor U18202 (N_18202,N_16232,N_16740);
nor U18203 (N_18203,N_17130,N_16947);
nand U18204 (N_18204,N_17558,N_16247);
or U18205 (N_18205,N_17486,N_16920);
xnor U18206 (N_18206,N_17979,N_16210);
nor U18207 (N_18207,N_17367,N_17447);
and U18208 (N_18208,N_16396,N_17375);
xor U18209 (N_18209,N_17352,N_17359);
or U18210 (N_18210,N_17645,N_17182);
or U18211 (N_18211,N_17953,N_16574);
nand U18212 (N_18212,N_17737,N_16182);
xor U18213 (N_18213,N_16499,N_17733);
and U18214 (N_18214,N_16490,N_16478);
nand U18215 (N_18215,N_17089,N_16965);
xnor U18216 (N_18216,N_16112,N_16174);
nand U18217 (N_18217,N_17831,N_17325);
or U18218 (N_18218,N_17567,N_16891);
and U18219 (N_18219,N_16521,N_17955);
nand U18220 (N_18220,N_17048,N_17068);
xnor U18221 (N_18221,N_17631,N_17058);
or U18222 (N_18222,N_17416,N_17338);
and U18223 (N_18223,N_16884,N_16328);
nor U18224 (N_18224,N_16077,N_17405);
or U18225 (N_18225,N_17782,N_17963);
or U18226 (N_18226,N_16671,N_17050);
xor U18227 (N_18227,N_16880,N_17368);
and U18228 (N_18228,N_17872,N_17877);
xnor U18229 (N_18229,N_16038,N_17180);
nor U18230 (N_18230,N_16878,N_16296);
and U18231 (N_18231,N_16691,N_16986);
or U18232 (N_18232,N_17213,N_17345);
or U18233 (N_18233,N_17356,N_17824);
nand U18234 (N_18234,N_16994,N_17559);
and U18235 (N_18235,N_17941,N_16846);
and U18236 (N_18236,N_16406,N_16198);
and U18237 (N_18237,N_16123,N_16051);
nor U18238 (N_18238,N_16075,N_17775);
nand U18239 (N_18239,N_16017,N_16238);
nand U18240 (N_18240,N_16458,N_17449);
and U18241 (N_18241,N_16261,N_17599);
or U18242 (N_18242,N_17566,N_17942);
and U18243 (N_18243,N_16941,N_16689);
xor U18244 (N_18244,N_17232,N_17746);
or U18245 (N_18245,N_16841,N_16913);
and U18246 (N_18246,N_17803,N_17668);
and U18247 (N_18247,N_16766,N_16613);
nand U18248 (N_18248,N_17500,N_17701);
and U18249 (N_18249,N_17790,N_16226);
xor U18250 (N_18250,N_16372,N_16892);
and U18251 (N_18251,N_16448,N_17648);
or U18252 (N_18252,N_16154,N_17372);
and U18253 (N_18253,N_17311,N_16677);
xor U18254 (N_18254,N_17217,N_16708);
nand U18255 (N_18255,N_16678,N_16813);
and U18256 (N_18256,N_17159,N_17880);
or U18257 (N_18257,N_16271,N_17465);
and U18258 (N_18258,N_16160,N_16467);
nor U18259 (N_18259,N_16046,N_16936);
and U18260 (N_18260,N_16844,N_17185);
or U18261 (N_18261,N_17090,N_16771);
nor U18262 (N_18262,N_17384,N_17262);
xnor U18263 (N_18263,N_17560,N_17191);
or U18264 (N_18264,N_17851,N_17734);
nand U18265 (N_18265,N_17227,N_17118);
and U18266 (N_18266,N_16872,N_17918);
nand U18267 (N_18267,N_16366,N_16888);
nor U18268 (N_18268,N_16217,N_17526);
nand U18269 (N_18269,N_17684,N_17835);
nand U18270 (N_18270,N_17820,N_16120);
nor U18271 (N_18271,N_16234,N_16577);
and U18272 (N_18272,N_16509,N_17265);
or U18273 (N_18273,N_17921,N_16183);
nand U18274 (N_18274,N_16472,N_16443);
and U18275 (N_18275,N_17353,N_16096);
xor U18276 (N_18276,N_16565,N_17010);
nand U18277 (N_18277,N_16963,N_16722);
and U18278 (N_18278,N_16688,N_16715);
nor U18279 (N_18279,N_16020,N_16228);
or U18280 (N_18280,N_16293,N_17551);
nand U18281 (N_18281,N_17402,N_16466);
nand U18282 (N_18282,N_16049,N_16770);
nand U18283 (N_18283,N_16133,N_17369);
nand U18284 (N_18284,N_16650,N_16631);
and U18285 (N_18285,N_17209,N_17105);
nor U18286 (N_18286,N_17505,N_16206);
and U18287 (N_18287,N_17458,N_17894);
nand U18288 (N_18288,N_17691,N_16356);
xnor U18289 (N_18289,N_17934,N_16346);
nor U18290 (N_18290,N_17021,N_17268);
xor U18291 (N_18291,N_17142,N_17269);
nand U18292 (N_18292,N_17022,N_16644);
nor U18293 (N_18293,N_17487,N_16475);
nor U18294 (N_18294,N_17905,N_16268);
xor U18295 (N_18295,N_17730,N_16731);
nand U18296 (N_18296,N_17664,N_17243);
and U18297 (N_18297,N_16736,N_17552);
xnor U18298 (N_18298,N_16071,N_16056);
nand U18299 (N_18299,N_16656,N_17069);
xnor U18300 (N_18300,N_16000,N_17484);
nand U18301 (N_18301,N_17053,N_16585);
or U18302 (N_18302,N_17721,N_16286);
xor U18303 (N_18303,N_17537,N_17308);
xor U18304 (N_18304,N_16753,N_16917);
or U18305 (N_18305,N_17771,N_17827);
xor U18306 (N_18306,N_16150,N_16483);
or U18307 (N_18307,N_16042,N_17187);
or U18308 (N_18308,N_16163,N_16204);
nand U18309 (N_18309,N_17494,N_17717);
and U18310 (N_18310,N_17507,N_16216);
and U18311 (N_18311,N_16280,N_17671);
nand U18312 (N_18312,N_17629,N_16875);
or U18313 (N_18313,N_16103,N_16194);
nand U18314 (N_18314,N_16240,N_16450);
xnor U18315 (N_18315,N_17127,N_17697);
xnor U18316 (N_18316,N_17284,N_17572);
nand U18317 (N_18317,N_17817,N_17502);
or U18318 (N_18318,N_16395,N_17299);
nand U18319 (N_18319,N_16486,N_16350);
and U18320 (N_18320,N_16193,N_16024);
xnor U18321 (N_18321,N_17225,N_17530);
xnor U18322 (N_18322,N_16816,N_17920);
xnor U18323 (N_18323,N_17329,N_16782);
and U18324 (N_18324,N_16854,N_16324);
nor U18325 (N_18325,N_17461,N_16680);
nand U18326 (N_18326,N_17642,N_16543);
nor U18327 (N_18327,N_17890,N_16568);
nor U18328 (N_18328,N_17576,N_16526);
xnor U18329 (N_18329,N_16700,N_16611);
or U18330 (N_18330,N_16062,N_16570);
nand U18331 (N_18331,N_17205,N_17843);
or U18332 (N_18332,N_17478,N_16571);
and U18333 (N_18333,N_16223,N_17808);
nand U18334 (N_18334,N_17832,N_16348);
and U18335 (N_18335,N_17712,N_16713);
nor U18336 (N_18336,N_16207,N_16380);
and U18337 (N_18337,N_16322,N_16564);
xnor U18338 (N_18338,N_17155,N_17914);
and U18339 (N_18339,N_17003,N_16800);
nor U18340 (N_18340,N_17000,N_17574);
xnor U18341 (N_18341,N_16849,N_17289);
and U18342 (N_18342,N_17641,N_16145);
nor U18343 (N_18343,N_16014,N_17043);
and U18344 (N_18344,N_16951,N_17398);
xnor U18345 (N_18345,N_16319,N_17907);
nor U18346 (N_18346,N_16338,N_17957);
nand U18347 (N_18347,N_16701,N_17423);
and U18348 (N_18348,N_16528,N_16977);
and U18349 (N_18349,N_16542,N_17241);
or U18350 (N_18350,N_16524,N_16546);
or U18351 (N_18351,N_16980,N_16137);
or U18352 (N_18352,N_17866,N_16714);
xnor U18353 (N_18353,N_17365,N_16454);
nand U18354 (N_18354,N_16808,N_16034);
xor U18355 (N_18355,N_16733,N_16525);
or U18356 (N_18356,N_17871,N_16052);
nand U18357 (N_18357,N_17340,N_16144);
and U18358 (N_18358,N_16659,N_17131);
or U18359 (N_18359,N_17926,N_17233);
and U18360 (N_18360,N_16116,N_17001);
or U18361 (N_18361,N_17627,N_16002);
xnor U18362 (N_18362,N_16461,N_16010);
xnor U18363 (N_18363,N_17910,N_17873);
nor U18364 (N_18364,N_17703,N_17997);
nor U18365 (N_18365,N_17230,N_17203);
xnor U18366 (N_18366,N_17736,N_16186);
and U18367 (N_18367,N_17214,N_17363);
nor U18368 (N_18368,N_17377,N_17063);
xnor U18369 (N_18369,N_17344,N_17488);
and U18370 (N_18370,N_17897,N_16364);
xor U18371 (N_18371,N_17636,N_17121);
nor U18372 (N_18372,N_17207,N_16969);
or U18373 (N_18373,N_16764,N_17463);
xnor U18374 (N_18374,N_17093,N_17188);
nand U18375 (N_18375,N_17157,N_16902);
or U18376 (N_18376,N_17524,N_17472);
or U18377 (N_18377,N_17666,N_16692);
and U18378 (N_18378,N_16201,N_16928);
nor U18379 (N_18379,N_17860,N_17318);
xnor U18380 (N_18380,N_16119,N_17693);
or U18381 (N_18381,N_17473,N_17435);
nor U18382 (N_18382,N_16398,N_16676);
and U18383 (N_18383,N_17343,N_16429);
or U18384 (N_18384,N_16547,N_17088);
and U18385 (N_18385,N_16428,N_16517);
nand U18386 (N_18386,N_17716,N_16751);
nand U18387 (N_18387,N_16789,N_17211);
nand U18388 (N_18388,N_16074,N_16755);
and U18389 (N_18389,N_16529,N_16784);
or U18390 (N_18390,N_17961,N_16876);
and U18391 (N_18391,N_16698,N_16684);
xnor U18392 (N_18392,N_17816,N_16909);
or U18393 (N_18393,N_16278,N_16363);
nor U18394 (N_18394,N_16349,N_17153);
nor U18395 (N_18395,N_16720,N_16817);
nand U18396 (N_18396,N_16505,N_17747);
xnor U18397 (N_18397,N_16161,N_16615);
or U18398 (N_18398,N_17119,N_16069);
and U18399 (N_18399,N_16850,N_17171);
or U18400 (N_18400,N_16744,N_16538);
xor U18401 (N_18401,N_16427,N_17982);
nor U18402 (N_18402,N_17933,N_16110);
nand U18403 (N_18403,N_16622,N_16215);
nor U18404 (N_18404,N_17019,N_16031);
nor U18405 (N_18405,N_17391,N_16520);
xor U18406 (N_18406,N_17767,N_17075);
nor U18407 (N_18407,N_16132,N_17967);
xnor U18408 (N_18408,N_16625,N_16606);
nor U18409 (N_18409,N_17177,N_16890);
nor U18410 (N_18410,N_17624,N_17374);
xor U18411 (N_18411,N_16067,N_17428);
and U18412 (N_18412,N_17702,N_16581);
or U18413 (N_18413,N_17640,N_16783);
and U18414 (N_18414,N_17715,N_16449);
nor U18415 (N_18415,N_17134,N_17381);
and U18416 (N_18416,N_16359,N_17023);
nor U18417 (N_18417,N_17223,N_17445);
nor U18418 (N_18418,N_17726,N_16165);
and U18419 (N_18419,N_17899,N_16230);
nor U18420 (N_18420,N_17609,N_17497);
or U18421 (N_18421,N_17313,N_17389);
nand U18422 (N_18422,N_17888,N_16862);
xor U18423 (N_18423,N_16737,N_17595);
or U18424 (N_18424,N_17651,N_17833);
or U18425 (N_18425,N_16982,N_16584);
and U18426 (N_18426,N_17490,N_16379);
or U18427 (N_18427,N_16162,N_16325);
nand U18428 (N_18428,N_17301,N_17783);
and U18429 (N_18429,N_16015,N_16297);
xnor U18430 (N_18430,N_17320,N_17577);
xor U18431 (N_18431,N_17973,N_17208);
nor U18432 (N_18432,N_17553,N_17244);
nand U18433 (N_18433,N_16390,N_16041);
or U18434 (N_18434,N_17809,N_17793);
xnor U18435 (N_18435,N_16662,N_17917);
xor U18436 (N_18436,N_16361,N_16605);
or U18437 (N_18437,N_17228,N_17072);
xor U18438 (N_18438,N_16822,N_17723);
xnor U18439 (N_18439,N_17672,N_16311);
and U18440 (N_18440,N_16926,N_16370);
nand U18441 (N_18441,N_17635,N_16342);
and U18442 (N_18442,N_17030,N_16468);
or U18443 (N_18443,N_16196,N_16453);
or U18444 (N_18444,N_17988,N_16670);
and U18445 (N_18445,N_17229,N_16516);
and U18446 (N_18446,N_16385,N_16494);
or U18447 (N_18447,N_16308,N_16113);
nor U18448 (N_18448,N_16820,N_16353);
or U18449 (N_18449,N_16237,N_16136);
or U18450 (N_18450,N_17240,N_17234);
or U18451 (N_18451,N_16369,N_16738);
and U18452 (N_18452,N_17383,N_17762);
and U18453 (N_18453,N_16421,N_17026);
xnor U18454 (N_18454,N_16885,N_16242);
nor U18455 (N_18455,N_17791,N_17235);
and U18456 (N_18456,N_17120,N_16633);
xor U18457 (N_18457,N_16887,N_17334);
or U18458 (N_18458,N_16661,N_16444);
nor U18459 (N_18459,N_17770,N_16382);
and U18460 (N_18460,N_17695,N_16460);
xor U18461 (N_18461,N_16968,N_16863);
xor U18462 (N_18462,N_16265,N_17698);
xnor U18463 (N_18463,N_16674,N_17427);
nand U18464 (N_18464,N_16595,N_16180);
nor U18465 (N_18465,N_16548,N_17278);
xor U18466 (N_18466,N_16420,N_17527);
nor U18467 (N_18467,N_16776,N_16006);
and U18468 (N_18468,N_17819,N_16569);
and U18469 (N_18469,N_16009,N_17007);
nor U18470 (N_18470,N_17923,N_16043);
nand U18471 (N_18471,N_16867,N_16612);
nand U18472 (N_18472,N_16593,N_16527);
and U18473 (N_18473,N_17806,N_17432);
xor U18474 (N_18474,N_16940,N_17959);
nor U18475 (N_18475,N_16896,N_17501);
xor U18476 (N_18476,N_16115,N_17360);
nor U18477 (N_18477,N_16233,N_17434);
or U18478 (N_18478,N_16904,N_17900);
xor U18479 (N_18479,N_17795,N_16893);
nor U18480 (N_18480,N_16164,N_17760);
or U18481 (N_18481,N_17288,N_16575);
and U18482 (N_18482,N_16866,N_17788);
xor U18483 (N_18483,N_16405,N_17807);
or U18484 (N_18484,N_16403,N_16754);
nor U18485 (N_18485,N_16590,N_16847);
xnor U18486 (N_18486,N_17138,N_16070);
or U18487 (N_18487,N_16386,N_17694);
nor U18488 (N_18488,N_16531,N_16638);
nor U18489 (N_18489,N_16306,N_17324);
nand U18490 (N_18490,N_17380,N_16030);
nor U18491 (N_18491,N_16774,N_17557);
xor U18492 (N_18492,N_17433,N_17714);
nor U18493 (N_18493,N_16649,N_16029);
nand U18494 (N_18494,N_16567,N_16729);
xnor U18495 (N_18495,N_17204,N_17222);
nand U18496 (N_18496,N_17425,N_16047);
or U18497 (N_18497,N_16922,N_17597);
nand U18498 (N_18498,N_17682,N_16139);
and U18499 (N_18499,N_17588,N_16932);
nand U18500 (N_18500,N_16185,N_16785);
nor U18501 (N_18501,N_16970,N_16860);
nor U18502 (N_18502,N_17471,N_16710);
nor U18503 (N_18503,N_17655,N_17467);
or U18504 (N_18504,N_16099,N_16843);
and U18505 (N_18505,N_17778,N_17906);
or U18506 (N_18506,N_16859,N_17798);
or U18507 (N_18507,N_16063,N_16480);
xor U18508 (N_18508,N_17878,N_16111);
xnor U18509 (N_18509,N_16879,N_17312);
nand U18510 (N_18510,N_16537,N_17102);
nor U18511 (N_18511,N_16344,N_16697);
or U18512 (N_18512,N_17455,N_16518);
or U18513 (N_18513,N_16387,N_16239);
nand U18514 (N_18514,N_16826,N_17621);
nand U18515 (N_18515,N_16642,N_16657);
nand U18516 (N_18516,N_16231,N_16422);
xnor U18517 (N_18517,N_16830,N_16257);
or U18518 (N_18518,N_16149,N_16243);
and U18519 (N_18519,N_16279,N_17137);
xor U18520 (N_18520,N_17960,N_16558);
or U18521 (N_18521,N_17061,N_17135);
nand U18522 (N_18522,N_17274,N_17183);
nand U18523 (N_18523,N_17838,N_17869);
xor U18524 (N_18524,N_16497,N_16362);
or U18525 (N_18525,N_16646,N_17128);
nor U18526 (N_18526,N_16147,N_17547);
or U18527 (N_18527,N_17498,N_16533);
xnor U18528 (N_18528,N_16787,N_16759);
and U18529 (N_18529,N_16864,N_16779);
xnor U18530 (N_18530,N_16682,N_16532);
or U18531 (N_18531,N_16651,N_17256);
nand U18532 (N_18532,N_16672,N_16610);
nand U18533 (N_18533,N_16959,N_17700);
nor U18534 (N_18534,N_16260,N_17895);
and U18535 (N_18535,N_17006,N_17863);
and U18536 (N_18536,N_17748,N_16307);
xnor U18537 (N_18537,N_17419,N_17594);
or U18538 (N_18538,N_16495,N_17935);
and U18539 (N_18539,N_17283,N_16900);
or U18540 (N_18540,N_16189,N_16995);
or U18541 (N_18541,N_16459,N_16381);
nand U18542 (N_18542,N_17785,N_17789);
and U18543 (N_18543,N_17876,N_17113);
nor U18544 (N_18544,N_17516,N_17829);
nand U18545 (N_18545,N_17290,N_17168);
or U18546 (N_18546,N_16976,N_17271);
or U18547 (N_18547,N_16221,N_16469);
and U18548 (N_18548,N_17786,N_16806);
and U18549 (N_18549,N_17011,N_16918);
nand U18550 (N_18550,N_17104,N_17291);
and U18551 (N_18551,N_17768,N_17885);
xnor U18552 (N_18552,N_16934,N_17731);
and U18553 (N_18553,N_16653,N_16775);
nand U18554 (N_18554,N_17056,N_16340);
or U18555 (N_18555,N_16447,N_17300);
and U18556 (N_18556,N_17985,N_17328);
and U18557 (N_18557,N_16792,N_17669);
nor U18558 (N_18558,N_17912,N_16375);
xor U18559 (N_18559,N_16769,N_17287);
nand U18560 (N_18560,N_16222,N_16906);
nor U18561 (N_18561,N_16107,N_17310);
xnor U18562 (N_18562,N_17752,N_17247);
nand U18563 (N_18563,N_16551,N_17865);
nand U18564 (N_18564,N_17390,N_16410);
and U18565 (N_18565,N_16578,N_16953);
nor U18566 (N_18566,N_16718,N_17751);
xnor U18567 (N_18567,N_17315,N_16954);
xnor U18568 (N_18568,N_16739,N_17529);
or U18569 (N_18569,N_17565,N_17462);
nor U18570 (N_18570,N_16192,N_17083);
xnor U18571 (N_18571,N_17499,N_17718);
and U18572 (N_18572,N_16637,N_17676);
or U18573 (N_18573,N_16392,N_17219);
xnor U18574 (N_18574,N_16760,N_16143);
and U18575 (N_18575,N_16446,N_16794);
xor U18576 (N_18576,N_16492,N_16176);
and U18577 (N_18577,N_17251,N_17870);
or U18578 (N_18578,N_16451,N_16937);
nor U18579 (N_18579,N_16660,N_17335);
xnor U18580 (N_18580,N_16999,N_17166);
xor U18581 (N_18581,N_16081,N_17073);
nand U18582 (N_18582,N_16903,N_17140);
nand U18583 (N_18583,N_17663,N_16975);
nand U18584 (N_18584,N_16856,N_16078);
nor U18585 (N_18585,N_16168,N_16786);
nand U18586 (N_18586,N_17525,N_16762);
or U18587 (N_18587,N_16973,N_17417);
or U18588 (N_18588,N_17969,N_17755);
and U18589 (N_18589,N_16415,N_17675);
xor U18590 (N_18590,N_16402,N_16252);
or U18591 (N_18591,N_17250,N_16858);
or U18592 (N_18592,N_16624,N_17456);
xnor U18593 (N_18593,N_16313,N_17351);
xnor U18594 (N_18594,N_16282,N_16833);
xnor U18595 (N_18595,N_16050,N_17518);
or U18596 (N_18596,N_17867,N_17238);
and U18597 (N_18597,N_17686,N_16128);
xnor U18598 (N_18598,N_17279,N_16321);
nand U18599 (N_18599,N_17074,N_16435);
and U18600 (N_18600,N_16805,N_17314);
or U18601 (N_18601,N_17100,N_16040);
xnor U18602 (N_18602,N_17652,N_16685);
or U18603 (N_18603,N_17990,N_17991);
nand U18604 (N_18604,N_17254,N_17647);
nand U18605 (N_18605,N_16886,N_17741);
or U18606 (N_18606,N_17508,N_16632);
xnor U18607 (N_18607,N_17810,N_16635);
xnor U18608 (N_18608,N_16440,N_16270);
nand U18609 (N_18609,N_17282,N_17496);
and U18610 (N_18610,N_17305,N_17679);
xor U18611 (N_18611,N_17307,N_17103);
nor U18612 (N_18612,N_16211,N_17713);
nand U18613 (N_18613,N_16910,N_16304);
nand U18614 (N_18614,N_16620,N_17882);
nor U18615 (N_18615,N_17792,N_16088);
and U18616 (N_18616,N_17049,N_16436);
and U18617 (N_18617,N_17841,N_17410);
and U18618 (N_18618,N_17618,N_17108);
xor U18619 (N_18619,N_17678,N_16559);
or U18620 (N_18620,N_16142,N_17457);
or U18621 (N_18621,N_17996,N_17779);
and U18622 (N_18622,N_17370,N_16942);
and U18623 (N_18623,N_16266,N_17388);
and U18624 (N_18624,N_16413,N_17008);
nand U18625 (N_18625,N_16129,N_16118);
or U18626 (N_18626,N_16706,N_17275);
and U18627 (N_18627,N_17092,N_16838);
nand U18628 (N_18628,N_16523,N_16273);
nand U18629 (N_18629,N_17306,N_16200);
xnor U18630 (N_18630,N_16673,N_17644);
nor U18631 (N_18631,N_17839,N_16345);
and U18632 (N_18632,N_16439,N_16530);
and U18633 (N_18633,N_17032,N_16961);
xnor U18634 (N_18634,N_16493,N_17440);
xnor U18635 (N_18635,N_17415,N_17587);
nand U18636 (N_18636,N_17915,N_16501);
nand U18637 (N_18637,N_17688,N_16057);
nor U18638 (N_18638,N_17149,N_16178);
and U18639 (N_18639,N_16007,N_16323);
nand U18640 (N_18640,N_17850,N_17638);
and U18641 (N_18641,N_17596,N_16384);
nor U18642 (N_18642,N_16834,N_16972);
or U18643 (N_18643,N_17522,N_17548);
xor U18644 (N_18644,N_16609,N_17141);
or U18645 (N_18645,N_17115,N_16848);
nor U18646 (N_18646,N_16295,N_16540);
and U18647 (N_18647,N_16869,N_16275);
or U18648 (N_18648,N_16795,N_17606);
nand U18649 (N_18649,N_16507,N_17893);
nand U18650 (N_18650,N_16033,N_16032);
or U18651 (N_18651,N_17110,N_16172);
nand U18652 (N_18652,N_16861,N_17327);
and U18653 (N_18653,N_17099,N_16868);
or U18654 (N_18654,N_17862,N_17673);
or U18655 (N_18655,N_17276,N_17450);
xnor U18656 (N_18656,N_17634,N_16219);
xor U18657 (N_18657,N_16085,N_16683);
nor U18658 (N_18658,N_17571,N_17902);
nand U18659 (N_18659,N_16905,N_17881);
and U18660 (N_18660,N_16248,N_17084);
nand U18661 (N_18661,N_17781,N_17346);
or U18662 (N_18662,N_16246,N_17909);
nor U18663 (N_18663,N_16984,N_17492);
xor U18664 (N_18664,N_16923,N_17009);
or U18665 (N_18665,N_17231,N_16907);
nor U18666 (N_18666,N_16227,N_17681);
nor U18667 (N_18667,N_16245,N_17358);
xnor U18668 (N_18668,N_17085,N_17757);
nand U18669 (N_18669,N_17366,N_16874);
nand U18670 (N_18670,N_16292,N_16510);
nand U18671 (N_18671,N_16456,N_16373);
and U18672 (N_18672,N_16619,N_17929);
or U18673 (N_18673,N_16512,N_17954);
or U18674 (N_18674,N_16011,N_16716);
xor U18675 (N_18675,N_17950,N_16462);
and U18676 (N_18676,N_16068,N_16899);
xor U18677 (N_18677,N_16135,N_16989);
and U18678 (N_18678,N_17354,N_16811);
nor U18679 (N_18679,N_16339,N_17535);
or U18680 (N_18680,N_17735,N_17993);
xor U18681 (N_18681,N_16374,N_16990);
or U18682 (N_18682,N_16709,N_17016);
xnor U18683 (N_18683,N_16544,N_16073);
nand U18684 (N_18684,N_16272,N_16285);
xnor U18685 (N_18685,N_17293,N_17943);
nor U18686 (N_18686,N_17875,N_16997);
xnor U18687 (N_18687,N_16930,N_17538);
nand U18688 (N_18688,N_17946,N_16654);
and U18689 (N_18689,N_16967,N_16262);
xor U18690 (N_18690,N_17855,N_17495);
nand U18691 (N_18691,N_16351,N_16005);
or U18692 (N_18692,N_17842,N_17218);
nand U18693 (N_18693,N_16284,N_17710);
nand U18694 (N_18694,N_16576,N_17503);
and U18695 (N_18695,N_17330,N_17031);
xor U18696 (N_18696,N_17107,N_16594);
nor U18697 (N_18697,N_16839,N_16473);
and U18698 (N_18698,N_17476,N_16249);
or U18699 (N_18699,N_17884,N_16742);
nor U18700 (N_18700,N_17309,N_16500);
nor U18701 (N_18701,N_17774,N_17095);
nand U18702 (N_18702,N_16173,N_16915);
and U18703 (N_18703,N_16746,N_17987);
nand U18704 (N_18704,N_16303,N_16244);
and U18705 (N_18705,N_17513,N_16401);
nor U18706 (N_18706,N_16114,N_16023);
or U18707 (N_18707,N_16318,N_16681);
nor U18708 (N_18708,N_17317,N_16522);
or U18709 (N_18709,N_16557,N_16580);
nor U18710 (N_18710,N_16334,N_16190);
nand U18711 (N_18711,N_17922,N_17272);
and U18712 (N_18712,N_17889,N_16727);
or U18713 (N_18713,N_17429,N_16315);
nor U18714 (N_18714,N_16944,N_16090);
and U18715 (N_18715,N_17094,N_16426);
nand U18716 (N_18716,N_17739,N_16425);
xor U18717 (N_18717,N_17556,N_16832);
or U18718 (N_18718,N_16895,N_17622);
nand U18719 (N_18719,N_16179,N_16218);
nor U18720 (N_18720,N_17925,N_17176);
nor U18721 (N_18721,N_17133,N_16124);
nand U18722 (N_18722,N_17592,N_17080);
and U18723 (N_18723,N_17590,N_16743);
nand U18724 (N_18724,N_16487,N_16812);
nor U18725 (N_18725,N_17371,N_16645);
nand U18726 (N_18726,N_17901,N_17285);
or U18727 (N_18727,N_17836,N_16368);
and U18728 (N_18728,N_16949,N_17096);
nand U18729 (N_18729,N_17804,N_16254);
nand U18730 (N_18730,N_17637,N_17280);
and U18731 (N_18731,N_17562,N_16664);
xor U18732 (N_18732,N_17485,N_16288);
or U18733 (N_18733,N_17589,N_16255);
and U18734 (N_18734,N_17297,N_17740);
xnor U18735 (N_18735,N_16703,N_16044);
xnor U18736 (N_18736,N_16778,N_16290);
or U18737 (N_18737,N_17614,N_16797);
nor U18738 (N_18738,N_16108,N_16310);
nor U18739 (N_18739,N_17625,N_17515);
xor U18740 (N_18740,N_16857,N_16092);
or U18741 (N_18741,N_17098,N_17430);
nor U18742 (N_18742,N_17834,N_17554);
xnor U18743 (N_18743,N_16202,N_17145);
and U18744 (N_18744,N_17117,N_17586);
nor U18745 (N_18745,N_17938,N_17025);
xor U18746 (N_18746,N_16083,N_17568);
nor U18747 (N_18747,N_17725,N_16485);
nand U18748 (N_18748,N_17984,N_16535);
xor U18749 (N_18749,N_16725,N_16780);
xor U18750 (N_18750,N_17239,N_17028);
xnor U18751 (N_18751,N_16601,N_16589);
or U18752 (N_18752,N_16851,N_17964);
and U18753 (N_18753,N_16705,N_16734);
xnor U18754 (N_18754,N_17692,N_16957);
xor U18755 (N_18755,N_17167,N_16962);
nor U18756 (N_18756,N_17580,N_16148);
and U18757 (N_18757,N_16481,N_17685);
xor U18758 (N_18758,N_16911,N_16629);
or U18759 (N_18759,N_16424,N_17193);
xor U18760 (N_18760,N_17066,N_17412);
xnor U18761 (N_18761,N_16562,N_16264);
or U18762 (N_18762,N_16341,N_16471);
or U18763 (N_18763,N_16355,N_16901);
nor U18764 (N_18764,N_17847,N_17253);
and U18765 (N_18765,N_16064,N_16702);
or U18766 (N_18766,N_16883,N_17569);
and U18767 (N_18767,N_17362,N_16981);
nor U18768 (N_18768,N_16276,N_17215);
nor U18769 (N_18769,N_17533,N_16019);
nand U18770 (N_18770,N_16195,N_17483);
nor U18771 (N_18771,N_17144,N_16993);
nand U18772 (N_18772,N_16640,N_17683);
nor U18773 (N_18773,N_16299,N_17939);
nor U18774 (N_18774,N_16602,N_16496);
xor U18775 (N_18775,N_17722,N_17706);
and U18776 (N_18776,N_17555,N_17052);
and U18777 (N_18777,N_16793,N_16084);
xnor U18778 (N_18778,N_16607,N_17339);
xor U18779 (N_18779,N_17220,N_17612);
nand U18780 (N_18780,N_16757,N_17598);
nand U18781 (N_18781,N_16690,N_17469);
or U18782 (N_18782,N_16199,N_17945);
or U18783 (N_18783,N_17754,N_16767);
xor U18784 (N_18784,N_16156,N_16668);
nand U18785 (N_18785,N_16209,N_17662);
or U18786 (N_18786,N_16663,N_17184);
and U18787 (N_18787,N_16404,N_16717);
nor U18788 (N_18788,N_16840,N_17994);
and U18789 (N_18789,N_16127,N_16573);
xor U18790 (N_18790,N_16790,N_17475);
and U18791 (N_18791,N_16087,N_16696);
and U18792 (N_18792,N_17659,N_17087);
nand U18793 (N_18793,N_17919,N_17321);
and U18794 (N_18794,N_16294,N_16437);
nor U18795 (N_18795,N_17654,N_16241);
and U18796 (N_18796,N_17583,N_16824);
nand U18797 (N_18797,N_17029,N_16960);
nor U18798 (N_18798,N_16515,N_17846);
or U18799 (N_18799,N_17146,N_16121);
and U18800 (N_18800,N_17689,N_17489);
xnor U18801 (N_18801,N_16819,N_17690);
and U18802 (N_18802,N_17474,N_16897);
xnor U18803 (N_18803,N_17845,N_16545);
or U18804 (N_18804,N_17403,N_17611);
nor U18805 (N_18805,N_17122,N_17777);
or U18806 (N_18806,N_16474,N_17212);
or U18807 (N_18807,N_17523,N_17756);
xor U18808 (N_18808,N_16001,N_17020);
or U18809 (N_18809,N_17081,N_17575);
or U18810 (N_18810,N_16314,N_16503);
or U18811 (N_18811,N_16929,N_17892);
xor U18812 (N_18812,N_16125,N_17055);
or U18813 (N_18813,N_16686,N_16818);
xnor U18814 (N_18814,N_16803,N_17602);
or U18815 (N_18815,N_16935,N_17521);
nand U18816 (N_18816,N_16013,N_17298);
xor U18817 (N_18817,N_16441,N_16109);
nor U18818 (N_18818,N_16931,N_17949);
or U18819 (N_18819,N_16730,N_16549);
nor U18820 (N_18820,N_16556,N_16829);
and U18821 (N_18821,N_17067,N_16138);
xor U18822 (N_18822,N_16331,N_16539);
xor U18823 (N_18823,N_17178,N_16093);
or U18824 (N_18824,N_16191,N_16140);
nand U18825 (N_18825,N_16807,N_16750);
xnor U18826 (N_18826,N_16591,N_17769);
and U18827 (N_18827,N_17510,N_16925);
nand U18828 (N_18828,N_17708,N_16788);
or U18829 (N_18829,N_16618,N_16337);
nor U18830 (N_18830,N_16105,N_16335);
nand U18831 (N_18831,N_17764,N_17540);
or U18832 (N_18832,N_16721,N_17543);
nand U18833 (N_18833,N_16921,N_16130);
or U18834 (N_18834,N_17034,N_16153);
nor U18835 (N_18835,N_17823,N_17281);
or U18836 (N_18836,N_17459,N_17582);
or U18837 (N_18837,N_17750,N_16695);
and U18838 (N_18838,N_17015,N_17002);
nand U18839 (N_18839,N_17970,N_16758);
nand U18840 (N_18840,N_17674,N_16416);
or U18841 (N_18841,N_16302,N_17392);
and U18842 (N_18842,N_17442,N_16988);
nand U18843 (N_18843,N_17013,N_17620);
xnor U18844 (N_18844,N_16058,N_17742);
or U18845 (N_18845,N_17236,N_16298);
nor U18846 (N_18846,N_16821,N_17773);
nand U18847 (N_18847,N_16666,N_16596);
and U18848 (N_18848,N_16352,N_16966);
nand U18849 (N_18849,N_17027,N_17528);
xnor U18850 (N_18850,N_16045,N_17696);
or U18851 (N_18851,N_17794,N_16012);
nor U18852 (N_18852,N_16964,N_17259);
or U18853 (N_18853,N_17163,N_16377);
nand U18854 (N_18854,N_16735,N_17584);
nor U18855 (N_18855,N_16274,N_17753);
nor U18856 (N_18856,N_17198,N_16235);
or U18857 (N_18857,N_16916,N_17041);
nand U18858 (N_18858,N_17585,N_16008);
xnor U18859 (N_18859,N_16236,N_17387);
or U18860 (N_18860,N_16391,N_16036);
and U18861 (N_18861,N_17541,N_16655);
and U18862 (N_18862,N_17650,N_16648);
or U18863 (N_18863,N_17446,N_16732);
nand U18864 (N_18864,N_17822,N_17179);
or U18865 (N_18865,N_16106,N_17071);
or U18866 (N_18866,N_17292,N_16511);
and U18867 (N_18867,N_17514,N_17813);
nor U18868 (N_18868,N_16079,N_17273);
xor U18869 (N_18869,N_17062,N_16371);
and U18870 (N_18870,N_16898,N_17414);
and U18871 (N_18871,N_17542,N_16214);
nor U18872 (N_18872,N_17936,N_16508);
nand U18873 (N_18873,N_16831,N_17971);
xnor U18874 (N_18874,N_17468,N_16810);
and U18875 (N_18875,N_17156,N_17948);
or U18876 (N_18876,N_16608,N_17077);
xnor U18877 (N_18877,N_16842,N_16171);
xnor U18878 (N_18878,N_16419,N_16283);
or U18879 (N_18879,N_17139,N_16513);
and U18880 (N_18880,N_16059,N_17591);
nand U18881 (N_18881,N_17148,N_16205);
nand U18882 (N_18882,N_16117,N_16061);
or U18883 (N_18883,N_16745,N_17126);
and U18884 (N_18884,N_17891,N_17709);
nand U18885 (N_18885,N_16157,N_17194);
or U18886 (N_18886,N_17546,N_16865);
and U18887 (N_18887,N_17190,N_16104);
nor U18888 (N_18888,N_16652,N_17844);
nand U18889 (N_18889,N_16853,N_16220);
nor U18890 (N_18890,N_17464,N_16748);
nor U18891 (N_18891,N_16586,N_17998);
or U18892 (N_18892,N_16992,N_16555);
nor U18893 (N_18893,N_17729,N_17656);
and U18894 (N_18894,N_17966,N_17913);
and U18895 (N_18895,N_17512,N_17114);
and U18896 (N_18896,N_16938,N_16151);
xor U18897 (N_18897,N_17975,N_16561);
nor U18898 (N_18898,N_17451,N_17258);
and U18899 (N_18899,N_17270,N_16504);
and U18900 (N_18900,N_16170,N_16101);
nand U18901 (N_18901,N_17436,N_16408);
and U18902 (N_18902,N_17357,N_16823);
and U18903 (N_18903,N_16155,N_17047);
nand U18904 (N_18904,N_16636,N_16724);
nor U18905 (N_18905,N_17161,N_17337);
nand U18906 (N_18906,N_16097,N_16167);
nor U18907 (N_18907,N_16711,N_16882);
xnor U18908 (N_18908,N_16791,N_16301);
nor U18909 (N_18909,N_17444,N_17361);
or U18910 (N_18910,N_16699,N_16291);
xnor U18911 (N_18911,N_17393,N_16599);
or U18912 (N_18912,N_17210,N_16287);
nand U18913 (N_18913,N_16399,N_17801);
and U18914 (N_18914,N_17376,N_17780);
nand U18915 (N_18915,N_16376,N_16836);
nand U18916 (N_18916,N_17017,N_16592);
nand U18917 (N_18917,N_16082,N_17687);
and U18918 (N_18918,N_16360,N_17174);
and U18919 (N_18919,N_17151,N_16694);
nand U18920 (N_18920,N_16312,N_16025);
nand U18921 (N_18921,N_17097,N_16768);
xor U18922 (N_18922,N_17012,N_16667);
and U18923 (N_18923,N_17479,N_17976);
nor U18924 (N_18924,N_17937,N_17460);
or U18925 (N_18925,N_16281,N_16919);
nand U18926 (N_18926,N_17981,N_17226);
xor U18927 (N_18927,N_16498,N_16756);
xor U18928 (N_18928,N_16587,N_16614);
and U18929 (N_18929,N_16224,N_16747);
nor U18930 (N_18930,N_17421,N_17962);
nor U18931 (N_18931,N_17350,N_16250);
or U18932 (N_18932,N_17036,N_17797);
and U18933 (N_18933,N_16251,N_16457);
xor U18934 (N_18934,N_17261,N_16080);
nor U18935 (N_18935,N_17202,N_17745);
or U18936 (N_18936,N_16604,N_17018);
and U18937 (N_18937,N_16582,N_17719);
and U18938 (N_18938,N_17799,N_16343);
and U18939 (N_18939,N_17197,N_16208);
nand U18940 (N_18940,N_16955,N_17765);
nand U18941 (N_18941,N_17175,N_16326);
nor U18942 (N_18942,N_17727,N_16773);
nand U18943 (N_18943,N_16572,N_16126);
or U18944 (N_18944,N_17619,N_17728);
xor U18945 (N_18945,N_16418,N_17342);
xor U18946 (N_18946,N_17160,N_16579);
nor U18947 (N_18947,N_17255,N_17064);
xor U18948 (N_18948,N_17482,N_17776);
and U18949 (N_18949,N_17221,N_17811);
nor U18950 (N_18950,N_17348,N_16881);
nand U18951 (N_18951,N_17581,N_16519);
and U18952 (N_18952,N_17437,N_17886);
nand U18953 (N_18953,N_16134,N_16566);
xor U18954 (N_18954,N_16203,N_17784);
nand U18955 (N_18955,N_16430,N_16181);
nand U18956 (N_18956,N_17802,N_16213);
or U18957 (N_18957,N_17677,N_16158);
xnor U18958 (N_18958,N_17326,N_17150);
and U18959 (N_18959,N_16560,N_17848);
xnor U18960 (N_18960,N_16835,N_17260);
or U18961 (N_18961,N_17242,N_17162);
or U18962 (N_18962,N_17224,N_17453);
xor U18963 (N_18963,N_17060,N_17610);
nand U18964 (N_18964,N_17152,N_16639);
and U18965 (N_18965,N_17199,N_16763);
and U18966 (N_18966,N_17763,N_16777);
xnor U18967 (N_18967,N_17452,N_17578);
and U18968 (N_18968,N_16358,N_17125);
nor U18969 (N_18969,N_16131,N_17123);
and U18970 (N_18970,N_17544,N_17014);
xnor U18971 (N_18971,N_17506,N_16184);
nor U18972 (N_18972,N_17536,N_17908);
xnor U18973 (N_18973,N_17441,N_17129);
or U18974 (N_18974,N_16985,N_17623);
xnor U18975 (N_18975,N_17443,N_17382);
xor U18976 (N_18976,N_17766,N_17759);
nand U18977 (N_18977,N_17422,N_17189);
and U18978 (N_18978,N_17883,N_17874);
xnor U18979 (N_18979,N_17604,N_17743);
and U18980 (N_18980,N_17649,N_16098);
xnor U18981 (N_18981,N_17201,N_16630);
nand U18982 (N_18982,N_17091,N_16781);
nand U18983 (N_18983,N_17980,N_17927);
nor U18984 (N_18984,N_17264,N_17665);
nand U18985 (N_18985,N_16798,N_17154);
nor U18986 (N_18986,N_17992,N_16804);
and U18987 (N_18987,N_16412,N_17549);
nand U18988 (N_18988,N_16397,N_17109);
or U18989 (N_18989,N_17531,N_16583);
nor U18990 (N_18990,N_17887,N_16188);
and U18991 (N_18991,N_16146,N_17720);
or U18992 (N_18992,N_17070,N_17840);
nor U18993 (N_18993,N_17200,N_16978);
nand U18994 (N_18994,N_17172,N_17295);
and U18995 (N_18995,N_17928,N_17828);
nor U18996 (N_18996,N_16550,N_16028);
and U18997 (N_18997,N_16873,N_16588);
nand U18998 (N_18998,N_16600,N_17005);
xnor U18999 (N_18999,N_16393,N_16998);
or U19000 (N_19000,N_17940,N_17878);
or U19001 (N_19001,N_17216,N_17992);
nand U19002 (N_19002,N_16265,N_16946);
nor U19003 (N_19003,N_17533,N_16416);
and U19004 (N_19004,N_16075,N_16478);
xor U19005 (N_19005,N_17908,N_16293);
and U19006 (N_19006,N_16748,N_17961);
nor U19007 (N_19007,N_16365,N_16118);
nand U19008 (N_19008,N_16311,N_17455);
and U19009 (N_19009,N_16316,N_16127);
nand U19010 (N_19010,N_17810,N_16514);
xor U19011 (N_19011,N_16613,N_17304);
nor U19012 (N_19012,N_16780,N_17372);
nor U19013 (N_19013,N_16072,N_17838);
and U19014 (N_19014,N_16258,N_17532);
and U19015 (N_19015,N_17851,N_17854);
and U19016 (N_19016,N_17007,N_16293);
or U19017 (N_19017,N_16587,N_16627);
or U19018 (N_19018,N_17562,N_16262);
and U19019 (N_19019,N_16578,N_16321);
or U19020 (N_19020,N_16915,N_17735);
or U19021 (N_19021,N_16236,N_16801);
and U19022 (N_19022,N_17257,N_17293);
nor U19023 (N_19023,N_17418,N_17905);
nand U19024 (N_19024,N_17725,N_16942);
nor U19025 (N_19025,N_16181,N_16734);
nor U19026 (N_19026,N_17432,N_17284);
nor U19027 (N_19027,N_16675,N_16967);
or U19028 (N_19028,N_17728,N_16491);
nor U19029 (N_19029,N_17114,N_17846);
or U19030 (N_19030,N_17780,N_17191);
or U19031 (N_19031,N_16355,N_16706);
or U19032 (N_19032,N_16416,N_16560);
nor U19033 (N_19033,N_17262,N_16616);
nand U19034 (N_19034,N_17382,N_17539);
and U19035 (N_19035,N_16307,N_17734);
and U19036 (N_19036,N_16010,N_17576);
xor U19037 (N_19037,N_17759,N_17007);
or U19038 (N_19038,N_16317,N_16249);
nor U19039 (N_19039,N_17149,N_17102);
nand U19040 (N_19040,N_16496,N_17861);
xor U19041 (N_19041,N_16906,N_16580);
or U19042 (N_19042,N_16374,N_16758);
xnor U19043 (N_19043,N_17101,N_17161);
xor U19044 (N_19044,N_16536,N_16729);
nor U19045 (N_19045,N_16463,N_16439);
nand U19046 (N_19046,N_16099,N_17258);
xor U19047 (N_19047,N_16283,N_16866);
nand U19048 (N_19048,N_17227,N_16644);
xor U19049 (N_19049,N_17778,N_16913);
nand U19050 (N_19050,N_16083,N_17808);
xnor U19051 (N_19051,N_17126,N_16366);
xor U19052 (N_19052,N_16009,N_16114);
nand U19053 (N_19053,N_17142,N_16274);
and U19054 (N_19054,N_17503,N_16804);
nor U19055 (N_19055,N_17958,N_17378);
or U19056 (N_19056,N_17378,N_17994);
and U19057 (N_19057,N_16066,N_16011);
nand U19058 (N_19058,N_17766,N_17806);
or U19059 (N_19059,N_17186,N_16897);
nor U19060 (N_19060,N_17426,N_17283);
nand U19061 (N_19061,N_16220,N_17963);
nand U19062 (N_19062,N_16060,N_17283);
nor U19063 (N_19063,N_16193,N_17903);
nand U19064 (N_19064,N_16047,N_16788);
and U19065 (N_19065,N_16748,N_17672);
xor U19066 (N_19066,N_17325,N_17457);
xnor U19067 (N_19067,N_17284,N_16316);
nand U19068 (N_19068,N_16323,N_16944);
and U19069 (N_19069,N_17824,N_16574);
nand U19070 (N_19070,N_16179,N_17617);
or U19071 (N_19071,N_17387,N_16860);
or U19072 (N_19072,N_16401,N_16706);
xor U19073 (N_19073,N_17635,N_16265);
or U19074 (N_19074,N_16922,N_16633);
nand U19075 (N_19075,N_17084,N_16168);
or U19076 (N_19076,N_17561,N_16518);
nor U19077 (N_19077,N_16026,N_17093);
nor U19078 (N_19078,N_17002,N_17775);
and U19079 (N_19079,N_17269,N_16269);
and U19080 (N_19080,N_17111,N_16953);
and U19081 (N_19081,N_16796,N_17192);
or U19082 (N_19082,N_17546,N_17429);
nor U19083 (N_19083,N_17489,N_16113);
nand U19084 (N_19084,N_17987,N_16163);
xor U19085 (N_19085,N_16555,N_16553);
nand U19086 (N_19086,N_17720,N_16583);
xnor U19087 (N_19087,N_17417,N_16517);
nor U19088 (N_19088,N_16305,N_16930);
nand U19089 (N_19089,N_17149,N_17511);
or U19090 (N_19090,N_17451,N_17231);
nand U19091 (N_19091,N_17136,N_16108);
nand U19092 (N_19092,N_17080,N_16053);
xor U19093 (N_19093,N_16854,N_17951);
xor U19094 (N_19094,N_17382,N_17321);
nor U19095 (N_19095,N_16654,N_16226);
and U19096 (N_19096,N_16727,N_17940);
xor U19097 (N_19097,N_17046,N_17477);
or U19098 (N_19098,N_17381,N_17789);
xnor U19099 (N_19099,N_17962,N_17772);
xor U19100 (N_19100,N_17879,N_16689);
nand U19101 (N_19101,N_16861,N_16491);
or U19102 (N_19102,N_17843,N_16930);
xor U19103 (N_19103,N_17881,N_16631);
xor U19104 (N_19104,N_16016,N_17625);
and U19105 (N_19105,N_17215,N_16331);
or U19106 (N_19106,N_16334,N_16292);
xor U19107 (N_19107,N_17739,N_17566);
xor U19108 (N_19108,N_17488,N_17831);
nand U19109 (N_19109,N_16714,N_17166);
or U19110 (N_19110,N_16348,N_16714);
nand U19111 (N_19111,N_17786,N_16278);
nand U19112 (N_19112,N_16517,N_17618);
or U19113 (N_19113,N_16107,N_17891);
or U19114 (N_19114,N_16762,N_16277);
or U19115 (N_19115,N_17559,N_16924);
nor U19116 (N_19116,N_16131,N_17075);
and U19117 (N_19117,N_17084,N_16255);
or U19118 (N_19118,N_17423,N_16835);
or U19119 (N_19119,N_17759,N_16471);
or U19120 (N_19120,N_17421,N_16886);
or U19121 (N_19121,N_17831,N_17228);
nand U19122 (N_19122,N_16247,N_17300);
xor U19123 (N_19123,N_16887,N_16210);
nand U19124 (N_19124,N_16346,N_16110);
nor U19125 (N_19125,N_16843,N_16359);
nand U19126 (N_19126,N_17297,N_17128);
nand U19127 (N_19127,N_16184,N_16695);
nor U19128 (N_19128,N_17744,N_16071);
or U19129 (N_19129,N_17259,N_16811);
or U19130 (N_19130,N_16452,N_16304);
nand U19131 (N_19131,N_16896,N_17505);
xor U19132 (N_19132,N_16772,N_17415);
and U19133 (N_19133,N_16887,N_17744);
xor U19134 (N_19134,N_17564,N_16070);
nor U19135 (N_19135,N_17927,N_16150);
nor U19136 (N_19136,N_17360,N_16650);
nand U19137 (N_19137,N_16631,N_17638);
and U19138 (N_19138,N_17866,N_16062);
xor U19139 (N_19139,N_16608,N_17556);
xnor U19140 (N_19140,N_17935,N_16621);
or U19141 (N_19141,N_17456,N_17131);
nor U19142 (N_19142,N_17323,N_16321);
xnor U19143 (N_19143,N_16774,N_16964);
nor U19144 (N_19144,N_17733,N_16670);
xnor U19145 (N_19145,N_17564,N_16873);
and U19146 (N_19146,N_16285,N_17515);
or U19147 (N_19147,N_17358,N_16323);
or U19148 (N_19148,N_17904,N_17310);
and U19149 (N_19149,N_17793,N_17525);
and U19150 (N_19150,N_16982,N_16402);
nand U19151 (N_19151,N_16315,N_16863);
nor U19152 (N_19152,N_17928,N_16011);
nor U19153 (N_19153,N_17170,N_16496);
and U19154 (N_19154,N_16986,N_17712);
and U19155 (N_19155,N_16386,N_16844);
nor U19156 (N_19156,N_16211,N_17392);
xor U19157 (N_19157,N_16189,N_16290);
or U19158 (N_19158,N_16752,N_16292);
and U19159 (N_19159,N_17223,N_16904);
or U19160 (N_19160,N_16828,N_17569);
xnor U19161 (N_19161,N_17100,N_17748);
xor U19162 (N_19162,N_16716,N_16249);
nor U19163 (N_19163,N_16347,N_16399);
or U19164 (N_19164,N_16339,N_16485);
nor U19165 (N_19165,N_17814,N_16374);
xor U19166 (N_19166,N_17229,N_16179);
and U19167 (N_19167,N_16422,N_16969);
nor U19168 (N_19168,N_17404,N_16595);
xor U19169 (N_19169,N_17418,N_16997);
and U19170 (N_19170,N_17184,N_16751);
and U19171 (N_19171,N_16838,N_16009);
nor U19172 (N_19172,N_16329,N_17452);
or U19173 (N_19173,N_16764,N_17344);
or U19174 (N_19174,N_16474,N_17607);
nand U19175 (N_19175,N_17432,N_16903);
or U19176 (N_19176,N_16517,N_17950);
or U19177 (N_19177,N_17019,N_17525);
nor U19178 (N_19178,N_16013,N_17431);
nand U19179 (N_19179,N_16607,N_17334);
nor U19180 (N_19180,N_17349,N_16714);
and U19181 (N_19181,N_16330,N_17578);
nor U19182 (N_19182,N_16977,N_17105);
xnor U19183 (N_19183,N_16894,N_16278);
nand U19184 (N_19184,N_16031,N_16248);
nor U19185 (N_19185,N_17500,N_16413);
or U19186 (N_19186,N_16676,N_17453);
nor U19187 (N_19187,N_16392,N_16910);
or U19188 (N_19188,N_16628,N_17261);
and U19189 (N_19189,N_17472,N_16054);
nand U19190 (N_19190,N_17047,N_17408);
and U19191 (N_19191,N_16637,N_17995);
xnor U19192 (N_19192,N_16405,N_16138);
or U19193 (N_19193,N_16587,N_16098);
xnor U19194 (N_19194,N_17243,N_16532);
nand U19195 (N_19195,N_17291,N_16071);
xnor U19196 (N_19196,N_16198,N_16361);
xor U19197 (N_19197,N_16642,N_17134);
nor U19198 (N_19198,N_17468,N_17577);
xor U19199 (N_19199,N_16763,N_16945);
nor U19200 (N_19200,N_17372,N_16598);
nand U19201 (N_19201,N_17813,N_16850);
xnor U19202 (N_19202,N_16293,N_16866);
or U19203 (N_19203,N_16220,N_16499);
xor U19204 (N_19204,N_17025,N_16290);
or U19205 (N_19205,N_17232,N_17125);
or U19206 (N_19206,N_17636,N_16154);
or U19207 (N_19207,N_16832,N_16247);
or U19208 (N_19208,N_17344,N_17147);
nor U19209 (N_19209,N_17087,N_16975);
nor U19210 (N_19210,N_17406,N_17726);
and U19211 (N_19211,N_17825,N_17125);
and U19212 (N_19212,N_16220,N_17892);
nand U19213 (N_19213,N_17667,N_16520);
or U19214 (N_19214,N_17626,N_17788);
nor U19215 (N_19215,N_16227,N_16346);
xor U19216 (N_19216,N_17327,N_16111);
or U19217 (N_19217,N_17956,N_17166);
xor U19218 (N_19218,N_17407,N_16537);
xor U19219 (N_19219,N_17361,N_17246);
and U19220 (N_19220,N_16921,N_17326);
and U19221 (N_19221,N_17623,N_16928);
xnor U19222 (N_19222,N_17248,N_16902);
xor U19223 (N_19223,N_17539,N_17742);
or U19224 (N_19224,N_17280,N_17380);
xnor U19225 (N_19225,N_16223,N_16249);
or U19226 (N_19226,N_17303,N_17215);
and U19227 (N_19227,N_16325,N_16577);
nand U19228 (N_19228,N_17705,N_17505);
xnor U19229 (N_19229,N_17451,N_17393);
or U19230 (N_19230,N_16185,N_17199);
and U19231 (N_19231,N_17235,N_16520);
xor U19232 (N_19232,N_16526,N_17173);
and U19233 (N_19233,N_17037,N_16867);
nor U19234 (N_19234,N_16390,N_17555);
nand U19235 (N_19235,N_17072,N_16067);
nor U19236 (N_19236,N_16070,N_17355);
nand U19237 (N_19237,N_17541,N_17848);
nand U19238 (N_19238,N_16607,N_17324);
xor U19239 (N_19239,N_16289,N_16803);
and U19240 (N_19240,N_16894,N_17672);
xnor U19241 (N_19241,N_16792,N_16020);
nand U19242 (N_19242,N_17158,N_16163);
nor U19243 (N_19243,N_17591,N_17715);
nand U19244 (N_19244,N_16629,N_16547);
xor U19245 (N_19245,N_17173,N_16208);
nor U19246 (N_19246,N_17745,N_16000);
xor U19247 (N_19247,N_17204,N_17643);
nor U19248 (N_19248,N_17681,N_17240);
nand U19249 (N_19249,N_17526,N_17556);
or U19250 (N_19250,N_16624,N_16105);
or U19251 (N_19251,N_16768,N_17370);
and U19252 (N_19252,N_16905,N_16542);
nor U19253 (N_19253,N_16667,N_16155);
nor U19254 (N_19254,N_17057,N_16018);
or U19255 (N_19255,N_17428,N_16517);
nor U19256 (N_19256,N_17129,N_16536);
and U19257 (N_19257,N_17343,N_17703);
nor U19258 (N_19258,N_16654,N_17190);
xor U19259 (N_19259,N_16641,N_17376);
nand U19260 (N_19260,N_17906,N_17372);
nand U19261 (N_19261,N_16756,N_17733);
nor U19262 (N_19262,N_16881,N_17040);
and U19263 (N_19263,N_17472,N_16339);
or U19264 (N_19264,N_16043,N_16964);
xor U19265 (N_19265,N_17672,N_16643);
or U19266 (N_19266,N_17381,N_17888);
nand U19267 (N_19267,N_17720,N_16904);
nor U19268 (N_19268,N_16963,N_17579);
xnor U19269 (N_19269,N_17957,N_17481);
nor U19270 (N_19270,N_17232,N_16222);
nor U19271 (N_19271,N_17390,N_17935);
and U19272 (N_19272,N_16724,N_17961);
nor U19273 (N_19273,N_17098,N_16370);
or U19274 (N_19274,N_16740,N_17521);
xnor U19275 (N_19275,N_16099,N_17040);
nor U19276 (N_19276,N_16797,N_17822);
nand U19277 (N_19277,N_17490,N_16732);
or U19278 (N_19278,N_16993,N_16951);
xor U19279 (N_19279,N_16747,N_16347);
or U19280 (N_19280,N_17147,N_16728);
and U19281 (N_19281,N_16591,N_17690);
nand U19282 (N_19282,N_16866,N_17108);
xor U19283 (N_19283,N_16009,N_16775);
nor U19284 (N_19284,N_17051,N_17571);
and U19285 (N_19285,N_17390,N_16542);
nor U19286 (N_19286,N_17461,N_16848);
and U19287 (N_19287,N_17368,N_16180);
nand U19288 (N_19288,N_16264,N_16283);
nand U19289 (N_19289,N_17532,N_17225);
or U19290 (N_19290,N_17697,N_16476);
or U19291 (N_19291,N_17163,N_16970);
nor U19292 (N_19292,N_16355,N_17178);
nand U19293 (N_19293,N_17590,N_17063);
nor U19294 (N_19294,N_16728,N_16591);
and U19295 (N_19295,N_17959,N_17547);
nand U19296 (N_19296,N_16806,N_17402);
nand U19297 (N_19297,N_16329,N_16585);
or U19298 (N_19298,N_16738,N_17875);
nand U19299 (N_19299,N_16550,N_17856);
xor U19300 (N_19300,N_16413,N_16111);
nand U19301 (N_19301,N_17748,N_16543);
or U19302 (N_19302,N_17388,N_17879);
or U19303 (N_19303,N_17683,N_16936);
nor U19304 (N_19304,N_16379,N_17525);
or U19305 (N_19305,N_17810,N_16161);
xnor U19306 (N_19306,N_16676,N_17256);
or U19307 (N_19307,N_17081,N_16625);
xnor U19308 (N_19308,N_16248,N_17001);
and U19309 (N_19309,N_16642,N_17827);
nor U19310 (N_19310,N_16093,N_17473);
and U19311 (N_19311,N_17165,N_17972);
nor U19312 (N_19312,N_16154,N_17755);
nand U19313 (N_19313,N_17968,N_16981);
and U19314 (N_19314,N_17454,N_16323);
nor U19315 (N_19315,N_17603,N_16790);
xnor U19316 (N_19316,N_17737,N_16869);
and U19317 (N_19317,N_16776,N_16164);
nor U19318 (N_19318,N_17926,N_17469);
nor U19319 (N_19319,N_16244,N_17915);
and U19320 (N_19320,N_17174,N_16160);
nand U19321 (N_19321,N_16286,N_17616);
or U19322 (N_19322,N_17291,N_16843);
and U19323 (N_19323,N_16725,N_17633);
nor U19324 (N_19324,N_17931,N_17935);
and U19325 (N_19325,N_16792,N_17802);
or U19326 (N_19326,N_16154,N_17156);
nand U19327 (N_19327,N_17959,N_16456);
and U19328 (N_19328,N_17838,N_17241);
xnor U19329 (N_19329,N_17646,N_17696);
nand U19330 (N_19330,N_17992,N_17563);
nand U19331 (N_19331,N_16310,N_17888);
or U19332 (N_19332,N_16270,N_16221);
or U19333 (N_19333,N_16650,N_16141);
and U19334 (N_19334,N_17219,N_16891);
and U19335 (N_19335,N_16419,N_17351);
xnor U19336 (N_19336,N_17528,N_17544);
xnor U19337 (N_19337,N_17375,N_16406);
or U19338 (N_19338,N_17653,N_17230);
or U19339 (N_19339,N_16897,N_17473);
or U19340 (N_19340,N_17559,N_16574);
nor U19341 (N_19341,N_16380,N_17124);
nand U19342 (N_19342,N_17640,N_16774);
and U19343 (N_19343,N_17227,N_17551);
nand U19344 (N_19344,N_16994,N_17956);
nor U19345 (N_19345,N_16658,N_16079);
or U19346 (N_19346,N_16036,N_16410);
nand U19347 (N_19347,N_16932,N_16718);
nor U19348 (N_19348,N_16671,N_16895);
nand U19349 (N_19349,N_17949,N_16381);
xor U19350 (N_19350,N_16605,N_17142);
nand U19351 (N_19351,N_16310,N_16705);
xor U19352 (N_19352,N_16455,N_16242);
and U19353 (N_19353,N_16130,N_16887);
nor U19354 (N_19354,N_16044,N_16281);
or U19355 (N_19355,N_17847,N_17617);
or U19356 (N_19356,N_16350,N_16002);
or U19357 (N_19357,N_17016,N_17627);
nand U19358 (N_19358,N_16785,N_17784);
nor U19359 (N_19359,N_17593,N_16867);
nor U19360 (N_19360,N_17636,N_16811);
xor U19361 (N_19361,N_16726,N_16718);
or U19362 (N_19362,N_17688,N_17690);
nand U19363 (N_19363,N_16025,N_17953);
or U19364 (N_19364,N_17153,N_16135);
nand U19365 (N_19365,N_17545,N_17593);
or U19366 (N_19366,N_16834,N_17722);
nand U19367 (N_19367,N_16004,N_17192);
nor U19368 (N_19368,N_16115,N_17605);
or U19369 (N_19369,N_16988,N_17560);
nor U19370 (N_19370,N_16300,N_16555);
or U19371 (N_19371,N_16452,N_16362);
xnor U19372 (N_19372,N_17792,N_17169);
nand U19373 (N_19373,N_17436,N_16360);
nor U19374 (N_19374,N_16759,N_16140);
nand U19375 (N_19375,N_17675,N_16267);
xnor U19376 (N_19376,N_16237,N_16027);
or U19377 (N_19377,N_17261,N_16738);
and U19378 (N_19378,N_16541,N_16815);
and U19379 (N_19379,N_17127,N_16000);
nand U19380 (N_19380,N_16658,N_16037);
or U19381 (N_19381,N_16486,N_17385);
nand U19382 (N_19382,N_16122,N_16187);
and U19383 (N_19383,N_17293,N_17523);
nand U19384 (N_19384,N_17423,N_16874);
nand U19385 (N_19385,N_16891,N_16587);
nor U19386 (N_19386,N_17525,N_17966);
and U19387 (N_19387,N_16056,N_17382);
nand U19388 (N_19388,N_16885,N_16995);
or U19389 (N_19389,N_17152,N_16017);
and U19390 (N_19390,N_17579,N_16713);
or U19391 (N_19391,N_16804,N_17099);
nand U19392 (N_19392,N_17029,N_17097);
xnor U19393 (N_19393,N_17599,N_17031);
and U19394 (N_19394,N_16438,N_17473);
nand U19395 (N_19395,N_17792,N_16499);
and U19396 (N_19396,N_17727,N_16910);
nor U19397 (N_19397,N_16245,N_16178);
and U19398 (N_19398,N_16108,N_17029);
and U19399 (N_19399,N_16571,N_17940);
nor U19400 (N_19400,N_16476,N_17467);
or U19401 (N_19401,N_16642,N_17705);
xnor U19402 (N_19402,N_17272,N_17643);
nor U19403 (N_19403,N_16840,N_17396);
nand U19404 (N_19404,N_17558,N_16687);
nor U19405 (N_19405,N_17846,N_16468);
xor U19406 (N_19406,N_16728,N_16033);
nand U19407 (N_19407,N_16126,N_16031);
nor U19408 (N_19408,N_17253,N_16038);
nand U19409 (N_19409,N_17329,N_17557);
nand U19410 (N_19410,N_17210,N_16641);
or U19411 (N_19411,N_17901,N_17569);
xor U19412 (N_19412,N_17132,N_16113);
nand U19413 (N_19413,N_17513,N_16570);
and U19414 (N_19414,N_17410,N_17161);
or U19415 (N_19415,N_16683,N_16621);
and U19416 (N_19416,N_17714,N_17598);
nor U19417 (N_19417,N_17234,N_17734);
and U19418 (N_19418,N_16119,N_16037);
nand U19419 (N_19419,N_16959,N_16155);
xnor U19420 (N_19420,N_16450,N_16488);
and U19421 (N_19421,N_16785,N_17123);
and U19422 (N_19422,N_16792,N_17068);
xor U19423 (N_19423,N_16136,N_16665);
nor U19424 (N_19424,N_17524,N_16624);
nand U19425 (N_19425,N_16526,N_17969);
nor U19426 (N_19426,N_16471,N_16714);
and U19427 (N_19427,N_17073,N_16638);
or U19428 (N_19428,N_16972,N_17092);
nand U19429 (N_19429,N_17982,N_16887);
and U19430 (N_19430,N_16018,N_16776);
and U19431 (N_19431,N_17974,N_17712);
nand U19432 (N_19432,N_17949,N_17890);
xnor U19433 (N_19433,N_16460,N_16515);
nand U19434 (N_19434,N_17509,N_17069);
nand U19435 (N_19435,N_16752,N_16519);
nand U19436 (N_19436,N_17374,N_17101);
xor U19437 (N_19437,N_16676,N_17671);
or U19438 (N_19438,N_16724,N_16819);
or U19439 (N_19439,N_17137,N_17459);
and U19440 (N_19440,N_17722,N_17073);
nor U19441 (N_19441,N_16793,N_17026);
nand U19442 (N_19442,N_16512,N_16749);
or U19443 (N_19443,N_16134,N_16092);
nand U19444 (N_19444,N_17085,N_17986);
and U19445 (N_19445,N_16231,N_17894);
xnor U19446 (N_19446,N_16069,N_16730);
nand U19447 (N_19447,N_17143,N_17250);
nand U19448 (N_19448,N_16020,N_16184);
and U19449 (N_19449,N_17095,N_17413);
nor U19450 (N_19450,N_17023,N_16200);
and U19451 (N_19451,N_16528,N_16881);
or U19452 (N_19452,N_17180,N_16363);
and U19453 (N_19453,N_16375,N_16821);
or U19454 (N_19454,N_16190,N_16754);
nand U19455 (N_19455,N_16631,N_17240);
and U19456 (N_19456,N_16081,N_16938);
or U19457 (N_19457,N_16178,N_16978);
nand U19458 (N_19458,N_17025,N_17889);
and U19459 (N_19459,N_16060,N_16893);
nand U19460 (N_19460,N_17600,N_16666);
or U19461 (N_19461,N_17744,N_17734);
or U19462 (N_19462,N_17262,N_16597);
nand U19463 (N_19463,N_17820,N_17423);
xnor U19464 (N_19464,N_16286,N_16244);
nor U19465 (N_19465,N_16787,N_17411);
or U19466 (N_19466,N_16050,N_17983);
nand U19467 (N_19467,N_16744,N_16237);
and U19468 (N_19468,N_16510,N_16447);
nor U19469 (N_19469,N_16603,N_17804);
nor U19470 (N_19470,N_16246,N_17801);
nor U19471 (N_19471,N_16152,N_16509);
and U19472 (N_19472,N_17761,N_16262);
nor U19473 (N_19473,N_16641,N_17410);
or U19474 (N_19474,N_17638,N_16732);
xnor U19475 (N_19475,N_16545,N_17094);
xor U19476 (N_19476,N_16222,N_17472);
nor U19477 (N_19477,N_17857,N_17641);
and U19478 (N_19478,N_16993,N_17930);
nand U19479 (N_19479,N_17666,N_16591);
and U19480 (N_19480,N_16601,N_17430);
nor U19481 (N_19481,N_17330,N_16119);
xor U19482 (N_19482,N_17221,N_16322);
xnor U19483 (N_19483,N_17157,N_16459);
or U19484 (N_19484,N_16106,N_16491);
or U19485 (N_19485,N_16492,N_17634);
nand U19486 (N_19486,N_17400,N_16341);
xnor U19487 (N_19487,N_16255,N_16073);
nor U19488 (N_19488,N_17359,N_16574);
or U19489 (N_19489,N_17585,N_16534);
and U19490 (N_19490,N_16808,N_17565);
or U19491 (N_19491,N_16207,N_16824);
xor U19492 (N_19492,N_16599,N_17276);
nor U19493 (N_19493,N_16146,N_16052);
or U19494 (N_19494,N_17774,N_17523);
or U19495 (N_19495,N_17164,N_16374);
xor U19496 (N_19496,N_17522,N_17693);
or U19497 (N_19497,N_16472,N_16389);
nand U19498 (N_19498,N_16335,N_16092);
or U19499 (N_19499,N_16328,N_16538);
xnor U19500 (N_19500,N_16922,N_17403);
and U19501 (N_19501,N_16050,N_17742);
nor U19502 (N_19502,N_16444,N_17250);
nor U19503 (N_19503,N_17191,N_17392);
and U19504 (N_19504,N_16205,N_17189);
and U19505 (N_19505,N_16902,N_16335);
nor U19506 (N_19506,N_17861,N_17949);
nand U19507 (N_19507,N_16687,N_16797);
nor U19508 (N_19508,N_16334,N_17347);
and U19509 (N_19509,N_17787,N_16269);
nor U19510 (N_19510,N_16789,N_17536);
nand U19511 (N_19511,N_17913,N_16158);
and U19512 (N_19512,N_17332,N_17075);
nor U19513 (N_19513,N_17500,N_16892);
nor U19514 (N_19514,N_16308,N_17844);
and U19515 (N_19515,N_17749,N_16046);
and U19516 (N_19516,N_16118,N_16196);
nand U19517 (N_19517,N_16287,N_17660);
xor U19518 (N_19518,N_17860,N_16346);
or U19519 (N_19519,N_17810,N_17664);
nor U19520 (N_19520,N_16802,N_16042);
nor U19521 (N_19521,N_17234,N_17664);
nand U19522 (N_19522,N_16541,N_16141);
or U19523 (N_19523,N_16922,N_16259);
or U19524 (N_19524,N_17703,N_17631);
xor U19525 (N_19525,N_17529,N_16102);
or U19526 (N_19526,N_17719,N_17710);
xnor U19527 (N_19527,N_17156,N_17119);
nor U19528 (N_19528,N_17006,N_16441);
nor U19529 (N_19529,N_17251,N_17024);
xor U19530 (N_19530,N_16325,N_17336);
and U19531 (N_19531,N_17249,N_17798);
and U19532 (N_19532,N_16307,N_17090);
or U19533 (N_19533,N_17447,N_17827);
xnor U19534 (N_19534,N_16755,N_16974);
nand U19535 (N_19535,N_17629,N_17767);
nor U19536 (N_19536,N_16175,N_16774);
nand U19537 (N_19537,N_17774,N_17675);
nor U19538 (N_19538,N_17260,N_17088);
xnor U19539 (N_19539,N_16066,N_17413);
xor U19540 (N_19540,N_16578,N_16940);
or U19541 (N_19541,N_17126,N_16446);
or U19542 (N_19542,N_17239,N_17286);
xnor U19543 (N_19543,N_16081,N_16176);
or U19544 (N_19544,N_16123,N_16263);
and U19545 (N_19545,N_16134,N_17098);
and U19546 (N_19546,N_17682,N_16076);
nand U19547 (N_19547,N_17598,N_16684);
or U19548 (N_19548,N_17691,N_16503);
and U19549 (N_19549,N_17570,N_17487);
xnor U19550 (N_19550,N_16140,N_16659);
nand U19551 (N_19551,N_16212,N_16791);
nor U19552 (N_19552,N_16334,N_16424);
xor U19553 (N_19553,N_16374,N_17944);
nand U19554 (N_19554,N_16630,N_16946);
nor U19555 (N_19555,N_17820,N_17664);
nor U19556 (N_19556,N_16083,N_16032);
nor U19557 (N_19557,N_17691,N_17924);
xor U19558 (N_19558,N_17283,N_16029);
or U19559 (N_19559,N_16785,N_16660);
nand U19560 (N_19560,N_16069,N_17574);
nand U19561 (N_19561,N_17943,N_16833);
xnor U19562 (N_19562,N_16876,N_16620);
or U19563 (N_19563,N_16289,N_16461);
xor U19564 (N_19564,N_16253,N_16596);
xor U19565 (N_19565,N_17768,N_17251);
or U19566 (N_19566,N_17897,N_17533);
and U19567 (N_19567,N_16241,N_17692);
or U19568 (N_19568,N_16003,N_17562);
nand U19569 (N_19569,N_17853,N_17961);
nor U19570 (N_19570,N_16049,N_16609);
xor U19571 (N_19571,N_16897,N_17273);
and U19572 (N_19572,N_17757,N_17896);
or U19573 (N_19573,N_17976,N_16853);
xnor U19574 (N_19574,N_16878,N_17077);
xnor U19575 (N_19575,N_17538,N_17708);
or U19576 (N_19576,N_16154,N_16803);
nand U19577 (N_19577,N_16268,N_16719);
nand U19578 (N_19578,N_17662,N_16477);
xnor U19579 (N_19579,N_17154,N_16811);
xnor U19580 (N_19580,N_17665,N_16033);
and U19581 (N_19581,N_17078,N_16602);
nor U19582 (N_19582,N_17643,N_16590);
or U19583 (N_19583,N_17074,N_16305);
nand U19584 (N_19584,N_16940,N_16599);
xor U19585 (N_19585,N_17778,N_17916);
nor U19586 (N_19586,N_17023,N_17076);
xnor U19587 (N_19587,N_16781,N_16971);
nand U19588 (N_19588,N_17643,N_17398);
xnor U19589 (N_19589,N_17435,N_16381);
nor U19590 (N_19590,N_17067,N_17007);
nand U19591 (N_19591,N_17322,N_16241);
and U19592 (N_19592,N_16067,N_16877);
xnor U19593 (N_19593,N_16272,N_17310);
xor U19594 (N_19594,N_16423,N_17039);
xnor U19595 (N_19595,N_16623,N_17324);
nand U19596 (N_19596,N_17600,N_17779);
nand U19597 (N_19597,N_17141,N_17430);
and U19598 (N_19598,N_16935,N_17365);
nor U19599 (N_19599,N_16571,N_17994);
nor U19600 (N_19600,N_17282,N_16266);
and U19601 (N_19601,N_16825,N_17530);
nand U19602 (N_19602,N_17448,N_17670);
and U19603 (N_19603,N_17160,N_16466);
or U19604 (N_19604,N_16512,N_16437);
nand U19605 (N_19605,N_17719,N_16153);
nand U19606 (N_19606,N_17926,N_17198);
and U19607 (N_19607,N_16410,N_16718);
or U19608 (N_19608,N_16431,N_16487);
and U19609 (N_19609,N_17620,N_17985);
nor U19610 (N_19610,N_17049,N_16197);
nor U19611 (N_19611,N_17222,N_16487);
xor U19612 (N_19612,N_17188,N_17524);
xnor U19613 (N_19613,N_16858,N_16657);
xor U19614 (N_19614,N_16728,N_16376);
and U19615 (N_19615,N_17824,N_17943);
and U19616 (N_19616,N_17846,N_17709);
nor U19617 (N_19617,N_17906,N_17890);
nor U19618 (N_19618,N_16128,N_17986);
nand U19619 (N_19619,N_16612,N_17740);
nor U19620 (N_19620,N_16923,N_16466);
and U19621 (N_19621,N_17284,N_17010);
or U19622 (N_19622,N_16610,N_16705);
and U19623 (N_19623,N_16713,N_17634);
xnor U19624 (N_19624,N_16226,N_17933);
xnor U19625 (N_19625,N_17437,N_16554);
and U19626 (N_19626,N_16358,N_17762);
or U19627 (N_19627,N_16986,N_17784);
and U19628 (N_19628,N_17008,N_17455);
xnor U19629 (N_19629,N_17098,N_16157);
nand U19630 (N_19630,N_16616,N_16326);
and U19631 (N_19631,N_16211,N_16461);
xor U19632 (N_19632,N_16765,N_16039);
nor U19633 (N_19633,N_16978,N_16832);
and U19634 (N_19634,N_17349,N_16101);
and U19635 (N_19635,N_16347,N_16883);
xnor U19636 (N_19636,N_16648,N_17145);
and U19637 (N_19637,N_16390,N_17746);
and U19638 (N_19638,N_16866,N_16521);
nor U19639 (N_19639,N_16320,N_17610);
xor U19640 (N_19640,N_17592,N_16190);
or U19641 (N_19641,N_17447,N_17276);
or U19642 (N_19642,N_16714,N_16139);
or U19643 (N_19643,N_17956,N_16856);
and U19644 (N_19644,N_16037,N_17756);
and U19645 (N_19645,N_17943,N_17907);
and U19646 (N_19646,N_16884,N_17381);
nand U19647 (N_19647,N_16749,N_16675);
nor U19648 (N_19648,N_17558,N_17799);
and U19649 (N_19649,N_16521,N_17497);
and U19650 (N_19650,N_16086,N_16650);
or U19651 (N_19651,N_17647,N_17277);
and U19652 (N_19652,N_16847,N_16934);
xnor U19653 (N_19653,N_16822,N_17537);
and U19654 (N_19654,N_17157,N_17244);
nand U19655 (N_19655,N_16486,N_17225);
nand U19656 (N_19656,N_16791,N_16096);
or U19657 (N_19657,N_16484,N_17978);
or U19658 (N_19658,N_16330,N_16816);
xnor U19659 (N_19659,N_17485,N_17437);
or U19660 (N_19660,N_16198,N_16898);
nor U19661 (N_19661,N_16567,N_17233);
and U19662 (N_19662,N_16316,N_16856);
xnor U19663 (N_19663,N_17388,N_17461);
nand U19664 (N_19664,N_17346,N_17194);
nand U19665 (N_19665,N_16972,N_17018);
or U19666 (N_19666,N_17746,N_16907);
and U19667 (N_19667,N_16164,N_17896);
and U19668 (N_19668,N_17420,N_17122);
and U19669 (N_19669,N_17390,N_16132);
nand U19670 (N_19670,N_16092,N_17802);
or U19671 (N_19671,N_16726,N_17718);
and U19672 (N_19672,N_16957,N_17773);
nor U19673 (N_19673,N_17499,N_17800);
and U19674 (N_19674,N_16302,N_17327);
xor U19675 (N_19675,N_16529,N_16902);
nor U19676 (N_19676,N_17025,N_17586);
and U19677 (N_19677,N_17264,N_17450);
nand U19678 (N_19678,N_17454,N_16614);
nor U19679 (N_19679,N_17313,N_16772);
xor U19680 (N_19680,N_17037,N_17150);
nand U19681 (N_19681,N_16423,N_17216);
nor U19682 (N_19682,N_16991,N_17144);
and U19683 (N_19683,N_17703,N_17512);
nor U19684 (N_19684,N_17732,N_17007);
or U19685 (N_19685,N_17507,N_16836);
nor U19686 (N_19686,N_16681,N_16554);
xnor U19687 (N_19687,N_17989,N_17138);
nand U19688 (N_19688,N_17175,N_17267);
and U19689 (N_19689,N_16719,N_16107);
nand U19690 (N_19690,N_17142,N_16255);
or U19691 (N_19691,N_16251,N_16662);
nand U19692 (N_19692,N_17857,N_16226);
and U19693 (N_19693,N_17000,N_16116);
or U19694 (N_19694,N_17618,N_16355);
nor U19695 (N_19695,N_16043,N_17408);
nor U19696 (N_19696,N_17017,N_16830);
nand U19697 (N_19697,N_17656,N_16365);
nor U19698 (N_19698,N_17274,N_16070);
xnor U19699 (N_19699,N_17275,N_16891);
or U19700 (N_19700,N_17640,N_17520);
nand U19701 (N_19701,N_17313,N_16992);
xor U19702 (N_19702,N_17317,N_16144);
xnor U19703 (N_19703,N_17378,N_17815);
nor U19704 (N_19704,N_17171,N_17270);
or U19705 (N_19705,N_17016,N_17339);
and U19706 (N_19706,N_17502,N_16205);
and U19707 (N_19707,N_17473,N_17111);
xnor U19708 (N_19708,N_17354,N_16921);
xor U19709 (N_19709,N_17174,N_16994);
nor U19710 (N_19710,N_16614,N_16269);
or U19711 (N_19711,N_17483,N_16203);
and U19712 (N_19712,N_16949,N_16988);
and U19713 (N_19713,N_17440,N_16008);
nand U19714 (N_19714,N_17336,N_17575);
nor U19715 (N_19715,N_16365,N_16393);
or U19716 (N_19716,N_16597,N_17348);
nor U19717 (N_19717,N_16647,N_16268);
nor U19718 (N_19718,N_17013,N_16268);
nor U19719 (N_19719,N_17782,N_17371);
nand U19720 (N_19720,N_16923,N_16963);
or U19721 (N_19721,N_16345,N_17726);
and U19722 (N_19722,N_16760,N_16464);
nor U19723 (N_19723,N_17112,N_17812);
nand U19724 (N_19724,N_17385,N_17834);
and U19725 (N_19725,N_16618,N_17737);
nor U19726 (N_19726,N_16896,N_16005);
nand U19727 (N_19727,N_16306,N_17937);
xor U19728 (N_19728,N_16146,N_17544);
xor U19729 (N_19729,N_16565,N_17629);
nand U19730 (N_19730,N_16025,N_16728);
xnor U19731 (N_19731,N_16681,N_17584);
or U19732 (N_19732,N_16323,N_17015);
or U19733 (N_19733,N_16700,N_16729);
xor U19734 (N_19734,N_16588,N_16505);
or U19735 (N_19735,N_17036,N_16806);
nand U19736 (N_19736,N_17474,N_17005);
and U19737 (N_19737,N_17048,N_17018);
or U19738 (N_19738,N_16423,N_16324);
and U19739 (N_19739,N_17192,N_16847);
xor U19740 (N_19740,N_17717,N_16136);
nand U19741 (N_19741,N_16729,N_17340);
and U19742 (N_19742,N_16883,N_16692);
nor U19743 (N_19743,N_17690,N_16511);
nor U19744 (N_19744,N_16347,N_16333);
xnor U19745 (N_19745,N_16304,N_16016);
or U19746 (N_19746,N_17337,N_16506);
xnor U19747 (N_19747,N_17282,N_16005);
xor U19748 (N_19748,N_17157,N_17250);
xnor U19749 (N_19749,N_16389,N_16178);
nor U19750 (N_19750,N_16166,N_17516);
xor U19751 (N_19751,N_16633,N_17530);
nand U19752 (N_19752,N_16753,N_17649);
nand U19753 (N_19753,N_17702,N_16331);
nor U19754 (N_19754,N_16893,N_17203);
nand U19755 (N_19755,N_17315,N_16943);
nand U19756 (N_19756,N_16332,N_16073);
nor U19757 (N_19757,N_17000,N_16093);
or U19758 (N_19758,N_17842,N_17729);
nand U19759 (N_19759,N_17288,N_17713);
or U19760 (N_19760,N_17837,N_16788);
and U19761 (N_19761,N_17294,N_16497);
xor U19762 (N_19762,N_16927,N_16191);
nor U19763 (N_19763,N_17755,N_16113);
or U19764 (N_19764,N_16989,N_17545);
nand U19765 (N_19765,N_17010,N_17845);
or U19766 (N_19766,N_17242,N_16533);
xor U19767 (N_19767,N_16861,N_17860);
nand U19768 (N_19768,N_17370,N_17750);
nor U19769 (N_19769,N_16544,N_17774);
nor U19770 (N_19770,N_16081,N_16254);
xor U19771 (N_19771,N_16888,N_17187);
or U19772 (N_19772,N_17188,N_16319);
nand U19773 (N_19773,N_17736,N_17311);
nand U19774 (N_19774,N_17692,N_16843);
and U19775 (N_19775,N_17419,N_16832);
and U19776 (N_19776,N_16647,N_17862);
nor U19777 (N_19777,N_16253,N_16084);
nand U19778 (N_19778,N_16165,N_17373);
and U19779 (N_19779,N_17946,N_17148);
nand U19780 (N_19780,N_17875,N_17837);
and U19781 (N_19781,N_16221,N_16077);
xor U19782 (N_19782,N_17635,N_16568);
xnor U19783 (N_19783,N_16510,N_17002);
xor U19784 (N_19784,N_16751,N_16424);
or U19785 (N_19785,N_17937,N_17073);
nand U19786 (N_19786,N_17646,N_17588);
xor U19787 (N_19787,N_16468,N_16346);
and U19788 (N_19788,N_17279,N_16903);
or U19789 (N_19789,N_17157,N_16954);
xor U19790 (N_19790,N_17862,N_17579);
nand U19791 (N_19791,N_17198,N_17807);
nand U19792 (N_19792,N_17912,N_17322);
nor U19793 (N_19793,N_16600,N_17806);
and U19794 (N_19794,N_16278,N_17561);
nor U19795 (N_19795,N_17143,N_16190);
nand U19796 (N_19796,N_17133,N_16072);
nor U19797 (N_19797,N_16664,N_16747);
xor U19798 (N_19798,N_17685,N_17626);
nand U19799 (N_19799,N_16837,N_16628);
and U19800 (N_19800,N_16539,N_16501);
xor U19801 (N_19801,N_17257,N_16357);
nand U19802 (N_19802,N_17236,N_16760);
nor U19803 (N_19803,N_17029,N_17173);
nand U19804 (N_19804,N_16537,N_17450);
nor U19805 (N_19805,N_17372,N_16532);
nand U19806 (N_19806,N_16431,N_17647);
nand U19807 (N_19807,N_16286,N_17746);
and U19808 (N_19808,N_17969,N_16585);
and U19809 (N_19809,N_16085,N_16009);
or U19810 (N_19810,N_17852,N_16895);
and U19811 (N_19811,N_17978,N_16042);
xnor U19812 (N_19812,N_17070,N_16467);
or U19813 (N_19813,N_17660,N_16845);
or U19814 (N_19814,N_17351,N_17889);
nand U19815 (N_19815,N_17447,N_16464);
xor U19816 (N_19816,N_16812,N_16893);
nand U19817 (N_19817,N_17015,N_16909);
or U19818 (N_19818,N_16443,N_16359);
nor U19819 (N_19819,N_16089,N_17084);
xnor U19820 (N_19820,N_17043,N_17178);
or U19821 (N_19821,N_17186,N_16578);
xor U19822 (N_19822,N_16643,N_16534);
or U19823 (N_19823,N_16616,N_16622);
and U19824 (N_19824,N_17598,N_16159);
and U19825 (N_19825,N_16204,N_17987);
or U19826 (N_19826,N_17570,N_16188);
xnor U19827 (N_19827,N_17026,N_16205);
nand U19828 (N_19828,N_16180,N_17424);
nor U19829 (N_19829,N_16637,N_16716);
nor U19830 (N_19830,N_16293,N_16784);
and U19831 (N_19831,N_17973,N_17844);
and U19832 (N_19832,N_17574,N_16572);
nand U19833 (N_19833,N_17416,N_16558);
and U19834 (N_19834,N_16179,N_16080);
or U19835 (N_19835,N_17620,N_16312);
nand U19836 (N_19836,N_17607,N_17801);
nand U19837 (N_19837,N_16418,N_16103);
nand U19838 (N_19838,N_16493,N_16169);
xor U19839 (N_19839,N_16641,N_17595);
xor U19840 (N_19840,N_16798,N_16806);
nor U19841 (N_19841,N_17774,N_16335);
or U19842 (N_19842,N_17027,N_16676);
or U19843 (N_19843,N_16462,N_16624);
xor U19844 (N_19844,N_16404,N_17108);
or U19845 (N_19845,N_16789,N_17445);
nand U19846 (N_19846,N_16037,N_17436);
or U19847 (N_19847,N_17071,N_17322);
nor U19848 (N_19848,N_17844,N_17133);
nand U19849 (N_19849,N_16196,N_16430);
or U19850 (N_19850,N_17525,N_17849);
nand U19851 (N_19851,N_16246,N_16985);
nand U19852 (N_19852,N_16014,N_16162);
or U19853 (N_19853,N_16254,N_17142);
xnor U19854 (N_19854,N_16115,N_16293);
nor U19855 (N_19855,N_16338,N_17422);
or U19856 (N_19856,N_17467,N_17637);
nand U19857 (N_19857,N_17622,N_17053);
nand U19858 (N_19858,N_16683,N_17948);
xnor U19859 (N_19859,N_16363,N_16547);
nand U19860 (N_19860,N_16824,N_16261);
and U19861 (N_19861,N_17474,N_17365);
xor U19862 (N_19862,N_16084,N_17001);
and U19863 (N_19863,N_17907,N_17485);
xnor U19864 (N_19864,N_17953,N_17959);
nor U19865 (N_19865,N_16961,N_17388);
or U19866 (N_19866,N_17608,N_17839);
and U19867 (N_19867,N_17279,N_16303);
and U19868 (N_19868,N_16096,N_16369);
nand U19869 (N_19869,N_16071,N_16093);
nor U19870 (N_19870,N_16419,N_17322);
nor U19871 (N_19871,N_17604,N_16773);
nor U19872 (N_19872,N_17251,N_16725);
nand U19873 (N_19873,N_17524,N_17734);
nor U19874 (N_19874,N_16928,N_16058);
nand U19875 (N_19875,N_16714,N_17983);
nand U19876 (N_19876,N_17032,N_17592);
xor U19877 (N_19877,N_16492,N_16177);
xnor U19878 (N_19878,N_17504,N_16154);
or U19879 (N_19879,N_17750,N_16561);
xnor U19880 (N_19880,N_17731,N_17465);
nand U19881 (N_19881,N_16762,N_16010);
xnor U19882 (N_19882,N_16254,N_17875);
nand U19883 (N_19883,N_16102,N_16306);
or U19884 (N_19884,N_16710,N_17585);
and U19885 (N_19885,N_17089,N_17984);
xnor U19886 (N_19886,N_17477,N_17914);
and U19887 (N_19887,N_16722,N_16991);
xnor U19888 (N_19888,N_16230,N_17022);
or U19889 (N_19889,N_16692,N_16687);
xnor U19890 (N_19890,N_16966,N_16084);
and U19891 (N_19891,N_17711,N_17923);
nand U19892 (N_19892,N_17774,N_16568);
nor U19893 (N_19893,N_16167,N_16409);
and U19894 (N_19894,N_17363,N_16495);
and U19895 (N_19895,N_16729,N_16045);
nand U19896 (N_19896,N_17584,N_16163);
nand U19897 (N_19897,N_17497,N_17627);
and U19898 (N_19898,N_16366,N_16979);
nor U19899 (N_19899,N_16420,N_16775);
xnor U19900 (N_19900,N_16751,N_17032);
or U19901 (N_19901,N_17595,N_17562);
nor U19902 (N_19902,N_16562,N_16905);
and U19903 (N_19903,N_17028,N_17959);
nor U19904 (N_19904,N_17700,N_17254);
or U19905 (N_19905,N_17253,N_16694);
and U19906 (N_19906,N_17946,N_17421);
xor U19907 (N_19907,N_16491,N_16162);
and U19908 (N_19908,N_16838,N_16706);
nor U19909 (N_19909,N_16497,N_17637);
or U19910 (N_19910,N_16381,N_17925);
nor U19911 (N_19911,N_17319,N_16050);
and U19912 (N_19912,N_17289,N_16830);
nor U19913 (N_19913,N_17921,N_16390);
and U19914 (N_19914,N_16642,N_17070);
and U19915 (N_19915,N_16958,N_17596);
xor U19916 (N_19916,N_17663,N_16276);
nor U19917 (N_19917,N_17196,N_16698);
nor U19918 (N_19918,N_16491,N_16100);
xnor U19919 (N_19919,N_17253,N_17386);
nand U19920 (N_19920,N_17158,N_16817);
and U19921 (N_19921,N_16689,N_17868);
or U19922 (N_19922,N_17945,N_16798);
xnor U19923 (N_19923,N_17386,N_17657);
or U19924 (N_19924,N_16865,N_17359);
xnor U19925 (N_19925,N_17790,N_16274);
and U19926 (N_19926,N_17553,N_17492);
and U19927 (N_19927,N_16206,N_17735);
xnor U19928 (N_19928,N_16158,N_16139);
and U19929 (N_19929,N_16076,N_17176);
or U19930 (N_19930,N_17781,N_17411);
nand U19931 (N_19931,N_16097,N_16377);
nor U19932 (N_19932,N_17642,N_17477);
or U19933 (N_19933,N_17579,N_17588);
xnor U19934 (N_19934,N_17761,N_16464);
nand U19935 (N_19935,N_16421,N_17332);
xnor U19936 (N_19936,N_17042,N_16522);
nand U19937 (N_19937,N_16737,N_17823);
nor U19938 (N_19938,N_16811,N_17716);
nor U19939 (N_19939,N_16607,N_16437);
xor U19940 (N_19940,N_16524,N_17747);
and U19941 (N_19941,N_17094,N_17410);
nand U19942 (N_19942,N_17162,N_16108);
and U19943 (N_19943,N_17429,N_16691);
nand U19944 (N_19944,N_16210,N_16542);
xor U19945 (N_19945,N_16694,N_16619);
and U19946 (N_19946,N_16263,N_16656);
or U19947 (N_19947,N_17590,N_16116);
and U19948 (N_19948,N_16646,N_17078);
or U19949 (N_19949,N_16327,N_17285);
xnor U19950 (N_19950,N_16538,N_17149);
nand U19951 (N_19951,N_17848,N_16561);
xnor U19952 (N_19952,N_16624,N_16464);
nor U19953 (N_19953,N_17646,N_16590);
nor U19954 (N_19954,N_16232,N_16145);
and U19955 (N_19955,N_17494,N_16935);
or U19956 (N_19956,N_16100,N_17870);
nor U19957 (N_19957,N_17250,N_16057);
nor U19958 (N_19958,N_16609,N_17286);
xor U19959 (N_19959,N_16800,N_16919);
and U19960 (N_19960,N_17931,N_17707);
xnor U19961 (N_19961,N_17753,N_17426);
or U19962 (N_19962,N_17553,N_17162);
nor U19963 (N_19963,N_17986,N_16075);
nand U19964 (N_19964,N_16942,N_16506);
nand U19965 (N_19965,N_16516,N_17661);
or U19966 (N_19966,N_17064,N_16164);
nand U19967 (N_19967,N_16842,N_17339);
nor U19968 (N_19968,N_16771,N_17829);
and U19969 (N_19969,N_16087,N_17416);
and U19970 (N_19970,N_17154,N_17390);
nor U19971 (N_19971,N_16109,N_17916);
and U19972 (N_19972,N_16678,N_16929);
and U19973 (N_19973,N_17271,N_17768);
and U19974 (N_19974,N_17613,N_17177);
xnor U19975 (N_19975,N_16621,N_17862);
xor U19976 (N_19976,N_17140,N_16031);
or U19977 (N_19977,N_17986,N_16144);
nand U19978 (N_19978,N_17225,N_17587);
xnor U19979 (N_19979,N_16823,N_17281);
and U19980 (N_19980,N_17366,N_17161);
nand U19981 (N_19981,N_17551,N_17665);
xnor U19982 (N_19982,N_16210,N_17482);
nand U19983 (N_19983,N_16985,N_17459);
or U19984 (N_19984,N_16658,N_17422);
xor U19985 (N_19985,N_17358,N_16661);
nand U19986 (N_19986,N_17969,N_16271);
nand U19987 (N_19987,N_16217,N_16237);
nor U19988 (N_19988,N_16060,N_17550);
and U19989 (N_19989,N_16755,N_16727);
nor U19990 (N_19990,N_16859,N_16771);
nand U19991 (N_19991,N_16953,N_17101);
or U19992 (N_19992,N_17390,N_16683);
or U19993 (N_19993,N_16421,N_16711);
xnor U19994 (N_19994,N_16996,N_16344);
or U19995 (N_19995,N_17865,N_16242);
xnor U19996 (N_19996,N_16041,N_17380);
and U19997 (N_19997,N_17206,N_16978);
or U19998 (N_19998,N_16571,N_17894);
or U19999 (N_19999,N_17126,N_16602);
and U20000 (N_20000,N_18868,N_18404);
nor U20001 (N_20001,N_18063,N_19189);
and U20002 (N_20002,N_19357,N_19377);
nor U20003 (N_20003,N_19919,N_18183);
and U20004 (N_20004,N_18441,N_19153);
xor U20005 (N_20005,N_18204,N_19121);
and U20006 (N_20006,N_18167,N_19315);
nand U20007 (N_20007,N_19604,N_19943);
nor U20008 (N_20008,N_19055,N_19216);
xnor U20009 (N_20009,N_19209,N_19676);
and U20010 (N_20010,N_19348,N_19924);
xor U20011 (N_20011,N_18541,N_19131);
nor U20012 (N_20012,N_18994,N_18826);
nor U20013 (N_20013,N_18170,N_18087);
nor U20014 (N_20014,N_18844,N_19244);
xnor U20015 (N_20015,N_19561,N_19213);
nor U20016 (N_20016,N_18388,N_19869);
and U20017 (N_20017,N_18394,N_18982);
and U20018 (N_20018,N_19148,N_19436);
and U20019 (N_20019,N_19163,N_19104);
or U20020 (N_20020,N_19840,N_19035);
nor U20021 (N_20021,N_19280,N_19159);
and U20022 (N_20022,N_19015,N_19753);
nand U20023 (N_20023,N_19132,N_18772);
xor U20024 (N_20024,N_19842,N_19651);
nand U20025 (N_20025,N_18535,N_18593);
nor U20026 (N_20026,N_19663,N_18788);
and U20027 (N_20027,N_19766,N_18075);
xor U20028 (N_20028,N_19728,N_18693);
nor U20029 (N_20029,N_19721,N_19633);
xor U20030 (N_20030,N_19788,N_19609);
nand U20031 (N_20031,N_19971,N_19220);
nand U20032 (N_20032,N_18106,N_18780);
xnor U20033 (N_20033,N_19563,N_19374);
nor U20034 (N_20034,N_19022,N_18897);
nor U20035 (N_20035,N_18481,N_18933);
nand U20036 (N_20036,N_19558,N_18948);
nor U20037 (N_20037,N_19725,N_18177);
nor U20038 (N_20038,N_18711,N_19152);
xnor U20039 (N_20039,N_19301,N_19618);
nand U20040 (N_20040,N_19265,N_19960);
or U20041 (N_20041,N_18281,N_19577);
xor U20042 (N_20042,N_19202,N_19020);
and U20043 (N_20043,N_19331,N_19136);
xnor U20044 (N_20044,N_19076,N_18040);
or U20045 (N_20045,N_19901,N_19297);
and U20046 (N_20046,N_19461,N_19142);
nor U20047 (N_20047,N_19729,N_19645);
xnor U20048 (N_20048,N_18910,N_19776);
nor U20049 (N_20049,N_18963,N_18611);
nand U20050 (N_20050,N_19113,N_19895);
and U20051 (N_20051,N_18052,N_18907);
nand U20052 (N_20052,N_19524,N_18280);
nand U20053 (N_20053,N_18960,N_18661);
or U20054 (N_20054,N_19476,N_18520);
or U20055 (N_20055,N_19654,N_18952);
xor U20056 (N_20056,N_18208,N_18721);
nand U20057 (N_20057,N_18483,N_19726);
or U20058 (N_20058,N_18526,N_18327);
or U20059 (N_20059,N_18150,N_19617);
and U20060 (N_20060,N_19748,N_19719);
or U20061 (N_20061,N_19143,N_18207);
and U20062 (N_20062,N_19855,N_18786);
nand U20063 (N_20063,N_18456,N_18572);
and U20064 (N_20064,N_19289,N_18166);
and U20065 (N_20065,N_19079,N_18057);
nand U20066 (N_20066,N_19591,N_18973);
and U20067 (N_20067,N_18013,N_19581);
xnor U20068 (N_20068,N_19211,N_19448);
and U20069 (N_20069,N_18479,N_19046);
nor U20070 (N_20070,N_19320,N_18220);
and U20071 (N_20071,N_18882,N_18002);
nor U20072 (N_20072,N_18333,N_18854);
xnor U20073 (N_20073,N_19481,N_18551);
nand U20074 (N_20074,N_19554,N_19905);
nand U20075 (N_20075,N_19629,N_18161);
nor U20076 (N_20076,N_19829,N_18311);
nor U20077 (N_20077,N_19061,N_18054);
nor U20078 (N_20078,N_19731,N_19797);
and U20079 (N_20079,N_18471,N_19918);
and U20080 (N_20080,N_19162,N_19953);
and U20081 (N_20081,N_18127,N_18368);
or U20082 (N_20082,N_19077,N_19067);
nand U20083 (N_20083,N_19050,N_18128);
or U20084 (N_20084,N_19590,N_18046);
nor U20085 (N_20085,N_18188,N_18294);
xor U20086 (N_20086,N_19307,N_19816);
and U20087 (N_20087,N_18930,N_19112);
nand U20088 (N_20088,N_19866,N_18631);
nand U20089 (N_20089,N_18009,N_19045);
or U20090 (N_20090,N_18972,N_19096);
nor U20091 (N_20091,N_19780,N_19459);
or U20092 (N_20092,N_19026,N_19256);
xnor U20093 (N_20093,N_19553,N_19527);
or U20094 (N_20094,N_18752,N_18407);
nand U20095 (N_20095,N_19120,N_18084);
xor U20096 (N_20096,N_18648,N_18888);
xor U20097 (N_20097,N_19469,N_18286);
and U20098 (N_20098,N_19942,N_18676);
xnor U20099 (N_20099,N_18640,N_18097);
nand U20100 (N_20100,N_18793,N_18146);
nand U20101 (N_20101,N_19087,N_18737);
nand U20102 (N_20102,N_18011,N_18957);
xor U20103 (N_20103,N_18026,N_18397);
or U20104 (N_20104,N_19705,N_18937);
or U20105 (N_20105,N_18792,N_18812);
nor U20106 (N_20106,N_19360,N_18839);
xor U20107 (N_20107,N_19813,N_19212);
or U20108 (N_20108,N_19048,N_18119);
xnor U20109 (N_20109,N_18382,N_19182);
xnor U20110 (N_20110,N_19976,N_19123);
nand U20111 (N_20111,N_19779,N_18134);
nor U20112 (N_20112,N_18914,N_18159);
xor U20113 (N_20113,N_18513,N_18978);
nand U20114 (N_20114,N_19820,N_19992);
nand U20115 (N_20115,N_18224,N_18408);
xnor U20116 (N_20116,N_19327,N_18303);
xnor U20117 (N_20117,N_19007,N_19827);
or U20118 (N_20118,N_19785,N_18453);
nor U20119 (N_20119,N_19429,N_18396);
xor U20120 (N_20120,N_18024,N_19004);
xnor U20121 (N_20121,N_19513,N_19756);
or U20122 (N_20122,N_19997,N_18015);
nor U20123 (N_20123,N_18317,N_18504);
nand U20124 (N_20124,N_19266,N_19303);
or U20125 (N_20125,N_19125,N_19199);
and U20126 (N_20126,N_19023,N_18964);
or U20127 (N_20127,N_18925,N_18626);
nor U20128 (N_20128,N_18210,N_18810);
nor U20129 (N_20129,N_19847,N_18262);
nand U20130 (N_20130,N_18216,N_19296);
nand U20131 (N_20131,N_18918,N_18472);
xnor U20132 (N_20132,N_18831,N_18320);
and U20133 (N_20133,N_18450,N_19789);
or U20134 (N_20134,N_19340,N_18719);
or U20135 (N_20135,N_19305,N_19547);
and U20136 (N_20136,N_19945,N_19674);
xnor U20137 (N_20137,N_19947,N_19562);
and U20138 (N_20138,N_18527,N_18860);
xor U20139 (N_20139,N_18079,N_19958);
and U20140 (N_20140,N_19188,N_18496);
nor U20141 (N_20141,N_18385,N_18427);
nor U20142 (N_20142,N_19065,N_19767);
nand U20143 (N_20143,N_19759,N_18096);
and U20144 (N_20144,N_18039,N_18044);
or U20145 (N_20145,N_19086,N_18098);
and U20146 (N_20146,N_19453,N_18981);
xnor U20147 (N_20147,N_18567,N_19402);
nor U20148 (N_20148,N_18126,N_18085);
or U20149 (N_20149,N_19528,N_18628);
and U20150 (N_20150,N_19846,N_18494);
or U20151 (N_20151,N_19187,N_19423);
xnor U20152 (N_20152,N_19384,N_18765);
nor U20153 (N_20153,N_19106,N_18191);
and U20154 (N_20154,N_19929,N_19304);
nand U20155 (N_20155,N_19990,N_19183);
or U20156 (N_20156,N_18345,N_18244);
and U20157 (N_20157,N_19248,N_19276);
nand U20158 (N_20158,N_18474,N_18668);
and U20159 (N_20159,N_18423,N_19295);
and U20160 (N_20160,N_18185,N_19229);
or U20161 (N_20161,N_19956,N_18334);
nand U20162 (N_20162,N_19603,N_18139);
nor U20163 (N_20163,N_18381,N_18199);
and U20164 (N_20164,N_18068,N_19412);
or U20165 (N_20165,N_18832,N_19791);
or U20166 (N_20166,N_18885,N_18708);
nor U20167 (N_20167,N_18621,N_18258);
and U20168 (N_20168,N_19578,N_18563);
and U20169 (N_20169,N_18249,N_19251);
nand U20170 (N_20170,N_19105,N_18393);
xnor U20171 (N_20171,N_19530,N_18947);
nor U20172 (N_20172,N_19777,N_19405);
nor U20173 (N_20173,N_19963,N_19675);
and U20174 (N_20174,N_19806,N_19477);
nand U20175 (N_20175,N_18148,N_18919);
xor U20176 (N_20176,N_18598,N_18218);
or U20177 (N_20177,N_19443,N_19544);
nand U20178 (N_20178,N_18709,N_18614);
nor U20179 (N_20179,N_18715,N_19566);
and U20180 (N_20180,N_19854,N_18647);
nand U20181 (N_20181,N_18547,N_18966);
and U20182 (N_20182,N_18997,N_19636);
nand U20183 (N_20183,N_19912,N_18877);
xor U20184 (N_20184,N_18935,N_18587);
nor U20185 (N_20185,N_19907,N_18739);
and U20186 (N_20186,N_18798,N_19385);
or U20187 (N_20187,N_19630,N_18817);
xor U20188 (N_20188,N_19100,N_19422);
nand U20189 (N_20189,N_19972,N_18078);
nor U20190 (N_20190,N_18617,N_19040);
or U20191 (N_20191,N_19093,N_19964);
nor U20192 (N_20192,N_18946,N_18880);
nor U20193 (N_20193,N_18705,N_18510);
or U20194 (N_20194,N_18575,N_18319);
or U20195 (N_20195,N_19946,N_18559);
and U20196 (N_20196,N_18645,N_19393);
or U20197 (N_20197,N_19445,N_19730);
xnor U20198 (N_20198,N_18515,N_18686);
nor U20199 (N_20199,N_19580,N_19804);
or U20200 (N_20200,N_18646,N_19338);
xor U20201 (N_20201,N_18665,N_19696);
xnor U20202 (N_20202,N_18245,N_18770);
nand U20203 (N_20203,N_18895,N_19662);
or U20204 (N_20204,N_19955,N_18321);
xor U20205 (N_20205,N_19710,N_19814);
and U20206 (N_20206,N_18934,N_19667);
or U20207 (N_20207,N_19999,N_18901);
or U20208 (N_20208,N_18414,N_18767);
and U20209 (N_20209,N_18082,N_19049);
or U20210 (N_20210,N_18499,N_19287);
nor U20211 (N_20211,N_18996,N_19416);
or U20212 (N_20212,N_19574,N_18674);
nand U20213 (N_20213,N_18833,N_18346);
xor U20214 (N_20214,N_18279,N_18552);
nor U20215 (N_20215,N_18763,N_19966);
and U20216 (N_20216,N_19682,N_18361);
nand U20217 (N_20217,N_19382,N_18400);
and U20218 (N_20218,N_18523,N_19885);
nand U20219 (N_20219,N_19364,N_18487);
and U20220 (N_20220,N_19775,N_19889);
or U20221 (N_20221,N_19826,N_18958);
or U20222 (N_20222,N_18736,N_18256);
xnor U20223 (N_20223,N_18603,N_19157);
nor U20224 (N_20224,N_19118,N_18298);
nor U20225 (N_20225,N_19768,N_18250);
or U20226 (N_20226,N_18909,N_19463);
or U20227 (N_20227,N_18942,N_19134);
or U20228 (N_20228,N_18500,N_19832);
xor U20229 (N_20229,N_18790,N_19986);
xnor U20230 (N_20230,N_19551,N_19274);
or U20231 (N_20231,N_18461,N_19882);
or U20232 (N_20232,N_18517,N_18025);
or U20233 (N_20233,N_19738,N_18519);
nand U20234 (N_20234,N_18858,N_19160);
nor U20235 (N_20235,N_18991,N_18437);
xor U20236 (N_20236,N_19593,N_18666);
and U20237 (N_20237,N_19127,N_19559);
xnor U20238 (N_20238,N_19088,N_18373);
or U20239 (N_20239,N_18440,N_18089);
and U20240 (N_20240,N_18112,N_18350);
and U20241 (N_20241,N_19631,N_18124);
nand U20242 (N_20242,N_19601,N_19568);
or U20243 (N_20243,N_18444,N_18337);
and U20244 (N_20244,N_19746,N_19458);
and U20245 (N_20245,N_18660,N_19437);
or U20246 (N_20246,N_19899,N_19720);
nand U20247 (N_20247,N_18446,N_19491);
and U20248 (N_20248,N_18168,N_18105);
xnor U20249 (N_20249,N_18067,N_19115);
nand U20250 (N_20250,N_18384,N_19242);
and U20251 (N_20251,N_18092,N_18390);
or U20252 (N_20252,N_18564,N_18402);
nor U20253 (N_20253,N_19383,N_19981);
and U20254 (N_20254,N_19390,N_18181);
nor U20255 (N_20255,N_18584,N_19008);
and U20256 (N_20256,N_19786,N_19692);
and U20257 (N_20257,N_18622,N_18269);
nand U20258 (N_20258,N_19537,N_18612);
and U20259 (N_20259,N_18042,N_18050);
xnor U20260 (N_20260,N_19161,N_19937);
nor U20261 (N_20261,N_19170,N_19980);
nand U20262 (N_20262,N_19039,N_19736);
xnor U20263 (N_20263,N_18623,N_18031);
and U20264 (N_20264,N_19498,N_19688);
xor U20265 (N_20265,N_18338,N_19896);
xor U20266 (N_20266,N_19397,N_19614);
nor U20267 (N_20267,N_19197,N_18689);
nor U20268 (N_20268,N_19910,N_19925);
and U20269 (N_20269,N_19515,N_18302);
xnor U20270 (N_20270,N_19583,N_19246);
nor U20271 (N_20271,N_19613,N_19119);
xnor U20272 (N_20272,N_19927,N_18577);
or U20273 (N_20273,N_19932,N_19703);
or U20274 (N_20274,N_18690,N_19595);
nor U20275 (N_20275,N_19582,N_19169);
xnor U20276 (N_20276,N_18071,N_18549);
or U20277 (N_20277,N_18945,N_18620);
and U20278 (N_20278,N_18787,N_19054);
or U20279 (N_20279,N_18634,N_19316);
and U20280 (N_20280,N_19363,N_19350);
xor U20281 (N_20281,N_18743,N_19634);
or U20282 (N_20282,N_18399,N_18285);
and U20283 (N_20283,N_18475,N_18682);
and U20284 (N_20284,N_19933,N_19478);
and U20285 (N_20285,N_19761,N_19178);
or U20286 (N_20286,N_19407,N_18953);
nor U20287 (N_20287,N_18016,N_18331);
nor U20288 (N_20288,N_19347,N_19455);
xnor U20289 (N_20289,N_18458,N_18114);
or U20290 (N_20290,N_19438,N_19639);
xor U20291 (N_20291,N_18506,N_19749);
nor U20292 (N_20292,N_18247,N_19569);
xnor U20293 (N_20293,N_19998,N_18955);
and U20294 (N_20294,N_18902,N_18041);
nand U20295 (N_20295,N_19424,N_18539);
or U20296 (N_20296,N_19668,N_18136);
nor U20297 (N_20297,N_19260,N_18217);
nand U20298 (N_20298,N_19264,N_19179);
xor U20299 (N_20299,N_18169,N_18903);
or U20300 (N_20300,N_19712,N_19754);
nand U20301 (N_20301,N_19403,N_19611);
or U20302 (N_20302,N_19859,N_18211);
xor U20303 (N_20303,N_19091,N_19800);
and U20304 (N_20304,N_18132,N_18196);
and U20305 (N_20305,N_19865,N_18176);
nand U20306 (N_20306,N_19095,N_18702);
or U20307 (N_20307,N_18429,N_19967);
nand U20308 (N_20308,N_18275,N_18754);
xor U20309 (N_20309,N_19074,N_18744);
nand U20310 (N_20310,N_18943,N_19241);
xnor U20311 (N_20311,N_19965,N_19042);
nand U20312 (N_20312,N_19223,N_18284);
xor U20313 (N_20313,N_19334,N_18123);
xnor U20314 (N_20314,N_19312,N_18579);
and U20315 (N_20315,N_19394,N_18581);
xor U20316 (N_20316,N_19451,N_19745);
nand U20317 (N_20317,N_18491,N_18649);
nor U20318 (N_20318,N_19621,N_19339);
xnor U20319 (N_20319,N_19520,N_18894);
xor U20320 (N_20320,N_19158,N_19870);
xnor U20321 (N_20321,N_19669,N_18795);
xnor U20322 (N_20322,N_18929,N_18254);
nor U20323 (N_20323,N_19763,N_19573);
and U20324 (N_20324,N_19253,N_18264);
or U20325 (N_20325,N_18814,N_18799);
nor U20326 (N_20326,N_18435,N_18460);
and U20327 (N_20327,N_19322,N_19534);
xor U20328 (N_20328,N_19431,N_19683);
and U20329 (N_20329,N_18422,N_18234);
and U20330 (N_20330,N_19979,N_19092);
and U20331 (N_20331,N_18652,N_19864);
nor U20332 (N_20332,N_18347,N_18323);
xnor U20333 (N_20333,N_19625,N_18418);
nor U20334 (N_20334,N_18706,N_19129);
or U20335 (N_20335,N_18111,N_18724);
and U20336 (N_20336,N_18887,N_18490);
or U20337 (N_20337,N_18202,N_18687);
nand U20338 (N_20338,N_18241,N_18508);
nand U20339 (N_20339,N_18349,N_18941);
or U20340 (N_20340,N_19888,N_18876);
and U20341 (N_20341,N_19677,N_18488);
xor U20342 (N_20342,N_18379,N_18029);
and U20343 (N_20343,N_19516,N_18805);
and U20344 (N_20344,N_19641,N_18610);
xnor U20345 (N_20345,N_19219,N_19724);
nor U20346 (N_20346,N_18650,N_18825);
xor U20347 (N_20347,N_19444,N_18701);
nand U20348 (N_20348,N_18354,N_18670);
and U20349 (N_20349,N_18607,N_18525);
or U20350 (N_20350,N_18365,N_19281);
or U20351 (N_20351,N_19485,N_18766);
nand U20352 (N_20352,N_18073,N_18273);
nand U20353 (N_20353,N_18055,N_19030);
nor U20354 (N_20354,N_19466,N_19743);
nand U20355 (N_20355,N_18533,N_19540);
xor U20356 (N_20356,N_18228,N_19319);
xor U20357 (N_20357,N_19146,N_19576);
or U20358 (N_20358,N_19679,N_19156);
and U20359 (N_20359,N_19388,N_18803);
and U20360 (N_20360,N_18233,N_19906);
xor U20361 (N_20361,N_19757,N_18624);
and U20362 (N_20362,N_19037,N_19311);
or U20363 (N_20363,N_19329,N_19435);
nand U20364 (N_20364,N_19313,N_19849);
xor U20365 (N_20365,N_18027,N_19068);
xnor U20366 (N_20366,N_18608,N_19411);
nand U20367 (N_20367,N_19828,N_18900);
or U20368 (N_20368,N_18434,N_18424);
or U20369 (N_20369,N_18184,N_18147);
nor U20370 (N_20370,N_18299,N_18657);
nor U20371 (N_20371,N_18113,N_19509);
nor U20372 (N_20372,N_19765,N_18033);
or U20373 (N_20373,N_18443,N_19542);
xnor U20374 (N_20374,N_19860,N_18118);
and U20375 (N_20375,N_18703,N_19492);
or U20376 (N_20376,N_18751,N_19508);
nor U20377 (N_20377,N_19755,N_18242);
xnor U20378 (N_20378,N_19543,N_19588);
xor U20379 (N_20379,N_18229,N_18616);
nand U20380 (N_20380,N_18100,N_19911);
nand U20381 (N_20381,N_19367,N_19273);
or U20382 (N_20382,N_19151,N_18305);
and U20383 (N_20383,N_18681,N_18420);
nand U20384 (N_20384,N_19505,N_18197);
and U20385 (N_20385,N_19016,N_18753);
and U20386 (N_20386,N_19701,N_18821);
nor U20387 (N_20387,N_18238,N_18664);
nor U20388 (N_20388,N_18728,N_18516);
or U20389 (N_20389,N_18130,N_18369);
nand U20390 (N_20390,N_18153,N_19380);
and U20391 (N_20391,N_19839,N_19936);
and U20392 (N_20392,N_19570,N_19638);
nand U20393 (N_20393,N_18590,N_19939);
nor U20394 (N_20394,N_19231,N_19805);
or U20395 (N_20395,N_18090,N_18193);
xor U20396 (N_20396,N_19880,N_19333);
nand U20397 (N_20397,N_18975,N_18117);
or U20398 (N_20398,N_18142,N_18095);
nand U20399 (N_20399,N_18292,N_19984);
or U20400 (N_20400,N_18066,N_18149);
or U20401 (N_20401,N_19970,N_19531);
xor U20402 (N_20402,N_19934,N_18988);
xnor U20403 (N_20403,N_19834,N_19200);
or U20404 (N_20404,N_18749,N_18309);
nor U20405 (N_20405,N_18034,N_18362);
nor U20406 (N_20406,N_19195,N_18008);
or U20407 (N_20407,N_18047,N_18524);
nand U20408 (N_20408,N_18398,N_18746);
and U20409 (N_20409,N_19019,N_18058);
or U20410 (N_20410,N_19954,N_18174);
nor U20411 (N_20411,N_19815,N_18561);
nor U20412 (N_20412,N_18061,N_18679);
nor U20413 (N_20413,N_18760,N_19798);
or U20414 (N_20414,N_19973,N_19841);
nand U20415 (N_20415,N_19252,N_19747);
nor U20416 (N_20416,N_18014,N_18389);
xor U20417 (N_20417,N_18849,N_19949);
xor U20418 (N_20418,N_19099,N_19326);
nand U20419 (N_20419,N_19191,N_18954);
xor U20420 (N_20420,N_18949,N_18846);
nor U20421 (N_20421,N_19270,N_18023);
or U20422 (N_20422,N_19109,N_18921);
xor U20423 (N_20423,N_18619,N_19519);
xor U20424 (N_20424,N_19005,N_19982);
and U20425 (N_20425,N_19318,N_19894);
and U20426 (N_20426,N_18195,N_19698);
xor U20427 (N_20427,N_19472,N_19400);
or U20428 (N_20428,N_18053,N_18295);
nand U20429 (N_20429,N_18554,N_18036);
nand U20430 (N_20430,N_18406,N_19552);
nand U20431 (N_20431,N_19389,N_18121);
nor U20432 (N_20432,N_18722,N_18392);
xor U20433 (N_20433,N_18951,N_19468);
and U20434 (N_20434,N_19186,N_19632);
nor U20435 (N_20435,N_19361,N_19454);
and U20436 (N_20436,N_19664,N_18571);
nand U20437 (N_20437,N_19830,N_18695);
and U20438 (N_20438,N_18143,N_18223);
or U20439 (N_20439,N_18872,N_19752);
or U20440 (N_20440,N_19103,N_19369);
xnor U20441 (N_20441,N_18120,N_18125);
nor U20442 (N_20442,N_18530,N_19793);
nor U20443 (N_20443,N_19494,N_18971);
nand U20444 (N_20444,N_19233,N_18932);
nor U20445 (N_20445,N_18529,N_18357);
nand U20446 (N_20446,N_19951,N_19072);
xnor U20447 (N_20447,N_18538,N_18940);
nor U20448 (N_20448,N_18864,N_18822);
or U20449 (N_20449,N_19822,N_18629);
xor U20450 (N_20450,N_19130,N_19332);
or U20451 (N_20451,N_18696,N_19323);
and U20452 (N_20452,N_18246,N_18771);
nor U20453 (N_20453,N_19330,N_18837);
or U20454 (N_20454,N_19300,N_18534);
nand U20455 (N_20455,N_19473,N_18080);
xor U20456 (N_20456,N_19877,N_18847);
or U20457 (N_20457,N_19717,N_18778);
or U20458 (N_20458,N_19760,N_19047);
or U20459 (N_20459,N_18677,N_18578);
or U20460 (N_20460,N_19395,N_18678);
or U20461 (N_20461,N_18099,N_19575);
nor U20462 (N_20462,N_19439,N_19011);
and U20463 (N_20463,N_18521,N_18824);
or U20464 (N_20464,N_19950,N_19009);
or U20465 (N_20465,N_19298,N_19107);
nand U20466 (N_20466,N_19607,N_19511);
nand U20467 (N_20467,N_18905,N_19837);
nand U20468 (N_20468,N_18540,N_19602);
nor U20469 (N_20469,N_18162,N_19781);
nor U20470 (N_20470,N_19057,N_18758);
xnor U20471 (N_20471,N_19628,N_19886);
nand U20472 (N_20472,N_18796,N_18301);
xnor U20473 (N_20473,N_18859,N_18409);
nand U20474 (N_20474,N_19584,N_18818);
xnor U20475 (N_20475,N_19802,N_18278);
nor U20476 (N_20476,N_19051,N_19337);
nor U20477 (N_20477,N_18850,N_18038);
nand U20478 (N_20478,N_19764,N_18155);
or U20479 (N_20479,N_19887,N_18899);
nor U20480 (N_20480,N_18447,N_18733);
or U20481 (N_20481,N_19379,N_19640);
nand U20482 (N_20482,N_19487,N_18465);
nand U20483 (N_20483,N_18003,N_19892);
and U20484 (N_20484,N_18801,N_18802);
or U20485 (N_20485,N_18852,N_19240);
or U20486 (N_20486,N_19139,N_19867);
and U20487 (N_20487,N_18315,N_19672);
nor U20488 (N_20488,N_19401,N_18353);
or U20489 (N_20489,N_18293,N_19145);
nand U20490 (N_20490,N_18820,N_18727);
or U20491 (N_20491,N_18830,N_19184);
nor U20492 (N_20492,N_18944,N_19975);
xor U20493 (N_20493,N_18720,N_19450);
nand U20494 (N_20494,N_19643,N_19938);
nand U20495 (N_20495,N_18144,N_19483);
nor U20496 (N_20496,N_19741,N_19824);
nor U20497 (N_20497,N_19456,N_19655);
nor U20498 (N_20498,N_18187,N_18667);
nand U20499 (N_20499,N_18339,N_18742);
and U20500 (N_20500,N_18175,N_19852);
nor U20501 (N_20501,N_19670,N_19387);
nor U20502 (N_20502,N_18477,N_18137);
or U20503 (N_20503,N_18342,N_18757);
and U20504 (N_20504,N_19166,N_18922);
and U20505 (N_20505,N_19522,N_18276);
nand U20506 (N_20506,N_19174,N_18359);
nor U20507 (N_20507,N_18005,N_19606);
nand U20508 (N_20508,N_19644,N_19546);
xnor U20509 (N_20509,N_18747,N_19038);
and U20510 (N_20510,N_18848,N_18138);
nor U20511 (N_20511,N_18340,N_19708);
and U20512 (N_20512,N_18669,N_19060);
nand U20513 (N_20513,N_19545,N_18020);
nor U20514 (N_20514,N_18378,N_19321);
nor U20515 (N_20515,N_18904,N_18512);
or U20516 (N_20516,N_19373,N_19267);
nand U20517 (N_20517,N_19269,N_19495);
xor U20518 (N_20518,N_18920,N_18289);
and U20519 (N_20519,N_19883,N_18486);
nand U20520 (N_20520,N_18088,N_18001);
and U20521 (N_20521,N_19714,N_18683);
xor U20522 (N_20522,N_18692,N_18738);
and U20523 (N_20523,N_19926,N_19902);
nand U20524 (N_20524,N_19490,N_18697);
and U20525 (N_20525,N_19836,N_19921);
xor U20526 (N_20526,N_19723,N_18186);
and U20527 (N_20527,N_19758,N_19996);
or U20528 (N_20528,N_18680,N_19245);
nor U20529 (N_20529,N_19001,N_18939);
or U20530 (N_20530,N_19850,N_19176);
nand U20531 (N_20531,N_18635,N_19623);
or U20532 (N_20532,N_18135,N_18641);
or U20533 (N_20533,N_18253,N_18566);
and U20534 (N_20534,N_18454,N_18898);
nand U20535 (N_20535,N_19175,N_18545);
and U20536 (N_20536,N_18656,N_19352);
xor U20537 (N_20537,N_18358,N_19908);
nor U20538 (N_20538,N_18808,N_19795);
and U20539 (N_20539,N_18252,N_18430);
nor U20540 (N_20540,N_19263,N_19154);
and U20541 (N_20541,N_19711,N_18049);
nand U20542 (N_20542,N_18959,N_18700);
nand U20543 (N_20543,N_19961,N_18511);
or U20544 (N_20544,N_18428,N_18606);
nand U20545 (N_20545,N_18355,N_18268);
and U20546 (N_20546,N_19235,N_19727);
nor U20547 (N_20547,N_19881,N_19697);
xor U20548 (N_20548,N_18102,N_18911);
or U20549 (N_20549,N_19108,N_19126);
or U20550 (N_20550,N_19733,N_18028);
xnor U20551 (N_20551,N_18867,N_19831);
and U20552 (N_20552,N_18694,N_19594);
nor U20553 (N_20553,N_19567,N_18573);
or U20554 (N_20554,N_19681,N_19739);
and U20555 (N_20555,N_18007,N_18857);
and U20556 (N_20556,N_19036,N_19482);
nor U20557 (N_20557,N_19598,N_19735);
xor U20558 (N_20558,N_18596,N_19722);
nor U20559 (N_20559,N_18189,N_18531);
xnor U20560 (N_20560,N_19770,N_18591);
nand U20561 (N_20561,N_18615,N_18889);
xnor U20562 (N_20562,N_18734,N_19003);
nand U20563 (N_20563,N_18870,N_19336);
or U20564 (N_20564,N_19230,N_19294);
nor U20565 (N_20565,N_18618,N_18190);
nor U20566 (N_20566,N_18260,N_18426);
or U20567 (N_20567,N_19426,N_19610);
or U20568 (N_20568,N_18783,N_19507);
and U20569 (N_20569,N_19657,N_19155);
and U20570 (N_20570,N_18449,N_18663);
xor U20571 (N_20571,N_18784,N_18809);
and U20572 (N_20572,N_18230,N_19597);
nor U20573 (N_20573,N_18077,N_19916);
nor U20574 (N_20574,N_18731,N_18764);
nor U20575 (N_20575,N_18048,N_19787);
nand U20576 (N_20576,N_19133,N_19532);
xnor U20577 (N_20577,N_19278,N_19440);
nand U20578 (N_20578,N_18562,N_18827);
xor U20579 (N_20579,N_19658,N_18755);
or U20580 (N_20580,N_18726,N_19744);
nand U20581 (N_20581,N_19599,N_19053);
nand U20582 (N_20582,N_18201,N_19066);
or U20583 (N_20583,N_19917,N_18655);
and U20584 (N_20584,N_18432,N_19441);
and U20585 (N_20585,N_19396,N_19349);
nor U20586 (N_20586,N_19417,N_18891);
xnor U20587 (N_20587,N_18936,N_18745);
nor U20588 (N_20588,N_18021,N_18171);
nand U20589 (N_20589,N_18698,N_19432);
and U20590 (N_20590,N_19879,N_19168);
xnor U20591 (N_20591,N_18917,N_18732);
nor U20592 (N_20592,N_18987,N_19706);
nor U20593 (N_20593,N_18324,N_19328);
nand U20594 (N_20594,N_19094,N_18503);
nand U20595 (N_20595,N_18962,N_19234);
and U20596 (N_20596,N_18462,N_19434);
nand U20597 (N_20597,N_19283,N_19605);
and U20598 (N_20598,N_19271,N_19488);
nand U20599 (N_20599,N_18865,N_18270);
or U20600 (N_20600,N_19693,N_19968);
xor U20601 (N_20601,N_19557,N_19923);
nand U20602 (N_20602,N_19844,N_19056);
or U20603 (N_20603,N_18627,N_19272);
xnor U20604 (N_20604,N_19533,N_19541);
or U20605 (N_20605,N_19351,N_19974);
or U20606 (N_20606,N_19616,N_19034);
nor U20607 (N_20607,N_18967,N_18644);
or U20608 (N_20608,N_18344,N_18828);
nor U20609 (N_20609,N_18231,N_19117);
xor U20610 (N_20610,N_18886,N_19716);
and U20611 (N_20611,N_18718,N_18308);
xor U20612 (N_20612,N_18928,N_18411);
nand U20613 (N_20613,N_19002,N_19381);
or U20614 (N_20614,N_18445,N_18586);
nand U20615 (N_20615,N_18457,N_18257);
nand U20616 (N_20616,N_18480,N_19427);
xor U20617 (N_20617,N_19518,N_18555);
and U20618 (N_20618,N_18060,N_19539);
nor U20619 (N_20619,N_19420,N_18501);
nand U20620 (N_20620,N_18845,N_18602);
and U20621 (N_20621,N_18151,N_19718);
nor U20622 (N_20622,N_18377,N_19635);
nand U20623 (N_20623,N_19089,N_19208);
nor U20624 (N_20624,N_19782,N_19774);
or U20625 (N_20625,N_18759,N_19375);
nor U20626 (N_20626,N_19875,N_19884);
and U20627 (N_20627,N_18375,N_18588);
and U20628 (N_20628,N_19771,N_18160);
and U20629 (N_20629,N_18307,N_19988);
xnor U20630 (N_20630,N_18543,N_18158);
xor U20631 (N_20631,N_19368,N_19608);
or U20632 (N_20632,N_18671,N_19442);
or U20633 (N_20633,N_19025,N_19962);
nor U20634 (N_20634,N_19665,N_18582);
nand U20635 (N_20635,N_19783,N_18464);
nand U20636 (N_20636,N_18568,N_19957);
nand U20637 (N_20637,N_19069,N_18115);
or U20638 (N_20638,N_19408,N_18156);
nand U20639 (N_20639,N_18522,N_19288);
xor U20640 (N_20640,N_18438,N_19732);
xor U20641 (N_20641,N_18756,N_19671);
or U20642 (N_20642,N_18896,N_18869);
and U20643 (N_20643,N_18604,N_18974);
or U20644 (N_20644,N_19876,N_19171);
nand U20645 (N_20645,N_19062,N_18351);
xnor U20646 (N_20646,N_18267,N_18636);
nor U20647 (N_20647,N_19512,N_19194);
or U20648 (N_20648,N_19414,N_19275);
xor U20649 (N_20649,N_18283,N_19406);
nand U20650 (N_20650,N_18992,N_19243);
and U20651 (N_20651,N_18425,N_18421);
nor U20652 (N_20652,N_19279,N_19666);
and U20653 (N_20653,N_19149,N_19821);
and U20654 (N_20654,N_18570,N_18851);
or U20655 (N_20655,N_19470,N_19650);
or U20656 (N_20656,N_18492,N_18259);
or U20657 (N_20657,N_18083,N_19457);
and U20658 (N_20658,N_18537,N_18658);
nand U20659 (N_20659,N_19823,N_19144);
nor U20660 (N_20660,N_19648,N_18352);
or U20661 (N_20661,N_18871,N_19354);
xor U20662 (N_20662,N_19215,N_19415);
or U20663 (N_20663,N_18300,N_19993);
nor U20664 (N_20664,N_18750,N_18835);
nand U20665 (N_20665,N_18415,N_18227);
and U20666 (N_20666,N_19858,N_19900);
nand U20667 (N_20667,N_19843,N_18017);
xor U20668 (N_20668,N_19430,N_19222);
nand U20669 (N_20669,N_18019,N_18916);
and U20670 (N_20670,N_19110,N_18630);
nor U20671 (N_20671,N_19225,N_19941);
and U20672 (N_20672,N_18712,N_19863);
and U20673 (N_20673,N_18482,N_18413);
nand U20674 (N_20674,N_19228,N_18985);
nor U20675 (N_20675,N_18813,N_18200);
and U20676 (N_20676,N_18979,N_18065);
or U20677 (N_20677,N_19309,N_18730);
xnor U20678 (N_20678,N_18370,N_18192);
xnor U20679 (N_20679,N_19044,N_18495);
nand U20680 (N_20680,N_19803,N_19615);
and U20681 (N_20681,N_19000,N_18194);
xor U20682 (N_20682,N_18326,N_18371);
nor U20683 (N_20683,N_18152,N_19206);
nor U20684 (N_20684,N_19474,N_19812);
nand U20685 (N_20685,N_19501,N_18819);
nor U20686 (N_20686,N_19237,N_18514);
and U20687 (N_20687,N_18209,N_19122);
and U20688 (N_20688,N_18583,N_19922);
nor U20689 (N_20689,N_19291,N_18823);
and U20690 (N_20690,N_18129,N_19913);
nor U20691 (N_20691,N_18672,N_18470);
xor U20692 (N_20692,N_18360,N_18673);
nor U20693 (N_20693,N_19794,N_19024);
nor U20694 (N_20694,N_18010,N_19250);
nor U20695 (N_20695,N_18557,N_19335);
nand U20696 (N_20696,N_19249,N_19646);
xnor U20697 (N_20697,N_19903,N_19102);
nand U20698 (N_20698,N_18287,N_18141);
xnor U20699 (N_20699,N_19032,N_18405);
xnor U20700 (N_20700,N_18576,N_19499);
xor U20701 (N_20701,N_19114,N_18806);
nor U20702 (N_20702,N_19399,N_19833);
nand U20703 (N_20703,N_18178,N_18688);
nor U20704 (N_20704,N_19475,N_19935);
and U20705 (N_20705,N_19535,N_18632);
xnor U20706 (N_20706,N_18006,N_19715);
and U20707 (N_20707,N_18059,N_19262);
xnor U20708 (N_20708,N_19493,N_19699);
nor U20709 (N_20709,N_19504,N_18804);
nor U20710 (N_20710,N_19525,N_19090);
nand U20711 (N_20711,N_18601,N_18383);
xor U20712 (N_20712,N_18548,N_18998);
nor U20713 (N_20713,N_19897,N_19128);
nor U20714 (N_20714,N_19028,N_18072);
and U20715 (N_20715,N_18318,N_18716);
nor U20716 (N_20716,N_18977,N_19257);
or U20717 (N_20717,N_18165,N_19346);
or U20718 (N_20718,N_19201,N_18198);
and U20719 (N_20719,N_18633,N_19734);
or U20720 (N_20720,N_18110,N_18391);
xor U20721 (N_20721,N_19642,N_18416);
nand U20722 (N_20722,N_18993,N_19586);
or U20723 (N_20723,N_19856,N_19686);
and U20724 (N_20724,N_18609,N_19261);
nand U20725 (N_20725,N_19536,N_18840);
or U20726 (N_20726,N_19376,N_19324);
xnor U20727 (N_20727,N_18507,N_19700);
nand U20728 (N_20728,N_19872,N_18862);
nand U20729 (N_20729,N_19799,N_19418);
xor U20730 (N_20730,N_18030,N_18995);
nand U20731 (N_20731,N_18794,N_18774);
nand U20732 (N_20732,N_19465,N_18968);
nand U20733 (N_20733,N_19521,N_19226);
nand U20734 (N_20734,N_18497,N_19310);
xor U20735 (N_20735,N_18542,N_19769);
nand U20736 (N_20736,N_18182,N_18314);
nor U20737 (N_20737,N_18580,N_19571);
nor U20738 (N_20738,N_18237,N_19255);
and U20739 (N_20739,N_18297,N_18707);
nor U20740 (N_20740,N_18489,N_19549);
or U20741 (N_20741,N_18163,N_19500);
and U20742 (N_20742,N_19041,N_18970);
xor U20743 (N_20743,N_19819,N_19709);
and U20744 (N_20744,N_19198,N_18325);
xnor U20745 (N_20745,N_19660,N_19914);
or U20746 (N_20746,N_18861,N_19073);
or U20747 (N_20747,N_18272,N_19523);
nand U20748 (N_20748,N_19685,N_19286);
or U20749 (N_20749,N_18841,N_19560);
nor U20750 (N_20750,N_19810,N_18597);
or U20751 (N_20751,N_19239,N_19386);
and U20752 (N_20752,N_19619,N_19983);
or U20753 (N_20753,N_18226,N_18714);
xor U20754 (N_20754,N_19707,N_19064);
or U20755 (N_20755,N_18713,N_19070);
and U20756 (N_20756,N_19344,N_19135);
nand U20757 (N_20757,N_19101,N_18364);
xor U20758 (N_20758,N_19355,N_18829);
nor U20759 (N_20759,N_18131,N_18544);
or U20760 (N_20760,N_19285,N_18938);
or U20761 (N_20761,N_18550,N_19704);
or U20762 (N_20762,N_18717,N_19299);
or U20763 (N_20763,N_18710,N_19678);
or U20764 (N_20764,N_18335,N_18498);
or U20765 (N_20765,N_19773,N_19713);
nand U20766 (N_20766,N_19624,N_18485);
or U20767 (N_20767,N_18735,N_18691);
or U20768 (N_20768,N_19081,N_18243);
and U20769 (N_20769,N_19204,N_18263);
xor U20770 (N_20770,N_19995,N_18843);
or U20771 (N_20771,N_18908,N_19012);
or U20772 (N_20772,N_19173,N_18403);
and U20773 (N_20773,N_18466,N_18873);
xnor U20774 (N_20774,N_19817,N_19684);
xor U20775 (N_20775,N_18372,N_18704);
and U20776 (N_20776,N_18986,N_19514);
nand U20777 (N_20777,N_19147,N_19221);
and U20778 (N_20778,N_18069,N_18893);
and U20779 (N_20779,N_19111,N_19600);
and U20780 (N_20780,N_19138,N_18232);
or U20781 (N_20781,N_19930,N_19447);
xnor U20782 (N_20782,N_19071,N_19193);
or U20783 (N_20783,N_18740,N_19172);
nor U20784 (N_20784,N_18222,N_18103);
xor U20785 (N_20785,N_19987,N_18459);
nor U20786 (N_20786,N_18779,N_19317);
and U20787 (N_20787,N_18387,N_18206);
nor U20788 (N_20788,N_19021,N_18505);
or U20789 (N_20789,N_18274,N_18255);
and U20790 (N_20790,N_19314,N_19078);
or U20791 (N_20791,N_19409,N_18140);
nand U20792 (N_20792,N_19506,N_19548);
or U20793 (N_20793,N_19029,N_18931);
nand U20794 (N_20794,N_18502,N_18874);
nor U20795 (N_20795,N_18592,N_18685);
xnor U20796 (N_20796,N_19909,N_18915);
xor U20797 (N_20797,N_18348,N_19510);
nor U20798 (N_20798,N_18419,N_18729);
nand U20799 (N_20799,N_18412,N_18776);
nor U20800 (N_20800,N_18642,N_19503);
nand U20801 (N_20801,N_19464,N_19370);
nand U20802 (N_20802,N_18956,N_18093);
nor U20803 (N_20803,N_19217,N_19140);
and U20804 (N_20804,N_19277,N_19928);
and U20805 (N_20805,N_18468,N_18180);
nand U20806 (N_20806,N_19378,N_19449);
and U20807 (N_20807,N_19224,N_18558);
or U20808 (N_20808,N_18277,N_19063);
nand U20809 (N_20809,N_18266,N_18296);
nor U20810 (N_20810,N_19550,N_19835);
or U20811 (N_20811,N_19661,N_19433);
nand U20812 (N_20812,N_19893,N_19293);
xor U20813 (N_20813,N_19177,N_18109);
nor U20814 (N_20814,N_18145,N_19419);
nand U20815 (N_20815,N_18313,N_18172);
nor U20816 (N_20816,N_19807,N_19421);
and U20817 (N_20817,N_18546,N_18961);
nand U20818 (N_20818,N_19565,N_19952);
nor U20819 (N_20819,N_19371,N_19862);
and U20820 (N_20820,N_18056,N_18431);
xnor U20821 (N_20821,N_18074,N_18467);
nand U20822 (N_20822,N_19236,N_19462);
nand U20823 (N_20823,N_18741,N_19043);
nand U20824 (N_20824,N_18589,N_19868);
nor U20825 (N_20825,N_19751,N_18875);
nand U20826 (N_20826,N_19694,N_19977);
and U20827 (N_20827,N_18881,N_18363);
and U20828 (N_20828,N_18157,N_19526);
nand U20829 (N_20829,N_18164,N_19341);
xnor U20830 (N_20830,N_19622,N_18639);
or U20831 (N_20831,N_18773,N_18225);
nand U20832 (N_20832,N_19207,N_19167);
and U20833 (N_20833,N_18653,N_19796);
and U20834 (N_20834,N_19467,N_19762);
xnor U20835 (N_20835,N_18594,N_18565);
and U20836 (N_20836,N_18769,N_18556);
nand U20837 (N_20837,N_19284,N_19425);
nand U20838 (N_20838,N_18595,N_18203);
nand U20839 (N_20839,N_19254,N_18469);
nand U20840 (N_20840,N_18984,N_18834);
xor U20841 (N_20841,N_18380,N_18290);
nand U20842 (N_20842,N_19342,N_18781);
or U20843 (N_20843,N_18768,N_19680);
and U20844 (N_20844,N_19150,N_18035);
xor U20845 (N_20845,N_19989,N_19838);
xnor U20846 (N_20846,N_19080,N_19428);
nor U20847 (N_20847,N_19027,N_19258);
and U20848 (N_20848,N_19811,N_18261);
nor U20849 (N_20849,N_19861,N_18493);
nor U20850 (N_20850,N_18600,N_18913);
or U20851 (N_20851,N_19247,N_18417);
xor U20852 (N_20852,N_18304,N_18980);
and U20853 (N_20853,N_19181,N_18912);
xnor U20854 (N_20854,N_19792,N_19058);
and U20855 (N_20855,N_18569,N_18213);
and U20856 (N_20856,N_18574,N_18037);
nand U20857 (N_20857,N_18212,N_18761);
xor U20858 (N_20858,N_18675,N_19413);
nand U20859 (N_20859,N_18328,N_18251);
and U20860 (N_20860,N_19052,N_19302);
or U20861 (N_20861,N_18051,N_18855);
nand U20862 (N_20862,N_18215,N_19589);
nor U20863 (N_20863,N_18282,N_19673);
xnor U20864 (N_20864,N_18043,N_18343);
nor U20865 (N_20865,N_19471,N_18965);
or U20866 (N_20866,N_18800,N_18310);
and U20867 (N_20867,N_18341,N_18291);
nand U20868 (N_20868,N_18990,N_19083);
nor U20869 (N_20869,N_19010,N_18045);
nor U20870 (N_20870,N_18842,N_19164);
nand U20871 (N_20871,N_18585,N_19502);
xor U20872 (N_20872,N_19210,N_18086);
nand U20873 (N_20873,N_19853,N_18863);
xnor U20874 (N_20874,N_18892,N_18439);
or U20875 (N_20875,N_19898,N_19116);
and U20876 (N_20876,N_18062,N_19353);
xnor U20877 (N_20877,N_19689,N_19059);
or U20878 (N_20878,N_19227,N_19345);
or U20879 (N_20879,N_19592,N_18599);
and U20880 (N_20880,N_18976,N_19587);
nand U20881 (N_20881,N_18883,N_19098);
xor U20882 (N_20882,N_18725,N_18651);
and U20883 (N_20883,N_18560,N_19084);
nand U20884 (N_20884,N_18476,N_18236);
or U20885 (N_20885,N_18926,N_19014);
nand U20886 (N_20886,N_19808,N_19612);
xnor U20887 (N_20887,N_18923,N_19737);
or U20888 (N_20888,N_18070,N_18638);
nor U20889 (N_20889,N_18376,N_18332);
or U20890 (N_20890,N_18329,N_18625);
and U20891 (N_20891,N_18878,N_18999);
xnor U20892 (N_20892,N_18094,N_18000);
xor U20893 (N_20893,N_18811,N_18081);
and U20894 (N_20894,N_19460,N_19978);
or U20895 (N_20895,N_18064,N_19366);
or U20896 (N_20896,N_19784,N_18924);
xor U20897 (N_20897,N_18452,N_19878);
xor U20898 (N_20898,N_18173,N_18518);
or U20899 (N_20899,N_18484,N_19497);
xor U20900 (N_20900,N_18782,N_18532);
or U20901 (N_20901,N_18473,N_19306);
xor U20902 (N_20902,N_19238,N_18312);
and U20903 (N_20903,N_18356,N_18536);
xnor U20904 (N_20904,N_18012,N_19750);
xor U20905 (N_20905,N_18410,N_18032);
nor U20906 (N_20906,N_18605,N_19652);
nand U20907 (N_20907,N_18235,N_19874);
nand U20908 (N_20908,N_18950,N_19626);
or U20909 (N_20909,N_19690,N_19017);
xor U20910 (N_20910,N_18336,N_19290);
nand U20911 (N_20911,N_19137,N_18108);
and U20912 (N_20912,N_19653,N_19165);
xnor U20913 (N_20913,N_18785,N_19801);
and U20914 (N_20914,N_19018,N_18775);
nor U20915 (N_20915,N_18448,N_18927);
or U20916 (N_20916,N_19985,N_18879);
xnor U20917 (N_20917,N_19097,N_18451);
and U20918 (N_20918,N_19790,N_18395);
nor U20919 (N_20919,N_19848,N_18983);
nor U20920 (N_20920,N_18374,N_18637);
or U20921 (N_20921,N_19259,N_19904);
and U20922 (N_20922,N_18613,N_19659);
xnor U20923 (N_20923,N_19818,N_18478);
nor U20924 (N_20924,N_18866,N_19185);
xor U20925 (N_20925,N_19991,N_19033);
xor U20926 (N_20926,N_19564,N_18853);
or U20927 (N_20927,N_18662,N_19452);
nand U20928 (N_20928,N_18442,N_18723);
xor U20929 (N_20929,N_19931,N_19075);
nand U20930 (N_20930,N_18509,N_18104);
xor U20931 (N_20931,N_19218,N_19596);
and U20932 (N_20932,N_19479,N_18076);
nor U20933 (N_20933,N_19282,N_18969);
and U20934 (N_20934,N_19496,N_18271);
nor U20935 (N_20935,N_19702,N_19778);
or U20936 (N_20936,N_19948,N_19085);
nor U20937 (N_20937,N_19205,N_19873);
nand U20938 (N_20938,N_19082,N_19940);
and U20939 (N_20939,N_19871,N_18154);
and U20940 (N_20940,N_18791,N_18322);
and U20941 (N_20941,N_18433,N_18815);
xor U20942 (N_20942,N_19398,N_18684);
nor U20943 (N_20943,N_19556,N_19656);
and U20944 (N_20944,N_18699,N_19141);
or U20945 (N_20945,N_19325,N_19358);
xnor U20946 (N_20946,N_19579,N_19480);
xor U20947 (N_20947,N_19687,N_18101);
xor U20948 (N_20948,N_18214,N_18553);
nand U20949 (N_20949,N_18133,N_19031);
and U20950 (N_20950,N_19292,N_18463);
and U20951 (N_20951,N_19362,N_18330);
nand U20952 (N_20952,N_18366,N_19620);
nor U20953 (N_20953,N_19969,N_19196);
xor U20954 (N_20954,N_19006,N_18179);
or U20955 (N_20955,N_19308,N_19268);
nor U20956 (N_20956,N_18455,N_19742);
xnor U20957 (N_20957,N_19809,N_18240);
or U20958 (N_20958,N_19203,N_18643);
xor U20959 (N_20959,N_18884,N_19124);
nand U20960 (N_20960,N_19404,N_18401);
and U20961 (N_20961,N_19845,N_18018);
or U20962 (N_20962,N_19851,N_19343);
nor U20963 (N_20963,N_19486,N_18856);
xor U20964 (N_20964,N_19920,N_18316);
nand U20965 (N_20965,N_19944,N_19585);
xnor U20966 (N_20966,N_19649,N_19691);
and U20967 (N_20967,N_19391,N_19637);
nand U20968 (N_20968,N_18248,N_18797);
nor U20969 (N_20969,N_18004,N_19410);
xnor U20970 (N_20970,N_19446,N_18265);
xnor U20971 (N_20971,N_18748,N_19740);
or U20972 (N_20972,N_18306,N_19915);
xor U20973 (N_20973,N_18221,N_19959);
and U20974 (N_20974,N_19232,N_18816);
xor U20975 (N_20975,N_18762,N_19517);
and U20976 (N_20976,N_18386,N_18789);
xnor U20977 (N_20977,N_19359,N_19013);
nand U20978 (N_20978,N_19695,N_18122);
xnor U20979 (N_20979,N_18239,N_19190);
xor U20980 (N_20980,N_19857,N_19825);
nor U20981 (N_20981,N_18022,N_18436);
nand U20982 (N_20982,N_18777,N_19214);
nor U20983 (N_20983,N_18659,N_18528);
and U20984 (N_20984,N_18205,N_19365);
nor U20985 (N_20985,N_18989,N_19392);
or U20986 (N_20986,N_19484,N_18838);
xnor U20987 (N_20987,N_19538,N_19192);
nand U20988 (N_20988,N_18906,N_19180);
and U20989 (N_20989,N_19555,N_19627);
nand U20990 (N_20990,N_18654,N_18107);
nor U20991 (N_20991,N_19647,N_19489);
or U20992 (N_20992,N_18890,N_19772);
and U20993 (N_20993,N_18091,N_19994);
xor U20994 (N_20994,N_18367,N_18116);
nand U20995 (N_20995,N_19891,N_18219);
and U20996 (N_20996,N_19529,N_18836);
xor U20997 (N_20997,N_19372,N_18807);
or U20998 (N_20998,N_18288,N_19572);
nor U20999 (N_20999,N_19890,N_19356);
or U21000 (N_21000,N_19105,N_18750);
and U21001 (N_21001,N_19764,N_19850);
nor U21002 (N_21002,N_19721,N_18515);
and U21003 (N_21003,N_19116,N_19846);
xnor U21004 (N_21004,N_19024,N_19202);
nand U21005 (N_21005,N_19559,N_19229);
xnor U21006 (N_21006,N_19117,N_18848);
and U21007 (N_21007,N_18262,N_19304);
xnor U21008 (N_21008,N_19359,N_19349);
and U21009 (N_21009,N_19584,N_19799);
and U21010 (N_21010,N_18983,N_18773);
xor U21011 (N_21011,N_18317,N_18322);
or U21012 (N_21012,N_18980,N_19213);
and U21013 (N_21013,N_18896,N_19052);
nand U21014 (N_21014,N_19119,N_19454);
nand U21015 (N_21015,N_19581,N_18205);
nor U21016 (N_21016,N_19038,N_18984);
and U21017 (N_21017,N_18417,N_19947);
nor U21018 (N_21018,N_18129,N_19382);
nand U21019 (N_21019,N_18245,N_18976);
or U21020 (N_21020,N_19302,N_19490);
nand U21021 (N_21021,N_18939,N_19976);
or U21022 (N_21022,N_19420,N_18692);
or U21023 (N_21023,N_18162,N_18132);
nor U21024 (N_21024,N_18497,N_18294);
nand U21025 (N_21025,N_18384,N_19912);
or U21026 (N_21026,N_19662,N_18747);
nand U21027 (N_21027,N_18081,N_18480);
or U21028 (N_21028,N_18644,N_18358);
and U21029 (N_21029,N_19649,N_19861);
nand U21030 (N_21030,N_18144,N_19224);
or U21031 (N_21031,N_19336,N_18537);
nor U21032 (N_21032,N_19899,N_18094);
nand U21033 (N_21033,N_18812,N_19472);
or U21034 (N_21034,N_18763,N_18075);
xor U21035 (N_21035,N_18286,N_19986);
nand U21036 (N_21036,N_19105,N_19438);
nand U21037 (N_21037,N_19590,N_18174);
xor U21038 (N_21038,N_19482,N_19117);
and U21039 (N_21039,N_18200,N_18249);
nand U21040 (N_21040,N_19539,N_19197);
and U21041 (N_21041,N_19970,N_19181);
or U21042 (N_21042,N_18341,N_19786);
xnor U21043 (N_21043,N_18468,N_18336);
and U21044 (N_21044,N_19029,N_19874);
nor U21045 (N_21045,N_19152,N_18111);
or U21046 (N_21046,N_18530,N_19955);
nor U21047 (N_21047,N_18484,N_19445);
nand U21048 (N_21048,N_19613,N_19440);
nand U21049 (N_21049,N_19631,N_18445);
xor U21050 (N_21050,N_19415,N_18689);
or U21051 (N_21051,N_18559,N_18280);
xnor U21052 (N_21052,N_19040,N_19306);
nand U21053 (N_21053,N_19762,N_18693);
nor U21054 (N_21054,N_18498,N_19137);
and U21055 (N_21055,N_19751,N_18867);
nor U21056 (N_21056,N_18972,N_18343);
nand U21057 (N_21057,N_19171,N_18671);
nand U21058 (N_21058,N_19607,N_18918);
nor U21059 (N_21059,N_18592,N_19700);
nor U21060 (N_21060,N_18384,N_18447);
and U21061 (N_21061,N_18857,N_19281);
nand U21062 (N_21062,N_18880,N_19077);
and U21063 (N_21063,N_19737,N_18339);
nand U21064 (N_21064,N_19510,N_19967);
or U21065 (N_21065,N_19628,N_19195);
or U21066 (N_21066,N_18312,N_18865);
nor U21067 (N_21067,N_18415,N_19186);
nor U21068 (N_21068,N_18703,N_18041);
or U21069 (N_21069,N_18339,N_18830);
and U21070 (N_21070,N_19005,N_19576);
or U21071 (N_21071,N_19963,N_18329);
nand U21072 (N_21072,N_19364,N_18325);
or U21073 (N_21073,N_18418,N_18457);
nor U21074 (N_21074,N_19760,N_19958);
nor U21075 (N_21075,N_18986,N_19991);
nor U21076 (N_21076,N_19964,N_19858);
xor U21077 (N_21077,N_19805,N_18721);
or U21078 (N_21078,N_18471,N_18598);
nand U21079 (N_21079,N_18226,N_18937);
xor U21080 (N_21080,N_18384,N_18535);
and U21081 (N_21081,N_18958,N_19827);
nor U21082 (N_21082,N_19125,N_19653);
nor U21083 (N_21083,N_19776,N_18180);
nand U21084 (N_21084,N_18470,N_18372);
or U21085 (N_21085,N_18018,N_19703);
xor U21086 (N_21086,N_19166,N_18278);
nor U21087 (N_21087,N_19197,N_19731);
and U21088 (N_21088,N_18085,N_18592);
nor U21089 (N_21089,N_19389,N_18556);
and U21090 (N_21090,N_19943,N_19895);
xor U21091 (N_21091,N_19973,N_18827);
xor U21092 (N_21092,N_18646,N_18366);
and U21093 (N_21093,N_18814,N_18395);
and U21094 (N_21094,N_18420,N_18504);
or U21095 (N_21095,N_18240,N_19269);
nand U21096 (N_21096,N_19010,N_19508);
and U21097 (N_21097,N_18686,N_18544);
nor U21098 (N_21098,N_19399,N_18546);
xnor U21099 (N_21099,N_19726,N_18535);
nand U21100 (N_21100,N_18065,N_19413);
or U21101 (N_21101,N_19616,N_19712);
and U21102 (N_21102,N_19818,N_19481);
xor U21103 (N_21103,N_19804,N_19022);
and U21104 (N_21104,N_19305,N_18057);
xnor U21105 (N_21105,N_18541,N_19763);
nand U21106 (N_21106,N_19728,N_19757);
or U21107 (N_21107,N_19310,N_18780);
nand U21108 (N_21108,N_19217,N_18871);
nand U21109 (N_21109,N_19952,N_18524);
xnor U21110 (N_21110,N_18494,N_18715);
or U21111 (N_21111,N_18228,N_19937);
nand U21112 (N_21112,N_19853,N_18115);
xor U21113 (N_21113,N_18277,N_18133);
or U21114 (N_21114,N_19299,N_18489);
nor U21115 (N_21115,N_18642,N_19550);
and U21116 (N_21116,N_19269,N_19252);
nand U21117 (N_21117,N_19543,N_19016);
nand U21118 (N_21118,N_19804,N_18161);
nand U21119 (N_21119,N_19391,N_18643);
or U21120 (N_21120,N_19971,N_18401);
or U21121 (N_21121,N_19327,N_19390);
or U21122 (N_21122,N_18215,N_19907);
and U21123 (N_21123,N_19295,N_19894);
nand U21124 (N_21124,N_19164,N_18926);
and U21125 (N_21125,N_19300,N_19314);
and U21126 (N_21126,N_18230,N_19171);
nand U21127 (N_21127,N_19593,N_19097);
or U21128 (N_21128,N_18675,N_18391);
xnor U21129 (N_21129,N_18384,N_19266);
xor U21130 (N_21130,N_19895,N_19823);
nand U21131 (N_21131,N_19898,N_19482);
xnor U21132 (N_21132,N_18566,N_18813);
nand U21133 (N_21133,N_18245,N_18294);
xor U21134 (N_21134,N_18137,N_18279);
nand U21135 (N_21135,N_18334,N_18694);
or U21136 (N_21136,N_19646,N_19123);
nand U21137 (N_21137,N_18087,N_18529);
xor U21138 (N_21138,N_18014,N_19088);
nand U21139 (N_21139,N_18224,N_19926);
xnor U21140 (N_21140,N_18310,N_18724);
nand U21141 (N_21141,N_18843,N_19760);
and U21142 (N_21142,N_18918,N_19933);
nor U21143 (N_21143,N_18932,N_18993);
and U21144 (N_21144,N_19791,N_19701);
xor U21145 (N_21145,N_19825,N_19885);
nand U21146 (N_21146,N_19380,N_18624);
nor U21147 (N_21147,N_19441,N_18595);
nor U21148 (N_21148,N_19547,N_19513);
nand U21149 (N_21149,N_18168,N_18839);
nand U21150 (N_21150,N_19088,N_19447);
xor U21151 (N_21151,N_18925,N_18786);
nor U21152 (N_21152,N_18051,N_19275);
nor U21153 (N_21153,N_19156,N_18358);
or U21154 (N_21154,N_18982,N_19430);
nand U21155 (N_21155,N_18296,N_18896);
and U21156 (N_21156,N_19632,N_19706);
xor U21157 (N_21157,N_18469,N_18197);
or U21158 (N_21158,N_19455,N_18075);
or U21159 (N_21159,N_18814,N_18492);
and U21160 (N_21160,N_18004,N_18834);
xor U21161 (N_21161,N_19824,N_18491);
and U21162 (N_21162,N_18530,N_18905);
or U21163 (N_21163,N_19891,N_19328);
xnor U21164 (N_21164,N_19417,N_18645);
or U21165 (N_21165,N_19759,N_19099);
xor U21166 (N_21166,N_18843,N_18837);
and U21167 (N_21167,N_19960,N_18674);
and U21168 (N_21168,N_19720,N_19933);
xnor U21169 (N_21169,N_18714,N_19843);
xor U21170 (N_21170,N_19451,N_19763);
nor U21171 (N_21171,N_19322,N_18995);
or U21172 (N_21172,N_19613,N_18855);
nand U21173 (N_21173,N_18484,N_18622);
or U21174 (N_21174,N_18238,N_18018);
nand U21175 (N_21175,N_18829,N_19778);
xor U21176 (N_21176,N_19860,N_18911);
nor U21177 (N_21177,N_18839,N_18364);
nand U21178 (N_21178,N_18784,N_19844);
and U21179 (N_21179,N_19253,N_19438);
xnor U21180 (N_21180,N_18149,N_19243);
and U21181 (N_21181,N_18186,N_18801);
or U21182 (N_21182,N_18002,N_18186);
nand U21183 (N_21183,N_18518,N_18822);
nand U21184 (N_21184,N_18038,N_18518);
nor U21185 (N_21185,N_18251,N_19404);
or U21186 (N_21186,N_18490,N_18472);
or U21187 (N_21187,N_19533,N_18309);
nand U21188 (N_21188,N_18774,N_18886);
nand U21189 (N_21189,N_18666,N_19446);
or U21190 (N_21190,N_19882,N_18604);
nor U21191 (N_21191,N_18077,N_19986);
nand U21192 (N_21192,N_19868,N_18453);
or U21193 (N_21193,N_19317,N_18008);
xor U21194 (N_21194,N_18692,N_18844);
nand U21195 (N_21195,N_19482,N_18853);
and U21196 (N_21196,N_18713,N_18241);
nor U21197 (N_21197,N_19851,N_19122);
and U21198 (N_21198,N_19644,N_19448);
nor U21199 (N_21199,N_19826,N_18831);
and U21200 (N_21200,N_19890,N_18562);
nor U21201 (N_21201,N_19658,N_19831);
and U21202 (N_21202,N_18979,N_18765);
nand U21203 (N_21203,N_18606,N_18792);
or U21204 (N_21204,N_18228,N_19025);
and U21205 (N_21205,N_19481,N_19915);
and U21206 (N_21206,N_18732,N_19224);
xnor U21207 (N_21207,N_19905,N_19177);
xor U21208 (N_21208,N_18751,N_19097);
nor U21209 (N_21209,N_19923,N_18865);
nand U21210 (N_21210,N_19188,N_19954);
nand U21211 (N_21211,N_19673,N_19559);
xnor U21212 (N_21212,N_18536,N_19709);
or U21213 (N_21213,N_19666,N_19082);
nand U21214 (N_21214,N_18250,N_18117);
and U21215 (N_21215,N_19101,N_19811);
nand U21216 (N_21216,N_18336,N_19791);
xor U21217 (N_21217,N_18361,N_19853);
and U21218 (N_21218,N_19063,N_19753);
nand U21219 (N_21219,N_18567,N_18662);
nor U21220 (N_21220,N_19166,N_19940);
or U21221 (N_21221,N_18095,N_18837);
and U21222 (N_21222,N_18647,N_19149);
nand U21223 (N_21223,N_19955,N_18383);
nor U21224 (N_21224,N_18343,N_19224);
or U21225 (N_21225,N_18510,N_19461);
and U21226 (N_21226,N_19407,N_19371);
nand U21227 (N_21227,N_19720,N_18576);
nand U21228 (N_21228,N_18386,N_19743);
nor U21229 (N_21229,N_18788,N_19710);
nor U21230 (N_21230,N_19894,N_19599);
nand U21231 (N_21231,N_18730,N_18990);
or U21232 (N_21232,N_19757,N_18329);
xnor U21233 (N_21233,N_18160,N_19649);
or U21234 (N_21234,N_19947,N_19153);
and U21235 (N_21235,N_18028,N_19013);
or U21236 (N_21236,N_18169,N_19305);
nor U21237 (N_21237,N_19013,N_19901);
and U21238 (N_21238,N_19750,N_18591);
nor U21239 (N_21239,N_18685,N_19539);
nand U21240 (N_21240,N_18274,N_18433);
nand U21241 (N_21241,N_19147,N_19654);
and U21242 (N_21242,N_18152,N_19825);
or U21243 (N_21243,N_18342,N_18642);
nand U21244 (N_21244,N_19607,N_18699);
nor U21245 (N_21245,N_19000,N_19502);
nand U21246 (N_21246,N_19867,N_18867);
xnor U21247 (N_21247,N_19592,N_18370);
nand U21248 (N_21248,N_19132,N_18488);
or U21249 (N_21249,N_19721,N_19718);
and U21250 (N_21250,N_19266,N_18460);
or U21251 (N_21251,N_19528,N_19159);
nor U21252 (N_21252,N_18802,N_19702);
nand U21253 (N_21253,N_19269,N_19300);
and U21254 (N_21254,N_19615,N_19244);
or U21255 (N_21255,N_18595,N_19347);
or U21256 (N_21256,N_18252,N_18587);
nand U21257 (N_21257,N_19692,N_18420);
and U21258 (N_21258,N_18973,N_19842);
or U21259 (N_21259,N_19127,N_18639);
nor U21260 (N_21260,N_19868,N_18283);
nand U21261 (N_21261,N_18585,N_18904);
or U21262 (N_21262,N_19588,N_18068);
xnor U21263 (N_21263,N_19582,N_18587);
and U21264 (N_21264,N_19675,N_19749);
nor U21265 (N_21265,N_18878,N_18645);
or U21266 (N_21266,N_19724,N_18981);
and U21267 (N_21267,N_18555,N_19288);
and U21268 (N_21268,N_18531,N_19907);
or U21269 (N_21269,N_19805,N_19553);
nand U21270 (N_21270,N_19970,N_18558);
or U21271 (N_21271,N_19389,N_19219);
nor U21272 (N_21272,N_19201,N_19519);
xor U21273 (N_21273,N_19084,N_19029);
nor U21274 (N_21274,N_18492,N_18769);
or U21275 (N_21275,N_18237,N_19385);
nor U21276 (N_21276,N_19510,N_18622);
or U21277 (N_21277,N_18398,N_19199);
xnor U21278 (N_21278,N_19346,N_19870);
or U21279 (N_21279,N_18210,N_19605);
nor U21280 (N_21280,N_19446,N_18512);
nand U21281 (N_21281,N_19860,N_18628);
nand U21282 (N_21282,N_19447,N_18770);
and U21283 (N_21283,N_19800,N_19717);
xnor U21284 (N_21284,N_19915,N_19719);
nor U21285 (N_21285,N_18852,N_19403);
and U21286 (N_21286,N_19380,N_18522);
nor U21287 (N_21287,N_19956,N_18498);
xnor U21288 (N_21288,N_18984,N_18381);
nand U21289 (N_21289,N_19437,N_18817);
nor U21290 (N_21290,N_18557,N_19481);
nand U21291 (N_21291,N_19408,N_19050);
nand U21292 (N_21292,N_18747,N_18522);
or U21293 (N_21293,N_19413,N_18821);
and U21294 (N_21294,N_18698,N_19771);
nand U21295 (N_21295,N_19369,N_19030);
nor U21296 (N_21296,N_19717,N_19477);
nor U21297 (N_21297,N_18917,N_18715);
xor U21298 (N_21298,N_19887,N_18695);
and U21299 (N_21299,N_19721,N_19380);
xor U21300 (N_21300,N_19158,N_19847);
xnor U21301 (N_21301,N_19016,N_18313);
or U21302 (N_21302,N_19457,N_19304);
and U21303 (N_21303,N_18964,N_19371);
nand U21304 (N_21304,N_19462,N_18489);
and U21305 (N_21305,N_18868,N_19935);
nor U21306 (N_21306,N_19938,N_18320);
and U21307 (N_21307,N_19006,N_18260);
xor U21308 (N_21308,N_19486,N_19019);
or U21309 (N_21309,N_18242,N_18937);
nor U21310 (N_21310,N_18530,N_19811);
or U21311 (N_21311,N_19210,N_19379);
nand U21312 (N_21312,N_18261,N_18596);
xnor U21313 (N_21313,N_18527,N_18058);
and U21314 (N_21314,N_18617,N_19759);
xnor U21315 (N_21315,N_19042,N_18498);
nor U21316 (N_21316,N_18334,N_18841);
nand U21317 (N_21317,N_19722,N_18495);
xnor U21318 (N_21318,N_19975,N_18934);
or U21319 (N_21319,N_18609,N_18465);
or U21320 (N_21320,N_19854,N_18098);
nand U21321 (N_21321,N_18948,N_19324);
or U21322 (N_21322,N_19230,N_19227);
nand U21323 (N_21323,N_19677,N_18564);
nor U21324 (N_21324,N_19733,N_19101);
nand U21325 (N_21325,N_19753,N_19606);
nor U21326 (N_21326,N_18113,N_19780);
nand U21327 (N_21327,N_19707,N_19692);
nand U21328 (N_21328,N_19943,N_19070);
nor U21329 (N_21329,N_18486,N_19191);
nor U21330 (N_21330,N_19615,N_19906);
nand U21331 (N_21331,N_18255,N_19704);
xor U21332 (N_21332,N_19586,N_19929);
or U21333 (N_21333,N_19043,N_18115);
xnor U21334 (N_21334,N_19689,N_19543);
and U21335 (N_21335,N_18366,N_19595);
or U21336 (N_21336,N_19145,N_19122);
nand U21337 (N_21337,N_19630,N_19956);
or U21338 (N_21338,N_19610,N_18776);
nor U21339 (N_21339,N_18421,N_18492);
nand U21340 (N_21340,N_18780,N_18963);
nand U21341 (N_21341,N_18659,N_19106);
nand U21342 (N_21342,N_18627,N_19955);
and U21343 (N_21343,N_19402,N_18514);
xnor U21344 (N_21344,N_18700,N_18167);
and U21345 (N_21345,N_18655,N_19367);
or U21346 (N_21346,N_18901,N_18274);
xnor U21347 (N_21347,N_18840,N_19291);
xor U21348 (N_21348,N_19900,N_18916);
nand U21349 (N_21349,N_18836,N_18209);
and U21350 (N_21350,N_19643,N_18842);
nor U21351 (N_21351,N_19217,N_18542);
xnor U21352 (N_21352,N_19541,N_18258);
nand U21353 (N_21353,N_18652,N_18566);
nand U21354 (N_21354,N_19246,N_18328);
or U21355 (N_21355,N_19163,N_19067);
nand U21356 (N_21356,N_18241,N_18971);
xnor U21357 (N_21357,N_19880,N_19726);
nand U21358 (N_21358,N_18209,N_18994);
nor U21359 (N_21359,N_19831,N_18439);
and U21360 (N_21360,N_18893,N_18349);
nand U21361 (N_21361,N_18874,N_18988);
xnor U21362 (N_21362,N_19001,N_19598);
nor U21363 (N_21363,N_18696,N_19587);
nor U21364 (N_21364,N_19573,N_18281);
nand U21365 (N_21365,N_18388,N_19830);
nor U21366 (N_21366,N_19056,N_18556);
nor U21367 (N_21367,N_18133,N_18927);
nand U21368 (N_21368,N_18708,N_18646);
nor U21369 (N_21369,N_19883,N_19172);
and U21370 (N_21370,N_19290,N_18923);
nor U21371 (N_21371,N_18489,N_18968);
nand U21372 (N_21372,N_18165,N_19569);
and U21373 (N_21373,N_19325,N_18810);
nand U21374 (N_21374,N_19881,N_19820);
and U21375 (N_21375,N_18988,N_19197);
and U21376 (N_21376,N_19716,N_19268);
nor U21377 (N_21377,N_18583,N_19871);
nor U21378 (N_21378,N_18524,N_19293);
xor U21379 (N_21379,N_18572,N_18194);
or U21380 (N_21380,N_18106,N_19651);
xor U21381 (N_21381,N_18233,N_18269);
nand U21382 (N_21382,N_19748,N_18783);
and U21383 (N_21383,N_19212,N_19788);
xor U21384 (N_21384,N_19770,N_18570);
nand U21385 (N_21385,N_18391,N_18180);
nand U21386 (N_21386,N_18089,N_18834);
nand U21387 (N_21387,N_18996,N_19735);
nand U21388 (N_21388,N_19222,N_19393);
nand U21389 (N_21389,N_19753,N_19378);
nand U21390 (N_21390,N_18223,N_19536);
nand U21391 (N_21391,N_19814,N_19038);
or U21392 (N_21392,N_19337,N_18758);
xor U21393 (N_21393,N_18696,N_18916);
or U21394 (N_21394,N_18053,N_18709);
and U21395 (N_21395,N_19778,N_18310);
nor U21396 (N_21396,N_19758,N_19427);
nor U21397 (N_21397,N_19469,N_19572);
and U21398 (N_21398,N_18372,N_18607);
nor U21399 (N_21399,N_19282,N_18039);
or U21400 (N_21400,N_18884,N_18367);
nor U21401 (N_21401,N_19116,N_18804);
nor U21402 (N_21402,N_19525,N_18565);
xor U21403 (N_21403,N_18508,N_18062);
nor U21404 (N_21404,N_18029,N_18986);
nor U21405 (N_21405,N_18238,N_19868);
nor U21406 (N_21406,N_18510,N_18731);
xnor U21407 (N_21407,N_18913,N_18689);
xnor U21408 (N_21408,N_19009,N_18372);
xnor U21409 (N_21409,N_19636,N_18365);
nor U21410 (N_21410,N_18443,N_18408);
and U21411 (N_21411,N_19065,N_19859);
and U21412 (N_21412,N_18311,N_19911);
or U21413 (N_21413,N_18041,N_18438);
nand U21414 (N_21414,N_19221,N_19783);
xor U21415 (N_21415,N_18171,N_18249);
nand U21416 (N_21416,N_18617,N_19528);
nor U21417 (N_21417,N_19004,N_19541);
and U21418 (N_21418,N_18846,N_18054);
nor U21419 (N_21419,N_19902,N_19033);
or U21420 (N_21420,N_19816,N_18046);
nor U21421 (N_21421,N_18733,N_19239);
nand U21422 (N_21422,N_18107,N_18358);
or U21423 (N_21423,N_18538,N_19252);
nand U21424 (N_21424,N_18718,N_19455);
nand U21425 (N_21425,N_18974,N_18128);
and U21426 (N_21426,N_18638,N_19729);
and U21427 (N_21427,N_19949,N_19017);
and U21428 (N_21428,N_18160,N_18476);
and U21429 (N_21429,N_19078,N_19045);
nor U21430 (N_21430,N_19696,N_18891);
or U21431 (N_21431,N_18996,N_19839);
xnor U21432 (N_21432,N_19004,N_19661);
nor U21433 (N_21433,N_18558,N_18642);
nand U21434 (N_21434,N_18125,N_19254);
nor U21435 (N_21435,N_19786,N_19655);
or U21436 (N_21436,N_18574,N_19367);
or U21437 (N_21437,N_18478,N_19134);
and U21438 (N_21438,N_19281,N_18297);
nand U21439 (N_21439,N_19715,N_19395);
nor U21440 (N_21440,N_18891,N_18978);
xor U21441 (N_21441,N_18869,N_19920);
xor U21442 (N_21442,N_18150,N_18576);
or U21443 (N_21443,N_18749,N_18802);
xor U21444 (N_21444,N_18666,N_19610);
xnor U21445 (N_21445,N_18246,N_19716);
and U21446 (N_21446,N_18634,N_19259);
nor U21447 (N_21447,N_18906,N_18693);
and U21448 (N_21448,N_18526,N_18181);
nand U21449 (N_21449,N_18220,N_19724);
nand U21450 (N_21450,N_19557,N_19879);
and U21451 (N_21451,N_18038,N_18665);
nand U21452 (N_21452,N_19253,N_18675);
or U21453 (N_21453,N_18838,N_18230);
xnor U21454 (N_21454,N_18676,N_19369);
xor U21455 (N_21455,N_19259,N_18159);
xnor U21456 (N_21456,N_18037,N_18987);
xor U21457 (N_21457,N_18854,N_18827);
nor U21458 (N_21458,N_19693,N_19700);
or U21459 (N_21459,N_18868,N_18143);
or U21460 (N_21460,N_19375,N_18662);
or U21461 (N_21461,N_18326,N_19972);
nand U21462 (N_21462,N_19386,N_19785);
or U21463 (N_21463,N_19841,N_19352);
nand U21464 (N_21464,N_18194,N_18361);
xor U21465 (N_21465,N_19510,N_18388);
nor U21466 (N_21466,N_19006,N_19102);
or U21467 (N_21467,N_19277,N_19282);
nand U21468 (N_21468,N_19468,N_19811);
or U21469 (N_21469,N_19763,N_18514);
or U21470 (N_21470,N_18571,N_18049);
xor U21471 (N_21471,N_18548,N_18870);
nand U21472 (N_21472,N_19701,N_18479);
xnor U21473 (N_21473,N_19211,N_18570);
nand U21474 (N_21474,N_19017,N_18479);
or U21475 (N_21475,N_18675,N_19660);
nand U21476 (N_21476,N_19912,N_18814);
or U21477 (N_21477,N_18664,N_19530);
xnor U21478 (N_21478,N_18759,N_18193);
nor U21479 (N_21479,N_18104,N_18390);
xnor U21480 (N_21480,N_18505,N_19406);
or U21481 (N_21481,N_18750,N_18344);
nand U21482 (N_21482,N_19987,N_19777);
xor U21483 (N_21483,N_18760,N_18781);
xor U21484 (N_21484,N_19037,N_19997);
nand U21485 (N_21485,N_18897,N_19624);
or U21486 (N_21486,N_19051,N_18610);
or U21487 (N_21487,N_18162,N_19671);
xor U21488 (N_21488,N_18748,N_19832);
or U21489 (N_21489,N_18056,N_18118);
nor U21490 (N_21490,N_18818,N_19200);
nand U21491 (N_21491,N_18575,N_19253);
nand U21492 (N_21492,N_18093,N_19492);
nand U21493 (N_21493,N_18544,N_18677);
xor U21494 (N_21494,N_18691,N_19520);
nor U21495 (N_21495,N_18180,N_19874);
and U21496 (N_21496,N_19112,N_19114);
nand U21497 (N_21497,N_19180,N_19367);
xnor U21498 (N_21498,N_18397,N_19150);
nor U21499 (N_21499,N_18511,N_19394);
xor U21500 (N_21500,N_18882,N_18267);
nand U21501 (N_21501,N_18055,N_19078);
xnor U21502 (N_21502,N_18540,N_19680);
nor U21503 (N_21503,N_18514,N_18969);
xor U21504 (N_21504,N_18652,N_19924);
or U21505 (N_21505,N_18682,N_18384);
or U21506 (N_21506,N_18534,N_19427);
or U21507 (N_21507,N_18466,N_18858);
nor U21508 (N_21508,N_18995,N_18553);
nor U21509 (N_21509,N_18698,N_19858);
xnor U21510 (N_21510,N_18132,N_18465);
nor U21511 (N_21511,N_19025,N_19383);
nand U21512 (N_21512,N_19412,N_18418);
or U21513 (N_21513,N_19138,N_18354);
and U21514 (N_21514,N_19926,N_18346);
or U21515 (N_21515,N_19629,N_18646);
xor U21516 (N_21516,N_19902,N_19205);
and U21517 (N_21517,N_18493,N_18020);
or U21518 (N_21518,N_19624,N_19949);
xor U21519 (N_21519,N_18267,N_19635);
and U21520 (N_21520,N_19161,N_18432);
and U21521 (N_21521,N_18807,N_18448);
nand U21522 (N_21522,N_19126,N_18620);
or U21523 (N_21523,N_19420,N_19119);
nand U21524 (N_21524,N_19449,N_19726);
and U21525 (N_21525,N_18501,N_18647);
nor U21526 (N_21526,N_19321,N_18997);
and U21527 (N_21527,N_18435,N_19044);
or U21528 (N_21528,N_18539,N_18274);
nor U21529 (N_21529,N_18098,N_19075);
nand U21530 (N_21530,N_19991,N_19184);
xnor U21531 (N_21531,N_18954,N_18246);
and U21532 (N_21532,N_19510,N_19495);
xor U21533 (N_21533,N_18404,N_19202);
or U21534 (N_21534,N_18765,N_19115);
and U21535 (N_21535,N_19304,N_19096);
xnor U21536 (N_21536,N_18884,N_19732);
or U21537 (N_21537,N_19646,N_18848);
or U21538 (N_21538,N_19916,N_19320);
and U21539 (N_21539,N_18533,N_18698);
or U21540 (N_21540,N_19918,N_18920);
or U21541 (N_21541,N_19449,N_19157);
nand U21542 (N_21542,N_18312,N_18394);
and U21543 (N_21543,N_19024,N_18652);
nand U21544 (N_21544,N_18448,N_19332);
nand U21545 (N_21545,N_18612,N_18562);
and U21546 (N_21546,N_19615,N_18892);
nor U21547 (N_21547,N_19016,N_18896);
nand U21548 (N_21548,N_18382,N_18568);
xor U21549 (N_21549,N_19576,N_19025);
xor U21550 (N_21550,N_18264,N_19294);
or U21551 (N_21551,N_19919,N_18522);
nand U21552 (N_21552,N_19420,N_18221);
and U21553 (N_21553,N_18620,N_19375);
nor U21554 (N_21554,N_18143,N_18042);
and U21555 (N_21555,N_18707,N_18020);
xnor U21556 (N_21556,N_19828,N_18115);
nor U21557 (N_21557,N_19524,N_19285);
or U21558 (N_21558,N_19705,N_18951);
nand U21559 (N_21559,N_19257,N_18429);
or U21560 (N_21560,N_18086,N_19759);
and U21561 (N_21561,N_19665,N_18619);
and U21562 (N_21562,N_19470,N_18684);
xor U21563 (N_21563,N_18842,N_18506);
or U21564 (N_21564,N_18265,N_19729);
and U21565 (N_21565,N_19307,N_18014);
nand U21566 (N_21566,N_19669,N_19997);
xor U21567 (N_21567,N_19343,N_19117);
xor U21568 (N_21568,N_19853,N_19361);
and U21569 (N_21569,N_19449,N_19468);
nor U21570 (N_21570,N_19707,N_18680);
and U21571 (N_21571,N_19497,N_19786);
nand U21572 (N_21572,N_18581,N_18219);
nand U21573 (N_21573,N_18398,N_19605);
nand U21574 (N_21574,N_18583,N_18169);
xor U21575 (N_21575,N_19554,N_19709);
xnor U21576 (N_21576,N_19555,N_18936);
xnor U21577 (N_21577,N_18122,N_18561);
nand U21578 (N_21578,N_18087,N_19206);
or U21579 (N_21579,N_19773,N_19284);
nand U21580 (N_21580,N_19940,N_18591);
nand U21581 (N_21581,N_18900,N_19002);
or U21582 (N_21582,N_19691,N_18900);
or U21583 (N_21583,N_18561,N_18570);
nor U21584 (N_21584,N_18206,N_19582);
nor U21585 (N_21585,N_19175,N_18450);
xor U21586 (N_21586,N_19358,N_19624);
nand U21587 (N_21587,N_19038,N_19759);
or U21588 (N_21588,N_18195,N_19979);
nand U21589 (N_21589,N_18860,N_19392);
and U21590 (N_21590,N_18241,N_18479);
nor U21591 (N_21591,N_18738,N_18831);
and U21592 (N_21592,N_19522,N_19598);
and U21593 (N_21593,N_18464,N_19968);
nor U21594 (N_21594,N_19929,N_18689);
or U21595 (N_21595,N_19033,N_18729);
and U21596 (N_21596,N_19856,N_18430);
xnor U21597 (N_21597,N_19069,N_19984);
nand U21598 (N_21598,N_19886,N_19442);
nor U21599 (N_21599,N_19834,N_18545);
nand U21600 (N_21600,N_19086,N_19463);
nand U21601 (N_21601,N_18533,N_19350);
nor U21602 (N_21602,N_18441,N_18892);
xnor U21603 (N_21603,N_18213,N_19682);
nand U21604 (N_21604,N_19469,N_19208);
and U21605 (N_21605,N_18437,N_19140);
or U21606 (N_21606,N_18022,N_18184);
nand U21607 (N_21607,N_19112,N_19047);
or U21608 (N_21608,N_19538,N_19950);
or U21609 (N_21609,N_18540,N_19587);
nor U21610 (N_21610,N_18786,N_18383);
nor U21611 (N_21611,N_19576,N_19630);
xnor U21612 (N_21612,N_19913,N_18710);
and U21613 (N_21613,N_19447,N_19378);
xnor U21614 (N_21614,N_18725,N_19547);
and U21615 (N_21615,N_19614,N_19807);
and U21616 (N_21616,N_18614,N_18372);
nor U21617 (N_21617,N_18828,N_19933);
or U21618 (N_21618,N_19158,N_18716);
nor U21619 (N_21619,N_19776,N_19372);
or U21620 (N_21620,N_18335,N_19387);
nor U21621 (N_21621,N_18123,N_19683);
nor U21622 (N_21622,N_18397,N_19907);
and U21623 (N_21623,N_19798,N_18070);
nand U21624 (N_21624,N_18001,N_18047);
xor U21625 (N_21625,N_19086,N_18274);
or U21626 (N_21626,N_19129,N_18138);
nor U21627 (N_21627,N_18672,N_19513);
xor U21628 (N_21628,N_18743,N_18082);
or U21629 (N_21629,N_18860,N_19178);
nor U21630 (N_21630,N_19324,N_19794);
xor U21631 (N_21631,N_18447,N_18251);
and U21632 (N_21632,N_19164,N_18256);
and U21633 (N_21633,N_19957,N_18971);
nor U21634 (N_21634,N_18158,N_19502);
or U21635 (N_21635,N_18717,N_19186);
nand U21636 (N_21636,N_18566,N_18169);
nor U21637 (N_21637,N_18509,N_19737);
or U21638 (N_21638,N_19855,N_19983);
or U21639 (N_21639,N_18474,N_19935);
or U21640 (N_21640,N_18613,N_19573);
nor U21641 (N_21641,N_18525,N_18795);
or U21642 (N_21642,N_18638,N_18154);
nand U21643 (N_21643,N_19573,N_18208);
and U21644 (N_21644,N_18933,N_18385);
or U21645 (N_21645,N_18697,N_18618);
and U21646 (N_21646,N_18577,N_19053);
nand U21647 (N_21647,N_18618,N_18143);
xor U21648 (N_21648,N_19399,N_19312);
and U21649 (N_21649,N_19804,N_18083);
nand U21650 (N_21650,N_18018,N_19809);
nor U21651 (N_21651,N_19641,N_18580);
and U21652 (N_21652,N_18034,N_18482);
and U21653 (N_21653,N_19003,N_19298);
and U21654 (N_21654,N_18333,N_18280);
or U21655 (N_21655,N_18610,N_19159);
nand U21656 (N_21656,N_19608,N_18738);
nor U21657 (N_21657,N_19350,N_18073);
nor U21658 (N_21658,N_19865,N_18406);
or U21659 (N_21659,N_18240,N_18083);
nor U21660 (N_21660,N_18694,N_18923);
nand U21661 (N_21661,N_19432,N_19060);
xnor U21662 (N_21662,N_19038,N_18973);
nand U21663 (N_21663,N_19561,N_19638);
and U21664 (N_21664,N_19446,N_18556);
and U21665 (N_21665,N_18320,N_18477);
and U21666 (N_21666,N_18359,N_18785);
nand U21667 (N_21667,N_19910,N_19862);
and U21668 (N_21668,N_18497,N_18849);
or U21669 (N_21669,N_19231,N_18456);
and U21670 (N_21670,N_19513,N_19377);
nor U21671 (N_21671,N_18455,N_18509);
xor U21672 (N_21672,N_18283,N_18567);
xnor U21673 (N_21673,N_19533,N_19015);
xnor U21674 (N_21674,N_18768,N_18102);
nand U21675 (N_21675,N_19517,N_19678);
or U21676 (N_21676,N_18734,N_19433);
nor U21677 (N_21677,N_18955,N_19923);
nand U21678 (N_21678,N_18643,N_18123);
xnor U21679 (N_21679,N_18758,N_19742);
or U21680 (N_21680,N_18722,N_18893);
and U21681 (N_21681,N_19230,N_19364);
and U21682 (N_21682,N_19094,N_19451);
nor U21683 (N_21683,N_19167,N_18678);
nor U21684 (N_21684,N_19649,N_19599);
or U21685 (N_21685,N_19993,N_18361);
nand U21686 (N_21686,N_19728,N_18453);
and U21687 (N_21687,N_18079,N_18843);
xor U21688 (N_21688,N_18125,N_19303);
xnor U21689 (N_21689,N_19106,N_19293);
nand U21690 (N_21690,N_18485,N_18114);
and U21691 (N_21691,N_19662,N_18210);
and U21692 (N_21692,N_19464,N_19139);
nand U21693 (N_21693,N_19404,N_18873);
nor U21694 (N_21694,N_18919,N_19693);
nor U21695 (N_21695,N_18253,N_18562);
or U21696 (N_21696,N_18738,N_18502);
nor U21697 (N_21697,N_19967,N_19545);
and U21698 (N_21698,N_18136,N_18022);
and U21699 (N_21699,N_18516,N_18310);
or U21700 (N_21700,N_19972,N_18802);
nand U21701 (N_21701,N_18324,N_19636);
and U21702 (N_21702,N_19994,N_19938);
nor U21703 (N_21703,N_19234,N_18967);
and U21704 (N_21704,N_18110,N_18779);
nand U21705 (N_21705,N_18957,N_18482);
xor U21706 (N_21706,N_18117,N_19917);
nor U21707 (N_21707,N_18191,N_19863);
or U21708 (N_21708,N_18980,N_18113);
or U21709 (N_21709,N_19727,N_19140);
nand U21710 (N_21710,N_18456,N_18920);
nand U21711 (N_21711,N_19862,N_19145);
and U21712 (N_21712,N_19106,N_19495);
xor U21713 (N_21713,N_18729,N_19164);
or U21714 (N_21714,N_19458,N_19622);
or U21715 (N_21715,N_19632,N_19875);
xnor U21716 (N_21716,N_19751,N_18496);
nor U21717 (N_21717,N_19186,N_19189);
or U21718 (N_21718,N_19069,N_19806);
or U21719 (N_21719,N_19314,N_18318);
nand U21720 (N_21720,N_18881,N_18378);
xor U21721 (N_21721,N_19086,N_19758);
nor U21722 (N_21722,N_19091,N_18827);
or U21723 (N_21723,N_19323,N_18196);
and U21724 (N_21724,N_18485,N_18253);
nor U21725 (N_21725,N_18364,N_19701);
nor U21726 (N_21726,N_19921,N_18526);
and U21727 (N_21727,N_19520,N_19481);
nand U21728 (N_21728,N_19791,N_19722);
or U21729 (N_21729,N_18680,N_19141);
and U21730 (N_21730,N_18788,N_18709);
nand U21731 (N_21731,N_19412,N_18466);
nand U21732 (N_21732,N_19663,N_19076);
or U21733 (N_21733,N_18638,N_18558);
and U21734 (N_21734,N_19596,N_19813);
and U21735 (N_21735,N_19975,N_18940);
nor U21736 (N_21736,N_18332,N_18756);
nor U21737 (N_21737,N_19556,N_18359);
nand U21738 (N_21738,N_19112,N_18382);
or U21739 (N_21739,N_18180,N_18108);
and U21740 (N_21740,N_18523,N_18673);
nor U21741 (N_21741,N_19435,N_19788);
or U21742 (N_21742,N_19046,N_19556);
nor U21743 (N_21743,N_18072,N_18859);
nor U21744 (N_21744,N_18399,N_19104);
nand U21745 (N_21745,N_19863,N_18720);
xnor U21746 (N_21746,N_18458,N_19967);
xor U21747 (N_21747,N_19179,N_19905);
xor U21748 (N_21748,N_19806,N_19220);
nor U21749 (N_21749,N_18132,N_19456);
and U21750 (N_21750,N_19965,N_18759);
nor U21751 (N_21751,N_19084,N_18936);
nand U21752 (N_21752,N_18791,N_19923);
nand U21753 (N_21753,N_18769,N_18805);
nand U21754 (N_21754,N_18306,N_18055);
nor U21755 (N_21755,N_18096,N_19188);
xor U21756 (N_21756,N_18462,N_19398);
nor U21757 (N_21757,N_18246,N_19733);
xor U21758 (N_21758,N_19093,N_19868);
and U21759 (N_21759,N_19496,N_18971);
nand U21760 (N_21760,N_18516,N_18475);
xor U21761 (N_21761,N_18577,N_19422);
nand U21762 (N_21762,N_19937,N_19376);
nand U21763 (N_21763,N_18275,N_19388);
nor U21764 (N_21764,N_18107,N_18083);
or U21765 (N_21765,N_18548,N_18481);
nand U21766 (N_21766,N_19519,N_19595);
or U21767 (N_21767,N_19679,N_18672);
or U21768 (N_21768,N_19911,N_18281);
and U21769 (N_21769,N_18327,N_18567);
or U21770 (N_21770,N_18717,N_18269);
nand U21771 (N_21771,N_19305,N_19922);
or U21772 (N_21772,N_19091,N_19093);
nand U21773 (N_21773,N_18977,N_19866);
or U21774 (N_21774,N_19994,N_18384);
nor U21775 (N_21775,N_18111,N_18387);
and U21776 (N_21776,N_18864,N_18055);
or U21777 (N_21777,N_18164,N_19331);
xor U21778 (N_21778,N_19466,N_19441);
and U21779 (N_21779,N_19800,N_18855);
xor U21780 (N_21780,N_19254,N_19659);
and U21781 (N_21781,N_18893,N_19102);
nand U21782 (N_21782,N_18448,N_18515);
nor U21783 (N_21783,N_19641,N_18697);
and U21784 (N_21784,N_18928,N_18907);
nand U21785 (N_21785,N_19193,N_18911);
and U21786 (N_21786,N_18317,N_19735);
nand U21787 (N_21787,N_18421,N_19032);
xnor U21788 (N_21788,N_18433,N_19677);
and U21789 (N_21789,N_18083,N_18769);
and U21790 (N_21790,N_19369,N_18300);
xor U21791 (N_21791,N_19600,N_19578);
nand U21792 (N_21792,N_18157,N_19758);
xnor U21793 (N_21793,N_18024,N_19502);
nand U21794 (N_21794,N_19845,N_18300);
nand U21795 (N_21795,N_19363,N_19376);
nand U21796 (N_21796,N_18733,N_18962);
or U21797 (N_21797,N_19952,N_19574);
nor U21798 (N_21798,N_19466,N_18200);
or U21799 (N_21799,N_19518,N_19114);
nand U21800 (N_21800,N_18950,N_18806);
xnor U21801 (N_21801,N_18646,N_18051);
nand U21802 (N_21802,N_19434,N_19785);
and U21803 (N_21803,N_18131,N_18662);
or U21804 (N_21804,N_18414,N_18037);
or U21805 (N_21805,N_18057,N_18160);
and U21806 (N_21806,N_19983,N_18406);
xor U21807 (N_21807,N_18658,N_19043);
and U21808 (N_21808,N_18264,N_19458);
nand U21809 (N_21809,N_18750,N_19995);
or U21810 (N_21810,N_18742,N_18951);
and U21811 (N_21811,N_19744,N_18939);
or U21812 (N_21812,N_19967,N_19164);
xnor U21813 (N_21813,N_19068,N_18946);
nand U21814 (N_21814,N_19609,N_19583);
or U21815 (N_21815,N_19809,N_19734);
and U21816 (N_21816,N_19552,N_18989);
nand U21817 (N_21817,N_18063,N_18260);
or U21818 (N_21818,N_19352,N_19362);
or U21819 (N_21819,N_19469,N_19404);
or U21820 (N_21820,N_18426,N_18548);
nor U21821 (N_21821,N_19932,N_18946);
xor U21822 (N_21822,N_19814,N_19538);
xor U21823 (N_21823,N_18707,N_19093);
or U21824 (N_21824,N_18537,N_18890);
or U21825 (N_21825,N_18737,N_19947);
and U21826 (N_21826,N_19255,N_18392);
and U21827 (N_21827,N_18638,N_18425);
nor U21828 (N_21828,N_19666,N_18610);
nand U21829 (N_21829,N_19071,N_18659);
nor U21830 (N_21830,N_18464,N_19715);
and U21831 (N_21831,N_19451,N_18894);
nor U21832 (N_21832,N_18556,N_18080);
or U21833 (N_21833,N_18473,N_18216);
xnor U21834 (N_21834,N_19133,N_18924);
xor U21835 (N_21835,N_19700,N_18843);
or U21836 (N_21836,N_19947,N_19684);
and U21837 (N_21837,N_18859,N_18280);
and U21838 (N_21838,N_19573,N_18331);
nor U21839 (N_21839,N_19291,N_19744);
and U21840 (N_21840,N_18929,N_19791);
nor U21841 (N_21841,N_18514,N_19810);
nand U21842 (N_21842,N_19224,N_18312);
or U21843 (N_21843,N_18970,N_18831);
or U21844 (N_21844,N_19571,N_18409);
xnor U21845 (N_21845,N_19644,N_18703);
nor U21846 (N_21846,N_18732,N_19387);
and U21847 (N_21847,N_19109,N_19358);
nor U21848 (N_21848,N_18974,N_19243);
xor U21849 (N_21849,N_19059,N_19310);
nand U21850 (N_21850,N_19926,N_19006);
nor U21851 (N_21851,N_19382,N_19269);
nor U21852 (N_21852,N_18765,N_19451);
nor U21853 (N_21853,N_19499,N_19884);
or U21854 (N_21854,N_19641,N_18470);
nand U21855 (N_21855,N_19427,N_19280);
xnor U21856 (N_21856,N_18376,N_18897);
or U21857 (N_21857,N_19825,N_19058);
nor U21858 (N_21858,N_19713,N_19124);
nor U21859 (N_21859,N_19607,N_19550);
nand U21860 (N_21860,N_18172,N_19081);
nor U21861 (N_21861,N_19123,N_18397);
nor U21862 (N_21862,N_19045,N_18733);
or U21863 (N_21863,N_18652,N_18713);
and U21864 (N_21864,N_18734,N_18837);
or U21865 (N_21865,N_19043,N_19514);
or U21866 (N_21866,N_19170,N_18816);
nand U21867 (N_21867,N_19185,N_19330);
nor U21868 (N_21868,N_18674,N_19425);
nand U21869 (N_21869,N_18802,N_18399);
nand U21870 (N_21870,N_18208,N_19095);
nor U21871 (N_21871,N_19882,N_19572);
or U21872 (N_21872,N_18779,N_18452);
and U21873 (N_21873,N_19795,N_19104);
and U21874 (N_21874,N_18043,N_19691);
and U21875 (N_21875,N_18095,N_18113);
nor U21876 (N_21876,N_19734,N_19302);
or U21877 (N_21877,N_18032,N_19963);
nand U21878 (N_21878,N_18638,N_19559);
nor U21879 (N_21879,N_18931,N_18078);
nand U21880 (N_21880,N_18498,N_18787);
nand U21881 (N_21881,N_19655,N_19275);
xor U21882 (N_21882,N_19842,N_19359);
nand U21883 (N_21883,N_18458,N_18994);
and U21884 (N_21884,N_18184,N_19961);
xor U21885 (N_21885,N_18481,N_19217);
xor U21886 (N_21886,N_19802,N_18782);
or U21887 (N_21887,N_19117,N_19928);
or U21888 (N_21888,N_19740,N_18820);
xor U21889 (N_21889,N_19786,N_19754);
or U21890 (N_21890,N_18987,N_19927);
or U21891 (N_21891,N_18784,N_18571);
xor U21892 (N_21892,N_19555,N_19297);
xor U21893 (N_21893,N_19181,N_18640);
nand U21894 (N_21894,N_18297,N_18788);
nand U21895 (N_21895,N_18481,N_18504);
xor U21896 (N_21896,N_18200,N_18366);
nor U21897 (N_21897,N_18706,N_18491);
or U21898 (N_21898,N_19167,N_18376);
nand U21899 (N_21899,N_18971,N_18892);
nand U21900 (N_21900,N_18138,N_19124);
nor U21901 (N_21901,N_19437,N_18218);
nor U21902 (N_21902,N_18629,N_18239);
or U21903 (N_21903,N_18624,N_18473);
and U21904 (N_21904,N_19713,N_19468);
or U21905 (N_21905,N_18791,N_18302);
nor U21906 (N_21906,N_18516,N_18105);
nand U21907 (N_21907,N_18011,N_18082);
nand U21908 (N_21908,N_19209,N_18712);
nor U21909 (N_21909,N_18555,N_19467);
xnor U21910 (N_21910,N_18126,N_18128);
and U21911 (N_21911,N_19720,N_19033);
and U21912 (N_21912,N_19328,N_18815);
xnor U21913 (N_21913,N_18757,N_18826);
xor U21914 (N_21914,N_18500,N_18726);
nor U21915 (N_21915,N_19408,N_19888);
xnor U21916 (N_21916,N_19687,N_19247);
nand U21917 (N_21917,N_18594,N_18323);
or U21918 (N_21918,N_19757,N_18392);
xor U21919 (N_21919,N_18422,N_18923);
nand U21920 (N_21920,N_19391,N_18036);
nand U21921 (N_21921,N_18148,N_19574);
nor U21922 (N_21922,N_19260,N_19102);
xor U21923 (N_21923,N_19931,N_18380);
nand U21924 (N_21924,N_18227,N_19826);
or U21925 (N_21925,N_19108,N_18138);
and U21926 (N_21926,N_19245,N_19026);
nor U21927 (N_21927,N_18501,N_19502);
xor U21928 (N_21928,N_19508,N_18613);
or U21929 (N_21929,N_19291,N_19380);
or U21930 (N_21930,N_19022,N_18177);
and U21931 (N_21931,N_19741,N_18880);
or U21932 (N_21932,N_19241,N_19902);
nor U21933 (N_21933,N_19522,N_19877);
nand U21934 (N_21934,N_19937,N_18075);
or U21935 (N_21935,N_18380,N_18103);
nand U21936 (N_21936,N_19308,N_18752);
and U21937 (N_21937,N_19081,N_18501);
or U21938 (N_21938,N_18163,N_18580);
xor U21939 (N_21939,N_18353,N_19070);
or U21940 (N_21940,N_19056,N_19159);
nor U21941 (N_21941,N_18683,N_19987);
xor U21942 (N_21942,N_19276,N_19440);
nor U21943 (N_21943,N_19411,N_18252);
nand U21944 (N_21944,N_18325,N_18526);
nor U21945 (N_21945,N_18557,N_19048);
or U21946 (N_21946,N_18533,N_18276);
xnor U21947 (N_21947,N_19581,N_18241);
and U21948 (N_21948,N_19284,N_19313);
or U21949 (N_21949,N_18241,N_18292);
and U21950 (N_21950,N_18342,N_19193);
nor U21951 (N_21951,N_19736,N_18394);
nand U21952 (N_21952,N_19743,N_19376);
and U21953 (N_21953,N_18119,N_19770);
xnor U21954 (N_21954,N_19866,N_18209);
nand U21955 (N_21955,N_19893,N_18293);
nand U21956 (N_21956,N_19317,N_18299);
nand U21957 (N_21957,N_18261,N_19803);
nor U21958 (N_21958,N_18514,N_19022);
nand U21959 (N_21959,N_19737,N_18916);
nor U21960 (N_21960,N_19551,N_19285);
and U21961 (N_21961,N_18283,N_18207);
xnor U21962 (N_21962,N_19802,N_19064);
nand U21963 (N_21963,N_18226,N_19514);
and U21964 (N_21964,N_19769,N_18859);
nand U21965 (N_21965,N_18250,N_19466);
nand U21966 (N_21966,N_19517,N_19866);
nand U21967 (N_21967,N_19838,N_19109);
or U21968 (N_21968,N_19809,N_19723);
nand U21969 (N_21969,N_19152,N_18228);
nor U21970 (N_21970,N_19374,N_19488);
nor U21971 (N_21971,N_18542,N_19470);
nand U21972 (N_21972,N_19626,N_18197);
nor U21973 (N_21973,N_19285,N_19682);
nor U21974 (N_21974,N_18537,N_19826);
or U21975 (N_21975,N_18435,N_19551);
and U21976 (N_21976,N_19282,N_18578);
nand U21977 (N_21977,N_19226,N_19509);
xor U21978 (N_21978,N_18177,N_18846);
and U21979 (N_21979,N_18391,N_18668);
xnor U21980 (N_21980,N_19237,N_18026);
or U21981 (N_21981,N_18731,N_18639);
xor U21982 (N_21982,N_18036,N_19256);
nor U21983 (N_21983,N_19379,N_18216);
or U21984 (N_21984,N_18017,N_18687);
or U21985 (N_21985,N_19626,N_18195);
xor U21986 (N_21986,N_19220,N_18392);
and U21987 (N_21987,N_18843,N_19033);
or U21988 (N_21988,N_18023,N_18442);
nand U21989 (N_21989,N_19269,N_18164);
nand U21990 (N_21990,N_18252,N_19401);
and U21991 (N_21991,N_19692,N_19993);
nand U21992 (N_21992,N_19525,N_18755);
nand U21993 (N_21993,N_19509,N_18747);
nor U21994 (N_21994,N_18773,N_19039);
or U21995 (N_21995,N_19678,N_19639);
nor U21996 (N_21996,N_19224,N_18350);
xnor U21997 (N_21997,N_18516,N_19281);
and U21998 (N_21998,N_19113,N_18273);
and U21999 (N_21999,N_19893,N_18007);
nor U22000 (N_22000,N_20920,N_20633);
or U22001 (N_22001,N_20083,N_20637);
and U22002 (N_22002,N_21061,N_20426);
xor U22003 (N_22003,N_21157,N_21120);
and U22004 (N_22004,N_20794,N_20451);
nand U22005 (N_22005,N_20846,N_21555);
nand U22006 (N_22006,N_20461,N_20068);
xor U22007 (N_22007,N_21199,N_21067);
nor U22008 (N_22008,N_21860,N_20375);
nor U22009 (N_22009,N_21978,N_21069);
nor U22010 (N_22010,N_20561,N_21723);
and U22011 (N_22011,N_20191,N_20378);
nor U22012 (N_22012,N_21689,N_21164);
nor U22013 (N_22013,N_20285,N_20389);
or U22014 (N_22014,N_20326,N_21329);
xnor U22015 (N_22015,N_20455,N_21317);
nor U22016 (N_22016,N_21380,N_21141);
nand U22017 (N_22017,N_20419,N_21287);
nand U22018 (N_22018,N_21298,N_20799);
nand U22019 (N_22019,N_20614,N_20370);
or U22020 (N_22020,N_21919,N_21969);
and U22021 (N_22021,N_21290,N_21614);
and U22022 (N_22022,N_20296,N_20317);
xor U22023 (N_22023,N_20662,N_21535);
nor U22024 (N_22024,N_20825,N_21872);
xnor U22025 (N_22025,N_21558,N_21469);
xor U22026 (N_22026,N_21055,N_20893);
xor U22027 (N_22027,N_21642,N_21001);
or U22028 (N_22028,N_21678,N_21637);
or U22029 (N_22029,N_20157,N_21435);
xor U22030 (N_22030,N_21064,N_20175);
nand U22031 (N_22031,N_21753,N_20705);
nand U22032 (N_22032,N_20536,N_20025);
or U22033 (N_22033,N_21700,N_20756);
xnor U22034 (N_22034,N_20562,N_21022);
or U22035 (N_22035,N_21262,N_21253);
nor U22036 (N_22036,N_21887,N_20476);
and U22037 (N_22037,N_20380,N_20650);
xor U22038 (N_22038,N_20813,N_20257);
and U22039 (N_22039,N_21395,N_21673);
nand U22040 (N_22040,N_20119,N_21154);
nand U22041 (N_22041,N_21431,N_20155);
xor U22042 (N_22042,N_20167,N_21534);
or U22043 (N_22043,N_20140,N_20356);
xnor U22044 (N_22044,N_20982,N_21994);
nand U22045 (N_22045,N_20355,N_21252);
and U22046 (N_22046,N_20905,N_20332);
and U22047 (N_22047,N_20160,N_20070);
and U22048 (N_22048,N_20395,N_20703);
nand U22049 (N_22049,N_21636,N_21100);
xor U22050 (N_22050,N_21714,N_20887);
nand U22051 (N_22051,N_20979,N_21312);
nand U22052 (N_22052,N_20344,N_21268);
nand U22053 (N_22053,N_21722,N_21648);
nor U22054 (N_22054,N_21833,N_21118);
nor U22055 (N_22055,N_20172,N_21800);
and U22056 (N_22056,N_21852,N_20425);
and U22057 (N_22057,N_20037,N_20351);
nand U22058 (N_22058,N_20041,N_20886);
xor U22059 (N_22059,N_20774,N_20897);
or U22060 (N_22060,N_21039,N_21237);
nand U22061 (N_22061,N_21938,N_20837);
nor U22062 (N_22062,N_21146,N_21179);
and U22063 (N_22063,N_21606,N_21956);
and U22064 (N_22064,N_20619,N_21948);
and U22065 (N_22065,N_20605,N_21242);
and U22066 (N_22066,N_21200,N_20544);
nand U22067 (N_22067,N_20632,N_21779);
nor U22068 (N_22068,N_20929,N_20401);
xor U22069 (N_22069,N_21822,N_21145);
nor U22070 (N_22070,N_20361,N_21964);
xor U22071 (N_22071,N_21679,N_21041);
and U22072 (N_22072,N_21984,N_20875);
nand U22073 (N_22073,N_20953,N_21198);
and U22074 (N_22074,N_21805,N_20397);
xnor U22075 (N_22075,N_21304,N_21052);
or U22076 (N_22076,N_20655,N_20470);
or U22077 (N_22077,N_20610,N_20376);
or U22078 (N_22078,N_20696,N_20797);
xor U22079 (N_22079,N_20453,N_21615);
or U22080 (N_22080,N_21772,N_20881);
or U22081 (N_22081,N_20024,N_21485);
nand U22082 (N_22082,N_21197,N_21655);
and U22083 (N_22083,N_21131,N_21657);
nand U22084 (N_22084,N_21214,N_21296);
xor U22085 (N_22085,N_21128,N_21640);
and U22086 (N_22086,N_21213,N_20940);
nand U22087 (N_22087,N_20579,N_21040);
and U22088 (N_22088,N_20008,N_21260);
or U22089 (N_22089,N_20297,N_21479);
or U22090 (N_22090,N_21092,N_20729);
xnor U22091 (N_22091,N_21936,N_20670);
nand U22092 (N_22092,N_21488,N_21434);
nor U22093 (N_22093,N_21433,N_20082);
xnor U22094 (N_22094,N_21259,N_21263);
xor U22095 (N_22095,N_20842,N_21907);
nand U22096 (N_22096,N_21160,N_20934);
nand U22097 (N_22097,N_20429,N_21560);
xnor U22098 (N_22098,N_21927,N_21357);
nand U22099 (N_22099,N_21439,N_21997);
nor U22100 (N_22100,N_20485,N_20061);
or U22101 (N_22101,N_20494,N_21085);
nor U22102 (N_22102,N_21462,N_20118);
nor U22103 (N_22103,N_20381,N_21114);
nor U22104 (N_22104,N_21946,N_20987);
and U22105 (N_22105,N_20968,N_21084);
nand U22106 (N_22106,N_21397,N_21788);
or U22107 (N_22107,N_21804,N_21945);
nand U22108 (N_22108,N_20798,N_20036);
nand U22109 (N_22109,N_21882,N_21471);
and U22110 (N_22110,N_20221,N_21587);
or U22111 (N_22111,N_20993,N_21011);
nand U22112 (N_22112,N_20571,N_20568);
nor U22113 (N_22113,N_21775,N_20438);
and U22114 (N_22114,N_20151,N_21241);
nand U22115 (N_22115,N_21638,N_20598);
nor U22116 (N_22116,N_20829,N_21531);
and U22117 (N_22117,N_21266,N_21561);
and U22118 (N_22118,N_20618,N_21697);
or U22119 (N_22119,N_20391,N_21342);
xor U22120 (N_22120,N_21062,N_21631);
nor U22121 (N_22121,N_21047,N_20955);
nor U22122 (N_22122,N_20984,N_21668);
nor U22123 (N_22123,N_20279,N_20806);
nand U22124 (N_22124,N_21592,N_20314);
nor U22125 (N_22125,N_21992,N_20882);
or U22126 (N_22126,N_21617,N_20033);
nand U22127 (N_22127,N_21542,N_21742);
or U22128 (N_22128,N_20493,N_21325);
xnor U22129 (N_22129,N_20246,N_21720);
xnor U22130 (N_22130,N_20908,N_21906);
and U22131 (N_22131,N_20564,N_20647);
or U22132 (N_22132,N_21201,N_21184);
nor U22133 (N_22133,N_20029,N_21394);
nand U22134 (N_22134,N_21239,N_20657);
and U22135 (N_22135,N_20345,N_21499);
xnor U22136 (N_22136,N_21327,N_21578);
and U22137 (N_22137,N_20138,N_20683);
xnor U22138 (N_22138,N_20002,N_21959);
or U22139 (N_22139,N_21427,N_20767);
and U22140 (N_22140,N_21862,N_21600);
and U22141 (N_22141,N_20126,N_20810);
nor U22142 (N_22142,N_21144,N_21713);
or U22143 (N_22143,N_20613,N_20483);
xnor U22144 (N_22144,N_21096,N_21349);
xor U22145 (N_22145,N_21225,N_20511);
nand U22146 (N_22146,N_20522,N_21937);
nand U22147 (N_22147,N_20324,N_20856);
nand U22148 (N_22148,N_20256,N_20871);
nor U22149 (N_22149,N_21307,N_20185);
and U22150 (N_22150,N_21299,N_21653);
nor U22151 (N_22151,N_20125,N_20433);
or U22152 (N_22152,N_21760,N_20414);
nor U22153 (N_22153,N_20520,N_20689);
nor U22154 (N_22154,N_21492,N_20552);
nor U22155 (N_22155,N_21687,N_20134);
nand U22156 (N_22156,N_21113,N_21140);
nor U22157 (N_22157,N_20644,N_21091);
and U22158 (N_22158,N_21767,N_20665);
and U22159 (N_22159,N_21831,N_21894);
or U22160 (N_22160,N_21962,N_20964);
nand U22161 (N_22161,N_21740,N_20708);
nor U22162 (N_22162,N_20570,N_20555);
xor U22163 (N_22163,N_21725,N_21881);
nand U22164 (N_22164,N_20962,N_21010);
nand U22165 (N_22165,N_20109,N_20527);
nor U22166 (N_22166,N_21690,N_20442);
or U22167 (N_22167,N_21686,N_21777);
nand U22168 (N_22168,N_21811,N_21078);
and U22169 (N_22169,N_20745,N_21633);
and U22170 (N_22170,N_20468,N_21981);
and U22171 (N_22171,N_21098,N_21979);
nor U22172 (N_22172,N_21147,N_20830);
and U22173 (N_22173,N_20075,N_21019);
xnor U22174 (N_22174,N_20459,N_21621);
nor U22175 (N_22175,N_20092,N_21797);
or U22176 (N_22176,N_20275,N_21837);
and U22177 (N_22177,N_21383,N_20110);
and U22178 (N_22178,N_21014,N_21584);
or U22179 (N_22179,N_20251,N_20349);
nor U22180 (N_22180,N_20835,N_20688);
xor U22181 (N_22181,N_21544,N_20515);
nor U22182 (N_22182,N_20178,N_21889);
nor U22183 (N_22183,N_20482,N_21046);
xor U22184 (N_22184,N_20142,N_21088);
nor U22185 (N_22185,N_21413,N_20712);
or U22186 (N_22186,N_20194,N_21191);
nor U22187 (N_22187,N_21366,N_20867);
nand U22188 (N_22188,N_21798,N_20937);
and U22189 (N_22189,N_21130,N_20150);
or U22190 (N_22190,N_21824,N_21963);
xnor U22191 (N_22191,N_20874,N_21481);
xnor U22192 (N_22192,N_21842,N_21138);
or U22193 (N_22193,N_21372,N_21928);
or U22194 (N_22194,N_21955,N_20081);
or U22195 (N_22195,N_21202,N_20519);
and U22196 (N_22196,N_21746,N_20186);
nor U22197 (N_22197,N_21109,N_20546);
or U22198 (N_22198,N_20864,N_20305);
xnor U22199 (N_22199,N_20673,N_20888);
or U22200 (N_22200,N_20838,N_20087);
or U22201 (N_22201,N_20720,N_20101);
and U22202 (N_22202,N_21368,N_21156);
and U22203 (N_22203,N_20898,N_20006);
nor U22204 (N_22204,N_20437,N_20085);
or U22205 (N_22205,N_20402,N_21950);
nor U22206 (N_22206,N_21111,N_21459);
and U22207 (N_22207,N_20734,N_20566);
nor U22208 (N_22208,N_20427,N_21495);
nor U22209 (N_22209,N_21170,N_20135);
xor U22210 (N_22210,N_21731,N_20592);
xnor U22211 (N_22211,N_21283,N_21497);
and U22212 (N_22212,N_20959,N_21574);
or U22213 (N_22213,N_20034,N_21051);
or U22214 (N_22214,N_21878,N_21244);
xnor U22215 (N_22215,N_20280,N_21013);
nor U22216 (N_22216,N_20885,N_20911);
nor U22217 (N_22217,N_20469,N_20782);
or U22218 (N_22218,N_20889,N_21579);
xor U22219 (N_22219,N_21134,N_20554);
nor U22220 (N_22220,N_20728,N_21384);
and U22221 (N_22221,N_21604,N_20058);
nor U22222 (N_22222,N_21338,N_21404);
xor U22223 (N_22223,N_20685,N_21457);
nand U22224 (N_22224,N_21566,N_21119);
or U22225 (N_22225,N_20393,N_20909);
xnor U22226 (N_22226,N_20635,N_21626);
and U22227 (N_22227,N_20558,N_21487);
nor U22228 (N_22228,N_21038,N_21844);
xnor U22229 (N_22229,N_20047,N_20541);
and U22230 (N_22230,N_21733,N_21515);
nor U22231 (N_22231,N_20211,N_21719);
and U22232 (N_22232,N_20724,N_21980);
or U22233 (N_22233,N_20112,N_21449);
nor U22234 (N_22234,N_21958,N_21988);
or U22235 (N_22235,N_21549,N_21786);
nand U22236 (N_22236,N_21059,N_21738);
or U22237 (N_22237,N_21890,N_20241);
and U22238 (N_22238,N_20809,N_21972);
and U22239 (N_22239,N_21586,N_21993);
nand U22240 (N_22240,N_21175,N_21904);
nand U22241 (N_22241,N_21908,N_21974);
and U22242 (N_22242,N_21539,N_21694);
nor U22243 (N_22243,N_20475,N_21334);
xnor U22244 (N_22244,N_21909,N_20026);
nor U22245 (N_22245,N_20808,N_20583);
xnor U22246 (N_22246,N_21185,N_20607);
xnor U22247 (N_22247,N_21647,N_20660);
xor U22248 (N_22248,N_20018,N_21356);
nor U22249 (N_22249,N_21828,N_20050);
nor U22250 (N_22250,N_21153,N_20702);
or U22251 (N_22251,N_20051,N_21400);
xor U22252 (N_22252,N_20645,N_21095);
or U22253 (N_22253,N_21149,N_21503);
or U22254 (N_22254,N_21483,N_20823);
nor U22255 (N_22255,N_21744,N_20396);
xor U22256 (N_22256,N_20141,N_20652);
xnor U22257 (N_22257,N_21204,N_20741);
nor U22258 (N_22258,N_21875,N_20323);
xor U22259 (N_22259,N_20342,N_21684);
nand U22260 (N_22260,N_21514,N_20479);
nor U22261 (N_22261,N_21915,N_20139);
and U22262 (N_22262,N_21220,N_20740);
nor U22263 (N_22263,N_20406,N_21231);
and U22264 (N_22264,N_20096,N_21521);
nor U22265 (N_22265,N_21794,N_21171);
xnor U22266 (N_22266,N_20748,N_20298);
xnor U22267 (N_22267,N_21953,N_21169);
nand U22268 (N_22268,N_20307,N_20352);
nand U22269 (N_22269,N_20668,N_21219);
xnor U22270 (N_22270,N_20675,N_21311);
and U22271 (N_22271,N_20590,N_21581);
xnor U22272 (N_22272,N_21387,N_20236);
nand U22273 (N_22273,N_21174,N_20099);
nand U22274 (N_22274,N_21693,N_21925);
or U22275 (N_22275,N_21821,N_20732);
xnor U22276 (N_22276,N_20507,N_20073);
nor U22277 (N_22277,N_20980,N_21310);
nor U22278 (N_22278,N_21105,N_21303);
or U22279 (N_22279,N_21099,N_20289);
xor U22280 (N_22280,N_20625,N_20664);
nor U22281 (N_22281,N_20303,N_20248);
nor U22282 (N_22282,N_20616,N_21522);
nor U22283 (N_22283,N_21801,N_21865);
nor U22284 (N_22284,N_21309,N_21627);
xor U22285 (N_22285,N_20832,N_20173);
or U22286 (N_22286,N_21278,N_20327);
nand U22287 (N_22287,N_21123,N_20384);
nand U22288 (N_22288,N_21461,N_21257);
and U22289 (N_22289,N_21848,N_20300);
and U22290 (N_22290,N_20709,N_21256);
nor U22291 (N_22291,N_20472,N_21618);
nor U22292 (N_22292,N_21757,N_21264);
or U22293 (N_22293,N_20267,N_20222);
nor U22294 (N_22294,N_20557,N_20563);
or U22295 (N_22295,N_20517,N_21269);
and U22296 (N_22296,N_21795,N_20834);
or U22297 (N_22297,N_20772,N_20430);
nand U22298 (N_22298,N_21077,N_20264);
nand U22299 (N_22299,N_21122,N_21208);
or U22300 (N_22300,N_20462,N_21331);
xnor U22301 (N_22301,N_20080,N_20692);
or U22302 (N_22302,N_20952,N_21892);
nor U22303 (N_22303,N_21705,N_21437);
nor U22304 (N_22304,N_20115,N_21300);
or U22305 (N_22305,N_21289,N_21093);
xnor U22306 (N_22306,N_21851,N_20739);
xnor U22307 (N_22307,N_21859,N_20777);
nor U22308 (N_22308,N_21158,N_21048);
and U22309 (N_22309,N_20775,N_21820);
nor U22310 (N_22310,N_20106,N_21918);
nand U22311 (N_22311,N_21594,N_21065);
and U22312 (N_22312,N_20977,N_21165);
xor U22313 (N_22313,N_21405,N_20945);
or U22314 (N_22314,N_20330,N_21965);
nor U22315 (N_22315,N_20052,N_20725);
or U22316 (N_22316,N_21335,N_21768);
nand U22317 (N_22317,N_20181,N_20481);
nor U22318 (N_22318,N_20053,N_21546);
and U22319 (N_22319,N_20713,N_20946);
nor U22320 (N_22320,N_21599,N_21698);
and U22321 (N_22321,N_21590,N_20512);
and U22322 (N_22322,N_20346,N_20184);
or U22323 (N_22323,N_20918,N_21447);
or U22324 (N_22324,N_20770,N_20902);
xor U22325 (N_22325,N_20254,N_21454);
nand U22326 (N_22326,N_20045,N_21796);
nor U22327 (N_22327,N_21502,N_20271);
xor U22328 (N_22328,N_20362,N_20622);
nor U22329 (N_22329,N_21739,N_21094);
and U22330 (N_22330,N_20572,N_20363);
xnor U22331 (N_22331,N_20667,N_21444);
and U22332 (N_22332,N_20210,N_20228);
nor U22333 (N_22333,N_21498,N_20319);
nand U22334 (N_22334,N_21803,N_20177);
or U22335 (N_22335,N_21110,N_21491);
and U22336 (N_22336,N_21205,N_21931);
nor U22337 (N_22337,N_21658,N_20057);
or U22338 (N_22338,N_21871,N_20392);
xnor U22339 (N_22339,N_20484,N_20761);
nand U22340 (N_22340,N_20726,N_20405);
nor U22341 (N_22341,N_21752,N_21006);
or U22342 (N_22342,N_21846,N_20532);
nor U22343 (N_22343,N_21509,N_20016);
xnor U22344 (N_22344,N_20857,N_21629);
nor U22345 (N_22345,N_20743,N_21417);
or U22346 (N_22346,N_21605,N_20957);
and U22347 (N_22347,N_21445,N_21090);
nand U22348 (N_22348,N_21947,N_20730);
or U22349 (N_22349,N_20258,N_21027);
nand U22350 (N_22350,N_21553,N_20684);
xnor U22351 (N_22351,N_20860,N_20078);
or U22352 (N_22352,N_21050,N_21858);
or U22353 (N_22353,N_21438,N_20366);
or U22354 (N_22354,N_20338,N_21359);
xnor U22355 (N_22355,N_21216,N_20997);
xor U22356 (N_22356,N_20400,N_21070);
nand U22357 (N_22357,N_20498,N_21369);
nor U22358 (N_22358,N_20711,N_21762);
xnor U22359 (N_22359,N_21576,N_21301);
xnor U22360 (N_22360,N_21813,N_20436);
nand U22361 (N_22361,N_21362,N_20521);
nand U22362 (N_22362,N_21996,N_20649);
xnor U22363 (N_22363,N_21814,N_20434);
and U22364 (N_22364,N_20615,N_20269);
or U22365 (N_22365,N_21044,N_20360);
and U22366 (N_22366,N_20274,N_21624);
or U22367 (N_22367,N_21643,N_20506);
nor U22368 (N_22368,N_20152,N_21973);
and U22369 (N_22369,N_21832,N_20411);
xnor U22370 (N_22370,N_20093,N_20913);
nor U22371 (N_22371,N_20304,N_21913);
nand U22372 (N_22372,N_21823,N_21516);
nor U22373 (N_22373,N_20930,N_20877);
or U22374 (N_22374,N_20503,N_20721);
xnor U22375 (N_22375,N_21364,N_21328);
or U22376 (N_22376,N_21215,N_21810);
and U22377 (N_22377,N_21282,N_21494);
xor U22378 (N_22378,N_20648,N_20188);
xnor U22379 (N_22379,N_20373,N_20900);
or U22380 (N_22380,N_21506,N_20315);
and U22381 (N_22381,N_20293,N_20238);
xor U22382 (N_22382,N_20364,N_20233);
and U22383 (N_22383,N_20680,N_21607);
xnor U22384 (N_22384,N_21363,N_20738);
nand U22385 (N_22385,N_21224,N_20672);
and U22386 (N_22386,N_20003,N_21025);
or U22387 (N_22387,N_20714,N_20883);
xnor U22388 (N_22388,N_20535,N_21567);
and U22389 (N_22389,N_21068,N_20477);
xor U22390 (N_22390,N_21505,N_21408);
nor U22391 (N_22391,N_21007,N_21281);
nand U22392 (N_22392,N_21670,N_20377);
and U22393 (N_22393,N_20587,N_21452);
xnor U22394 (N_22394,N_20731,N_21385);
or U22395 (N_22395,N_21843,N_20801);
nand U22396 (N_22396,N_21559,N_20956);
and U22397 (N_22397,N_20056,N_21911);
nor U22398 (N_22398,N_21671,N_20145);
nand U22399 (N_22399,N_21735,N_21270);
or U22400 (N_22400,N_20634,N_21773);
nor U22401 (N_22401,N_20754,N_20795);
or U22402 (N_22402,N_20146,N_20450);
nor U22403 (N_22403,N_20128,N_21030);
or U22404 (N_22404,N_21511,N_21707);
nor U22405 (N_22405,N_20223,N_20944);
nor U22406 (N_22406,N_21751,N_20925);
nand U22407 (N_22407,N_21337,N_21883);
nor U22408 (N_22408,N_21769,N_20624);
nand U22409 (N_22409,N_21961,N_20951);
or U22410 (N_22410,N_20302,N_20369);
nand U22411 (N_22411,N_20578,N_21275);
and U22412 (N_22412,N_20490,N_21935);
xnor U22413 (N_22413,N_20677,N_21692);
xor U22414 (N_22414,N_21489,N_20884);
and U22415 (N_22415,N_20910,N_20408);
nor U22416 (N_22416,N_21473,N_21551);
and U22417 (N_22417,N_20965,N_21023);
or U22418 (N_22418,N_20213,N_20382);
nor U22419 (N_22419,N_21021,N_21162);
nor U22420 (N_22420,N_20687,N_21343);
nand U22421 (N_22421,N_21957,N_20460);
or U22422 (N_22422,N_21125,N_20240);
and U22423 (N_22423,N_21132,N_21856);
or U22424 (N_22424,N_21152,N_21401);
or U22425 (N_22425,N_20591,N_21058);
xor U22426 (N_22426,N_21480,N_20876);
xor U22427 (N_22427,N_21718,N_20394);
nor U22428 (N_22428,N_21227,N_21054);
and U22429 (N_22429,N_20301,N_20379);
nand U22430 (N_22430,N_20963,N_20387);
nor U22431 (N_22431,N_20077,N_21172);
and U22432 (N_22432,N_21180,N_21209);
and U22433 (N_22433,N_21819,N_21274);
nor U22434 (N_22434,N_20499,N_20784);
xor U22435 (N_22435,N_20757,N_20901);
xor U22436 (N_22436,N_21129,N_20147);
and U22437 (N_22437,N_20844,N_21748);
or U22438 (N_22438,N_21650,N_20441);
nand U22439 (N_22439,N_21507,N_20751);
xor U22440 (N_22440,N_21321,N_21009);
xor U22441 (N_22441,N_21986,N_21921);
nor U22442 (N_22442,N_20028,N_21834);
xnor U22443 (N_22443,N_21108,N_20694);
nor U22444 (N_22444,N_20495,N_21178);
nand U22445 (N_22445,N_20584,N_20852);
xnor U22446 (N_22446,N_20432,N_21166);
nor U22447 (N_22447,N_20851,N_20800);
nand U22448 (N_22448,N_20638,N_20074);
xor U22449 (N_22449,N_20286,N_21016);
nor U22450 (N_22450,N_20574,N_21024);
nor U22451 (N_22451,N_20180,N_20203);
and U22452 (N_22452,N_20773,N_21482);
xnor U22453 (N_22453,N_21367,N_20200);
or U22454 (N_22454,N_21721,N_21939);
or U22455 (N_22455,N_21370,N_21563);
nand U22456 (N_22456,N_21285,N_21681);
or U22457 (N_22457,N_20537,N_20048);
and U22458 (N_22458,N_20621,N_20698);
and U22459 (N_22459,N_20596,N_20162);
and U22460 (N_22460,N_20065,N_21675);
xnor U22461 (N_22461,N_20833,N_20431);
and U22462 (N_22462,N_21035,N_21525);
and U22463 (N_22463,N_20961,N_20939);
xor U22464 (N_22464,N_21127,N_20320);
and U22465 (N_22465,N_21189,N_20144);
nor U22466 (N_22466,N_20932,N_20284);
xnor U22467 (N_22467,N_21635,N_21573);
nand U22468 (N_22468,N_20793,N_20385);
and U22469 (N_22469,N_21730,N_20950);
or U22470 (N_22470,N_21151,N_20153);
and U22471 (N_22471,N_21799,N_20127);
nand U22472 (N_22472,N_20448,N_21926);
nor U22473 (N_22473,N_21541,N_20473);
or U22474 (N_22474,N_21711,N_21273);
xnor U22475 (N_22475,N_21429,N_21176);
and U22476 (N_22476,N_21912,N_21371);
and U22477 (N_22477,N_20249,N_21806);
xor U22478 (N_22478,N_21916,N_20534);
nand U22479 (N_22479,N_20287,N_21641);
and U22480 (N_22480,N_21468,N_21893);
and U22481 (N_22481,N_20446,N_20010);
or U22482 (N_22482,N_20924,N_21954);
nand U22483 (N_22483,N_20130,N_21139);
or U22484 (N_22484,N_20113,N_21376);
xor U22485 (N_22485,N_21398,N_20543);
or U22486 (N_22486,N_20066,N_21570);
or U22487 (N_22487,N_20681,N_21998);
nand U22488 (N_22488,N_20005,N_20824);
or U22489 (N_22489,N_21729,N_20371);
nand U22490 (N_22490,N_20969,N_20600);
or U22491 (N_22491,N_20158,N_21258);
nor U22492 (N_22492,N_20513,N_20179);
xor U22493 (N_22493,N_20779,N_21308);
nor U22494 (N_22494,N_20669,N_21580);
xor U22495 (N_22495,N_21701,N_21695);
nand U22496 (N_22496,N_20359,N_21082);
or U22497 (N_22497,N_20231,N_20581);
and U22498 (N_22498,N_21428,N_21591);
and U22499 (N_22499,N_21333,N_20294);
nand U22500 (N_22500,N_21161,N_21419);
nor U22501 (N_22501,N_20548,N_20253);
or U22502 (N_22502,N_20055,N_21830);
and U22503 (N_22503,N_21853,N_21332);
or U22504 (N_22504,N_20076,N_21106);
xor U22505 (N_22505,N_21870,N_21774);
nor U22506 (N_22506,N_20084,N_20752);
nand U22507 (N_22507,N_21324,N_20654);
xnor U22508 (N_22508,N_20547,N_21029);
or U22509 (N_22509,N_21571,N_20991);
nor U22510 (N_22510,N_20019,N_21873);
nor U22511 (N_22511,N_20701,N_21717);
and U22512 (N_22512,N_21465,N_20896);
xor U22513 (N_22513,N_20971,N_21791);
nand U22514 (N_22514,N_20299,N_20755);
nor U22515 (N_22515,N_21233,N_21540);
or U22516 (N_22516,N_21975,N_20915);
nand U22517 (N_22517,N_21952,N_20102);
or U22518 (N_22518,N_20530,N_20593);
nor U22519 (N_22519,N_21361,N_21905);
xnor U22520 (N_22520,N_20148,N_20524);
nor U22521 (N_22521,N_20291,N_20465);
or U22522 (N_22522,N_21042,N_20707);
nor U22523 (N_22523,N_21243,N_21877);
or U22524 (N_22524,N_20197,N_20133);
and U22525 (N_22525,N_20805,N_20727);
and U22526 (N_22526,N_20780,N_20325);
and U22527 (N_22527,N_20447,N_21593);
xnor U22528 (N_22528,N_20204,N_20164);
or U22529 (N_22529,N_20042,N_21386);
nand U22530 (N_22530,N_21876,N_21267);
xnor U22531 (N_22531,N_21142,N_21240);
and U22532 (N_22532,N_21864,N_21995);
or U22533 (N_22533,N_21839,N_20281);
nand U22534 (N_22534,N_20658,N_21949);
and U22535 (N_22535,N_21608,N_20972);
xnor U22536 (N_22536,N_21451,N_21137);
and U22537 (N_22537,N_20020,N_21886);
or U22538 (N_22538,N_21143,N_20424);
nor U22539 (N_22539,N_20348,N_21470);
xnor U22540 (N_22540,N_20095,N_21982);
and U22541 (N_22541,N_20283,N_21808);
and U22542 (N_22542,N_21914,N_20329);
and U22543 (N_22543,N_20399,N_21217);
or U22544 (N_22544,N_21922,N_21622);
nor U22545 (N_22545,N_21076,N_20131);
nor U22546 (N_22546,N_20717,N_21478);
xor U22547 (N_22547,N_21902,N_20021);
and U22548 (N_22548,N_20661,N_21003);
and U22549 (N_22549,N_21183,N_21351);
or U22550 (N_22550,N_21989,N_20816);
nand U22551 (N_22551,N_21341,N_21530);
and U22552 (N_22552,N_20035,N_21818);
nor U22553 (N_22553,N_20586,N_20868);
xnor U22554 (N_22554,N_20089,N_21442);
xor U22555 (N_22555,N_20609,N_21743);
nand U22556 (N_22556,N_21815,N_21280);
and U22557 (N_22557,N_21087,N_20904);
nor U22558 (N_22558,N_21203,N_21418);
and U22559 (N_22559,N_20859,N_21903);
nor U22560 (N_22560,N_20567,N_20778);
xor U22561 (N_22561,N_21603,N_20216);
or U22562 (N_22562,N_21532,N_20478);
or U22563 (N_22563,N_21812,N_21682);
nor U22564 (N_22564,N_20710,N_21450);
nand U22565 (N_22565,N_20166,N_21787);
nor U22566 (N_22566,N_20252,N_20892);
and U22567 (N_22567,N_21318,N_21841);
nor U22568 (N_22568,N_20814,N_20261);
xnor U22569 (N_22569,N_20407,N_21374);
and U22570 (N_22570,N_20640,N_21245);
nor U22571 (N_22571,N_20195,N_21382);
nand U22572 (N_22572,N_21940,N_20091);
xnor U22573 (N_22573,N_21920,N_20230);
and U22574 (N_22574,N_21868,N_21232);
nand U22575 (N_22575,N_21229,N_21410);
nand U22576 (N_22576,N_20423,N_21086);
or U22577 (N_22577,N_20803,N_21547);
xnor U22578 (N_22578,N_20998,N_20011);
nor U22579 (N_22579,N_20219,N_20027);
xnor U22580 (N_22580,N_20207,N_20855);
nand U22581 (N_22581,N_21218,N_21284);
and U22582 (N_22582,N_20699,N_21550);
xor U22583 (N_22583,N_20193,N_20313);
xnor U22584 (N_22584,N_20242,N_21971);
or U22585 (N_22585,N_21569,N_21323);
nand U22586 (N_22586,N_20454,N_21664);
and U22587 (N_22587,N_21667,N_21601);
nand U22588 (N_22588,N_21770,N_20812);
or U22589 (N_22589,N_20422,N_21562);
nor U22590 (N_22590,N_20626,N_21536);
or U22591 (N_22591,N_20540,N_21855);
nand U22592 (N_22592,N_21467,N_21741);
and U22593 (N_22593,N_20783,N_20653);
nand U22594 (N_22594,N_20492,N_21436);
xor U22595 (N_22595,N_21596,N_21691);
nor U22596 (N_22596,N_20290,N_21020);
or U22597 (N_22597,N_20388,N_20604);
and U22598 (N_22598,N_21809,N_21453);
or U22599 (N_22599,N_20718,N_21501);
or U22600 (N_22600,N_21703,N_21857);
xor U22601 (N_22601,N_20268,N_21115);
nand U22602 (N_22602,N_21246,N_21472);
nand U22603 (N_22603,N_21005,N_21117);
nand U22604 (N_22604,N_21517,N_20989);
xnor U22605 (N_22605,N_21750,N_21103);
nor U22606 (N_22606,N_20012,N_21758);
and U22607 (N_22607,N_21838,N_21709);
nand U22608 (N_22608,N_21339,N_20308);
or U22609 (N_22609,N_21543,N_20215);
or U22610 (N_22610,N_20769,N_21754);
xnor U22611 (N_22611,N_20533,N_20518);
nand U22612 (N_22612,N_20981,N_20217);
nor U22613 (N_22613,N_21985,N_20819);
nor U22614 (N_22614,N_21031,N_20060);
nor U22615 (N_22615,N_20818,N_20390);
nor U22616 (N_22616,N_21314,N_20791);
and U22617 (N_22617,N_20733,N_21699);
or U22618 (N_22618,N_20768,N_21389);
nand U22619 (N_22619,N_21789,N_20182);
and U22620 (N_22620,N_21415,N_21737);
nand U22621 (N_22621,N_20737,N_20322);
nand U22622 (N_22622,N_21347,N_21411);
and U22623 (N_22623,N_20510,N_20457);
or U22624 (N_22624,N_21545,N_20266);
nor U22625 (N_22625,N_21970,N_20403);
nor U22626 (N_22626,N_20573,N_21840);
xnor U22627 (N_22627,N_21867,N_21736);
or U22628 (N_22628,N_21783,N_21967);
and U22629 (N_22629,N_21286,N_21625);
nand U22630 (N_22630,N_20154,N_20311);
nand U22631 (N_22631,N_20165,N_21350);
or U22632 (N_22632,N_20505,N_21255);
nor U22633 (N_22633,N_20629,N_21619);
xor U22634 (N_22634,N_20295,N_20603);
nor U22635 (N_22635,N_20504,N_20386);
and U22636 (N_22636,N_21782,N_21523);
xor U22637 (N_22637,N_20923,N_20415);
or U22638 (N_22638,N_21230,N_20220);
nor U22639 (N_22639,N_21526,N_20891);
or U22640 (N_22640,N_20679,N_21210);
xor U22641 (N_22641,N_21330,N_20580);
and U22642 (N_22642,N_21424,N_20265);
or U22643 (N_22643,N_20079,N_20107);
nor U22644 (N_22644,N_20440,N_20758);
xnor U22645 (N_22645,N_20023,N_21097);
or U22646 (N_22646,N_20232,N_21440);
and U22647 (N_22647,N_21829,N_20659);
xor U22648 (N_22648,N_20817,N_20059);
xor U22649 (N_22649,N_20974,N_21089);
xor U22650 (N_22650,N_20214,N_21432);
or U22651 (N_22651,N_21316,N_21421);
nand U22652 (N_22652,N_20870,N_20966);
nand U22653 (N_22653,N_20700,N_21173);
nor U22654 (N_22654,N_20270,N_21836);
nand U22655 (N_22655,N_21977,N_20528);
nand U22656 (N_22656,N_20722,N_21315);
xnor U22657 (N_22657,N_21373,N_20922);
nand U22658 (N_22658,N_20038,N_20559);
and U22659 (N_22659,N_21645,N_20843);
xor U22660 (N_22660,N_20189,N_20122);
nand U22661 (N_22661,N_21017,N_21595);
nand U22662 (N_22662,N_20094,N_21168);
xnor U22663 (N_22663,N_20014,N_20365);
xor U22664 (N_22664,N_20435,N_20418);
nand U22665 (N_22665,N_20636,N_20651);
xor U22666 (N_22666,N_20553,N_20260);
and U22667 (N_22667,N_21941,N_20334);
and U22668 (N_22668,N_21207,N_20716);
nor U22669 (N_22669,N_21403,N_21726);
nor U22670 (N_22670,N_21685,N_20353);
nand U22671 (N_22671,N_21083,N_20347);
xnor U22672 (N_22672,N_21177,N_21817);
nor U22673 (N_22673,N_20606,N_20862);
and U22674 (N_22674,N_21360,N_20620);
or U22675 (N_22675,N_20994,N_21651);
nor U22676 (N_22676,N_21080,N_20421);
or U22677 (N_22677,N_20497,N_20331);
xnor U22678 (N_22678,N_20117,N_21602);
nand U22679 (N_22679,N_20686,N_20811);
and U22680 (N_22680,N_21486,N_20337);
nand U22681 (N_22681,N_21518,N_21669);
or U22682 (N_22682,N_21182,N_20556);
nand U22683 (N_22683,N_21354,N_20226);
xor U22684 (N_22684,N_21223,N_21226);
nor U22685 (N_22685,N_21508,N_21513);
nand U22686 (N_22686,N_21930,N_20973);
and U22687 (N_22687,N_21597,N_21662);
nand U22688 (N_22688,N_20903,N_20880);
nor U22689 (N_22689,N_20273,N_21529);
and U22690 (N_22690,N_21426,N_20764);
and U22691 (N_22691,N_21460,N_21079);
nor U22692 (N_22692,N_20639,N_21288);
and U22693 (N_22693,N_21399,N_21628);
nor U22694 (N_22694,N_20890,N_20350);
nand U22695 (N_22695,N_21960,N_20628);
or U22696 (N_22696,N_21033,N_20156);
nand U22697 (N_22697,N_21402,N_20978);
or U22698 (N_22698,N_20602,N_20858);
or U22699 (N_22699,N_21761,N_21422);
nand U22700 (N_22700,N_21238,N_21654);
nand U22701 (N_22701,N_21568,N_21524);
or U22702 (N_22702,N_20747,N_21072);
nor U22703 (N_22703,N_20137,N_20502);
nand U22704 (N_22704,N_21126,N_20072);
nor U22705 (N_22705,N_21732,N_20272);
xnor U22706 (N_22706,N_21656,N_20071);
and U22707 (N_22707,N_21763,N_20187);
and U22708 (N_22708,N_20551,N_21032);
nand U22709 (N_22709,N_21261,N_21991);
or U22710 (N_22710,N_20372,N_20333);
xor U22711 (N_22711,N_20192,N_20168);
and U22712 (N_22712,N_20086,N_21923);
xor U22713 (N_22713,N_21552,N_20617);
xnor U22714 (N_22714,N_21012,N_20250);
nor U22715 (N_22715,N_21704,N_20227);
and U22716 (N_22716,N_20936,N_20143);
nor U22717 (N_22717,N_20577,N_20970);
nor U22718 (N_22718,N_21344,N_20209);
nand U22719 (N_22719,N_20341,N_21790);
xnor U22720 (N_22720,N_21966,N_20542);
nand U22721 (N_22721,N_21056,N_20866);
nand U22722 (N_22722,N_21577,N_20212);
nor U22723 (N_22723,N_20169,N_21136);
nand U22724 (N_22724,N_20199,N_21898);
nand U22725 (N_22725,N_21102,N_20919);
and U22726 (N_22726,N_20336,N_20921);
xnor U22727 (N_22727,N_20030,N_21066);
or U22728 (N_22728,N_20671,N_21816);
and U22729 (N_22729,N_20149,N_21565);
or U22730 (N_22730,N_20785,N_20736);
and U22731 (N_22731,N_21781,N_21510);
nand U22732 (N_22732,N_21807,N_20802);
nand U22733 (N_22733,N_21696,N_21932);
or U22734 (N_22734,N_21715,N_21375);
and U22735 (N_22735,N_20043,N_20456);
nor U22736 (N_22736,N_20879,N_20032);
xor U22737 (N_22737,N_21827,N_21441);
and U22738 (N_22738,N_20312,N_21104);
nor U22739 (N_22739,N_21416,N_21910);
xnor U22740 (N_22740,N_20225,N_21880);
or U22741 (N_22741,N_20960,N_20763);
xor U22742 (N_22742,N_20933,N_21672);
and U22743 (N_22743,N_21924,N_21015);
nor U22744 (N_22744,N_20310,N_20863);
nand U22745 (N_22745,N_20049,N_20682);
and U22746 (N_22746,N_21271,N_20067);
and U22747 (N_22747,N_21747,N_20288);
and U22748 (N_22748,N_21026,N_20318);
nand U22749 (N_22749,N_20306,N_20853);
nor U22750 (N_22750,N_20040,N_21352);
nor U22751 (N_22751,N_21322,N_21247);
nor U22752 (N_22752,N_21458,N_20488);
nand U22753 (N_22753,N_21388,N_20259);
nand U22754 (N_22754,N_21135,N_20744);
or U22755 (N_22755,N_21148,N_20539);
xnor U22756 (N_22756,N_21727,N_21291);
nand U22757 (N_22757,N_21455,N_21825);
or U22758 (N_22758,N_20914,N_21420);
and U22759 (N_22759,N_20121,N_20009);
nor U22760 (N_22760,N_20815,N_21885);
xnor U22761 (N_22761,N_20983,N_21326);
nand U22762 (N_22762,N_21538,N_20693);
nor U22763 (N_22763,N_20412,N_20235);
nor U22764 (N_22764,N_20525,N_21381);
nand U22765 (N_22765,N_21107,N_21036);
or U22766 (N_22766,N_21112,N_20508);
nand U22767 (N_22767,N_20463,N_21652);
nand U22768 (N_22768,N_21004,N_21406);
or U22769 (N_22769,N_21073,N_21133);
and U22770 (N_22770,N_20975,N_21850);
and U22771 (N_22771,N_20938,N_21588);
and U22772 (N_22772,N_20514,N_20208);
nand U22773 (N_22773,N_20691,N_20069);
xnor U22774 (N_22774,N_21045,N_20569);
xor U22775 (N_22775,N_20486,N_20988);
nand U22776 (N_22776,N_20646,N_20111);
and U22777 (N_22777,N_21702,N_20899);
nor U22778 (N_22778,N_20004,N_21644);
or U22779 (N_22779,N_21463,N_20100);
xor U22780 (N_22780,N_21520,N_20443);
and U22781 (N_22781,N_20398,N_20827);
and U22782 (N_22782,N_21292,N_20458);
and U22783 (N_22783,N_20762,N_21060);
or U22784 (N_22784,N_21983,N_20792);
nand U22785 (N_22785,N_20695,N_21968);
nor U22786 (N_22786,N_20958,N_20031);
xnor U22787 (N_22787,N_20202,N_20174);
nor U22788 (N_22788,N_20719,N_21272);
nor U22789 (N_22789,N_20608,N_20723);
xnor U22790 (N_22790,N_20529,N_20309);
and U22791 (N_22791,N_20976,N_21646);
and U22792 (N_22792,N_21780,N_21771);
nor U22793 (N_22793,N_21319,N_20046);
and U22794 (N_22794,N_21081,N_21683);
nand U22795 (N_22795,N_21377,N_21446);
nand U22796 (N_22796,N_21295,N_20947);
and U22797 (N_22797,N_21378,N_20516);
xnor U22798 (N_22798,N_20277,N_21712);
or U22799 (N_22799,N_21124,N_20845);
nand U22800 (N_22800,N_21874,N_20383);
nor U22801 (N_22801,N_20480,N_21228);
nor U22802 (N_22802,N_21765,N_20576);
nand U22803 (N_22803,N_21785,N_20663);
and U22804 (N_22804,N_21348,N_20420);
nand U22805 (N_22805,N_20869,N_20358);
nand U22806 (N_22806,N_21665,N_20064);
nor U22807 (N_22807,N_20044,N_21407);
nor U22808 (N_22808,N_21392,N_20183);
nand U22809 (N_22809,N_20623,N_20943);
and U22810 (N_22810,N_20585,N_20007);
nor U22811 (N_22811,N_21784,N_21490);
or U22812 (N_22812,N_20449,N_21313);
xnor U22813 (N_22813,N_20413,N_20917);
nand U22814 (N_22814,N_21847,N_20771);
or U22815 (N_22815,N_20781,N_20746);
xnor U22816 (N_22816,N_21716,N_21897);
and U22817 (N_22817,N_21512,N_20263);
xor U22818 (N_22818,N_21101,N_21663);
xnor U22819 (N_22819,N_20907,N_21884);
and U22820 (N_22820,N_20247,N_20804);
nand U22821 (N_22821,N_21934,N_20218);
nor U22822 (N_22822,N_20753,N_20159);
nand U22823 (N_22823,N_21396,N_21464);
nor U22824 (N_22824,N_21466,N_20039);
nor U22825 (N_22825,N_21265,N_21556);
and U22826 (N_22826,N_21706,N_21917);
xor U22827 (N_22827,N_21674,N_21879);
and U22828 (N_22828,N_20839,N_20062);
nor U22829 (N_22829,N_20224,N_21708);
and U22830 (N_22830,N_21759,N_21251);
or U22831 (N_22831,N_21234,N_21212);
and U22832 (N_22832,N_20916,N_21053);
xor U22833 (N_22833,N_21896,N_20912);
nor U22834 (N_22834,N_20595,N_20927);
or U22835 (N_22835,N_20865,N_20643);
nor U22836 (N_22836,N_21504,N_20205);
and U22837 (N_22837,N_20985,N_21476);
or U22838 (N_22838,N_20996,N_21835);
and U22839 (N_22839,N_20840,N_21776);
xnor U22840 (N_22840,N_20656,N_21194);
or U22841 (N_22841,N_21630,N_21305);
nor U22842 (N_22842,N_21206,N_21710);
nor U22843 (N_22843,N_20416,N_20895);
and U22844 (N_22844,N_20196,N_20750);
or U22845 (N_22845,N_21018,N_21456);
xor U22846 (N_22846,N_20786,N_21734);
xnor U22847 (N_22847,N_20097,N_21063);
and U22848 (N_22848,N_20790,N_20796);
nor U22849 (N_22849,N_20749,N_21346);
and U22850 (N_22850,N_20627,N_20452);
nand U22851 (N_22851,N_20116,N_20706);
and U22852 (N_22852,N_21167,N_20831);
and U22853 (N_22853,N_21676,N_21583);
nand U22854 (N_22854,N_20105,N_20690);
xor U22855 (N_22855,N_20599,N_21159);
or U22856 (N_22856,N_21409,N_21609);
or U22857 (N_22857,N_20935,N_21116);
nor U22858 (N_22858,N_21942,N_21493);
nor U22859 (N_22859,N_20942,N_20565);
and U22860 (N_22860,N_20631,N_21659);
or U22861 (N_22861,N_21528,N_20471);
and U22862 (N_22862,N_21613,N_21196);
xnor U22863 (N_22863,N_21900,N_21649);
nor U22864 (N_22864,N_21236,N_21639);
nor U22865 (N_22865,N_21792,N_20104);
nand U22866 (N_22866,N_21358,N_20704);
or U22867 (N_22867,N_20594,N_20873);
nor U22868 (N_22868,N_20339,N_21484);
or U22869 (N_22869,N_20239,N_20015);
xnor U22870 (N_22870,N_20276,N_21793);
or U22871 (N_22871,N_21320,N_20171);
or U22872 (N_22872,N_20549,N_20787);
nor U22873 (N_22873,N_21987,N_21186);
nand U22874 (N_22874,N_21474,N_20526);
nand U22875 (N_22875,N_20697,N_21620);
and U22876 (N_22876,N_21430,N_20190);
and U22877 (N_22877,N_21755,N_20340);
and U22878 (N_22878,N_20129,N_20001);
xor U22879 (N_22879,N_21999,N_21564);
nand U22880 (N_22880,N_21193,N_21680);
nand U22881 (N_22881,N_21002,N_21190);
nand U22882 (N_22882,N_21944,N_20161);
nand U22883 (N_22883,N_20560,N_21745);
and U22884 (N_22884,N_20828,N_20878);
nand U22885 (N_22885,N_20409,N_20941);
or U22886 (N_22886,N_20229,N_20807);
nor U22887 (N_22887,N_20464,N_21951);
or U22888 (N_22888,N_20847,N_20822);
nor U22889 (N_22889,N_20354,N_20597);
nand U22890 (N_22890,N_20417,N_20103);
and U22891 (N_22891,N_20931,N_20501);
or U22892 (N_22892,N_20906,N_20368);
nand U22893 (N_22893,N_21861,N_21990);
or U22894 (N_22894,N_20986,N_20545);
nand U22895 (N_22895,N_20496,N_21756);
and U22896 (N_22896,N_21379,N_21293);
and U22897 (N_22897,N_20163,N_21034);
or U22898 (N_22898,N_20531,N_21943);
nor U22899 (N_22899,N_20054,N_21623);
nor U22900 (N_22900,N_21849,N_21611);
or U22901 (N_22901,N_20500,N_21572);
nor U22902 (N_22902,N_20234,N_20201);
or U22903 (N_22903,N_21632,N_21888);
or U22904 (N_22904,N_20894,N_21895);
xnor U22905 (N_22905,N_21355,N_20278);
and U22906 (N_22906,N_21393,N_20170);
xor U22907 (N_22907,N_21075,N_21276);
and U22908 (N_22908,N_20367,N_20742);
or U22909 (N_22909,N_20090,N_21533);
xor U22910 (N_22910,N_20439,N_21181);
and U22911 (N_22911,N_21279,N_20132);
nand U22912 (N_22912,N_20611,N_21688);
or U22913 (N_22913,N_20836,N_21150);
or U22914 (N_22914,N_20642,N_21412);
and U22915 (N_22915,N_20374,N_21527);
and U22916 (N_22916,N_20245,N_21869);
xor U22917 (N_22917,N_21634,N_21391);
nand U22918 (N_22918,N_21443,N_20949);
nand U22919 (N_22919,N_20760,N_20491);
xor U22920 (N_22920,N_20466,N_21302);
nor U22921 (N_22921,N_20666,N_20013);
nor U22922 (N_22922,N_20321,N_21250);
xnor U22923 (N_22923,N_21901,N_21345);
and U22924 (N_22924,N_20641,N_20674);
or U22925 (N_22925,N_21074,N_20612);
nor U22926 (N_22926,N_20108,N_20735);
xor U22927 (N_22927,N_21071,N_20715);
nor U22928 (N_22928,N_20098,N_21933);
nor U22929 (N_22929,N_20841,N_21582);
nand U22930 (N_22930,N_20120,N_21802);
nand U22931 (N_22931,N_20114,N_21192);
xor U22932 (N_22932,N_20995,N_20136);
nor U22933 (N_22933,N_20410,N_20123);
and U22934 (N_22934,N_20948,N_21423);
nor U22935 (N_22935,N_21826,N_21187);
or U22936 (N_22936,N_21866,N_20759);
xor U22937 (N_22937,N_21306,N_20854);
xnor U22938 (N_22938,N_21548,N_20678);
nor U22939 (N_22939,N_20262,N_21610);
or U22940 (N_22940,N_21248,N_20255);
and U22941 (N_22941,N_21188,N_20765);
xor U22942 (N_22942,N_21661,N_21336);
xor U22943 (N_22943,N_21854,N_21297);
or U22944 (N_22944,N_20343,N_20928);
nand U22945 (N_22945,N_20428,N_20849);
or U22946 (N_22946,N_20848,N_21589);
xnor U22947 (N_22947,N_20776,N_20282);
xor U22948 (N_22948,N_20206,N_21353);
and U22949 (N_22949,N_21277,N_20237);
and U22950 (N_22950,N_20088,N_21929);
nor U22951 (N_22951,N_20017,N_21000);
and U22952 (N_22952,N_20335,N_20467);
or U22953 (N_22953,N_20872,N_20820);
nand U22954 (N_22954,N_20198,N_20990);
nand U22955 (N_22955,N_20861,N_21254);
and U22956 (N_22956,N_21585,N_21028);
or U22957 (N_22957,N_20789,N_20589);
and U22958 (N_22958,N_21557,N_21448);
xnor U22959 (N_22959,N_20926,N_20523);
nand U22960 (N_22960,N_21899,N_21049);
nor U22961 (N_22961,N_21425,N_20176);
or U22962 (N_22962,N_21155,N_20601);
nand U22963 (N_22963,N_20550,N_21766);
nor U22964 (N_22964,N_21764,N_21728);
nor U22965 (N_22965,N_21496,N_20575);
xor U22966 (N_22966,N_21612,N_20244);
and U22967 (N_22967,N_20850,N_20992);
and U22968 (N_22968,N_20022,N_20954);
nand U22969 (N_22969,N_20509,N_21163);
xor U22970 (N_22970,N_20582,N_20357);
and U22971 (N_22971,N_20474,N_20999);
xor U22972 (N_22972,N_21477,N_20404);
xor U22973 (N_22973,N_20630,N_21537);
nand U22974 (N_22974,N_21340,N_20489);
xor U22975 (N_22975,N_21519,N_21778);
nand U22976 (N_22976,N_20445,N_20444);
and U22977 (N_22977,N_20292,N_21976);
or U22978 (N_22978,N_21365,N_21554);
and U22979 (N_22979,N_21390,N_20766);
and U22980 (N_22980,N_21235,N_20967);
or U22981 (N_22981,N_21863,N_20328);
nand U22982 (N_22982,N_20538,N_21294);
nand U22983 (N_22983,N_21211,N_20821);
nor U22984 (N_22984,N_20316,N_21598);
xor U22985 (N_22985,N_21249,N_20487);
and U22986 (N_22986,N_21221,N_21222);
or U22987 (N_22987,N_21845,N_21616);
and U22988 (N_22988,N_21660,N_21891);
xnor U22989 (N_22989,N_21057,N_20000);
xor U22990 (N_22990,N_21500,N_21121);
nor U22991 (N_22991,N_21195,N_20788);
xor U22992 (N_22992,N_21666,N_20588);
nor U22993 (N_22993,N_21037,N_21008);
and U22994 (N_22994,N_21677,N_20826);
nand U22995 (N_22995,N_21749,N_20243);
nor U22996 (N_22996,N_20124,N_20676);
nand U22997 (N_22997,N_21043,N_21414);
nand U22998 (N_22998,N_21724,N_21575);
nand U22999 (N_22999,N_20063,N_21475);
nor U23000 (N_23000,N_20817,N_21608);
nor U23001 (N_23001,N_21885,N_20465);
nor U23002 (N_23002,N_21924,N_21994);
xnor U23003 (N_23003,N_20034,N_20400);
nand U23004 (N_23004,N_20115,N_21220);
xnor U23005 (N_23005,N_21549,N_21215);
xor U23006 (N_23006,N_20233,N_21219);
nor U23007 (N_23007,N_20511,N_20429);
nand U23008 (N_23008,N_20479,N_20862);
or U23009 (N_23009,N_20395,N_21882);
or U23010 (N_23010,N_21939,N_21370);
xnor U23011 (N_23011,N_20180,N_21782);
nor U23012 (N_23012,N_21244,N_21379);
nand U23013 (N_23013,N_21464,N_20317);
xor U23014 (N_23014,N_20264,N_21482);
xor U23015 (N_23015,N_20962,N_21124);
or U23016 (N_23016,N_21553,N_20404);
nor U23017 (N_23017,N_20169,N_21646);
xnor U23018 (N_23018,N_20603,N_20742);
or U23019 (N_23019,N_21718,N_21567);
xnor U23020 (N_23020,N_21806,N_21168);
nor U23021 (N_23021,N_20463,N_21211);
nor U23022 (N_23022,N_21165,N_21071);
or U23023 (N_23023,N_20323,N_20724);
or U23024 (N_23024,N_21709,N_21161);
nand U23025 (N_23025,N_21232,N_21443);
nor U23026 (N_23026,N_21916,N_21042);
nand U23027 (N_23027,N_21690,N_20913);
nor U23028 (N_23028,N_21806,N_21914);
or U23029 (N_23029,N_21445,N_21054);
xnor U23030 (N_23030,N_20669,N_20235);
xnor U23031 (N_23031,N_20505,N_21167);
nor U23032 (N_23032,N_21481,N_20525);
nand U23033 (N_23033,N_20605,N_20152);
or U23034 (N_23034,N_21286,N_21911);
xnor U23035 (N_23035,N_21515,N_21037);
and U23036 (N_23036,N_20990,N_20203);
nand U23037 (N_23037,N_21571,N_20257);
xnor U23038 (N_23038,N_20424,N_20699);
nor U23039 (N_23039,N_21598,N_21037);
and U23040 (N_23040,N_21747,N_20489);
and U23041 (N_23041,N_20732,N_20350);
or U23042 (N_23042,N_21706,N_20768);
and U23043 (N_23043,N_20484,N_21436);
nor U23044 (N_23044,N_21158,N_21919);
and U23045 (N_23045,N_21413,N_21813);
nor U23046 (N_23046,N_21718,N_20816);
and U23047 (N_23047,N_21043,N_21765);
xnor U23048 (N_23048,N_21546,N_20732);
nand U23049 (N_23049,N_20234,N_21584);
or U23050 (N_23050,N_21281,N_20810);
and U23051 (N_23051,N_21687,N_20568);
nor U23052 (N_23052,N_20954,N_21909);
and U23053 (N_23053,N_21871,N_20563);
nor U23054 (N_23054,N_20822,N_20960);
nand U23055 (N_23055,N_20144,N_21509);
nand U23056 (N_23056,N_20489,N_20285);
nand U23057 (N_23057,N_20260,N_20370);
nand U23058 (N_23058,N_21219,N_21048);
xor U23059 (N_23059,N_21916,N_21896);
nor U23060 (N_23060,N_21853,N_21899);
nor U23061 (N_23061,N_21411,N_21219);
and U23062 (N_23062,N_20740,N_21156);
or U23063 (N_23063,N_21880,N_21657);
and U23064 (N_23064,N_20505,N_21992);
nor U23065 (N_23065,N_20006,N_20195);
or U23066 (N_23066,N_20110,N_20473);
and U23067 (N_23067,N_21899,N_20799);
xor U23068 (N_23068,N_21230,N_20744);
xor U23069 (N_23069,N_21762,N_21557);
or U23070 (N_23070,N_21388,N_21329);
nor U23071 (N_23071,N_20546,N_21958);
nor U23072 (N_23072,N_21659,N_20540);
and U23073 (N_23073,N_20625,N_21894);
nand U23074 (N_23074,N_20648,N_20987);
or U23075 (N_23075,N_21436,N_21267);
nand U23076 (N_23076,N_20017,N_21489);
or U23077 (N_23077,N_21481,N_20238);
or U23078 (N_23078,N_21195,N_21527);
or U23079 (N_23079,N_21188,N_21120);
nor U23080 (N_23080,N_21688,N_20277);
xor U23081 (N_23081,N_20084,N_20138);
and U23082 (N_23082,N_21403,N_20204);
or U23083 (N_23083,N_20834,N_20639);
nand U23084 (N_23084,N_20181,N_20275);
xor U23085 (N_23085,N_21258,N_20966);
nor U23086 (N_23086,N_20904,N_21674);
or U23087 (N_23087,N_21119,N_21320);
nor U23088 (N_23088,N_21504,N_20972);
nor U23089 (N_23089,N_21111,N_20615);
or U23090 (N_23090,N_20205,N_21961);
and U23091 (N_23091,N_21613,N_21113);
xor U23092 (N_23092,N_21337,N_20487);
or U23093 (N_23093,N_20326,N_21567);
nor U23094 (N_23094,N_21505,N_21179);
xnor U23095 (N_23095,N_21723,N_20455);
and U23096 (N_23096,N_20065,N_21445);
nand U23097 (N_23097,N_20904,N_20504);
nand U23098 (N_23098,N_21804,N_21647);
and U23099 (N_23099,N_20249,N_20350);
and U23100 (N_23100,N_21699,N_21594);
xnor U23101 (N_23101,N_21716,N_21762);
xnor U23102 (N_23102,N_21597,N_20582);
xnor U23103 (N_23103,N_21441,N_20774);
or U23104 (N_23104,N_20555,N_20471);
and U23105 (N_23105,N_21733,N_20676);
xnor U23106 (N_23106,N_20942,N_20301);
xnor U23107 (N_23107,N_21985,N_20739);
nand U23108 (N_23108,N_21007,N_20194);
nor U23109 (N_23109,N_20659,N_21220);
xnor U23110 (N_23110,N_21341,N_21151);
nor U23111 (N_23111,N_20802,N_20884);
nor U23112 (N_23112,N_21158,N_20047);
nor U23113 (N_23113,N_21694,N_20055);
and U23114 (N_23114,N_20482,N_21798);
and U23115 (N_23115,N_21576,N_21245);
xnor U23116 (N_23116,N_21639,N_20114);
xor U23117 (N_23117,N_21481,N_20721);
nor U23118 (N_23118,N_20982,N_20458);
or U23119 (N_23119,N_21117,N_20223);
nand U23120 (N_23120,N_21407,N_21225);
nor U23121 (N_23121,N_21521,N_21340);
and U23122 (N_23122,N_21791,N_20477);
or U23123 (N_23123,N_21264,N_20331);
or U23124 (N_23124,N_20835,N_21884);
and U23125 (N_23125,N_21932,N_20448);
xnor U23126 (N_23126,N_20932,N_21383);
and U23127 (N_23127,N_21663,N_21374);
or U23128 (N_23128,N_20136,N_20425);
and U23129 (N_23129,N_21789,N_21116);
nor U23130 (N_23130,N_21655,N_20636);
nand U23131 (N_23131,N_21491,N_20078);
nor U23132 (N_23132,N_21657,N_21585);
and U23133 (N_23133,N_21742,N_20794);
nor U23134 (N_23134,N_21726,N_21350);
xnor U23135 (N_23135,N_20217,N_21803);
nor U23136 (N_23136,N_21140,N_21850);
nor U23137 (N_23137,N_21057,N_20843);
xor U23138 (N_23138,N_21725,N_20129);
or U23139 (N_23139,N_20188,N_20808);
and U23140 (N_23140,N_20778,N_21444);
and U23141 (N_23141,N_20070,N_21061);
or U23142 (N_23142,N_20930,N_20110);
and U23143 (N_23143,N_20039,N_21124);
nand U23144 (N_23144,N_21998,N_21800);
nor U23145 (N_23145,N_20012,N_21964);
nand U23146 (N_23146,N_20813,N_21877);
xor U23147 (N_23147,N_20182,N_21035);
nor U23148 (N_23148,N_20483,N_20413);
or U23149 (N_23149,N_20045,N_20839);
xor U23150 (N_23150,N_21043,N_20896);
and U23151 (N_23151,N_20291,N_20235);
or U23152 (N_23152,N_20847,N_20533);
xnor U23153 (N_23153,N_21941,N_20281);
and U23154 (N_23154,N_21694,N_21293);
nand U23155 (N_23155,N_21850,N_20260);
nand U23156 (N_23156,N_21114,N_21208);
nand U23157 (N_23157,N_21256,N_20843);
nand U23158 (N_23158,N_20809,N_20338);
xor U23159 (N_23159,N_21941,N_20500);
nand U23160 (N_23160,N_21163,N_21725);
and U23161 (N_23161,N_20917,N_21395);
and U23162 (N_23162,N_21905,N_21612);
nand U23163 (N_23163,N_21530,N_21627);
or U23164 (N_23164,N_21108,N_21023);
nand U23165 (N_23165,N_20484,N_20794);
or U23166 (N_23166,N_21187,N_21110);
nand U23167 (N_23167,N_20616,N_21347);
or U23168 (N_23168,N_21523,N_20125);
xnor U23169 (N_23169,N_20231,N_20852);
and U23170 (N_23170,N_21857,N_20751);
or U23171 (N_23171,N_21285,N_20274);
nor U23172 (N_23172,N_20719,N_20012);
or U23173 (N_23173,N_21819,N_21557);
and U23174 (N_23174,N_20047,N_20211);
xor U23175 (N_23175,N_21988,N_21736);
or U23176 (N_23176,N_20926,N_20425);
xnor U23177 (N_23177,N_20574,N_21041);
nor U23178 (N_23178,N_20289,N_20279);
xnor U23179 (N_23179,N_20483,N_20247);
nor U23180 (N_23180,N_21316,N_21482);
or U23181 (N_23181,N_20656,N_21691);
and U23182 (N_23182,N_20602,N_21721);
and U23183 (N_23183,N_20936,N_20718);
and U23184 (N_23184,N_21107,N_20755);
nor U23185 (N_23185,N_21895,N_20926);
xnor U23186 (N_23186,N_20317,N_21589);
nand U23187 (N_23187,N_20441,N_21059);
nor U23188 (N_23188,N_21320,N_21071);
nand U23189 (N_23189,N_21986,N_21974);
and U23190 (N_23190,N_20436,N_20243);
xnor U23191 (N_23191,N_21055,N_21100);
and U23192 (N_23192,N_20228,N_21820);
nor U23193 (N_23193,N_21351,N_21378);
or U23194 (N_23194,N_20732,N_20173);
nand U23195 (N_23195,N_20210,N_21562);
xnor U23196 (N_23196,N_21150,N_21237);
nor U23197 (N_23197,N_20036,N_21943);
xnor U23198 (N_23198,N_20083,N_20116);
nor U23199 (N_23199,N_21115,N_20361);
xor U23200 (N_23200,N_20036,N_20989);
nand U23201 (N_23201,N_21682,N_21145);
and U23202 (N_23202,N_20825,N_21581);
nor U23203 (N_23203,N_20405,N_20229);
and U23204 (N_23204,N_20678,N_20096);
or U23205 (N_23205,N_20743,N_21779);
nand U23206 (N_23206,N_21894,N_21995);
or U23207 (N_23207,N_21357,N_21868);
nand U23208 (N_23208,N_21788,N_20055);
xor U23209 (N_23209,N_21749,N_21394);
nand U23210 (N_23210,N_20974,N_21320);
xnor U23211 (N_23211,N_20282,N_21536);
nor U23212 (N_23212,N_20913,N_20120);
xnor U23213 (N_23213,N_21740,N_20295);
or U23214 (N_23214,N_20923,N_21754);
nand U23215 (N_23215,N_21784,N_20985);
xnor U23216 (N_23216,N_21992,N_20684);
xor U23217 (N_23217,N_20219,N_21647);
nand U23218 (N_23218,N_21223,N_21337);
nand U23219 (N_23219,N_20769,N_21118);
nand U23220 (N_23220,N_21525,N_20351);
or U23221 (N_23221,N_21210,N_20722);
xor U23222 (N_23222,N_21206,N_21681);
xor U23223 (N_23223,N_20292,N_20664);
xor U23224 (N_23224,N_20026,N_21303);
and U23225 (N_23225,N_20163,N_21373);
nand U23226 (N_23226,N_21787,N_20635);
nand U23227 (N_23227,N_20414,N_21240);
nor U23228 (N_23228,N_20918,N_20756);
nand U23229 (N_23229,N_20330,N_21586);
nand U23230 (N_23230,N_20135,N_20880);
and U23231 (N_23231,N_21037,N_21636);
nand U23232 (N_23232,N_20597,N_21087);
xor U23233 (N_23233,N_21149,N_20925);
xnor U23234 (N_23234,N_20484,N_21850);
xnor U23235 (N_23235,N_21616,N_21354);
nand U23236 (N_23236,N_21230,N_20920);
xnor U23237 (N_23237,N_20385,N_21285);
xnor U23238 (N_23238,N_21799,N_20208);
and U23239 (N_23239,N_21009,N_20256);
nor U23240 (N_23240,N_21853,N_20925);
nor U23241 (N_23241,N_20363,N_20616);
nor U23242 (N_23242,N_21409,N_21867);
and U23243 (N_23243,N_21543,N_21459);
or U23244 (N_23244,N_20316,N_21982);
xor U23245 (N_23245,N_21468,N_20791);
and U23246 (N_23246,N_20144,N_20661);
xor U23247 (N_23247,N_20866,N_20381);
xnor U23248 (N_23248,N_20360,N_21009);
and U23249 (N_23249,N_21466,N_20086);
nor U23250 (N_23250,N_21355,N_20808);
xnor U23251 (N_23251,N_21374,N_21969);
xnor U23252 (N_23252,N_20461,N_21330);
nand U23253 (N_23253,N_21230,N_20371);
or U23254 (N_23254,N_20358,N_20093);
and U23255 (N_23255,N_20332,N_21104);
or U23256 (N_23256,N_20576,N_20414);
nor U23257 (N_23257,N_21836,N_21692);
nor U23258 (N_23258,N_21563,N_21873);
nand U23259 (N_23259,N_21614,N_20623);
xnor U23260 (N_23260,N_20730,N_20821);
and U23261 (N_23261,N_20584,N_21464);
and U23262 (N_23262,N_20225,N_21046);
and U23263 (N_23263,N_20054,N_20978);
or U23264 (N_23264,N_21614,N_20604);
nor U23265 (N_23265,N_21373,N_21010);
nor U23266 (N_23266,N_21049,N_20588);
or U23267 (N_23267,N_21749,N_21330);
or U23268 (N_23268,N_21861,N_20358);
nor U23269 (N_23269,N_20316,N_20626);
nor U23270 (N_23270,N_21741,N_21992);
nand U23271 (N_23271,N_21632,N_20151);
and U23272 (N_23272,N_20374,N_20410);
xnor U23273 (N_23273,N_20168,N_21562);
xor U23274 (N_23274,N_20556,N_20172);
and U23275 (N_23275,N_21349,N_21305);
xnor U23276 (N_23276,N_21312,N_20390);
nand U23277 (N_23277,N_20647,N_21207);
xnor U23278 (N_23278,N_21477,N_20519);
nor U23279 (N_23279,N_20722,N_21005);
nor U23280 (N_23280,N_20919,N_20159);
xnor U23281 (N_23281,N_21157,N_20869);
and U23282 (N_23282,N_21948,N_20280);
nor U23283 (N_23283,N_21221,N_21245);
nor U23284 (N_23284,N_20809,N_20423);
or U23285 (N_23285,N_21201,N_21956);
and U23286 (N_23286,N_21210,N_21989);
and U23287 (N_23287,N_20485,N_20133);
xor U23288 (N_23288,N_20816,N_20251);
or U23289 (N_23289,N_21513,N_20450);
xor U23290 (N_23290,N_21429,N_20607);
nand U23291 (N_23291,N_21616,N_21941);
nand U23292 (N_23292,N_21350,N_20883);
nor U23293 (N_23293,N_20912,N_20627);
and U23294 (N_23294,N_21304,N_21715);
xor U23295 (N_23295,N_20468,N_20976);
xor U23296 (N_23296,N_20078,N_21573);
nand U23297 (N_23297,N_20107,N_21978);
nand U23298 (N_23298,N_20876,N_21174);
xor U23299 (N_23299,N_20780,N_20307);
xor U23300 (N_23300,N_21908,N_21950);
nor U23301 (N_23301,N_21064,N_21306);
and U23302 (N_23302,N_21529,N_20308);
or U23303 (N_23303,N_21358,N_20651);
xor U23304 (N_23304,N_20261,N_21241);
xor U23305 (N_23305,N_21285,N_20365);
and U23306 (N_23306,N_20755,N_20318);
or U23307 (N_23307,N_21155,N_21960);
xor U23308 (N_23308,N_21401,N_20961);
nor U23309 (N_23309,N_21550,N_21195);
xor U23310 (N_23310,N_20726,N_21512);
xnor U23311 (N_23311,N_20216,N_21125);
or U23312 (N_23312,N_21566,N_21684);
nor U23313 (N_23313,N_20259,N_20191);
nor U23314 (N_23314,N_20877,N_20495);
xor U23315 (N_23315,N_21132,N_21040);
and U23316 (N_23316,N_21522,N_21888);
or U23317 (N_23317,N_20256,N_21986);
nand U23318 (N_23318,N_21510,N_20027);
or U23319 (N_23319,N_21542,N_20961);
nor U23320 (N_23320,N_21797,N_20669);
nand U23321 (N_23321,N_21457,N_20752);
xnor U23322 (N_23322,N_21836,N_21007);
or U23323 (N_23323,N_20828,N_21312);
nand U23324 (N_23324,N_21685,N_20769);
nor U23325 (N_23325,N_20420,N_20773);
xnor U23326 (N_23326,N_20434,N_21977);
nor U23327 (N_23327,N_20408,N_20902);
xor U23328 (N_23328,N_20697,N_21224);
xor U23329 (N_23329,N_21566,N_20454);
and U23330 (N_23330,N_21097,N_20959);
xor U23331 (N_23331,N_20556,N_20755);
or U23332 (N_23332,N_20871,N_21640);
nor U23333 (N_23333,N_20098,N_20721);
and U23334 (N_23334,N_21852,N_21147);
nand U23335 (N_23335,N_21867,N_20882);
xor U23336 (N_23336,N_21572,N_20681);
or U23337 (N_23337,N_20959,N_21862);
nand U23338 (N_23338,N_20175,N_20150);
and U23339 (N_23339,N_20822,N_20582);
and U23340 (N_23340,N_20535,N_20196);
nor U23341 (N_23341,N_21220,N_20875);
nand U23342 (N_23342,N_21323,N_21856);
or U23343 (N_23343,N_20707,N_21222);
or U23344 (N_23344,N_21894,N_20344);
nor U23345 (N_23345,N_20528,N_20681);
and U23346 (N_23346,N_21154,N_21791);
or U23347 (N_23347,N_20060,N_20755);
nor U23348 (N_23348,N_21930,N_21753);
nor U23349 (N_23349,N_21776,N_21197);
or U23350 (N_23350,N_20533,N_21880);
xor U23351 (N_23351,N_20768,N_20247);
nor U23352 (N_23352,N_21571,N_21975);
nor U23353 (N_23353,N_21119,N_21992);
xor U23354 (N_23354,N_20562,N_20719);
nor U23355 (N_23355,N_21444,N_21790);
xnor U23356 (N_23356,N_20944,N_21261);
or U23357 (N_23357,N_21327,N_20333);
or U23358 (N_23358,N_20411,N_21960);
nor U23359 (N_23359,N_20049,N_20220);
or U23360 (N_23360,N_21367,N_20011);
and U23361 (N_23361,N_21106,N_21144);
nor U23362 (N_23362,N_20580,N_20542);
and U23363 (N_23363,N_21586,N_20662);
nor U23364 (N_23364,N_20235,N_20800);
xor U23365 (N_23365,N_20555,N_20104);
nand U23366 (N_23366,N_21548,N_20641);
or U23367 (N_23367,N_20482,N_20708);
and U23368 (N_23368,N_20462,N_21206);
xor U23369 (N_23369,N_21667,N_21357);
xnor U23370 (N_23370,N_20012,N_20181);
nor U23371 (N_23371,N_21459,N_21457);
xor U23372 (N_23372,N_21436,N_21729);
xor U23373 (N_23373,N_20843,N_20020);
nand U23374 (N_23374,N_20340,N_21597);
or U23375 (N_23375,N_21756,N_20096);
nand U23376 (N_23376,N_21800,N_20933);
nand U23377 (N_23377,N_21798,N_21360);
xnor U23378 (N_23378,N_20193,N_20123);
and U23379 (N_23379,N_21321,N_20366);
nor U23380 (N_23380,N_20439,N_20565);
xor U23381 (N_23381,N_21632,N_21506);
nand U23382 (N_23382,N_20388,N_21539);
or U23383 (N_23383,N_21505,N_20018);
xor U23384 (N_23384,N_21325,N_20812);
nand U23385 (N_23385,N_20310,N_20243);
and U23386 (N_23386,N_21189,N_21860);
and U23387 (N_23387,N_20108,N_21458);
and U23388 (N_23388,N_21264,N_21207);
and U23389 (N_23389,N_21751,N_21770);
and U23390 (N_23390,N_21966,N_20490);
xor U23391 (N_23391,N_21549,N_21124);
nor U23392 (N_23392,N_20212,N_21511);
nand U23393 (N_23393,N_21911,N_21782);
nand U23394 (N_23394,N_20595,N_20201);
nor U23395 (N_23395,N_21396,N_21592);
and U23396 (N_23396,N_20401,N_20438);
nor U23397 (N_23397,N_20600,N_21208);
nor U23398 (N_23398,N_21620,N_21426);
and U23399 (N_23399,N_21115,N_20202);
or U23400 (N_23400,N_21105,N_20750);
nor U23401 (N_23401,N_21344,N_21181);
xnor U23402 (N_23402,N_20070,N_21223);
and U23403 (N_23403,N_20844,N_21381);
nor U23404 (N_23404,N_20079,N_21214);
or U23405 (N_23405,N_20316,N_20450);
nor U23406 (N_23406,N_21948,N_20732);
or U23407 (N_23407,N_21546,N_20866);
xor U23408 (N_23408,N_20928,N_20514);
and U23409 (N_23409,N_21747,N_21680);
or U23410 (N_23410,N_21473,N_21902);
or U23411 (N_23411,N_21735,N_21042);
and U23412 (N_23412,N_20805,N_21181);
or U23413 (N_23413,N_21423,N_20821);
and U23414 (N_23414,N_21280,N_21661);
xor U23415 (N_23415,N_21943,N_21593);
xnor U23416 (N_23416,N_20022,N_21205);
and U23417 (N_23417,N_21950,N_20797);
nor U23418 (N_23418,N_20615,N_21112);
and U23419 (N_23419,N_21725,N_20580);
xor U23420 (N_23420,N_21586,N_20863);
xor U23421 (N_23421,N_21531,N_20525);
and U23422 (N_23422,N_20629,N_21329);
nand U23423 (N_23423,N_21040,N_20646);
and U23424 (N_23424,N_20905,N_20326);
xnor U23425 (N_23425,N_20099,N_21362);
xnor U23426 (N_23426,N_20340,N_20446);
nand U23427 (N_23427,N_21530,N_21628);
xor U23428 (N_23428,N_20786,N_20276);
or U23429 (N_23429,N_21895,N_20838);
nand U23430 (N_23430,N_21619,N_20344);
xnor U23431 (N_23431,N_21333,N_21661);
and U23432 (N_23432,N_20877,N_21917);
and U23433 (N_23433,N_21591,N_20448);
nor U23434 (N_23434,N_20129,N_21980);
nand U23435 (N_23435,N_21203,N_21182);
nor U23436 (N_23436,N_20622,N_21942);
nor U23437 (N_23437,N_21155,N_20258);
nand U23438 (N_23438,N_21239,N_21738);
nand U23439 (N_23439,N_20245,N_21112);
nor U23440 (N_23440,N_21824,N_21698);
or U23441 (N_23441,N_20216,N_20476);
or U23442 (N_23442,N_20402,N_21701);
nand U23443 (N_23443,N_21625,N_20734);
nand U23444 (N_23444,N_21092,N_21173);
nand U23445 (N_23445,N_21280,N_21225);
xnor U23446 (N_23446,N_21627,N_21010);
nor U23447 (N_23447,N_21323,N_20801);
and U23448 (N_23448,N_21004,N_21319);
nor U23449 (N_23449,N_20649,N_21766);
nand U23450 (N_23450,N_20296,N_21799);
xnor U23451 (N_23451,N_20473,N_21717);
nor U23452 (N_23452,N_20184,N_20277);
nand U23453 (N_23453,N_21541,N_20311);
and U23454 (N_23454,N_21370,N_21672);
nor U23455 (N_23455,N_21210,N_21903);
and U23456 (N_23456,N_20458,N_20812);
xor U23457 (N_23457,N_20634,N_20467);
and U23458 (N_23458,N_20169,N_20476);
xnor U23459 (N_23459,N_20514,N_20473);
nand U23460 (N_23460,N_20581,N_21001);
and U23461 (N_23461,N_21074,N_20500);
and U23462 (N_23462,N_20937,N_20712);
and U23463 (N_23463,N_21117,N_21182);
nand U23464 (N_23464,N_21094,N_20153);
nor U23465 (N_23465,N_21816,N_20924);
nor U23466 (N_23466,N_20322,N_20344);
nand U23467 (N_23467,N_20812,N_20723);
and U23468 (N_23468,N_21506,N_20381);
and U23469 (N_23469,N_21016,N_21440);
xor U23470 (N_23470,N_21563,N_21706);
or U23471 (N_23471,N_20034,N_20288);
nor U23472 (N_23472,N_20757,N_20180);
xor U23473 (N_23473,N_21356,N_21456);
xor U23474 (N_23474,N_20017,N_21660);
nand U23475 (N_23475,N_21940,N_20686);
or U23476 (N_23476,N_21430,N_20920);
nand U23477 (N_23477,N_21025,N_20847);
xor U23478 (N_23478,N_20881,N_21201);
and U23479 (N_23479,N_21392,N_20750);
or U23480 (N_23480,N_20533,N_20871);
and U23481 (N_23481,N_20961,N_21900);
nor U23482 (N_23482,N_20283,N_21020);
or U23483 (N_23483,N_20577,N_21009);
nand U23484 (N_23484,N_21138,N_20576);
and U23485 (N_23485,N_20361,N_20543);
or U23486 (N_23486,N_20956,N_20619);
nor U23487 (N_23487,N_20690,N_21932);
or U23488 (N_23488,N_21171,N_20547);
xnor U23489 (N_23489,N_20034,N_20103);
nor U23490 (N_23490,N_20886,N_21335);
and U23491 (N_23491,N_20655,N_20693);
or U23492 (N_23492,N_20905,N_21854);
nor U23493 (N_23493,N_21255,N_20569);
nand U23494 (N_23494,N_21144,N_20045);
and U23495 (N_23495,N_21510,N_20891);
nor U23496 (N_23496,N_20283,N_20939);
nor U23497 (N_23497,N_21154,N_20734);
nand U23498 (N_23498,N_20991,N_20647);
xnor U23499 (N_23499,N_20589,N_20244);
and U23500 (N_23500,N_21920,N_20318);
nor U23501 (N_23501,N_20274,N_21935);
and U23502 (N_23502,N_21878,N_21043);
nand U23503 (N_23503,N_20993,N_21062);
and U23504 (N_23504,N_20769,N_20794);
and U23505 (N_23505,N_20287,N_20962);
nor U23506 (N_23506,N_20773,N_21457);
xnor U23507 (N_23507,N_21137,N_20098);
nand U23508 (N_23508,N_21290,N_20408);
and U23509 (N_23509,N_21609,N_20990);
or U23510 (N_23510,N_21195,N_21857);
xor U23511 (N_23511,N_21375,N_21532);
xor U23512 (N_23512,N_21729,N_21632);
nor U23513 (N_23513,N_21267,N_20356);
xnor U23514 (N_23514,N_21841,N_20784);
nor U23515 (N_23515,N_21970,N_21680);
nor U23516 (N_23516,N_20826,N_21585);
nor U23517 (N_23517,N_20054,N_20797);
and U23518 (N_23518,N_21247,N_20512);
nand U23519 (N_23519,N_21814,N_21636);
xor U23520 (N_23520,N_21786,N_21130);
nand U23521 (N_23521,N_21728,N_21087);
and U23522 (N_23522,N_21999,N_21206);
xor U23523 (N_23523,N_20927,N_20590);
or U23524 (N_23524,N_21851,N_21431);
and U23525 (N_23525,N_20560,N_20634);
and U23526 (N_23526,N_21139,N_21158);
or U23527 (N_23527,N_20577,N_21008);
xnor U23528 (N_23528,N_21259,N_21553);
nor U23529 (N_23529,N_21376,N_21081);
nand U23530 (N_23530,N_21031,N_21520);
nand U23531 (N_23531,N_20833,N_20483);
nor U23532 (N_23532,N_21614,N_21344);
or U23533 (N_23533,N_21542,N_20934);
nor U23534 (N_23534,N_20662,N_21706);
nand U23535 (N_23535,N_21932,N_20855);
nand U23536 (N_23536,N_21097,N_20411);
nor U23537 (N_23537,N_20109,N_21153);
xor U23538 (N_23538,N_20891,N_21250);
nor U23539 (N_23539,N_20923,N_21599);
nand U23540 (N_23540,N_21029,N_21282);
nor U23541 (N_23541,N_21757,N_20134);
nor U23542 (N_23542,N_21889,N_21753);
and U23543 (N_23543,N_21503,N_21341);
nor U23544 (N_23544,N_21563,N_21121);
nand U23545 (N_23545,N_21766,N_21706);
nand U23546 (N_23546,N_21812,N_20497);
nor U23547 (N_23547,N_20103,N_21398);
or U23548 (N_23548,N_21073,N_20135);
or U23549 (N_23549,N_21146,N_21747);
nor U23550 (N_23550,N_21459,N_20538);
nand U23551 (N_23551,N_21757,N_21673);
nor U23552 (N_23552,N_21890,N_21830);
nor U23553 (N_23553,N_21527,N_21765);
xor U23554 (N_23554,N_20180,N_21980);
and U23555 (N_23555,N_20911,N_21257);
and U23556 (N_23556,N_20725,N_21470);
or U23557 (N_23557,N_21878,N_21298);
and U23558 (N_23558,N_20450,N_20394);
or U23559 (N_23559,N_21064,N_21386);
and U23560 (N_23560,N_21751,N_20678);
nor U23561 (N_23561,N_20860,N_20656);
xor U23562 (N_23562,N_20587,N_21441);
or U23563 (N_23563,N_21015,N_21258);
nor U23564 (N_23564,N_21882,N_21724);
nand U23565 (N_23565,N_21200,N_20941);
xor U23566 (N_23566,N_20995,N_20578);
nand U23567 (N_23567,N_21298,N_21731);
xor U23568 (N_23568,N_21096,N_21672);
xor U23569 (N_23569,N_20334,N_20753);
xnor U23570 (N_23570,N_20824,N_21198);
or U23571 (N_23571,N_21729,N_21643);
and U23572 (N_23572,N_21367,N_20817);
and U23573 (N_23573,N_21010,N_21317);
or U23574 (N_23574,N_20209,N_21900);
nor U23575 (N_23575,N_21730,N_21563);
xnor U23576 (N_23576,N_21345,N_20101);
and U23577 (N_23577,N_21552,N_21429);
nand U23578 (N_23578,N_20160,N_21294);
nand U23579 (N_23579,N_21602,N_21448);
xor U23580 (N_23580,N_20231,N_21389);
nand U23581 (N_23581,N_20063,N_20236);
nor U23582 (N_23582,N_21588,N_21154);
and U23583 (N_23583,N_21649,N_21493);
nor U23584 (N_23584,N_20981,N_20496);
nor U23585 (N_23585,N_20236,N_20580);
nor U23586 (N_23586,N_20601,N_21910);
or U23587 (N_23587,N_20195,N_21346);
nand U23588 (N_23588,N_21905,N_21639);
and U23589 (N_23589,N_20592,N_21586);
nand U23590 (N_23590,N_20717,N_21585);
and U23591 (N_23591,N_20613,N_21451);
nor U23592 (N_23592,N_21808,N_20979);
and U23593 (N_23593,N_20960,N_21000);
nor U23594 (N_23594,N_21366,N_21700);
nor U23595 (N_23595,N_20135,N_20725);
nor U23596 (N_23596,N_20114,N_20785);
nor U23597 (N_23597,N_21329,N_21338);
or U23598 (N_23598,N_21536,N_21927);
xor U23599 (N_23599,N_21643,N_20539);
or U23600 (N_23600,N_20289,N_21669);
and U23601 (N_23601,N_20318,N_21381);
or U23602 (N_23602,N_20157,N_21761);
or U23603 (N_23603,N_21139,N_21209);
or U23604 (N_23604,N_20108,N_20519);
and U23605 (N_23605,N_21504,N_21731);
nand U23606 (N_23606,N_21765,N_21420);
nor U23607 (N_23607,N_21067,N_21744);
nor U23608 (N_23608,N_20391,N_20186);
and U23609 (N_23609,N_21585,N_21751);
or U23610 (N_23610,N_20204,N_21278);
xnor U23611 (N_23611,N_21085,N_21173);
and U23612 (N_23612,N_21310,N_20442);
or U23613 (N_23613,N_20781,N_21692);
nor U23614 (N_23614,N_20244,N_21599);
nand U23615 (N_23615,N_20871,N_20344);
nor U23616 (N_23616,N_20394,N_21266);
xnor U23617 (N_23617,N_21997,N_21918);
nand U23618 (N_23618,N_21773,N_21345);
and U23619 (N_23619,N_20239,N_21156);
and U23620 (N_23620,N_21153,N_21915);
nor U23621 (N_23621,N_20645,N_20558);
nand U23622 (N_23622,N_20437,N_20376);
nor U23623 (N_23623,N_20350,N_21627);
or U23624 (N_23624,N_20920,N_20800);
nand U23625 (N_23625,N_21039,N_20773);
xor U23626 (N_23626,N_21005,N_20810);
and U23627 (N_23627,N_20845,N_21781);
nand U23628 (N_23628,N_21108,N_21531);
or U23629 (N_23629,N_21550,N_20983);
nor U23630 (N_23630,N_21471,N_20351);
and U23631 (N_23631,N_20475,N_21554);
or U23632 (N_23632,N_21154,N_21911);
and U23633 (N_23633,N_21901,N_21414);
and U23634 (N_23634,N_20488,N_21291);
nor U23635 (N_23635,N_21127,N_20313);
nand U23636 (N_23636,N_20900,N_21164);
nand U23637 (N_23637,N_20443,N_20236);
nand U23638 (N_23638,N_21736,N_20328);
nor U23639 (N_23639,N_20354,N_20718);
or U23640 (N_23640,N_21396,N_21126);
or U23641 (N_23641,N_21814,N_20619);
nand U23642 (N_23642,N_21783,N_21785);
xnor U23643 (N_23643,N_21733,N_20747);
nor U23644 (N_23644,N_20457,N_21786);
or U23645 (N_23645,N_20598,N_21648);
or U23646 (N_23646,N_21646,N_20701);
nor U23647 (N_23647,N_20516,N_20756);
xnor U23648 (N_23648,N_20305,N_20976);
and U23649 (N_23649,N_20700,N_20080);
nand U23650 (N_23650,N_21513,N_20188);
or U23651 (N_23651,N_20479,N_20520);
nor U23652 (N_23652,N_20706,N_20876);
nand U23653 (N_23653,N_20676,N_20905);
nor U23654 (N_23654,N_20812,N_21912);
nor U23655 (N_23655,N_20133,N_21117);
or U23656 (N_23656,N_21111,N_21168);
xnor U23657 (N_23657,N_21402,N_20176);
nand U23658 (N_23658,N_20293,N_21649);
or U23659 (N_23659,N_20980,N_20284);
nor U23660 (N_23660,N_20713,N_20951);
nand U23661 (N_23661,N_20589,N_21641);
and U23662 (N_23662,N_21769,N_20845);
and U23663 (N_23663,N_20153,N_21755);
or U23664 (N_23664,N_20969,N_21537);
xor U23665 (N_23665,N_20226,N_21269);
nand U23666 (N_23666,N_20888,N_20423);
nand U23667 (N_23667,N_21258,N_20888);
xnor U23668 (N_23668,N_21029,N_20066);
or U23669 (N_23669,N_21629,N_20563);
nor U23670 (N_23670,N_20724,N_20623);
or U23671 (N_23671,N_20349,N_21861);
xor U23672 (N_23672,N_20672,N_21932);
or U23673 (N_23673,N_21971,N_20494);
and U23674 (N_23674,N_20756,N_21217);
nand U23675 (N_23675,N_21864,N_21396);
or U23676 (N_23676,N_21996,N_20577);
and U23677 (N_23677,N_21768,N_20535);
nand U23678 (N_23678,N_21377,N_21701);
nor U23679 (N_23679,N_20398,N_21739);
nor U23680 (N_23680,N_21976,N_21835);
and U23681 (N_23681,N_20949,N_21272);
or U23682 (N_23682,N_21742,N_21859);
nand U23683 (N_23683,N_20139,N_20906);
and U23684 (N_23684,N_21294,N_20033);
nor U23685 (N_23685,N_21435,N_21793);
xnor U23686 (N_23686,N_20929,N_21819);
nor U23687 (N_23687,N_21847,N_20807);
xnor U23688 (N_23688,N_20543,N_21268);
xnor U23689 (N_23689,N_21242,N_20888);
nor U23690 (N_23690,N_20253,N_20639);
or U23691 (N_23691,N_21800,N_20094);
and U23692 (N_23692,N_21228,N_21258);
or U23693 (N_23693,N_20065,N_21658);
xor U23694 (N_23694,N_20703,N_20091);
nor U23695 (N_23695,N_21904,N_20701);
or U23696 (N_23696,N_20987,N_20353);
or U23697 (N_23697,N_20767,N_20299);
nor U23698 (N_23698,N_21004,N_21576);
and U23699 (N_23699,N_20473,N_21373);
nor U23700 (N_23700,N_21604,N_20492);
and U23701 (N_23701,N_21868,N_21645);
nand U23702 (N_23702,N_20179,N_20644);
or U23703 (N_23703,N_21707,N_21084);
xor U23704 (N_23704,N_20281,N_21918);
nand U23705 (N_23705,N_21762,N_21902);
xnor U23706 (N_23706,N_21003,N_21615);
nand U23707 (N_23707,N_20411,N_20004);
or U23708 (N_23708,N_20468,N_21964);
nor U23709 (N_23709,N_21043,N_20947);
xnor U23710 (N_23710,N_20649,N_20261);
nand U23711 (N_23711,N_21185,N_20354);
xor U23712 (N_23712,N_20100,N_20160);
nor U23713 (N_23713,N_21480,N_20834);
nor U23714 (N_23714,N_20275,N_21317);
xor U23715 (N_23715,N_20116,N_20031);
xor U23716 (N_23716,N_20937,N_21784);
or U23717 (N_23717,N_20369,N_20874);
nand U23718 (N_23718,N_21083,N_21801);
and U23719 (N_23719,N_20403,N_20631);
nor U23720 (N_23720,N_21876,N_21437);
nand U23721 (N_23721,N_20760,N_20041);
nor U23722 (N_23722,N_21161,N_20093);
nor U23723 (N_23723,N_20636,N_21130);
xor U23724 (N_23724,N_20534,N_20990);
or U23725 (N_23725,N_20111,N_21452);
or U23726 (N_23726,N_21883,N_21148);
nor U23727 (N_23727,N_21157,N_21114);
nand U23728 (N_23728,N_21853,N_20672);
or U23729 (N_23729,N_20192,N_21194);
or U23730 (N_23730,N_21570,N_20050);
nand U23731 (N_23731,N_21980,N_20021);
or U23732 (N_23732,N_20516,N_20022);
xnor U23733 (N_23733,N_20557,N_21746);
xor U23734 (N_23734,N_21348,N_21155);
and U23735 (N_23735,N_21767,N_20125);
nand U23736 (N_23736,N_20369,N_21385);
nor U23737 (N_23737,N_21081,N_20183);
xor U23738 (N_23738,N_20868,N_20520);
and U23739 (N_23739,N_20709,N_20383);
and U23740 (N_23740,N_20348,N_20411);
nor U23741 (N_23741,N_20281,N_20693);
and U23742 (N_23742,N_21910,N_21560);
xnor U23743 (N_23743,N_20071,N_20284);
xor U23744 (N_23744,N_21301,N_21909);
xor U23745 (N_23745,N_20026,N_20272);
or U23746 (N_23746,N_20123,N_21112);
or U23747 (N_23747,N_20949,N_21714);
and U23748 (N_23748,N_20692,N_21294);
nand U23749 (N_23749,N_20501,N_21888);
nor U23750 (N_23750,N_20574,N_20501);
and U23751 (N_23751,N_20803,N_21802);
xor U23752 (N_23752,N_20132,N_20198);
xnor U23753 (N_23753,N_21031,N_20995);
and U23754 (N_23754,N_21716,N_21522);
xnor U23755 (N_23755,N_20742,N_21137);
and U23756 (N_23756,N_20442,N_21570);
or U23757 (N_23757,N_21674,N_20611);
and U23758 (N_23758,N_21788,N_21014);
and U23759 (N_23759,N_20395,N_20433);
or U23760 (N_23760,N_21527,N_20440);
nor U23761 (N_23761,N_21080,N_21316);
xnor U23762 (N_23762,N_20489,N_21063);
xnor U23763 (N_23763,N_20603,N_20881);
xor U23764 (N_23764,N_21184,N_20757);
and U23765 (N_23765,N_21253,N_20774);
and U23766 (N_23766,N_20711,N_21325);
and U23767 (N_23767,N_21931,N_20252);
or U23768 (N_23768,N_20804,N_20149);
nand U23769 (N_23769,N_21549,N_21592);
and U23770 (N_23770,N_20004,N_21632);
nand U23771 (N_23771,N_20899,N_20477);
nand U23772 (N_23772,N_20438,N_20421);
and U23773 (N_23773,N_20283,N_21923);
nor U23774 (N_23774,N_20412,N_20470);
nand U23775 (N_23775,N_20871,N_21429);
nand U23776 (N_23776,N_20866,N_21858);
or U23777 (N_23777,N_20618,N_21898);
xor U23778 (N_23778,N_20600,N_21842);
nand U23779 (N_23779,N_21439,N_21808);
and U23780 (N_23780,N_20158,N_21776);
or U23781 (N_23781,N_20364,N_20063);
nor U23782 (N_23782,N_21925,N_20248);
or U23783 (N_23783,N_21962,N_20202);
or U23784 (N_23784,N_21117,N_21183);
nand U23785 (N_23785,N_21168,N_21407);
or U23786 (N_23786,N_21569,N_20689);
and U23787 (N_23787,N_21362,N_21209);
or U23788 (N_23788,N_20334,N_20027);
nand U23789 (N_23789,N_20698,N_21018);
nand U23790 (N_23790,N_20920,N_20397);
nand U23791 (N_23791,N_20500,N_21921);
and U23792 (N_23792,N_21409,N_20216);
xnor U23793 (N_23793,N_21597,N_21208);
nand U23794 (N_23794,N_21294,N_20746);
and U23795 (N_23795,N_20326,N_20484);
and U23796 (N_23796,N_21689,N_21667);
nand U23797 (N_23797,N_21793,N_20618);
or U23798 (N_23798,N_20642,N_21120);
nand U23799 (N_23799,N_20174,N_20287);
nand U23800 (N_23800,N_20492,N_20494);
nand U23801 (N_23801,N_20903,N_20560);
nand U23802 (N_23802,N_20324,N_21757);
and U23803 (N_23803,N_21991,N_21577);
nor U23804 (N_23804,N_21499,N_20798);
xor U23805 (N_23805,N_21652,N_21140);
nor U23806 (N_23806,N_21840,N_21649);
nand U23807 (N_23807,N_20607,N_21555);
xor U23808 (N_23808,N_21756,N_20212);
nor U23809 (N_23809,N_21127,N_20202);
nor U23810 (N_23810,N_21255,N_20360);
and U23811 (N_23811,N_20288,N_20286);
and U23812 (N_23812,N_21056,N_21511);
or U23813 (N_23813,N_21129,N_20902);
nor U23814 (N_23814,N_20414,N_20410);
nand U23815 (N_23815,N_21630,N_21856);
xnor U23816 (N_23816,N_21050,N_21927);
nand U23817 (N_23817,N_20436,N_21427);
xor U23818 (N_23818,N_21006,N_21364);
nand U23819 (N_23819,N_21843,N_21996);
nor U23820 (N_23820,N_21575,N_20444);
nor U23821 (N_23821,N_20586,N_21934);
nor U23822 (N_23822,N_20991,N_21542);
nor U23823 (N_23823,N_21796,N_20113);
or U23824 (N_23824,N_20006,N_20395);
nand U23825 (N_23825,N_21664,N_20736);
nor U23826 (N_23826,N_21018,N_20043);
and U23827 (N_23827,N_21207,N_21997);
or U23828 (N_23828,N_20243,N_20020);
and U23829 (N_23829,N_21895,N_20421);
or U23830 (N_23830,N_20913,N_20184);
nand U23831 (N_23831,N_21270,N_20657);
nor U23832 (N_23832,N_21485,N_20604);
nand U23833 (N_23833,N_21285,N_20392);
xnor U23834 (N_23834,N_21576,N_21557);
and U23835 (N_23835,N_20174,N_20303);
xnor U23836 (N_23836,N_20533,N_20789);
or U23837 (N_23837,N_21504,N_20937);
xnor U23838 (N_23838,N_21803,N_20284);
xor U23839 (N_23839,N_20394,N_21293);
nand U23840 (N_23840,N_21105,N_20598);
nor U23841 (N_23841,N_20800,N_20769);
xnor U23842 (N_23842,N_21584,N_20127);
or U23843 (N_23843,N_21877,N_20168);
nand U23844 (N_23844,N_21779,N_21829);
and U23845 (N_23845,N_21400,N_20832);
nor U23846 (N_23846,N_20245,N_20484);
nor U23847 (N_23847,N_20967,N_20635);
nand U23848 (N_23848,N_21696,N_21503);
or U23849 (N_23849,N_20251,N_21551);
xor U23850 (N_23850,N_21690,N_21912);
or U23851 (N_23851,N_21430,N_21572);
and U23852 (N_23852,N_21865,N_21712);
nand U23853 (N_23853,N_21742,N_20694);
nor U23854 (N_23854,N_20030,N_20264);
or U23855 (N_23855,N_20953,N_21886);
nor U23856 (N_23856,N_20911,N_21873);
or U23857 (N_23857,N_21821,N_21613);
and U23858 (N_23858,N_20442,N_21163);
xor U23859 (N_23859,N_20137,N_20435);
or U23860 (N_23860,N_20626,N_20575);
or U23861 (N_23861,N_20781,N_20488);
or U23862 (N_23862,N_21306,N_21241);
or U23863 (N_23863,N_21404,N_20462);
and U23864 (N_23864,N_20714,N_20394);
xnor U23865 (N_23865,N_20987,N_20193);
or U23866 (N_23866,N_20923,N_21311);
and U23867 (N_23867,N_21546,N_21416);
xnor U23868 (N_23868,N_21334,N_21014);
nor U23869 (N_23869,N_21410,N_20240);
nand U23870 (N_23870,N_21267,N_20852);
nand U23871 (N_23871,N_20449,N_20062);
or U23872 (N_23872,N_20690,N_20355);
nor U23873 (N_23873,N_21578,N_20593);
or U23874 (N_23874,N_20203,N_20703);
xor U23875 (N_23875,N_21489,N_20745);
or U23876 (N_23876,N_21376,N_21223);
xor U23877 (N_23877,N_20896,N_21201);
nand U23878 (N_23878,N_21025,N_20022);
nand U23879 (N_23879,N_20509,N_20802);
nand U23880 (N_23880,N_21261,N_21671);
nand U23881 (N_23881,N_21996,N_20008);
nand U23882 (N_23882,N_20361,N_20410);
and U23883 (N_23883,N_20967,N_21308);
xnor U23884 (N_23884,N_20972,N_20671);
xor U23885 (N_23885,N_21317,N_21356);
xor U23886 (N_23886,N_21775,N_20077);
nor U23887 (N_23887,N_20667,N_21313);
nor U23888 (N_23888,N_20107,N_20020);
nand U23889 (N_23889,N_21083,N_21346);
and U23890 (N_23890,N_20668,N_20872);
or U23891 (N_23891,N_21835,N_20742);
nand U23892 (N_23892,N_21161,N_21795);
xnor U23893 (N_23893,N_20618,N_20995);
or U23894 (N_23894,N_20437,N_21892);
nand U23895 (N_23895,N_20532,N_20317);
nand U23896 (N_23896,N_20842,N_20581);
and U23897 (N_23897,N_20247,N_21427);
nor U23898 (N_23898,N_20923,N_21746);
nor U23899 (N_23899,N_21851,N_20709);
xor U23900 (N_23900,N_20772,N_21076);
nand U23901 (N_23901,N_21554,N_20778);
and U23902 (N_23902,N_21893,N_20487);
nand U23903 (N_23903,N_21717,N_20156);
nor U23904 (N_23904,N_21202,N_20740);
or U23905 (N_23905,N_20929,N_20543);
nor U23906 (N_23906,N_20894,N_20646);
nand U23907 (N_23907,N_20935,N_21235);
or U23908 (N_23908,N_20224,N_21528);
or U23909 (N_23909,N_20983,N_21160);
xor U23910 (N_23910,N_21436,N_21647);
nand U23911 (N_23911,N_20968,N_21364);
and U23912 (N_23912,N_20080,N_20632);
nand U23913 (N_23913,N_20131,N_20407);
and U23914 (N_23914,N_20108,N_20712);
xnor U23915 (N_23915,N_20969,N_20454);
xnor U23916 (N_23916,N_21887,N_21067);
nand U23917 (N_23917,N_20616,N_20239);
nand U23918 (N_23918,N_20455,N_21432);
and U23919 (N_23919,N_21788,N_21486);
nor U23920 (N_23920,N_21065,N_20596);
xor U23921 (N_23921,N_21453,N_21257);
nand U23922 (N_23922,N_21750,N_20177);
nand U23923 (N_23923,N_20627,N_20372);
or U23924 (N_23924,N_21238,N_20982);
nand U23925 (N_23925,N_20922,N_20779);
nand U23926 (N_23926,N_20446,N_21352);
nor U23927 (N_23927,N_21045,N_20448);
or U23928 (N_23928,N_21144,N_21232);
nand U23929 (N_23929,N_21306,N_20092);
and U23930 (N_23930,N_21401,N_21766);
xnor U23931 (N_23931,N_21960,N_21650);
nor U23932 (N_23932,N_20924,N_21328);
nand U23933 (N_23933,N_21372,N_20951);
or U23934 (N_23934,N_20022,N_21005);
nand U23935 (N_23935,N_20691,N_21509);
and U23936 (N_23936,N_20018,N_20026);
and U23937 (N_23937,N_21512,N_21615);
nor U23938 (N_23938,N_20168,N_20062);
xnor U23939 (N_23939,N_21869,N_21563);
nor U23940 (N_23940,N_21819,N_21214);
or U23941 (N_23941,N_21427,N_21434);
and U23942 (N_23942,N_21688,N_21941);
or U23943 (N_23943,N_21471,N_20360);
nand U23944 (N_23944,N_21719,N_21535);
xnor U23945 (N_23945,N_20251,N_21582);
and U23946 (N_23946,N_21719,N_20175);
xor U23947 (N_23947,N_20543,N_21479);
and U23948 (N_23948,N_21743,N_20406);
nor U23949 (N_23949,N_20989,N_21329);
nor U23950 (N_23950,N_21930,N_21515);
and U23951 (N_23951,N_21411,N_20060);
nor U23952 (N_23952,N_20655,N_21313);
xnor U23953 (N_23953,N_20075,N_21238);
xnor U23954 (N_23954,N_21904,N_21271);
xnor U23955 (N_23955,N_21457,N_21208);
nor U23956 (N_23956,N_20828,N_21181);
nor U23957 (N_23957,N_20513,N_20909);
nand U23958 (N_23958,N_21599,N_21485);
or U23959 (N_23959,N_21208,N_21270);
or U23960 (N_23960,N_21476,N_20455);
nand U23961 (N_23961,N_21969,N_21533);
xor U23962 (N_23962,N_20891,N_20384);
nand U23963 (N_23963,N_20163,N_20969);
nor U23964 (N_23964,N_20275,N_21708);
and U23965 (N_23965,N_21287,N_20695);
or U23966 (N_23966,N_20373,N_21172);
and U23967 (N_23967,N_21852,N_21256);
nor U23968 (N_23968,N_20316,N_21233);
nand U23969 (N_23969,N_20484,N_21486);
and U23970 (N_23970,N_21304,N_20122);
and U23971 (N_23971,N_21004,N_20276);
nand U23972 (N_23972,N_20233,N_21729);
xnor U23973 (N_23973,N_21583,N_20721);
and U23974 (N_23974,N_21214,N_20409);
xor U23975 (N_23975,N_20452,N_21882);
nand U23976 (N_23976,N_21578,N_20148);
and U23977 (N_23977,N_21389,N_21186);
or U23978 (N_23978,N_20560,N_21885);
and U23979 (N_23979,N_20981,N_20890);
xnor U23980 (N_23980,N_21785,N_20543);
or U23981 (N_23981,N_20293,N_20476);
nand U23982 (N_23982,N_21562,N_20430);
nand U23983 (N_23983,N_21979,N_20846);
or U23984 (N_23984,N_20818,N_21082);
xor U23985 (N_23985,N_20276,N_20275);
nand U23986 (N_23986,N_20097,N_21834);
nor U23987 (N_23987,N_20339,N_21665);
and U23988 (N_23988,N_20681,N_20572);
or U23989 (N_23989,N_20155,N_20366);
nand U23990 (N_23990,N_21427,N_20980);
or U23991 (N_23991,N_20319,N_21023);
nand U23992 (N_23992,N_21940,N_21832);
or U23993 (N_23993,N_20674,N_20395);
or U23994 (N_23994,N_20511,N_21196);
xnor U23995 (N_23995,N_21877,N_21792);
and U23996 (N_23996,N_21778,N_21465);
and U23997 (N_23997,N_20821,N_21191);
nand U23998 (N_23998,N_20471,N_21068);
and U23999 (N_23999,N_21922,N_20345);
nor U24000 (N_24000,N_23110,N_22083);
nor U24001 (N_24001,N_23730,N_23539);
nor U24002 (N_24002,N_23326,N_23302);
or U24003 (N_24003,N_22625,N_22041);
and U24004 (N_24004,N_22744,N_23363);
xor U24005 (N_24005,N_22296,N_23499);
xnor U24006 (N_24006,N_22954,N_23025);
or U24007 (N_24007,N_23323,N_23941);
nand U24008 (N_24008,N_22000,N_22366);
nor U24009 (N_24009,N_23868,N_22938);
and U24010 (N_24010,N_23999,N_22817);
nand U24011 (N_24011,N_22726,N_23954);
xor U24012 (N_24012,N_22654,N_22620);
nor U24013 (N_24013,N_22202,N_23918);
nor U24014 (N_24014,N_23117,N_22847);
or U24015 (N_24015,N_22866,N_22788);
xor U24016 (N_24016,N_22660,N_22405);
and U24017 (N_24017,N_22646,N_23344);
nand U24018 (N_24018,N_23938,N_23692);
nor U24019 (N_24019,N_22207,N_22250);
or U24020 (N_24020,N_22926,N_22306);
and U24021 (N_24021,N_22699,N_22843);
nor U24022 (N_24022,N_22570,N_23542);
or U24023 (N_24023,N_23257,N_22786);
and U24024 (N_24024,N_22868,N_23787);
or U24025 (N_24025,N_23811,N_22446);
nor U24026 (N_24026,N_22059,N_23501);
nor U24027 (N_24027,N_22171,N_23333);
and U24028 (N_24028,N_23669,N_23582);
or U24029 (N_24029,N_23906,N_23545);
nor U24030 (N_24030,N_23482,N_22696);
xnor U24031 (N_24031,N_23795,N_23554);
nand U24032 (N_24032,N_23822,N_23907);
nor U24033 (N_24033,N_22402,N_23076);
nor U24034 (N_24034,N_23672,N_22193);
nand U24035 (N_24035,N_22502,N_22476);
nor U24036 (N_24036,N_22747,N_22679);
and U24037 (N_24037,N_22604,N_23518);
nor U24038 (N_24038,N_23424,N_23088);
or U24039 (N_24039,N_22712,N_22731);
nand U24040 (N_24040,N_22451,N_22822);
nor U24041 (N_24041,N_23712,N_22203);
or U24042 (N_24042,N_23421,N_22267);
and U24043 (N_24043,N_23320,N_22572);
and U24044 (N_24044,N_22839,N_22629);
xnor U24045 (N_24045,N_23523,N_23564);
xor U24046 (N_24046,N_23022,N_22903);
xor U24047 (N_24047,N_22997,N_22720);
or U24048 (N_24048,N_23119,N_22020);
nor U24049 (N_24049,N_23782,N_23218);
or U24050 (N_24050,N_22481,N_23816);
nand U24051 (N_24051,N_22634,N_22872);
nand U24052 (N_24052,N_23735,N_22040);
or U24053 (N_24053,N_23940,N_23338);
and U24054 (N_24054,N_23580,N_22915);
nor U24055 (N_24055,N_22844,N_22790);
or U24056 (N_24056,N_22220,N_23736);
and U24057 (N_24057,N_23574,N_23280);
and U24058 (N_24058,N_22281,N_23139);
nand U24059 (N_24059,N_22167,N_22319);
nor U24060 (N_24060,N_23885,N_23001);
or U24061 (N_24061,N_22079,N_23312);
nand U24062 (N_24062,N_23707,N_22136);
nand U24063 (N_24063,N_23030,N_22180);
nor U24064 (N_24064,N_23521,N_23528);
and U24065 (N_24065,N_22454,N_23975);
nor U24066 (N_24066,N_22687,N_23206);
and U24067 (N_24067,N_22586,N_23503);
nand U24068 (N_24068,N_22461,N_23910);
nand U24069 (N_24069,N_23045,N_23190);
or U24070 (N_24070,N_22673,N_22653);
nand U24071 (N_24071,N_23679,N_23274);
or U24072 (N_24072,N_22854,N_23487);
nand U24073 (N_24073,N_23357,N_23824);
or U24074 (N_24074,N_23814,N_22980);
and U24075 (N_24075,N_23087,N_23802);
xor U24076 (N_24076,N_22999,N_22116);
or U24077 (N_24077,N_22173,N_23095);
nand U24078 (N_24078,N_23255,N_22739);
xor U24079 (N_24079,N_23075,N_23540);
and U24080 (N_24080,N_23207,N_23792);
or U24081 (N_24081,N_23310,N_23226);
or U24082 (N_24082,N_23931,N_23447);
and U24083 (N_24083,N_22514,N_23055);
or U24084 (N_24084,N_23929,N_22266);
nor U24085 (N_24085,N_22569,N_23498);
xor U24086 (N_24086,N_22480,N_22327);
xnor U24087 (N_24087,N_23519,N_23400);
xnor U24088 (N_24088,N_23094,N_22871);
nand U24089 (N_24089,N_23883,N_23683);
nand U24090 (N_24090,N_23556,N_23149);
nand U24091 (N_24091,N_22565,N_23586);
xnor U24092 (N_24092,N_22691,N_23548);
nor U24093 (N_24093,N_22450,N_22588);
nor U24094 (N_24094,N_23308,N_23838);
xnor U24095 (N_24095,N_23111,N_22609);
or U24096 (N_24096,N_22800,N_23983);
and U24097 (N_24097,N_22897,N_23874);
and U24098 (N_24098,N_22426,N_23164);
or U24099 (N_24099,N_22354,N_23151);
nand U24100 (N_24100,N_23711,N_22917);
nand U24101 (N_24101,N_22096,N_22486);
xor U24102 (N_24102,N_22335,N_22210);
nor U24103 (N_24103,N_23209,N_23834);
nor U24104 (N_24104,N_23432,N_22380);
and U24105 (N_24105,N_23279,N_23296);
nand U24106 (N_24106,N_22891,N_22975);
and U24107 (N_24107,N_22114,N_23685);
nor U24108 (N_24108,N_22365,N_22928);
xnor U24109 (N_24109,N_23057,N_22432);
or U24110 (N_24110,N_23973,N_23301);
nor U24111 (N_24111,N_23856,N_23861);
nand U24112 (N_24112,N_22017,N_23125);
and U24113 (N_24113,N_23364,N_22295);
xnor U24114 (N_24114,N_22492,N_22236);
and U24115 (N_24115,N_22259,N_23143);
xor U24116 (N_24116,N_22692,N_23851);
and U24117 (N_24117,N_23474,N_23407);
nand U24118 (N_24118,N_23618,N_22342);
nor U24119 (N_24119,N_23442,N_23924);
and U24120 (N_24120,N_22904,N_22242);
and U24121 (N_24121,N_22766,N_22881);
or U24122 (N_24122,N_23056,N_22746);
nor U24123 (N_24123,N_23131,N_23794);
nor U24124 (N_24124,N_22802,N_22183);
nor U24125 (N_24125,N_22248,N_23073);
nor U24126 (N_24126,N_23713,N_22665);
nor U24127 (N_24127,N_23675,N_22793);
xor U24128 (N_24128,N_22924,N_23452);
or U24129 (N_24129,N_22853,N_22467);
or U24130 (N_24130,N_22910,N_22069);
or U24131 (N_24131,N_23242,N_23163);
or U24132 (N_24132,N_22715,N_22389);
or U24133 (N_24133,N_22400,N_23642);
nor U24134 (N_24134,N_22166,N_23021);
nand U24135 (N_24135,N_23461,N_22995);
and U24136 (N_24136,N_22035,N_22320);
nor U24137 (N_24137,N_23522,N_22907);
or U24138 (N_24138,N_22876,N_22846);
or U24139 (N_24139,N_23342,N_22716);
xor U24140 (N_24140,N_22721,N_23705);
xor U24141 (N_24141,N_23661,N_23568);
nand U24142 (N_24142,N_23750,N_23646);
and U24143 (N_24143,N_23516,N_22919);
xor U24144 (N_24144,N_23557,N_23616);
and U24145 (N_24145,N_23146,N_22663);
nand U24146 (N_24146,N_22247,N_23463);
nand U24147 (N_24147,N_23024,N_22753);
or U24148 (N_24148,N_22632,N_23555);
xnor U24149 (N_24149,N_23283,N_23815);
nand U24150 (N_24150,N_22285,N_22869);
nor U24151 (N_24151,N_23352,N_23145);
or U24152 (N_24152,N_23598,N_23531);
xnor U24153 (N_24153,N_23903,N_22593);
and U24154 (N_24154,N_23112,N_23784);
nor U24155 (N_24155,N_22559,N_23901);
nor U24156 (N_24156,N_23657,N_22120);
or U24157 (N_24157,N_23478,N_23199);
xnor U24158 (N_24158,N_23168,N_23437);
nand U24159 (N_24159,N_23416,N_22656);
nand U24160 (N_24160,N_23169,N_23157);
or U24161 (N_24161,N_22381,N_22641);
nor U24162 (N_24162,N_23476,N_22666);
nor U24163 (N_24163,N_22398,N_22765);
or U24164 (N_24164,N_22277,N_22602);
and U24165 (N_24165,N_22226,N_23742);
and U24166 (N_24166,N_22914,N_22782);
xor U24167 (N_24167,N_22889,N_22951);
or U24168 (N_24168,N_22592,N_22707);
nor U24169 (N_24169,N_22425,N_23912);
nor U24170 (N_24170,N_22087,N_23253);
nor U24171 (N_24171,N_23917,N_23664);
nand U24172 (N_24172,N_22316,N_23434);
or U24173 (N_24173,N_23547,N_23197);
xor U24174 (N_24174,N_22482,N_23028);
nand U24175 (N_24175,N_23063,N_23272);
nand U24176 (N_24176,N_23099,N_22594);
xor U24177 (N_24177,N_22374,N_22900);
and U24178 (N_24178,N_23454,N_22192);
and U24179 (N_24179,N_22470,N_22159);
nand U24180 (N_24180,N_22612,N_22194);
xor U24181 (N_24181,N_23881,N_23541);
xor U24182 (N_24182,N_22263,N_22291);
xnor U24183 (N_24183,N_23699,N_22090);
and U24184 (N_24184,N_22735,N_23789);
and U24185 (N_24185,N_23409,N_22168);
nand U24186 (N_24186,N_22803,N_23827);
or U24187 (N_24187,N_22540,N_23697);
and U24188 (N_24188,N_23018,N_23295);
nand U24189 (N_24189,N_22410,N_23488);
nor U24190 (N_24190,N_22912,N_23093);
nand U24191 (N_24191,N_22045,N_22145);
nand U24192 (N_24192,N_23769,N_23061);
and U24193 (N_24193,N_23285,N_22784);
nor U24194 (N_24194,N_22464,N_22819);
nand U24195 (N_24195,N_23059,N_23037);
xor U24196 (N_24196,N_22104,N_22066);
or U24197 (N_24197,N_22574,N_23069);
nor U24198 (N_24198,N_22538,N_23167);
xor U24199 (N_24199,N_22761,N_23029);
nor U24200 (N_24200,N_22440,N_23041);
nor U24201 (N_24201,N_23777,N_23708);
nor U24202 (N_24202,N_23191,N_23264);
or U24203 (N_24203,N_23966,N_22187);
nor U24204 (N_24204,N_22658,N_23989);
and U24205 (N_24205,N_23311,N_23804);
or U24206 (N_24206,N_23104,N_22579);
or U24207 (N_24207,N_23902,N_23126);
nand U24208 (N_24208,N_22528,N_22393);
xor U24209 (N_24209,N_23821,N_23597);
or U24210 (N_24210,N_23876,N_23064);
xor U24211 (N_24211,N_22829,N_22982);
and U24212 (N_24212,N_22471,N_23982);
xnor U24213 (N_24213,N_22275,N_23443);
nor U24214 (N_24214,N_22206,N_23774);
and U24215 (N_24215,N_23819,N_23397);
nand U24216 (N_24216,N_23993,N_22190);
or U24217 (N_24217,N_23000,N_23512);
xnor U24218 (N_24218,N_23172,N_22345);
nor U24219 (N_24219,N_23241,N_23919);
nor U24220 (N_24220,N_22082,N_22644);
or U24221 (N_24221,N_23263,N_22227);
and U24222 (N_24222,N_22274,N_23863);
and U24223 (N_24223,N_23674,N_23778);
nor U24224 (N_24224,N_23309,N_22830);
nor U24225 (N_24225,N_23201,N_22969);
nand U24226 (N_24226,N_23402,N_23622);
nand U24227 (N_24227,N_22027,N_23106);
xor U24228 (N_24228,N_23549,N_22386);
and U24229 (N_24229,N_22585,N_22621);
and U24230 (N_24230,N_23445,N_22456);
nand U24231 (N_24231,N_22775,N_22430);
xnor U24232 (N_24232,N_22947,N_23992);
nor U24233 (N_24233,N_22616,N_23174);
or U24234 (N_24234,N_22519,N_23273);
nand U24235 (N_24235,N_22649,N_23590);
nor U24236 (N_24236,N_22028,N_23985);
nand U24237 (N_24237,N_22751,N_23974);
and U24238 (N_24238,N_22169,N_22521);
nand U24239 (N_24239,N_23765,N_22051);
or U24240 (N_24240,N_22010,N_22332);
xor U24241 (N_24241,N_22610,N_22029);
nor U24242 (N_24242,N_23517,N_22060);
or U24243 (N_24243,N_23886,N_22003);
or U24244 (N_24244,N_23897,N_22391);
nand U24245 (N_24245,N_23566,N_22534);
xor U24246 (N_24246,N_23007,N_22163);
xor U24247 (N_24247,N_22055,N_23998);
nand U24248 (N_24248,N_23004,N_22283);
xor U24249 (N_24249,N_23734,N_22061);
and U24250 (N_24250,N_22763,N_22182);
nand U24251 (N_24251,N_23219,N_22966);
and U24252 (N_24252,N_23298,N_22408);
or U24253 (N_24253,N_23757,N_22578);
xnor U24254 (N_24254,N_23529,N_22189);
xnor U24255 (N_24255,N_23150,N_23494);
nand U24256 (N_24256,N_22036,N_23714);
nand U24257 (N_24257,N_23072,N_22068);
xnor U24258 (N_24258,N_23722,N_22262);
or U24259 (N_24259,N_23505,N_23645);
nor U24260 (N_24260,N_23842,N_22209);
or U24261 (N_24261,N_23438,N_22600);
nor U24262 (N_24262,N_23136,N_23603);
or U24263 (N_24263,N_23185,N_23155);
or U24264 (N_24264,N_22501,N_22049);
nand U24265 (N_24265,N_23888,N_23160);
or U24266 (N_24266,N_23133,N_22895);
or U24267 (N_24267,N_23412,N_23335);
or U24268 (N_24268,N_23915,N_22706);
or U24269 (N_24269,N_22297,N_23455);
nand U24270 (N_24270,N_23943,N_22932);
nand U24271 (N_24271,N_22799,N_23620);
xnor U24272 (N_24272,N_22740,N_23508);
nand U24273 (N_24273,N_22328,N_23640);
nor U24274 (N_24274,N_23567,N_22271);
nor U24275 (N_24275,N_22734,N_23395);
nor U24276 (N_24276,N_23147,N_22360);
nor U24277 (N_24277,N_23823,N_22221);
nor U24278 (N_24278,N_23835,N_23132);
nand U24279 (N_24279,N_23062,N_22085);
and U24280 (N_24280,N_23944,N_22089);
or U24281 (N_24281,N_22418,N_22264);
or U24282 (N_24282,N_22640,N_23922);
and U24283 (N_24283,N_22823,N_23891);
nand U24284 (N_24284,N_23444,N_23570);
and U24285 (N_24285,N_23629,N_23080);
xor U24286 (N_24286,N_23847,N_23404);
nor U24287 (N_24287,N_23319,N_22124);
or U24288 (N_24288,N_23808,N_23798);
xor U24289 (N_24289,N_22630,N_23391);
nor U24290 (N_24290,N_22048,N_23953);
and U24291 (N_24291,N_23621,N_22896);
xnor U24292 (N_24292,N_22109,N_22902);
nor U24293 (N_24293,N_23336,N_23754);
and U24294 (N_24294,N_22222,N_23451);
or U24295 (N_24295,N_22535,N_23889);
or U24296 (N_24296,N_23228,N_23020);
or U24297 (N_24297,N_22395,N_22973);
nand U24298 (N_24298,N_22195,N_22898);
xnor U24299 (N_24299,N_23643,N_23949);
and U24300 (N_24300,N_23562,N_23392);
nand U24301 (N_24301,N_22280,N_23036);
or U24302 (N_24302,N_23384,N_22860);
nand U24303 (N_24303,N_23232,N_23102);
nor U24304 (N_24304,N_22708,N_23995);
nor U24305 (N_24305,N_23939,N_23745);
xnor U24306 (N_24306,N_23159,N_23698);
and U24307 (N_24307,N_23610,N_23702);
nor U24308 (N_24308,N_22694,N_22967);
xor U24309 (N_24309,N_23581,N_23042);
and U24310 (N_24310,N_22922,N_22032);
and U24311 (N_24311,N_22322,N_23739);
nand U24312 (N_24312,N_23857,N_22596);
nand U24313 (N_24313,N_22346,N_22628);
nand U24314 (N_24314,N_22546,N_23238);
or U24315 (N_24315,N_23513,N_23532);
or U24316 (N_24316,N_22774,N_23372);
nor U24317 (N_24317,N_22133,N_22243);
xor U24318 (N_24318,N_23783,N_22934);
xnor U24319 (N_24319,N_22479,N_22942);
or U24320 (N_24320,N_23079,N_22619);
xor U24321 (N_24321,N_22827,N_22305);
nor U24322 (N_24322,N_23458,N_23246);
or U24323 (N_24323,N_23179,N_23192);
nor U24324 (N_24324,N_22228,N_22552);
or U24325 (N_24325,N_22458,N_23085);
xnor U24326 (N_24326,N_22416,N_22901);
nand U24327 (N_24327,N_22230,N_22930);
and U24328 (N_24328,N_22121,N_23256);
nor U24329 (N_24329,N_22867,N_23208);
or U24330 (N_24330,N_23654,N_23920);
nor U24331 (N_24331,N_22008,N_23233);
xnor U24332 (N_24332,N_22125,N_22359);
xnor U24333 (N_24333,N_23429,N_23759);
nor U24334 (N_24334,N_22437,N_23636);
xor U24335 (N_24335,N_23457,N_22288);
nand U24336 (N_24336,N_22452,N_22870);
nor U24337 (N_24337,N_23221,N_22575);
nand U24338 (N_24338,N_22545,N_22181);
and U24339 (N_24339,N_23978,N_23909);
nand U24340 (N_24340,N_22598,N_23362);
xnor U24341 (N_24341,N_22996,N_23089);
nand U24342 (N_24342,N_23666,N_22377);
nand U24343 (N_24343,N_22567,N_22057);
or U24344 (N_24344,N_22836,N_22564);
nand U24345 (N_24345,N_22750,N_22353);
nand U24346 (N_24346,N_22518,N_23313);
nor U24347 (N_24347,N_23710,N_23958);
xnor U24348 (N_24348,N_23423,N_23282);
nand U24349 (N_24349,N_23040,N_23373);
xor U24350 (N_24350,N_23044,N_23930);
nand U24351 (N_24351,N_23656,N_22568);
nand U24352 (N_24352,N_23700,N_22561);
and U24353 (N_24353,N_23760,N_22812);
or U24354 (N_24354,N_23623,N_23252);
nand U24355 (N_24355,N_23230,N_23872);
and U24356 (N_24356,N_23011,N_22092);
or U24357 (N_24357,N_23606,N_22196);
nor U24358 (N_24358,N_23514,N_23895);
nor U24359 (N_24359,N_23398,N_22376);
and U24360 (N_24360,N_23977,N_23096);
nand U24361 (N_24361,N_23047,N_23422);
and U24362 (N_24362,N_23236,N_23459);
nand U24363 (N_24363,N_22358,N_22058);
xor U24364 (N_24364,N_22608,N_22815);
nand U24365 (N_24365,N_22674,N_23970);
and U24366 (N_24366,N_23709,N_22433);
nor U24367 (N_24367,N_23376,N_23287);
nand U24368 (N_24368,N_23748,N_22965);
and U24369 (N_24369,N_23859,N_23043);
xnor U24370 (N_24370,N_22558,N_22018);
xnor U24371 (N_24371,N_23492,N_22804);
xnor U24372 (N_24372,N_22798,N_22583);
or U24373 (N_24373,N_22094,N_22704);
nor U24374 (N_24374,N_23306,N_22968);
nor U24375 (N_24375,N_22931,N_23904);
nor U24376 (N_24376,N_23994,N_23187);
nor U24377 (N_24377,N_23186,N_22873);
and U24378 (N_24378,N_23177,N_23976);
or U24379 (N_24379,N_22841,N_22474);
or U24380 (N_24380,N_22979,N_22762);
xnor U24381 (N_24381,N_23617,N_23873);
and U24382 (N_24382,N_23936,N_23399);
nor U24383 (N_24383,N_22490,N_22427);
or U24384 (N_24384,N_22255,N_23641);
xor U24385 (N_24385,N_22727,N_22088);
nor U24386 (N_24386,N_23969,N_23611);
and U24387 (N_24387,N_22445,N_23563);
or U24388 (N_24388,N_22796,N_22789);
nor U24389 (N_24389,N_23942,N_22547);
xor U24390 (N_24390,N_22582,N_22807);
xor U24391 (N_24391,N_22184,N_23440);
nor U24392 (N_24392,N_23571,N_23317);
nand U24393 (N_24393,N_22864,N_23171);
xor U24394 (N_24394,N_22429,N_22256);
nand U24395 (N_24395,N_22019,N_23653);
and U24396 (N_24396,N_22677,N_22991);
nand U24397 (N_24397,N_23741,N_23552);
nor U24398 (N_24398,N_22507,N_22858);
and U24399 (N_24399,N_22053,N_22606);
nand U24400 (N_24400,N_23587,N_22152);
nand U24401 (N_24401,N_23984,N_22899);
or U24402 (N_24402,N_22394,N_22818);
xor U24403 (N_24403,N_23500,N_22941);
nand U24404 (N_24404,N_22517,N_23229);
nand U24405 (N_24405,N_23196,N_23776);
nor U24406 (N_24406,N_22964,N_22955);
nand U24407 (N_24407,N_23170,N_23963);
and U24408 (N_24408,N_22729,N_23880);
nor U24409 (N_24409,N_23659,N_23204);
nand U24410 (N_24410,N_23138,N_23905);
nor U24411 (N_24411,N_23465,N_23866);
or U24412 (N_24412,N_22300,N_23369);
or U24413 (N_24413,N_22080,N_23947);
or U24414 (N_24414,N_23052,N_23758);
nor U24415 (N_24415,N_23845,N_22333);
or U24416 (N_24416,N_23247,N_22397);
nor U24417 (N_24417,N_23428,N_22075);
and U24418 (N_24418,N_23202,N_23351);
nand U24419 (N_24419,N_22378,N_22741);
xnor U24420 (N_24420,N_23810,N_22343);
or U24421 (N_24421,N_23694,N_22496);
xnor U24422 (N_24422,N_23430,N_23359);
nor U24423 (N_24423,N_22537,N_23812);
and U24424 (N_24424,N_23875,N_22257);
and U24425 (N_24425,N_23123,N_23358);
xnor U24426 (N_24426,N_22161,N_23544);
and U24427 (N_24427,N_23934,N_22229);
or U24428 (N_24428,N_23354,N_23533);
xor U24429 (N_24429,N_23321,N_23182);
nand U24430 (N_24430,N_23250,N_23225);
nor U24431 (N_24431,N_22801,N_22856);
nand U24432 (N_24432,N_22805,N_23585);
xor U24433 (N_24433,N_23594,N_23584);
and U24434 (N_24434,N_23775,N_22056);
xor U24435 (N_24435,N_22218,N_23850);
nor U24436 (N_24436,N_23378,N_23829);
or U24437 (N_24437,N_22444,N_23871);
nand U24438 (N_24438,N_23050,N_22587);
and U24439 (N_24439,N_23740,N_22671);
and U24440 (N_24440,N_22617,N_23367);
nor U24441 (N_24441,N_23176,N_23141);
or U24442 (N_24442,N_22052,N_23738);
nor U24443 (N_24443,N_22773,N_22006);
nand U24444 (N_24444,N_23109,N_23331);
nor U24445 (N_24445,N_22007,N_22755);
nand U24446 (N_24446,N_22212,N_23009);
nor U24447 (N_24447,N_22334,N_23377);
or U24448 (N_24448,N_23054,N_23341);
and U24449 (N_24449,N_22011,N_22005);
and U24450 (N_24450,N_23092,N_23527);
and U24451 (N_24451,N_23945,N_23026);
or U24452 (N_24452,N_23771,N_22406);
or U24453 (N_24453,N_22613,N_22690);
and U24454 (N_24454,N_23216,N_22806);
or U24455 (N_24455,N_23806,N_23375);
or U24456 (N_24456,N_23781,N_23725);
nor U24457 (N_24457,N_22488,N_22315);
or U24458 (N_24458,N_22350,N_22178);
nor U24459 (N_24459,N_23879,N_22701);
and U24460 (N_24460,N_22920,N_22703);
and U24461 (N_24461,N_23220,N_23010);
or U24462 (N_24462,N_22764,N_22441);
or U24463 (N_24463,N_22883,N_22664);
and U24464 (N_24464,N_22711,N_23788);
and U24465 (N_24465,N_22667,N_23419);
or U24466 (N_24466,N_23667,N_22214);
and U24467 (N_24467,N_22893,N_23014);
nand U24468 (N_24468,N_22463,N_22832);
xnor U24469 (N_24469,N_22639,N_23628);
nor U24470 (N_24470,N_23270,N_22944);
and U24471 (N_24471,N_22555,N_22208);
and U24472 (N_24472,N_23148,N_22369);
and U24473 (N_24473,N_22787,N_23393);
xor U24474 (N_24474,N_22179,N_22652);
and U24475 (N_24475,N_23865,N_22287);
and U24476 (N_24476,N_23217,N_22820);
and U24477 (N_24477,N_23870,N_23962);
or U24478 (N_24478,N_23933,N_23837);
nor U24479 (N_24479,N_22270,N_22945);
xor U24480 (N_24480,N_22299,N_22984);
and U24481 (N_24481,N_23660,N_23908);
xnor U24482 (N_24482,N_22279,N_22730);
nand U24483 (N_24483,N_22099,N_23413);
and U24484 (N_24484,N_22713,N_22185);
nand U24485 (N_24485,N_22372,N_23153);
xor U24486 (N_24486,N_22754,N_22106);
nand U24487 (N_24487,N_22525,N_23003);
and U24488 (N_24488,N_23715,N_23224);
xnor U24489 (N_24489,N_23695,N_22137);
or U24490 (N_24490,N_22216,N_23913);
and U24491 (N_24491,N_23275,N_22795);
or U24492 (N_24492,N_22064,N_22105);
or U24493 (N_24493,N_22175,N_23979);
xor U24494 (N_24494,N_23923,N_23403);
and U24495 (N_24495,N_22199,N_22526);
nor U24496 (N_24496,N_22536,N_22842);
or U24497 (N_24497,N_22863,N_22067);
xnor U24498 (N_24498,N_22529,N_23107);
or U24499 (N_24499,N_23361,N_22158);
nand U24500 (N_24500,N_23205,N_23633);
or U24501 (N_24501,N_22384,N_22781);
nor U24502 (N_24502,N_22331,N_23718);
xor U24503 (N_24503,N_23595,N_22623);
and U24504 (N_24504,N_23086,N_23479);
nor U24505 (N_24505,N_23801,N_23350);
xor U24506 (N_24506,N_22102,N_22542);
or U24507 (N_24507,N_22577,N_22268);
nor U24508 (N_24508,N_22645,N_23832);
and U24509 (N_24509,N_22323,N_23634);
nand U24510 (N_24510,N_23997,N_22845);
and U24511 (N_24511,N_22510,N_22417);
nand U24512 (N_24512,N_23480,N_22307);
and U24513 (N_24513,N_23383,N_22809);
or U24514 (N_24514,N_22543,N_22043);
and U24515 (N_24515,N_23294,N_22246);
nor U24516 (N_24516,N_22531,N_23858);
nor U24517 (N_24517,N_22258,N_22071);
or U24518 (N_24518,N_22004,N_23878);
nor U24519 (N_24519,N_22714,N_22757);
and U24520 (N_24520,N_23243,N_23921);
xnor U24521 (N_24521,N_22878,N_23198);
or U24522 (N_24522,N_23178,N_22855);
and U24523 (N_24523,N_23462,N_22493);
nand U24524 (N_24524,N_22352,N_23388);
nand U24525 (N_24525,N_22367,N_23005);
or U24526 (N_24526,N_22252,N_23188);
and U24527 (N_24527,N_23791,N_22201);
and U24528 (N_24528,N_22118,N_22356);
nand U24529 (N_24529,N_23506,N_23729);
and U24530 (N_24530,N_22491,N_22992);
xnor U24531 (N_24531,N_22508,N_23410);
xnor U24532 (N_24532,N_22312,N_23716);
xor U24533 (N_24533,N_22962,N_23988);
nor U24534 (N_24534,N_22217,N_22780);
and U24535 (N_24535,N_22689,N_23387);
xnor U24536 (N_24536,N_23200,N_22117);
or U24537 (N_24537,N_23892,N_23818);
xnor U24538 (N_24538,N_22100,N_22308);
and U24539 (N_24539,N_23530,N_23577);
nand U24540 (N_24540,N_22046,N_23964);
nor U24541 (N_24541,N_23752,N_23955);
and U24542 (N_24542,N_23896,N_22407);
xnor U24543 (N_24543,N_23386,N_22413);
or U24544 (N_24544,N_23483,N_22563);
and U24545 (N_24545,N_22723,N_23248);
and U24546 (N_24546,N_22457,N_23670);
nor U24547 (N_24547,N_22970,N_22240);
xor U24548 (N_24548,N_22357,N_22756);
and U24549 (N_24549,N_23632,N_22160);
or U24550 (N_24550,N_22211,N_22177);
or U24551 (N_24551,N_22489,N_23100);
or U24552 (N_24552,N_23166,N_22669);
xnor U24553 (N_24553,N_22937,N_23360);
and U24554 (N_24554,N_22198,N_22509);
or U24555 (N_24555,N_22940,N_23763);
nor U24556 (N_24556,N_22157,N_23593);
nor U24557 (N_24557,N_23601,N_22553);
nand U24558 (N_24558,N_22993,N_23278);
and U24559 (N_24559,N_23749,N_22115);
xnor U24560 (N_24560,N_22810,N_23103);
xnor U24561 (N_24561,N_22560,N_22419);
xnor U24562 (N_24562,N_22143,N_22505);
or U24563 (N_24563,N_23848,N_22001);
xor U24564 (N_24564,N_23626,N_22235);
nand U24565 (N_24565,N_23604,N_22550);
and U24566 (N_24566,N_23405,N_22825);
or U24567 (N_24567,N_23124,N_22424);
and U24568 (N_24568,N_22478,N_22301);
xor U24569 (N_24569,N_22745,N_23382);
xnor U24570 (N_24570,N_22977,N_23495);
or U24571 (N_24571,N_23926,N_22717);
nand U24572 (N_24572,N_22379,N_23390);
nor U24573 (N_24573,N_23578,N_22821);
or U24574 (N_24574,N_22439,N_22859);
nand U24575 (N_24575,N_23453,N_22956);
and U24576 (N_24576,N_23292,N_23596);
and U24577 (N_24577,N_22385,N_23469);
or U24578 (N_24578,N_22146,N_23786);
or U24579 (N_24579,N_23304,N_23460);
nand U24580 (N_24580,N_22344,N_23662);
nand U24581 (N_24581,N_22998,N_22779);
and U24582 (N_24582,N_23189,N_22144);
or U24583 (N_24583,N_23510,N_22742);
or U24584 (N_24584,N_23678,N_22336);
nor U24585 (N_24585,N_22953,N_22072);
and U24586 (N_24586,N_23986,N_22111);
and U24587 (N_24587,N_23316,N_22548);
and U24588 (N_24588,N_23589,N_22434);
xnor U24589 (N_24589,N_23237,N_22453);
nor U24590 (N_24590,N_23446,N_22324);
xor U24591 (N_24591,N_22777,N_23751);
nand U24592 (N_24592,N_22562,N_22607);
or U24593 (N_24593,N_22831,N_22091);
xor U24594 (N_24594,N_23299,N_23862);
xor U24595 (N_24595,N_23340,N_23053);
and U24596 (N_24596,N_22081,N_23546);
nand U24597 (N_24597,N_22086,N_22544);
xor U24598 (N_24598,N_22792,N_23535);
or U24599 (N_24599,N_23033,N_23550);
xor U24600 (N_24600,N_22874,N_23433);
nand U24601 (N_24601,N_22498,N_22961);
nor U24602 (N_24602,N_22348,N_22292);
nor U24603 (N_24603,N_23673,N_23251);
and U24604 (N_24604,N_22465,N_23173);
and U24605 (N_24605,N_22329,N_23212);
and U24606 (N_24606,N_22948,N_23766);
or U24607 (N_24607,N_23952,N_22244);
and U24608 (N_24608,N_23129,N_23693);
nand U24609 (N_24609,N_22554,N_22338);
nor U24610 (N_24610,N_23613,N_22626);
xnor U24611 (N_24611,N_23864,N_22943);
nand U24612 (N_24612,N_22659,N_23082);
and U24613 (N_24613,N_23509,N_23265);
nand U24614 (N_24614,N_23401,N_22317);
nand U24615 (N_24615,N_22785,N_23677);
or U24616 (N_24616,N_22294,N_23687);
xor U24617 (N_24617,N_22718,N_22172);
nand U24618 (N_24618,N_23799,N_23262);
or U24619 (N_24619,N_22680,N_23140);
xor U24620 (N_24620,N_22204,N_23411);
xor U24621 (N_24621,N_23485,N_23091);
and U24622 (N_24622,N_22373,N_23254);
nor U24623 (N_24623,N_23743,N_23266);
and U24624 (N_24624,N_23614,N_23849);
and U24625 (N_24625,N_23293,N_23034);
nor U24626 (N_24626,N_22885,N_23303);
and U24627 (N_24627,N_22772,N_23240);
xor U24628 (N_24628,N_22026,N_22431);
and U24629 (N_24629,N_22404,N_22282);
nand U24630 (N_24630,N_23481,N_22850);
nand U24631 (N_24631,N_22880,N_22098);
and U24632 (N_24632,N_23900,N_23127);
or U24633 (N_24633,N_22523,N_22527);
xor U24634 (N_24634,N_23817,N_23882);
or U24635 (N_24635,N_22728,N_22783);
and U24636 (N_24636,N_23520,N_23841);
nor U24637 (N_24637,N_22078,N_22797);
nand U24638 (N_24638,N_22215,N_23569);
and U24639 (N_24639,N_23490,N_22390);
and U24640 (N_24640,N_22065,N_23625);
nor U24641 (N_24641,N_22399,N_23836);
nor U24642 (N_24642,N_22473,N_22581);
xnor U24643 (N_24643,N_22131,N_22848);
nor U24644 (N_24644,N_23701,N_22905);
xor U24645 (N_24645,N_23065,N_23008);
xor U24646 (N_24646,N_23222,N_23418);
or U24647 (N_24647,N_22813,N_23925);
xor U24648 (N_24648,N_22877,N_23048);
nor U24649 (N_24649,N_22513,N_22683);
xor U24650 (N_24650,N_22599,N_23753);
and U24651 (N_24651,N_22392,N_22650);
and U24652 (N_24652,N_22989,N_23049);
and U24653 (N_24653,N_22918,N_23639);
or U24654 (N_24654,N_22615,N_23068);
nand U24655 (N_24655,N_22293,N_22097);
nor U24656 (N_24656,N_23526,N_22732);
nor U24657 (N_24657,N_23561,N_22363);
and U24658 (N_24658,N_22449,N_23118);
nor U24659 (N_24659,N_22835,N_23860);
nand U24660 (N_24660,N_22241,N_23961);
and U24661 (N_24661,N_23472,N_23668);
and U24662 (N_24662,N_22156,N_23630);
and U24663 (N_24663,N_23648,N_22139);
and U24664 (N_24664,N_22110,N_23627);
nor U24665 (N_24665,N_23796,N_23475);
and U24666 (N_24666,N_22808,N_22459);
nand U24667 (N_24667,N_22814,N_22573);
and U24668 (N_24668,N_22362,N_22678);
xor U24669 (N_24669,N_23846,N_23426);
and U24670 (N_24670,N_22504,N_23496);
or U24671 (N_24671,N_22637,N_23015);
xnor U24672 (N_24672,N_22571,N_22511);
nor U24673 (N_24673,N_23869,N_22261);
nor U24674 (N_24674,N_23833,N_23213);
xor U24675 (N_24675,N_23504,N_22495);
and U24676 (N_24676,N_22254,N_22186);
or U24677 (N_24677,N_23558,N_22840);
and U24678 (N_24678,N_23258,N_23070);
xor U24679 (N_24679,N_23142,N_22884);
and U24680 (N_24680,N_22382,N_23414);
xor U24681 (N_24681,N_22811,N_23853);
and U24682 (N_24682,N_22927,N_23450);
and U24683 (N_24683,N_22475,N_22648);
nor U24684 (N_24684,N_23467,N_22054);
or U24685 (N_24685,N_23655,N_23764);
or U24686 (N_24686,N_23877,N_23971);
and U24687 (N_24687,N_23337,N_23560);
and U24688 (N_24688,N_23058,N_22443);
nand U24689 (N_24689,N_23719,N_22122);
and U24690 (N_24690,N_22462,N_23600);
and U24691 (N_24691,N_23746,N_23803);
and U24692 (N_24692,N_22484,N_23477);
xor U24693 (N_24693,N_22983,N_23637);
nand U24694 (N_24694,N_22128,N_22468);
nand U24695 (N_24695,N_22313,N_22760);
nand U24696 (N_24696,N_23380,N_23259);
xor U24697 (N_24697,N_22015,N_23502);
nor U24698 (N_24698,N_23038,N_22076);
or U24699 (N_24699,N_22584,N_22595);
and U24700 (N_24700,N_23884,N_23473);
or U24701 (N_24701,N_23957,N_22769);
or U24702 (N_24702,N_22129,N_22661);
nor U24703 (N_24703,N_22047,N_23762);
or U24704 (N_24704,N_23355,N_22415);
nor U24705 (N_24705,N_23470,N_23647);
nand U24706 (N_24706,N_22232,N_22153);
xnor U24707 (N_24707,N_23793,N_22530);
or U24708 (N_24708,N_23195,N_22174);
nor U24709 (N_24709,N_23348,N_22865);
xnor U24710 (N_24710,N_23035,N_22736);
or U24711 (N_24711,N_23830,N_23019);
xor U24712 (N_24712,N_23334,N_22682);
xor U24713 (N_24713,N_22401,N_23731);
or U24714 (N_24714,N_22239,N_22093);
nand U24715 (N_24715,N_23649,N_22635);
nor U24716 (N_24716,N_23346,N_22532);
nor U24717 (N_24717,N_22705,N_22733);
or U24718 (N_24718,N_23016,N_22123);
or U24719 (N_24719,N_23768,N_22950);
xnor U24720 (N_24720,N_23175,N_23511);
nor U24721 (N_24721,N_23867,N_22771);
or U24722 (N_24722,N_23854,N_23307);
and U24723 (N_24723,N_22188,N_22958);
nand U24724 (N_24724,N_23223,N_23396);
nand U24725 (N_24725,N_22073,N_23394);
and U24726 (N_24726,N_23565,N_23417);
nand U24727 (N_24727,N_23928,N_23932);
or U24728 (N_24728,N_22002,N_22994);
xnor U24729 (N_24729,N_22290,N_23987);
xnor U24730 (N_24730,N_23572,N_23315);
or U24731 (N_24731,N_23305,N_23244);
xor U24732 (N_24732,N_23724,N_22633);
nor U24733 (N_24733,N_22908,N_22421);
xnor U24734 (N_24734,N_23156,N_22888);
xor U24735 (N_24735,N_22833,N_22963);
nand U24736 (N_24736,N_22298,N_23427);
nand U24737 (N_24737,N_23898,N_23980);
xor U24738 (N_24738,N_22063,N_23755);
nand U24739 (N_24739,N_22126,N_22886);
and U24740 (N_24740,N_22719,N_22791);
xor U24741 (N_24741,N_22314,N_23322);
and U24742 (N_24742,N_23680,N_22487);
nand U24743 (N_24743,N_23090,N_22024);
or U24744 (N_24744,N_22636,N_22725);
xnor U24745 (N_24745,N_23468,N_23894);
nor U24746 (N_24746,N_22890,N_23608);
and U24747 (N_24747,N_23619,N_22824);
nor U24748 (N_24748,N_22589,N_23493);
nand U24749 (N_24749,N_23899,N_22909);
nand U24750 (N_24750,N_22233,N_23773);
xor U24751 (N_24751,N_22147,N_22494);
nor U24752 (N_24752,N_23152,N_22025);
nand U24753 (N_24753,N_23579,N_23039);
xor U24754 (N_24754,N_23211,N_22077);
and U24755 (N_24755,N_23536,N_22709);
and U24756 (N_24756,N_22412,N_23449);
xor U24757 (N_24757,N_23767,N_23023);
xnor U24758 (N_24758,N_22119,N_23431);
and U24759 (N_24759,N_23074,N_22921);
nor U24760 (N_24760,N_22219,N_23366);
nor U24761 (N_24761,N_22698,N_22935);
and U24762 (N_24762,N_22768,N_22276);
xnor U24763 (N_24763,N_23852,N_23573);
nor U24764 (N_24764,N_22141,N_22722);
nand U24765 (N_24765,N_22084,N_22310);
nand U24766 (N_24766,N_22107,N_22170);
nand U24767 (N_24767,N_23733,N_22355);
or U24768 (N_24768,N_23612,N_23193);
nor U24769 (N_24769,N_23120,N_23855);
and U24770 (N_24770,N_22500,N_22759);
and U24771 (N_24771,N_23330,N_23785);
nand U24772 (N_24772,N_22155,N_23239);
and U24773 (N_24773,N_22981,N_22388);
xnor U24774 (N_24774,N_22828,N_23184);
xor U24775 (N_24775,N_22364,N_22148);
xor U24776 (N_24776,N_22485,N_22265);
or U24777 (N_24777,N_23543,N_22436);
and U24778 (N_24778,N_22949,N_22566);
nand U24779 (N_24779,N_23231,N_22447);
xor U24780 (N_24780,N_22455,N_23721);
and U24781 (N_24781,N_23644,N_23772);
and U24782 (N_24782,N_22770,N_23820);
and U24783 (N_24783,N_23890,N_22668);
xnor U24784 (N_24784,N_23605,N_23286);
nor U24785 (N_24785,N_22601,N_22403);
nor U24786 (N_24786,N_22611,N_22684);
nand U24787 (N_24787,N_22976,N_23084);
or U24788 (N_24788,N_23105,N_22516);
xor U24789 (N_24789,N_22330,N_23635);
or U24790 (N_24790,N_22326,N_22936);
nand U24791 (N_24791,N_22162,N_22681);
nor U24792 (N_24792,N_22438,N_23911);
nor U24793 (N_24793,N_22016,N_22985);
xor U24794 (N_24794,N_23276,N_23466);
nor U24795 (N_24795,N_22340,N_22794);
and U24796 (N_24796,N_23327,N_23651);
xnor U24797 (N_24797,N_22879,N_22978);
nor U24798 (N_24798,N_22557,N_22030);
nand U24799 (N_24799,N_22409,N_23113);
nand U24800 (N_24800,N_23194,N_23583);
nand U24801 (N_24801,N_22238,N_22710);
xor U24802 (N_24802,N_22197,N_22012);
or U24803 (N_24803,N_22213,N_23756);
or U24804 (N_24804,N_22245,N_23368);
nand U24805 (N_24805,N_22923,N_23732);
or U24806 (N_24806,N_23329,N_23813);
nor U24807 (N_24807,N_22039,N_22414);
or U24808 (N_24808,N_22150,N_22289);
xor U24809 (N_24809,N_23215,N_22894);
nor U24810 (N_24810,N_23385,N_22988);
and U24811 (N_24811,N_22834,N_23347);
nand U24812 (N_24812,N_22368,N_23831);
xor U24813 (N_24813,N_22127,N_23325);
nor U24814 (N_24814,N_22946,N_22164);
nand U24815 (N_24815,N_23937,N_22371);
nor U24816 (N_24816,N_23779,N_23797);
nand U24817 (N_24817,N_23704,N_22676);
nand U24818 (N_24818,N_23744,N_22466);
nor U24819 (N_24819,N_22349,N_22752);
xnor U24820 (N_24820,N_22070,N_23101);
xnor U24821 (N_24821,N_23013,N_22135);
xor U24822 (N_24822,N_23650,N_23599);
nand U24823 (N_24823,N_22038,N_23314);
or U24824 (N_24824,N_22685,N_23663);
and U24825 (N_24825,N_23281,N_23843);
nand U24826 (N_24826,N_22686,N_23374);
or U24827 (N_24827,N_22875,N_22700);
nor U24828 (N_24828,N_23356,N_22442);
nor U24829 (N_24829,N_22549,N_23290);
nand U24830 (N_24830,N_22370,N_23723);
or U24831 (N_24831,N_23538,N_23968);
or U24832 (N_24832,N_23203,N_22411);
and U24833 (N_24833,N_23002,N_23249);
nor U24834 (N_24834,N_22095,N_23515);
and U24835 (N_24835,N_22837,N_23727);
nor U24836 (N_24836,N_23017,N_22520);
or U24837 (N_24837,N_23682,N_22375);
xor U24838 (N_24838,N_22112,N_22631);
xnor U24839 (N_24839,N_23720,N_22225);
nor U24840 (N_24840,N_23991,N_23728);
or U24841 (N_24841,N_22556,N_23805);
nor U24842 (N_24842,N_23435,N_23245);
nand U24843 (N_24843,N_22031,N_22651);
and U24844 (N_24844,N_23415,N_22205);
nor U24845 (N_24845,N_22972,N_22062);
or U24846 (N_24846,N_22816,N_23525);
xor U24847 (N_24847,N_23706,N_23420);
and U24848 (N_24848,N_22670,N_22108);
nor U24849 (N_24849,N_22339,N_22023);
and U24850 (N_24850,N_22435,N_23381);
and U24851 (N_24851,N_22200,N_23615);
xor U24852 (N_24852,N_22624,N_23981);
nor U24853 (N_24853,N_22273,N_22013);
or U24854 (N_24854,N_22477,N_22448);
nor U24855 (N_24855,N_22672,N_23676);
or U24856 (N_24856,N_23115,N_22272);
or U24857 (N_24857,N_23956,N_22657);
and U24858 (N_24858,N_22034,N_23078);
nor U24859 (N_24859,N_23051,N_23951);
or U24860 (N_24860,N_23343,N_22990);
or U24861 (N_24861,N_23371,N_23349);
xor U24862 (N_24862,N_23291,N_23689);
or U24863 (N_24863,N_22906,N_23379);
xnor U24864 (N_24864,N_23914,N_23800);
nor U24865 (N_24865,N_23227,N_22939);
nor U24866 (N_24866,N_22149,N_22191);
and U24867 (N_24867,N_23032,N_22882);
xor U24868 (N_24868,N_23098,N_23916);
xnor U24869 (N_24869,N_22234,N_23439);
and U24870 (N_24870,N_23345,N_23006);
and U24871 (N_24871,N_22724,N_22021);
and U24872 (N_24872,N_23534,N_23624);
or U24873 (N_24873,N_23108,N_23559);
nor U24874 (N_24874,N_22341,N_22849);
xnor U24875 (N_24875,N_23747,N_23840);
xor U24876 (N_24876,N_23959,N_22347);
nand U24877 (N_24877,N_23665,N_22580);
or U24878 (N_24878,N_23128,N_23761);
nand U24879 (N_24879,N_22042,N_23288);
or U24880 (N_24880,N_23060,N_23353);
or U24881 (N_24881,N_23114,N_22913);
or U24882 (N_24882,N_23972,N_23134);
nor U24883 (N_24883,N_23690,N_22675);
xor U24884 (N_24884,N_23116,N_22351);
nand U24885 (N_24885,N_22605,N_23893);
or U24886 (N_24886,N_22887,N_23284);
xor U24887 (N_24887,N_22541,N_23688);
and U24888 (N_24888,N_23012,N_23297);
and U24889 (N_24889,N_23609,N_23370);
nand U24890 (N_24890,N_23081,N_22396);
or U24891 (N_24891,N_22986,N_22460);
nor U24892 (N_24892,N_22260,N_22304);
nor U24893 (N_24893,N_22269,N_23489);
xor U24894 (N_24894,N_23318,N_22132);
nand U24895 (N_24895,N_23161,N_22318);
or U24896 (N_24896,N_23130,N_23214);
xor U24897 (N_24897,N_22361,N_23464);
and U24898 (N_24898,N_23839,N_23162);
nand U24899 (N_24899,N_22224,N_23537);
nor U24900 (N_24900,N_22165,N_23471);
and U24901 (N_24901,N_22857,N_22851);
xnor U24902 (N_24902,N_23807,N_23486);
xnor U24903 (N_24903,N_23591,N_23365);
xnor U24904 (N_24904,N_22512,N_22590);
and U24905 (N_24905,N_23607,N_22524);
nand U24906 (N_24906,N_22286,N_23448);
nand U24907 (N_24907,N_22647,N_23083);
xor U24908 (N_24908,N_23825,N_23602);
or U24909 (N_24909,N_22638,N_22697);
and U24910 (N_24910,N_23696,N_23031);
xor U24911 (N_24911,N_22852,N_23681);
nand U24912 (N_24912,N_23234,N_22151);
nor U24913 (N_24913,N_22506,N_23553);
xnor U24914 (N_24914,N_22957,N_23703);
xor U24915 (N_24915,N_23339,N_22778);
or U24916 (N_24916,N_22387,N_22952);
and U24917 (N_24917,N_23967,N_22737);
nand U24918 (N_24918,N_22037,N_23684);
nand U24919 (N_24919,N_23990,N_22551);
nor U24920 (N_24920,N_23261,N_22603);
nor U24921 (N_24921,N_23121,N_22693);
xor U24922 (N_24922,N_23137,N_23165);
and U24923 (N_24923,N_23576,N_22695);
and U24924 (N_24924,N_22748,N_23267);
nand U24925 (N_24925,N_22916,N_23066);
nor U24926 (N_24926,N_22014,N_23671);
or U24927 (N_24927,N_22422,N_23269);
xor U24928 (N_24928,N_22142,N_23077);
or U24929 (N_24929,N_23551,N_23271);
and U24930 (N_24930,N_23097,N_23631);
or U24931 (N_24931,N_23686,N_22767);
nand U24932 (N_24932,N_23652,N_23158);
nor U24933 (N_24933,N_22130,N_22383);
nor U24934 (N_24934,N_23638,N_22959);
nand U24935 (N_24935,N_22176,N_22925);
and U24936 (N_24936,N_22325,N_22428);
xnor U24937 (N_24937,N_22758,N_22911);
or U24938 (N_24938,N_23960,N_23497);
and U24939 (N_24939,N_22929,N_23183);
nor U24940 (N_24940,N_23948,N_22420);
or U24941 (N_24941,N_22892,N_22044);
and U24942 (N_24942,N_23726,N_22688);
xnor U24943 (N_24943,N_22337,N_22503);
nor U24944 (N_24944,N_22591,N_22253);
nand U24945 (N_24945,N_23328,N_22113);
and U24946 (N_24946,N_23181,N_22472);
and U24947 (N_24947,N_22321,N_23524);
or U24948 (N_24948,N_22251,N_23441);
xnor U24949 (N_24949,N_22533,N_23927);
and U24950 (N_24950,N_22655,N_23144);
xor U24951 (N_24951,N_23737,N_23122);
nor U24952 (N_24952,N_22576,N_23950);
xor U24953 (N_24953,N_22469,N_23406);
nor U24954 (N_24954,N_22960,N_22987);
or U24955 (N_24955,N_22284,N_22515);
or U24956 (N_24956,N_22101,N_23300);
nor U24957 (N_24957,N_22614,N_23389);
nor U24958 (N_24958,N_22154,N_22303);
xor U24959 (N_24959,N_22237,N_23027);
or U24960 (N_24960,N_23717,N_23588);
xor U24961 (N_24961,N_23235,N_22050);
nand U24962 (N_24962,N_23996,N_22702);
and U24963 (N_24963,N_23408,N_22103);
xor U24964 (N_24964,N_22074,N_22776);
nor U24965 (N_24965,N_23965,N_22223);
nand U24966 (N_24966,N_22627,N_22597);
nor U24967 (N_24967,N_23154,N_22738);
and U24968 (N_24968,N_23491,N_23067);
and U24969 (N_24969,N_23507,N_22311);
nand U24970 (N_24970,N_22838,N_23046);
or U24971 (N_24971,N_23826,N_22309);
or U24972 (N_24972,N_22249,N_22933);
or U24973 (N_24973,N_23935,N_23180);
and U24974 (N_24974,N_23691,N_22622);
or U24975 (N_24975,N_22826,N_23592);
or U24976 (N_24976,N_23324,N_23780);
xor U24977 (N_24977,N_22033,N_23770);
and U24978 (N_24978,N_22278,N_22302);
xnor U24979 (N_24979,N_22231,N_23260);
and U24980 (N_24980,N_22618,N_22138);
nor U24981 (N_24981,N_23484,N_23436);
nand U24982 (N_24982,N_23425,N_22022);
nor U24983 (N_24983,N_23135,N_22861);
xor U24984 (N_24984,N_23809,N_22971);
and U24985 (N_24985,N_23844,N_22643);
and U24986 (N_24986,N_23790,N_22743);
nor U24987 (N_24987,N_22642,N_23887);
nand U24988 (N_24988,N_22140,N_22134);
nor U24989 (N_24989,N_22423,N_22974);
xnor U24990 (N_24990,N_22009,N_22499);
xor U24991 (N_24991,N_23268,N_22497);
nor U24992 (N_24992,N_23575,N_23277);
or U24993 (N_24993,N_23658,N_22522);
nor U24994 (N_24994,N_22862,N_23946);
or U24995 (N_24995,N_23210,N_22662);
nand U24996 (N_24996,N_23289,N_22749);
nand U24997 (N_24997,N_22539,N_22483);
and U24998 (N_24998,N_23828,N_23071);
or U24999 (N_24999,N_23332,N_23456);
xnor U25000 (N_25000,N_23352,N_22232);
and U25001 (N_25001,N_23418,N_22242);
or U25002 (N_25002,N_23293,N_23862);
nor U25003 (N_25003,N_22684,N_22159);
nor U25004 (N_25004,N_23021,N_23541);
and U25005 (N_25005,N_23064,N_22314);
and U25006 (N_25006,N_22763,N_22999);
nor U25007 (N_25007,N_23746,N_22051);
nand U25008 (N_25008,N_22676,N_23215);
xnor U25009 (N_25009,N_22452,N_23325);
nand U25010 (N_25010,N_22031,N_22823);
xor U25011 (N_25011,N_23147,N_23355);
xnor U25012 (N_25012,N_23609,N_23512);
xor U25013 (N_25013,N_22698,N_23266);
xor U25014 (N_25014,N_23946,N_23968);
nor U25015 (N_25015,N_23329,N_23398);
xor U25016 (N_25016,N_23699,N_22719);
xnor U25017 (N_25017,N_23762,N_22886);
nand U25018 (N_25018,N_22142,N_22876);
xor U25019 (N_25019,N_22730,N_23025);
xnor U25020 (N_25020,N_23235,N_22573);
nand U25021 (N_25021,N_22007,N_23925);
and U25022 (N_25022,N_23933,N_23684);
xnor U25023 (N_25023,N_23948,N_23565);
or U25024 (N_25024,N_23995,N_23963);
or U25025 (N_25025,N_23698,N_22675);
and U25026 (N_25026,N_23415,N_23987);
and U25027 (N_25027,N_23123,N_22499);
or U25028 (N_25028,N_22309,N_22843);
xor U25029 (N_25029,N_22022,N_23178);
and U25030 (N_25030,N_23627,N_22687);
nor U25031 (N_25031,N_23146,N_23377);
nor U25032 (N_25032,N_23376,N_22070);
or U25033 (N_25033,N_22277,N_23076);
xnor U25034 (N_25034,N_22644,N_23277);
nor U25035 (N_25035,N_23611,N_23865);
or U25036 (N_25036,N_22873,N_22368);
and U25037 (N_25037,N_23745,N_22365);
and U25038 (N_25038,N_23414,N_22753);
nand U25039 (N_25039,N_22613,N_22299);
nor U25040 (N_25040,N_23748,N_23269);
and U25041 (N_25041,N_23915,N_23430);
xor U25042 (N_25042,N_23892,N_22593);
or U25043 (N_25043,N_23567,N_22070);
and U25044 (N_25044,N_23013,N_22923);
nor U25045 (N_25045,N_23290,N_23954);
xnor U25046 (N_25046,N_23382,N_22859);
nand U25047 (N_25047,N_22340,N_23104);
or U25048 (N_25048,N_22887,N_23798);
xor U25049 (N_25049,N_23637,N_22119);
or U25050 (N_25050,N_23910,N_23841);
nand U25051 (N_25051,N_23156,N_22223);
and U25052 (N_25052,N_22910,N_22797);
or U25053 (N_25053,N_23411,N_23852);
or U25054 (N_25054,N_22075,N_23315);
xnor U25055 (N_25055,N_23077,N_23401);
nand U25056 (N_25056,N_23084,N_22382);
nand U25057 (N_25057,N_23879,N_23308);
or U25058 (N_25058,N_22988,N_23519);
xnor U25059 (N_25059,N_23005,N_22280);
nand U25060 (N_25060,N_23397,N_23389);
nand U25061 (N_25061,N_22064,N_23789);
and U25062 (N_25062,N_22377,N_23249);
nand U25063 (N_25063,N_23744,N_23032);
and U25064 (N_25064,N_23376,N_22321);
xnor U25065 (N_25065,N_23481,N_22625);
xnor U25066 (N_25066,N_22581,N_23729);
or U25067 (N_25067,N_23877,N_22215);
or U25068 (N_25068,N_23756,N_23900);
xor U25069 (N_25069,N_22684,N_23976);
and U25070 (N_25070,N_22023,N_22244);
nor U25071 (N_25071,N_23353,N_22816);
nand U25072 (N_25072,N_22781,N_23594);
or U25073 (N_25073,N_22857,N_23077);
nor U25074 (N_25074,N_22975,N_22608);
nand U25075 (N_25075,N_23665,N_22940);
or U25076 (N_25076,N_23845,N_22177);
nor U25077 (N_25077,N_23634,N_23199);
or U25078 (N_25078,N_23569,N_23036);
nand U25079 (N_25079,N_23264,N_23948);
xor U25080 (N_25080,N_23115,N_23306);
and U25081 (N_25081,N_23830,N_23795);
nand U25082 (N_25082,N_22036,N_22129);
xor U25083 (N_25083,N_23314,N_23376);
or U25084 (N_25084,N_23259,N_22701);
xnor U25085 (N_25085,N_23106,N_23740);
nand U25086 (N_25086,N_22645,N_22417);
or U25087 (N_25087,N_22451,N_23906);
xor U25088 (N_25088,N_23668,N_22412);
nand U25089 (N_25089,N_22537,N_22400);
or U25090 (N_25090,N_23888,N_22011);
nand U25091 (N_25091,N_22116,N_23374);
or U25092 (N_25092,N_22192,N_23853);
xor U25093 (N_25093,N_22959,N_23679);
xnor U25094 (N_25094,N_22565,N_23963);
xor U25095 (N_25095,N_23438,N_22321);
and U25096 (N_25096,N_23207,N_22857);
or U25097 (N_25097,N_22192,N_22418);
xor U25098 (N_25098,N_23842,N_23782);
or U25099 (N_25099,N_23394,N_23160);
nand U25100 (N_25100,N_23467,N_23700);
xor U25101 (N_25101,N_23680,N_22814);
xor U25102 (N_25102,N_23326,N_23431);
xnor U25103 (N_25103,N_22210,N_23623);
nor U25104 (N_25104,N_23678,N_23021);
and U25105 (N_25105,N_23318,N_23432);
xor U25106 (N_25106,N_23884,N_23753);
nand U25107 (N_25107,N_23458,N_23302);
and U25108 (N_25108,N_23434,N_22119);
nor U25109 (N_25109,N_22733,N_23240);
and U25110 (N_25110,N_23832,N_23039);
and U25111 (N_25111,N_22766,N_22682);
xnor U25112 (N_25112,N_22065,N_23656);
nor U25113 (N_25113,N_22647,N_22813);
nand U25114 (N_25114,N_22207,N_22903);
or U25115 (N_25115,N_22641,N_23921);
nor U25116 (N_25116,N_23034,N_22739);
xor U25117 (N_25117,N_22147,N_23864);
or U25118 (N_25118,N_22537,N_22117);
nand U25119 (N_25119,N_22698,N_23170);
xnor U25120 (N_25120,N_22033,N_22126);
nand U25121 (N_25121,N_22028,N_22960);
nor U25122 (N_25122,N_23071,N_22488);
and U25123 (N_25123,N_23582,N_22385);
or U25124 (N_25124,N_23618,N_22899);
xor U25125 (N_25125,N_22096,N_22193);
nand U25126 (N_25126,N_23491,N_23502);
or U25127 (N_25127,N_22352,N_22156);
nor U25128 (N_25128,N_22078,N_23651);
or U25129 (N_25129,N_23476,N_23330);
or U25130 (N_25130,N_22118,N_22802);
nand U25131 (N_25131,N_22348,N_23434);
xnor U25132 (N_25132,N_22783,N_22913);
or U25133 (N_25133,N_23616,N_22049);
xnor U25134 (N_25134,N_22328,N_23955);
and U25135 (N_25135,N_23029,N_22077);
nor U25136 (N_25136,N_23738,N_22366);
nand U25137 (N_25137,N_23655,N_23766);
xor U25138 (N_25138,N_23205,N_23439);
nand U25139 (N_25139,N_23089,N_23271);
and U25140 (N_25140,N_23039,N_22760);
xor U25141 (N_25141,N_22916,N_22314);
xnor U25142 (N_25142,N_23513,N_23249);
and U25143 (N_25143,N_22863,N_23537);
nand U25144 (N_25144,N_23879,N_22554);
xnor U25145 (N_25145,N_23377,N_23106);
nand U25146 (N_25146,N_22538,N_22696);
or U25147 (N_25147,N_23182,N_23492);
nor U25148 (N_25148,N_23212,N_22534);
and U25149 (N_25149,N_23929,N_22844);
xor U25150 (N_25150,N_22459,N_23841);
nor U25151 (N_25151,N_23826,N_22445);
or U25152 (N_25152,N_22124,N_22830);
nor U25153 (N_25153,N_22383,N_23653);
or U25154 (N_25154,N_22540,N_22578);
nand U25155 (N_25155,N_22724,N_23966);
xnor U25156 (N_25156,N_23750,N_23021);
xor U25157 (N_25157,N_22476,N_22358);
xnor U25158 (N_25158,N_23240,N_23309);
or U25159 (N_25159,N_22661,N_23647);
or U25160 (N_25160,N_23418,N_23378);
nor U25161 (N_25161,N_23839,N_22932);
xor U25162 (N_25162,N_22424,N_22737);
and U25163 (N_25163,N_23463,N_22451);
nand U25164 (N_25164,N_22691,N_23751);
or U25165 (N_25165,N_23373,N_22125);
or U25166 (N_25166,N_22492,N_22239);
and U25167 (N_25167,N_23840,N_23963);
or U25168 (N_25168,N_23585,N_23935);
and U25169 (N_25169,N_23845,N_22794);
xnor U25170 (N_25170,N_22993,N_23934);
nor U25171 (N_25171,N_22363,N_23844);
and U25172 (N_25172,N_22445,N_22636);
or U25173 (N_25173,N_22349,N_22785);
and U25174 (N_25174,N_23244,N_23444);
nor U25175 (N_25175,N_23975,N_22976);
or U25176 (N_25176,N_23291,N_23094);
nand U25177 (N_25177,N_23480,N_22626);
or U25178 (N_25178,N_22893,N_22046);
xnor U25179 (N_25179,N_22430,N_22950);
or U25180 (N_25180,N_23986,N_23101);
or U25181 (N_25181,N_22802,N_23591);
and U25182 (N_25182,N_23354,N_22262);
and U25183 (N_25183,N_22657,N_23716);
nand U25184 (N_25184,N_23915,N_23280);
xnor U25185 (N_25185,N_22996,N_22721);
nand U25186 (N_25186,N_23088,N_22387);
and U25187 (N_25187,N_23849,N_22079);
or U25188 (N_25188,N_23551,N_22341);
or U25189 (N_25189,N_23263,N_22622);
nand U25190 (N_25190,N_23243,N_23738);
xnor U25191 (N_25191,N_22348,N_22102);
nand U25192 (N_25192,N_22440,N_23630);
xor U25193 (N_25193,N_23459,N_23783);
nand U25194 (N_25194,N_22125,N_22748);
or U25195 (N_25195,N_22954,N_22337);
xnor U25196 (N_25196,N_23460,N_23333);
nor U25197 (N_25197,N_22757,N_23556);
xnor U25198 (N_25198,N_22513,N_23655);
xor U25199 (N_25199,N_22228,N_23006);
nor U25200 (N_25200,N_23033,N_22660);
and U25201 (N_25201,N_23396,N_22480);
and U25202 (N_25202,N_23854,N_23630);
xor U25203 (N_25203,N_23167,N_23153);
and U25204 (N_25204,N_23103,N_22111);
nor U25205 (N_25205,N_23659,N_23775);
xor U25206 (N_25206,N_22717,N_23827);
xnor U25207 (N_25207,N_23518,N_23826);
nor U25208 (N_25208,N_23897,N_23816);
nand U25209 (N_25209,N_23192,N_22414);
xor U25210 (N_25210,N_22275,N_22833);
xor U25211 (N_25211,N_22102,N_22689);
nor U25212 (N_25212,N_23140,N_22578);
xor U25213 (N_25213,N_22079,N_22231);
nand U25214 (N_25214,N_22868,N_22296);
nand U25215 (N_25215,N_23703,N_23054);
nor U25216 (N_25216,N_22038,N_23968);
xor U25217 (N_25217,N_23759,N_23823);
nand U25218 (N_25218,N_22849,N_23991);
xnor U25219 (N_25219,N_23783,N_23182);
nand U25220 (N_25220,N_22163,N_22224);
xnor U25221 (N_25221,N_23775,N_22752);
and U25222 (N_25222,N_23801,N_23583);
nor U25223 (N_25223,N_22062,N_22549);
nand U25224 (N_25224,N_23551,N_23288);
nand U25225 (N_25225,N_23217,N_23059);
nor U25226 (N_25226,N_23130,N_22655);
nand U25227 (N_25227,N_23353,N_23703);
nor U25228 (N_25228,N_22778,N_22253);
nor U25229 (N_25229,N_22460,N_23146);
nor U25230 (N_25230,N_22593,N_22564);
nor U25231 (N_25231,N_23835,N_23872);
xor U25232 (N_25232,N_22032,N_23865);
and U25233 (N_25233,N_23290,N_22176);
nor U25234 (N_25234,N_22418,N_23277);
and U25235 (N_25235,N_22764,N_22840);
and U25236 (N_25236,N_22197,N_23354);
nand U25237 (N_25237,N_23178,N_23514);
nor U25238 (N_25238,N_23550,N_23173);
and U25239 (N_25239,N_23543,N_22424);
or U25240 (N_25240,N_22461,N_23671);
nand U25241 (N_25241,N_22033,N_23338);
xor U25242 (N_25242,N_23399,N_22730);
nand U25243 (N_25243,N_23344,N_22484);
or U25244 (N_25244,N_23389,N_22425);
nand U25245 (N_25245,N_22152,N_23868);
nand U25246 (N_25246,N_23518,N_22411);
and U25247 (N_25247,N_22155,N_22159);
or U25248 (N_25248,N_22654,N_23211);
nand U25249 (N_25249,N_23890,N_23432);
or U25250 (N_25250,N_22701,N_23586);
nor U25251 (N_25251,N_23691,N_22280);
and U25252 (N_25252,N_22842,N_23599);
nand U25253 (N_25253,N_23721,N_22319);
and U25254 (N_25254,N_22235,N_22170);
xnor U25255 (N_25255,N_23679,N_22366);
and U25256 (N_25256,N_23899,N_23255);
or U25257 (N_25257,N_23266,N_22593);
nand U25258 (N_25258,N_23420,N_22094);
and U25259 (N_25259,N_22903,N_23284);
nor U25260 (N_25260,N_22896,N_22064);
and U25261 (N_25261,N_22969,N_23431);
nand U25262 (N_25262,N_22180,N_22216);
or U25263 (N_25263,N_23907,N_23413);
nand U25264 (N_25264,N_22520,N_22312);
nand U25265 (N_25265,N_22581,N_22866);
and U25266 (N_25266,N_23795,N_22792);
or U25267 (N_25267,N_23258,N_23386);
nor U25268 (N_25268,N_22481,N_23828);
nor U25269 (N_25269,N_22806,N_22078);
or U25270 (N_25270,N_23913,N_22861);
nand U25271 (N_25271,N_22220,N_23080);
nand U25272 (N_25272,N_23468,N_22716);
nor U25273 (N_25273,N_23530,N_22899);
xnor U25274 (N_25274,N_23470,N_22419);
nor U25275 (N_25275,N_22167,N_23830);
xnor U25276 (N_25276,N_22581,N_22270);
or U25277 (N_25277,N_23736,N_22349);
nand U25278 (N_25278,N_23662,N_23094);
and U25279 (N_25279,N_22166,N_23751);
nand U25280 (N_25280,N_23631,N_23123);
or U25281 (N_25281,N_23928,N_23103);
and U25282 (N_25282,N_23156,N_23996);
nor U25283 (N_25283,N_23287,N_22115);
nor U25284 (N_25284,N_22744,N_23548);
nor U25285 (N_25285,N_22912,N_23785);
xor U25286 (N_25286,N_23688,N_22598);
and U25287 (N_25287,N_23522,N_22421);
xor U25288 (N_25288,N_23756,N_22770);
nor U25289 (N_25289,N_22998,N_23814);
nor U25290 (N_25290,N_22783,N_22501);
xnor U25291 (N_25291,N_23584,N_23101);
and U25292 (N_25292,N_22129,N_23419);
nor U25293 (N_25293,N_23243,N_22303);
nand U25294 (N_25294,N_23166,N_23895);
xor U25295 (N_25295,N_22427,N_22651);
nand U25296 (N_25296,N_22190,N_23677);
xnor U25297 (N_25297,N_23569,N_23455);
nand U25298 (N_25298,N_22887,N_23183);
or U25299 (N_25299,N_23394,N_23685);
and U25300 (N_25300,N_22359,N_23946);
or U25301 (N_25301,N_22663,N_23961);
xor U25302 (N_25302,N_23771,N_23307);
xnor U25303 (N_25303,N_23872,N_23792);
xor U25304 (N_25304,N_22215,N_22145);
xnor U25305 (N_25305,N_23115,N_22128);
xnor U25306 (N_25306,N_22209,N_23318);
and U25307 (N_25307,N_23093,N_22990);
or U25308 (N_25308,N_23489,N_22003);
xnor U25309 (N_25309,N_22948,N_23063);
or U25310 (N_25310,N_23120,N_22152);
nand U25311 (N_25311,N_23682,N_23835);
xor U25312 (N_25312,N_22193,N_22922);
nand U25313 (N_25313,N_23260,N_23286);
or U25314 (N_25314,N_22963,N_22504);
and U25315 (N_25315,N_23340,N_23818);
nand U25316 (N_25316,N_23870,N_23451);
nor U25317 (N_25317,N_22284,N_22612);
or U25318 (N_25318,N_23685,N_22933);
nand U25319 (N_25319,N_23216,N_23109);
or U25320 (N_25320,N_22351,N_23776);
nand U25321 (N_25321,N_22495,N_22294);
or U25322 (N_25322,N_22073,N_23540);
or U25323 (N_25323,N_23980,N_22472);
nor U25324 (N_25324,N_23862,N_22985);
nand U25325 (N_25325,N_22273,N_22861);
or U25326 (N_25326,N_22307,N_22554);
xor U25327 (N_25327,N_22279,N_23964);
or U25328 (N_25328,N_23572,N_23790);
nand U25329 (N_25329,N_22450,N_23919);
or U25330 (N_25330,N_23099,N_23132);
and U25331 (N_25331,N_23697,N_22015);
xnor U25332 (N_25332,N_22132,N_23350);
and U25333 (N_25333,N_23992,N_23881);
or U25334 (N_25334,N_22356,N_23119);
and U25335 (N_25335,N_22146,N_22654);
xnor U25336 (N_25336,N_23786,N_22256);
or U25337 (N_25337,N_22608,N_22481);
nand U25338 (N_25338,N_23697,N_22949);
and U25339 (N_25339,N_23372,N_22341);
or U25340 (N_25340,N_22664,N_22818);
nor U25341 (N_25341,N_23373,N_22006);
or U25342 (N_25342,N_23658,N_23619);
and U25343 (N_25343,N_23357,N_23140);
or U25344 (N_25344,N_22241,N_23240);
or U25345 (N_25345,N_23298,N_22897);
nor U25346 (N_25346,N_23026,N_22890);
xnor U25347 (N_25347,N_23487,N_22883);
or U25348 (N_25348,N_23183,N_23746);
or U25349 (N_25349,N_23132,N_23182);
or U25350 (N_25350,N_22212,N_22773);
nand U25351 (N_25351,N_23807,N_22539);
xnor U25352 (N_25352,N_23026,N_22369);
nand U25353 (N_25353,N_23116,N_22433);
nand U25354 (N_25354,N_22593,N_22007);
nand U25355 (N_25355,N_23203,N_22657);
nand U25356 (N_25356,N_22410,N_22916);
and U25357 (N_25357,N_22055,N_23936);
nand U25358 (N_25358,N_23168,N_22008);
and U25359 (N_25359,N_22041,N_22695);
nand U25360 (N_25360,N_22211,N_22759);
xor U25361 (N_25361,N_22750,N_22650);
and U25362 (N_25362,N_23809,N_22397);
nand U25363 (N_25363,N_22100,N_22945);
nand U25364 (N_25364,N_23019,N_22592);
nor U25365 (N_25365,N_22603,N_23681);
and U25366 (N_25366,N_23996,N_23145);
nor U25367 (N_25367,N_22063,N_22289);
nor U25368 (N_25368,N_23538,N_22957);
and U25369 (N_25369,N_23297,N_22948);
nand U25370 (N_25370,N_22145,N_22007);
nand U25371 (N_25371,N_23052,N_22736);
nand U25372 (N_25372,N_23566,N_23626);
and U25373 (N_25373,N_22142,N_23787);
nand U25374 (N_25374,N_22440,N_22018);
and U25375 (N_25375,N_23041,N_22348);
nor U25376 (N_25376,N_23959,N_22349);
and U25377 (N_25377,N_23961,N_23832);
or U25378 (N_25378,N_22731,N_22788);
and U25379 (N_25379,N_22031,N_22147);
nor U25380 (N_25380,N_22265,N_22644);
nand U25381 (N_25381,N_22320,N_23925);
nand U25382 (N_25382,N_23038,N_23374);
nor U25383 (N_25383,N_22607,N_23797);
and U25384 (N_25384,N_22403,N_22495);
and U25385 (N_25385,N_23421,N_22140);
nor U25386 (N_25386,N_23383,N_22220);
and U25387 (N_25387,N_22523,N_22953);
nor U25388 (N_25388,N_22640,N_22895);
nand U25389 (N_25389,N_23452,N_23022);
nand U25390 (N_25390,N_22869,N_23024);
and U25391 (N_25391,N_23622,N_22769);
xor U25392 (N_25392,N_23656,N_22103);
nor U25393 (N_25393,N_22783,N_22438);
nand U25394 (N_25394,N_23223,N_22264);
xor U25395 (N_25395,N_23235,N_22183);
nand U25396 (N_25396,N_22137,N_22828);
nand U25397 (N_25397,N_22050,N_22427);
and U25398 (N_25398,N_22963,N_23281);
xor U25399 (N_25399,N_23609,N_22903);
and U25400 (N_25400,N_22067,N_23996);
nand U25401 (N_25401,N_22126,N_23735);
or U25402 (N_25402,N_22876,N_22912);
nor U25403 (N_25403,N_23990,N_23559);
or U25404 (N_25404,N_22271,N_23779);
nor U25405 (N_25405,N_22194,N_22179);
or U25406 (N_25406,N_22718,N_22474);
or U25407 (N_25407,N_22109,N_23032);
nand U25408 (N_25408,N_22752,N_23796);
nor U25409 (N_25409,N_23145,N_22727);
nor U25410 (N_25410,N_22968,N_23609);
xnor U25411 (N_25411,N_22303,N_23312);
or U25412 (N_25412,N_22545,N_22040);
xor U25413 (N_25413,N_23032,N_22360);
nand U25414 (N_25414,N_23972,N_23099);
and U25415 (N_25415,N_22886,N_22304);
nand U25416 (N_25416,N_23920,N_22655);
and U25417 (N_25417,N_22549,N_22867);
or U25418 (N_25418,N_23683,N_22451);
nor U25419 (N_25419,N_22729,N_22569);
nor U25420 (N_25420,N_23921,N_23425);
xnor U25421 (N_25421,N_22500,N_23811);
and U25422 (N_25422,N_23378,N_22710);
xor U25423 (N_25423,N_23727,N_22347);
xnor U25424 (N_25424,N_22373,N_22536);
or U25425 (N_25425,N_23279,N_23248);
nand U25426 (N_25426,N_22826,N_22011);
or U25427 (N_25427,N_22861,N_22216);
or U25428 (N_25428,N_22865,N_23480);
and U25429 (N_25429,N_23557,N_23417);
and U25430 (N_25430,N_22028,N_23217);
nand U25431 (N_25431,N_23403,N_23389);
nor U25432 (N_25432,N_22342,N_23868);
nor U25433 (N_25433,N_23043,N_23097);
xnor U25434 (N_25434,N_22588,N_22542);
nand U25435 (N_25435,N_22285,N_23659);
or U25436 (N_25436,N_23474,N_22444);
nor U25437 (N_25437,N_22721,N_23419);
or U25438 (N_25438,N_23407,N_23921);
or U25439 (N_25439,N_22981,N_23946);
or U25440 (N_25440,N_23564,N_23418);
or U25441 (N_25441,N_23897,N_23561);
nand U25442 (N_25442,N_23973,N_22351);
xnor U25443 (N_25443,N_23908,N_22241);
nor U25444 (N_25444,N_23143,N_23371);
xnor U25445 (N_25445,N_23030,N_23120);
nand U25446 (N_25446,N_23543,N_22683);
xor U25447 (N_25447,N_22430,N_22686);
nor U25448 (N_25448,N_22429,N_22265);
or U25449 (N_25449,N_22408,N_22406);
nand U25450 (N_25450,N_22422,N_22371);
and U25451 (N_25451,N_23320,N_23631);
nand U25452 (N_25452,N_22423,N_23297);
and U25453 (N_25453,N_23010,N_23637);
nor U25454 (N_25454,N_22958,N_22330);
nor U25455 (N_25455,N_23514,N_23878);
nand U25456 (N_25456,N_23572,N_23865);
or U25457 (N_25457,N_22174,N_22822);
and U25458 (N_25458,N_22889,N_22723);
or U25459 (N_25459,N_23348,N_23988);
nor U25460 (N_25460,N_22044,N_22945);
xnor U25461 (N_25461,N_22113,N_23555);
nor U25462 (N_25462,N_23886,N_22538);
nand U25463 (N_25463,N_23034,N_22136);
nand U25464 (N_25464,N_23981,N_23718);
or U25465 (N_25465,N_22715,N_22403);
nand U25466 (N_25466,N_22384,N_23561);
xor U25467 (N_25467,N_22096,N_22337);
nand U25468 (N_25468,N_22205,N_23452);
xnor U25469 (N_25469,N_23362,N_23085);
xnor U25470 (N_25470,N_22135,N_22501);
xor U25471 (N_25471,N_23343,N_22910);
nand U25472 (N_25472,N_22837,N_22942);
and U25473 (N_25473,N_22406,N_23070);
or U25474 (N_25474,N_22293,N_22176);
xor U25475 (N_25475,N_22798,N_23566);
nand U25476 (N_25476,N_22005,N_23318);
nand U25477 (N_25477,N_23864,N_23636);
or U25478 (N_25478,N_22492,N_22048);
or U25479 (N_25479,N_23472,N_22405);
nor U25480 (N_25480,N_23446,N_23986);
nor U25481 (N_25481,N_22488,N_23978);
nand U25482 (N_25482,N_23399,N_23546);
nor U25483 (N_25483,N_23489,N_23863);
or U25484 (N_25484,N_22130,N_22137);
xnor U25485 (N_25485,N_22027,N_23817);
nand U25486 (N_25486,N_22250,N_23322);
xnor U25487 (N_25487,N_23140,N_23389);
nor U25488 (N_25488,N_22189,N_22613);
nor U25489 (N_25489,N_22177,N_23884);
nor U25490 (N_25490,N_22071,N_23789);
nand U25491 (N_25491,N_22364,N_22438);
nand U25492 (N_25492,N_22794,N_22234);
and U25493 (N_25493,N_22089,N_22263);
xor U25494 (N_25494,N_22517,N_23432);
or U25495 (N_25495,N_23536,N_22582);
and U25496 (N_25496,N_23502,N_22913);
nand U25497 (N_25497,N_23848,N_22453);
and U25498 (N_25498,N_23106,N_23860);
or U25499 (N_25499,N_23907,N_23598);
nor U25500 (N_25500,N_22693,N_22330);
nand U25501 (N_25501,N_22382,N_22059);
nand U25502 (N_25502,N_23704,N_23290);
or U25503 (N_25503,N_23846,N_23775);
and U25504 (N_25504,N_23003,N_22816);
nand U25505 (N_25505,N_23470,N_22998);
nand U25506 (N_25506,N_22709,N_22164);
nor U25507 (N_25507,N_23721,N_23647);
and U25508 (N_25508,N_23490,N_22093);
nor U25509 (N_25509,N_23503,N_22136);
and U25510 (N_25510,N_22985,N_22720);
or U25511 (N_25511,N_22542,N_22838);
and U25512 (N_25512,N_22227,N_23261);
nand U25513 (N_25513,N_23543,N_22573);
xnor U25514 (N_25514,N_22866,N_23139);
and U25515 (N_25515,N_22863,N_23678);
xnor U25516 (N_25516,N_22238,N_22102);
nor U25517 (N_25517,N_22415,N_23698);
and U25518 (N_25518,N_23615,N_22094);
nand U25519 (N_25519,N_22024,N_22779);
xnor U25520 (N_25520,N_22752,N_22531);
or U25521 (N_25521,N_22335,N_22948);
or U25522 (N_25522,N_23835,N_22436);
and U25523 (N_25523,N_22234,N_23583);
or U25524 (N_25524,N_22414,N_22413);
or U25525 (N_25525,N_22460,N_23936);
nand U25526 (N_25526,N_22781,N_23958);
and U25527 (N_25527,N_23463,N_23826);
or U25528 (N_25528,N_23755,N_23686);
and U25529 (N_25529,N_22069,N_22542);
nor U25530 (N_25530,N_23538,N_23609);
nand U25531 (N_25531,N_22275,N_23348);
xor U25532 (N_25532,N_23970,N_23472);
and U25533 (N_25533,N_23018,N_23508);
xor U25534 (N_25534,N_23644,N_23525);
or U25535 (N_25535,N_23210,N_23720);
nand U25536 (N_25536,N_22852,N_23406);
or U25537 (N_25537,N_23143,N_23254);
and U25538 (N_25538,N_23047,N_23558);
and U25539 (N_25539,N_23402,N_22501);
or U25540 (N_25540,N_23786,N_23129);
xor U25541 (N_25541,N_23234,N_22069);
nor U25542 (N_25542,N_22827,N_22337);
or U25543 (N_25543,N_22292,N_22652);
and U25544 (N_25544,N_23947,N_23971);
and U25545 (N_25545,N_23065,N_22065);
and U25546 (N_25546,N_22659,N_23535);
nand U25547 (N_25547,N_22243,N_23460);
or U25548 (N_25548,N_23113,N_23183);
nor U25549 (N_25549,N_23927,N_23419);
and U25550 (N_25550,N_23948,N_22137);
xor U25551 (N_25551,N_22674,N_23027);
nand U25552 (N_25552,N_23554,N_23970);
and U25553 (N_25553,N_23818,N_22645);
and U25554 (N_25554,N_22562,N_23547);
nor U25555 (N_25555,N_23666,N_22201);
or U25556 (N_25556,N_23165,N_23921);
xnor U25557 (N_25557,N_23487,N_23232);
or U25558 (N_25558,N_23345,N_22498);
nor U25559 (N_25559,N_22807,N_22059);
nand U25560 (N_25560,N_22560,N_22998);
nor U25561 (N_25561,N_22008,N_23704);
nor U25562 (N_25562,N_22350,N_22534);
xor U25563 (N_25563,N_23257,N_23801);
nand U25564 (N_25564,N_23126,N_23973);
nand U25565 (N_25565,N_22094,N_23664);
and U25566 (N_25566,N_22830,N_22885);
or U25567 (N_25567,N_23306,N_23446);
or U25568 (N_25568,N_22764,N_22159);
or U25569 (N_25569,N_22686,N_23698);
nor U25570 (N_25570,N_23261,N_23788);
nor U25571 (N_25571,N_23496,N_23159);
nor U25572 (N_25572,N_23374,N_23319);
nand U25573 (N_25573,N_22278,N_22611);
xnor U25574 (N_25574,N_23910,N_23074);
nand U25575 (N_25575,N_22331,N_22694);
nand U25576 (N_25576,N_22602,N_22609);
or U25577 (N_25577,N_22043,N_23695);
or U25578 (N_25578,N_22703,N_22306);
or U25579 (N_25579,N_23163,N_23918);
and U25580 (N_25580,N_22819,N_23236);
or U25581 (N_25581,N_23782,N_22184);
xor U25582 (N_25582,N_22538,N_22877);
xnor U25583 (N_25583,N_22973,N_22442);
xor U25584 (N_25584,N_22720,N_22948);
or U25585 (N_25585,N_23984,N_23695);
xnor U25586 (N_25586,N_23702,N_22881);
xor U25587 (N_25587,N_23321,N_22141);
nand U25588 (N_25588,N_23448,N_23501);
and U25589 (N_25589,N_23912,N_22900);
nand U25590 (N_25590,N_23591,N_23708);
nor U25591 (N_25591,N_23685,N_23468);
nor U25592 (N_25592,N_22136,N_22608);
and U25593 (N_25593,N_22980,N_23942);
and U25594 (N_25594,N_22069,N_22596);
or U25595 (N_25595,N_22273,N_22118);
and U25596 (N_25596,N_23653,N_23440);
xor U25597 (N_25597,N_22663,N_23559);
xor U25598 (N_25598,N_22714,N_22766);
and U25599 (N_25599,N_23998,N_23777);
and U25600 (N_25600,N_23760,N_23898);
nand U25601 (N_25601,N_22076,N_22126);
or U25602 (N_25602,N_23058,N_23274);
and U25603 (N_25603,N_22884,N_23959);
and U25604 (N_25604,N_23537,N_23861);
or U25605 (N_25605,N_22866,N_23513);
xnor U25606 (N_25606,N_23439,N_23032);
and U25607 (N_25607,N_23236,N_23848);
nand U25608 (N_25608,N_22253,N_23219);
xnor U25609 (N_25609,N_22301,N_23695);
and U25610 (N_25610,N_23697,N_22294);
nor U25611 (N_25611,N_23021,N_22568);
or U25612 (N_25612,N_23998,N_22622);
or U25613 (N_25613,N_23756,N_23374);
nor U25614 (N_25614,N_22560,N_23960);
nor U25615 (N_25615,N_22556,N_22434);
or U25616 (N_25616,N_22399,N_22330);
nor U25617 (N_25617,N_23638,N_23473);
xnor U25618 (N_25618,N_23191,N_23984);
and U25619 (N_25619,N_22587,N_22356);
and U25620 (N_25620,N_22702,N_23398);
xor U25621 (N_25621,N_23082,N_22741);
nand U25622 (N_25622,N_23060,N_22782);
or U25623 (N_25623,N_22362,N_22294);
xor U25624 (N_25624,N_23951,N_22487);
nand U25625 (N_25625,N_23790,N_22616);
xor U25626 (N_25626,N_23794,N_23665);
nand U25627 (N_25627,N_22906,N_22293);
and U25628 (N_25628,N_23886,N_22896);
or U25629 (N_25629,N_22092,N_22188);
nand U25630 (N_25630,N_22797,N_22535);
nand U25631 (N_25631,N_23741,N_23864);
and U25632 (N_25632,N_22581,N_22813);
nor U25633 (N_25633,N_22164,N_22358);
nand U25634 (N_25634,N_23648,N_23285);
and U25635 (N_25635,N_23929,N_23230);
xor U25636 (N_25636,N_22816,N_22714);
nor U25637 (N_25637,N_22489,N_23972);
or U25638 (N_25638,N_22452,N_23626);
and U25639 (N_25639,N_22095,N_23731);
nor U25640 (N_25640,N_23424,N_22465);
nand U25641 (N_25641,N_23822,N_22364);
or U25642 (N_25642,N_22864,N_23689);
and U25643 (N_25643,N_22856,N_22186);
xor U25644 (N_25644,N_23876,N_22451);
xnor U25645 (N_25645,N_22090,N_23035);
and U25646 (N_25646,N_23723,N_22074);
nand U25647 (N_25647,N_22298,N_22500);
nor U25648 (N_25648,N_22896,N_22009);
and U25649 (N_25649,N_22884,N_22936);
xor U25650 (N_25650,N_22700,N_22362);
nor U25651 (N_25651,N_23016,N_22043);
or U25652 (N_25652,N_22288,N_22147);
nor U25653 (N_25653,N_23600,N_22858);
nor U25654 (N_25654,N_23541,N_23767);
and U25655 (N_25655,N_22970,N_22666);
nor U25656 (N_25656,N_22300,N_23651);
or U25657 (N_25657,N_23743,N_23541);
nor U25658 (N_25658,N_23485,N_23194);
xnor U25659 (N_25659,N_23271,N_22642);
nand U25660 (N_25660,N_22993,N_22332);
nor U25661 (N_25661,N_23277,N_22260);
nor U25662 (N_25662,N_22758,N_22394);
xnor U25663 (N_25663,N_23068,N_23462);
nand U25664 (N_25664,N_22136,N_23712);
and U25665 (N_25665,N_23953,N_23264);
nor U25666 (N_25666,N_22152,N_23985);
nand U25667 (N_25667,N_23222,N_23210);
nand U25668 (N_25668,N_22784,N_23900);
or U25669 (N_25669,N_22606,N_22345);
nand U25670 (N_25670,N_22209,N_22540);
nand U25671 (N_25671,N_22781,N_22077);
xnor U25672 (N_25672,N_22113,N_23163);
nand U25673 (N_25673,N_22912,N_23543);
and U25674 (N_25674,N_22765,N_22749);
and U25675 (N_25675,N_22372,N_23800);
xnor U25676 (N_25676,N_23450,N_22162);
xor U25677 (N_25677,N_23456,N_23778);
xnor U25678 (N_25678,N_22238,N_23133);
and U25679 (N_25679,N_23292,N_22281);
and U25680 (N_25680,N_22681,N_22471);
or U25681 (N_25681,N_22033,N_22865);
xor U25682 (N_25682,N_22811,N_22167);
or U25683 (N_25683,N_23875,N_23464);
nand U25684 (N_25684,N_23670,N_22157);
and U25685 (N_25685,N_23260,N_22997);
or U25686 (N_25686,N_23758,N_23841);
xnor U25687 (N_25687,N_22613,N_23751);
nor U25688 (N_25688,N_23151,N_23332);
xnor U25689 (N_25689,N_22760,N_22198);
or U25690 (N_25690,N_23888,N_22018);
or U25691 (N_25691,N_22474,N_22656);
xnor U25692 (N_25692,N_23334,N_22544);
or U25693 (N_25693,N_22861,N_23964);
xnor U25694 (N_25694,N_23364,N_22013);
or U25695 (N_25695,N_22302,N_23850);
nand U25696 (N_25696,N_22383,N_23980);
nand U25697 (N_25697,N_23815,N_22629);
or U25698 (N_25698,N_23709,N_22651);
nor U25699 (N_25699,N_23168,N_22265);
nor U25700 (N_25700,N_23068,N_22110);
xor U25701 (N_25701,N_22238,N_23178);
or U25702 (N_25702,N_23245,N_23135);
nor U25703 (N_25703,N_22275,N_23586);
nand U25704 (N_25704,N_22832,N_23858);
nand U25705 (N_25705,N_22475,N_22882);
and U25706 (N_25706,N_23207,N_23322);
nand U25707 (N_25707,N_22341,N_23393);
nand U25708 (N_25708,N_22357,N_23969);
xor U25709 (N_25709,N_23526,N_22555);
or U25710 (N_25710,N_23845,N_23981);
nand U25711 (N_25711,N_23162,N_23004);
nor U25712 (N_25712,N_23111,N_22236);
and U25713 (N_25713,N_22446,N_23308);
xor U25714 (N_25714,N_22958,N_23749);
nor U25715 (N_25715,N_22687,N_22998);
or U25716 (N_25716,N_23522,N_22454);
nor U25717 (N_25717,N_23243,N_23616);
or U25718 (N_25718,N_22412,N_22939);
or U25719 (N_25719,N_23510,N_23315);
nor U25720 (N_25720,N_22935,N_22825);
and U25721 (N_25721,N_23325,N_23576);
and U25722 (N_25722,N_22192,N_23118);
and U25723 (N_25723,N_23966,N_22703);
and U25724 (N_25724,N_23704,N_22948);
nand U25725 (N_25725,N_23370,N_23757);
nand U25726 (N_25726,N_23047,N_23299);
nand U25727 (N_25727,N_23366,N_23777);
xor U25728 (N_25728,N_22925,N_22321);
nor U25729 (N_25729,N_23306,N_23374);
nand U25730 (N_25730,N_22724,N_22203);
or U25731 (N_25731,N_23893,N_22204);
and U25732 (N_25732,N_22389,N_23188);
or U25733 (N_25733,N_23719,N_23721);
nor U25734 (N_25734,N_22934,N_23932);
and U25735 (N_25735,N_23473,N_22001);
nand U25736 (N_25736,N_22633,N_22455);
nor U25737 (N_25737,N_22091,N_23443);
and U25738 (N_25738,N_23429,N_23374);
nand U25739 (N_25739,N_22434,N_23047);
xor U25740 (N_25740,N_23637,N_22244);
nand U25741 (N_25741,N_23318,N_23072);
nor U25742 (N_25742,N_23951,N_23136);
xnor U25743 (N_25743,N_23752,N_22397);
and U25744 (N_25744,N_22379,N_22313);
or U25745 (N_25745,N_23798,N_23564);
xor U25746 (N_25746,N_23952,N_23714);
nor U25747 (N_25747,N_22064,N_23165);
nand U25748 (N_25748,N_22319,N_23736);
nor U25749 (N_25749,N_22595,N_22850);
nor U25750 (N_25750,N_22291,N_23417);
nand U25751 (N_25751,N_22240,N_22416);
nor U25752 (N_25752,N_23663,N_23197);
nor U25753 (N_25753,N_23219,N_22662);
or U25754 (N_25754,N_23319,N_22927);
or U25755 (N_25755,N_23999,N_22255);
nand U25756 (N_25756,N_23465,N_23983);
nor U25757 (N_25757,N_23077,N_22594);
xnor U25758 (N_25758,N_23954,N_22843);
nor U25759 (N_25759,N_22469,N_22150);
and U25760 (N_25760,N_22504,N_23820);
nor U25761 (N_25761,N_23338,N_22566);
and U25762 (N_25762,N_23359,N_22715);
nand U25763 (N_25763,N_22511,N_22955);
nand U25764 (N_25764,N_23013,N_23319);
xor U25765 (N_25765,N_23383,N_22052);
and U25766 (N_25766,N_23135,N_22731);
nor U25767 (N_25767,N_22832,N_22002);
xnor U25768 (N_25768,N_23411,N_22071);
or U25769 (N_25769,N_23190,N_22790);
nor U25770 (N_25770,N_23124,N_22770);
nand U25771 (N_25771,N_23813,N_22309);
or U25772 (N_25772,N_22200,N_23379);
xnor U25773 (N_25773,N_22417,N_22795);
xnor U25774 (N_25774,N_22247,N_23720);
and U25775 (N_25775,N_23848,N_23932);
or U25776 (N_25776,N_22998,N_23308);
xnor U25777 (N_25777,N_22025,N_23139);
or U25778 (N_25778,N_23530,N_23350);
nand U25779 (N_25779,N_23645,N_22126);
nor U25780 (N_25780,N_23114,N_23851);
nand U25781 (N_25781,N_23399,N_22807);
and U25782 (N_25782,N_22653,N_22502);
nor U25783 (N_25783,N_23621,N_22680);
nor U25784 (N_25784,N_22766,N_22433);
and U25785 (N_25785,N_22719,N_23274);
or U25786 (N_25786,N_22634,N_22388);
or U25787 (N_25787,N_23082,N_22440);
or U25788 (N_25788,N_22254,N_23293);
nand U25789 (N_25789,N_22345,N_23426);
xor U25790 (N_25790,N_23044,N_23823);
nand U25791 (N_25791,N_22692,N_22163);
xor U25792 (N_25792,N_23763,N_23941);
and U25793 (N_25793,N_23183,N_22318);
xnor U25794 (N_25794,N_22083,N_22422);
xor U25795 (N_25795,N_23467,N_23154);
nor U25796 (N_25796,N_22296,N_23331);
and U25797 (N_25797,N_23865,N_23117);
xnor U25798 (N_25798,N_23267,N_23342);
or U25799 (N_25799,N_22937,N_22249);
nor U25800 (N_25800,N_22726,N_22205);
and U25801 (N_25801,N_22922,N_23967);
nand U25802 (N_25802,N_23449,N_22418);
xor U25803 (N_25803,N_22946,N_23654);
xor U25804 (N_25804,N_22349,N_23152);
and U25805 (N_25805,N_23724,N_23273);
xor U25806 (N_25806,N_22536,N_23239);
nand U25807 (N_25807,N_22327,N_22714);
xnor U25808 (N_25808,N_22321,N_22046);
nand U25809 (N_25809,N_22211,N_23609);
nor U25810 (N_25810,N_23639,N_22378);
nand U25811 (N_25811,N_23917,N_23851);
nand U25812 (N_25812,N_22870,N_23912);
or U25813 (N_25813,N_22654,N_22406);
nand U25814 (N_25814,N_22178,N_22257);
nor U25815 (N_25815,N_22627,N_22109);
xor U25816 (N_25816,N_23586,N_22633);
nand U25817 (N_25817,N_22547,N_22999);
or U25818 (N_25818,N_22790,N_22623);
or U25819 (N_25819,N_22749,N_23333);
or U25820 (N_25820,N_22222,N_23631);
and U25821 (N_25821,N_22226,N_23072);
or U25822 (N_25822,N_22183,N_22826);
nor U25823 (N_25823,N_23170,N_22237);
nand U25824 (N_25824,N_22231,N_23314);
nand U25825 (N_25825,N_22183,N_23804);
xor U25826 (N_25826,N_22345,N_22990);
nor U25827 (N_25827,N_23141,N_22756);
nor U25828 (N_25828,N_23074,N_22883);
xor U25829 (N_25829,N_23113,N_22646);
nand U25830 (N_25830,N_22500,N_22435);
xnor U25831 (N_25831,N_22244,N_22111);
nand U25832 (N_25832,N_23525,N_22468);
nor U25833 (N_25833,N_22857,N_22590);
xnor U25834 (N_25834,N_22374,N_23570);
xnor U25835 (N_25835,N_22759,N_23896);
or U25836 (N_25836,N_22867,N_22145);
and U25837 (N_25837,N_22233,N_23495);
xor U25838 (N_25838,N_22316,N_23561);
or U25839 (N_25839,N_22282,N_22977);
nor U25840 (N_25840,N_23341,N_23280);
xnor U25841 (N_25841,N_23710,N_23546);
xnor U25842 (N_25842,N_22303,N_22978);
xor U25843 (N_25843,N_23405,N_22702);
or U25844 (N_25844,N_22781,N_22912);
or U25845 (N_25845,N_23907,N_22875);
xnor U25846 (N_25846,N_22847,N_23466);
and U25847 (N_25847,N_22615,N_22118);
and U25848 (N_25848,N_22867,N_23231);
and U25849 (N_25849,N_22873,N_23446);
nor U25850 (N_25850,N_23054,N_23504);
nor U25851 (N_25851,N_22928,N_22829);
or U25852 (N_25852,N_22352,N_22371);
nand U25853 (N_25853,N_23736,N_23864);
or U25854 (N_25854,N_23284,N_23922);
and U25855 (N_25855,N_23602,N_22893);
or U25856 (N_25856,N_23649,N_22040);
nor U25857 (N_25857,N_23416,N_22099);
nor U25858 (N_25858,N_22103,N_22215);
nand U25859 (N_25859,N_22064,N_22403);
or U25860 (N_25860,N_23281,N_23815);
nor U25861 (N_25861,N_23503,N_23414);
and U25862 (N_25862,N_23421,N_23649);
nor U25863 (N_25863,N_23172,N_23960);
nand U25864 (N_25864,N_22089,N_23145);
and U25865 (N_25865,N_22240,N_22131);
and U25866 (N_25866,N_22939,N_22920);
or U25867 (N_25867,N_23225,N_23171);
and U25868 (N_25868,N_23995,N_22510);
nor U25869 (N_25869,N_22559,N_23255);
nand U25870 (N_25870,N_23053,N_23273);
xor U25871 (N_25871,N_23489,N_23985);
nor U25872 (N_25872,N_22858,N_23942);
nand U25873 (N_25873,N_22282,N_23996);
nand U25874 (N_25874,N_22365,N_23151);
or U25875 (N_25875,N_23752,N_23630);
and U25876 (N_25876,N_23999,N_23509);
or U25877 (N_25877,N_23433,N_22272);
and U25878 (N_25878,N_22570,N_22220);
or U25879 (N_25879,N_23536,N_22133);
and U25880 (N_25880,N_22413,N_22008);
and U25881 (N_25881,N_23978,N_23492);
xnor U25882 (N_25882,N_23807,N_22077);
or U25883 (N_25883,N_23641,N_22871);
nand U25884 (N_25884,N_22833,N_22617);
nand U25885 (N_25885,N_23172,N_23570);
and U25886 (N_25886,N_23768,N_22569);
nor U25887 (N_25887,N_22091,N_23647);
nand U25888 (N_25888,N_22233,N_22111);
nor U25889 (N_25889,N_22781,N_23338);
nand U25890 (N_25890,N_22455,N_22846);
nand U25891 (N_25891,N_22352,N_22234);
xnor U25892 (N_25892,N_23459,N_23771);
nor U25893 (N_25893,N_23180,N_23455);
and U25894 (N_25894,N_22190,N_23929);
or U25895 (N_25895,N_22805,N_23269);
or U25896 (N_25896,N_23573,N_23098);
xnor U25897 (N_25897,N_23355,N_22113);
xor U25898 (N_25898,N_22475,N_22043);
nand U25899 (N_25899,N_23093,N_22004);
or U25900 (N_25900,N_23981,N_22454);
xor U25901 (N_25901,N_22248,N_23021);
or U25902 (N_25902,N_22682,N_23350);
nand U25903 (N_25903,N_22738,N_23608);
xor U25904 (N_25904,N_22425,N_23619);
or U25905 (N_25905,N_22945,N_23208);
nand U25906 (N_25906,N_23042,N_22524);
xnor U25907 (N_25907,N_23951,N_22020);
nor U25908 (N_25908,N_22888,N_22711);
and U25909 (N_25909,N_22930,N_22339);
xor U25910 (N_25910,N_23653,N_23135);
and U25911 (N_25911,N_23376,N_23153);
or U25912 (N_25912,N_23439,N_22175);
and U25913 (N_25913,N_23465,N_22240);
nor U25914 (N_25914,N_23797,N_22514);
and U25915 (N_25915,N_22627,N_23722);
and U25916 (N_25916,N_23461,N_23761);
and U25917 (N_25917,N_22676,N_23152);
nand U25918 (N_25918,N_22571,N_22301);
xnor U25919 (N_25919,N_22289,N_22633);
nor U25920 (N_25920,N_23340,N_23377);
nor U25921 (N_25921,N_23849,N_23686);
and U25922 (N_25922,N_23016,N_23129);
or U25923 (N_25923,N_22646,N_22926);
nand U25924 (N_25924,N_23471,N_23443);
xor U25925 (N_25925,N_23030,N_22239);
nand U25926 (N_25926,N_23955,N_22479);
nand U25927 (N_25927,N_22012,N_22311);
nor U25928 (N_25928,N_22631,N_22348);
nand U25929 (N_25929,N_23200,N_23207);
nand U25930 (N_25930,N_22309,N_22688);
or U25931 (N_25931,N_22466,N_22230);
or U25932 (N_25932,N_23315,N_23919);
nand U25933 (N_25933,N_22499,N_22979);
or U25934 (N_25934,N_23104,N_23230);
or U25935 (N_25935,N_23464,N_22289);
or U25936 (N_25936,N_23706,N_23541);
nand U25937 (N_25937,N_23341,N_23755);
nand U25938 (N_25938,N_22322,N_23072);
and U25939 (N_25939,N_23567,N_23115);
nor U25940 (N_25940,N_23578,N_23291);
xor U25941 (N_25941,N_23873,N_23427);
and U25942 (N_25942,N_22847,N_23435);
nand U25943 (N_25943,N_22234,N_23406);
or U25944 (N_25944,N_22554,N_23529);
nor U25945 (N_25945,N_22719,N_23104);
or U25946 (N_25946,N_22645,N_22494);
and U25947 (N_25947,N_22131,N_22555);
and U25948 (N_25948,N_23451,N_23964);
or U25949 (N_25949,N_22319,N_23913);
nand U25950 (N_25950,N_22891,N_22339);
xor U25951 (N_25951,N_22518,N_23436);
xor U25952 (N_25952,N_22328,N_23238);
nor U25953 (N_25953,N_22522,N_22990);
nor U25954 (N_25954,N_23787,N_22333);
xnor U25955 (N_25955,N_23567,N_23126);
and U25956 (N_25956,N_22341,N_23970);
nor U25957 (N_25957,N_22803,N_22847);
xor U25958 (N_25958,N_22568,N_23587);
and U25959 (N_25959,N_22782,N_23600);
nand U25960 (N_25960,N_22800,N_23218);
and U25961 (N_25961,N_23997,N_23217);
nor U25962 (N_25962,N_23861,N_22708);
or U25963 (N_25963,N_23807,N_22546);
or U25964 (N_25964,N_23758,N_23086);
and U25965 (N_25965,N_22276,N_23164);
xnor U25966 (N_25966,N_22080,N_22841);
or U25967 (N_25967,N_23561,N_22681);
and U25968 (N_25968,N_23751,N_23221);
xnor U25969 (N_25969,N_23552,N_22643);
or U25970 (N_25970,N_23325,N_23801);
xnor U25971 (N_25971,N_23479,N_23362);
nor U25972 (N_25972,N_23931,N_23784);
or U25973 (N_25973,N_22860,N_23601);
nor U25974 (N_25974,N_22112,N_23412);
nor U25975 (N_25975,N_23023,N_23358);
or U25976 (N_25976,N_22262,N_23027);
nor U25977 (N_25977,N_23464,N_23599);
nor U25978 (N_25978,N_22858,N_22934);
xnor U25979 (N_25979,N_22451,N_22849);
nor U25980 (N_25980,N_22893,N_23000);
and U25981 (N_25981,N_22336,N_22799);
nor U25982 (N_25982,N_22736,N_22590);
nand U25983 (N_25983,N_22158,N_23371);
or U25984 (N_25984,N_23540,N_23104);
nor U25985 (N_25985,N_22244,N_23263);
nor U25986 (N_25986,N_22168,N_22952);
xnor U25987 (N_25987,N_23672,N_22140);
and U25988 (N_25988,N_23735,N_22545);
nor U25989 (N_25989,N_23986,N_23437);
nor U25990 (N_25990,N_22218,N_23282);
nand U25991 (N_25991,N_23269,N_22758);
nor U25992 (N_25992,N_23693,N_22324);
nor U25993 (N_25993,N_22621,N_22914);
and U25994 (N_25994,N_22522,N_23089);
and U25995 (N_25995,N_23757,N_23741);
nor U25996 (N_25996,N_23728,N_22815);
and U25997 (N_25997,N_23135,N_23157);
nor U25998 (N_25998,N_23147,N_22386);
xnor U25999 (N_25999,N_23999,N_22050);
or U26000 (N_26000,N_25423,N_24232);
or U26001 (N_26001,N_25328,N_24855);
and U26002 (N_26002,N_24079,N_25789);
nand U26003 (N_26003,N_24828,N_25231);
nor U26004 (N_26004,N_25071,N_25192);
and U26005 (N_26005,N_24992,N_24517);
or U26006 (N_26006,N_25548,N_24612);
nor U26007 (N_26007,N_24868,N_24241);
nor U26008 (N_26008,N_25927,N_24212);
nand U26009 (N_26009,N_25700,N_24845);
or U26010 (N_26010,N_25667,N_24599);
xor U26011 (N_26011,N_24162,N_24821);
or U26012 (N_26012,N_25591,N_24980);
or U26013 (N_26013,N_24383,N_25246);
nor U26014 (N_26014,N_25010,N_25310);
and U26015 (N_26015,N_25908,N_24959);
xnor U26016 (N_26016,N_24720,N_24535);
xnor U26017 (N_26017,N_24319,N_25422);
and U26018 (N_26018,N_25498,N_24370);
xnor U26019 (N_26019,N_25777,N_25191);
and U26020 (N_26020,N_25783,N_25032);
and U26021 (N_26021,N_24905,N_25823);
nand U26022 (N_26022,N_25483,N_24401);
nand U26023 (N_26023,N_25638,N_24406);
xnor U26024 (N_26024,N_25386,N_24938);
or U26025 (N_26025,N_25069,N_24777);
or U26026 (N_26026,N_25523,N_24113);
nor U26027 (N_26027,N_24875,N_25121);
xnor U26028 (N_26028,N_25558,N_25126);
nor U26029 (N_26029,N_25346,N_25016);
and U26030 (N_26030,N_24615,N_24862);
or U26031 (N_26031,N_25366,N_25172);
nor U26032 (N_26032,N_25274,N_24687);
nand U26033 (N_26033,N_24904,N_25288);
and U26034 (N_26034,N_25299,N_24671);
or U26035 (N_26035,N_25444,N_25578);
or U26036 (N_26036,N_25023,N_24657);
nor U26037 (N_26037,N_25350,N_24903);
xnor U26038 (N_26038,N_25182,N_25045);
or U26039 (N_26039,N_24573,N_24758);
nand U26040 (N_26040,N_24709,N_25799);
or U26041 (N_26041,N_25384,N_24073);
xnor U26042 (N_26042,N_24591,N_25501);
nand U26043 (N_26043,N_25096,N_24545);
nor U26044 (N_26044,N_25547,N_25780);
xnor U26045 (N_26045,N_25695,N_24864);
nand U26046 (N_26046,N_24397,N_25321);
or U26047 (N_26047,N_25183,N_25124);
nor U26048 (N_26048,N_25961,N_24306);
and U26049 (N_26049,N_25987,N_24295);
nand U26050 (N_26050,N_24956,N_25719);
nor U26051 (N_26051,N_25786,N_25872);
nand U26052 (N_26052,N_24963,N_24813);
xnor U26053 (N_26053,N_24568,N_24128);
xor U26054 (N_26054,N_24784,N_24254);
xor U26055 (N_26055,N_24613,N_24100);
nand U26056 (N_26056,N_24165,N_24153);
and U26057 (N_26057,N_24267,N_25448);
nor U26058 (N_26058,N_25820,N_24861);
nand U26059 (N_26059,N_24769,N_24891);
nand U26060 (N_26060,N_24061,N_25929);
nor U26061 (N_26061,N_24550,N_24327);
and U26062 (N_26062,N_24863,N_24393);
xor U26063 (N_26063,N_25199,N_24432);
and U26064 (N_26064,N_24754,N_25136);
and U26065 (N_26065,N_25073,N_24735);
nor U26066 (N_26066,N_25742,N_24378);
xnor U26067 (N_26067,N_24399,N_25038);
or U26068 (N_26068,N_25099,N_24848);
xnor U26069 (N_26069,N_25062,N_25259);
nor U26070 (N_26070,N_25382,N_25280);
nor U26071 (N_26071,N_24625,N_24317);
nor U26072 (N_26072,N_25112,N_24690);
and U26073 (N_26073,N_24194,N_25014);
nand U26074 (N_26074,N_24936,N_24227);
or U26075 (N_26075,N_24071,N_24453);
nor U26076 (N_26076,N_24078,N_24357);
xor U26077 (N_26077,N_25919,N_25075);
and U26078 (N_26078,N_24592,N_25909);
or U26079 (N_26079,N_24626,N_24792);
and U26080 (N_26080,N_24260,N_25019);
nor U26081 (N_26081,N_24977,N_24638);
nand U26082 (N_26082,N_24482,N_25599);
xor U26083 (N_26083,N_24567,N_25995);
nor U26084 (N_26084,N_25171,N_24576);
nand U26085 (N_26085,N_25204,N_25686);
and U26086 (N_26086,N_24301,N_25287);
or U26087 (N_26087,N_25392,N_24135);
nand U26088 (N_26088,N_25178,N_24070);
nor U26089 (N_26089,N_25602,N_25035);
and U26090 (N_26090,N_24964,N_25074);
xnor U26091 (N_26091,N_24400,N_24452);
xor U26092 (N_26092,N_25922,N_25911);
nor U26093 (N_26093,N_25736,N_24055);
nor U26094 (N_26094,N_25738,N_24705);
and U26095 (N_26095,N_24297,N_24202);
or U26096 (N_26096,N_24674,N_25026);
nor U26097 (N_26097,N_25962,N_25141);
and U26098 (N_26098,N_24971,N_24494);
and U26099 (N_26099,N_24003,N_24985);
nor U26100 (N_26100,N_25974,N_24666);
nand U26101 (N_26101,N_24640,N_24693);
nand U26102 (N_26102,N_24058,N_25406);
or U26103 (N_26103,N_24827,N_24802);
and U26104 (N_26104,N_24919,N_24787);
xor U26105 (N_26105,N_24990,N_25330);
or U26106 (N_26106,N_25201,N_24531);
xor U26107 (N_26107,N_25557,N_25085);
xnor U26108 (N_26108,N_25507,N_25898);
or U26109 (N_26109,N_24222,N_24155);
nand U26110 (N_26110,N_24385,N_24818);
nand U26111 (N_26111,N_25242,N_24087);
xor U26112 (N_26112,N_25505,N_25748);
nor U26113 (N_26113,N_24470,N_24923);
nand U26114 (N_26114,N_25939,N_25568);
and U26115 (N_26115,N_24477,N_24747);
nand U26116 (N_26116,N_25882,N_24487);
nand U26117 (N_26117,N_25292,N_24391);
nand U26118 (N_26118,N_25776,N_24791);
xor U26119 (N_26119,N_25362,N_25395);
nor U26120 (N_26120,N_25093,N_25671);
nand U26121 (N_26121,N_24285,N_25077);
and U26122 (N_26122,N_25132,N_25130);
and U26123 (N_26123,N_25825,N_25262);
and U26124 (N_26124,N_25159,N_24252);
and U26125 (N_26125,N_24525,N_25969);
xnor U26126 (N_26126,N_25434,N_24463);
and U26127 (N_26127,N_25937,N_24051);
xnor U26128 (N_26128,N_25743,N_25570);
nor U26129 (N_26129,N_25270,N_24719);
nand U26130 (N_26130,N_24121,N_25670);
or U26131 (N_26131,N_25691,N_24253);
xor U26132 (N_26132,N_25404,N_25796);
and U26133 (N_26133,N_25012,N_25369);
and U26134 (N_26134,N_25463,N_25488);
xor U26135 (N_26135,N_24352,N_25164);
and U26136 (N_26136,N_24586,N_24617);
nand U26137 (N_26137,N_24793,N_25834);
xor U26138 (N_26138,N_25646,N_24553);
nor U26139 (N_26139,N_24819,N_25980);
or U26140 (N_26140,N_24530,N_24644);
nand U26141 (N_26141,N_25542,N_25795);
nand U26142 (N_26142,N_24398,N_24384);
nor U26143 (N_26143,N_25835,N_25869);
nor U26144 (N_26144,N_25539,N_24095);
xnor U26145 (N_26145,N_24603,N_25530);
nand U26146 (N_26146,N_24271,N_24018);
and U26147 (N_26147,N_24105,N_24523);
nor U26148 (N_26148,N_24217,N_24506);
nor U26149 (N_26149,N_25689,N_25326);
xor U26150 (N_26150,N_24433,N_24094);
and U26151 (N_26151,N_24449,N_25146);
and U26152 (N_26152,N_24129,N_25137);
xor U26153 (N_26153,N_24972,N_24918);
and U26154 (N_26154,N_25634,N_25913);
or U26155 (N_26155,N_25286,N_25057);
nor U26156 (N_26156,N_24560,N_25458);
or U26157 (N_26157,N_24824,N_24526);
nor U26158 (N_26158,N_24011,N_24724);
nor U26159 (N_26159,N_25531,N_25829);
nor U26160 (N_26160,N_25865,N_24369);
or U26161 (N_26161,N_24697,N_25678);
nor U26162 (N_26162,N_25847,N_24218);
nor U26163 (N_26163,N_25416,N_25128);
nor U26164 (N_26164,N_25561,N_24542);
nor U26165 (N_26165,N_25639,N_24286);
xor U26166 (N_26166,N_24092,N_25914);
xor U26167 (N_26167,N_25772,N_25732);
or U26168 (N_26168,N_25197,N_24275);
and U26169 (N_26169,N_25936,N_25848);
nor U26170 (N_26170,N_25915,N_25988);
and U26171 (N_26171,N_25094,N_25791);
nor U26172 (N_26172,N_24368,N_25526);
nor U26173 (N_26173,N_25443,N_25475);
or U26174 (N_26174,N_25515,N_25902);
nand U26175 (N_26175,N_24839,N_24420);
nand U26176 (N_26176,N_25187,N_25767);
nor U26177 (N_26177,N_25842,N_25439);
nor U26178 (N_26178,N_25592,N_25029);
or U26179 (N_26179,N_25756,N_24009);
xor U26180 (N_26180,N_25389,N_25863);
and U26181 (N_26181,N_25473,N_24069);
or U26182 (N_26182,N_25903,N_25618);
or U26183 (N_26183,N_24183,N_24474);
nand U26184 (N_26184,N_24151,N_25880);
xor U26185 (N_26185,N_24686,N_25682);
or U26186 (N_26186,N_24587,N_25857);
nand U26187 (N_26187,N_25712,N_24302);
xor U26188 (N_26188,N_25413,N_25143);
or U26189 (N_26189,N_24388,N_25904);
nor U26190 (N_26190,N_24380,N_24130);
nor U26191 (N_26191,N_25551,N_25455);
xor U26192 (N_26192,N_25427,N_25418);
or U26193 (N_26193,N_24220,N_24326);
xnor U26194 (N_26194,N_25387,N_25556);
or U26195 (N_26195,N_24046,N_25749);
xor U26196 (N_26196,N_24975,N_24173);
nand U26197 (N_26197,N_24081,N_25658);
and U26198 (N_26198,N_24499,N_24473);
nand U26199 (N_26199,N_25706,N_25153);
nand U26200 (N_26200,N_24334,N_25604);
nand U26201 (N_26201,N_24331,N_24034);
nand U26202 (N_26202,N_25946,N_24226);
xor U26203 (N_26203,N_24781,N_24283);
nor U26204 (N_26204,N_24888,N_24027);
nand U26205 (N_26205,N_25173,N_25065);
xnor U26206 (N_26206,N_25209,N_25399);
or U26207 (N_26207,N_25202,N_25367);
and U26208 (N_26208,N_25603,N_24846);
xor U26209 (N_26209,N_25643,N_25131);
nor U26210 (N_26210,N_25268,N_24880);
or U26211 (N_26211,N_25868,N_24858);
nor U26212 (N_26212,N_25521,N_25812);
xor U26213 (N_26213,N_24702,N_24795);
and U26214 (N_26214,N_24480,N_24161);
or U26215 (N_26215,N_24414,N_25572);
and U26216 (N_26216,N_25745,N_25849);
or U26217 (N_26217,N_25345,N_25968);
or U26218 (N_26218,N_24157,N_25291);
and U26219 (N_26219,N_24873,N_24083);
nor U26220 (N_26220,N_25709,N_24665);
or U26221 (N_26221,N_24757,N_25105);
or U26222 (N_26222,N_24916,N_25705);
nand U26223 (N_26223,N_24108,N_25648);
or U26224 (N_26224,N_25664,N_25398);
or U26225 (N_26225,N_25657,N_24219);
and U26226 (N_26226,N_25773,N_25456);
or U26227 (N_26227,N_25821,N_25725);
or U26228 (N_26228,N_24973,N_24900);
nand U26229 (N_26229,N_24355,N_25368);
nor U26230 (N_26230,N_24475,N_25798);
and U26231 (N_26231,N_24547,N_25930);
nand U26232 (N_26232,N_25598,N_25840);
or U26233 (N_26233,N_24251,N_24596);
or U26234 (N_26234,N_24736,N_25138);
xnor U26235 (N_26235,N_24635,N_25302);
xor U26236 (N_26236,N_25763,N_25650);
nor U26237 (N_26237,N_25471,N_25170);
and U26238 (N_26238,N_24656,N_24539);
xor U26239 (N_26239,N_25619,N_25497);
nor U26240 (N_26240,N_24269,N_24765);
nand U26241 (N_26241,N_24159,N_25831);
or U26242 (N_26242,N_25947,N_25309);
and U26243 (N_26243,N_25436,N_25317);
nor U26244 (N_26244,N_24325,N_25943);
nand U26245 (N_26245,N_25324,N_24688);
nand U26246 (N_26246,N_25994,N_25335);
nor U26247 (N_26247,N_25500,N_25466);
and U26248 (N_26248,N_25008,N_24060);
or U26249 (N_26249,N_25021,N_25890);
nor U26250 (N_26250,N_25666,N_25605);
and U26251 (N_26251,N_25396,N_24960);
and U26252 (N_26252,N_25900,N_24750);
nor U26253 (N_26253,N_25213,N_25190);
or U26254 (N_26254,N_24659,N_24440);
xor U26255 (N_26255,N_24210,N_25043);
xor U26256 (N_26256,N_25429,N_25990);
and U26257 (N_26257,N_25460,N_25577);
and U26258 (N_26258,N_25050,N_25692);
or U26259 (N_26259,N_25690,N_24978);
nor U26260 (N_26260,N_24176,N_24174);
nand U26261 (N_26261,N_25221,N_25977);
nand U26262 (N_26262,N_24419,N_25104);
xor U26263 (N_26263,N_24021,N_25472);
or U26264 (N_26264,N_24571,N_25533);
and U26265 (N_26265,N_25952,N_25703);
or U26266 (N_26266,N_25726,N_25824);
or U26267 (N_26267,N_24941,N_25668);
nor U26268 (N_26268,N_24200,N_24059);
and U26269 (N_26269,N_25119,N_24091);
xor U26270 (N_26270,N_24318,N_24853);
nor U26271 (N_26271,N_24281,N_24867);
nor U26272 (N_26272,N_25140,N_24387);
nor U26273 (N_26273,N_24538,N_25985);
nor U26274 (N_26274,N_24955,N_25319);
xnor U26275 (N_26275,N_24122,N_25079);
nor U26276 (N_26276,N_24294,N_25967);
xnor U26277 (N_26277,N_25240,N_24168);
nor U26278 (N_26278,N_24367,N_25710);
nand U26279 (N_26279,N_24023,N_24277);
xor U26280 (N_26280,N_25724,N_24831);
and U26281 (N_26281,N_25964,N_25470);
and U26282 (N_26282,N_25573,N_24407);
nor U26283 (N_26283,N_24564,N_24685);
nand U26284 (N_26284,N_24945,N_25254);
xnor U26285 (N_26285,N_25516,N_25447);
and U26286 (N_26286,N_25134,N_25185);
and U26287 (N_26287,N_25744,N_25402);
and U26288 (N_26288,N_25051,N_24928);
or U26289 (N_26289,N_25469,N_24887);
nor U26290 (N_26290,N_24692,N_25255);
xnor U26291 (N_26291,N_25256,N_25906);
or U26292 (N_26292,N_24158,N_24590);
and U26293 (N_26293,N_24837,N_25243);
and U26294 (N_26294,N_25654,N_25624);
and U26295 (N_26295,N_24057,N_24483);
nand U26296 (N_26296,N_24050,N_24698);
nand U26297 (N_26297,N_25269,N_25801);
xnor U26298 (N_26298,N_25597,N_25923);
and U26299 (N_26299,N_24810,N_24225);
nand U26300 (N_26300,N_25839,N_24607);
xor U26301 (N_26301,N_24486,N_25337);
xor U26302 (N_26302,N_24409,N_24361);
and U26303 (N_26303,N_25973,N_25549);
and U26304 (N_26304,N_24313,N_24125);
nand U26305 (N_26305,N_24583,N_24365);
or U26306 (N_26306,N_25478,N_24363);
nand U26307 (N_26307,N_24537,N_25347);
or U26308 (N_26308,N_25740,N_25778);
or U26309 (N_26309,N_25275,N_25933);
and U26310 (N_26310,N_24184,N_25247);
xor U26311 (N_26311,N_24230,N_24460);
nand U26312 (N_26312,N_25295,N_24982);
xor U26313 (N_26313,N_24330,N_25411);
xnor U26314 (N_26314,N_24072,N_25587);
or U26315 (N_26315,N_25217,N_25815);
nor U26316 (N_26316,N_24714,N_25152);
and U26317 (N_26317,N_25163,N_24191);
nand U26318 (N_26318,N_25215,N_24910);
and U26319 (N_26319,N_25855,N_24658);
nor U26320 (N_26320,N_24426,N_24213);
xor U26321 (N_26321,N_25941,N_24580);
xor U26322 (N_26322,N_25734,N_25737);
nand U26323 (N_26323,N_24934,N_25098);
nor U26324 (N_26324,N_24233,N_24731);
nand U26325 (N_26325,N_24006,N_25252);
xor U26326 (N_26326,N_25306,N_25688);
nand U26327 (N_26327,N_24907,N_24236);
nand U26328 (N_26328,N_24981,N_25109);
or U26329 (N_26329,N_25063,N_24013);
nand U26330 (N_26330,N_25177,N_24834);
or U26331 (N_26331,N_25965,N_25800);
and U26332 (N_26332,N_24504,N_24146);
and U26333 (N_26333,N_25064,N_24700);
nor U26334 (N_26334,N_25450,N_24639);
nand U26335 (N_26335,N_24348,N_25838);
or U26336 (N_26336,N_25342,N_25087);
xor U26337 (N_26337,N_25226,N_24737);
nor U26338 (N_26338,N_25499,N_25788);
nand U26339 (N_26339,N_25996,N_25708);
nand U26340 (N_26340,N_25462,N_25176);
and U26341 (N_26341,N_24287,N_25316);
or U26342 (N_26342,N_24117,N_24708);
nor U26343 (N_26343,N_25544,N_25258);
or U26344 (N_26344,N_25856,N_24570);
and U26345 (N_26345,N_24175,N_25509);
xor U26346 (N_26346,N_24142,N_24628);
and U26347 (N_26347,N_24669,N_25510);
nand U26348 (N_26348,N_25566,N_24373);
nor U26349 (N_26349,N_25633,N_24386);
nand U26350 (N_26350,N_25179,N_25804);
and U26351 (N_26351,N_24002,N_25145);
xor U26352 (N_26352,N_24138,N_24825);
nor U26353 (N_26353,N_25858,N_24478);
nand U26354 (N_26354,N_25030,N_24065);
or U26355 (N_26355,N_24534,N_24788);
nand U26356 (N_26356,N_25753,N_24771);
xnor U26357 (N_26357,N_24624,N_25283);
xor U26358 (N_26358,N_25149,N_24554);
or U26359 (N_26359,N_25477,N_24322);
or U26360 (N_26360,N_25931,N_24798);
xnor U26361 (N_26361,N_25200,N_25110);
xor U26362 (N_26362,N_24033,N_24717);
and U26363 (N_26363,N_24991,N_24048);
xor U26364 (N_26364,N_25151,N_24304);
or U26365 (N_26365,N_25101,N_25056);
and U26366 (N_26366,N_24767,N_24120);
nor U26367 (N_26367,N_24169,N_25590);
and U26368 (N_26368,N_24090,N_24497);
or U26369 (N_26369,N_25660,N_24776);
nor U26370 (N_26370,N_25139,N_24779);
nand U26371 (N_26371,N_24962,N_25876);
or U26372 (N_26372,N_25000,N_25942);
or U26373 (N_26373,N_25066,N_25078);
nand U26374 (N_26374,N_25955,N_25645);
xor U26375 (N_26375,N_24512,N_24421);
xor U26376 (N_26376,N_25918,N_25060);
xnor U26377 (N_26377,N_24282,N_24925);
nor U26378 (N_26378,N_25759,N_25340);
xor U26379 (N_26379,N_25721,N_25752);
nor U26380 (N_26380,N_24595,N_25267);
nand U26381 (N_26381,N_24682,N_24284);
and U26382 (N_26382,N_25966,N_24608);
nor U26383 (N_26383,N_25612,N_24366);
xor U26384 (N_26384,N_25891,N_24240);
nor U26385 (N_26385,N_24300,N_25926);
or U26386 (N_26386,N_25632,N_25092);
nand U26387 (N_26387,N_25949,N_24997);
nor U26388 (N_26388,N_24642,N_24604);
and U26389 (N_26389,N_25963,N_25527);
and U26390 (N_26390,N_24636,N_24239);
xnor U26391 (N_26391,N_24623,N_24773);
or U26392 (N_26392,N_24299,N_24783);
nand U26393 (N_26393,N_25257,N_25741);
xnor U26394 (N_26394,N_25899,N_25626);
nand U26395 (N_26395,N_24376,N_24118);
or U26396 (N_26396,N_25365,N_24501);
or U26397 (N_26397,N_25385,N_25728);
or U26398 (N_26398,N_24970,N_24948);
or U26399 (N_26399,N_24351,N_25672);
nor U26400 (N_26400,N_25115,N_24620);
xnor U26401 (N_26401,N_24246,N_25341);
or U26402 (N_26402,N_24223,N_25641);
and U26403 (N_26403,N_24789,N_25120);
or U26404 (N_26404,N_25610,N_24641);
xnor U26405 (N_26405,N_24524,N_25797);
nand U26406 (N_26406,N_24311,N_25532);
xor U26407 (N_26407,N_25581,N_25495);
nand U26408 (N_26408,N_25249,N_24766);
xor U26409 (N_26409,N_24883,N_24242);
or U26410 (N_26410,N_24468,N_25397);
nand U26411 (N_26411,N_24946,N_25054);
xnor U26412 (N_26412,N_24262,N_25278);
or U26413 (N_26413,N_24953,N_25729);
nor U26414 (N_26414,N_25198,N_24618);
nand U26415 (N_26415,N_25046,N_25219);
xor U26416 (N_26416,N_25156,N_25596);
nand U26417 (N_26417,N_25053,N_25860);
or U26418 (N_26418,N_24681,N_24585);
or U26419 (N_26419,N_25956,N_24866);
and U26420 (N_26420,N_25517,N_25600);
nor U26421 (N_26421,N_24143,N_24298);
and U26422 (N_26422,N_24780,N_25895);
xnor U26423 (N_26423,N_25334,N_25363);
and U26424 (N_26424,N_25793,N_25622);
or U26425 (N_26425,N_25364,N_24790);
or U26426 (N_26426,N_25579,N_25113);
and U26427 (N_26427,N_24832,N_24593);
xor U26428 (N_26428,N_24235,N_24661);
xnor U26429 (N_26429,N_25512,N_25580);
xnor U26430 (N_26430,N_24633,N_25883);
nand U26431 (N_26431,N_24958,N_25764);
xnor U26432 (N_26432,N_25454,N_24133);
nand U26433 (N_26433,N_24514,N_24805);
nand U26434 (N_26434,N_24876,N_24711);
nand U26435 (N_26435,N_25784,N_25493);
xnor U26436 (N_26436,N_25771,N_25511);
or U26437 (N_26437,N_24707,N_24012);
nor U26438 (N_26438,N_25055,N_24152);
xor U26439 (N_26439,N_24303,N_25285);
nor U26440 (N_26440,N_25559,N_24548);
and U26441 (N_26441,N_25885,N_25308);
xnor U26442 (N_26442,N_24649,N_24049);
nor U26443 (N_26443,N_25059,N_24416);
nand U26444 (N_26444,N_24182,N_25656);
xor U26445 (N_26445,N_25205,N_25787);
and U26446 (N_26446,N_25912,N_25117);
or U26447 (N_26447,N_25676,N_25575);
nand U26448 (N_26448,N_25601,N_24256);
xor U26449 (N_26449,N_25984,N_24752);
nor U26450 (N_26450,N_24276,N_24672);
or U26451 (N_26451,N_25161,N_24696);
xor U26452 (N_26452,N_24631,N_24605);
nand U26453 (N_26453,N_24101,N_25730);
and U26454 (N_26454,N_24307,N_24575);
xor U26455 (N_26455,N_25723,N_24339);
nand U26456 (N_26456,N_25699,N_24668);
or U26457 (N_26457,N_25589,N_24247);
and U26458 (N_26458,N_24446,N_24461);
or U26459 (N_26459,N_25529,N_24292);
or U26460 (N_26460,N_25220,N_25374);
xor U26461 (N_26461,N_24746,N_25372);
nor U26462 (N_26462,N_25513,N_25216);
nand U26463 (N_26463,N_24485,N_24296);
nand U26464 (N_26464,N_25100,N_24106);
nor U26465 (N_26465,N_24836,N_25158);
xor U26466 (N_26466,N_24350,N_24753);
and U26467 (N_26467,N_25250,N_25222);
or U26468 (N_26468,N_24663,N_25355);
and U26469 (N_26469,N_25028,N_24577);
nor U26470 (N_26470,N_25166,N_25044);
xnor U26471 (N_26471,N_25896,N_24878);
xor U26472 (N_26472,N_24578,N_24043);
nor U26473 (N_26473,N_24343,N_25613);
and U26474 (N_26474,N_25123,N_24341);
xor U26475 (N_26475,N_24544,N_24140);
nand U26476 (N_26476,N_24803,N_25464);
nor U26477 (N_26477,N_24085,N_25453);
and U26478 (N_26478,N_25503,N_24969);
nor U26479 (N_26479,N_24931,N_25675);
xnor U26480 (N_26480,N_24609,N_25272);
xor U26481 (N_26481,N_24715,N_24216);
or U26482 (N_26482,N_24986,N_24541);
nand U26483 (N_26483,N_24199,N_25805);
and U26484 (N_26484,N_24847,N_25430);
xnor U26485 (N_26485,N_25538,N_24229);
nand U26486 (N_26486,N_25212,N_25090);
xnor U26487 (N_26487,N_24646,N_25870);
xnor U26488 (N_26488,N_24056,N_25024);
nor U26489 (N_26489,N_25625,N_24774);
and U26490 (N_26490,N_25718,N_24908);
and U26491 (N_26491,N_24392,N_24914);
nand U26492 (N_26492,N_25606,N_24346);
and U26493 (N_26493,N_24481,N_25614);
xnor U26494 (N_26494,N_24424,N_24823);
nand U26495 (N_26495,N_25571,N_24505);
and U26496 (N_26496,N_24812,N_24134);
or U26497 (N_26497,N_25953,N_24842);
or U26498 (N_26498,N_25441,N_24987);
nand U26499 (N_26499,N_25349,N_24053);
and U26500 (N_26500,N_25681,N_25907);
nand U26501 (N_26501,N_24148,N_24431);
and U26502 (N_26502,N_25852,N_24224);
xor U26503 (N_26503,N_24912,N_24951);
and U26504 (N_26504,N_24495,N_25320);
xnor U26505 (N_26505,N_25630,N_25281);
xnor U26506 (N_26506,N_24415,N_24290);
nand U26507 (N_26507,N_24589,N_24305);
and U26508 (N_26508,N_24807,N_24451);
or U26509 (N_26509,N_24532,N_25554);
nand U26510 (N_26510,N_25843,N_25111);
and U26511 (N_26511,N_24762,N_24906);
xnor U26512 (N_26512,N_25388,N_25877);
nand U26513 (N_26513,N_25958,N_24683);
nor U26514 (N_26514,N_24337,N_24154);
nand U26515 (N_26515,N_25144,N_25449);
or U26516 (N_26516,N_24111,N_24555);
xnor U26517 (N_26517,N_24565,N_25811);
nand U26518 (N_26518,N_25662,N_24949);
xnor U26519 (N_26519,N_24008,N_25583);
nand U26520 (N_26520,N_25218,N_25251);
or U26521 (N_26521,N_24729,N_24231);
xor U26522 (N_26522,N_24885,N_24450);
nand U26523 (N_26523,N_25461,N_24288);
nand U26524 (N_26524,N_25631,N_25356);
or U26525 (N_26525,N_24775,N_25420);
and U26526 (N_26526,N_25022,N_24259);
nor U26527 (N_26527,N_25304,N_25207);
nor U26528 (N_26528,N_24250,N_25168);
xor U26529 (N_26529,N_25394,N_25864);
and U26530 (N_26530,N_25241,N_24924);
or U26531 (N_26531,N_25802,N_25978);
nand U26532 (N_26532,N_24435,N_24456);
nor U26533 (N_26533,N_25041,N_24364);
xor U26534 (N_26534,N_25307,N_24263);
xnor U26535 (N_26535,N_25379,N_24265);
or U26536 (N_26536,N_25935,N_24749);
and U26537 (N_26537,N_24438,N_25844);
or U26538 (N_26538,N_25313,N_24974);
xor U26539 (N_26539,N_25628,N_25298);
or U26540 (N_26540,N_24801,N_24833);
and U26541 (N_26541,N_24172,N_25034);
or U26542 (N_26542,N_25361,N_24965);
nor U26543 (N_26543,N_24209,N_24741);
xnor U26544 (N_26544,N_25236,N_25264);
nor U26545 (N_26545,N_24042,N_24115);
and U26546 (N_26546,N_24733,N_24112);
xnor U26547 (N_26547,N_25289,N_24562);
and U26548 (N_26548,N_24160,N_24019);
and U26549 (N_26549,N_25623,N_24028);
or U26550 (N_26550,N_25520,N_24865);
or U26551 (N_26551,N_24279,N_24838);
xor U26552 (N_26552,N_25537,N_24718);
xnor U26553 (N_26553,N_24660,N_24574);
nand U26554 (N_26554,N_24099,N_24000);
nor U26555 (N_26555,N_25203,N_25301);
nand U26556 (N_26556,N_24770,N_25862);
or U26557 (N_26557,N_25822,N_25003);
and U26558 (N_26558,N_25514,N_25889);
or U26559 (N_26559,N_24389,N_24871);
xor U26560 (N_26560,N_25186,N_24312);
and U26561 (N_26561,N_25157,N_24040);
nor U26562 (N_26562,N_25196,N_25331);
nand U26563 (N_26563,N_25103,N_24448);
xor U26564 (N_26564,N_25426,N_24835);
xnor U26565 (N_26565,N_25116,N_24132);
xnor U26566 (N_26566,N_25564,N_24748);
and U26567 (N_26567,N_25762,N_24543);
nor U26568 (N_26568,N_24856,N_25524);
and U26569 (N_26569,N_25897,N_24315);
and U26570 (N_26570,N_24509,N_24404);
xnor U26571 (N_26571,N_25754,N_24084);
or U26572 (N_26572,N_25944,N_25871);
nor U26573 (N_26573,N_24163,N_25576);
nor U26574 (N_26574,N_24881,N_24204);
or U26575 (N_26575,N_24654,N_25037);
xor U26576 (N_26576,N_24248,N_24124);
nor U26577 (N_26577,N_25981,N_24679);
nand U26578 (N_26578,N_24884,N_24257);
and U26579 (N_26579,N_24976,N_25950);
or U26580 (N_26580,N_24519,N_24425);
or U26581 (N_26581,N_25325,N_25817);
xor U26582 (N_26582,N_24933,N_25409);
and U26583 (N_26583,N_24632,N_25794);
nor U26584 (N_26584,N_25989,N_24484);
nor U26585 (N_26585,N_24358,N_24309);
nor U26586 (N_26586,N_24098,N_24728);
and U26587 (N_26587,N_25983,N_24727);
xnor U26588 (N_26588,N_24342,N_25414);
or U26589 (N_26589,N_25481,N_24954);
xor U26590 (N_26590,N_25832,N_25960);
and U26591 (N_26591,N_24177,N_24264);
or U26592 (N_26592,N_25574,N_25233);
nand U26593 (N_26593,N_24338,N_24270);
nor U26594 (N_26594,N_24944,N_24622);
nand U26595 (N_26595,N_24274,N_25005);
nand U26596 (N_26596,N_24740,N_24394);
xor U26597 (N_26597,N_24064,N_24913);
xnor U26598 (N_26598,N_25640,N_24520);
nand U26599 (N_26599,N_24581,N_24614);
and U26600 (N_26600,N_25940,N_25184);
xor U26601 (N_26601,N_24063,N_25188);
or U26602 (N_26602,N_24915,N_24441);
xnor U26603 (N_26603,N_24966,N_24540);
and U26604 (N_26604,N_24187,N_25265);
nand U26605 (N_26605,N_25417,N_24742);
nand U26606 (N_26606,N_25751,N_25765);
or U26607 (N_26607,N_24335,N_24503);
and U26608 (N_26608,N_25490,N_25391);
xor U26609 (N_26609,N_25679,N_24675);
and U26610 (N_26610,N_24911,N_24527);
or U26611 (N_26611,N_24651,N_25582);
xor U26612 (N_26612,N_24507,N_25167);
and U26613 (N_26613,N_24652,N_24511);
nor U26614 (N_26614,N_25400,N_24479);
nor U26615 (N_26615,N_25147,N_24751);
and U26616 (N_26616,N_24897,N_24455);
xor U26617 (N_26617,N_24390,N_25318);
or U26618 (N_26618,N_24476,N_24498);
nor U26619 (N_26619,N_25586,N_25181);
nand U26620 (N_26620,N_24860,N_24020);
nor U26621 (N_26621,N_25816,N_25540);
or U26622 (N_26622,N_24588,N_25025);
and U26623 (N_26623,N_24694,N_24759);
nor U26624 (N_26624,N_25790,N_24080);
nor U26625 (N_26625,N_25659,N_24127);
or U26626 (N_26626,N_24546,N_24680);
and U26627 (N_26627,N_24678,N_24428);
and U26628 (N_26628,N_25616,N_24984);
xnor U26629 (N_26629,N_25986,N_25133);
xor U26630 (N_26630,N_25792,N_25339);
nand U26631 (N_26631,N_24137,N_25194);
and U26632 (N_26632,N_25343,N_24237);
or U26633 (N_26633,N_24600,N_25694);
and U26634 (N_26634,N_24826,N_25175);
or U26635 (N_26635,N_24324,N_24886);
nand U26636 (N_26636,N_24922,N_24490);
xnor U26637 (N_26637,N_24859,N_25522);
xor U26638 (N_26638,N_24075,N_24732);
or U26639 (N_26639,N_25480,N_24206);
and U26640 (N_26640,N_25836,N_25001);
nor U26641 (N_26641,N_25410,N_24830);
nand U26642 (N_26642,N_24333,N_24413);
xnor U26643 (N_26643,N_24145,N_25371);
nand U26644 (N_26644,N_25245,N_24382);
and U26645 (N_26645,N_24308,N_25348);
or U26646 (N_26646,N_25084,N_25680);
xnor U26647 (N_26647,N_24344,N_24345);
xnor U26648 (N_26648,N_25042,N_24381);
nor U26649 (N_26649,N_24465,N_24141);
or U26650 (N_26650,N_24109,N_25808);
nor U26651 (N_26651,N_24947,N_25867);
nand U26652 (N_26652,N_25433,N_25390);
xnor U26653 (N_26653,N_24114,N_24466);
nor U26654 (N_26654,N_25518,N_25845);
nand U26655 (N_26655,N_24052,N_24268);
xor U26656 (N_26656,N_24932,N_24238);
xor U26657 (N_26657,N_24332,N_25750);
xor U26658 (N_26658,N_25948,N_24722);
nor U26659 (N_26659,N_25859,N_25438);
nand U26660 (N_26660,N_25296,N_24653);
xnor U26661 (N_26661,N_24536,N_25358);
xnor U26662 (N_26662,N_24768,N_25615);
or U26663 (N_26663,N_25484,N_25476);
or U26664 (N_26664,N_25180,N_24336);
nor U26665 (N_26665,N_25588,N_25826);
nor U26666 (N_26666,N_25160,N_24349);
nand U26667 (N_26667,N_25785,N_24123);
or U26668 (N_26668,N_24961,N_24598);
or U26669 (N_26669,N_24797,N_24062);
xor U26670 (N_26670,N_24667,N_25106);
xnor U26671 (N_26671,N_24458,N_24195);
and U26672 (N_26672,N_25048,N_24627);
nand U26673 (N_26673,N_25550,N_25114);
or U26674 (N_26674,N_25655,N_24935);
or U26675 (N_26675,N_24695,N_24150);
xor U26676 (N_26676,N_25260,N_24522);
or U26677 (N_26677,N_24418,N_25803);
xnor U26678 (N_26678,N_25020,N_25874);
or U26679 (N_26679,N_24786,N_24809);
or U26680 (N_26680,N_24551,N_25716);
or U26681 (N_26681,N_25553,N_24434);
and U26682 (N_26682,N_24249,N_24761);
or U26683 (N_26683,N_25373,N_24619);
or U26684 (N_26684,N_24328,N_25300);
nand U26685 (N_26685,N_25957,N_24353);
nor U26686 (N_26686,N_24890,N_24340);
or U26687 (N_26687,N_24026,N_24273);
or U26688 (N_26688,N_25432,N_25758);
nand U26689 (N_26689,N_24879,N_25206);
xnor U26690 (N_26690,N_25351,N_25155);
nand U26691 (N_26691,N_24186,N_25841);
and U26692 (N_26692,N_24077,N_25881);
or U26693 (N_26693,N_24179,N_24995);
and U26694 (N_26694,N_25421,N_24178);
and U26695 (N_26695,N_24025,N_25129);
and U26696 (N_26696,N_24601,N_25594);
nor U26697 (N_26697,N_24804,N_24808);
and U26698 (N_26698,N_25828,N_24457);
or U26699 (N_26699,N_24926,N_25091);
nor U26700 (N_26700,N_25714,N_25727);
or U26701 (N_26701,N_24611,N_25061);
or U26702 (N_26702,N_24756,N_24844);
and U26703 (N_26703,N_24869,N_24074);
xor U26704 (N_26704,N_25665,N_25118);
and U26705 (N_26705,N_24500,N_25127);
and U26706 (N_26706,N_25519,N_24726);
and U26707 (N_26707,N_25536,N_25380);
or U26708 (N_26708,N_24621,N_25621);
and U26709 (N_26709,N_25068,N_24929);
xor U26710 (N_26710,N_24467,N_25818);
and U26711 (N_26711,N_24244,N_25928);
nor U26712 (N_26712,N_24131,N_24896);
and U26713 (N_26713,N_25711,N_24515);
nand U26714 (N_26714,N_24558,N_25336);
and U26715 (N_26715,N_25381,N_24243);
nand U26716 (N_26716,N_24234,N_24829);
nand U26717 (N_26717,N_24513,N_25921);
nand U26718 (N_26718,N_25154,N_24894);
or U26719 (N_26719,N_25076,N_24203);
nand U26720 (N_26720,N_24447,N_24508);
and U26721 (N_26721,N_25642,N_24968);
nand U26722 (N_26722,N_25924,N_25070);
nand U26723 (N_26723,N_25669,N_25440);
and U26724 (N_26724,N_24650,N_24067);
xnor U26725 (N_26725,N_24375,N_24716);
xnor U26726 (N_26726,N_25338,N_25378);
nor U26727 (N_26727,N_25122,N_25565);
xnor U26728 (N_26728,N_25653,N_25235);
xnor U26729 (N_26729,N_24047,N_24410);
and U26730 (N_26730,N_24939,N_25543);
and U26731 (N_26731,N_24197,N_25506);
xnor U26732 (N_26732,N_25761,N_25609);
nor U26733 (N_26733,N_24817,N_24196);
xor U26734 (N_26734,N_25311,N_25887);
and U26735 (N_26735,N_24016,N_25407);
or U26736 (N_26736,N_25314,N_24899);
xnor U26737 (N_26737,N_24266,N_25174);
and U26738 (N_26738,N_25951,N_24895);
xor U26739 (N_26739,N_24725,N_25629);
nor U26740 (N_26740,N_24054,N_25684);
nand U26741 (N_26741,N_24967,N_24430);
nor U26742 (N_26742,N_24979,N_25552);
xor U26743 (N_26743,N_25617,N_25698);
xnor U26744 (N_26744,N_24730,N_25782);
or U26745 (N_26745,N_25879,N_25303);
nor U26746 (N_26746,N_24566,N_25276);
nor U26747 (N_26747,N_25305,N_24940);
nor U26748 (N_26748,N_24278,N_24102);
nand U26749 (N_26749,N_25332,N_24502);
nand U26750 (N_26750,N_25383,N_24745);
nand U26751 (N_26751,N_24999,N_25894);
nor U26752 (N_26752,N_25401,N_24412);
nor U26753 (N_26753,N_25428,N_25344);
and U26754 (N_26754,N_25297,N_24272);
or U26755 (N_26755,N_24822,N_24068);
or U26756 (N_26756,N_24491,N_25607);
xnor U26757 (N_26757,N_25489,N_24211);
and U26758 (N_26758,N_24528,N_25567);
xnor U26759 (N_26759,N_24316,N_25095);
and U26760 (N_26760,N_25261,N_24898);
xnor U26761 (N_26761,N_24921,N_25735);
nand U26762 (N_26762,N_24289,N_25393);
xnor U26763 (N_26763,N_24901,N_24193);
nand U26764 (N_26764,N_24374,N_25819);
xor U26765 (N_26765,N_24988,N_24602);
xnor U26766 (N_26766,N_25359,N_25693);
xnor U26767 (N_26767,N_25125,N_24677);
nand U26768 (N_26768,N_24606,N_24181);
or U26769 (N_26769,N_25412,N_24763);
or U26770 (N_26770,N_24723,N_24215);
nand U26771 (N_26771,N_24321,N_24439);
xor U26772 (N_26772,N_25993,N_24082);
and U26773 (N_26773,N_24557,N_25006);
nand U26774 (N_26774,N_24310,N_25294);
xnor U26775 (N_26775,N_24755,N_25781);
nor U26776 (N_26776,N_25437,N_25058);
xor U26777 (N_26777,N_25408,N_24937);
nor U26778 (N_26778,N_25673,N_24291);
and U26779 (N_26779,N_25081,N_25651);
or U26780 (N_26780,N_24794,N_25009);
or U26781 (N_26781,N_25972,N_24038);
nand U26782 (N_26782,N_25039,N_25925);
xor U26783 (N_26783,N_25492,N_25991);
xor U26784 (N_26784,N_25677,N_24086);
xnor U26785 (N_26785,N_24170,N_25479);
and U26786 (N_26786,N_24872,N_25446);
and U26787 (N_26787,N_24104,N_24030);
xnor U26788 (N_26788,N_25886,N_24371);
nand U26789 (N_26789,N_25148,N_25040);
and U26790 (N_26790,N_24800,N_24429);
or U26791 (N_26791,N_24610,N_25833);
xnor U26792 (N_26792,N_25354,N_24706);
nor U26793 (N_26793,N_25807,N_24024);
and U26794 (N_26794,N_25747,N_25713);
xnor U26795 (N_26795,N_25722,N_25775);
xor U26796 (N_26796,N_25697,N_24594);
nor U26797 (N_26797,N_24662,N_25223);
and U26798 (N_26798,N_24942,N_25884);
nor U26799 (N_26799,N_25452,N_24670);
xor U26800 (N_26800,N_25563,N_25237);
xnor U26801 (N_26801,N_24796,N_25720);
nand U26802 (N_26802,N_25107,N_25916);
nand U26803 (N_26803,N_24472,N_24721);
or U26804 (N_26804,N_25528,N_25403);
nand U26805 (N_26805,N_24629,N_25353);
nand U26806 (N_26806,N_24093,N_24516);
or U26807 (N_26807,N_24044,N_24840);
nand U26808 (N_26808,N_25253,N_25701);
xnor U26809 (N_26809,N_25424,N_25370);
xnor U26810 (N_26810,N_24462,N_25017);
or U26811 (N_26811,N_25018,N_25435);
nor U26812 (N_26812,N_24643,N_25866);
xnor U26813 (N_26813,N_25731,N_24360);
or U26814 (N_26814,N_25569,N_24764);
or U26815 (N_26815,N_24395,N_25696);
nand U26816 (N_26816,N_25704,N_25238);
nor U26817 (N_26817,N_24096,N_24320);
and U26818 (N_26818,N_25636,N_25755);
xor U26819 (N_26819,N_25135,N_25760);
xnor U26820 (N_26820,N_24192,N_25504);
xnor U26821 (N_26821,N_24645,N_25779);
nand U26822 (N_26822,N_25873,N_25663);
or U26823 (N_26823,N_24045,N_24459);
nand U26824 (N_26824,N_24471,N_25715);
nor U26825 (N_26825,N_24442,N_25277);
and U26826 (N_26826,N_25047,N_25323);
nor U26827 (N_26827,N_25938,N_24088);
nand U26828 (N_26828,N_25945,N_24738);
and U26829 (N_26829,N_25830,N_25998);
nor U26830 (N_26830,N_24874,N_25644);
xor U26831 (N_26831,N_25049,N_25502);
or U26832 (N_26832,N_25901,N_25999);
nand U26833 (N_26833,N_24144,N_24772);
xor U26834 (N_26834,N_25230,N_24841);
and U26835 (N_26835,N_24569,N_25263);
xor U26836 (N_26836,N_25333,N_24097);
and U26837 (N_26837,N_25465,N_24634);
or U26838 (N_26838,N_25608,N_24902);
xnor U26839 (N_26839,N_25982,N_25850);
xnor U26840 (N_26840,N_24035,N_24207);
and U26841 (N_26841,N_24379,N_24323);
nand U26842 (N_26842,N_25766,N_24004);
nand U26843 (N_26843,N_25227,N_24584);
xnor U26844 (N_26844,N_24760,N_25494);
nor U26845 (N_26845,N_25089,N_24703);
nor U26846 (N_26846,N_25485,N_24037);
or U26847 (N_26847,N_25611,N_24655);
xnor U26848 (N_26848,N_24983,N_25707);
xor U26849 (N_26849,N_24518,N_25097);
xnor U26850 (N_26850,N_24362,N_25482);
and U26851 (N_26851,N_25228,N_25685);
nand U26852 (N_26852,N_25496,N_24022);
nand U26853 (N_26853,N_24396,N_24529);
nand U26854 (N_26854,N_25142,N_24356);
and U26855 (N_26855,N_24699,N_25975);
nand U26856 (N_26856,N_25086,N_25377);
nand U26857 (N_26857,N_24579,N_24103);
or U26858 (N_26858,N_25474,N_25293);
or U26859 (N_26859,N_25674,N_24676);
xnor U26860 (N_26860,N_24684,N_25108);
and U26861 (N_26861,N_25649,N_24208);
nor U26862 (N_26862,N_24496,N_25687);
nor U26863 (N_26863,N_25232,N_25002);
xnor U26864 (N_26864,N_25004,N_25282);
nor U26865 (N_26865,N_24010,N_24559);
xnor U26866 (N_26866,N_24372,N_24782);
xor U26867 (N_26867,N_24359,N_25769);
or U26868 (N_26868,N_24561,N_25419);
or U26869 (N_26869,N_24549,N_24816);
and U26870 (N_26870,N_25193,N_25892);
and U26871 (N_26871,N_24815,N_25920);
nor U26872 (N_26872,N_25067,N_24806);
xor U26873 (N_26873,N_24119,N_25733);
or U26874 (N_26874,N_25585,N_24039);
and U26875 (N_26875,N_25661,N_25702);
xnor U26876 (N_26876,N_24423,N_24850);
nor U26877 (N_26877,N_24701,N_25893);
nor U26878 (N_26878,N_25970,N_25229);
xor U26879 (N_26879,N_25266,N_25210);
or U26880 (N_26880,N_24552,N_25195);
or U26881 (N_26881,N_24255,N_24139);
nand U26882 (N_26882,N_24889,N_25491);
xnor U26883 (N_26883,N_24201,N_24422);
or U26884 (N_26884,N_25534,N_24354);
nor U26885 (N_26885,N_24556,N_25224);
nor U26886 (N_26886,N_25225,N_24843);
or U26887 (N_26887,N_24166,N_24637);
xnor U26888 (N_26888,N_24521,N_24205);
and U26889 (N_26889,N_25033,N_25757);
nand U26890 (N_26890,N_24001,N_24228);
xnor U26891 (N_26891,N_25445,N_24464);
and U26892 (N_26892,N_25683,N_25878);
nand U26893 (N_26893,N_25813,N_24417);
and U26894 (N_26894,N_25211,N_25717);
nand U26895 (N_26895,N_25169,N_25635);
and U26896 (N_26896,N_24882,N_24811);
and U26897 (N_26897,N_25290,N_24293);
xor U26898 (N_26898,N_25910,N_24408);
xnor U26899 (N_26899,N_24185,N_25165);
xnor U26900 (N_26900,N_24744,N_24996);
nand U26901 (N_26901,N_25083,N_25036);
nor U26902 (N_26902,N_25468,N_25627);
nand U26903 (N_26903,N_24245,N_24704);
nor U26904 (N_26904,N_25853,N_24673);
or U26905 (N_26905,N_25647,N_24189);
nand U26906 (N_26906,N_24147,N_24031);
xor U26907 (N_26907,N_25992,N_25327);
xor U26908 (N_26908,N_24126,N_24950);
xor U26909 (N_26909,N_24136,N_25315);
nor U26910 (N_26910,N_24989,N_24563);
nand U26911 (N_26911,N_25875,N_24994);
nor U26912 (N_26912,N_24849,N_25545);
nor U26913 (N_26913,N_24998,N_25271);
and U26914 (N_26914,N_25375,N_24076);
and U26915 (N_26915,N_24171,N_25954);
or U26916 (N_26916,N_24852,N_25768);
nor U26917 (N_26917,N_25934,N_24180);
nor U26918 (N_26918,N_24089,N_24778);
or U26919 (N_26919,N_25971,N_24405);
nand U26920 (N_26920,N_25770,N_24036);
nor U26921 (N_26921,N_25234,N_25329);
or U26922 (N_26922,N_25352,N_25541);
nor U26923 (N_26923,N_24017,N_24329);
nand U26924 (N_26924,N_25244,N_25102);
xnor U26925 (N_26925,N_25979,N_24597);
or U26926 (N_26926,N_25584,N_25976);
xor U26927 (N_26927,N_25031,N_25535);
nand U26928 (N_26928,N_24713,N_25072);
xor U26929 (N_26929,N_24014,N_25959);
nor U26930 (N_26930,N_24164,N_25451);
nor U26931 (N_26931,N_24469,N_25273);
or U26932 (N_26932,N_24444,N_25415);
nand U26933 (N_26933,N_24739,N_24188);
xnor U26934 (N_26934,N_24107,N_25997);
and U26935 (N_26935,N_25457,N_24648);
and U26936 (N_26936,N_25248,N_24533);
and U26937 (N_26937,N_25011,N_25027);
xor U26938 (N_26938,N_24993,N_24156);
xnor U26939 (N_26939,N_24493,N_24007);
nor U26940 (N_26940,N_24957,N_24149);
and U26941 (N_26941,N_24743,N_24427);
xnor U26942 (N_26942,N_24893,N_25814);
xor U26943 (N_26943,N_24734,N_24854);
nor U26944 (N_26944,N_25851,N_25810);
or U26945 (N_26945,N_25431,N_24041);
nand U26946 (N_26946,N_24489,N_24198);
nand U26947 (N_26947,N_25052,N_25357);
xnor U26948 (N_26948,N_24066,N_25739);
or U26949 (N_26949,N_25620,N_24402);
xor U26950 (N_26950,N_25360,N_25405);
or U26951 (N_26951,N_25007,N_25487);
xnor U26952 (N_26952,N_24032,N_24909);
and U26953 (N_26953,N_24437,N_24280);
nand U26954 (N_26954,N_25162,N_24015);
or U26955 (N_26955,N_24029,N_24488);
nor U26956 (N_26956,N_25239,N_25279);
nand U26957 (N_26957,N_25013,N_24857);
or U26958 (N_26958,N_24630,N_24920);
nand U26959 (N_26959,N_24785,N_25846);
nand U26960 (N_26960,N_24190,N_24851);
or U26961 (N_26961,N_24799,N_25637);
and U26962 (N_26962,N_24943,N_25932);
or U26963 (N_26963,N_24443,N_24917);
xor U26964 (N_26964,N_25774,N_25905);
xnor U26965 (N_26965,N_24572,N_25560);
nor U26966 (N_26966,N_24814,N_25015);
xnor U26967 (N_26967,N_25425,N_25189);
nor U26968 (N_26968,N_24261,N_25088);
nand U26969 (N_26969,N_24691,N_24689);
nand U26970 (N_26970,N_25861,N_24712);
and U26971 (N_26971,N_25546,N_24005);
or U26972 (N_26972,N_24167,N_25459);
and U26973 (N_26973,N_24411,N_25809);
nand U26974 (N_26974,N_25442,N_24647);
nand U26975 (N_26975,N_24214,N_25562);
and U26976 (N_26976,N_25746,N_25508);
nand U26977 (N_26977,N_24952,N_24258);
or U26978 (N_26978,N_25150,N_24492);
xor U26979 (N_26979,N_25214,N_25322);
nand U26980 (N_26980,N_24870,N_24927);
nand U26981 (N_26981,N_24664,N_24347);
xor U26982 (N_26982,N_25888,N_25837);
and U26983 (N_26983,N_25525,N_25806);
xnor U26984 (N_26984,N_24221,N_24436);
and U26985 (N_26985,N_25080,N_24877);
xnor U26986 (N_26986,N_25917,N_24445);
or U26987 (N_26987,N_24820,N_24892);
and U26988 (N_26988,N_25284,N_25376);
nor U26989 (N_26989,N_24930,N_24710);
and U26990 (N_26990,N_24454,N_25082);
or U26991 (N_26991,N_24616,N_24110);
and U26992 (N_26992,N_25854,N_25467);
xnor U26993 (N_26993,N_24314,N_24377);
or U26994 (N_26994,N_25593,N_24116);
or U26995 (N_26995,N_25652,N_24582);
and U26996 (N_26996,N_25486,N_25555);
nand U26997 (N_26997,N_24510,N_25827);
nor U26998 (N_26998,N_25208,N_25312);
or U26999 (N_26999,N_24403,N_25595);
and U27000 (N_27000,N_25241,N_24446);
nor U27001 (N_27001,N_24810,N_25346);
or U27002 (N_27002,N_24643,N_25864);
xnor U27003 (N_27003,N_25262,N_24537);
nor U27004 (N_27004,N_24288,N_24502);
or U27005 (N_27005,N_24496,N_25838);
or U27006 (N_27006,N_24704,N_25805);
xor U27007 (N_27007,N_24787,N_25281);
and U27008 (N_27008,N_25433,N_24641);
nor U27009 (N_27009,N_25919,N_25953);
xnor U27010 (N_27010,N_25343,N_25170);
and U27011 (N_27011,N_24742,N_25290);
xnor U27012 (N_27012,N_24269,N_25491);
and U27013 (N_27013,N_24617,N_25270);
nand U27014 (N_27014,N_25281,N_25118);
or U27015 (N_27015,N_25635,N_25989);
xnor U27016 (N_27016,N_25027,N_24061);
nor U27017 (N_27017,N_24380,N_25558);
xor U27018 (N_27018,N_25611,N_25505);
nor U27019 (N_27019,N_24334,N_24942);
nand U27020 (N_27020,N_25109,N_25861);
xor U27021 (N_27021,N_24428,N_24454);
nor U27022 (N_27022,N_25245,N_24535);
nor U27023 (N_27023,N_24949,N_24460);
xor U27024 (N_27024,N_24281,N_24607);
nor U27025 (N_27025,N_24474,N_25263);
and U27026 (N_27026,N_25411,N_24693);
and U27027 (N_27027,N_24808,N_25812);
or U27028 (N_27028,N_24658,N_24888);
and U27029 (N_27029,N_24447,N_25131);
nand U27030 (N_27030,N_24663,N_24863);
nand U27031 (N_27031,N_24951,N_25774);
nand U27032 (N_27032,N_24686,N_24484);
nor U27033 (N_27033,N_24099,N_24414);
xor U27034 (N_27034,N_25806,N_24524);
nor U27035 (N_27035,N_25178,N_24728);
nor U27036 (N_27036,N_24046,N_24938);
and U27037 (N_27037,N_24956,N_24604);
xor U27038 (N_27038,N_25998,N_25793);
or U27039 (N_27039,N_25528,N_24610);
and U27040 (N_27040,N_25097,N_25062);
xor U27041 (N_27041,N_25476,N_25126);
or U27042 (N_27042,N_25256,N_24438);
xor U27043 (N_27043,N_24113,N_24647);
or U27044 (N_27044,N_24649,N_24670);
and U27045 (N_27045,N_24414,N_24156);
nor U27046 (N_27046,N_24510,N_24900);
xnor U27047 (N_27047,N_24424,N_24459);
nor U27048 (N_27048,N_25775,N_24603);
or U27049 (N_27049,N_24187,N_25884);
xnor U27050 (N_27050,N_25322,N_25590);
or U27051 (N_27051,N_24455,N_24979);
nor U27052 (N_27052,N_24478,N_25528);
nand U27053 (N_27053,N_24823,N_25061);
xor U27054 (N_27054,N_24099,N_25014);
nor U27055 (N_27055,N_24426,N_25905);
and U27056 (N_27056,N_25623,N_24258);
or U27057 (N_27057,N_24794,N_25467);
nand U27058 (N_27058,N_25627,N_25422);
and U27059 (N_27059,N_25682,N_24332);
nor U27060 (N_27060,N_24669,N_25233);
nor U27061 (N_27061,N_25084,N_24359);
and U27062 (N_27062,N_25898,N_24773);
nor U27063 (N_27063,N_24896,N_25429);
or U27064 (N_27064,N_25302,N_24943);
nor U27065 (N_27065,N_24305,N_24947);
nor U27066 (N_27066,N_24585,N_25258);
nor U27067 (N_27067,N_25699,N_25930);
or U27068 (N_27068,N_25814,N_24319);
xnor U27069 (N_27069,N_24793,N_25049);
xnor U27070 (N_27070,N_24761,N_25305);
or U27071 (N_27071,N_24092,N_24348);
nor U27072 (N_27072,N_25717,N_24950);
nand U27073 (N_27073,N_25362,N_25894);
xor U27074 (N_27074,N_24647,N_25944);
or U27075 (N_27075,N_24793,N_25403);
or U27076 (N_27076,N_24930,N_24954);
or U27077 (N_27077,N_24861,N_25536);
nand U27078 (N_27078,N_24108,N_24243);
and U27079 (N_27079,N_24475,N_24035);
xnor U27080 (N_27080,N_24850,N_25429);
xnor U27081 (N_27081,N_25406,N_24037);
xor U27082 (N_27082,N_24287,N_25840);
xor U27083 (N_27083,N_25794,N_25592);
nand U27084 (N_27084,N_25804,N_25262);
nor U27085 (N_27085,N_25172,N_25372);
or U27086 (N_27086,N_24383,N_25925);
or U27087 (N_27087,N_24111,N_24461);
or U27088 (N_27088,N_25733,N_25308);
nor U27089 (N_27089,N_25233,N_24736);
or U27090 (N_27090,N_25255,N_25924);
and U27091 (N_27091,N_24258,N_24937);
or U27092 (N_27092,N_25805,N_25134);
nor U27093 (N_27093,N_25226,N_24100);
and U27094 (N_27094,N_24844,N_24366);
xnor U27095 (N_27095,N_25694,N_24920);
and U27096 (N_27096,N_24071,N_25874);
xor U27097 (N_27097,N_24584,N_25826);
nand U27098 (N_27098,N_25231,N_24842);
xor U27099 (N_27099,N_24456,N_24985);
nand U27100 (N_27100,N_25433,N_24639);
xnor U27101 (N_27101,N_24588,N_24010);
nor U27102 (N_27102,N_25327,N_25019);
and U27103 (N_27103,N_24669,N_24250);
nand U27104 (N_27104,N_25746,N_25382);
xor U27105 (N_27105,N_25890,N_25953);
nand U27106 (N_27106,N_24345,N_25432);
nand U27107 (N_27107,N_24766,N_25686);
xnor U27108 (N_27108,N_24685,N_25102);
or U27109 (N_27109,N_25373,N_25351);
or U27110 (N_27110,N_24365,N_25071);
nor U27111 (N_27111,N_24571,N_24848);
xor U27112 (N_27112,N_25192,N_24872);
nand U27113 (N_27113,N_24823,N_24838);
nor U27114 (N_27114,N_24837,N_25112);
xor U27115 (N_27115,N_25026,N_25895);
nand U27116 (N_27116,N_24450,N_24249);
nor U27117 (N_27117,N_24482,N_24292);
nor U27118 (N_27118,N_25783,N_25467);
or U27119 (N_27119,N_24817,N_24394);
and U27120 (N_27120,N_24481,N_25194);
or U27121 (N_27121,N_24132,N_24294);
nor U27122 (N_27122,N_24170,N_24871);
nand U27123 (N_27123,N_24536,N_25080);
and U27124 (N_27124,N_25784,N_25160);
xnor U27125 (N_27125,N_24089,N_25200);
nand U27126 (N_27126,N_24689,N_24528);
nor U27127 (N_27127,N_24165,N_25288);
nand U27128 (N_27128,N_24641,N_25242);
and U27129 (N_27129,N_24495,N_24867);
xnor U27130 (N_27130,N_25116,N_25793);
or U27131 (N_27131,N_24949,N_24644);
nor U27132 (N_27132,N_24964,N_25292);
and U27133 (N_27133,N_24900,N_25402);
nand U27134 (N_27134,N_25666,N_24908);
and U27135 (N_27135,N_25589,N_25876);
xnor U27136 (N_27136,N_25416,N_25067);
and U27137 (N_27137,N_25436,N_25975);
and U27138 (N_27138,N_24996,N_25725);
nand U27139 (N_27139,N_24676,N_25664);
or U27140 (N_27140,N_24174,N_25331);
or U27141 (N_27141,N_25475,N_24754);
nor U27142 (N_27142,N_25230,N_25211);
and U27143 (N_27143,N_24688,N_25898);
and U27144 (N_27144,N_24843,N_25598);
or U27145 (N_27145,N_24498,N_25417);
or U27146 (N_27146,N_24837,N_25608);
or U27147 (N_27147,N_25807,N_24224);
nand U27148 (N_27148,N_24713,N_25101);
xor U27149 (N_27149,N_24953,N_24931);
xnor U27150 (N_27150,N_25005,N_24883);
and U27151 (N_27151,N_24402,N_25439);
xnor U27152 (N_27152,N_24000,N_25826);
or U27153 (N_27153,N_25777,N_25530);
nor U27154 (N_27154,N_25510,N_24666);
and U27155 (N_27155,N_24218,N_25196);
or U27156 (N_27156,N_24174,N_24895);
nand U27157 (N_27157,N_25211,N_25348);
or U27158 (N_27158,N_25279,N_25705);
xor U27159 (N_27159,N_25464,N_25489);
or U27160 (N_27160,N_25631,N_25610);
and U27161 (N_27161,N_24269,N_25487);
and U27162 (N_27162,N_24774,N_25266);
nand U27163 (N_27163,N_25324,N_24780);
xor U27164 (N_27164,N_24384,N_25076);
or U27165 (N_27165,N_25538,N_25887);
or U27166 (N_27166,N_25189,N_24880);
nor U27167 (N_27167,N_24478,N_24384);
nor U27168 (N_27168,N_24821,N_25030);
and U27169 (N_27169,N_25237,N_24086);
and U27170 (N_27170,N_25580,N_24288);
and U27171 (N_27171,N_24404,N_25456);
nor U27172 (N_27172,N_24058,N_25131);
nand U27173 (N_27173,N_24850,N_25141);
nor U27174 (N_27174,N_24234,N_25864);
or U27175 (N_27175,N_24591,N_24992);
nor U27176 (N_27176,N_24840,N_24751);
or U27177 (N_27177,N_25021,N_24756);
nand U27178 (N_27178,N_25223,N_25989);
nand U27179 (N_27179,N_25241,N_24717);
xnor U27180 (N_27180,N_24774,N_24464);
and U27181 (N_27181,N_25875,N_24825);
xor U27182 (N_27182,N_24171,N_25405);
nor U27183 (N_27183,N_25107,N_24860);
or U27184 (N_27184,N_25163,N_25384);
and U27185 (N_27185,N_24062,N_25235);
or U27186 (N_27186,N_25954,N_25759);
or U27187 (N_27187,N_25977,N_24457);
and U27188 (N_27188,N_25193,N_24043);
nand U27189 (N_27189,N_25836,N_25450);
nand U27190 (N_27190,N_24087,N_25710);
or U27191 (N_27191,N_24148,N_24695);
nor U27192 (N_27192,N_25014,N_25052);
xor U27193 (N_27193,N_25696,N_24678);
nor U27194 (N_27194,N_25601,N_24787);
and U27195 (N_27195,N_24689,N_25184);
nand U27196 (N_27196,N_25428,N_24884);
nand U27197 (N_27197,N_24376,N_25995);
and U27198 (N_27198,N_24601,N_24191);
xnor U27199 (N_27199,N_24500,N_25419);
nand U27200 (N_27200,N_25191,N_24904);
and U27201 (N_27201,N_24136,N_25379);
and U27202 (N_27202,N_24095,N_25014);
nand U27203 (N_27203,N_25621,N_24807);
nor U27204 (N_27204,N_25606,N_24951);
or U27205 (N_27205,N_24997,N_24121);
nor U27206 (N_27206,N_25258,N_24586);
nand U27207 (N_27207,N_25431,N_25356);
and U27208 (N_27208,N_24352,N_25305);
nor U27209 (N_27209,N_24387,N_25456);
or U27210 (N_27210,N_25847,N_24405);
and U27211 (N_27211,N_25366,N_25533);
nand U27212 (N_27212,N_25761,N_25039);
nor U27213 (N_27213,N_25617,N_25957);
and U27214 (N_27214,N_24465,N_25785);
and U27215 (N_27215,N_24093,N_24823);
xor U27216 (N_27216,N_24965,N_24134);
or U27217 (N_27217,N_25132,N_24067);
and U27218 (N_27218,N_25151,N_24039);
xor U27219 (N_27219,N_24607,N_25955);
and U27220 (N_27220,N_24694,N_25879);
or U27221 (N_27221,N_24072,N_25212);
and U27222 (N_27222,N_24439,N_25474);
nor U27223 (N_27223,N_25557,N_24162);
and U27224 (N_27224,N_24944,N_24984);
and U27225 (N_27225,N_25812,N_25256);
nand U27226 (N_27226,N_25846,N_25336);
xor U27227 (N_27227,N_24632,N_25047);
or U27228 (N_27228,N_25667,N_25321);
and U27229 (N_27229,N_24565,N_24636);
nand U27230 (N_27230,N_25944,N_24121);
nand U27231 (N_27231,N_25859,N_25490);
and U27232 (N_27232,N_24690,N_25431);
xor U27233 (N_27233,N_24169,N_24446);
xor U27234 (N_27234,N_24984,N_25619);
xor U27235 (N_27235,N_25384,N_25710);
nand U27236 (N_27236,N_25021,N_24897);
xnor U27237 (N_27237,N_24861,N_25224);
or U27238 (N_27238,N_24454,N_24342);
and U27239 (N_27239,N_24587,N_25814);
and U27240 (N_27240,N_24017,N_25982);
and U27241 (N_27241,N_25449,N_24086);
and U27242 (N_27242,N_25640,N_25791);
xnor U27243 (N_27243,N_25878,N_25944);
nand U27244 (N_27244,N_24792,N_24775);
xor U27245 (N_27245,N_24763,N_25718);
xnor U27246 (N_27246,N_24538,N_25466);
nor U27247 (N_27247,N_25246,N_24821);
or U27248 (N_27248,N_25101,N_25789);
or U27249 (N_27249,N_24279,N_24281);
xnor U27250 (N_27250,N_24276,N_24383);
nor U27251 (N_27251,N_24535,N_24126);
or U27252 (N_27252,N_24147,N_24069);
xnor U27253 (N_27253,N_25456,N_25797);
xnor U27254 (N_27254,N_25950,N_24529);
and U27255 (N_27255,N_24081,N_24583);
xnor U27256 (N_27256,N_25647,N_24751);
xnor U27257 (N_27257,N_24298,N_24149);
or U27258 (N_27258,N_25258,N_25889);
xor U27259 (N_27259,N_25818,N_25548);
or U27260 (N_27260,N_25983,N_24331);
nand U27261 (N_27261,N_25339,N_24818);
nand U27262 (N_27262,N_25874,N_25943);
and U27263 (N_27263,N_25023,N_24201);
or U27264 (N_27264,N_24074,N_24893);
nor U27265 (N_27265,N_25964,N_24711);
and U27266 (N_27266,N_25074,N_25214);
and U27267 (N_27267,N_25038,N_25770);
nand U27268 (N_27268,N_24155,N_24763);
or U27269 (N_27269,N_24497,N_25511);
nand U27270 (N_27270,N_24097,N_24605);
nor U27271 (N_27271,N_25632,N_24871);
or U27272 (N_27272,N_25745,N_25374);
nand U27273 (N_27273,N_24377,N_25777);
and U27274 (N_27274,N_24849,N_24050);
and U27275 (N_27275,N_24153,N_24280);
and U27276 (N_27276,N_25804,N_25539);
or U27277 (N_27277,N_24558,N_25733);
or U27278 (N_27278,N_25892,N_25882);
xnor U27279 (N_27279,N_24911,N_24496);
xnor U27280 (N_27280,N_25815,N_24201);
nand U27281 (N_27281,N_24591,N_24246);
nand U27282 (N_27282,N_24161,N_25485);
nor U27283 (N_27283,N_25744,N_24125);
xnor U27284 (N_27284,N_25674,N_25178);
nor U27285 (N_27285,N_24612,N_24786);
nand U27286 (N_27286,N_24350,N_24496);
xor U27287 (N_27287,N_24833,N_25832);
and U27288 (N_27288,N_25445,N_24917);
and U27289 (N_27289,N_25114,N_25689);
and U27290 (N_27290,N_25224,N_24784);
nand U27291 (N_27291,N_24473,N_25059);
nand U27292 (N_27292,N_25680,N_24774);
or U27293 (N_27293,N_24128,N_25100);
xor U27294 (N_27294,N_24258,N_25961);
nor U27295 (N_27295,N_25509,N_25377);
nand U27296 (N_27296,N_25308,N_25298);
nand U27297 (N_27297,N_25435,N_24167);
and U27298 (N_27298,N_25576,N_25622);
nor U27299 (N_27299,N_25570,N_25811);
nand U27300 (N_27300,N_24911,N_25900);
or U27301 (N_27301,N_24458,N_24813);
nor U27302 (N_27302,N_25945,N_24629);
xor U27303 (N_27303,N_24901,N_24293);
or U27304 (N_27304,N_24901,N_25049);
nand U27305 (N_27305,N_25106,N_24284);
and U27306 (N_27306,N_24229,N_25070);
and U27307 (N_27307,N_25327,N_25935);
nand U27308 (N_27308,N_25670,N_25906);
or U27309 (N_27309,N_24544,N_25849);
xor U27310 (N_27310,N_24478,N_25184);
and U27311 (N_27311,N_24325,N_24174);
and U27312 (N_27312,N_25536,N_25180);
and U27313 (N_27313,N_25549,N_24973);
nand U27314 (N_27314,N_25353,N_24333);
xnor U27315 (N_27315,N_24121,N_24862);
nand U27316 (N_27316,N_24947,N_25725);
nor U27317 (N_27317,N_25216,N_24276);
nand U27318 (N_27318,N_25102,N_25647);
and U27319 (N_27319,N_24105,N_24939);
and U27320 (N_27320,N_25998,N_25244);
xor U27321 (N_27321,N_25976,N_24671);
nand U27322 (N_27322,N_25793,N_24307);
nand U27323 (N_27323,N_24568,N_24623);
and U27324 (N_27324,N_24430,N_25041);
nor U27325 (N_27325,N_24154,N_24312);
nand U27326 (N_27326,N_25361,N_25666);
nor U27327 (N_27327,N_24266,N_25456);
nor U27328 (N_27328,N_25477,N_25300);
and U27329 (N_27329,N_24880,N_24555);
or U27330 (N_27330,N_24014,N_25118);
xnor U27331 (N_27331,N_25151,N_24903);
nand U27332 (N_27332,N_24391,N_25152);
nand U27333 (N_27333,N_25119,N_24760);
nor U27334 (N_27334,N_24446,N_25680);
nand U27335 (N_27335,N_25975,N_25268);
and U27336 (N_27336,N_24307,N_25051);
xnor U27337 (N_27337,N_25048,N_24295);
nor U27338 (N_27338,N_25087,N_24957);
nor U27339 (N_27339,N_25578,N_24933);
or U27340 (N_27340,N_25574,N_25187);
or U27341 (N_27341,N_25560,N_24399);
nand U27342 (N_27342,N_25098,N_25703);
xnor U27343 (N_27343,N_24576,N_25599);
and U27344 (N_27344,N_25200,N_25429);
nor U27345 (N_27345,N_24485,N_24824);
nor U27346 (N_27346,N_24862,N_24506);
nor U27347 (N_27347,N_24709,N_25328);
nand U27348 (N_27348,N_24123,N_25120);
nand U27349 (N_27349,N_25917,N_24934);
nor U27350 (N_27350,N_25231,N_25174);
xor U27351 (N_27351,N_24540,N_24158);
xnor U27352 (N_27352,N_25743,N_24777);
xor U27353 (N_27353,N_25595,N_25759);
nand U27354 (N_27354,N_25457,N_24651);
or U27355 (N_27355,N_24063,N_25097);
nand U27356 (N_27356,N_24634,N_24349);
nor U27357 (N_27357,N_24462,N_24331);
and U27358 (N_27358,N_24764,N_24303);
nand U27359 (N_27359,N_25344,N_25945);
and U27360 (N_27360,N_24489,N_25105);
xnor U27361 (N_27361,N_24653,N_24857);
or U27362 (N_27362,N_24254,N_24415);
or U27363 (N_27363,N_25101,N_25310);
or U27364 (N_27364,N_24157,N_25209);
nand U27365 (N_27365,N_25245,N_25478);
nand U27366 (N_27366,N_25537,N_24253);
xnor U27367 (N_27367,N_24544,N_25422);
nor U27368 (N_27368,N_25032,N_24239);
nand U27369 (N_27369,N_24811,N_25653);
or U27370 (N_27370,N_25993,N_25659);
nor U27371 (N_27371,N_24030,N_24864);
xnor U27372 (N_27372,N_24978,N_24697);
nand U27373 (N_27373,N_25760,N_24060);
and U27374 (N_27374,N_24610,N_25646);
nand U27375 (N_27375,N_24184,N_24461);
or U27376 (N_27376,N_24713,N_24246);
xor U27377 (N_27377,N_25177,N_24134);
nor U27378 (N_27378,N_24526,N_25147);
xor U27379 (N_27379,N_24365,N_24462);
xnor U27380 (N_27380,N_24540,N_24783);
nor U27381 (N_27381,N_24677,N_24057);
or U27382 (N_27382,N_24467,N_24836);
nor U27383 (N_27383,N_25350,N_24318);
nand U27384 (N_27384,N_24459,N_25087);
nor U27385 (N_27385,N_24657,N_24936);
or U27386 (N_27386,N_24527,N_24594);
nand U27387 (N_27387,N_25421,N_24098);
xor U27388 (N_27388,N_24353,N_25797);
nor U27389 (N_27389,N_25764,N_24913);
xor U27390 (N_27390,N_24291,N_24388);
nor U27391 (N_27391,N_24443,N_24223);
xnor U27392 (N_27392,N_24048,N_24068);
or U27393 (N_27393,N_24202,N_25894);
nand U27394 (N_27394,N_24993,N_24169);
xnor U27395 (N_27395,N_25927,N_24087);
or U27396 (N_27396,N_25365,N_25592);
xnor U27397 (N_27397,N_24129,N_24136);
nor U27398 (N_27398,N_24039,N_24786);
and U27399 (N_27399,N_24135,N_24892);
nand U27400 (N_27400,N_25968,N_24798);
or U27401 (N_27401,N_24464,N_25875);
and U27402 (N_27402,N_24283,N_25247);
xnor U27403 (N_27403,N_25643,N_25318);
and U27404 (N_27404,N_25490,N_24311);
or U27405 (N_27405,N_24211,N_24592);
xnor U27406 (N_27406,N_25033,N_24248);
nor U27407 (N_27407,N_25562,N_24794);
and U27408 (N_27408,N_25286,N_24346);
xnor U27409 (N_27409,N_24985,N_24856);
and U27410 (N_27410,N_24369,N_24586);
or U27411 (N_27411,N_24008,N_25055);
or U27412 (N_27412,N_25108,N_25886);
or U27413 (N_27413,N_25169,N_24245);
or U27414 (N_27414,N_25251,N_24413);
or U27415 (N_27415,N_25187,N_24203);
xor U27416 (N_27416,N_25659,N_24794);
nand U27417 (N_27417,N_25570,N_24260);
nor U27418 (N_27418,N_24474,N_25881);
nor U27419 (N_27419,N_24010,N_25425);
nand U27420 (N_27420,N_25414,N_25163);
and U27421 (N_27421,N_25959,N_25496);
or U27422 (N_27422,N_24156,N_24055);
or U27423 (N_27423,N_24366,N_25482);
or U27424 (N_27424,N_25109,N_25531);
or U27425 (N_27425,N_25335,N_24852);
nor U27426 (N_27426,N_24839,N_25188);
nor U27427 (N_27427,N_25935,N_24168);
and U27428 (N_27428,N_25214,N_25088);
nor U27429 (N_27429,N_24561,N_24330);
or U27430 (N_27430,N_25649,N_25387);
or U27431 (N_27431,N_25023,N_24325);
nand U27432 (N_27432,N_25563,N_24084);
nand U27433 (N_27433,N_24981,N_24861);
xnor U27434 (N_27434,N_25557,N_24392);
nand U27435 (N_27435,N_24968,N_25719);
nand U27436 (N_27436,N_25782,N_25310);
or U27437 (N_27437,N_24828,N_25254);
and U27438 (N_27438,N_25795,N_24056);
xnor U27439 (N_27439,N_25726,N_24508);
or U27440 (N_27440,N_24532,N_24519);
xnor U27441 (N_27441,N_24779,N_24601);
nor U27442 (N_27442,N_24326,N_24517);
and U27443 (N_27443,N_25056,N_24437);
or U27444 (N_27444,N_24628,N_25488);
or U27445 (N_27445,N_24156,N_25014);
and U27446 (N_27446,N_25146,N_25605);
or U27447 (N_27447,N_24846,N_25150);
nand U27448 (N_27448,N_24591,N_25878);
nor U27449 (N_27449,N_24263,N_25119);
and U27450 (N_27450,N_25285,N_24730);
or U27451 (N_27451,N_24043,N_24277);
nor U27452 (N_27452,N_24927,N_25878);
or U27453 (N_27453,N_24400,N_24632);
nand U27454 (N_27454,N_25044,N_24573);
or U27455 (N_27455,N_24401,N_25299);
and U27456 (N_27456,N_24148,N_25234);
xnor U27457 (N_27457,N_24468,N_24135);
xor U27458 (N_27458,N_25205,N_25330);
nand U27459 (N_27459,N_24530,N_25425);
or U27460 (N_27460,N_24349,N_25431);
xnor U27461 (N_27461,N_24951,N_25349);
or U27462 (N_27462,N_25057,N_24879);
nor U27463 (N_27463,N_24602,N_24231);
xnor U27464 (N_27464,N_25757,N_25514);
and U27465 (N_27465,N_24439,N_24434);
nand U27466 (N_27466,N_25515,N_25975);
xnor U27467 (N_27467,N_25521,N_25014);
xor U27468 (N_27468,N_24754,N_24181);
nand U27469 (N_27469,N_24339,N_24528);
xnor U27470 (N_27470,N_24183,N_25915);
nor U27471 (N_27471,N_25518,N_25828);
or U27472 (N_27472,N_24889,N_25892);
nand U27473 (N_27473,N_24055,N_24324);
and U27474 (N_27474,N_24800,N_25634);
and U27475 (N_27475,N_25341,N_25407);
xnor U27476 (N_27476,N_24569,N_25271);
nor U27477 (N_27477,N_24499,N_24288);
xnor U27478 (N_27478,N_24876,N_25540);
or U27479 (N_27479,N_25728,N_24248);
nor U27480 (N_27480,N_24929,N_25241);
or U27481 (N_27481,N_25382,N_25514);
and U27482 (N_27482,N_24046,N_24962);
nor U27483 (N_27483,N_25233,N_25665);
and U27484 (N_27484,N_25207,N_25603);
xor U27485 (N_27485,N_25502,N_25072);
nor U27486 (N_27486,N_25873,N_24873);
nor U27487 (N_27487,N_24815,N_24547);
nor U27488 (N_27488,N_24165,N_24102);
xor U27489 (N_27489,N_25513,N_25420);
nand U27490 (N_27490,N_24129,N_25337);
nor U27491 (N_27491,N_24345,N_25728);
or U27492 (N_27492,N_25408,N_24150);
or U27493 (N_27493,N_24904,N_25091);
xor U27494 (N_27494,N_24589,N_25542);
nand U27495 (N_27495,N_25435,N_25719);
or U27496 (N_27496,N_25009,N_24713);
or U27497 (N_27497,N_25827,N_24212);
or U27498 (N_27498,N_25780,N_25004);
or U27499 (N_27499,N_24602,N_25673);
nand U27500 (N_27500,N_24966,N_25774);
and U27501 (N_27501,N_25398,N_24437);
xnor U27502 (N_27502,N_25109,N_25556);
and U27503 (N_27503,N_25476,N_24159);
or U27504 (N_27504,N_24028,N_25556);
and U27505 (N_27505,N_25448,N_25367);
or U27506 (N_27506,N_25233,N_25872);
nor U27507 (N_27507,N_25056,N_24300);
nand U27508 (N_27508,N_25393,N_24319);
xnor U27509 (N_27509,N_25659,N_25797);
xnor U27510 (N_27510,N_24182,N_25641);
xor U27511 (N_27511,N_25507,N_24594);
nand U27512 (N_27512,N_24405,N_25308);
or U27513 (N_27513,N_25766,N_25770);
nor U27514 (N_27514,N_25769,N_24875);
or U27515 (N_27515,N_24126,N_24479);
nand U27516 (N_27516,N_25113,N_24236);
nor U27517 (N_27517,N_24921,N_25393);
or U27518 (N_27518,N_24186,N_25084);
xnor U27519 (N_27519,N_25750,N_25972);
nor U27520 (N_27520,N_24616,N_25586);
or U27521 (N_27521,N_24273,N_24802);
xor U27522 (N_27522,N_25451,N_24589);
or U27523 (N_27523,N_24456,N_24236);
and U27524 (N_27524,N_25058,N_25069);
xor U27525 (N_27525,N_25887,N_25534);
or U27526 (N_27526,N_25718,N_24657);
nor U27527 (N_27527,N_25457,N_24080);
nand U27528 (N_27528,N_25067,N_24553);
nand U27529 (N_27529,N_25174,N_24923);
and U27530 (N_27530,N_24716,N_24045);
nand U27531 (N_27531,N_24697,N_25839);
nor U27532 (N_27532,N_25335,N_24628);
or U27533 (N_27533,N_25447,N_25788);
or U27534 (N_27534,N_25735,N_24570);
nand U27535 (N_27535,N_24230,N_25296);
or U27536 (N_27536,N_25501,N_24369);
and U27537 (N_27537,N_24174,N_25715);
and U27538 (N_27538,N_25875,N_24002);
and U27539 (N_27539,N_24020,N_25293);
or U27540 (N_27540,N_24750,N_24547);
nor U27541 (N_27541,N_24419,N_24392);
or U27542 (N_27542,N_25896,N_25211);
xnor U27543 (N_27543,N_25307,N_25384);
or U27544 (N_27544,N_24762,N_24327);
or U27545 (N_27545,N_25323,N_25035);
and U27546 (N_27546,N_25909,N_25190);
nand U27547 (N_27547,N_24566,N_25034);
nand U27548 (N_27548,N_24042,N_24005);
nor U27549 (N_27549,N_24241,N_24941);
nor U27550 (N_27550,N_24382,N_24637);
xor U27551 (N_27551,N_24441,N_25358);
or U27552 (N_27552,N_25734,N_25024);
nor U27553 (N_27553,N_24236,N_24102);
and U27554 (N_27554,N_25540,N_25566);
or U27555 (N_27555,N_24780,N_25452);
or U27556 (N_27556,N_25740,N_24825);
nand U27557 (N_27557,N_25223,N_25277);
xor U27558 (N_27558,N_25710,N_25373);
nor U27559 (N_27559,N_24155,N_25539);
and U27560 (N_27560,N_25679,N_24160);
nor U27561 (N_27561,N_25321,N_25004);
xor U27562 (N_27562,N_24074,N_24436);
xor U27563 (N_27563,N_24053,N_24327);
and U27564 (N_27564,N_24735,N_25263);
and U27565 (N_27565,N_24415,N_25780);
nor U27566 (N_27566,N_24192,N_25586);
nor U27567 (N_27567,N_25355,N_24500);
or U27568 (N_27568,N_24357,N_24696);
or U27569 (N_27569,N_25657,N_25185);
xor U27570 (N_27570,N_24072,N_24366);
and U27571 (N_27571,N_25806,N_24520);
xor U27572 (N_27572,N_25311,N_25168);
nand U27573 (N_27573,N_25009,N_25549);
xnor U27574 (N_27574,N_25038,N_24652);
and U27575 (N_27575,N_24256,N_24235);
nor U27576 (N_27576,N_25311,N_25533);
xor U27577 (N_27577,N_25313,N_25138);
xor U27578 (N_27578,N_25233,N_24813);
and U27579 (N_27579,N_25815,N_25492);
or U27580 (N_27580,N_24051,N_25665);
and U27581 (N_27581,N_24825,N_24004);
xor U27582 (N_27582,N_25320,N_25425);
and U27583 (N_27583,N_25041,N_25228);
xnor U27584 (N_27584,N_25656,N_24394);
or U27585 (N_27585,N_25095,N_25228);
and U27586 (N_27586,N_25358,N_24721);
or U27587 (N_27587,N_24883,N_24359);
or U27588 (N_27588,N_24344,N_24278);
and U27589 (N_27589,N_25237,N_24573);
xnor U27590 (N_27590,N_25384,N_24205);
or U27591 (N_27591,N_24483,N_24526);
nand U27592 (N_27592,N_24532,N_25297);
and U27593 (N_27593,N_25416,N_24296);
xnor U27594 (N_27594,N_25344,N_25776);
and U27595 (N_27595,N_25032,N_24491);
nor U27596 (N_27596,N_25293,N_24177);
and U27597 (N_27597,N_25852,N_25517);
xnor U27598 (N_27598,N_25954,N_24606);
nor U27599 (N_27599,N_24106,N_24783);
or U27600 (N_27600,N_25162,N_24923);
xnor U27601 (N_27601,N_25822,N_24555);
and U27602 (N_27602,N_25254,N_24917);
nor U27603 (N_27603,N_24818,N_25967);
xnor U27604 (N_27604,N_24308,N_25509);
nor U27605 (N_27605,N_24147,N_24815);
or U27606 (N_27606,N_24644,N_25149);
xnor U27607 (N_27607,N_24748,N_24171);
nor U27608 (N_27608,N_24526,N_24656);
and U27609 (N_27609,N_24171,N_24561);
xnor U27610 (N_27610,N_24496,N_24385);
nor U27611 (N_27611,N_24325,N_25084);
xor U27612 (N_27612,N_24969,N_24372);
and U27613 (N_27613,N_25797,N_25957);
and U27614 (N_27614,N_25937,N_25985);
nand U27615 (N_27615,N_24997,N_25335);
and U27616 (N_27616,N_24792,N_24055);
or U27617 (N_27617,N_25247,N_24993);
xnor U27618 (N_27618,N_24457,N_24027);
nor U27619 (N_27619,N_24476,N_25955);
or U27620 (N_27620,N_24132,N_24164);
nand U27621 (N_27621,N_25261,N_24901);
and U27622 (N_27622,N_25204,N_24630);
and U27623 (N_27623,N_25453,N_24061);
xnor U27624 (N_27624,N_25517,N_24416);
nor U27625 (N_27625,N_25036,N_24053);
or U27626 (N_27626,N_25308,N_24417);
xnor U27627 (N_27627,N_25527,N_24120);
and U27628 (N_27628,N_25453,N_24671);
nand U27629 (N_27629,N_25928,N_24272);
or U27630 (N_27630,N_25378,N_24023);
or U27631 (N_27631,N_24177,N_25017);
and U27632 (N_27632,N_24291,N_25597);
and U27633 (N_27633,N_25901,N_25487);
nand U27634 (N_27634,N_25428,N_25463);
nor U27635 (N_27635,N_24210,N_25719);
xor U27636 (N_27636,N_25117,N_25580);
nor U27637 (N_27637,N_25285,N_25056);
nor U27638 (N_27638,N_24894,N_24608);
nor U27639 (N_27639,N_24115,N_25512);
or U27640 (N_27640,N_25445,N_25588);
nor U27641 (N_27641,N_24976,N_24756);
or U27642 (N_27642,N_24487,N_25942);
xnor U27643 (N_27643,N_24681,N_25703);
and U27644 (N_27644,N_25568,N_25969);
nand U27645 (N_27645,N_24540,N_24857);
or U27646 (N_27646,N_25490,N_24560);
nand U27647 (N_27647,N_25739,N_25465);
or U27648 (N_27648,N_24124,N_24471);
nor U27649 (N_27649,N_25666,N_25839);
xnor U27650 (N_27650,N_25545,N_24779);
or U27651 (N_27651,N_25364,N_25315);
and U27652 (N_27652,N_25061,N_24439);
xnor U27653 (N_27653,N_24075,N_24624);
or U27654 (N_27654,N_24323,N_25173);
or U27655 (N_27655,N_25559,N_25451);
nor U27656 (N_27656,N_25589,N_24505);
and U27657 (N_27657,N_24413,N_25131);
and U27658 (N_27658,N_24293,N_25221);
or U27659 (N_27659,N_25537,N_24519);
nand U27660 (N_27660,N_24598,N_25120);
and U27661 (N_27661,N_25285,N_24018);
xnor U27662 (N_27662,N_24261,N_24322);
xor U27663 (N_27663,N_24616,N_24040);
nand U27664 (N_27664,N_24461,N_25142);
and U27665 (N_27665,N_24127,N_24474);
or U27666 (N_27666,N_25185,N_25624);
nor U27667 (N_27667,N_25265,N_24205);
or U27668 (N_27668,N_24394,N_25014);
or U27669 (N_27669,N_24062,N_24003);
nand U27670 (N_27670,N_24476,N_25846);
or U27671 (N_27671,N_25709,N_25250);
and U27672 (N_27672,N_24029,N_24517);
and U27673 (N_27673,N_25771,N_24390);
nand U27674 (N_27674,N_24497,N_25574);
or U27675 (N_27675,N_24916,N_24261);
and U27676 (N_27676,N_24035,N_24405);
and U27677 (N_27677,N_25104,N_25351);
nor U27678 (N_27678,N_24189,N_25136);
and U27679 (N_27679,N_25294,N_25762);
or U27680 (N_27680,N_25004,N_24867);
nor U27681 (N_27681,N_24723,N_24812);
nand U27682 (N_27682,N_25045,N_25390);
nor U27683 (N_27683,N_25425,N_24462);
nor U27684 (N_27684,N_24015,N_25014);
xnor U27685 (N_27685,N_25284,N_24363);
and U27686 (N_27686,N_24460,N_25024);
nor U27687 (N_27687,N_24343,N_24353);
and U27688 (N_27688,N_24111,N_24142);
nand U27689 (N_27689,N_25293,N_24607);
or U27690 (N_27690,N_24862,N_24353);
nor U27691 (N_27691,N_24063,N_24739);
nand U27692 (N_27692,N_25735,N_25236);
xor U27693 (N_27693,N_24309,N_24953);
or U27694 (N_27694,N_24928,N_24134);
xnor U27695 (N_27695,N_24359,N_25409);
and U27696 (N_27696,N_25802,N_25768);
and U27697 (N_27697,N_24855,N_24713);
nand U27698 (N_27698,N_24025,N_24913);
nand U27699 (N_27699,N_24823,N_24322);
nand U27700 (N_27700,N_24149,N_24140);
nor U27701 (N_27701,N_25883,N_24827);
nor U27702 (N_27702,N_25230,N_25294);
nand U27703 (N_27703,N_25716,N_25381);
and U27704 (N_27704,N_24623,N_25302);
nor U27705 (N_27705,N_25344,N_25362);
xnor U27706 (N_27706,N_24339,N_25672);
or U27707 (N_27707,N_24438,N_25823);
or U27708 (N_27708,N_24472,N_24347);
xnor U27709 (N_27709,N_25442,N_25643);
and U27710 (N_27710,N_25899,N_24180);
xnor U27711 (N_27711,N_24657,N_24611);
or U27712 (N_27712,N_25884,N_25112);
and U27713 (N_27713,N_24509,N_25659);
or U27714 (N_27714,N_25312,N_25847);
nand U27715 (N_27715,N_25190,N_25919);
xor U27716 (N_27716,N_25214,N_24915);
nor U27717 (N_27717,N_24423,N_24362);
or U27718 (N_27718,N_24546,N_24001);
nor U27719 (N_27719,N_24330,N_25574);
or U27720 (N_27720,N_25056,N_24154);
nand U27721 (N_27721,N_24763,N_25760);
nor U27722 (N_27722,N_25233,N_25792);
nor U27723 (N_27723,N_24993,N_25819);
xnor U27724 (N_27724,N_24815,N_24297);
and U27725 (N_27725,N_24889,N_24298);
nand U27726 (N_27726,N_25236,N_24175);
nand U27727 (N_27727,N_25334,N_24387);
or U27728 (N_27728,N_24219,N_24224);
xnor U27729 (N_27729,N_24214,N_25388);
nand U27730 (N_27730,N_25406,N_24018);
xor U27731 (N_27731,N_24492,N_24093);
or U27732 (N_27732,N_25479,N_25616);
nand U27733 (N_27733,N_24298,N_25704);
nand U27734 (N_27734,N_25882,N_24391);
nor U27735 (N_27735,N_24772,N_25259);
xnor U27736 (N_27736,N_24047,N_25433);
and U27737 (N_27737,N_25589,N_25719);
xor U27738 (N_27738,N_24873,N_24092);
nand U27739 (N_27739,N_24770,N_25999);
or U27740 (N_27740,N_24146,N_25502);
nand U27741 (N_27741,N_24474,N_24850);
and U27742 (N_27742,N_25397,N_24698);
xnor U27743 (N_27743,N_24003,N_25445);
xnor U27744 (N_27744,N_24825,N_24850);
nand U27745 (N_27745,N_24782,N_25989);
nand U27746 (N_27746,N_24134,N_24278);
nor U27747 (N_27747,N_25535,N_25047);
nand U27748 (N_27748,N_24055,N_25036);
nor U27749 (N_27749,N_25648,N_25418);
or U27750 (N_27750,N_24605,N_25771);
xnor U27751 (N_27751,N_24918,N_24858);
nor U27752 (N_27752,N_24569,N_24351);
xor U27753 (N_27753,N_25798,N_24742);
nor U27754 (N_27754,N_24909,N_25779);
nand U27755 (N_27755,N_25651,N_24051);
nor U27756 (N_27756,N_25596,N_25016);
nand U27757 (N_27757,N_25557,N_24124);
nor U27758 (N_27758,N_24780,N_25905);
nor U27759 (N_27759,N_24839,N_24044);
nor U27760 (N_27760,N_25715,N_24798);
nor U27761 (N_27761,N_24960,N_25111);
and U27762 (N_27762,N_24545,N_25401);
and U27763 (N_27763,N_25290,N_25121);
nor U27764 (N_27764,N_24846,N_24381);
xor U27765 (N_27765,N_25599,N_24904);
nor U27766 (N_27766,N_24701,N_24302);
or U27767 (N_27767,N_24790,N_24518);
and U27768 (N_27768,N_25085,N_24344);
nand U27769 (N_27769,N_25382,N_25615);
or U27770 (N_27770,N_24945,N_25203);
nor U27771 (N_27771,N_24248,N_24509);
nor U27772 (N_27772,N_25257,N_25872);
and U27773 (N_27773,N_24138,N_25745);
or U27774 (N_27774,N_24061,N_25951);
or U27775 (N_27775,N_24547,N_25762);
nor U27776 (N_27776,N_25813,N_24479);
or U27777 (N_27777,N_25928,N_25620);
or U27778 (N_27778,N_25727,N_24272);
nand U27779 (N_27779,N_24929,N_24462);
or U27780 (N_27780,N_24684,N_25757);
nand U27781 (N_27781,N_24428,N_25598);
xor U27782 (N_27782,N_24498,N_25151);
nand U27783 (N_27783,N_24363,N_24283);
or U27784 (N_27784,N_24243,N_25713);
nor U27785 (N_27785,N_24797,N_25789);
xor U27786 (N_27786,N_24822,N_25966);
nor U27787 (N_27787,N_25587,N_25119);
nor U27788 (N_27788,N_24537,N_24853);
xnor U27789 (N_27789,N_24548,N_24373);
and U27790 (N_27790,N_24447,N_24881);
and U27791 (N_27791,N_25374,N_24229);
nor U27792 (N_27792,N_25262,N_25309);
or U27793 (N_27793,N_25892,N_25863);
nand U27794 (N_27794,N_25494,N_25347);
nand U27795 (N_27795,N_24262,N_24718);
and U27796 (N_27796,N_24637,N_25351);
nand U27797 (N_27797,N_25184,N_24988);
nor U27798 (N_27798,N_25423,N_25888);
nor U27799 (N_27799,N_25963,N_24616);
nor U27800 (N_27800,N_25119,N_24806);
nor U27801 (N_27801,N_24154,N_24923);
and U27802 (N_27802,N_24956,N_25334);
xor U27803 (N_27803,N_25658,N_24351);
xnor U27804 (N_27804,N_25908,N_24192);
or U27805 (N_27805,N_24746,N_25836);
nand U27806 (N_27806,N_24460,N_25243);
and U27807 (N_27807,N_25399,N_24762);
and U27808 (N_27808,N_24417,N_25670);
xnor U27809 (N_27809,N_25471,N_25354);
xor U27810 (N_27810,N_25177,N_25025);
nor U27811 (N_27811,N_25293,N_24287);
xnor U27812 (N_27812,N_25453,N_25211);
nand U27813 (N_27813,N_24954,N_25326);
nor U27814 (N_27814,N_25305,N_24830);
or U27815 (N_27815,N_25718,N_25481);
or U27816 (N_27816,N_25488,N_25640);
xnor U27817 (N_27817,N_25330,N_25179);
xnor U27818 (N_27818,N_25425,N_24488);
xor U27819 (N_27819,N_25917,N_25591);
xor U27820 (N_27820,N_24278,N_24211);
and U27821 (N_27821,N_25348,N_24319);
xor U27822 (N_27822,N_25348,N_24715);
xor U27823 (N_27823,N_24052,N_25480);
xnor U27824 (N_27824,N_24144,N_25579);
nor U27825 (N_27825,N_24383,N_24796);
or U27826 (N_27826,N_24358,N_24841);
xnor U27827 (N_27827,N_25817,N_25619);
nor U27828 (N_27828,N_24340,N_25544);
and U27829 (N_27829,N_24765,N_24846);
and U27830 (N_27830,N_24402,N_25634);
or U27831 (N_27831,N_24110,N_25689);
nand U27832 (N_27832,N_24188,N_25276);
or U27833 (N_27833,N_24449,N_24852);
or U27834 (N_27834,N_24914,N_25890);
or U27835 (N_27835,N_25353,N_24858);
nand U27836 (N_27836,N_25308,N_24589);
nand U27837 (N_27837,N_25391,N_24990);
or U27838 (N_27838,N_25754,N_25805);
and U27839 (N_27839,N_25980,N_24303);
xnor U27840 (N_27840,N_25550,N_25430);
and U27841 (N_27841,N_25916,N_25293);
xnor U27842 (N_27842,N_25454,N_24900);
nand U27843 (N_27843,N_25226,N_24801);
and U27844 (N_27844,N_24922,N_24712);
or U27845 (N_27845,N_25745,N_25764);
nor U27846 (N_27846,N_25273,N_25943);
or U27847 (N_27847,N_24335,N_24830);
or U27848 (N_27848,N_24150,N_24658);
nor U27849 (N_27849,N_24720,N_25128);
and U27850 (N_27850,N_25495,N_24784);
nand U27851 (N_27851,N_25491,N_25937);
xor U27852 (N_27852,N_25759,N_24138);
xor U27853 (N_27853,N_24613,N_24837);
nand U27854 (N_27854,N_25420,N_24730);
nand U27855 (N_27855,N_24694,N_25130);
nand U27856 (N_27856,N_25914,N_25343);
nand U27857 (N_27857,N_24410,N_25425);
xnor U27858 (N_27858,N_25648,N_25480);
and U27859 (N_27859,N_24433,N_25820);
xnor U27860 (N_27860,N_25441,N_24492);
nor U27861 (N_27861,N_25987,N_25192);
or U27862 (N_27862,N_25969,N_24019);
or U27863 (N_27863,N_24632,N_24100);
nor U27864 (N_27864,N_25329,N_24771);
and U27865 (N_27865,N_25324,N_24415);
or U27866 (N_27866,N_25883,N_24475);
or U27867 (N_27867,N_24243,N_24241);
xnor U27868 (N_27868,N_24686,N_25398);
xnor U27869 (N_27869,N_24581,N_24722);
nor U27870 (N_27870,N_24397,N_25404);
nor U27871 (N_27871,N_24420,N_25719);
nor U27872 (N_27872,N_25667,N_24527);
or U27873 (N_27873,N_24858,N_25174);
or U27874 (N_27874,N_25240,N_24926);
nand U27875 (N_27875,N_24433,N_24613);
nand U27876 (N_27876,N_24969,N_25154);
and U27877 (N_27877,N_24115,N_24706);
xor U27878 (N_27878,N_24571,N_24390);
and U27879 (N_27879,N_24726,N_25888);
and U27880 (N_27880,N_25025,N_25751);
xor U27881 (N_27881,N_25845,N_25169);
and U27882 (N_27882,N_25730,N_24700);
nor U27883 (N_27883,N_24812,N_25434);
nand U27884 (N_27884,N_25349,N_24819);
nor U27885 (N_27885,N_24066,N_25381);
nand U27886 (N_27886,N_24772,N_24767);
or U27887 (N_27887,N_25927,N_24532);
xor U27888 (N_27888,N_25986,N_25187);
and U27889 (N_27889,N_24279,N_25607);
nor U27890 (N_27890,N_25519,N_24862);
xnor U27891 (N_27891,N_25164,N_25201);
xor U27892 (N_27892,N_25811,N_25818);
nor U27893 (N_27893,N_25574,N_25760);
nor U27894 (N_27894,N_24103,N_24923);
or U27895 (N_27895,N_24920,N_25288);
nor U27896 (N_27896,N_24633,N_24338);
and U27897 (N_27897,N_24786,N_24193);
nor U27898 (N_27898,N_24858,N_25895);
nand U27899 (N_27899,N_24027,N_25249);
xor U27900 (N_27900,N_25411,N_25226);
nand U27901 (N_27901,N_24559,N_25030);
nor U27902 (N_27902,N_25009,N_25708);
nor U27903 (N_27903,N_24403,N_24567);
nand U27904 (N_27904,N_24510,N_25863);
nor U27905 (N_27905,N_24722,N_24743);
nor U27906 (N_27906,N_24533,N_24307);
xor U27907 (N_27907,N_24800,N_25756);
or U27908 (N_27908,N_24054,N_24485);
or U27909 (N_27909,N_24857,N_25160);
or U27910 (N_27910,N_24616,N_24924);
nand U27911 (N_27911,N_25169,N_24557);
nor U27912 (N_27912,N_25620,N_24613);
nor U27913 (N_27913,N_24934,N_24277);
or U27914 (N_27914,N_24983,N_24036);
nor U27915 (N_27915,N_25205,N_24985);
nor U27916 (N_27916,N_25951,N_25058);
nand U27917 (N_27917,N_25546,N_25564);
xnor U27918 (N_27918,N_24803,N_25846);
or U27919 (N_27919,N_24290,N_25379);
nand U27920 (N_27920,N_25998,N_25938);
nor U27921 (N_27921,N_25229,N_24678);
and U27922 (N_27922,N_24113,N_25364);
or U27923 (N_27923,N_25728,N_24276);
and U27924 (N_27924,N_24677,N_25843);
or U27925 (N_27925,N_25518,N_25133);
xor U27926 (N_27926,N_24005,N_25997);
xnor U27927 (N_27927,N_25939,N_24744);
and U27928 (N_27928,N_25082,N_24017);
xor U27929 (N_27929,N_24735,N_25969);
nand U27930 (N_27930,N_25672,N_24089);
or U27931 (N_27931,N_24244,N_25913);
or U27932 (N_27932,N_25473,N_24329);
nor U27933 (N_27933,N_24109,N_25505);
or U27934 (N_27934,N_25486,N_24627);
xor U27935 (N_27935,N_24446,N_25372);
nand U27936 (N_27936,N_25741,N_25021);
or U27937 (N_27937,N_25627,N_24391);
and U27938 (N_27938,N_25370,N_24657);
nor U27939 (N_27939,N_24033,N_25659);
and U27940 (N_27940,N_25315,N_25695);
nor U27941 (N_27941,N_25304,N_24158);
nand U27942 (N_27942,N_24756,N_24092);
nor U27943 (N_27943,N_25008,N_24842);
nand U27944 (N_27944,N_25188,N_24158);
nor U27945 (N_27945,N_24909,N_25821);
nand U27946 (N_27946,N_24735,N_25131);
nor U27947 (N_27947,N_24791,N_24568);
nand U27948 (N_27948,N_25755,N_25892);
nand U27949 (N_27949,N_24386,N_25686);
xor U27950 (N_27950,N_25802,N_25051);
or U27951 (N_27951,N_25913,N_24792);
nor U27952 (N_27952,N_24373,N_25509);
xnor U27953 (N_27953,N_24028,N_24917);
xnor U27954 (N_27954,N_25299,N_24681);
xnor U27955 (N_27955,N_24915,N_24658);
and U27956 (N_27956,N_25036,N_25175);
xnor U27957 (N_27957,N_24399,N_24049);
xor U27958 (N_27958,N_24423,N_24654);
xnor U27959 (N_27959,N_25476,N_24263);
xor U27960 (N_27960,N_24193,N_24214);
xor U27961 (N_27961,N_24632,N_24517);
or U27962 (N_27962,N_25695,N_25446);
or U27963 (N_27963,N_24241,N_24204);
and U27964 (N_27964,N_24474,N_24649);
nor U27965 (N_27965,N_24291,N_25264);
and U27966 (N_27966,N_25493,N_24686);
xor U27967 (N_27967,N_25920,N_25209);
and U27968 (N_27968,N_25884,N_24695);
or U27969 (N_27969,N_24179,N_25327);
and U27970 (N_27970,N_24598,N_25685);
xnor U27971 (N_27971,N_24690,N_25966);
xor U27972 (N_27972,N_24789,N_25369);
or U27973 (N_27973,N_24436,N_25102);
and U27974 (N_27974,N_24174,N_25072);
nor U27975 (N_27975,N_24394,N_24349);
or U27976 (N_27976,N_24221,N_25477);
or U27977 (N_27977,N_24634,N_25793);
nor U27978 (N_27978,N_24405,N_24564);
nor U27979 (N_27979,N_24659,N_24532);
or U27980 (N_27980,N_25914,N_25457);
or U27981 (N_27981,N_25320,N_24780);
or U27982 (N_27982,N_25880,N_25486);
or U27983 (N_27983,N_24868,N_25859);
and U27984 (N_27984,N_24852,N_25643);
nor U27985 (N_27985,N_25137,N_25796);
nor U27986 (N_27986,N_24383,N_25233);
nand U27987 (N_27987,N_25334,N_25346);
or U27988 (N_27988,N_24836,N_25339);
and U27989 (N_27989,N_25830,N_24245);
nor U27990 (N_27990,N_25595,N_25764);
or U27991 (N_27991,N_25935,N_25726);
nand U27992 (N_27992,N_25016,N_24046);
xnor U27993 (N_27993,N_25659,N_25349);
nand U27994 (N_27994,N_25465,N_24212);
or U27995 (N_27995,N_24911,N_24818);
and U27996 (N_27996,N_24031,N_24593);
nand U27997 (N_27997,N_25400,N_25959);
and U27998 (N_27998,N_24919,N_24640);
nor U27999 (N_27999,N_24384,N_24189);
and U28000 (N_28000,N_26445,N_26877);
nand U28001 (N_28001,N_27422,N_27835);
nor U28002 (N_28002,N_27715,N_26959);
and U28003 (N_28003,N_27397,N_27309);
or U28004 (N_28004,N_26148,N_27563);
nand U28005 (N_28005,N_27066,N_27853);
xor U28006 (N_28006,N_27510,N_26781);
or U28007 (N_28007,N_27122,N_26462);
nor U28008 (N_28008,N_26474,N_27773);
or U28009 (N_28009,N_26788,N_26806);
nor U28010 (N_28010,N_27026,N_26897);
and U28011 (N_28011,N_27148,N_26753);
xnor U28012 (N_28012,N_27185,N_26968);
nor U28013 (N_28013,N_27249,N_27246);
xor U28014 (N_28014,N_27513,N_27906);
or U28015 (N_28015,N_26096,N_27157);
and U28016 (N_28016,N_27613,N_26328);
or U28017 (N_28017,N_27478,N_27177);
nand U28018 (N_28018,N_27393,N_27031);
or U28019 (N_28019,N_26989,N_26286);
and U28020 (N_28020,N_26612,N_27044);
nor U28021 (N_28021,N_26186,N_27114);
or U28022 (N_28022,N_26130,N_27860);
nand U28023 (N_28023,N_27210,N_27964);
xnor U28024 (N_28024,N_27915,N_26925);
nand U28025 (N_28025,N_27310,N_27960);
xor U28026 (N_28026,N_27271,N_26343);
nor U28027 (N_28027,N_26229,N_27356);
and U28028 (N_28028,N_26205,N_27014);
nor U28029 (N_28029,N_27149,N_26718);
or U28030 (N_28030,N_27299,N_26681);
xnor U28031 (N_28031,N_26124,N_27697);
or U28032 (N_28032,N_26540,N_27743);
nor U28033 (N_28033,N_26087,N_26036);
nor U28034 (N_28034,N_26258,N_27601);
or U28035 (N_28035,N_27805,N_27237);
nand U28036 (N_28036,N_26280,N_27129);
xor U28037 (N_28037,N_27867,N_26845);
xnor U28038 (N_28038,N_27474,N_27575);
or U28039 (N_28039,N_27671,N_27231);
nor U28040 (N_28040,N_27099,N_26583);
or U28041 (N_28041,N_26090,N_27750);
nand U28042 (N_28042,N_26011,N_26965);
nor U28043 (N_28043,N_26425,N_26434);
and U28044 (N_28044,N_26340,N_26003);
xnor U28045 (N_28045,N_26240,N_27433);
nor U28046 (N_28046,N_26828,N_27387);
nor U28047 (N_28047,N_27100,N_26610);
and U28048 (N_28048,N_26734,N_27001);
xnor U28049 (N_28049,N_26043,N_27348);
nor U28050 (N_28050,N_27038,N_26476);
nor U28051 (N_28051,N_27968,N_26482);
xnor U28052 (N_28052,N_27747,N_27887);
nor U28053 (N_28053,N_27046,N_27179);
and U28054 (N_28054,N_27234,N_26008);
and U28055 (N_28055,N_27987,N_26893);
xnor U28056 (N_28056,N_26868,N_26715);
nand U28057 (N_28057,N_27399,N_26708);
nand U28058 (N_28058,N_27439,N_26267);
nor U28059 (N_28059,N_27998,N_27574);
and U28060 (N_28060,N_27430,N_26443);
or U28061 (N_28061,N_26074,N_27219);
and U28062 (N_28062,N_26201,N_26381);
xnor U28063 (N_28063,N_27334,N_26283);
nor U28064 (N_28064,N_27751,N_26935);
nor U28065 (N_28065,N_27760,N_27701);
or U28066 (N_28066,N_27153,N_26830);
and U28067 (N_28067,N_26131,N_27625);
or U28068 (N_28068,N_26707,N_27034);
or U28069 (N_28069,N_27212,N_26969);
nand U28070 (N_28070,N_27260,N_27322);
xnor U28071 (N_28071,N_27595,N_26547);
or U28072 (N_28072,N_27783,N_26360);
nand U28073 (N_28073,N_27838,N_27244);
xor U28074 (N_28074,N_26323,N_27257);
xor U28075 (N_28075,N_27067,N_26565);
and U28076 (N_28076,N_27446,N_27349);
nor U28077 (N_28077,N_27241,N_26883);
xnor U28078 (N_28078,N_26000,N_27431);
xor U28079 (N_28079,N_26566,N_27610);
or U28080 (N_28080,N_27909,N_27208);
nor U28081 (N_28081,N_26756,N_26878);
and U28082 (N_28082,N_26232,N_26386);
nor U28083 (N_28083,N_27343,N_26084);
xor U28084 (N_28084,N_27297,N_27593);
nor U28085 (N_28085,N_26789,N_27218);
nor U28086 (N_28086,N_26651,N_26791);
xnor U28087 (N_28087,N_27500,N_27776);
nor U28088 (N_28088,N_27082,N_26932);
nand U28089 (N_28089,N_27146,N_27583);
or U28090 (N_28090,N_27460,N_26273);
and U28091 (N_28091,N_27539,N_27351);
nand U28092 (N_28092,N_27102,N_27429);
or U28093 (N_28093,N_27742,N_27920);
nor U28094 (N_28094,N_26062,N_26370);
nand U28095 (N_28095,N_26295,N_26481);
nand U28096 (N_28096,N_27159,N_27418);
xor U28097 (N_28097,N_27373,N_26355);
xnor U28098 (N_28098,N_26534,N_27354);
nor U28099 (N_28099,N_27361,N_26220);
or U28100 (N_28100,N_26032,N_27489);
xor U28101 (N_28101,N_26354,N_27767);
and U28102 (N_28102,N_26910,N_26567);
nor U28103 (N_28103,N_27139,N_26271);
xnor U28104 (N_28104,N_26486,N_27926);
xor U28105 (N_28105,N_27766,N_26636);
and U28106 (N_28106,N_27426,N_26406);
xnor U28107 (N_28107,N_27062,N_26392);
and U28108 (N_28108,N_26147,N_26326);
and U28109 (N_28109,N_27746,N_26584);
and U28110 (N_28110,N_27878,N_27344);
xnor U28111 (N_28111,N_26203,N_26721);
nand U28112 (N_28112,N_26071,N_27092);
and U28113 (N_28113,N_26782,N_26176);
nor U28114 (N_28114,N_27358,N_26168);
or U28115 (N_28115,N_27285,N_26705);
and U28116 (N_28116,N_26912,N_27629);
and U28117 (N_28117,N_27956,N_26376);
xor U28118 (N_28118,N_27719,N_26843);
nor U28119 (N_28119,N_26563,N_27874);
xnor U28120 (N_28120,N_26160,N_26711);
nand U28121 (N_28121,N_26955,N_26094);
nand U28122 (N_28122,N_27190,N_27499);
nand U28123 (N_28123,N_27480,N_27068);
nand U28124 (N_28124,N_26654,N_27728);
or U28125 (N_28125,N_27947,N_27768);
nand U28126 (N_28126,N_26512,N_27658);
or U28127 (N_28127,N_27669,N_26763);
and U28128 (N_28128,N_26377,N_26042);
nor U28129 (N_28129,N_27592,N_27880);
or U28130 (N_28130,N_26790,N_26928);
nand U28131 (N_28131,N_27134,N_27955);
nor U28132 (N_28132,N_27492,N_27705);
nand U28133 (N_28133,N_27264,N_27869);
xor U28134 (N_28134,N_26467,N_27829);
xor U28135 (N_28135,N_26680,N_26246);
nand U28136 (N_28136,N_27603,N_27895);
nand U28137 (N_28137,N_27690,N_27424);
and U28138 (N_28138,N_26259,N_26743);
nor U28139 (N_28139,N_27542,N_27732);
nand U28140 (N_28140,N_27465,N_26542);
nand U28141 (N_28141,N_27999,N_26758);
xnor U28142 (N_28142,N_27951,N_27693);
or U28143 (N_28143,N_26416,N_27990);
and U28144 (N_28144,N_26662,N_26947);
and U28145 (N_28145,N_27565,N_26757);
or U28146 (N_28146,N_26300,N_27462);
xor U28147 (N_28147,N_27367,N_27858);
nor U28148 (N_28148,N_26449,N_27982);
nand U28149 (N_28149,N_27389,N_27220);
xnor U28150 (N_28150,N_27176,N_27006);
nand U28151 (N_28151,N_26568,N_26463);
xnor U28152 (N_28152,N_27657,N_27485);
nand U28153 (N_28153,N_26159,N_27479);
and U28154 (N_28154,N_26674,N_27338);
nand U28155 (N_28155,N_26458,N_27106);
xor U28156 (N_28156,N_27084,N_27455);
and U28157 (N_28157,N_26035,N_27847);
nor U28158 (N_28158,N_26344,N_26930);
xor U28159 (N_28159,N_27620,N_26053);
xor U28160 (N_28160,N_26864,N_27167);
nand U28161 (N_28161,N_27833,N_26817);
xnor U28162 (N_28162,N_27073,N_26438);
or U28163 (N_28163,N_27755,N_27248);
or U28164 (N_28164,N_27702,N_26498);
nand U28165 (N_28165,N_27971,N_27546);
and U28166 (N_28166,N_27250,N_27030);
nor U28167 (N_28167,N_27741,N_27298);
and U28168 (N_28168,N_26359,N_26531);
nor U28169 (N_28169,N_27556,N_26667);
and U28170 (N_28170,N_27568,N_26092);
nand U28171 (N_28171,N_27213,N_26039);
nor U28172 (N_28172,N_26703,N_26480);
xnor U28173 (N_28173,N_26621,N_26044);
and U28174 (N_28174,N_27180,N_26504);
and U28175 (N_28175,N_26915,N_26275);
and U28176 (N_28176,N_27059,N_26155);
nor U28177 (N_28177,N_26200,N_26898);
and U28178 (N_28178,N_26493,N_26597);
xor U28179 (N_28179,N_26279,N_26793);
or U28180 (N_28180,N_27929,N_26134);
xnor U28181 (N_28181,N_26632,N_27032);
xor U28182 (N_28182,N_26018,N_26551);
nand U28183 (N_28183,N_26952,N_26061);
and U28184 (N_28184,N_26146,N_27182);
xor U28185 (N_28185,N_27127,N_27614);
nor U28186 (N_28186,N_26666,N_27681);
and U28187 (N_28187,N_27475,N_26627);
nand U28188 (N_28188,N_27726,N_26500);
nand U28189 (N_28189,N_26809,N_26937);
nor U28190 (N_28190,N_27836,N_26922);
nand U28191 (N_28191,N_27071,N_26774);
nor U28192 (N_28192,N_26050,N_27405);
nand U28193 (N_28193,N_27882,N_27470);
and U28194 (N_28194,N_26016,N_27543);
or U28195 (N_28195,N_27305,N_27989);
nor U28196 (N_28196,N_26266,N_27181);
and U28197 (N_28197,N_26799,N_27227);
nor U28198 (N_28198,N_27709,N_26872);
and U28199 (N_28199,N_26698,N_26996);
or U28200 (N_28200,N_26423,N_26101);
and U28201 (N_28201,N_27997,N_26466);
and U28202 (N_28202,N_26410,N_26293);
or U28203 (N_28203,N_27296,N_27531);
xnor U28204 (N_28204,N_27816,N_27323);
nand U28205 (N_28205,N_26330,N_27894);
and U28206 (N_28206,N_26640,N_27827);
nand U28207 (N_28207,N_27799,N_26385);
nor U28208 (N_28208,N_26759,N_27457);
or U28209 (N_28209,N_26195,N_27434);
or U28210 (N_28210,N_27937,N_27118);
and U28211 (N_28211,N_27916,N_27441);
or U28212 (N_28212,N_27598,N_26836);
nor U28213 (N_28213,N_26859,N_26388);
xor U28214 (N_28214,N_27109,N_27377);
and U28215 (N_28215,N_26499,N_26987);
xnor U28216 (N_28216,N_27022,N_27004);
xnor U28217 (N_28217,N_26901,N_27198);
nor U28218 (N_28218,N_26672,N_27163);
nand U28219 (N_28219,N_26484,N_26119);
nand U28220 (N_28220,N_27504,N_26646);
nand U28221 (N_28221,N_27792,N_27024);
or U28222 (N_28222,N_27281,N_26825);
nor U28223 (N_28223,N_26982,N_27812);
nand U28224 (N_28224,N_26037,N_26616);
or U28225 (N_28225,N_26136,N_27640);
xnor U28226 (N_28226,N_27856,N_27581);
xor U28227 (N_28227,N_26489,N_26850);
and U28228 (N_28228,N_27537,N_27722);
or U28229 (N_28229,N_27079,N_27273);
xnor U28230 (N_28230,N_26145,N_27611);
nor U28231 (N_28231,N_27846,N_26902);
xor U28232 (N_28232,N_26847,N_26807);
xnor U28233 (N_28233,N_27253,N_26615);
nand U28234 (N_28234,N_26460,N_26545);
or U28235 (N_28235,N_26879,N_27739);
xnor U28236 (N_28236,N_26737,N_26236);
and U28237 (N_28237,N_26972,N_26917);
xnor U28238 (N_28238,N_27639,N_27223);
nor U28239 (N_28239,N_27394,N_26589);
nor U28240 (N_28240,N_27015,N_27011);
nor U28241 (N_28241,N_27501,N_27184);
and U28242 (N_28242,N_26752,N_26196);
xnor U28243 (N_28243,N_26960,N_27392);
nor U28244 (N_28244,N_27570,N_26193);
nor U28245 (N_28245,N_26369,N_26170);
xnor U28246 (N_28246,N_27884,N_26181);
or U28247 (N_28247,N_27400,N_27949);
or U28248 (N_28248,N_27301,N_27085);
xor U28249 (N_28249,N_27169,N_26574);
nand U28250 (N_28250,N_27345,N_26031);
nor U28251 (N_28251,N_27141,N_26390);
nor U28252 (N_28252,N_26317,N_27514);
and U28253 (N_28253,N_26310,N_26455);
nand U28254 (N_28254,N_27516,N_27521);
nor U28255 (N_28255,N_26931,N_27395);
or U28256 (N_28256,N_27633,N_26840);
xnor U28257 (N_28257,N_26550,N_27958);
and U28258 (N_28258,N_27936,N_27498);
nand U28259 (N_28259,N_26079,N_26783);
xor U28260 (N_28260,N_26338,N_27567);
and U28261 (N_28261,N_27547,N_26361);
or U28262 (N_28262,N_27113,N_26553);
xor U28263 (N_28263,N_26052,N_26978);
and U28264 (N_28264,N_26316,N_26730);
and U28265 (N_28265,N_27165,N_26066);
or U28266 (N_28266,N_26886,N_26576);
and U28267 (N_28267,N_27137,N_27037);
nand U28268 (N_28268,N_27421,N_26284);
and U28269 (N_28269,N_27938,N_26358);
nor U28270 (N_28270,N_27682,N_27597);
or U28271 (N_28271,N_27511,N_26080);
and U28272 (N_28272,N_27186,N_27590);
nor U28273 (N_28273,N_27152,N_27854);
nor U28274 (N_28274,N_27566,N_27585);
and U28275 (N_28275,N_26800,N_27676);
nor U28276 (N_28276,N_27054,N_26573);
nand U28277 (N_28277,N_27454,N_27379);
nand U28278 (N_28278,N_26473,N_27905);
nor U28279 (N_28279,N_27764,N_26884);
nor U28280 (N_28280,N_26848,N_26736);
nand U28281 (N_28281,N_26623,N_27781);
nand U28282 (N_28282,N_27005,N_27497);
and U28283 (N_28283,N_27950,N_26860);
and U28284 (N_28284,N_26165,N_26314);
nand U28285 (N_28285,N_27381,N_26810);
nand U28286 (N_28286,N_26239,N_26287);
nor U28287 (N_28287,N_26852,N_26318);
or U28288 (N_28288,N_27060,N_26126);
nand U28289 (N_28289,N_27790,N_27840);
nand U28290 (N_28290,N_27675,N_27370);
or U28291 (N_28291,N_27052,N_26532);
xor U28292 (N_28292,N_26792,N_27941);
and U28293 (N_28293,N_26535,N_27969);
and U28294 (N_28294,N_27890,N_27228);
nand U28295 (N_28295,N_26132,N_26953);
or U28296 (N_28296,N_27268,N_27923);
nor U28297 (N_28297,N_27484,N_26645);
nor U28298 (N_28298,N_26426,N_27983);
and U28299 (N_28299,N_26391,N_27573);
and U28300 (N_28300,N_27362,N_27138);
nand U28301 (N_28301,N_27368,N_26998);
nor U28302 (N_28302,N_27612,N_26888);
nand U28303 (N_28303,N_26109,N_26522);
xor U28304 (N_28304,N_27885,N_27467);
nand U28305 (N_28305,N_26268,N_27043);
xor U28306 (N_28306,N_27528,N_26822);
or U28307 (N_28307,N_26107,N_26161);
nand U28308 (N_28308,N_26421,N_26111);
xor U28309 (N_28309,N_26453,N_27132);
or U28310 (N_28310,N_26688,N_26784);
nor U28311 (N_28311,N_27041,N_27461);
nand U28312 (N_28312,N_27155,N_26140);
xor U28313 (N_28313,N_27889,N_26143);
xor U28314 (N_28314,N_26335,N_26400);
xor U28315 (N_28315,N_26729,N_27278);
xor U28316 (N_28316,N_26188,N_27404);
nor U28317 (N_28317,N_26638,N_26536);
and U28318 (N_28318,N_26562,N_26659);
xor U28319 (N_28319,N_27631,N_27782);
nand U28320 (N_28320,N_26511,N_27339);
xnor U28321 (N_28321,N_27723,N_26502);
xnor U28322 (N_28322,N_26577,N_26521);
and U28323 (N_28323,N_26308,N_27576);
or U28324 (N_28324,N_27518,N_26228);
nor U28325 (N_28325,N_27832,N_26276);
nor U28326 (N_28326,N_26732,N_26710);
nor U28327 (N_28327,N_26065,N_26301);
nand U28328 (N_28328,N_26078,N_26857);
and U28329 (N_28329,N_27282,N_27197);
xnor U28330 (N_28330,N_27939,N_26858);
and U28331 (N_28331,N_26387,N_26961);
and U28332 (N_28332,N_27793,N_26657);
or U28333 (N_28333,N_26346,N_26320);
nand U28334 (N_28334,N_26520,N_26395);
or U28335 (N_28335,N_26802,N_27189);
xor U28336 (N_28336,N_26115,N_27666);
or U28337 (N_28337,N_26837,N_27353);
nor U28338 (N_28338,N_26975,N_26207);
and U28339 (N_28339,N_26601,N_26285);
or U28340 (N_28340,N_27689,N_26327);
and U28341 (N_28341,N_26060,N_26288);
xnor U28342 (N_28342,N_26282,N_27770);
or U28343 (N_28343,N_26614,N_27333);
xnor U28344 (N_28344,N_26076,N_27774);
nand U28345 (N_28345,N_27789,N_26905);
nor U28346 (N_28346,N_26424,N_26208);
nand U28347 (N_28347,N_26999,N_26670);
nor U28348 (N_28348,N_27493,N_26988);
and U28349 (N_28349,N_27063,N_27944);
xnor U28350 (N_28350,N_27608,N_27850);
or U28351 (N_28351,N_27116,N_26838);
and U28352 (N_28352,N_27036,N_26334);
nor U28353 (N_28353,N_26189,N_26221);
and U28354 (N_28354,N_26816,N_26834);
nand U28355 (N_28355,N_27437,N_26613);
or U28356 (N_28356,N_27679,N_26471);
nor U28357 (N_28357,N_26786,N_26908);
and U28358 (N_28358,N_27626,N_27587);
nor U28359 (N_28359,N_26517,N_26448);
xnor U28360 (N_28360,N_27131,N_27506);
or U28361 (N_28361,N_26211,N_26639);
nand U28362 (N_28362,N_27788,N_27557);
and U28363 (N_28363,N_26559,N_27488);
nor U28364 (N_28364,N_26985,N_27865);
or U28365 (N_28365,N_27327,N_26957);
and U28366 (N_28366,N_26306,N_26501);
nor U28367 (N_28367,N_26167,N_26741);
or U28368 (N_28368,N_26541,N_26948);
and U28369 (N_28369,N_26673,N_27352);
nand U28370 (N_28370,N_27105,N_26997);
and U28371 (N_28371,N_27415,N_26768);
nand U28372 (N_28372,N_26557,N_26656);
and U28373 (N_28373,N_26637,N_27900);
and U28374 (N_28374,N_27391,N_27300);
or U28375 (N_28375,N_27209,N_26095);
nand U28376 (N_28376,N_27959,N_26812);
nand U28377 (N_28377,N_26649,N_26823);
xor U28378 (N_28378,N_27976,N_26029);
xnor U28379 (N_28379,N_27125,N_27494);
xor U28380 (N_28380,N_26977,N_26856);
or U28381 (N_28381,N_27718,N_27094);
nand U28382 (N_28382,N_27205,N_27495);
and U28383 (N_28383,N_26325,N_26761);
nor U28384 (N_28384,N_26525,N_26051);
nor U28385 (N_28385,N_26098,N_26776);
nand U28386 (N_28386,N_27048,N_26184);
xnor U28387 (N_28387,N_26122,N_27380);
xnor U28388 (N_28388,N_26315,N_26655);
or U28389 (N_28389,N_26920,N_26311);
nor U28390 (N_28390,N_27730,N_27053);
nand U28391 (N_28391,N_27193,N_26669);
nor U28392 (N_28392,N_26393,N_26202);
nor U28393 (N_28393,N_26144,N_26773);
xnor U28394 (N_28394,N_27445,N_27624);
nand U28395 (N_28395,N_26581,N_27617);
nand U28396 (N_28396,N_27552,N_26139);
or U28397 (N_28397,N_27056,N_26379);
nand U28398 (N_28398,N_27808,N_27098);
and U28399 (N_28399,N_26496,N_26151);
nor U28400 (N_28400,N_27126,N_27525);
or U28401 (N_28401,N_27215,N_26881);
xor U28402 (N_28402,N_26021,N_27069);
and U28403 (N_28403,N_26345,N_26223);
nor U28404 (N_28404,N_27725,N_26077);
and U28405 (N_28405,N_27680,N_27630);
and U28406 (N_28406,N_27256,N_27924);
xnor U28407 (N_28407,N_26093,N_26477);
or U28408 (N_28408,N_26863,N_26192);
nor U28409 (N_28409,N_26336,N_27444);
or U28410 (N_28410,N_26411,N_26070);
nor U28411 (N_28411,N_27435,N_26507);
or U28412 (N_28412,N_27794,N_27688);
or U28413 (N_28413,N_27385,N_27632);
or U28414 (N_28414,N_26628,N_27178);
nor U28415 (N_28415,N_27272,N_26055);
nand U28416 (N_28416,N_27819,N_26516);
or U28417 (N_28417,N_27233,N_27440);
and U28418 (N_28418,N_26794,N_26403);
and U28419 (N_28419,N_26396,N_27883);
nor U28420 (N_28420,N_27691,N_27161);
or U28421 (N_28421,N_26875,N_27487);
nand U28422 (N_28422,N_26924,N_27810);
nor U28423 (N_28423,N_27145,N_26779);
and U28424 (N_28424,N_27450,N_27979);
or U28425 (N_28425,N_26117,N_26352);
nand U28426 (N_28426,N_26771,N_27262);
xnor U28427 (N_28427,N_26257,N_26523);
or U28428 (N_28428,N_27779,N_26608);
or U28429 (N_28429,N_27628,N_27007);
and U28430 (N_28430,N_26775,N_27913);
and U28431 (N_28431,N_27003,N_27616);
nand U28432 (N_28432,N_26088,N_27110);
or U28433 (N_28433,N_26342,N_26141);
nand U28434 (N_28434,N_27403,N_26116);
nand U28435 (N_28435,N_27117,N_26735);
nand U28436 (N_28436,N_26896,N_27226);
and U28437 (N_28437,N_27710,N_26247);
and U28438 (N_28438,N_26772,N_26938);
nand U28439 (N_28439,N_27076,N_27121);
or U28440 (N_28440,N_27384,N_27919);
or U28441 (N_28441,N_27174,N_27505);
and U28442 (N_28442,N_27436,N_26097);
or U28443 (N_28443,N_26740,N_27606);
nand U28444 (N_28444,N_26091,N_26956);
nor U28445 (N_28445,N_27191,N_26372);
xnor U28446 (N_28446,N_27622,N_27623);
and U28447 (N_28447,N_26675,N_27419);
xor U28448 (N_28448,N_27965,N_26739);
nand U28449 (N_28449,N_26465,N_26609);
and U28450 (N_28450,N_27996,N_27533);
xnor U28451 (N_28451,N_26700,N_26665);
or U28452 (N_28452,N_26652,N_26487);
nor U28453 (N_28453,N_27315,N_26227);
nor U28454 (N_28454,N_26981,N_27873);
or U28455 (N_28455,N_26544,N_26238);
nor U28456 (N_28456,N_26446,N_26394);
and U28457 (N_28457,N_27033,N_26128);
nand U28458 (N_28458,N_27822,N_26578);
xor U28459 (N_28459,N_27861,N_26028);
and U28460 (N_28460,N_26015,N_26853);
nand U28461 (N_28461,N_27265,N_26733);
xnor U28462 (N_28462,N_26951,N_27780);
or U28463 (N_28463,N_27921,N_27762);
or U28464 (N_28464,N_27655,N_27376);
and U28465 (N_28465,N_27673,N_27758);
or U28466 (N_28466,N_27229,N_27107);
xnor U28467 (N_28467,N_27599,N_27548);
and U28468 (N_28468,N_26120,N_26222);
or U28469 (N_28469,N_26983,N_26949);
or U28470 (N_28470,N_26179,N_26605);
nand U28471 (N_28471,N_27330,N_26742);
or U28472 (N_28472,N_26252,N_27796);
nand U28473 (N_28473,N_26941,N_26475);
or U28474 (N_28474,N_27571,N_26180);
nor U28475 (N_28475,N_26019,N_26766);
xor U28476 (N_28476,N_26701,N_26591);
nand U28477 (N_28477,N_27160,N_26769);
or U28478 (N_28478,N_27759,N_26683);
nand U28479 (N_28479,N_26363,N_26679);
and U28480 (N_28480,N_27569,N_27605);
nor U28481 (N_28481,N_27420,N_26023);
xor U28482 (N_28482,N_27259,N_27809);
nor U28483 (N_28483,N_26904,N_27413);
nor U28484 (N_28484,N_27269,N_26641);
xor U28485 (N_28485,N_26650,N_26682);
nor U28486 (N_28486,N_26599,N_27642);
xnor U28487 (N_28487,N_27684,N_27195);
nand U28488 (N_28488,N_26013,N_26337);
nor U28489 (N_28489,N_27000,N_27294);
and U28490 (N_28490,N_27520,N_26291);
and U28491 (N_28491,N_27509,N_27992);
and U28492 (N_28492,N_26210,N_27279);
xor U28493 (N_28493,N_26720,N_27010);
xor U28494 (N_28494,N_26405,N_27787);
xor U28495 (N_28495,N_27332,N_26006);
or U28496 (N_28496,N_26307,N_27108);
or U28497 (N_28497,N_27307,N_26592);
nor U28498 (N_28498,N_26940,N_27096);
and U28499 (N_28499,N_27660,N_27903);
nor U28500 (N_28500,N_27897,N_27328);
nor U28501 (N_28501,N_27712,N_27649);
nand U28502 (N_28502,N_26692,N_26251);
nor U28503 (N_28503,N_26281,N_27687);
nor U28504 (N_28504,N_26414,N_26243);
xnor U28505 (N_28505,N_26313,N_26341);
nand U28506 (N_28506,N_26457,N_26891);
xnor U28507 (N_28507,N_26787,N_26580);
nor U28508 (N_28508,N_26745,N_27845);
and U28509 (N_28509,N_27876,N_27245);
nand U28510 (N_28510,N_27277,N_26913);
xnor U28511 (N_28511,N_26727,N_27324);
nand U28512 (N_28512,N_27283,N_26713);
nor U28513 (N_28513,N_27991,N_26086);
or U28514 (N_28514,N_26469,N_27217);
nor U28515 (N_28515,N_27733,N_27589);
or U28516 (N_28516,N_27111,N_26492);
or U28517 (N_28517,N_26110,N_26431);
nor U28518 (N_28518,N_27409,N_27945);
nor U28519 (N_28519,N_27097,N_26112);
xnor U28520 (N_28520,N_26495,N_26933);
and U28521 (N_28521,N_26054,N_26510);
and U28522 (N_28522,N_26558,N_27600);
nor U28523 (N_28523,N_27716,N_27677);
nand U28524 (N_28524,N_27147,N_27103);
nor U28525 (N_28525,N_27172,N_26127);
xor U28526 (N_28526,N_26105,N_26461);
nor U28527 (N_28527,N_26722,N_27636);
and U28528 (N_28528,N_27995,N_27040);
nor U28529 (N_28529,N_26538,N_27962);
or U28530 (N_28530,N_26777,N_26412);
or U28531 (N_28531,N_26764,N_27242);
nand U28532 (N_28532,N_26005,N_26647);
or U28533 (N_28533,N_27318,N_27656);
nand U28534 (N_28534,N_26242,N_26447);
nor U28535 (N_28535,N_27634,N_27586);
and U28536 (N_28536,N_26269,N_26135);
nand U28537 (N_28537,N_26604,N_26030);
xor U28538 (N_28538,N_26867,N_26724);
or U28539 (N_28539,N_26818,N_26690);
nor U28540 (N_28540,N_27483,N_26009);
or U28541 (N_28541,N_27469,N_26198);
nand U28542 (N_28542,N_26040,N_27175);
and U28543 (N_28543,N_26509,N_26687);
xnor U28544 (N_28544,N_27202,N_27477);
and U28545 (N_28545,N_26150,N_26422);
nor U28546 (N_28546,N_27154,N_27641);
or U28547 (N_28547,N_26261,N_27230);
or U28548 (N_28548,N_26420,N_27232);
nor U28549 (N_28549,N_26010,N_26755);
xor U28550 (N_28550,N_26404,N_26600);
nor U28551 (N_28551,N_26709,N_26844);
nand U28552 (N_28552,N_26876,N_27088);
xor U28553 (N_28553,N_27700,N_26911);
xor U28554 (N_28554,N_27252,N_27448);
and U28555 (N_28555,N_27047,N_27021);
nand U28556 (N_28556,N_27637,N_27375);
nor U28557 (N_28557,N_27164,N_26024);
nand U28558 (N_28558,N_26375,N_26506);
and U28559 (N_28559,N_27740,N_27872);
and U28560 (N_28560,N_27667,N_27527);
nor U28561 (N_28561,N_27855,N_26428);
or U28562 (N_28562,N_26841,N_27359);
and U28563 (N_28563,N_27517,N_26045);
nand U28564 (N_28564,N_26100,N_27130);
and U28565 (N_28565,N_27466,N_27280);
and U28566 (N_28566,N_27074,N_26603);
nor U28567 (N_28567,N_26272,N_27225);
and U28568 (N_28568,N_26767,N_26149);
and U28569 (N_28569,N_26607,N_27588);
xor U28570 (N_28570,N_27862,N_26513);
nand U28571 (N_28571,N_27150,N_26870);
and U28572 (N_28572,N_26152,N_27261);
nor U28573 (N_28573,N_27553,N_26444);
xnor U28574 (N_28574,N_27841,N_27550);
nor U28575 (N_28575,N_27627,N_26570);
xnor U28576 (N_28576,N_27643,N_26046);
nand U28577 (N_28577,N_26488,N_26785);
xor U28578 (N_28578,N_26164,N_27800);
nor U28579 (N_28579,N_27240,N_27236);
nand U28580 (N_28580,N_26518,N_27144);
nor U28581 (N_28581,N_27785,N_26831);
nor U28582 (N_28582,N_26163,N_26157);
or U28583 (N_28583,N_26846,N_26923);
or U28584 (N_28584,N_26322,N_27188);
and U28585 (N_28585,N_27859,N_26209);
nand U28586 (N_28586,N_26963,N_26069);
and U28587 (N_28587,N_26177,N_27002);
nand U28588 (N_28588,N_26629,N_27018);
nor U28589 (N_28589,N_26383,N_26468);
or U28590 (N_28590,N_26572,N_26778);
nand U28591 (N_28591,N_27123,N_26224);
nand U28592 (N_28592,N_26695,N_27647);
nor U28593 (N_28593,N_26439,N_26892);
or U28594 (N_28594,N_27025,N_26751);
and U28595 (N_28595,N_26068,N_26289);
nor U28596 (N_28596,N_27491,N_27258);
and U28597 (N_28597,N_26451,N_27974);
nor U28598 (N_28598,N_27128,N_26861);
nor U28599 (N_28599,N_26699,N_27761);
and U28600 (N_28600,N_26626,N_27112);
xor U28601 (N_28601,N_26974,N_27875);
nand U28602 (N_28602,N_27798,N_26217);
xor U28603 (N_28603,N_26658,N_27519);
and U28604 (N_28604,N_26374,N_27748);
xor U28605 (N_28605,N_27757,N_27778);
nor U28606 (N_28606,N_26356,N_27287);
xnor U28607 (N_28607,N_27879,N_27866);
or U28608 (N_28608,N_27532,N_27119);
or U28609 (N_28609,N_27238,N_27686);
xor U28610 (N_28610,N_26248,N_26265);
or U28611 (N_28611,N_27911,N_27891);
and U28612 (N_28612,N_27482,N_27443);
or U28613 (N_28613,N_27863,N_26380);
or U28614 (N_28614,N_26435,N_26805);
nor U28615 (N_28615,N_26539,N_26611);
nand U28616 (N_28616,N_27035,N_27672);
xor U28617 (N_28617,N_26397,N_27591);
nor U28618 (N_28618,N_26226,N_26663);
nor U28619 (N_28619,N_27645,N_26555);
and U28620 (N_28620,N_26824,N_26027);
nand U28621 (N_28621,N_27452,N_26552);
nand U28622 (N_28622,N_26644,N_26862);
or U28623 (N_28623,N_27276,N_27828);
or U28624 (N_28624,N_26185,N_27888);
or U28625 (N_28625,N_26804,N_26102);
nor U28626 (N_28626,N_26237,N_27724);
nand U28627 (N_28627,N_27187,N_27893);
or U28628 (N_28628,N_27158,N_26382);
nor U28629 (N_28629,N_27648,N_27670);
nand U28630 (N_28630,N_27745,N_27830);
nand U28631 (N_28631,N_27411,N_26292);
xnor U28632 (N_28632,N_27042,N_27507);
xor U28633 (N_28633,N_27703,N_26219);
or U28634 (N_28634,N_27142,N_27286);
or U28635 (N_28635,N_27317,N_27662);
xor U28636 (N_28636,N_26063,N_26664);
nand U28637 (N_28637,N_27077,N_27235);
nor U28638 (N_28638,N_27151,N_27817);
or U28639 (N_28639,N_26976,N_27051);
nor U28640 (N_28640,N_26528,N_26137);
nand U28641 (N_28641,N_27562,N_26204);
nor U28642 (N_28642,N_27156,N_26661);
nor U28643 (N_28643,N_27708,N_26241);
or U28644 (N_28644,N_26433,N_27961);
nand U28645 (N_28645,N_26133,N_26971);
or U28646 (N_28646,N_27306,N_26676);
and U28647 (N_28647,N_27290,N_26012);
xor U28648 (N_28648,N_27192,N_27549);
nor U28649 (N_28649,N_27912,N_26191);
nand U28650 (N_28650,N_27975,N_26808);
nor U28651 (N_28651,N_27771,N_27699);
and U28652 (N_28652,N_27346,N_26332);
and U28653 (N_28653,N_26505,N_27200);
or U28654 (N_28654,N_26801,N_26378);
nor U28655 (N_28655,N_26014,N_27196);
nand U28656 (N_28656,N_27374,N_27486);
xnor U28657 (N_28657,N_26263,N_27239);
xor U28658 (N_28658,N_26099,N_27206);
xor U28659 (N_28659,N_27752,N_26527);
xnor U28660 (N_28660,N_26072,N_26907);
nand U28661 (N_28661,N_27057,N_26579);
nor U28662 (N_28662,N_27694,N_26253);
and U28663 (N_28663,N_27402,N_26244);
nand U28664 (N_28664,N_26854,N_27303);
and U28665 (N_28665,N_27934,N_26606);
xnor U28666 (N_28666,N_26235,N_27698);
nand U28667 (N_28667,N_26648,N_26526);
xor U28668 (N_28668,N_27529,N_27815);
or U28669 (N_28669,N_26780,N_26617);
nand U28670 (N_28670,N_26530,N_27857);
nor U28671 (N_28671,N_26712,N_27806);
or U28672 (N_28672,N_27821,N_27496);
or U28673 (N_28673,N_27320,N_27104);
nand U28674 (N_28674,N_27943,N_27319);
xor U28675 (N_28675,N_26595,N_26125);
and U28676 (N_28676,N_27247,N_27027);
xor U28677 (N_28677,N_27653,N_27363);
nand U28678 (N_28678,N_26894,N_26408);
or U28679 (N_28679,N_27058,N_26437);
xnor U28680 (N_28680,N_26255,N_26890);
or U28681 (N_28681,N_26123,N_26642);
and U28682 (N_28682,N_27985,N_27023);
nand U28683 (N_28683,N_27136,N_27843);
and U28684 (N_28684,N_27803,N_27289);
xnor U28685 (N_28685,N_27902,N_27340);
and U28686 (N_28686,N_27336,N_27335);
nor U28687 (N_28687,N_26754,N_27834);
nand U28688 (N_28688,N_26138,N_27558);
nor U28689 (N_28689,N_26821,N_27646);
and U28690 (N_28690,N_26554,N_27288);
nor U28691 (N_28691,N_26819,N_26082);
xor U28692 (N_28692,N_26885,N_27966);
nor U28693 (N_28693,N_26260,N_26934);
or U28694 (N_28694,N_26689,N_27738);
and U28695 (N_28695,N_26873,N_27901);
xor U28696 (N_28696,N_26746,N_27967);
xnor U28697 (N_28697,N_27972,N_27678);
nor U28698 (N_28698,N_26921,N_26979);
or U28699 (N_28699,N_26297,N_26294);
nor U28700 (N_28700,N_26256,N_26660);
or U28701 (N_28701,N_27090,N_26025);
nor U28702 (N_28702,N_27737,N_27851);
xnor U28703 (N_28703,N_26725,N_27207);
or U28704 (N_28704,N_27842,N_27251);
and U28705 (N_28705,N_27388,N_26059);
xor U28706 (N_28706,N_27428,N_27652);
xnor U28707 (N_28707,N_27008,N_26479);
or U28708 (N_28708,N_27824,N_27898);
and U28709 (N_28709,N_27772,N_26472);
nand U28710 (N_28710,N_26245,N_27735);
xor U28711 (N_28711,N_26067,N_26106);
xor U28712 (N_28712,N_26075,N_27089);
and U28713 (N_28713,N_26350,N_27095);
nor U28714 (N_28714,N_26409,N_27615);
nand U28715 (N_28715,N_27115,N_27093);
nor U28716 (N_28716,N_27918,N_26587);
and U28717 (N_28717,N_27341,N_26942);
xor U28718 (N_28718,N_26716,N_26643);
nor U28719 (N_28719,N_27503,N_27017);
nor U28720 (N_28720,N_27254,N_27607);
xnor U28721 (N_28721,N_27892,N_26357);
or U28722 (N_28722,N_26413,N_27984);
and U28723 (N_28723,N_26329,N_27266);
nand U28724 (N_28724,N_26142,N_26197);
xnor U28725 (N_28725,N_26696,N_27442);
and U28726 (N_28726,N_26417,N_27382);
nand U28727 (N_28727,N_27904,N_27203);
and U28728 (N_28728,N_27314,N_27534);
nand U28729 (N_28729,N_27922,N_26728);
nor U28730 (N_28730,N_27410,N_27545);
nor U28731 (N_28731,N_27535,N_26866);
or U28732 (N_28732,N_26118,N_27416);
xnor U28733 (N_28733,N_26049,N_26849);
and U28734 (N_28734,N_27848,N_27928);
and U28735 (N_28735,N_26304,N_27383);
nand U28736 (N_28736,N_26602,N_27663);
nor U28737 (N_28737,N_27049,N_26958);
xnor U28738 (N_28738,N_27933,N_26571);
and U28739 (N_28739,N_27456,N_27618);
xor U28740 (N_28740,N_27713,N_27162);
xnor U28741 (N_28741,N_27826,N_26353);
nand U28742 (N_28742,N_27120,N_27871);
and U28743 (N_28743,N_27194,N_27818);
nor U28744 (N_28744,N_26296,N_27993);
and U28745 (N_28745,N_26839,N_26490);
nor U28746 (N_28746,N_27295,N_27086);
and U28747 (N_28747,N_27449,N_27414);
and U28748 (N_28748,N_26158,N_27580);
and U28749 (N_28749,N_27061,N_27784);
nor U28750 (N_28750,N_27070,N_26685);
nand U28751 (N_28751,N_27820,N_26312);
xor U28752 (N_28752,N_26470,N_26089);
nor U28753 (N_28753,N_26367,N_26869);
or U28754 (N_28754,N_27540,N_26114);
and U28755 (N_28755,N_26929,N_26903);
xnor U28756 (N_28756,N_27133,N_27432);
and U28757 (N_28757,N_26954,N_27408);
or U28758 (N_28758,N_26693,N_27870);
or U28759 (N_28759,N_26365,N_26519);
xnor U28760 (N_28760,N_27714,N_26795);
xor U28761 (N_28761,N_26770,N_26215);
xnor U28762 (N_28762,N_26895,N_27572);
and U28763 (N_28763,N_27406,N_26440);
nor U28764 (N_28764,N_27512,N_26218);
or U28765 (N_28765,N_26731,N_27347);
and U28766 (N_28766,N_27706,N_26714);
and U28767 (N_28767,N_27378,N_27211);
nor U28768 (N_28768,N_27201,N_26653);
or U28769 (N_28769,N_26366,N_27777);
nor U28770 (N_28770,N_27554,N_26832);
nand U28771 (N_28771,N_26169,N_26033);
nor U28772 (N_28772,N_26004,N_27515);
or U28773 (N_28773,N_27963,N_26491);
or U28774 (N_28774,N_26058,N_27577);
or U28775 (N_28775,N_26129,N_26214);
or U28776 (N_28776,N_27736,N_27564);
or U28777 (N_28777,N_26814,N_27357);
or U28778 (N_28778,N_27644,N_27342);
xor U28779 (N_28779,N_27355,N_26225);
and U28780 (N_28780,N_26034,N_27020);
xnor U28781 (N_28781,N_26748,N_26919);
and U28782 (N_28782,N_26995,N_26633);
nand U28783 (N_28783,N_26686,N_26939);
nand U28784 (N_28784,N_27407,N_26514);
and U28785 (N_28785,N_27331,N_26351);
nor U28786 (N_28786,N_26153,N_27293);
nand U28787 (N_28787,N_27530,N_26331);
xnor U28788 (N_28788,N_27316,N_27243);
or U28789 (N_28789,N_26865,N_26212);
xnor U28790 (N_28790,N_27216,N_26277);
nor U28791 (N_28791,N_27823,N_26156);
and U28792 (N_28792,N_26719,N_26085);
nor U28793 (N_28793,N_26909,N_27311);
and U28794 (N_28794,N_27604,N_27685);
and U28795 (N_28795,N_27555,N_26017);
or U28796 (N_28796,N_27401,N_26582);
nor U28797 (N_28797,N_26803,N_26984);
xor U28798 (N_28798,N_26450,N_26993);
xor U28799 (N_28799,N_26497,N_26586);
nand U28800 (N_28800,N_26172,N_26990);
and U28801 (N_28801,N_26407,N_26162);
nor U28802 (N_28802,N_27970,N_27012);
xor U28803 (N_28803,N_26950,N_27674);
xnor U28804 (N_28804,N_26048,N_27173);
xor U28805 (N_28805,N_27325,N_27802);
xnor U28806 (N_28806,N_26270,N_26702);
or U28807 (N_28807,N_26047,N_26194);
nor U28808 (N_28808,N_27977,N_27584);
and U28809 (N_28809,N_27953,N_27453);
xor U28810 (N_28810,N_26813,N_26103);
nor U28811 (N_28811,N_26401,N_26671);
nand U28812 (N_28812,N_26593,N_26073);
xor U28813 (N_28813,N_26402,N_27930);
xor U28814 (N_28814,N_26723,N_27321);
or U28815 (N_28815,N_27124,N_27329);
and U28816 (N_28816,N_27019,N_27721);
or U28817 (N_28817,N_27490,N_26635);
xor U28818 (N_28818,N_27396,N_27813);
xnor U28819 (N_28819,N_26190,N_26081);
nor U28820 (N_28820,N_27908,N_26298);
or U28821 (N_28821,N_26362,N_27143);
or U28822 (N_28822,N_26738,N_26973);
xor U28823 (N_28823,N_27753,N_27222);
nor U28824 (N_28824,N_26432,N_27302);
nor U28825 (N_28825,N_26927,N_27825);
nor U28826 (N_28826,N_27692,N_27561);
nand U28827 (N_28827,N_26419,N_26427);
and U28828 (N_28828,N_27072,N_26305);
or U28829 (N_28829,N_26691,N_26524);
nor U28830 (N_28830,N_27602,N_26750);
or U28831 (N_28831,N_26456,N_27412);
nand U28832 (N_28832,N_27814,N_27868);
or U28833 (N_28833,N_26944,N_26827);
and U28834 (N_28834,N_27523,N_26349);
or U28835 (N_28835,N_26717,N_26945);
and U28836 (N_28836,N_27650,N_26624);
and U28837 (N_28837,N_27952,N_27508);
nor U28838 (N_28838,N_26038,N_27594);
nand U28839 (N_28839,N_26943,N_26290);
or U28840 (N_28840,N_26249,N_27274);
and U28841 (N_28841,N_26348,N_26429);
nand U28842 (N_28842,N_27801,N_27704);
nand U28843 (N_28843,N_26452,N_27769);
or U28844 (N_28844,N_27925,N_27786);
nor U28845 (N_28845,N_26026,N_26324);
or U28846 (N_28846,N_26556,N_26234);
xor U28847 (N_28847,N_27831,N_27371);
xor U28848 (N_28848,N_26598,N_27981);
or U28849 (N_28849,N_26887,N_27914);
xor U28850 (N_28850,N_27744,N_27275);
xor U28851 (N_28851,N_26561,N_27837);
nor U28852 (N_28852,N_26529,N_26418);
nor U28853 (N_28853,N_27171,N_27907);
and U28854 (N_28854,N_26002,N_27308);
and U28855 (N_28855,N_26697,N_27427);
and U28856 (N_28856,N_26684,N_26967);
or U28857 (N_28857,N_26855,N_26590);
nand U28858 (N_28858,N_26515,N_26618);
and U28859 (N_28859,N_27270,N_26765);
nor U28860 (N_28860,N_26992,N_27459);
or U28861 (N_28861,N_27864,N_27596);
nor U28862 (N_28862,N_27609,N_26900);
nor U28863 (N_28863,N_27980,N_27988);
and U28864 (N_28864,N_26970,N_26630);
and U28865 (N_28865,N_26677,N_26622);
nor U28866 (N_28866,N_27683,N_26842);
or U28867 (N_28867,N_27039,N_27524);
nand U28868 (N_28868,N_26216,N_27013);
nand U28869 (N_28869,N_26262,N_26442);
and U28870 (N_28870,N_27101,N_26104);
or U28871 (N_28871,N_26113,N_27016);
nand U28872 (N_28872,N_26811,N_27386);
or U28873 (N_28873,N_27255,N_26483);
nand U28874 (N_28874,N_27168,N_26543);
xor U28875 (N_28875,N_27973,N_26183);
or U28876 (N_28876,N_26964,N_26454);
xnor U28877 (N_28877,N_26994,N_26368);
xnor U28878 (N_28878,N_27707,N_27659);
xor U28879 (N_28879,N_27621,N_27366);
nand U28880 (N_28880,N_27791,N_27438);
nand U28881 (N_28881,N_26619,N_27417);
and U28882 (N_28882,N_27292,N_26796);
and U28883 (N_28883,N_26199,N_26064);
or U28884 (N_28884,N_27468,N_26302);
xor U28885 (N_28885,N_26347,N_27917);
xnor U28886 (N_28886,N_27886,N_26962);
and U28887 (N_28887,N_27729,N_26882);
or U28888 (N_28888,N_26001,N_27811);
nand U28889 (N_28889,N_27423,N_27204);
nor U28890 (N_28890,N_26441,N_26946);
and U28891 (N_28891,N_26020,N_27471);
or U28892 (N_28892,N_26906,N_27978);
nand U28893 (N_28893,N_27087,N_27765);
nor U28894 (N_28894,N_27224,N_26309);
or U28895 (N_28895,N_26899,N_27390);
nand U28896 (N_28896,N_27582,N_27881);
nand U28897 (N_28897,N_26250,N_27717);
nor U28898 (N_28898,N_26459,N_27221);
xor U28899 (N_28899,N_26415,N_26926);
or U28900 (N_28900,N_26254,N_27559);
xnor U28901 (N_28901,N_27065,N_26625);
and U28902 (N_28902,N_27635,N_26230);
and U28903 (N_28903,N_26620,N_27425);
or U28904 (N_28904,N_27481,N_26041);
nor U28905 (N_28905,N_26278,N_27948);
nor U28906 (N_28906,N_26373,N_27775);
nor U28907 (N_28907,N_27029,N_27910);
nand U28908 (N_28908,N_26575,N_27931);
or U28909 (N_28909,N_26634,N_27170);
nor U28910 (N_28910,N_26057,N_27551);
nand U28911 (N_28911,N_26436,N_27804);
xnor U28912 (N_28912,N_26749,N_27807);
xnor U28913 (N_28913,N_26503,N_26880);
and U28914 (N_28914,N_26007,N_27350);
or U28915 (N_28915,N_27994,N_27214);
and U28916 (N_28916,N_27078,N_27045);
or U28917 (N_28917,N_27711,N_27055);
nor U28918 (N_28918,N_27754,N_26399);
and U28919 (N_28919,N_27064,N_26747);
xor U28920 (N_28920,N_27083,N_26264);
xor U28921 (N_28921,N_26537,N_27526);
nor U28922 (N_28922,N_26083,N_27695);
and U28923 (N_28923,N_27731,N_26564);
and U28924 (N_28924,N_26121,N_26174);
nor U28925 (N_28925,N_26533,N_26588);
nand U28926 (N_28926,N_26966,N_26384);
nor U28927 (N_28927,N_27749,N_26166);
nor U28928 (N_28928,N_26319,N_26494);
nor U28929 (N_28929,N_26833,N_26171);
and U28930 (N_28930,N_27304,N_26820);
xnor U28931 (N_28931,N_27080,N_26585);
nor U28932 (N_28932,N_26549,N_27696);
or U28933 (N_28933,N_26464,N_26206);
nor U28934 (N_28934,N_27464,N_26918);
nand U28935 (N_28935,N_27476,N_27337);
xnor U28936 (N_28936,N_26678,N_27957);
xnor U28937 (N_28937,N_26815,N_27619);
xor U28938 (N_28938,N_26704,N_27291);
and U28939 (N_28939,N_26056,N_27284);
nand U28940 (N_28940,N_27756,N_26175);
nor U28941 (N_28941,N_27927,N_26914);
nor U28942 (N_28942,N_27651,N_26478);
nand U28943 (N_28943,N_26274,N_26182);
nand U28944 (N_28944,N_27654,N_27720);
xor U28945 (N_28945,N_27398,N_27940);
and U28946 (N_28946,N_26762,N_27458);
or U28947 (N_28947,N_26835,N_27665);
or U28948 (N_28948,N_26760,N_27081);
nor U28949 (N_28949,N_27727,N_26173);
and U28950 (N_28950,N_27472,N_26871);
nor U28951 (N_28951,N_27028,N_26744);
or U28952 (N_28952,N_27661,N_27183);
nor U28953 (N_28953,N_26569,N_26594);
and U28954 (N_28954,N_26916,N_27849);
xor U28955 (N_28955,N_26980,N_26022);
nand U28956 (N_28956,N_26548,N_27852);
nor U28957 (N_28957,N_27447,N_26333);
and U28958 (N_28958,N_27839,N_26797);
nand U28959 (N_28959,N_27312,N_26874);
or U28960 (N_28960,N_26299,N_27091);
and U28961 (N_28961,N_26339,N_26829);
and U28962 (N_28962,N_27009,N_26826);
and U28963 (N_28963,N_27986,N_26389);
and U28964 (N_28964,N_27544,N_26178);
xnor U28965 (N_28965,N_27896,N_27522);
nand U28966 (N_28966,N_27797,N_26364);
xnor U28967 (N_28967,N_27451,N_27541);
xor U28968 (N_28968,N_27795,N_27932);
nor U28969 (N_28969,N_27946,N_27536);
xnor U28970 (N_28970,N_27365,N_26889);
nor U28971 (N_28971,N_26321,N_27267);
and U28972 (N_28972,N_27075,N_27560);
nor U28973 (N_28973,N_27579,N_26187);
and U28974 (N_28974,N_27638,N_27463);
and U28975 (N_28975,N_26108,N_26303);
nor U28976 (N_28976,N_27140,N_26398);
nand U28977 (N_28977,N_27263,N_26726);
nand U28978 (N_28978,N_26430,N_26233);
nor U28979 (N_28979,N_27538,N_26936);
nand U28980 (N_28980,N_26560,N_26213);
nand U28981 (N_28981,N_26485,N_26371);
nor U28982 (N_28982,N_27166,N_27369);
or U28983 (N_28983,N_26508,N_27954);
xor U28984 (N_28984,N_27899,N_27668);
and U28985 (N_28985,N_27502,N_27763);
xnor U28986 (N_28986,N_26986,N_26154);
and U28987 (N_28987,N_26631,N_26668);
or U28988 (N_28988,N_26851,N_27473);
nand U28989 (N_28989,N_26546,N_26991);
or U28990 (N_28990,N_27844,N_27578);
nor U28991 (N_28991,N_27199,N_26231);
and U28992 (N_28992,N_27877,N_27135);
xor U28993 (N_28993,N_27372,N_27734);
and U28994 (N_28994,N_26706,N_26694);
nand U28995 (N_28995,N_27360,N_27050);
nand U28996 (N_28996,N_27935,N_26596);
xor U28997 (N_28997,N_27326,N_26798);
or U28998 (N_28998,N_27942,N_27313);
nand U28999 (N_28999,N_27664,N_27364);
xor U29000 (N_29000,N_27898,N_26817);
nand U29001 (N_29001,N_26216,N_26892);
nor U29002 (N_29002,N_27000,N_26755);
and U29003 (N_29003,N_27133,N_26562);
nand U29004 (N_29004,N_27353,N_26278);
and U29005 (N_29005,N_27031,N_26393);
and U29006 (N_29006,N_27402,N_26057);
and U29007 (N_29007,N_26077,N_27966);
xnor U29008 (N_29008,N_27258,N_27411);
or U29009 (N_29009,N_26085,N_26259);
xor U29010 (N_29010,N_27222,N_26194);
nand U29011 (N_29011,N_26753,N_26247);
and U29012 (N_29012,N_27246,N_27665);
or U29013 (N_29013,N_26718,N_26353);
xor U29014 (N_29014,N_27249,N_26343);
nand U29015 (N_29015,N_26633,N_27839);
xor U29016 (N_29016,N_27904,N_27091);
or U29017 (N_29017,N_26082,N_27072);
nand U29018 (N_29018,N_27371,N_27640);
xor U29019 (N_29019,N_26930,N_27683);
or U29020 (N_29020,N_27286,N_26539);
and U29021 (N_29021,N_27314,N_26730);
or U29022 (N_29022,N_26926,N_26783);
or U29023 (N_29023,N_27834,N_27853);
xnor U29024 (N_29024,N_27065,N_26553);
nand U29025 (N_29025,N_27575,N_26119);
xnor U29026 (N_29026,N_27937,N_26985);
xnor U29027 (N_29027,N_26368,N_27300);
or U29028 (N_29028,N_27020,N_26143);
and U29029 (N_29029,N_26114,N_26237);
nand U29030 (N_29030,N_26322,N_27430);
and U29031 (N_29031,N_26597,N_27474);
or U29032 (N_29032,N_27711,N_27552);
or U29033 (N_29033,N_26965,N_26661);
xor U29034 (N_29034,N_27749,N_26200);
or U29035 (N_29035,N_27992,N_26252);
nor U29036 (N_29036,N_27678,N_27880);
nand U29037 (N_29037,N_27454,N_27817);
xnor U29038 (N_29038,N_27622,N_27384);
and U29039 (N_29039,N_27583,N_26169);
xnor U29040 (N_29040,N_26370,N_27118);
or U29041 (N_29041,N_26648,N_27674);
or U29042 (N_29042,N_26425,N_27627);
and U29043 (N_29043,N_27534,N_27790);
and U29044 (N_29044,N_26985,N_26886);
xnor U29045 (N_29045,N_27153,N_26854);
or U29046 (N_29046,N_26230,N_26182);
or U29047 (N_29047,N_27542,N_26769);
or U29048 (N_29048,N_27297,N_27736);
or U29049 (N_29049,N_26595,N_27044);
or U29050 (N_29050,N_27565,N_26766);
xnor U29051 (N_29051,N_26431,N_26742);
xor U29052 (N_29052,N_26680,N_26816);
xnor U29053 (N_29053,N_27887,N_27297);
xor U29054 (N_29054,N_27932,N_27939);
xor U29055 (N_29055,N_27220,N_27330);
or U29056 (N_29056,N_26706,N_26884);
xnor U29057 (N_29057,N_27958,N_26585);
and U29058 (N_29058,N_27969,N_26643);
nand U29059 (N_29059,N_27239,N_26406);
nand U29060 (N_29060,N_27205,N_27397);
or U29061 (N_29061,N_26224,N_26646);
nand U29062 (N_29062,N_26567,N_27298);
nor U29063 (N_29063,N_26653,N_26407);
nand U29064 (N_29064,N_27789,N_27662);
or U29065 (N_29065,N_27911,N_26736);
xnor U29066 (N_29066,N_26887,N_26522);
nand U29067 (N_29067,N_26801,N_26665);
or U29068 (N_29068,N_27576,N_27555);
or U29069 (N_29069,N_26979,N_27866);
nand U29070 (N_29070,N_27269,N_27604);
xnor U29071 (N_29071,N_26199,N_27716);
nand U29072 (N_29072,N_26969,N_27071);
and U29073 (N_29073,N_26316,N_27937);
xor U29074 (N_29074,N_27246,N_26064);
nor U29075 (N_29075,N_26806,N_27727);
nor U29076 (N_29076,N_27084,N_27748);
nor U29077 (N_29077,N_26396,N_27872);
nor U29078 (N_29078,N_27936,N_27477);
xor U29079 (N_29079,N_26362,N_26782);
nand U29080 (N_29080,N_26803,N_26339);
nand U29081 (N_29081,N_26115,N_27975);
and U29082 (N_29082,N_26722,N_27029);
or U29083 (N_29083,N_26308,N_26696);
nand U29084 (N_29084,N_26153,N_27416);
nand U29085 (N_29085,N_26282,N_27288);
or U29086 (N_29086,N_27005,N_26109);
nand U29087 (N_29087,N_26600,N_27246);
nor U29088 (N_29088,N_27673,N_27367);
nor U29089 (N_29089,N_27983,N_27525);
and U29090 (N_29090,N_27546,N_27816);
xnor U29091 (N_29091,N_26217,N_26447);
or U29092 (N_29092,N_26340,N_26079);
and U29093 (N_29093,N_27997,N_26533);
xnor U29094 (N_29094,N_26566,N_27829);
nor U29095 (N_29095,N_26024,N_27505);
and U29096 (N_29096,N_27694,N_27991);
xnor U29097 (N_29097,N_27886,N_27421);
nand U29098 (N_29098,N_26145,N_26943);
nor U29099 (N_29099,N_27423,N_26674);
and U29100 (N_29100,N_27008,N_27696);
or U29101 (N_29101,N_27355,N_26977);
nor U29102 (N_29102,N_27896,N_26917);
nor U29103 (N_29103,N_27079,N_27608);
or U29104 (N_29104,N_26887,N_26247);
xor U29105 (N_29105,N_26444,N_27724);
and U29106 (N_29106,N_26416,N_26957);
nor U29107 (N_29107,N_27470,N_27447);
nor U29108 (N_29108,N_26991,N_26027);
or U29109 (N_29109,N_27874,N_27325);
and U29110 (N_29110,N_26583,N_26671);
or U29111 (N_29111,N_26605,N_26423);
or U29112 (N_29112,N_27723,N_27474);
nand U29113 (N_29113,N_26536,N_26213);
nand U29114 (N_29114,N_26743,N_26345);
and U29115 (N_29115,N_26332,N_27655);
and U29116 (N_29116,N_26853,N_26141);
nor U29117 (N_29117,N_27521,N_27837);
nor U29118 (N_29118,N_27762,N_27102);
nor U29119 (N_29119,N_27375,N_26486);
xnor U29120 (N_29120,N_27662,N_27007);
nor U29121 (N_29121,N_27201,N_26079);
nor U29122 (N_29122,N_27776,N_27862);
and U29123 (N_29123,N_26367,N_26187);
xnor U29124 (N_29124,N_26629,N_26214);
nor U29125 (N_29125,N_27176,N_27002);
xnor U29126 (N_29126,N_26510,N_27921);
xor U29127 (N_29127,N_26464,N_26923);
nand U29128 (N_29128,N_27653,N_26177);
nor U29129 (N_29129,N_26054,N_26585);
xnor U29130 (N_29130,N_26044,N_27188);
xor U29131 (N_29131,N_27471,N_27133);
and U29132 (N_29132,N_26996,N_26876);
xor U29133 (N_29133,N_27815,N_27786);
nand U29134 (N_29134,N_27082,N_27134);
xnor U29135 (N_29135,N_26022,N_27774);
and U29136 (N_29136,N_26901,N_27492);
or U29137 (N_29137,N_27429,N_27094);
xnor U29138 (N_29138,N_26328,N_26459);
nor U29139 (N_29139,N_26873,N_27434);
or U29140 (N_29140,N_27523,N_27206);
xor U29141 (N_29141,N_27765,N_27948);
nand U29142 (N_29142,N_26253,N_27948);
nor U29143 (N_29143,N_26622,N_27530);
and U29144 (N_29144,N_27479,N_26250);
or U29145 (N_29145,N_26053,N_26723);
or U29146 (N_29146,N_26575,N_27291);
and U29147 (N_29147,N_27178,N_26755);
nor U29148 (N_29148,N_27906,N_27811);
and U29149 (N_29149,N_26072,N_26776);
nor U29150 (N_29150,N_27489,N_26329);
nand U29151 (N_29151,N_27782,N_27283);
and U29152 (N_29152,N_26694,N_26928);
nor U29153 (N_29153,N_26940,N_27246);
xnor U29154 (N_29154,N_27874,N_26997);
and U29155 (N_29155,N_26062,N_27241);
xor U29156 (N_29156,N_26898,N_26338);
nor U29157 (N_29157,N_26700,N_27340);
xor U29158 (N_29158,N_27339,N_26322);
nor U29159 (N_29159,N_27177,N_26683);
nor U29160 (N_29160,N_26138,N_27816);
xnor U29161 (N_29161,N_27276,N_27642);
nand U29162 (N_29162,N_27017,N_26007);
nand U29163 (N_29163,N_26416,N_27290);
nor U29164 (N_29164,N_26133,N_26253);
and U29165 (N_29165,N_27711,N_26434);
nand U29166 (N_29166,N_27430,N_26110);
nand U29167 (N_29167,N_26499,N_26650);
or U29168 (N_29168,N_26672,N_26408);
and U29169 (N_29169,N_27535,N_27373);
nor U29170 (N_29170,N_26052,N_26808);
nor U29171 (N_29171,N_27387,N_27498);
xor U29172 (N_29172,N_27074,N_27786);
xor U29173 (N_29173,N_26013,N_27136);
nand U29174 (N_29174,N_27825,N_27823);
or U29175 (N_29175,N_27816,N_26939);
nand U29176 (N_29176,N_26277,N_26693);
nor U29177 (N_29177,N_26448,N_27118);
and U29178 (N_29178,N_27131,N_26228);
nor U29179 (N_29179,N_26636,N_27127);
and U29180 (N_29180,N_27675,N_26947);
and U29181 (N_29181,N_26453,N_26713);
nor U29182 (N_29182,N_26998,N_26546);
nor U29183 (N_29183,N_27479,N_27694);
nor U29184 (N_29184,N_27478,N_27887);
or U29185 (N_29185,N_27063,N_27907);
nor U29186 (N_29186,N_26788,N_27905);
and U29187 (N_29187,N_26995,N_26779);
nand U29188 (N_29188,N_26865,N_27903);
or U29189 (N_29189,N_26971,N_26119);
xnor U29190 (N_29190,N_26379,N_26598);
xor U29191 (N_29191,N_27894,N_26930);
or U29192 (N_29192,N_26927,N_26364);
nand U29193 (N_29193,N_27036,N_27733);
nand U29194 (N_29194,N_27640,N_26706);
and U29195 (N_29195,N_27276,N_26314);
xnor U29196 (N_29196,N_26412,N_26992);
xor U29197 (N_29197,N_26709,N_26903);
xnor U29198 (N_29198,N_26415,N_27413);
xnor U29199 (N_29199,N_27489,N_26101);
nand U29200 (N_29200,N_27649,N_26871);
or U29201 (N_29201,N_27650,N_27818);
nor U29202 (N_29202,N_26701,N_27018);
or U29203 (N_29203,N_26221,N_26985);
nor U29204 (N_29204,N_27103,N_26857);
xnor U29205 (N_29205,N_26871,N_26666);
nor U29206 (N_29206,N_26729,N_27360);
nand U29207 (N_29207,N_26398,N_27428);
xnor U29208 (N_29208,N_26022,N_27591);
and U29209 (N_29209,N_26337,N_27280);
nor U29210 (N_29210,N_27936,N_26984);
or U29211 (N_29211,N_27875,N_27755);
nor U29212 (N_29212,N_26571,N_26099);
or U29213 (N_29213,N_27209,N_26122);
or U29214 (N_29214,N_27360,N_27996);
nand U29215 (N_29215,N_26502,N_26704);
or U29216 (N_29216,N_26523,N_27662);
or U29217 (N_29217,N_27876,N_26649);
and U29218 (N_29218,N_26086,N_27242);
or U29219 (N_29219,N_26454,N_27165);
nor U29220 (N_29220,N_26674,N_26193);
nor U29221 (N_29221,N_26453,N_27374);
or U29222 (N_29222,N_26913,N_27649);
nor U29223 (N_29223,N_27980,N_27502);
or U29224 (N_29224,N_27200,N_27573);
or U29225 (N_29225,N_27493,N_26749);
or U29226 (N_29226,N_26789,N_26425);
or U29227 (N_29227,N_26681,N_26700);
or U29228 (N_29228,N_27727,N_26716);
nand U29229 (N_29229,N_27068,N_27360);
nor U29230 (N_29230,N_27378,N_26780);
nand U29231 (N_29231,N_27330,N_27765);
and U29232 (N_29232,N_26042,N_27881);
and U29233 (N_29233,N_27638,N_27903);
xor U29234 (N_29234,N_26499,N_26683);
and U29235 (N_29235,N_27003,N_26358);
or U29236 (N_29236,N_27184,N_27543);
xnor U29237 (N_29237,N_27910,N_27536);
or U29238 (N_29238,N_27663,N_26092);
nor U29239 (N_29239,N_27395,N_27503);
nor U29240 (N_29240,N_27015,N_27359);
and U29241 (N_29241,N_27914,N_27130);
nor U29242 (N_29242,N_26588,N_27801);
or U29243 (N_29243,N_26620,N_27685);
xnor U29244 (N_29244,N_27423,N_26010);
nand U29245 (N_29245,N_26925,N_27981);
or U29246 (N_29246,N_26021,N_26832);
nor U29247 (N_29247,N_26954,N_26829);
nor U29248 (N_29248,N_26805,N_27250);
or U29249 (N_29249,N_27579,N_26581);
and U29250 (N_29250,N_27472,N_26553);
nand U29251 (N_29251,N_26372,N_26515);
xnor U29252 (N_29252,N_27686,N_27125);
nor U29253 (N_29253,N_26838,N_26363);
nor U29254 (N_29254,N_27570,N_27432);
xnor U29255 (N_29255,N_26733,N_27034);
xor U29256 (N_29256,N_27369,N_26437);
nand U29257 (N_29257,N_27510,N_26344);
nor U29258 (N_29258,N_27917,N_27276);
xnor U29259 (N_29259,N_26758,N_27548);
and U29260 (N_29260,N_27173,N_27698);
xnor U29261 (N_29261,N_27046,N_27073);
nand U29262 (N_29262,N_27443,N_27900);
xor U29263 (N_29263,N_26081,N_26409);
xor U29264 (N_29264,N_27088,N_27116);
or U29265 (N_29265,N_26264,N_26920);
and U29266 (N_29266,N_26387,N_26870);
nand U29267 (N_29267,N_27305,N_27013);
and U29268 (N_29268,N_26073,N_27903);
and U29269 (N_29269,N_27231,N_26358);
nand U29270 (N_29270,N_27768,N_27879);
and U29271 (N_29271,N_27049,N_27345);
nand U29272 (N_29272,N_26506,N_27607);
nand U29273 (N_29273,N_27098,N_26336);
xor U29274 (N_29274,N_27382,N_27825);
nor U29275 (N_29275,N_26449,N_26101);
nor U29276 (N_29276,N_27846,N_26943);
nand U29277 (N_29277,N_27229,N_27264);
nand U29278 (N_29278,N_27617,N_27149);
nor U29279 (N_29279,N_26113,N_27344);
xnor U29280 (N_29280,N_26295,N_27454);
nand U29281 (N_29281,N_27594,N_26407);
xnor U29282 (N_29282,N_27599,N_26624);
xnor U29283 (N_29283,N_26260,N_27476);
xnor U29284 (N_29284,N_26198,N_27921);
xor U29285 (N_29285,N_27914,N_26957);
or U29286 (N_29286,N_26441,N_27548);
xnor U29287 (N_29287,N_26497,N_26877);
nor U29288 (N_29288,N_27761,N_27594);
and U29289 (N_29289,N_27470,N_27595);
or U29290 (N_29290,N_26709,N_27352);
and U29291 (N_29291,N_27921,N_27131);
nand U29292 (N_29292,N_27970,N_26351);
and U29293 (N_29293,N_27251,N_26125);
nand U29294 (N_29294,N_26521,N_27498);
nand U29295 (N_29295,N_27208,N_26615);
nand U29296 (N_29296,N_27538,N_27055);
nor U29297 (N_29297,N_26469,N_27395);
and U29298 (N_29298,N_26000,N_26694);
or U29299 (N_29299,N_27576,N_27203);
or U29300 (N_29300,N_26833,N_26430);
xnor U29301 (N_29301,N_26719,N_26266);
nor U29302 (N_29302,N_26869,N_26244);
nor U29303 (N_29303,N_26923,N_27760);
nor U29304 (N_29304,N_27551,N_26234);
xnor U29305 (N_29305,N_27494,N_27937);
nand U29306 (N_29306,N_27364,N_26477);
and U29307 (N_29307,N_27599,N_27637);
nor U29308 (N_29308,N_27945,N_27632);
or U29309 (N_29309,N_26484,N_27537);
or U29310 (N_29310,N_27642,N_27943);
nor U29311 (N_29311,N_26403,N_27085);
xnor U29312 (N_29312,N_27975,N_26302);
nand U29313 (N_29313,N_27697,N_27549);
or U29314 (N_29314,N_26367,N_27006);
nand U29315 (N_29315,N_27728,N_27670);
nand U29316 (N_29316,N_26605,N_26909);
xnor U29317 (N_29317,N_26145,N_26887);
or U29318 (N_29318,N_26079,N_26958);
nor U29319 (N_29319,N_27065,N_26737);
nand U29320 (N_29320,N_27351,N_27040);
or U29321 (N_29321,N_26332,N_27808);
xor U29322 (N_29322,N_26975,N_26385);
and U29323 (N_29323,N_27538,N_27822);
nand U29324 (N_29324,N_26289,N_27849);
nor U29325 (N_29325,N_27916,N_27510);
or U29326 (N_29326,N_27943,N_27103);
or U29327 (N_29327,N_26160,N_27476);
or U29328 (N_29328,N_26187,N_27156);
xnor U29329 (N_29329,N_26733,N_27410);
xor U29330 (N_29330,N_26669,N_26782);
nand U29331 (N_29331,N_26130,N_27924);
nor U29332 (N_29332,N_26632,N_27825);
and U29333 (N_29333,N_27922,N_27434);
nor U29334 (N_29334,N_26451,N_27538);
or U29335 (N_29335,N_26689,N_27587);
and U29336 (N_29336,N_26947,N_26680);
nor U29337 (N_29337,N_26420,N_27596);
nand U29338 (N_29338,N_26383,N_26416);
xor U29339 (N_29339,N_26047,N_26388);
nand U29340 (N_29340,N_27771,N_26010);
nor U29341 (N_29341,N_27815,N_26396);
nor U29342 (N_29342,N_27163,N_26670);
nor U29343 (N_29343,N_26812,N_26931);
xor U29344 (N_29344,N_27260,N_27586);
and U29345 (N_29345,N_26186,N_27492);
nor U29346 (N_29346,N_26874,N_26530);
or U29347 (N_29347,N_27588,N_27239);
xor U29348 (N_29348,N_26110,N_26735);
nand U29349 (N_29349,N_27951,N_26187);
and U29350 (N_29350,N_27557,N_26821);
nand U29351 (N_29351,N_26417,N_27745);
and U29352 (N_29352,N_26571,N_27979);
xor U29353 (N_29353,N_26230,N_26479);
and U29354 (N_29354,N_26152,N_27409);
and U29355 (N_29355,N_26122,N_26762);
xor U29356 (N_29356,N_27321,N_26700);
and U29357 (N_29357,N_27378,N_26593);
xnor U29358 (N_29358,N_26965,N_27331);
nand U29359 (N_29359,N_27047,N_27380);
nand U29360 (N_29360,N_27753,N_27199);
and U29361 (N_29361,N_27144,N_27733);
and U29362 (N_29362,N_27355,N_27749);
nand U29363 (N_29363,N_27265,N_27881);
or U29364 (N_29364,N_27529,N_26832);
and U29365 (N_29365,N_26013,N_27310);
or U29366 (N_29366,N_26198,N_27347);
nand U29367 (N_29367,N_27550,N_26318);
nand U29368 (N_29368,N_27908,N_27872);
or U29369 (N_29369,N_26018,N_26587);
xnor U29370 (N_29370,N_27101,N_27359);
xnor U29371 (N_29371,N_26770,N_27533);
and U29372 (N_29372,N_27474,N_26295);
and U29373 (N_29373,N_27368,N_27933);
and U29374 (N_29374,N_27493,N_26002);
and U29375 (N_29375,N_27791,N_26899);
nor U29376 (N_29376,N_26944,N_26543);
xnor U29377 (N_29377,N_26928,N_27647);
nor U29378 (N_29378,N_27213,N_26275);
nand U29379 (N_29379,N_27584,N_27220);
nor U29380 (N_29380,N_27693,N_27798);
nand U29381 (N_29381,N_27387,N_27715);
or U29382 (N_29382,N_27355,N_27463);
and U29383 (N_29383,N_27602,N_26409);
nor U29384 (N_29384,N_27807,N_26085);
xnor U29385 (N_29385,N_27076,N_27900);
nor U29386 (N_29386,N_27963,N_26207);
nor U29387 (N_29387,N_27567,N_26078);
xor U29388 (N_29388,N_26396,N_27232);
and U29389 (N_29389,N_26781,N_26934);
xor U29390 (N_29390,N_26105,N_26123);
xor U29391 (N_29391,N_26171,N_27224);
nand U29392 (N_29392,N_27758,N_27123);
nand U29393 (N_29393,N_26712,N_26982);
and U29394 (N_29394,N_27490,N_27394);
and U29395 (N_29395,N_26521,N_26147);
nand U29396 (N_29396,N_26331,N_27847);
or U29397 (N_29397,N_26934,N_26301);
and U29398 (N_29398,N_26554,N_26857);
nor U29399 (N_29399,N_27445,N_27474);
and U29400 (N_29400,N_27301,N_27057);
xnor U29401 (N_29401,N_27002,N_27313);
and U29402 (N_29402,N_26414,N_27770);
xor U29403 (N_29403,N_27781,N_26979);
nor U29404 (N_29404,N_27106,N_27263);
xor U29405 (N_29405,N_26221,N_27971);
or U29406 (N_29406,N_26155,N_27045);
xor U29407 (N_29407,N_26213,N_27607);
and U29408 (N_29408,N_26396,N_27416);
nand U29409 (N_29409,N_26351,N_26940);
nor U29410 (N_29410,N_27520,N_27923);
nand U29411 (N_29411,N_26877,N_26123);
nor U29412 (N_29412,N_27656,N_26391);
or U29413 (N_29413,N_27907,N_26563);
xor U29414 (N_29414,N_27354,N_26842);
and U29415 (N_29415,N_26053,N_26311);
and U29416 (N_29416,N_27231,N_27985);
or U29417 (N_29417,N_27123,N_26079);
xor U29418 (N_29418,N_26547,N_27719);
or U29419 (N_29419,N_27078,N_26705);
or U29420 (N_29420,N_26098,N_26748);
or U29421 (N_29421,N_26883,N_26197);
and U29422 (N_29422,N_27530,N_26886);
nand U29423 (N_29423,N_27714,N_27967);
or U29424 (N_29424,N_27723,N_27162);
nor U29425 (N_29425,N_26727,N_26117);
or U29426 (N_29426,N_26098,N_27562);
xor U29427 (N_29427,N_26443,N_26318);
xor U29428 (N_29428,N_27345,N_26864);
nand U29429 (N_29429,N_27015,N_27805);
xnor U29430 (N_29430,N_26204,N_27841);
or U29431 (N_29431,N_27061,N_27894);
xor U29432 (N_29432,N_26129,N_26537);
nor U29433 (N_29433,N_27678,N_26536);
and U29434 (N_29434,N_26080,N_26402);
nor U29435 (N_29435,N_26409,N_27727);
nor U29436 (N_29436,N_27977,N_26479);
nor U29437 (N_29437,N_27528,N_27980);
nor U29438 (N_29438,N_26272,N_26166);
nor U29439 (N_29439,N_26078,N_26173);
nor U29440 (N_29440,N_27732,N_27885);
xnor U29441 (N_29441,N_26050,N_26666);
and U29442 (N_29442,N_27123,N_26981);
or U29443 (N_29443,N_26664,N_26545);
and U29444 (N_29444,N_26490,N_26097);
nor U29445 (N_29445,N_26171,N_26300);
xnor U29446 (N_29446,N_27715,N_26602);
or U29447 (N_29447,N_27775,N_27622);
xnor U29448 (N_29448,N_27656,N_26703);
nand U29449 (N_29449,N_27172,N_26196);
and U29450 (N_29450,N_27550,N_26940);
nand U29451 (N_29451,N_26535,N_27800);
and U29452 (N_29452,N_26314,N_27797);
and U29453 (N_29453,N_26367,N_27025);
xnor U29454 (N_29454,N_27465,N_27524);
or U29455 (N_29455,N_26552,N_27022);
and U29456 (N_29456,N_27697,N_26072);
and U29457 (N_29457,N_27049,N_26817);
nor U29458 (N_29458,N_26327,N_26342);
or U29459 (N_29459,N_26576,N_26151);
or U29460 (N_29460,N_27755,N_27599);
and U29461 (N_29461,N_26495,N_26190);
or U29462 (N_29462,N_27455,N_27182);
xor U29463 (N_29463,N_26481,N_26801);
nor U29464 (N_29464,N_26560,N_26714);
nand U29465 (N_29465,N_27042,N_26689);
or U29466 (N_29466,N_27401,N_27189);
xor U29467 (N_29467,N_26613,N_26217);
or U29468 (N_29468,N_27432,N_26909);
nand U29469 (N_29469,N_26920,N_26703);
nand U29470 (N_29470,N_27709,N_27484);
and U29471 (N_29471,N_27405,N_26274);
or U29472 (N_29472,N_27609,N_26346);
nor U29473 (N_29473,N_26795,N_27306);
nor U29474 (N_29474,N_27889,N_26869);
and U29475 (N_29475,N_27617,N_27937);
xor U29476 (N_29476,N_27693,N_27001);
nor U29477 (N_29477,N_27181,N_26952);
xnor U29478 (N_29478,N_26696,N_27280);
or U29479 (N_29479,N_27645,N_27125);
nand U29480 (N_29480,N_26580,N_27027);
or U29481 (N_29481,N_27011,N_26008);
nand U29482 (N_29482,N_27415,N_26007);
and U29483 (N_29483,N_26735,N_26249);
nor U29484 (N_29484,N_27644,N_26096);
and U29485 (N_29485,N_27902,N_27463);
nor U29486 (N_29486,N_27544,N_27529);
nand U29487 (N_29487,N_27441,N_27093);
xor U29488 (N_29488,N_27864,N_26516);
or U29489 (N_29489,N_26624,N_27087);
and U29490 (N_29490,N_27106,N_27381);
and U29491 (N_29491,N_27964,N_26570);
nor U29492 (N_29492,N_26634,N_26941);
or U29493 (N_29493,N_27723,N_27556);
nor U29494 (N_29494,N_26969,N_26004);
and U29495 (N_29495,N_27455,N_26250);
nor U29496 (N_29496,N_26624,N_27125);
nor U29497 (N_29497,N_27679,N_27991);
xor U29498 (N_29498,N_27047,N_27782);
xor U29499 (N_29499,N_26600,N_26104);
and U29500 (N_29500,N_26005,N_26544);
nand U29501 (N_29501,N_27326,N_26319);
and U29502 (N_29502,N_27122,N_27743);
nor U29503 (N_29503,N_26668,N_27809);
nor U29504 (N_29504,N_26927,N_26745);
nor U29505 (N_29505,N_26186,N_27670);
or U29506 (N_29506,N_26966,N_27252);
xor U29507 (N_29507,N_27493,N_27837);
and U29508 (N_29508,N_26375,N_26978);
xor U29509 (N_29509,N_27753,N_26457);
nor U29510 (N_29510,N_26907,N_26150);
xnor U29511 (N_29511,N_26304,N_26371);
xor U29512 (N_29512,N_27731,N_27188);
and U29513 (N_29513,N_27168,N_27876);
nand U29514 (N_29514,N_26526,N_26996);
and U29515 (N_29515,N_27516,N_26407);
and U29516 (N_29516,N_27233,N_26306);
nor U29517 (N_29517,N_27625,N_26690);
xnor U29518 (N_29518,N_27984,N_27521);
xnor U29519 (N_29519,N_26076,N_26797);
or U29520 (N_29520,N_26411,N_27506);
nor U29521 (N_29521,N_27321,N_26369);
and U29522 (N_29522,N_27880,N_26070);
nor U29523 (N_29523,N_27743,N_26503);
or U29524 (N_29524,N_27933,N_26427);
nor U29525 (N_29525,N_27486,N_27285);
nand U29526 (N_29526,N_27049,N_26783);
nor U29527 (N_29527,N_26804,N_27649);
xor U29528 (N_29528,N_27038,N_27205);
and U29529 (N_29529,N_26620,N_26158);
and U29530 (N_29530,N_27076,N_26588);
nand U29531 (N_29531,N_26266,N_26363);
and U29532 (N_29532,N_26658,N_27674);
and U29533 (N_29533,N_26516,N_26256);
or U29534 (N_29534,N_26253,N_27478);
and U29535 (N_29535,N_27312,N_27616);
and U29536 (N_29536,N_27372,N_27681);
or U29537 (N_29537,N_26881,N_26762);
xor U29538 (N_29538,N_27969,N_27523);
xnor U29539 (N_29539,N_27420,N_27224);
nand U29540 (N_29540,N_27032,N_26147);
nand U29541 (N_29541,N_27038,N_26046);
or U29542 (N_29542,N_26790,N_27628);
xor U29543 (N_29543,N_27724,N_27232);
nand U29544 (N_29544,N_26579,N_26297);
or U29545 (N_29545,N_27832,N_27454);
xnor U29546 (N_29546,N_27303,N_27944);
or U29547 (N_29547,N_26643,N_27172);
nand U29548 (N_29548,N_26994,N_26086);
nor U29549 (N_29549,N_27539,N_26811);
xor U29550 (N_29550,N_26557,N_26382);
nand U29551 (N_29551,N_27187,N_26890);
xor U29552 (N_29552,N_26775,N_27127);
nor U29553 (N_29553,N_26123,N_27139);
and U29554 (N_29554,N_26658,N_27535);
xor U29555 (N_29555,N_26988,N_26023);
xnor U29556 (N_29556,N_26413,N_26156);
nor U29557 (N_29557,N_26891,N_27227);
or U29558 (N_29558,N_27871,N_26346);
xor U29559 (N_29559,N_26408,N_26336);
and U29560 (N_29560,N_27844,N_26528);
or U29561 (N_29561,N_27437,N_27501);
nor U29562 (N_29562,N_27689,N_27763);
xnor U29563 (N_29563,N_26171,N_26773);
nand U29564 (N_29564,N_27172,N_26368);
nand U29565 (N_29565,N_27703,N_27790);
and U29566 (N_29566,N_27045,N_27764);
xnor U29567 (N_29567,N_26627,N_27569);
xnor U29568 (N_29568,N_27790,N_26135);
or U29569 (N_29569,N_26260,N_26489);
nor U29570 (N_29570,N_26006,N_26198);
and U29571 (N_29571,N_27503,N_26283);
or U29572 (N_29572,N_26870,N_27107);
nand U29573 (N_29573,N_27796,N_27143);
nand U29574 (N_29574,N_26507,N_27882);
nand U29575 (N_29575,N_26278,N_27314);
and U29576 (N_29576,N_27336,N_26791);
nor U29577 (N_29577,N_26920,N_27622);
nor U29578 (N_29578,N_27584,N_27003);
nor U29579 (N_29579,N_26475,N_26765);
xnor U29580 (N_29580,N_26501,N_27269);
nand U29581 (N_29581,N_26007,N_27366);
xor U29582 (N_29582,N_26049,N_27516);
or U29583 (N_29583,N_26846,N_26300);
xnor U29584 (N_29584,N_27380,N_26664);
nor U29585 (N_29585,N_27539,N_27247);
and U29586 (N_29586,N_26486,N_27855);
and U29587 (N_29587,N_27084,N_27334);
nand U29588 (N_29588,N_27673,N_26721);
xnor U29589 (N_29589,N_27106,N_27594);
xnor U29590 (N_29590,N_27108,N_26282);
nand U29591 (N_29591,N_27330,N_27250);
and U29592 (N_29592,N_27432,N_27756);
nand U29593 (N_29593,N_27695,N_27580);
and U29594 (N_29594,N_26900,N_26522);
and U29595 (N_29595,N_26796,N_27169);
nand U29596 (N_29596,N_26255,N_26591);
xnor U29597 (N_29597,N_26374,N_26250);
or U29598 (N_29598,N_26011,N_27214);
nand U29599 (N_29599,N_26543,N_26211);
and U29600 (N_29600,N_27404,N_27592);
nand U29601 (N_29601,N_27147,N_27793);
or U29602 (N_29602,N_27458,N_26855);
nor U29603 (N_29603,N_27823,N_27469);
xor U29604 (N_29604,N_27064,N_26092);
and U29605 (N_29605,N_26426,N_26211);
or U29606 (N_29606,N_26382,N_26832);
nand U29607 (N_29607,N_26887,N_26640);
or U29608 (N_29608,N_26769,N_26026);
nor U29609 (N_29609,N_26486,N_27826);
xor U29610 (N_29610,N_26296,N_26341);
nor U29611 (N_29611,N_26592,N_27376);
and U29612 (N_29612,N_27172,N_27323);
or U29613 (N_29613,N_27926,N_26941);
xor U29614 (N_29614,N_26160,N_27532);
or U29615 (N_29615,N_26557,N_27355);
nor U29616 (N_29616,N_26491,N_26818);
and U29617 (N_29617,N_27749,N_27494);
or U29618 (N_29618,N_27451,N_26407);
nand U29619 (N_29619,N_27592,N_27445);
nand U29620 (N_29620,N_26644,N_27712);
or U29621 (N_29621,N_26476,N_26512);
nand U29622 (N_29622,N_27753,N_27774);
xnor U29623 (N_29623,N_26976,N_27747);
xnor U29624 (N_29624,N_27090,N_27625);
nor U29625 (N_29625,N_26789,N_26723);
nand U29626 (N_29626,N_26921,N_27084);
nor U29627 (N_29627,N_27711,N_26751);
nor U29628 (N_29628,N_27536,N_26912);
or U29629 (N_29629,N_27496,N_27360);
nor U29630 (N_29630,N_26795,N_27879);
and U29631 (N_29631,N_26930,N_26486);
nand U29632 (N_29632,N_26727,N_26968);
nor U29633 (N_29633,N_26050,N_26392);
and U29634 (N_29634,N_27935,N_27822);
and U29635 (N_29635,N_27616,N_26896);
xnor U29636 (N_29636,N_27000,N_26256);
nand U29637 (N_29637,N_26665,N_27565);
xor U29638 (N_29638,N_26546,N_26196);
and U29639 (N_29639,N_27945,N_26006);
xnor U29640 (N_29640,N_26305,N_27789);
and U29641 (N_29641,N_27863,N_27668);
nand U29642 (N_29642,N_26197,N_27807);
xor U29643 (N_29643,N_26250,N_27554);
or U29644 (N_29644,N_27089,N_27979);
and U29645 (N_29645,N_27346,N_26731);
nand U29646 (N_29646,N_27897,N_27179);
xor U29647 (N_29647,N_26306,N_27840);
or U29648 (N_29648,N_27985,N_26672);
nor U29649 (N_29649,N_27384,N_27100);
or U29650 (N_29650,N_26341,N_26798);
and U29651 (N_29651,N_27287,N_27019);
xor U29652 (N_29652,N_27273,N_26112);
and U29653 (N_29653,N_26929,N_27944);
and U29654 (N_29654,N_27259,N_27025);
nand U29655 (N_29655,N_27101,N_26082);
xor U29656 (N_29656,N_26624,N_27716);
or U29657 (N_29657,N_26161,N_27315);
and U29658 (N_29658,N_27298,N_26973);
nand U29659 (N_29659,N_26623,N_26378);
nor U29660 (N_29660,N_26516,N_26875);
and U29661 (N_29661,N_26792,N_27006);
nand U29662 (N_29662,N_26547,N_27364);
and U29663 (N_29663,N_27416,N_26226);
and U29664 (N_29664,N_26498,N_27247);
xnor U29665 (N_29665,N_27483,N_27249);
and U29666 (N_29666,N_26950,N_26055);
nor U29667 (N_29667,N_26315,N_27586);
or U29668 (N_29668,N_26521,N_26096);
nor U29669 (N_29669,N_26748,N_27914);
and U29670 (N_29670,N_26848,N_27901);
nand U29671 (N_29671,N_27930,N_27588);
xnor U29672 (N_29672,N_26587,N_27117);
nor U29673 (N_29673,N_27289,N_26542);
nand U29674 (N_29674,N_27323,N_26117);
nor U29675 (N_29675,N_26664,N_26547);
nor U29676 (N_29676,N_27651,N_27910);
nor U29677 (N_29677,N_27611,N_26160);
nand U29678 (N_29678,N_26637,N_27631);
nor U29679 (N_29679,N_26319,N_27702);
xor U29680 (N_29680,N_26045,N_26787);
or U29681 (N_29681,N_26370,N_26056);
nand U29682 (N_29682,N_26438,N_26508);
xnor U29683 (N_29683,N_26634,N_27977);
xnor U29684 (N_29684,N_26671,N_26951);
and U29685 (N_29685,N_27266,N_26344);
xnor U29686 (N_29686,N_27572,N_27605);
nor U29687 (N_29687,N_26722,N_27136);
nor U29688 (N_29688,N_27933,N_27091);
xnor U29689 (N_29689,N_26236,N_26956);
and U29690 (N_29690,N_26873,N_27574);
or U29691 (N_29691,N_26686,N_26326);
and U29692 (N_29692,N_27989,N_27410);
nand U29693 (N_29693,N_26279,N_26055);
and U29694 (N_29694,N_27305,N_26652);
and U29695 (N_29695,N_26221,N_26053);
nand U29696 (N_29696,N_26577,N_26695);
nor U29697 (N_29697,N_26341,N_26162);
nor U29698 (N_29698,N_27888,N_27381);
or U29699 (N_29699,N_27072,N_26157);
nand U29700 (N_29700,N_27312,N_27787);
nor U29701 (N_29701,N_27992,N_26647);
or U29702 (N_29702,N_26360,N_26835);
or U29703 (N_29703,N_27328,N_26600);
or U29704 (N_29704,N_27209,N_26617);
nor U29705 (N_29705,N_26492,N_27912);
nor U29706 (N_29706,N_27804,N_27558);
xor U29707 (N_29707,N_26017,N_26511);
or U29708 (N_29708,N_26279,N_27371);
nor U29709 (N_29709,N_27591,N_26924);
nand U29710 (N_29710,N_26604,N_26037);
nor U29711 (N_29711,N_27924,N_26988);
or U29712 (N_29712,N_26085,N_26713);
xor U29713 (N_29713,N_27431,N_27467);
xnor U29714 (N_29714,N_27762,N_27311);
nor U29715 (N_29715,N_27400,N_27870);
nor U29716 (N_29716,N_27200,N_26569);
nand U29717 (N_29717,N_26949,N_27588);
nand U29718 (N_29718,N_26250,N_27337);
or U29719 (N_29719,N_26028,N_27144);
xor U29720 (N_29720,N_27928,N_26929);
and U29721 (N_29721,N_26518,N_27257);
nor U29722 (N_29722,N_27437,N_27557);
nand U29723 (N_29723,N_27318,N_27524);
nor U29724 (N_29724,N_26743,N_26848);
nand U29725 (N_29725,N_26238,N_26994);
nor U29726 (N_29726,N_27676,N_26096);
nand U29727 (N_29727,N_26126,N_26238);
nand U29728 (N_29728,N_27233,N_26289);
or U29729 (N_29729,N_27008,N_26523);
xnor U29730 (N_29730,N_27658,N_27394);
nand U29731 (N_29731,N_27774,N_27064);
or U29732 (N_29732,N_26308,N_27689);
or U29733 (N_29733,N_27854,N_27440);
xor U29734 (N_29734,N_26785,N_26863);
nor U29735 (N_29735,N_27250,N_27856);
or U29736 (N_29736,N_27876,N_26095);
nand U29737 (N_29737,N_27557,N_27533);
or U29738 (N_29738,N_26017,N_27707);
xor U29739 (N_29739,N_27809,N_26861);
nor U29740 (N_29740,N_26560,N_26071);
nor U29741 (N_29741,N_27333,N_27551);
and U29742 (N_29742,N_26942,N_27463);
xnor U29743 (N_29743,N_26942,N_26130);
and U29744 (N_29744,N_26706,N_26310);
nand U29745 (N_29745,N_27079,N_26890);
nor U29746 (N_29746,N_27769,N_26074);
and U29747 (N_29747,N_26975,N_26431);
nand U29748 (N_29748,N_27774,N_26546);
xor U29749 (N_29749,N_27009,N_26373);
nor U29750 (N_29750,N_26255,N_27494);
nand U29751 (N_29751,N_26866,N_26883);
xnor U29752 (N_29752,N_26298,N_27142);
xor U29753 (N_29753,N_26449,N_27945);
or U29754 (N_29754,N_26156,N_26483);
nand U29755 (N_29755,N_27428,N_26932);
nand U29756 (N_29756,N_27492,N_27741);
and U29757 (N_29757,N_26546,N_26784);
or U29758 (N_29758,N_27472,N_26710);
or U29759 (N_29759,N_26489,N_27230);
nor U29760 (N_29760,N_26382,N_27296);
and U29761 (N_29761,N_27302,N_27780);
or U29762 (N_29762,N_27860,N_26783);
and U29763 (N_29763,N_26960,N_26841);
or U29764 (N_29764,N_26789,N_27552);
nor U29765 (N_29765,N_26288,N_27157);
xnor U29766 (N_29766,N_26330,N_27209);
xnor U29767 (N_29767,N_27241,N_26687);
nand U29768 (N_29768,N_27568,N_26682);
and U29769 (N_29769,N_26295,N_27821);
nor U29770 (N_29770,N_27408,N_26142);
nand U29771 (N_29771,N_27929,N_27891);
and U29772 (N_29772,N_27620,N_26509);
nand U29773 (N_29773,N_27967,N_27375);
and U29774 (N_29774,N_26549,N_27122);
and U29775 (N_29775,N_27203,N_26005);
or U29776 (N_29776,N_26566,N_27287);
xor U29777 (N_29777,N_27248,N_26259);
nand U29778 (N_29778,N_27021,N_26975);
nand U29779 (N_29779,N_26806,N_26705);
and U29780 (N_29780,N_27218,N_26581);
xnor U29781 (N_29781,N_27530,N_26288);
nor U29782 (N_29782,N_27943,N_26647);
nand U29783 (N_29783,N_27192,N_27277);
xor U29784 (N_29784,N_26754,N_26753);
nand U29785 (N_29785,N_27771,N_26326);
and U29786 (N_29786,N_26433,N_26820);
nor U29787 (N_29787,N_26353,N_27289);
nor U29788 (N_29788,N_26367,N_26756);
nand U29789 (N_29789,N_26754,N_26282);
or U29790 (N_29790,N_27523,N_26848);
and U29791 (N_29791,N_27640,N_26360);
nor U29792 (N_29792,N_27611,N_27652);
and U29793 (N_29793,N_26094,N_26058);
xor U29794 (N_29794,N_27006,N_27548);
and U29795 (N_29795,N_27125,N_26067);
nand U29796 (N_29796,N_26285,N_27626);
nand U29797 (N_29797,N_27518,N_27983);
and U29798 (N_29798,N_27358,N_26894);
or U29799 (N_29799,N_26253,N_27416);
nor U29800 (N_29800,N_27446,N_27300);
nand U29801 (N_29801,N_26177,N_27816);
nand U29802 (N_29802,N_26294,N_27934);
or U29803 (N_29803,N_27076,N_27193);
and U29804 (N_29804,N_27457,N_27868);
xor U29805 (N_29805,N_27441,N_27116);
nand U29806 (N_29806,N_27014,N_27071);
and U29807 (N_29807,N_27786,N_26095);
nor U29808 (N_29808,N_26797,N_27192);
nor U29809 (N_29809,N_26726,N_27659);
nand U29810 (N_29810,N_27851,N_26481);
or U29811 (N_29811,N_26204,N_27024);
nand U29812 (N_29812,N_27196,N_26429);
xnor U29813 (N_29813,N_27763,N_27201);
nand U29814 (N_29814,N_27419,N_27122);
or U29815 (N_29815,N_26949,N_26451);
or U29816 (N_29816,N_26232,N_27376);
xor U29817 (N_29817,N_26601,N_27188);
xnor U29818 (N_29818,N_26797,N_26973);
xor U29819 (N_29819,N_27937,N_26023);
or U29820 (N_29820,N_26113,N_27644);
xnor U29821 (N_29821,N_26568,N_26340);
nor U29822 (N_29822,N_26768,N_27845);
or U29823 (N_29823,N_26133,N_26168);
and U29824 (N_29824,N_27045,N_26657);
xnor U29825 (N_29825,N_26281,N_27735);
xor U29826 (N_29826,N_26185,N_26063);
or U29827 (N_29827,N_27245,N_26539);
nand U29828 (N_29828,N_26146,N_27488);
nor U29829 (N_29829,N_26827,N_27110);
nand U29830 (N_29830,N_27627,N_27327);
xnor U29831 (N_29831,N_26660,N_27407);
nor U29832 (N_29832,N_26331,N_27097);
nand U29833 (N_29833,N_26861,N_27965);
or U29834 (N_29834,N_27868,N_27293);
and U29835 (N_29835,N_26352,N_26906);
or U29836 (N_29836,N_27981,N_27156);
nor U29837 (N_29837,N_26211,N_26466);
or U29838 (N_29838,N_27204,N_27671);
or U29839 (N_29839,N_26007,N_27889);
xnor U29840 (N_29840,N_26556,N_26505);
and U29841 (N_29841,N_26480,N_27492);
nand U29842 (N_29842,N_26488,N_27274);
xnor U29843 (N_29843,N_26857,N_27480);
and U29844 (N_29844,N_26470,N_26574);
and U29845 (N_29845,N_26610,N_27777);
or U29846 (N_29846,N_26216,N_27034);
xnor U29847 (N_29847,N_26402,N_26057);
and U29848 (N_29848,N_26567,N_27627);
nand U29849 (N_29849,N_26273,N_27439);
nor U29850 (N_29850,N_26539,N_27603);
or U29851 (N_29851,N_26802,N_26968);
nand U29852 (N_29852,N_27434,N_26369);
xnor U29853 (N_29853,N_27867,N_27380);
or U29854 (N_29854,N_27592,N_26103);
and U29855 (N_29855,N_26406,N_27399);
and U29856 (N_29856,N_26197,N_26843);
and U29857 (N_29857,N_27772,N_27959);
xnor U29858 (N_29858,N_27066,N_27631);
nand U29859 (N_29859,N_27174,N_26409);
or U29860 (N_29860,N_27357,N_27921);
xor U29861 (N_29861,N_27794,N_26191);
nor U29862 (N_29862,N_27892,N_26888);
nand U29863 (N_29863,N_26603,N_27399);
nand U29864 (N_29864,N_27383,N_26017);
nor U29865 (N_29865,N_26477,N_27506);
nand U29866 (N_29866,N_27641,N_27394);
or U29867 (N_29867,N_26980,N_26920);
nor U29868 (N_29868,N_26472,N_27959);
or U29869 (N_29869,N_26573,N_26909);
xor U29870 (N_29870,N_27788,N_27563);
xor U29871 (N_29871,N_27320,N_26529);
xor U29872 (N_29872,N_26542,N_27381);
nand U29873 (N_29873,N_26246,N_26017);
and U29874 (N_29874,N_27641,N_26597);
nor U29875 (N_29875,N_27799,N_26333);
or U29876 (N_29876,N_26531,N_26056);
or U29877 (N_29877,N_26592,N_27028);
or U29878 (N_29878,N_26593,N_26878);
and U29879 (N_29879,N_27759,N_27706);
or U29880 (N_29880,N_27259,N_27563);
and U29881 (N_29881,N_26586,N_26013);
and U29882 (N_29882,N_26473,N_27764);
nand U29883 (N_29883,N_27868,N_26796);
or U29884 (N_29884,N_27684,N_27781);
or U29885 (N_29885,N_27932,N_27624);
nor U29886 (N_29886,N_26174,N_26441);
nand U29887 (N_29887,N_26595,N_27416);
and U29888 (N_29888,N_27020,N_26860);
or U29889 (N_29889,N_26796,N_26028);
xor U29890 (N_29890,N_27751,N_27803);
and U29891 (N_29891,N_27286,N_26809);
nor U29892 (N_29892,N_26613,N_27722);
nand U29893 (N_29893,N_27281,N_26009);
nand U29894 (N_29894,N_27411,N_27218);
or U29895 (N_29895,N_27846,N_26383);
nor U29896 (N_29896,N_27564,N_26992);
nor U29897 (N_29897,N_27696,N_26964);
and U29898 (N_29898,N_26009,N_27991);
or U29899 (N_29899,N_26808,N_26295);
nor U29900 (N_29900,N_26349,N_26807);
nor U29901 (N_29901,N_26304,N_26819);
nor U29902 (N_29902,N_27586,N_26243);
and U29903 (N_29903,N_27067,N_26775);
xnor U29904 (N_29904,N_27274,N_27635);
nand U29905 (N_29905,N_26740,N_27572);
and U29906 (N_29906,N_27346,N_26313);
nand U29907 (N_29907,N_27936,N_26544);
and U29908 (N_29908,N_27290,N_27139);
nand U29909 (N_29909,N_27898,N_27831);
xnor U29910 (N_29910,N_26066,N_27360);
nor U29911 (N_29911,N_27969,N_27890);
nand U29912 (N_29912,N_26896,N_27099);
nor U29913 (N_29913,N_26032,N_27286);
xnor U29914 (N_29914,N_27360,N_27052);
nor U29915 (N_29915,N_27056,N_27996);
or U29916 (N_29916,N_26713,N_27334);
and U29917 (N_29917,N_26971,N_27252);
xor U29918 (N_29918,N_26649,N_26424);
nand U29919 (N_29919,N_27734,N_27925);
nor U29920 (N_29920,N_27012,N_26442);
nand U29921 (N_29921,N_27962,N_27376);
nand U29922 (N_29922,N_26040,N_26617);
or U29923 (N_29923,N_26054,N_26090);
and U29924 (N_29924,N_27886,N_27936);
xnor U29925 (N_29925,N_26439,N_26072);
or U29926 (N_29926,N_27121,N_26065);
and U29927 (N_29927,N_26198,N_27947);
and U29928 (N_29928,N_26041,N_26332);
and U29929 (N_29929,N_27332,N_26512);
nor U29930 (N_29930,N_27589,N_26645);
xnor U29931 (N_29931,N_26358,N_27841);
and U29932 (N_29932,N_27181,N_26922);
xnor U29933 (N_29933,N_27251,N_26055);
nor U29934 (N_29934,N_26337,N_26790);
or U29935 (N_29935,N_27130,N_26333);
nand U29936 (N_29936,N_26768,N_26714);
or U29937 (N_29937,N_26010,N_27361);
and U29938 (N_29938,N_27579,N_27095);
and U29939 (N_29939,N_26046,N_26912);
and U29940 (N_29940,N_27349,N_26174);
xor U29941 (N_29941,N_26741,N_26015);
nor U29942 (N_29942,N_26158,N_27172);
nand U29943 (N_29943,N_26844,N_27901);
and U29944 (N_29944,N_27374,N_26313);
and U29945 (N_29945,N_26398,N_26834);
or U29946 (N_29946,N_27773,N_27341);
or U29947 (N_29947,N_26897,N_26533);
nor U29948 (N_29948,N_26960,N_27186);
and U29949 (N_29949,N_27394,N_27267);
nand U29950 (N_29950,N_27160,N_27774);
nor U29951 (N_29951,N_26923,N_27873);
xnor U29952 (N_29952,N_27284,N_27918);
nand U29953 (N_29953,N_26954,N_27789);
nor U29954 (N_29954,N_27937,N_27133);
nand U29955 (N_29955,N_27118,N_27649);
or U29956 (N_29956,N_27830,N_26057);
nand U29957 (N_29957,N_27573,N_26736);
or U29958 (N_29958,N_27215,N_26111);
nand U29959 (N_29959,N_26683,N_27266);
or U29960 (N_29960,N_27561,N_27250);
and U29961 (N_29961,N_27987,N_27542);
xnor U29962 (N_29962,N_26634,N_26855);
and U29963 (N_29963,N_26043,N_26655);
nand U29964 (N_29964,N_26502,N_26274);
nor U29965 (N_29965,N_27319,N_26348);
or U29966 (N_29966,N_26344,N_27549);
nor U29967 (N_29967,N_27586,N_26398);
and U29968 (N_29968,N_26074,N_27138);
or U29969 (N_29969,N_26722,N_26118);
xnor U29970 (N_29970,N_26574,N_27440);
and U29971 (N_29971,N_27460,N_27062);
or U29972 (N_29972,N_27711,N_27234);
nor U29973 (N_29973,N_27202,N_26195);
or U29974 (N_29974,N_26853,N_26837);
and U29975 (N_29975,N_27070,N_26547);
nand U29976 (N_29976,N_26304,N_26188);
and U29977 (N_29977,N_27550,N_26360);
nand U29978 (N_29978,N_26675,N_27973);
nand U29979 (N_29979,N_26513,N_27961);
xor U29980 (N_29980,N_27228,N_27303);
or U29981 (N_29981,N_26922,N_27729);
or U29982 (N_29982,N_26504,N_26980);
nor U29983 (N_29983,N_26377,N_27052);
or U29984 (N_29984,N_27745,N_26423);
or U29985 (N_29985,N_27507,N_26936);
or U29986 (N_29986,N_26261,N_26339);
xnor U29987 (N_29987,N_26743,N_27471);
xor U29988 (N_29988,N_26401,N_26194);
or U29989 (N_29989,N_27860,N_26189);
nor U29990 (N_29990,N_27223,N_26750);
xor U29991 (N_29991,N_26916,N_27938);
or U29992 (N_29992,N_27534,N_26232);
nor U29993 (N_29993,N_26622,N_27504);
or U29994 (N_29994,N_27084,N_27104);
nor U29995 (N_29995,N_26716,N_26280);
xor U29996 (N_29996,N_26712,N_26230);
or U29997 (N_29997,N_27018,N_26531);
xnor U29998 (N_29998,N_26121,N_27180);
xnor U29999 (N_29999,N_26088,N_26093);
nand UO_0 (O_0,N_28373,N_28405);
nor UO_1 (O_1,N_28337,N_29692);
nor UO_2 (O_2,N_28657,N_28278);
and UO_3 (O_3,N_28848,N_28133);
or UO_4 (O_4,N_28751,N_29871);
nand UO_5 (O_5,N_29261,N_29666);
nor UO_6 (O_6,N_28924,N_28069);
xor UO_7 (O_7,N_29732,N_29371);
nor UO_8 (O_8,N_28461,N_29091);
nor UO_9 (O_9,N_29569,N_28703);
nand UO_10 (O_10,N_28729,N_29635);
nand UO_11 (O_11,N_29029,N_28186);
and UO_12 (O_12,N_29075,N_29134);
xnor UO_13 (O_13,N_28377,N_28802);
xnor UO_14 (O_14,N_28594,N_29094);
nand UO_15 (O_15,N_29342,N_29586);
and UO_16 (O_16,N_29731,N_28131);
nor UO_17 (O_17,N_29744,N_28570);
nand UO_18 (O_18,N_29647,N_29778);
nor UO_19 (O_19,N_29138,N_29409);
or UO_20 (O_20,N_29950,N_29881);
and UO_21 (O_21,N_29644,N_28125);
or UO_22 (O_22,N_29378,N_28296);
and UO_23 (O_23,N_29679,N_28564);
or UO_24 (O_24,N_28578,N_29956);
nor UO_25 (O_25,N_28053,N_29764);
or UO_26 (O_26,N_28937,N_29878);
xor UO_27 (O_27,N_29452,N_29701);
nand UO_28 (O_28,N_29031,N_29769);
nor UO_29 (O_29,N_28952,N_29303);
xnor UO_30 (O_30,N_29973,N_28107);
nor UO_31 (O_31,N_29114,N_28722);
nand UO_32 (O_32,N_29350,N_28718);
and UO_33 (O_33,N_28993,N_29844);
nor UO_34 (O_34,N_28506,N_29536);
and UO_35 (O_35,N_28095,N_28119);
and UO_36 (O_36,N_28584,N_29270);
and UO_37 (O_37,N_28241,N_29977);
xor UO_38 (O_38,N_29159,N_29135);
and UO_39 (O_39,N_28326,N_28558);
xor UO_40 (O_40,N_29634,N_28240);
xnor UO_41 (O_41,N_28650,N_29018);
nor UO_42 (O_42,N_28013,N_29405);
or UO_43 (O_43,N_28372,N_29641);
and UO_44 (O_44,N_28910,N_29605);
nand UO_45 (O_45,N_29408,N_28890);
and UO_46 (O_46,N_29406,N_28451);
and UO_47 (O_47,N_29760,N_29604);
nor UO_48 (O_48,N_28124,N_29723);
or UO_49 (O_49,N_28551,N_28087);
xnor UO_50 (O_50,N_29664,N_28479);
nor UO_51 (O_51,N_29804,N_29348);
and UO_52 (O_52,N_29838,N_28995);
or UO_53 (O_53,N_29815,N_29203);
nor UO_54 (O_54,N_28212,N_28475);
and UO_55 (O_55,N_28877,N_28407);
nand UO_56 (O_56,N_29200,N_28694);
and UO_57 (O_57,N_29868,N_28839);
and UO_58 (O_58,N_28561,N_28238);
nor UO_59 (O_59,N_29932,N_29889);
xnor UO_60 (O_60,N_28484,N_29898);
nand UO_61 (O_61,N_28324,N_29063);
xnor UO_62 (O_62,N_29433,N_28901);
or UO_63 (O_63,N_28550,N_28646);
nor UO_64 (O_64,N_28332,N_28209);
nand UO_65 (O_65,N_29376,N_29118);
or UO_66 (O_66,N_28968,N_28918);
nand UO_67 (O_67,N_28930,N_29776);
xor UO_68 (O_68,N_29689,N_28437);
or UO_69 (O_69,N_28350,N_28032);
nor UO_70 (O_70,N_29227,N_28772);
xnor UO_71 (O_71,N_28992,N_29799);
nand UO_72 (O_72,N_29122,N_28971);
xor UO_73 (O_73,N_28579,N_29811);
and UO_74 (O_74,N_29296,N_28222);
nor UO_75 (O_75,N_29566,N_28560);
nor UO_76 (O_76,N_28068,N_28431);
nand UO_77 (O_77,N_28428,N_29353);
nand UO_78 (O_78,N_29110,N_29882);
xor UO_79 (O_79,N_28433,N_29958);
or UO_80 (O_80,N_28298,N_29187);
or UO_81 (O_81,N_28641,N_28526);
and UO_82 (O_82,N_28953,N_29022);
or UO_83 (O_83,N_28299,N_29347);
nand UO_84 (O_84,N_28904,N_29624);
and UO_85 (O_85,N_28368,N_28605);
xor UO_86 (O_86,N_29496,N_29596);
or UO_87 (O_87,N_29235,N_29281);
nand UO_88 (O_88,N_29730,N_29365);
nand UO_89 (O_89,N_29665,N_28002);
xnor UO_90 (O_90,N_29089,N_29740);
nor UO_91 (O_91,N_29320,N_28757);
xnor UO_92 (O_92,N_29380,N_28736);
xor UO_93 (O_93,N_29886,N_29108);
nor UO_94 (O_94,N_28935,N_29663);
or UO_95 (O_95,N_29790,N_29323);
xnor UO_96 (O_96,N_28171,N_29116);
nand UO_97 (O_97,N_28192,N_29014);
nand UO_98 (O_98,N_28986,N_28341);
and UO_99 (O_99,N_28697,N_28670);
or UO_100 (O_100,N_28949,N_28478);
and UO_101 (O_101,N_28654,N_28911);
xnor UO_102 (O_102,N_29785,N_29792);
or UO_103 (O_103,N_28861,N_29854);
nand UO_104 (O_104,N_28141,N_29971);
or UO_105 (O_105,N_28712,N_28872);
xor UO_106 (O_106,N_29160,N_28319);
and UO_107 (O_107,N_29481,N_28283);
nand UO_108 (O_108,N_29289,N_28206);
or UO_109 (O_109,N_28616,N_28794);
xor UO_110 (O_110,N_28977,N_29263);
nand UO_111 (O_111,N_29593,N_28933);
or UO_112 (O_112,N_29193,N_29923);
nor UO_113 (O_113,N_29753,N_28259);
or UO_114 (O_114,N_28025,N_29309);
nand UO_115 (O_115,N_28860,N_29787);
nor UO_116 (O_116,N_28956,N_28155);
and UO_117 (O_117,N_29775,N_28389);
xor UO_118 (O_118,N_28793,N_28342);
nor UO_119 (O_119,N_28157,N_29057);
xnor UO_120 (O_120,N_28690,N_29646);
nor UO_121 (O_121,N_28850,N_28317);
nor UO_122 (O_122,N_28940,N_28434);
nand UO_123 (O_123,N_29738,N_29630);
and UO_124 (O_124,N_29890,N_28439);
xnor UO_125 (O_125,N_29062,N_28814);
or UO_126 (O_126,N_29954,N_29828);
nand UO_127 (O_127,N_29766,N_29332);
nand UO_128 (O_128,N_28826,N_29758);
xnor UO_129 (O_129,N_28493,N_29262);
xnor UO_130 (O_130,N_28181,N_29855);
or UO_131 (O_131,N_28246,N_29123);
nor UO_132 (O_132,N_29860,N_29456);
and UO_133 (O_133,N_29251,N_29511);
nand UO_134 (O_134,N_28339,N_28029);
nand UO_135 (O_135,N_28197,N_29970);
nand UO_136 (O_136,N_28836,N_29594);
nand UO_137 (O_137,N_29508,N_29652);
or UO_138 (O_138,N_29830,N_28159);
or UO_139 (O_139,N_28281,N_28914);
or UO_140 (O_140,N_28734,N_29754);
nor UO_141 (O_141,N_28618,N_29422);
xnor UO_142 (O_142,N_29927,N_28799);
or UO_143 (O_143,N_29237,N_29478);
nor UO_144 (O_144,N_29975,N_28783);
nand UO_145 (O_145,N_28282,N_29250);
xnor UO_146 (O_146,N_29117,N_28106);
nor UO_147 (O_147,N_29367,N_28533);
and UO_148 (O_148,N_29952,N_28233);
or UO_149 (O_149,N_29391,N_28041);
and UO_150 (O_150,N_28494,N_29243);
xnor UO_151 (O_151,N_28498,N_28989);
or UO_152 (O_152,N_28689,N_28922);
nand UO_153 (O_153,N_28130,N_29249);
nand UO_154 (O_154,N_28601,N_28661);
nand UO_155 (O_155,N_29542,N_29484);
nand UO_156 (O_156,N_28936,N_29084);
xor UO_157 (O_157,N_29726,N_28396);
xor UO_158 (O_158,N_29026,N_29382);
nor UO_159 (O_159,N_28292,N_28523);
or UO_160 (O_160,N_28459,N_29209);
nor UO_161 (O_161,N_29675,N_29182);
xor UO_162 (O_162,N_29255,N_28114);
or UO_163 (O_163,N_28932,N_29247);
and UO_164 (O_164,N_28400,N_28409);
xnor UO_165 (O_165,N_28800,N_29885);
nor UO_166 (O_166,N_29561,N_28969);
or UO_167 (O_167,N_29087,N_28682);
nand UO_168 (O_168,N_29821,N_29814);
and UO_169 (O_169,N_28062,N_29239);
or UO_170 (O_170,N_28955,N_28012);
and UO_171 (O_171,N_28047,N_29434);
nand UO_172 (O_172,N_29695,N_28672);
and UO_173 (O_173,N_29042,N_28684);
or UO_174 (O_174,N_28280,N_28685);
xnor UO_175 (O_175,N_28243,N_29514);
nor UO_176 (O_176,N_28820,N_29387);
and UO_177 (O_177,N_29290,N_29384);
nor UO_178 (O_178,N_29196,N_28028);
nor UO_179 (O_179,N_29872,N_29291);
and UO_180 (O_180,N_29083,N_29590);
and UO_181 (O_181,N_28176,N_28307);
nand UO_182 (O_182,N_28146,N_28998);
nand UO_183 (O_183,N_28410,N_28340);
or UO_184 (O_184,N_29512,N_28942);
xor UO_185 (O_185,N_28030,N_29517);
or UO_186 (O_186,N_28511,N_29992);
nor UO_187 (O_187,N_29500,N_28273);
nor UO_188 (O_188,N_29071,N_29749);
nor UO_189 (O_189,N_28815,N_28035);
nand UO_190 (O_190,N_28276,N_29276);
or UO_191 (O_191,N_28709,N_28929);
xnor UO_192 (O_192,N_28760,N_29498);
or UO_193 (O_193,N_29964,N_28336);
and UO_194 (O_194,N_29806,N_28122);
and UO_195 (O_195,N_28200,N_28158);
or UO_196 (O_196,N_29469,N_28809);
nand UO_197 (O_197,N_28797,N_29437);
or UO_198 (O_198,N_28662,N_28160);
and UO_199 (O_199,N_29836,N_29027);
nand UO_200 (O_200,N_28948,N_28589);
xnor UO_201 (O_201,N_28780,N_29941);
nand UO_202 (O_202,N_29951,N_28215);
nor UO_203 (O_203,N_29066,N_29366);
xnor UO_204 (O_204,N_29213,N_28590);
or UO_205 (O_205,N_28313,N_29313);
nand UO_206 (O_206,N_29254,N_29462);
and UO_207 (O_207,N_29712,N_29448);
xor UO_208 (O_208,N_28086,N_28825);
xor UO_209 (O_209,N_28333,N_28897);
nand UO_210 (O_210,N_29651,N_28599);
or UO_211 (O_211,N_28597,N_28194);
nand UO_212 (O_212,N_29155,N_29832);
nand UO_213 (O_213,N_29460,N_28142);
or UO_214 (O_214,N_29341,N_29335);
xnor UO_215 (O_215,N_29390,N_29172);
nand UO_216 (O_216,N_29673,N_28416);
or UO_217 (O_217,N_28453,N_28811);
nor UO_218 (O_218,N_28330,N_28738);
nand UO_219 (O_219,N_28521,N_29574);
nand UO_220 (O_220,N_28457,N_29761);
nand UO_221 (O_221,N_29346,N_28678);
and UO_222 (O_222,N_29592,N_28505);
and UO_223 (O_223,N_29337,N_29888);
and UO_224 (O_224,N_28585,N_28756);
and UO_225 (O_225,N_28345,N_28322);
nor UO_226 (O_226,N_29745,N_28039);
nor UO_227 (O_227,N_28666,N_29642);
or UO_228 (O_228,N_28656,N_29113);
or UO_229 (O_229,N_29924,N_28321);
nand UO_230 (O_230,N_28353,N_29614);
xnor UO_231 (O_231,N_28379,N_29611);
xor UO_232 (O_232,N_29615,N_29315);
nor UO_233 (O_233,N_28167,N_29685);
nor UO_234 (O_234,N_29497,N_29788);
nand UO_235 (O_235,N_29455,N_28175);
nor UO_236 (O_236,N_29426,N_29963);
nand UO_237 (O_237,N_28831,N_29714);
nor UO_238 (O_238,N_28027,N_29389);
nor UO_239 (O_239,N_29993,N_28294);
nand UO_240 (O_240,N_29283,N_29189);
nor UO_241 (O_241,N_29774,N_29333);
xnor UO_242 (O_242,N_28928,N_29300);
and UO_243 (O_243,N_29805,N_29543);
xor UO_244 (O_244,N_28329,N_28403);
nand UO_245 (O_245,N_29051,N_28824);
nand UO_246 (O_246,N_28821,N_29495);
nand UO_247 (O_247,N_29706,N_28126);
nor UO_248 (O_248,N_28978,N_29120);
and UO_249 (O_249,N_28205,N_28893);
nand UO_250 (O_250,N_28143,N_28208);
nand UO_251 (O_251,N_29866,N_28943);
or UO_252 (O_252,N_28745,N_28249);
or UO_253 (O_253,N_29962,N_29779);
and UO_254 (O_254,N_28213,N_29102);
and UO_255 (O_255,N_29528,N_28787);
nor UO_256 (O_256,N_28302,N_29076);
and UO_257 (O_257,N_29602,N_29232);
nand UO_258 (O_258,N_28174,N_29669);
or UO_259 (O_259,N_29539,N_28442);
nand UO_260 (O_260,N_28753,N_28856);
xor UO_261 (O_261,N_29677,N_28752);
nor UO_262 (O_262,N_28941,N_28145);
xor UO_263 (O_263,N_29648,N_28499);
nand UO_264 (O_264,N_28097,N_29450);
xnor UO_265 (O_265,N_29955,N_28868);
and UO_266 (O_266,N_28853,N_28483);
nand UO_267 (O_267,N_29395,N_29304);
nor UO_268 (O_268,N_28015,N_28885);
and UO_269 (O_269,N_29873,N_28362);
and UO_270 (O_270,N_29865,N_28845);
xnor UO_271 (O_271,N_28996,N_29229);
and UO_272 (O_272,N_28717,N_28369);
and UO_273 (O_273,N_29795,N_28529);
and UO_274 (O_274,N_28769,N_29430);
or UO_275 (O_275,N_29680,N_29894);
xnor UO_276 (O_276,N_28653,N_29241);
and UO_277 (O_277,N_29204,N_28128);
and UO_278 (O_278,N_29285,N_29912);
nand UO_279 (O_279,N_29392,N_29555);
or UO_280 (O_280,N_29937,N_29717);
xor UO_281 (O_281,N_29052,N_28468);
and UO_282 (O_282,N_28279,N_29710);
nand UO_283 (O_283,N_28303,N_29631);
nand UO_284 (O_284,N_28436,N_28184);
xor UO_285 (O_285,N_28572,N_28401);
nor UO_286 (O_286,N_29340,N_28083);
or UO_287 (O_287,N_28816,N_29576);
nor UO_288 (O_288,N_29794,N_29326);
xor UO_289 (O_289,N_29907,N_28520);
and UO_290 (O_290,N_29506,N_28406);
nand UO_291 (O_291,N_28554,N_29183);
or UO_292 (O_292,N_29741,N_28805);
or UO_293 (O_293,N_29041,N_29980);
and UO_294 (O_294,N_28180,N_28621);
xnor UO_295 (O_295,N_29253,N_29765);
or UO_296 (O_296,N_28611,N_28889);
nor UO_297 (O_297,N_29633,N_28471);
nor UO_298 (O_298,N_28228,N_29791);
nand UO_299 (O_299,N_29109,N_29823);
xor UO_300 (O_300,N_29097,N_28349);
nor UO_301 (O_301,N_28044,N_29899);
or UO_302 (O_302,N_29718,N_29208);
and UO_303 (O_303,N_29439,N_29150);
nor UO_304 (O_304,N_28144,N_28443);
nand UO_305 (O_305,N_28038,N_28739);
nand UO_306 (O_306,N_28883,N_29659);
or UO_307 (O_307,N_29021,N_28003);
nand UO_308 (O_308,N_29067,N_29394);
nor UO_309 (O_309,N_28876,N_29550);
xnor UO_310 (O_310,N_29529,N_28104);
or UO_311 (O_311,N_28430,N_28925);
or UO_312 (O_312,N_29880,N_29314);
nand UO_313 (O_313,N_29545,N_29195);
or UO_314 (O_314,N_29330,N_28573);
nor UO_315 (O_315,N_28545,N_29662);
nor UO_316 (O_316,N_28840,N_29006);
and UO_317 (O_317,N_29181,N_29672);
and UO_318 (O_318,N_29999,N_28927);
nand UO_319 (O_319,N_29709,N_29533);
nor UO_320 (O_320,N_29466,N_29928);
or UO_321 (O_321,N_29747,N_29085);
nand UO_322 (O_322,N_29361,N_28429);
and UO_323 (O_323,N_29997,N_29107);
xor UO_324 (O_324,N_29930,N_28659);
nor UO_325 (O_325,N_29205,N_29104);
and UO_326 (O_326,N_28852,N_28067);
xor UO_327 (O_327,N_29535,N_29683);
or UO_328 (O_328,N_28447,N_28587);
nand UO_329 (O_329,N_29591,N_28586);
nand UO_330 (O_330,N_28701,N_29442);
nand UO_331 (O_331,N_29445,N_28204);
nand UO_332 (O_332,N_28510,N_28488);
nor UO_333 (O_333,N_28151,N_28528);
nor UO_334 (O_334,N_28066,N_28486);
and UO_335 (O_335,N_28834,N_29064);
nor UO_336 (O_336,N_29186,N_28867);
nor UO_337 (O_337,N_28994,N_28542);
nor UO_338 (O_338,N_28301,N_28490);
xor UO_339 (O_339,N_29435,N_29280);
nand UO_340 (O_340,N_28531,N_29850);
xor UO_341 (O_341,N_29003,N_28424);
and UO_342 (O_342,N_29523,N_28256);
xor UO_343 (O_343,N_29998,N_29657);
xnor UO_344 (O_344,N_28822,N_29119);
or UO_345 (O_345,N_28093,N_28583);
nor UO_346 (O_346,N_28912,N_29972);
or UO_347 (O_347,N_28008,N_28365);
xnor UO_348 (O_348,N_29299,N_28525);
xnor UO_349 (O_349,N_29226,N_28325);
xor UO_350 (O_350,N_28726,N_28537);
nor UO_351 (O_351,N_29059,N_28593);
nand UO_352 (O_352,N_28767,N_28765);
or UO_353 (O_353,N_29883,N_29755);
xnor UO_354 (O_354,N_28744,N_28073);
nand UO_355 (O_355,N_28458,N_28908);
nor UO_356 (O_356,N_28612,N_28909);
and UO_357 (O_357,N_28713,N_29807);
or UO_358 (O_358,N_28725,N_28707);
and UO_359 (O_359,N_28818,N_29982);
and UO_360 (O_360,N_28556,N_28980);
nand UO_361 (O_361,N_29767,N_29893);
xnor UO_362 (O_362,N_29198,N_29967);
xnor UO_363 (O_363,N_28183,N_29820);
or UO_364 (O_364,N_29548,N_28134);
nor UO_365 (O_365,N_29218,N_29736);
and UO_366 (O_366,N_29349,N_29681);
nor UO_367 (O_367,N_29658,N_29454);
and UO_368 (O_368,N_29816,N_28636);
or UO_369 (O_369,N_28982,N_28764);
or UO_370 (O_370,N_28449,N_29343);
or UO_371 (O_371,N_29989,N_28177);
xnor UO_372 (O_372,N_29149,N_28919);
or UO_373 (O_373,N_28463,N_28637);
xor UO_374 (O_374,N_29260,N_29061);
nor UO_375 (O_375,N_29507,N_28762);
xor UO_376 (O_376,N_29271,N_29400);
nand UO_377 (O_377,N_28394,N_28951);
or UO_378 (O_378,N_29485,N_28371);
xor UO_379 (O_379,N_28673,N_29038);
or UO_380 (O_380,N_28984,N_28830);
and UO_381 (O_381,N_29474,N_28123);
nand UO_382 (O_382,N_28148,N_28967);
xor UO_383 (O_383,N_29733,N_28161);
and UO_384 (O_384,N_28733,N_29581);
nand UO_385 (O_385,N_29322,N_29040);
or UO_386 (O_386,N_29177,N_28231);
nor UO_387 (O_387,N_28366,N_29465);
and UO_388 (O_388,N_28864,N_29638);
nand UO_389 (O_389,N_28109,N_29098);
nor UO_390 (O_390,N_28380,N_29471);
nand UO_391 (O_391,N_28019,N_29050);
xor UO_392 (O_392,N_29070,N_29278);
xnor UO_393 (O_393,N_28837,N_28959);
nor UO_394 (O_394,N_29417,N_29655);
and UO_395 (O_395,N_28539,N_29476);
or UO_396 (O_396,N_28253,N_29024);
or UO_397 (O_397,N_28147,N_29704);
and UO_398 (O_398,N_28414,N_28346);
or UO_399 (O_399,N_28746,N_28859);
nand UO_400 (O_400,N_29944,N_28629);
and UO_401 (O_401,N_28724,N_29170);
or UO_402 (O_402,N_29707,N_28269);
and UO_403 (O_403,N_29858,N_28308);
xnor UO_404 (O_404,N_28686,N_29833);
xnor UO_405 (O_405,N_28367,N_29725);
and UO_406 (O_406,N_28440,N_29140);
and UO_407 (O_407,N_28732,N_28973);
and UO_408 (O_408,N_29876,N_29922);
or UO_409 (O_409,N_28644,N_28504);
xor UO_410 (O_410,N_28309,N_28896);
nor UO_411 (O_411,N_28633,N_28397);
nand UO_412 (O_412,N_28057,N_29988);
nor UO_413 (O_413,N_29424,N_28477);
and UO_414 (O_414,N_28966,N_29479);
xor UO_415 (O_415,N_29599,N_29169);
xor UO_416 (O_416,N_28515,N_28507);
xnor UO_417 (O_417,N_28121,N_28242);
xor UO_418 (O_418,N_29921,N_28516);
and UO_419 (O_419,N_28255,N_28105);
or UO_420 (O_420,N_28402,N_28214);
xor UO_421 (O_421,N_29046,N_28454);
xnor UO_422 (O_422,N_29151,N_29763);
nor UO_423 (O_423,N_29653,N_29115);
nor UO_424 (O_424,N_28944,N_28356);
nor UO_425 (O_425,N_29835,N_29617);
nor UO_426 (O_426,N_28318,N_28761);
nand UO_427 (O_427,N_29438,N_29661);
xnor UO_428 (O_428,N_28513,N_29938);
xor UO_429 (O_429,N_29579,N_29165);
xnor UO_430 (O_430,N_28750,N_29636);
nor UO_431 (O_431,N_29748,N_28687);
xnor UO_432 (O_432,N_28037,N_29489);
nor UO_433 (O_433,N_28985,N_28306);
nand UO_434 (O_434,N_29345,N_29443);
nand UO_435 (O_435,N_28335,N_28603);
nand UO_436 (O_436,N_29307,N_29933);
xor UO_437 (O_437,N_28775,N_28862);
nand UO_438 (O_438,N_28879,N_28884);
nand UO_439 (O_439,N_28404,N_29622);
nand UO_440 (O_440,N_29054,N_29477);
nand UO_441 (O_441,N_29722,N_28487);
nand UO_442 (O_442,N_28898,N_28216);
xor UO_443 (O_443,N_29267,N_28011);
xnor UO_444 (O_444,N_28153,N_29179);
or UO_445 (O_445,N_28700,N_29292);
or UO_446 (O_446,N_29246,N_28846);
and UO_447 (O_447,N_28323,N_28527);
or UO_448 (O_448,N_29377,N_28934);
xor UO_449 (O_449,N_29991,N_28286);
xor UO_450 (O_450,N_28524,N_28894);
nand UO_451 (O_451,N_29789,N_28835);
or UO_452 (O_452,N_28354,N_29800);
or UO_453 (O_453,N_28481,N_28849);
xor UO_454 (O_454,N_29441,N_28796);
nor UO_455 (O_455,N_29128,N_29667);
and UO_456 (O_456,N_29813,N_29143);
or UO_457 (O_457,N_29564,N_28263);
nand UO_458 (O_458,N_29568,N_29487);
nand UO_459 (O_459,N_28203,N_28696);
or UO_460 (O_460,N_29161,N_28748);
nand UO_461 (O_461,N_29793,N_28981);
nand UO_462 (O_462,N_28168,N_28310);
nor UO_463 (O_463,N_29856,N_28863);
or UO_464 (O_464,N_28500,N_29475);
nand UO_465 (O_465,N_28680,N_28359);
and UO_466 (O_466,N_29978,N_29065);
xor UO_467 (O_467,N_29095,N_28129);
nand UO_468 (O_468,N_28024,N_29688);
or UO_469 (O_469,N_29308,N_29570);
nor UO_470 (O_470,N_29185,N_28234);
nor UO_471 (O_471,N_29004,N_28731);
or UO_472 (O_472,N_29483,N_28219);
nor UO_473 (O_473,N_29124,N_29214);
nand UO_474 (O_474,N_28284,N_28888);
nor UO_475 (O_475,N_29310,N_29640);
xor UO_476 (O_476,N_29781,N_29735);
and UO_477 (O_477,N_28370,N_29413);
nor UO_478 (O_478,N_28508,N_28311);
nand UO_479 (O_479,N_28838,N_28266);
nand UO_480 (O_480,N_29412,N_29656);
xor UO_481 (O_481,N_28223,N_28625);
nand UO_482 (O_482,N_29874,N_28444);
nor UO_483 (O_483,N_29534,N_29895);
xor UO_484 (O_484,N_28950,N_29184);
nor UO_485 (O_485,N_29224,N_29520);
nand UO_486 (O_486,N_29399,N_28546);
xnor UO_487 (O_487,N_29163,N_29650);
xnor UO_488 (O_488,N_28999,N_28262);
xnor UO_489 (O_489,N_28169,N_28391);
xor UO_490 (O_490,N_28875,N_28679);
or UO_491 (O_491,N_29266,N_28006);
nor UO_492 (O_492,N_28399,N_28348);
or UO_493 (O_493,N_29277,N_28706);
xor UO_494 (O_494,N_28991,N_29002);
and UO_495 (O_495,N_28221,N_28381);
or UO_496 (O_496,N_29589,N_28923);
nand UO_497 (O_497,N_29691,N_29884);
and UO_498 (O_498,N_29803,N_29903);
or UO_499 (O_499,N_29859,N_28568);
nand UO_500 (O_500,N_28602,N_29086);
nand UO_501 (O_501,N_28163,N_29136);
and UO_502 (O_502,N_28608,N_28702);
nand UO_503 (O_503,N_28017,N_28534);
nand UO_504 (O_504,N_29510,N_28046);
xor UO_505 (O_505,N_28363,N_29969);
xor UO_506 (O_506,N_28492,N_29188);
and UO_507 (O_507,N_29558,N_29176);
nor UO_508 (O_508,N_29711,N_28947);
nor UO_509 (O_509,N_28913,N_29374);
or UO_510 (O_510,N_29913,N_29911);
nor UO_511 (O_511,N_28624,N_28334);
or UO_512 (O_512,N_29269,N_28675);
nand UO_513 (O_513,N_29137,N_28668);
nand UO_514 (O_514,N_28544,N_29034);
xor UO_515 (O_515,N_28865,N_28622);
nor UO_516 (O_516,N_28833,N_29777);
xor UO_517 (O_517,N_29696,N_29298);
or UO_518 (O_518,N_28828,N_28084);
xnor UO_519 (O_519,N_28275,N_29429);
and UO_520 (O_520,N_29639,N_28792);
and UO_521 (O_521,N_29142,N_29457);
xor UO_522 (O_522,N_28899,N_28615);
xnor UO_523 (O_523,N_29049,N_29228);
nor UO_524 (O_524,N_28020,N_29762);
nand UO_525 (O_525,N_28728,N_29464);
xor UO_526 (O_526,N_29105,N_28827);
nand UO_527 (O_527,N_29379,N_28620);
and UO_528 (O_528,N_29863,N_29920);
xor UO_529 (O_529,N_28462,N_28788);
nand UO_530 (O_530,N_29618,N_29219);
nor UO_531 (O_531,N_29017,N_29750);
xnor UO_532 (O_532,N_28411,N_29311);
and UO_533 (O_533,N_28387,N_29047);
nand UO_534 (O_534,N_29654,N_28248);
or UO_535 (O_535,N_28581,N_28552);
and UO_536 (O_536,N_29572,N_29771);
or UO_537 (O_537,N_28395,N_28001);
or UO_538 (O_538,N_29601,N_28665);
and UO_539 (O_539,N_28580,N_28218);
or UO_540 (O_540,N_28755,N_29431);
nor UO_541 (O_541,N_29575,N_28054);
or UO_542 (O_542,N_29223,N_28210);
or UO_543 (O_543,N_28789,N_29393);
nand UO_544 (O_544,N_28199,N_29995);
nor UO_545 (O_545,N_29106,N_28051);
nand UO_546 (O_546,N_29567,N_29428);
nand UO_547 (O_547,N_29547,N_29588);
and UO_548 (O_548,N_28450,N_28591);
and UO_549 (O_549,N_29949,N_28305);
and UO_550 (O_550,N_28768,N_28642);
nor UO_551 (O_551,N_29453,N_29363);
or UO_552 (O_552,N_29019,N_28136);
or UO_553 (O_553,N_29446,N_29145);
xnor UO_554 (O_554,N_29974,N_28819);
or UO_555 (O_555,N_29861,N_29557);
and UO_556 (O_556,N_29867,N_28031);
nor UO_557 (O_557,N_29053,N_29166);
nand UO_558 (O_558,N_29822,N_29282);
nand UO_559 (O_559,N_28466,N_29996);
nand UO_560 (O_560,N_28426,N_28979);
or UO_561 (O_561,N_29199,N_28094);
nor UO_562 (O_562,N_29519,N_29404);
xor UO_563 (O_563,N_28331,N_29334);
or UO_564 (O_564,N_29908,N_28727);
nand UO_565 (O_565,N_29501,N_29734);
or UO_566 (O_566,N_28771,N_28026);
or UO_567 (O_567,N_29147,N_28096);
nand UO_568 (O_568,N_28217,N_28740);
nor UO_569 (O_569,N_28588,N_28251);
nand UO_570 (O_570,N_28361,N_29001);
nor UO_571 (O_571,N_29968,N_29058);
xor UO_572 (O_572,N_29449,N_28598);
nand UO_573 (O_573,N_29925,N_29705);
and UO_574 (O_574,N_29981,N_28351);
nor UO_575 (O_575,N_29410,N_28080);
and UO_576 (O_576,N_29225,N_29957);
nor UO_577 (O_577,N_28419,N_28101);
xnor UO_578 (O_578,N_28632,N_29167);
xor UO_579 (O_579,N_28274,N_29211);
xnor UO_580 (O_580,N_28237,N_28674);
or UO_581 (O_581,N_29402,N_29286);
or UO_582 (O_582,N_28741,N_29328);
or UO_583 (O_583,N_28268,N_29467);
or UO_584 (O_584,N_29959,N_28055);
or UO_585 (O_585,N_28716,N_28548);
and UO_586 (O_586,N_29154,N_28220);
nor UO_587 (O_587,N_29397,N_29486);
or UO_588 (O_588,N_28881,N_29849);
nor UO_589 (O_589,N_29416,N_29383);
nand UO_590 (O_590,N_29096,N_28671);
xnor UO_591 (O_591,N_29129,N_28412);
nor UO_592 (O_592,N_29621,N_28711);
and UO_593 (O_593,N_29676,N_29060);
nor UO_594 (O_594,N_29005,N_29537);
nor UO_595 (O_595,N_28777,N_29491);
nor UO_596 (O_596,N_29197,N_28817);
nor UO_597 (O_597,N_29612,N_28997);
xor UO_598 (O_598,N_28074,N_28343);
or UO_599 (O_599,N_29532,N_28058);
nand UO_600 (O_600,N_29716,N_28116);
xor UO_601 (O_601,N_28392,N_29583);
xor UO_602 (O_602,N_29357,N_29111);
or UO_603 (O_603,N_29220,N_28514);
nand UO_604 (O_604,N_28502,N_29207);
xnor UO_605 (O_605,N_29628,N_29926);
xor UO_606 (O_606,N_28376,N_29942);
and UO_607 (O_607,N_29231,N_28415);
nand UO_608 (O_608,N_28735,N_28149);
nor UO_609 (O_609,N_28645,N_28315);
or UO_610 (O_610,N_29607,N_28596);
nand UO_611 (O_611,N_28631,N_29984);
nor UO_612 (O_612,N_29620,N_29013);
xnor UO_613 (O_613,N_28236,N_28569);
and UO_614 (O_614,N_28658,N_29273);
nor UO_615 (O_615,N_28651,N_29055);
nand UO_616 (O_616,N_29112,N_28166);
xnor UO_617 (O_617,N_28829,N_28988);
and UO_618 (O_618,N_29192,N_29202);
nand UO_619 (O_619,N_29423,N_28921);
and UO_620 (O_620,N_29259,N_29546);
and UO_621 (O_621,N_29221,N_28915);
xor UO_622 (O_622,N_29931,N_29164);
or UO_623 (O_623,N_28961,N_28976);
nand UO_624 (O_624,N_29783,N_28071);
and UO_625 (O_625,N_28737,N_28010);
xor UO_626 (O_626,N_28139,N_28785);
and UO_627 (O_627,N_29746,N_28352);
nor UO_628 (O_628,N_29162,N_28417);
nor UO_629 (O_629,N_28907,N_28823);
nand UO_630 (O_630,N_29918,N_29773);
xnor UO_631 (O_631,N_28791,N_28582);
nor UO_632 (O_632,N_28277,N_28547);
xor UO_633 (O_633,N_29101,N_28108);
or UO_634 (O_634,N_28938,N_28473);
nor UO_635 (O_635,N_29573,N_29362);
xor UO_636 (O_636,N_29801,N_29216);
and UO_637 (O_637,N_29036,N_28009);
and UO_638 (O_638,N_28188,N_29007);
nand UO_639 (O_639,N_29470,N_29339);
nor UO_640 (O_640,N_28132,N_29461);
xnor UO_641 (O_641,N_28446,N_28784);
and UO_642 (O_642,N_29072,N_28851);
nand UO_643 (O_643,N_28638,N_28619);
nor UO_644 (O_644,N_29915,N_29752);
and UO_645 (O_645,N_28489,N_29279);
and UO_646 (O_646,N_28699,N_29853);
xor UO_647 (O_647,N_29302,N_29274);
nor UO_648 (O_648,N_28413,N_29468);
nand UO_649 (O_649,N_29864,N_29321);
xor UO_650 (O_650,N_29902,N_29201);
xnor UO_651 (O_651,N_29919,N_28781);
and UO_652 (O_652,N_29619,N_28347);
nor UO_653 (O_653,N_28808,N_28627);
nand UO_654 (O_654,N_28187,N_28964);
nor UO_655 (O_655,N_28871,N_29358);
or UO_656 (O_656,N_28782,N_29606);
or UO_657 (O_657,N_28643,N_28398);
or UO_658 (O_658,N_29632,N_29324);
nand UO_659 (O_659,N_28190,N_29540);
and UO_660 (O_660,N_29180,N_28076);
nor UO_661 (O_661,N_28100,N_29088);
and UO_662 (O_662,N_28110,N_28448);
or UO_663 (O_663,N_29472,N_28975);
and UO_664 (O_664,N_29671,N_29940);
or UO_665 (O_665,N_28543,N_29016);
and UO_666 (O_666,N_29493,N_29258);
and UO_667 (O_667,N_28202,N_28247);
nor UO_668 (O_668,N_29396,N_28014);
xnor UO_669 (O_669,N_29505,N_28470);
xor UO_670 (O_670,N_28945,N_29598);
or UO_671 (O_671,N_28880,N_29458);
xnor UO_672 (O_672,N_29906,N_29073);
nor UO_673 (O_673,N_28747,N_29157);
nor UO_674 (O_674,N_29336,N_29503);
or UO_675 (O_675,N_28099,N_28072);
xor UO_676 (O_676,N_28295,N_29713);
or UO_677 (O_677,N_28795,N_28855);
nor UO_678 (O_678,N_29488,N_29325);
and UO_679 (O_679,N_29236,N_28007);
nand UO_680 (O_680,N_29432,N_29090);
and UO_681 (O_681,N_29824,N_29444);
nor UO_682 (O_682,N_28021,N_28338);
and UO_683 (O_683,N_29000,N_29174);
or UO_684 (O_684,N_28892,N_28847);
xnor UO_685 (O_685,N_29979,N_29877);
nor UO_686 (O_686,N_28060,N_29295);
nand UO_687 (O_687,N_29043,N_29414);
nand UO_688 (O_688,N_29553,N_29943);
or UO_689 (O_689,N_29896,N_28495);
or UO_690 (O_690,N_29562,N_29693);
or UO_691 (O_691,N_28691,N_29551);
nor UO_692 (O_692,N_28254,N_29351);
nand UO_693 (O_693,N_29039,N_29715);
nor UO_694 (O_694,N_28467,N_28052);
xnor UO_695 (O_695,N_29329,N_28882);
nand UO_696 (O_696,N_29388,N_28891);
xor UO_697 (O_697,N_28806,N_28469);
xnor UO_698 (O_698,N_29171,N_28595);
nand UO_699 (O_699,N_29316,N_28749);
nand UO_700 (O_700,N_29194,N_29025);
and UO_701 (O_701,N_29152,N_29851);
or UO_702 (O_702,N_29146,N_29780);
or UO_703 (O_703,N_28522,N_29288);
and UO_704 (O_704,N_29841,N_28669);
xnor UO_705 (O_705,N_29530,N_28535);
or UO_706 (O_706,N_28360,N_29834);
nand UO_707 (O_707,N_29284,N_29077);
and UO_708 (O_708,N_28258,N_29133);
nand UO_709 (O_709,N_29905,N_28115);
or UO_710 (O_710,N_28705,N_29595);
nand UO_711 (O_711,N_29264,N_28267);
xor UO_712 (O_712,N_29699,N_28456);
nor UO_713 (O_713,N_28695,N_28375);
or UO_714 (O_714,N_28610,N_29629);
and UO_715 (O_715,N_28090,N_28042);
nor UO_716 (O_716,N_29516,N_29265);
nand UO_717 (O_717,N_28162,N_28111);
or UO_718 (O_718,N_29862,N_28704);
and UO_719 (O_719,N_28900,N_29757);
and UO_720 (O_720,N_29668,N_29369);
or UO_721 (O_721,N_29272,N_28628);
and UO_722 (O_722,N_28465,N_28045);
nand UO_723 (O_723,N_28607,N_28574);
and UO_724 (O_724,N_29825,N_29032);
xnor UO_725 (O_725,N_29987,N_28623);
and UO_726 (O_726,N_28297,N_29625);
or UO_727 (O_727,N_29756,N_29010);
nand UO_728 (O_728,N_29153,N_29244);
nor UO_729 (O_729,N_28858,N_29421);
nor UO_730 (O_730,N_28983,N_28320);
nand UO_731 (O_731,N_28250,N_29141);
nor UO_732 (O_732,N_28571,N_28719);
nand UO_733 (O_733,N_29518,N_29103);
xnor UO_734 (O_734,N_29306,N_28113);
or UO_735 (O_735,N_28427,N_28137);
or UO_736 (O_736,N_28640,N_28265);
nor UO_737 (O_737,N_28832,N_28804);
and UO_738 (O_738,N_28290,N_29875);
xnor UO_739 (O_739,N_29100,N_28441);
nand UO_740 (O_740,N_29802,N_29772);
or UO_741 (O_741,N_29660,N_29427);
and UO_742 (O_742,N_28708,N_28195);
nand UO_743 (O_743,N_29020,N_29240);
or UO_744 (O_744,N_28150,N_28316);
and UO_745 (O_745,N_29904,N_28165);
nor UO_746 (O_746,N_29737,N_28807);
xor UO_747 (O_747,N_28917,N_28390);
nand UO_748 (O_748,N_29580,N_29645);
and UO_749 (O_749,N_29698,N_29009);
or UO_750 (O_750,N_28606,N_29419);
xor UO_751 (O_751,N_28358,N_29797);
xnor UO_752 (O_752,N_28786,N_28648);
nand UO_753 (O_753,N_28089,N_28617);
or UO_754 (O_754,N_28519,N_28423);
xor UO_755 (O_755,N_28482,N_29509);
or UO_756 (O_756,N_28422,N_28509);
and UO_757 (O_757,N_28344,N_29541);
nor UO_758 (O_758,N_29840,N_28714);
and UO_759 (O_759,N_29571,N_29947);
xor UO_760 (O_760,N_28232,N_29728);
and UO_761 (O_761,N_29577,N_29385);
and UO_762 (O_762,N_29727,N_28257);
xnor UO_763 (O_763,N_28497,N_28559);
nor UO_764 (O_764,N_29817,N_28474);
nand UO_765 (O_765,N_29494,N_29035);
nor UO_766 (O_766,N_29929,N_28312);
nand UO_767 (O_767,N_29770,N_29768);
xnor UO_768 (O_768,N_29934,N_28225);
xnor UO_769 (O_769,N_28655,N_28196);
or UO_770 (O_770,N_28743,N_28721);
xor UO_771 (O_771,N_28842,N_28532);
nor UO_772 (O_772,N_29897,N_29554);
and UO_773 (O_773,N_29502,N_28098);
nand UO_774 (O_774,N_28530,N_28271);
nor UO_775 (O_775,N_28464,N_28103);
or UO_776 (O_776,N_28903,N_29852);
and UO_777 (O_777,N_28112,N_29403);
xor UO_778 (O_778,N_29079,N_28634);
nand UO_779 (O_779,N_28566,N_29513);
nor UO_780 (O_780,N_28229,N_28287);
xor UO_781 (O_781,N_29724,N_29175);
and UO_782 (O_782,N_29674,N_29670);
xor UO_783 (O_783,N_29600,N_29965);
nor UO_784 (O_784,N_29178,N_29584);
nor UO_785 (O_785,N_28460,N_29275);
nand UO_786 (O_786,N_29011,N_28393);
nor UO_787 (O_787,N_28517,N_29415);
xor UO_788 (O_788,N_28920,N_28557);
xor UO_789 (O_789,N_29407,N_29686);
and UO_790 (O_790,N_28018,N_29212);
or UO_791 (O_791,N_28902,N_29869);
or UO_792 (O_792,N_28285,N_28435);
nor UO_793 (O_793,N_28803,N_28065);
nor UO_794 (O_794,N_28189,N_28120);
nor UO_795 (O_795,N_29044,N_28843);
nand UO_796 (O_796,N_29578,N_28245);
nand UO_797 (O_797,N_29819,N_29936);
or UO_798 (O_798,N_28926,N_28364);
xnor UO_799 (O_799,N_28178,N_28485);
xnor UO_800 (O_800,N_29368,N_28518);
and UO_801 (O_801,N_29515,N_29917);
and UO_802 (O_802,N_28425,N_29798);
nand UO_803 (O_803,N_28043,N_29843);
and UO_804 (O_804,N_28774,N_29729);
nor UO_805 (O_805,N_29751,N_28562);
or UO_806 (O_806,N_29909,N_28939);
and UO_807 (O_807,N_28990,N_28567);
nand UO_808 (O_808,N_29827,N_28873);
and UO_809 (O_809,N_29784,N_29626);
or UO_810 (O_810,N_28085,N_28496);
nor UO_811 (O_811,N_28235,N_29826);
and UO_812 (O_812,N_29268,N_28421);
nand UO_813 (O_813,N_28754,N_29191);
nor UO_814 (O_814,N_29125,N_28639);
or UO_815 (O_815,N_28575,N_28355);
nand UO_816 (O_816,N_29703,N_29356);
and UO_817 (O_817,N_28022,N_29891);
or UO_818 (O_818,N_29447,N_28118);
or UO_819 (O_819,N_29845,N_28059);
nand UO_820 (O_820,N_29870,N_28857);
nand UO_821 (O_821,N_29364,N_29623);
and UO_822 (O_822,N_28385,N_29582);
and UO_823 (O_823,N_28541,N_29948);
nand UO_824 (O_824,N_28081,N_29012);
nor UO_825 (O_825,N_28244,N_29708);
or UO_826 (O_826,N_29099,N_28801);
or UO_827 (O_827,N_28565,N_28878);
nand UO_828 (O_828,N_28683,N_28005);
and UO_829 (O_829,N_29983,N_29526);
and UO_830 (O_830,N_29525,N_28357);
nor UO_831 (O_831,N_29690,N_29786);
and UO_832 (O_832,N_28327,N_29451);
nand UO_833 (O_833,N_28382,N_29092);
or UO_834 (O_834,N_28386,N_29521);
nand UO_835 (O_835,N_28663,N_29045);
nand UO_836 (O_836,N_29720,N_28048);
or UO_837 (O_837,N_28264,N_28810);
and UO_838 (O_838,N_29809,N_28773);
xor UO_839 (O_839,N_28715,N_28270);
nand UO_840 (O_840,N_29354,N_28962);
nand UO_841 (O_841,N_29037,N_29082);
nor UO_842 (O_842,N_28692,N_29846);
xnor UO_843 (O_843,N_29234,N_28958);
nor UO_844 (O_844,N_29961,N_28201);
and UO_845 (O_845,N_28652,N_29960);
and UO_846 (O_846,N_29531,N_28779);
nand UO_847 (O_847,N_29837,N_29459);
and UO_848 (O_848,N_29742,N_29976);
and UO_849 (O_849,N_28040,N_29945);
or UO_850 (O_850,N_29210,N_28886);
xor UO_851 (O_851,N_29721,N_29482);
or UO_852 (O_852,N_29048,N_28577);
and UO_853 (O_853,N_28647,N_28538);
nor UO_854 (O_854,N_29490,N_29609);
xor UO_855 (O_855,N_29375,N_29613);
xor UO_856 (O_856,N_28156,N_29847);
or UO_857 (O_857,N_28770,N_29857);
nand UO_858 (O_858,N_28170,N_28869);
nand UO_859 (O_859,N_29687,N_29700);
nand UO_860 (O_860,N_29144,N_29318);
nor UO_861 (O_861,N_29697,N_28866);
and UO_862 (O_862,N_28844,N_28252);
and UO_863 (O_863,N_28905,N_29739);
nor UO_864 (O_864,N_29327,N_29440);
xnor UO_865 (O_865,N_29033,N_29215);
nand UO_866 (O_866,N_29879,N_29565);
nand UO_867 (O_867,N_28676,N_29217);
xor UO_868 (O_868,N_28501,N_28491);
nand UO_869 (O_869,N_29293,N_28445);
nand UO_870 (O_870,N_28895,N_29603);
nor UO_871 (O_871,N_29069,N_29829);
and UO_872 (O_872,N_28536,N_29544);
xnor UO_873 (O_873,N_28016,N_29242);
and UO_874 (O_874,N_28224,N_28193);
nor UO_875 (O_875,N_28776,N_28512);
or UO_876 (O_876,N_28763,N_29222);
nand UO_877 (O_877,N_29608,N_29678);
nor UO_878 (O_878,N_28677,N_29616);
or UO_879 (O_879,N_28211,N_29812);
or UO_880 (O_880,N_28418,N_28630);
nand UO_881 (O_881,N_29627,N_28600);
nand UO_882 (O_882,N_28613,N_29901);
and UO_883 (O_883,N_29702,N_28135);
or UO_884 (O_884,N_28314,N_28185);
xnor UO_885 (O_885,N_29524,N_28127);
nor UO_886 (O_886,N_28609,N_29808);
nor UO_887 (O_887,N_28227,N_29549);
nor UO_888 (O_888,N_29597,N_28592);
nand UO_889 (O_889,N_28563,N_29946);
and UO_890 (O_890,N_28152,N_29480);
xor UO_891 (O_891,N_29994,N_28798);
xnor UO_892 (O_892,N_29499,N_29552);
or UO_893 (O_893,N_29831,N_29436);
nand UO_894 (O_894,N_29317,N_29245);
or UO_895 (O_895,N_28452,N_29023);
nand UO_896 (O_896,N_28036,N_28555);
and UO_897 (O_897,N_29473,N_29492);
or UO_898 (O_898,N_29068,N_29939);
nand UO_899 (O_899,N_29559,N_28540);
and UO_900 (O_900,N_28182,N_29158);
xor UO_901 (O_901,N_29028,N_28472);
nor UO_902 (O_902,N_29121,N_28960);
nor UO_903 (O_903,N_28033,N_28289);
or UO_904 (O_904,N_28388,N_29256);
nor UO_905 (O_905,N_29463,N_28079);
nor UO_906 (O_906,N_29081,N_29990);
nor UO_907 (O_907,N_28854,N_29359);
xnor UO_908 (O_908,N_29230,N_28432);
and UO_909 (O_909,N_29411,N_29527);
nor UO_910 (O_910,N_29910,N_29297);
and UO_911 (O_911,N_29684,N_28374);
or UO_912 (O_912,N_28906,N_28140);
nand UO_913 (O_913,N_29008,N_28384);
nor UO_914 (O_914,N_29372,N_28974);
and UO_915 (O_915,N_28635,N_28681);
and UO_916 (O_916,N_28077,N_28064);
nand UO_917 (O_917,N_29206,N_29953);
or UO_918 (O_918,N_29130,N_28720);
or UO_919 (O_919,N_28070,N_29810);
nor UO_920 (O_920,N_28503,N_29694);
or UO_921 (O_921,N_29370,N_28664);
and UO_922 (O_922,N_28730,N_29818);
nor UO_923 (O_923,N_29649,N_29131);
or UO_924 (O_924,N_28963,N_28698);
or UO_925 (O_925,N_29168,N_29030);
or UO_926 (O_926,N_28778,N_29759);
nor UO_927 (O_927,N_29074,N_28693);
and UO_928 (O_928,N_29139,N_29344);
nand UO_929 (O_929,N_28293,N_29148);
nor UO_930 (O_930,N_28408,N_29233);
nor UO_931 (O_931,N_28023,N_28972);
or UO_932 (O_932,N_28138,N_28075);
or UO_933 (O_933,N_29386,N_29319);
nor UO_934 (O_934,N_29126,N_28710);
nand UO_935 (O_935,N_28553,N_28078);
nor UO_936 (O_936,N_29425,N_28061);
nor UO_937 (O_937,N_29556,N_29892);
xor UO_938 (O_938,N_28987,N_28088);
xnor UO_939 (O_939,N_29093,N_28604);
nor UO_940 (O_940,N_28957,N_29373);
and UO_941 (O_941,N_28091,N_29900);
and UO_942 (O_942,N_29305,N_29839);
and UO_943 (O_943,N_29355,N_28172);
nor UO_944 (O_944,N_28198,N_28614);
nor UO_945 (O_945,N_29078,N_28173);
nor UO_946 (O_946,N_29637,N_28758);
nor UO_947 (O_947,N_28455,N_28239);
nor UO_948 (O_948,N_29294,N_28049);
xnor UO_949 (O_949,N_29782,N_28813);
or UO_950 (O_950,N_28759,N_28000);
nand UO_951 (O_951,N_28300,N_29312);
nor UO_952 (O_952,N_28887,N_29916);
nand UO_953 (O_953,N_28576,N_29848);
xor UO_954 (O_954,N_28092,N_29538);
and UO_955 (O_955,N_29252,N_28226);
xor UO_956 (O_956,N_28667,N_28191);
xnor UO_957 (O_957,N_28954,N_29127);
nor UO_958 (O_958,N_29610,N_29352);
xor UO_959 (O_959,N_28082,N_29682);
xnor UO_960 (O_960,N_29257,N_29743);
nor UO_961 (O_961,N_28272,N_29719);
xnor UO_962 (O_962,N_29156,N_28261);
and UO_963 (O_963,N_29842,N_28034);
xor UO_964 (O_964,N_28164,N_29248);
nand UO_965 (O_965,N_28063,N_29238);
nor UO_966 (O_966,N_28304,N_29887);
xor UO_967 (O_967,N_28841,N_28260);
nand UO_968 (O_968,N_28438,N_29522);
xor UO_969 (O_969,N_28946,N_29056);
nand UO_970 (O_970,N_29585,N_28874);
or UO_971 (O_971,N_28480,N_28230);
xor UO_972 (O_972,N_28291,N_29643);
nand UO_973 (O_973,N_29914,N_29563);
nor UO_974 (O_974,N_28117,N_28812);
nand UO_975 (O_975,N_28102,N_28383);
and UO_976 (O_976,N_29985,N_28723);
and UO_977 (O_977,N_28688,N_29966);
or UO_978 (O_978,N_29381,N_29338);
and UO_979 (O_979,N_28931,N_28970);
or UO_980 (O_980,N_29331,N_28056);
nand UO_981 (O_981,N_28790,N_28378);
or UO_982 (O_982,N_29173,N_29398);
nor UO_983 (O_983,N_29587,N_29796);
nor UO_984 (O_984,N_28649,N_29360);
nand UO_985 (O_985,N_28179,N_29560);
nor UO_986 (O_986,N_29287,N_28476);
or UO_987 (O_987,N_28328,N_28004);
nor UO_988 (O_988,N_28660,N_29132);
and UO_989 (O_989,N_28965,N_28288);
xor UO_990 (O_990,N_29504,N_28050);
nand UO_991 (O_991,N_28549,N_29190);
and UO_992 (O_992,N_28420,N_28870);
nand UO_993 (O_993,N_29418,N_29401);
or UO_994 (O_994,N_28207,N_28766);
nor UO_995 (O_995,N_29015,N_28626);
and UO_996 (O_996,N_29935,N_28742);
and UO_997 (O_997,N_29080,N_29420);
or UO_998 (O_998,N_29301,N_28916);
nand UO_999 (O_999,N_29986,N_28154);
nand UO_1000 (O_1000,N_28411,N_29132);
and UO_1001 (O_1001,N_28258,N_28909);
and UO_1002 (O_1002,N_28153,N_28707);
nor UO_1003 (O_1003,N_28756,N_28673);
nand UO_1004 (O_1004,N_28611,N_28926);
or UO_1005 (O_1005,N_29929,N_28852);
and UO_1006 (O_1006,N_28180,N_28750);
nand UO_1007 (O_1007,N_29239,N_28716);
and UO_1008 (O_1008,N_29015,N_28261);
xor UO_1009 (O_1009,N_28124,N_29558);
xnor UO_1010 (O_1010,N_28220,N_29223);
xor UO_1011 (O_1011,N_29249,N_29420);
and UO_1012 (O_1012,N_28140,N_29030);
xor UO_1013 (O_1013,N_29616,N_28504);
nor UO_1014 (O_1014,N_28982,N_28694);
and UO_1015 (O_1015,N_29001,N_29364);
and UO_1016 (O_1016,N_29016,N_29957);
nand UO_1017 (O_1017,N_29562,N_28488);
or UO_1018 (O_1018,N_29682,N_29487);
nor UO_1019 (O_1019,N_29014,N_28915);
xor UO_1020 (O_1020,N_28870,N_29542);
or UO_1021 (O_1021,N_29411,N_28850);
nand UO_1022 (O_1022,N_28886,N_29181);
xor UO_1023 (O_1023,N_28598,N_28327);
nand UO_1024 (O_1024,N_28156,N_28516);
or UO_1025 (O_1025,N_29229,N_28268);
nand UO_1026 (O_1026,N_29037,N_29732);
nor UO_1027 (O_1027,N_29340,N_29679);
and UO_1028 (O_1028,N_29329,N_29756);
and UO_1029 (O_1029,N_29165,N_29961);
nor UO_1030 (O_1030,N_29643,N_28091);
nor UO_1031 (O_1031,N_29734,N_28725);
xnor UO_1032 (O_1032,N_28154,N_29740);
nand UO_1033 (O_1033,N_28828,N_28251);
nand UO_1034 (O_1034,N_29066,N_28181);
xor UO_1035 (O_1035,N_28190,N_29170);
nor UO_1036 (O_1036,N_28534,N_28196);
nor UO_1037 (O_1037,N_28999,N_29722);
or UO_1038 (O_1038,N_29284,N_29594);
or UO_1039 (O_1039,N_28451,N_28005);
nor UO_1040 (O_1040,N_29712,N_28647);
and UO_1041 (O_1041,N_29694,N_28454);
nor UO_1042 (O_1042,N_28855,N_28008);
and UO_1043 (O_1043,N_28599,N_29728);
xor UO_1044 (O_1044,N_29277,N_29700);
xnor UO_1045 (O_1045,N_29239,N_29949);
nand UO_1046 (O_1046,N_29888,N_29044);
xnor UO_1047 (O_1047,N_28517,N_29315);
nor UO_1048 (O_1048,N_28496,N_28203);
nor UO_1049 (O_1049,N_28463,N_29121);
or UO_1050 (O_1050,N_28479,N_29499);
or UO_1051 (O_1051,N_29440,N_28763);
nand UO_1052 (O_1052,N_28656,N_29485);
xnor UO_1053 (O_1053,N_28756,N_28215);
nand UO_1054 (O_1054,N_28805,N_28835);
and UO_1055 (O_1055,N_29781,N_29247);
or UO_1056 (O_1056,N_29034,N_28378);
nand UO_1057 (O_1057,N_29295,N_29929);
nand UO_1058 (O_1058,N_28374,N_28002);
and UO_1059 (O_1059,N_29139,N_28161);
xor UO_1060 (O_1060,N_29651,N_28443);
and UO_1061 (O_1061,N_29095,N_29737);
nor UO_1062 (O_1062,N_28225,N_29184);
nor UO_1063 (O_1063,N_28699,N_28799);
nor UO_1064 (O_1064,N_28501,N_29009);
or UO_1065 (O_1065,N_29252,N_29342);
or UO_1066 (O_1066,N_28396,N_29545);
nor UO_1067 (O_1067,N_28989,N_29418);
nor UO_1068 (O_1068,N_29285,N_29217);
or UO_1069 (O_1069,N_29445,N_28126);
and UO_1070 (O_1070,N_29439,N_29217);
nand UO_1071 (O_1071,N_29449,N_29217);
nand UO_1072 (O_1072,N_29073,N_28826);
and UO_1073 (O_1073,N_28147,N_29030);
and UO_1074 (O_1074,N_29149,N_28927);
and UO_1075 (O_1075,N_28966,N_29694);
nand UO_1076 (O_1076,N_29383,N_28513);
or UO_1077 (O_1077,N_28283,N_28422);
or UO_1078 (O_1078,N_28341,N_28685);
nor UO_1079 (O_1079,N_28703,N_29831);
or UO_1080 (O_1080,N_28330,N_28366);
or UO_1081 (O_1081,N_29168,N_29831);
nand UO_1082 (O_1082,N_29647,N_28747);
nand UO_1083 (O_1083,N_29901,N_29850);
nand UO_1084 (O_1084,N_29165,N_29135);
nand UO_1085 (O_1085,N_28470,N_29086);
xor UO_1086 (O_1086,N_29910,N_29524);
nand UO_1087 (O_1087,N_28260,N_29712);
nand UO_1088 (O_1088,N_28208,N_29160);
and UO_1089 (O_1089,N_29877,N_28186);
xnor UO_1090 (O_1090,N_28889,N_28261);
nand UO_1091 (O_1091,N_28748,N_28119);
nor UO_1092 (O_1092,N_28295,N_28758);
nor UO_1093 (O_1093,N_29624,N_29313);
nand UO_1094 (O_1094,N_28799,N_29568);
nor UO_1095 (O_1095,N_29135,N_28636);
nor UO_1096 (O_1096,N_28529,N_28734);
xnor UO_1097 (O_1097,N_29143,N_28110);
or UO_1098 (O_1098,N_29105,N_29925);
nand UO_1099 (O_1099,N_29097,N_28602);
and UO_1100 (O_1100,N_29529,N_28982);
nand UO_1101 (O_1101,N_29421,N_29774);
and UO_1102 (O_1102,N_28534,N_28287);
nor UO_1103 (O_1103,N_29540,N_29517);
nor UO_1104 (O_1104,N_29668,N_28138);
nand UO_1105 (O_1105,N_28175,N_29968);
nand UO_1106 (O_1106,N_29752,N_28388);
and UO_1107 (O_1107,N_29335,N_29504);
xor UO_1108 (O_1108,N_28280,N_29131);
xor UO_1109 (O_1109,N_29229,N_29224);
and UO_1110 (O_1110,N_28479,N_28185);
or UO_1111 (O_1111,N_28244,N_28081);
xor UO_1112 (O_1112,N_28603,N_28664);
xor UO_1113 (O_1113,N_29308,N_29964);
nor UO_1114 (O_1114,N_28227,N_29196);
and UO_1115 (O_1115,N_29465,N_28557);
nor UO_1116 (O_1116,N_28583,N_28508);
nor UO_1117 (O_1117,N_28361,N_28985);
xor UO_1118 (O_1118,N_28519,N_28976);
and UO_1119 (O_1119,N_28977,N_29816);
or UO_1120 (O_1120,N_29695,N_28471);
and UO_1121 (O_1121,N_28597,N_28841);
xor UO_1122 (O_1122,N_29679,N_28914);
xor UO_1123 (O_1123,N_29087,N_28368);
nand UO_1124 (O_1124,N_28874,N_28264);
nand UO_1125 (O_1125,N_28184,N_28535);
xor UO_1126 (O_1126,N_28491,N_28377);
xor UO_1127 (O_1127,N_29589,N_29302);
nand UO_1128 (O_1128,N_28467,N_28001);
nand UO_1129 (O_1129,N_28923,N_28460);
nor UO_1130 (O_1130,N_28460,N_29529);
nor UO_1131 (O_1131,N_28591,N_29201);
or UO_1132 (O_1132,N_29004,N_29036);
or UO_1133 (O_1133,N_29777,N_29241);
or UO_1134 (O_1134,N_28362,N_29352);
nor UO_1135 (O_1135,N_28794,N_29911);
and UO_1136 (O_1136,N_28479,N_29807);
nand UO_1137 (O_1137,N_28220,N_28741);
xnor UO_1138 (O_1138,N_28327,N_29847);
nor UO_1139 (O_1139,N_29947,N_29815);
nand UO_1140 (O_1140,N_29180,N_29913);
xnor UO_1141 (O_1141,N_28955,N_29982);
xnor UO_1142 (O_1142,N_28623,N_28603);
xnor UO_1143 (O_1143,N_29245,N_28123);
nand UO_1144 (O_1144,N_29176,N_29606);
nand UO_1145 (O_1145,N_28983,N_28966);
xor UO_1146 (O_1146,N_29419,N_28295);
or UO_1147 (O_1147,N_28365,N_28451);
nor UO_1148 (O_1148,N_29671,N_28275);
and UO_1149 (O_1149,N_28357,N_28412);
nor UO_1150 (O_1150,N_29884,N_29791);
and UO_1151 (O_1151,N_29557,N_29975);
xor UO_1152 (O_1152,N_28072,N_29909);
nor UO_1153 (O_1153,N_28817,N_29879);
nand UO_1154 (O_1154,N_29859,N_28186);
nand UO_1155 (O_1155,N_28409,N_29579);
nor UO_1156 (O_1156,N_29743,N_29721);
and UO_1157 (O_1157,N_29556,N_28097);
and UO_1158 (O_1158,N_29254,N_29661);
and UO_1159 (O_1159,N_29035,N_29277);
and UO_1160 (O_1160,N_28443,N_28308);
or UO_1161 (O_1161,N_28170,N_29889);
or UO_1162 (O_1162,N_29654,N_28821);
or UO_1163 (O_1163,N_28155,N_29995);
and UO_1164 (O_1164,N_29532,N_29407);
xnor UO_1165 (O_1165,N_28084,N_28844);
and UO_1166 (O_1166,N_28599,N_28376);
nand UO_1167 (O_1167,N_28503,N_29641);
nor UO_1168 (O_1168,N_28537,N_29459);
nor UO_1169 (O_1169,N_29086,N_29235);
nor UO_1170 (O_1170,N_29359,N_28119);
xnor UO_1171 (O_1171,N_28511,N_28880);
nand UO_1172 (O_1172,N_29692,N_29698);
nand UO_1173 (O_1173,N_29345,N_29653);
or UO_1174 (O_1174,N_29837,N_28098);
or UO_1175 (O_1175,N_28287,N_28676);
xor UO_1176 (O_1176,N_28656,N_28124);
nor UO_1177 (O_1177,N_29625,N_29540);
and UO_1178 (O_1178,N_29563,N_28856);
xnor UO_1179 (O_1179,N_28489,N_29884);
and UO_1180 (O_1180,N_28194,N_29609);
xnor UO_1181 (O_1181,N_29518,N_29917);
nand UO_1182 (O_1182,N_29149,N_29969);
xor UO_1183 (O_1183,N_28253,N_28872);
or UO_1184 (O_1184,N_28527,N_29917);
and UO_1185 (O_1185,N_29583,N_28067);
xor UO_1186 (O_1186,N_28408,N_29696);
nor UO_1187 (O_1187,N_28057,N_29132);
nand UO_1188 (O_1188,N_28235,N_29717);
xnor UO_1189 (O_1189,N_29290,N_29484);
nand UO_1190 (O_1190,N_29309,N_29091);
nor UO_1191 (O_1191,N_29809,N_28797);
nor UO_1192 (O_1192,N_28636,N_28629);
xnor UO_1193 (O_1193,N_28384,N_28039);
nor UO_1194 (O_1194,N_29785,N_29130);
or UO_1195 (O_1195,N_28097,N_28924);
nand UO_1196 (O_1196,N_28927,N_29579);
nand UO_1197 (O_1197,N_28971,N_28561);
and UO_1198 (O_1198,N_28251,N_29429);
nor UO_1199 (O_1199,N_28016,N_29577);
nand UO_1200 (O_1200,N_29158,N_28673);
nor UO_1201 (O_1201,N_28111,N_28923);
or UO_1202 (O_1202,N_28686,N_28670);
nor UO_1203 (O_1203,N_28733,N_29466);
nor UO_1204 (O_1204,N_29126,N_29235);
xnor UO_1205 (O_1205,N_29660,N_29373);
or UO_1206 (O_1206,N_28547,N_29950);
and UO_1207 (O_1207,N_29177,N_28829);
nand UO_1208 (O_1208,N_29905,N_28259);
nand UO_1209 (O_1209,N_28994,N_29458);
xor UO_1210 (O_1210,N_29955,N_28457);
nor UO_1211 (O_1211,N_28179,N_29438);
xnor UO_1212 (O_1212,N_28003,N_29053);
nor UO_1213 (O_1213,N_28702,N_29062);
xor UO_1214 (O_1214,N_28789,N_28662);
nand UO_1215 (O_1215,N_29609,N_28842);
or UO_1216 (O_1216,N_28082,N_29697);
and UO_1217 (O_1217,N_28720,N_28456);
nor UO_1218 (O_1218,N_28017,N_28572);
or UO_1219 (O_1219,N_28136,N_28745);
or UO_1220 (O_1220,N_28567,N_29044);
or UO_1221 (O_1221,N_28795,N_29532);
xor UO_1222 (O_1222,N_29866,N_28874);
and UO_1223 (O_1223,N_28797,N_29787);
nor UO_1224 (O_1224,N_28698,N_28854);
nand UO_1225 (O_1225,N_28615,N_29476);
and UO_1226 (O_1226,N_29843,N_28414);
and UO_1227 (O_1227,N_29182,N_29116);
xor UO_1228 (O_1228,N_29646,N_29898);
xnor UO_1229 (O_1229,N_28331,N_28475);
or UO_1230 (O_1230,N_28888,N_29800);
nor UO_1231 (O_1231,N_29713,N_28154);
nand UO_1232 (O_1232,N_28667,N_28571);
and UO_1233 (O_1233,N_28925,N_28600);
and UO_1234 (O_1234,N_28373,N_28840);
xnor UO_1235 (O_1235,N_28717,N_29121);
and UO_1236 (O_1236,N_29522,N_28297);
nor UO_1237 (O_1237,N_28017,N_29632);
nor UO_1238 (O_1238,N_29383,N_29272);
and UO_1239 (O_1239,N_28768,N_29639);
and UO_1240 (O_1240,N_29854,N_28824);
nor UO_1241 (O_1241,N_29491,N_28437);
nand UO_1242 (O_1242,N_28005,N_29052);
xnor UO_1243 (O_1243,N_29627,N_29514);
and UO_1244 (O_1244,N_28617,N_29602);
nand UO_1245 (O_1245,N_28134,N_29424);
and UO_1246 (O_1246,N_29112,N_29545);
and UO_1247 (O_1247,N_28527,N_29441);
and UO_1248 (O_1248,N_29648,N_28250);
and UO_1249 (O_1249,N_29345,N_29724);
xnor UO_1250 (O_1250,N_28923,N_28043);
xnor UO_1251 (O_1251,N_29945,N_28575);
and UO_1252 (O_1252,N_28310,N_29203);
or UO_1253 (O_1253,N_29342,N_28216);
nor UO_1254 (O_1254,N_28998,N_28074);
or UO_1255 (O_1255,N_29696,N_28597);
nor UO_1256 (O_1256,N_29718,N_28458);
or UO_1257 (O_1257,N_29472,N_29108);
or UO_1258 (O_1258,N_29570,N_29497);
nand UO_1259 (O_1259,N_29800,N_28682);
nand UO_1260 (O_1260,N_28174,N_28106);
nor UO_1261 (O_1261,N_28081,N_29956);
xnor UO_1262 (O_1262,N_29232,N_29124);
xnor UO_1263 (O_1263,N_28447,N_28958);
nor UO_1264 (O_1264,N_29146,N_28496);
and UO_1265 (O_1265,N_29866,N_29585);
and UO_1266 (O_1266,N_28307,N_29949);
xnor UO_1267 (O_1267,N_28840,N_29000);
or UO_1268 (O_1268,N_29323,N_28835);
and UO_1269 (O_1269,N_28190,N_29721);
or UO_1270 (O_1270,N_28398,N_28527);
nand UO_1271 (O_1271,N_29260,N_29945);
nor UO_1272 (O_1272,N_29517,N_28054);
or UO_1273 (O_1273,N_28154,N_29978);
xnor UO_1274 (O_1274,N_29797,N_29111);
nand UO_1275 (O_1275,N_29371,N_29482);
or UO_1276 (O_1276,N_28184,N_29679);
nor UO_1277 (O_1277,N_29238,N_28856);
nand UO_1278 (O_1278,N_29031,N_29874);
and UO_1279 (O_1279,N_28270,N_29298);
nor UO_1280 (O_1280,N_29583,N_29019);
or UO_1281 (O_1281,N_29829,N_29448);
xor UO_1282 (O_1282,N_28898,N_28290);
nor UO_1283 (O_1283,N_29073,N_29807);
or UO_1284 (O_1284,N_28758,N_29030);
nand UO_1285 (O_1285,N_28050,N_29829);
nor UO_1286 (O_1286,N_28752,N_28238);
nor UO_1287 (O_1287,N_29026,N_29312);
nor UO_1288 (O_1288,N_29847,N_29505);
nand UO_1289 (O_1289,N_28568,N_29095);
or UO_1290 (O_1290,N_29348,N_28567);
and UO_1291 (O_1291,N_28390,N_29292);
xor UO_1292 (O_1292,N_28189,N_29588);
nand UO_1293 (O_1293,N_29867,N_29286);
or UO_1294 (O_1294,N_28609,N_28279);
nand UO_1295 (O_1295,N_29156,N_28881);
or UO_1296 (O_1296,N_28269,N_28322);
nor UO_1297 (O_1297,N_29341,N_29227);
nor UO_1298 (O_1298,N_29888,N_29164);
nand UO_1299 (O_1299,N_29392,N_29197);
xor UO_1300 (O_1300,N_28060,N_29296);
nor UO_1301 (O_1301,N_28145,N_28854);
xnor UO_1302 (O_1302,N_28465,N_29050);
xnor UO_1303 (O_1303,N_29663,N_29349);
or UO_1304 (O_1304,N_29892,N_29430);
xnor UO_1305 (O_1305,N_28785,N_29131);
nand UO_1306 (O_1306,N_29301,N_29614);
or UO_1307 (O_1307,N_29465,N_28654);
and UO_1308 (O_1308,N_29983,N_29267);
nor UO_1309 (O_1309,N_29481,N_29019);
and UO_1310 (O_1310,N_29874,N_29202);
xnor UO_1311 (O_1311,N_29826,N_28161);
or UO_1312 (O_1312,N_28985,N_28867);
nand UO_1313 (O_1313,N_29251,N_28182);
nand UO_1314 (O_1314,N_29877,N_28140);
and UO_1315 (O_1315,N_29167,N_29738);
xnor UO_1316 (O_1316,N_28792,N_28442);
nand UO_1317 (O_1317,N_29239,N_28484);
nor UO_1318 (O_1318,N_28670,N_28171);
xnor UO_1319 (O_1319,N_28808,N_29101);
or UO_1320 (O_1320,N_28009,N_29204);
xnor UO_1321 (O_1321,N_29332,N_28221);
or UO_1322 (O_1322,N_29575,N_29974);
or UO_1323 (O_1323,N_28730,N_29752);
xnor UO_1324 (O_1324,N_29152,N_29110);
nand UO_1325 (O_1325,N_29506,N_29670);
nand UO_1326 (O_1326,N_28062,N_28533);
nor UO_1327 (O_1327,N_28110,N_28675);
xnor UO_1328 (O_1328,N_28133,N_28281);
xor UO_1329 (O_1329,N_28072,N_29593);
and UO_1330 (O_1330,N_28798,N_28965);
xnor UO_1331 (O_1331,N_28493,N_28990);
and UO_1332 (O_1332,N_28673,N_28024);
and UO_1333 (O_1333,N_28886,N_29709);
nor UO_1334 (O_1334,N_29270,N_28416);
nand UO_1335 (O_1335,N_29950,N_28117);
nand UO_1336 (O_1336,N_28691,N_29678);
nand UO_1337 (O_1337,N_29876,N_29544);
nand UO_1338 (O_1338,N_29330,N_28090);
and UO_1339 (O_1339,N_29141,N_29058);
xnor UO_1340 (O_1340,N_29400,N_28507);
nor UO_1341 (O_1341,N_29081,N_29699);
or UO_1342 (O_1342,N_28194,N_28078);
and UO_1343 (O_1343,N_29577,N_28075);
nand UO_1344 (O_1344,N_29363,N_28745);
or UO_1345 (O_1345,N_29844,N_28696);
and UO_1346 (O_1346,N_28800,N_29505);
nand UO_1347 (O_1347,N_29539,N_28977);
and UO_1348 (O_1348,N_28248,N_29957);
and UO_1349 (O_1349,N_29618,N_28616);
or UO_1350 (O_1350,N_28460,N_28219);
nand UO_1351 (O_1351,N_28835,N_29922);
xnor UO_1352 (O_1352,N_29643,N_29426);
nor UO_1353 (O_1353,N_29476,N_28155);
xnor UO_1354 (O_1354,N_28496,N_28813);
nor UO_1355 (O_1355,N_29906,N_28934);
and UO_1356 (O_1356,N_29608,N_29174);
and UO_1357 (O_1357,N_28327,N_28528);
nor UO_1358 (O_1358,N_29475,N_28845);
or UO_1359 (O_1359,N_29547,N_29342);
or UO_1360 (O_1360,N_28007,N_29130);
nor UO_1361 (O_1361,N_29963,N_29029);
and UO_1362 (O_1362,N_28401,N_29666);
xnor UO_1363 (O_1363,N_29396,N_28531);
xor UO_1364 (O_1364,N_29876,N_29743);
nor UO_1365 (O_1365,N_29112,N_29268);
xor UO_1366 (O_1366,N_28962,N_29121);
and UO_1367 (O_1367,N_28336,N_28664);
and UO_1368 (O_1368,N_29150,N_28118);
nand UO_1369 (O_1369,N_29579,N_29174);
nand UO_1370 (O_1370,N_29953,N_29536);
or UO_1371 (O_1371,N_28348,N_28629);
or UO_1372 (O_1372,N_29237,N_29263);
xnor UO_1373 (O_1373,N_29300,N_29521);
nor UO_1374 (O_1374,N_28610,N_28136);
nand UO_1375 (O_1375,N_29083,N_29918);
nor UO_1376 (O_1376,N_29390,N_29027);
nor UO_1377 (O_1377,N_29587,N_29963);
nand UO_1378 (O_1378,N_29514,N_29008);
or UO_1379 (O_1379,N_28879,N_29393);
nor UO_1380 (O_1380,N_28929,N_28370);
nor UO_1381 (O_1381,N_28546,N_29559);
and UO_1382 (O_1382,N_28339,N_29935);
xor UO_1383 (O_1383,N_29044,N_28696);
nor UO_1384 (O_1384,N_29201,N_29877);
nand UO_1385 (O_1385,N_29535,N_29473);
xor UO_1386 (O_1386,N_28894,N_28523);
nor UO_1387 (O_1387,N_29288,N_29353);
or UO_1388 (O_1388,N_29331,N_28277);
nand UO_1389 (O_1389,N_29898,N_29258);
nor UO_1390 (O_1390,N_29626,N_29122);
xor UO_1391 (O_1391,N_28321,N_29763);
nand UO_1392 (O_1392,N_28514,N_29578);
and UO_1393 (O_1393,N_29720,N_28299);
and UO_1394 (O_1394,N_29931,N_29192);
xor UO_1395 (O_1395,N_28927,N_29691);
nor UO_1396 (O_1396,N_29272,N_29131);
nand UO_1397 (O_1397,N_28138,N_28633);
and UO_1398 (O_1398,N_28106,N_29506);
xor UO_1399 (O_1399,N_28019,N_29950);
or UO_1400 (O_1400,N_29984,N_28687);
or UO_1401 (O_1401,N_28265,N_29986);
nor UO_1402 (O_1402,N_28736,N_28666);
and UO_1403 (O_1403,N_28183,N_29184);
nor UO_1404 (O_1404,N_28437,N_29058);
or UO_1405 (O_1405,N_29683,N_28098);
nor UO_1406 (O_1406,N_29900,N_28677);
nor UO_1407 (O_1407,N_28772,N_28714);
nor UO_1408 (O_1408,N_29978,N_28018);
or UO_1409 (O_1409,N_29135,N_29554);
nand UO_1410 (O_1410,N_28959,N_28305);
xor UO_1411 (O_1411,N_29758,N_29943);
nor UO_1412 (O_1412,N_29145,N_28941);
xor UO_1413 (O_1413,N_28642,N_29542);
nand UO_1414 (O_1414,N_28348,N_28604);
nand UO_1415 (O_1415,N_29010,N_29327);
nand UO_1416 (O_1416,N_29425,N_28966);
and UO_1417 (O_1417,N_28278,N_28417);
or UO_1418 (O_1418,N_29627,N_29274);
xor UO_1419 (O_1419,N_28330,N_28803);
xnor UO_1420 (O_1420,N_29425,N_29990);
nand UO_1421 (O_1421,N_29651,N_29660);
nand UO_1422 (O_1422,N_29209,N_28204);
xor UO_1423 (O_1423,N_29060,N_28779);
and UO_1424 (O_1424,N_28534,N_28197);
nor UO_1425 (O_1425,N_29176,N_29211);
nor UO_1426 (O_1426,N_28724,N_29532);
xnor UO_1427 (O_1427,N_29084,N_29569);
xnor UO_1428 (O_1428,N_29627,N_29626);
or UO_1429 (O_1429,N_29318,N_28820);
nand UO_1430 (O_1430,N_29734,N_29049);
and UO_1431 (O_1431,N_28357,N_29773);
nand UO_1432 (O_1432,N_28159,N_28401);
or UO_1433 (O_1433,N_29277,N_28926);
nand UO_1434 (O_1434,N_29675,N_28808);
xor UO_1435 (O_1435,N_29437,N_28774);
xnor UO_1436 (O_1436,N_29900,N_28656);
nor UO_1437 (O_1437,N_28932,N_29727);
xor UO_1438 (O_1438,N_28729,N_29860);
xor UO_1439 (O_1439,N_29932,N_29622);
or UO_1440 (O_1440,N_29100,N_29123);
and UO_1441 (O_1441,N_29845,N_28055);
or UO_1442 (O_1442,N_28161,N_29472);
nand UO_1443 (O_1443,N_28792,N_28369);
nand UO_1444 (O_1444,N_29501,N_28353);
nor UO_1445 (O_1445,N_29233,N_28801);
nor UO_1446 (O_1446,N_28119,N_28921);
nand UO_1447 (O_1447,N_28554,N_28919);
and UO_1448 (O_1448,N_28065,N_28596);
nand UO_1449 (O_1449,N_29109,N_29696);
and UO_1450 (O_1450,N_28069,N_28827);
nor UO_1451 (O_1451,N_29903,N_29451);
nand UO_1452 (O_1452,N_28683,N_28030);
or UO_1453 (O_1453,N_29758,N_28492);
xor UO_1454 (O_1454,N_28265,N_28051);
xnor UO_1455 (O_1455,N_29636,N_29577);
xor UO_1456 (O_1456,N_29624,N_28021);
nor UO_1457 (O_1457,N_28525,N_29176);
and UO_1458 (O_1458,N_28930,N_28511);
xnor UO_1459 (O_1459,N_28869,N_29312);
nor UO_1460 (O_1460,N_29229,N_29418);
xor UO_1461 (O_1461,N_29702,N_29939);
or UO_1462 (O_1462,N_28100,N_29624);
nor UO_1463 (O_1463,N_28880,N_28307);
nor UO_1464 (O_1464,N_29450,N_28722);
nor UO_1465 (O_1465,N_29504,N_28931);
and UO_1466 (O_1466,N_29612,N_28417);
xor UO_1467 (O_1467,N_29071,N_28256);
and UO_1468 (O_1468,N_28933,N_29599);
nor UO_1469 (O_1469,N_29228,N_28811);
or UO_1470 (O_1470,N_28278,N_29752);
nand UO_1471 (O_1471,N_28937,N_29618);
nand UO_1472 (O_1472,N_29557,N_28718);
xor UO_1473 (O_1473,N_29937,N_29769);
and UO_1474 (O_1474,N_28816,N_29857);
nand UO_1475 (O_1475,N_29221,N_28164);
nand UO_1476 (O_1476,N_29996,N_29816);
nor UO_1477 (O_1477,N_28209,N_28010);
and UO_1478 (O_1478,N_28602,N_28179);
nand UO_1479 (O_1479,N_29299,N_28914);
xnor UO_1480 (O_1480,N_29524,N_28797);
or UO_1481 (O_1481,N_29134,N_28521);
and UO_1482 (O_1482,N_29747,N_28832);
and UO_1483 (O_1483,N_28757,N_28467);
nor UO_1484 (O_1484,N_29904,N_29679);
nand UO_1485 (O_1485,N_28781,N_29126);
or UO_1486 (O_1486,N_29888,N_28394);
and UO_1487 (O_1487,N_29904,N_29165);
nand UO_1488 (O_1488,N_29286,N_28814);
nand UO_1489 (O_1489,N_28266,N_28884);
and UO_1490 (O_1490,N_29542,N_28603);
and UO_1491 (O_1491,N_29871,N_28888);
xnor UO_1492 (O_1492,N_28200,N_28410);
and UO_1493 (O_1493,N_28385,N_28356);
or UO_1494 (O_1494,N_28459,N_29745);
and UO_1495 (O_1495,N_29048,N_29783);
xnor UO_1496 (O_1496,N_29179,N_29983);
and UO_1497 (O_1497,N_28491,N_29878);
nand UO_1498 (O_1498,N_28928,N_29659);
nor UO_1499 (O_1499,N_29225,N_28400);
and UO_1500 (O_1500,N_28380,N_29933);
nand UO_1501 (O_1501,N_29280,N_28834);
xnor UO_1502 (O_1502,N_28673,N_28951);
nor UO_1503 (O_1503,N_28729,N_29548);
and UO_1504 (O_1504,N_29837,N_28073);
and UO_1505 (O_1505,N_28936,N_29683);
or UO_1506 (O_1506,N_29334,N_29896);
nor UO_1507 (O_1507,N_29784,N_28277);
and UO_1508 (O_1508,N_29762,N_29854);
xor UO_1509 (O_1509,N_28581,N_29753);
and UO_1510 (O_1510,N_29941,N_28014);
nor UO_1511 (O_1511,N_29517,N_28829);
or UO_1512 (O_1512,N_29890,N_29029);
xor UO_1513 (O_1513,N_28257,N_29208);
nor UO_1514 (O_1514,N_29753,N_29519);
and UO_1515 (O_1515,N_28946,N_29617);
nor UO_1516 (O_1516,N_29890,N_28483);
nand UO_1517 (O_1517,N_29702,N_28105);
nor UO_1518 (O_1518,N_29117,N_29411);
nor UO_1519 (O_1519,N_28316,N_29297);
and UO_1520 (O_1520,N_29659,N_29861);
xnor UO_1521 (O_1521,N_28523,N_28638);
xnor UO_1522 (O_1522,N_29320,N_28730);
xnor UO_1523 (O_1523,N_28642,N_28605);
and UO_1524 (O_1524,N_28172,N_28610);
or UO_1525 (O_1525,N_29434,N_29341);
xnor UO_1526 (O_1526,N_28900,N_28357);
and UO_1527 (O_1527,N_29554,N_28649);
nor UO_1528 (O_1528,N_29811,N_29999);
and UO_1529 (O_1529,N_28386,N_29279);
nand UO_1530 (O_1530,N_29957,N_29401);
or UO_1531 (O_1531,N_29489,N_28064);
nand UO_1532 (O_1532,N_29423,N_29675);
xor UO_1533 (O_1533,N_29809,N_28366);
or UO_1534 (O_1534,N_29251,N_29293);
and UO_1535 (O_1535,N_28995,N_29935);
or UO_1536 (O_1536,N_28726,N_28532);
nor UO_1537 (O_1537,N_28224,N_29147);
xor UO_1538 (O_1538,N_28344,N_29832);
nor UO_1539 (O_1539,N_29879,N_28802);
nor UO_1540 (O_1540,N_28632,N_29850);
nand UO_1541 (O_1541,N_29220,N_29067);
or UO_1542 (O_1542,N_28562,N_29634);
xnor UO_1543 (O_1543,N_28239,N_29751);
or UO_1544 (O_1544,N_28628,N_29437);
nor UO_1545 (O_1545,N_28902,N_28737);
nor UO_1546 (O_1546,N_29788,N_29054);
and UO_1547 (O_1547,N_28588,N_29336);
nand UO_1548 (O_1548,N_28110,N_28547);
or UO_1549 (O_1549,N_28595,N_28107);
and UO_1550 (O_1550,N_28140,N_29356);
nand UO_1551 (O_1551,N_28787,N_28803);
or UO_1552 (O_1552,N_28433,N_28413);
nand UO_1553 (O_1553,N_28862,N_29787);
or UO_1554 (O_1554,N_28840,N_28267);
or UO_1555 (O_1555,N_29861,N_28967);
nor UO_1556 (O_1556,N_29705,N_28169);
nand UO_1557 (O_1557,N_28413,N_29134);
or UO_1558 (O_1558,N_29656,N_29456);
xnor UO_1559 (O_1559,N_29178,N_28155);
and UO_1560 (O_1560,N_29414,N_29182);
or UO_1561 (O_1561,N_29883,N_28237);
nor UO_1562 (O_1562,N_29748,N_28583);
or UO_1563 (O_1563,N_28702,N_29007);
nand UO_1564 (O_1564,N_28271,N_29328);
nand UO_1565 (O_1565,N_29405,N_29211);
nor UO_1566 (O_1566,N_29989,N_28609);
xnor UO_1567 (O_1567,N_29476,N_29830);
nand UO_1568 (O_1568,N_28462,N_28050);
xnor UO_1569 (O_1569,N_29628,N_29577);
and UO_1570 (O_1570,N_28479,N_28903);
or UO_1571 (O_1571,N_28505,N_29684);
and UO_1572 (O_1572,N_28936,N_28973);
nor UO_1573 (O_1573,N_29320,N_28673);
or UO_1574 (O_1574,N_29476,N_28629);
nand UO_1575 (O_1575,N_29727,N_29892);
xnor UO_1576 (O_1576,N_29076,N_28670);
nor UO_1577 (O_1577,N_29346,N_28152);
xor UO_1578 (O_1578,N_29477,N_29642);
nand UO_1579 (O_1579,N_28792,N_28847);
nor UO_1580 (O_1580,N_29538,N_29063);
and UO_1581 (O_1581,N_28543,N_29007);
xor UO_1582 (O_1582,N_29132,N_29559);
and UO_1583 (O_1583,N_28878,N_29609);
or UO_1584 (O_1584,N_29319,N_28564);
or UO_1585 (O_1585,N_29592,N_29058);
nor UO_1586 (O_1586,N_29030,N_29270);
and UO_1587 (O_1587,N_28339,N_28943);
nand UO_1588 (O_1588,N_28917,N_29172);
nor UO_1589 (O_1589,N_28778,N_28753);
and UO_1590 (O_1590,N_28781,N_29514);
xor UO_1591 (O_1591,N_29751,N_28191);
and UO_1592 (O_1592,N_29437,N_28341);
and UO_1593 (O_1593,N_29386,N_28495);
nand UO_1594 (O_1594,N_29566,N_29896);
and UO_1595 (O_1595,N_28999,N_29466);
nor UO_1596 (O_1596,N_29045,N_28464);
and UO_1597 (O_1597,N_29964,N_29903);
or UO_1598 (O_1598,N_28536,N_29440);
nor UO_1599 (O_1599,N_28178,N_29713);
and UO_1600 (O_1600,N_28156,N_29555);
or UO_1601 (O_1601,N_28278,N_29270);
nor UO_1602 (O_1602,N_28762,N_29521);
nand UO_1603 (O_1603,N_29406,N_29436);
and UO_1604 (O_1604,N_28090,N_29412);
and UO_1605 (O_1605,N_29847,N_28113);
xor UO_1606 (O_1606,N_28795,N_28397);
nand UO_1607 (O_1607,N_29208,N_29280);
or UO_1608 (O_1608,N_29568,N_28557);
or UO_1609 (O_1609,N_29518,N_28435);
or UO_1610 (O_1610,N_29251,N_29060);
nand UO_1611 (O_1611,N_29856,N_29771);
nor UO_1612 (O_1612,N_28721,N_29326);
xnor UO_1613 (O_1613,N_28419,N_29063);
nor UO_1614 (O_1614,N_28629,N_29857);
or UO_1615 (O_1615,N_28190,N_29292);
xnor UO_1616 (O_1616,N_28190,N_28790);
and UO_1617 (O_1617,N_28671,N_28407);
or UO_1618 (O_1618,N_29969,N_28373);
xnor UO_1619 (O_1619,N_29942,N_29458);
or UO_1620 (O_1620,N_29764,N_28769);
or UO_1621 (O_1621,N_28171,N_28277);
and UO_1622 (O_1622,N_29640,N_28298);
xnor UO_1623 (O_1623,N_29627,N_29867);
xor UO_1624 (O_1624,N_29171,N_28149);
nand UO_1625 (O_1625,N_29874,N_29045);
xor UO_1626 (O_1626,N_28819,N_29200);
nor UO_1627 (O_1627,N_28668,N_29384);
xnor UO_1628 (O_1628,N_28392,N_28162);
nand UO_1629 (O_1629,N_29892,N_28657);
nor UO_1630 (O_1630,N_29345,N_29242);
and UO_1631 (O_1631,N_29748,N_29541);
nand UO_1632 (O_1632,N_28007,N_29118);
and UO_1633 (O_1633,N_28405,N_28304);
xor UO_1634 (O_1634,N_28998,N_29868);
and UO_1635 (O_1635,N_28090,N_29037);
xor UO_1636 (O_1636,N_29348,N_29056);
xor UO_1637 (O_1637,N_28572,N_29038);
xor UO_1638 (O_1638,N_29985,N_29177);
xor UO_1639 (O_1639,N_29385,N_28794);
nand UO_1640 (O_1640,N_28682,N_28196);
nor UO_1641 (O_1641,N_29717,N_28261);
nor UO_1642 (O_1642,N_28827,N_29119);
nor UO_1643 (O_1643,N_29902,N_28853);
nand UO_1644 (O_1644,N_29233,N_28094);
or UO_1645 (O_1645,N_28531,N_28716);
and UO_1646 (O_1646,N_28969,N_29166);
xor UO_1647 (O_1647,N_28405,N_29043);
nand UO_1648 (O_1648,N_29863,N_28583);
or UO_1649 (O_1649,N_28780,N_28326);
nand UO_1650 (O_1650,N_29557,N_29785);
or UO_1651 (O_1651,N_28240,N_29570);
xnor UO_1652 (O_1652,N_29574,N_29041);
or UO_1653 (O_1653,N_29850,N_29515);
nand UO_1654 (O_1654,N_29512,N_28048);
xnor UO_1655 (O_1655,N_29533,N_29717);
xor UO_1656 (O_1656,N_29206,N_28699);
or UO_1657 (O_1657,N_28577,N_29965);
xnor UO_1658 (O_1658,N_29541,N_28876);
xor UO_1659 (O_1659,N_28551,N_29124);
or UO_1660 (O_1660,N_28985,N_29518);
nor UO_1661 (O_1661,N_29325,N_29403);
and UO_1662 (O_1662,N_29039,N_28619);
or UO_1663 (O_1663,N_28131,N_29991);
nand UO_1664 (O_1664,N_29443,N_29966);
nand UO_1665 (O_1665,N_29530,N_29827);
nand UO_1666 (O_1666,N_28733,N_28295);
nand UO_1667 (O_1667,N_28215,N_29834);
xnor UO_1668 (O_1668,N_28219,N_28558);
nor UO_1669 (O_1669,N_28006,N_29824);
nand UO_1670 (O_1670,N_28157,N_29297);
nand UO_1671 (O_1671,N_29929,N_28765);
nand UO_1672 (O_1672,N_28610,N_29321);
xor UO_1673 (O_1673,N_29488,N_29139);
nor UO_1674 (O_1674,N_28893,N_28390);
nor UO_1675 (O_1675,N_29028,N_28782);
nor UO_1676 (O_1676,N_28896,N_28082);
xor UO_1677 (O_1677,N_28843,N_28935);
or UO_1678 (O_1678,N_28348,N_28217);
or UO_1679 (O_1679,N_29600,N_29374);
and UO_1680 (O_1680,N_29788,N_29743);
nor UO_1681 (O_1681,N_28847,N_29403);
xnor UO_1682 (O_1682,N_28058,N_29217);
nand UO_1683 (O_1683,N_29943,N_29158);
or UO_1684 (O_1684,N_29508,N_28267);
or UO_1685 (O_1685,N_28684,N_29519);
or UO_1686 (O_1686,N_29151,N_29021);
and UO_1687 (O_1687,N_29750,N_28083);
nor UO_1688 (O_1688,N_28928,N_28575);
or UO_1689 (O_1689,N_28595,N_28532);
and UO_1690 (O_1690,N_29963,N_29740);
and UO_1691 (O_1691,N_29656,N_28904);
nor UO_1692 (O_1692,N_28209,N_29869);
and UO_1693 (O_1693,N_29952,N_28416);
or UO_1694 (O_1694,N_29930,N_29279);
nand UO_1695 (O_1695,N_28678,N_29020);
nand UO_1696 (O_1696,N_29085,N_29637);
nand UO_1697 (O_1697,N_28164,N_29027);
or UO_1698 (O_1698,N_28051,N_29957);
or UO_1699 (O_1699,N_28910,N_29120);
nor UO_1700 (O_1700,N_29965,N_29137);
xnor UO_1701 (O_1701,N_28528,N_29898);
nor UO_1702 (O_1702,N_29405,N_28337);
nor UO_1703 (O_1703,N_28755,N_28450);
nand UO_1704 (O_1704,N_28645,N_29543);
xnor UO_1705 (O_1705,N_28305,N_29055);
nor UO_1706 (O_1706,N_28399,N_28799);
nand UO_1707 (O_1707,N_29420,N_29773);
or UO_1708 (O_1708,N_28200,N_28168);
and UO_1709 (O_1709,N_29077,N_29851);
or UO_1710 (O_1710,N_28649,N_29164);
xor UO_1711 (O_1711,N_28823,N_28769);
and UO_1712 (O_1712,N_29658,N_28456);
nor UO_1713 (O_1713,N_29102,N_28880);
and UO_1714 (O_1714,N_28605,N_28533);
xor UO_1715 (O_1715,N_29157,N_29394);
xnor UO_1716 (O_1716,N_28053,N_28490);
and UO_1717 (O_1717,N_28805,N_28968);
nand UO_1718 (O_1718,N_28020,N_28739);
and UO_1719 (O_1719,N_28597,N_29459);
nand UO_1720 (O_1720,N_29882,N_29118);
nor UO_1721 (O_1721,N_28181,N_29944);
or UO_1722 (O_1722,N_29313,N_29699);
nor UO_1723 (O_1723,N_28732,N_29199);
or UO_1724 (O_1724,N_28183,N_29523);
xor UO_1725 (O_1725,N_29759,N_28393);
and UO_1726 (O_1726,N_29581,N_29966);
nand UO_1727 (O_1727,N_28848,N_28580);
xor UO_1728 (O_1728,N_28257,N_28318);
or UO_1729 (O_1729,N_29630,N_28331);
and UO_1730 (O_1730,N_29664,N_29997);
nor UO_1731 (O_1731,N_29514,N_28449);
and UO_1732 (O_1732,N_29335,N_28869);
nand UO_1733 (O_1733,N_28207,N_29123);
nand UO_1734 (O_1734,N_28468,N_28206);
xnor UO_1735 (O_1735,N_28373,N_28275);
and UO_1736 (O_1736,N_28812,N_29321);
and UO_1737 (O_1737,N_28155,N_29015);
nor UO_1738 (O_1738,N_28623,N_28507);
xnor UO_1739 (O_1739,N_28696,N_29628);
and UO_1740 (O_1740,N_29924,N_29814);
and UO_1741 (O_1741,N_29754,N_28709);
nand UO_1742 (O_1742,N_28220,N_28215);
and UO_1743 (O_1743,N_29795,N_29440);
or UO_1744 (O_1744,N_28104,N_29404);
nor UO_1745 (O_1745,N_29385,N_28429);
nand UO_1746 (O_1746,N_28024,N_29566);
or UO_1747 (O_1747,N_29496,N_28327);
or UO_1748 (O_1748,N_29340,N_29444);
xnor UO_1749 (O_1749,N_28043,N_29840);
or UO_1750 (O_1750,N_28360,N_28978);
or UO_1751 (O_1751,N_29459,N_29981);
nor UO_1752 (O_1752,N_28525,N_29472);
nor UO_1753 (O_1753,N_28863,N_28105);
or UO_1754 (O_1754,N_28811,N_28930);
nand UO_1755 (O_1755,N_29060,N_28864);
or UO_1756 (O_1756,N_28365,N_29228);
and UO_1757 (O_1757,N_29215,N_29633);
nor UO_1758 (O_1758,N_29613,N_29019);
nand UO_1759 (O_1759,N_29258,N_28940);
or UO_1760 (O_1760,N_29450,N_28676);
and UO_1761 (O_1761,N_29828,N_29010);
or UO_1762 (O_1762,N_29129,N_29133);
and UO_1763 (O_1763,N_29690,N_28017);
xnor UO_1764 (O_1764,N_28764,N_28827);
nand UO_1765 (O_1765,N_28109,N_29553);
xor UO_1766 (O_1766,N_29426,N_28758);
and UO_1767 (O_1767,N_28130,N_29298);
nor UO_1768 (O_1768,N_28565,N_29155);
nand UO_1769 (O_1769,N_28822,N_28804);
nand UO_1770 (O_1770,N_29212,N_28483);
or UO_1771 (O_1771,N_28041,N_28161);
and UO_1772 (O_1772,N_29103,N_29465);
and UO_1773 (O_1773,N_28631,N_29333);
nand UO_1774 (O_1774,N_29565,N_28735);
and UO_1775 (O_1775,N_29434,N_28214);
nor UO_1776 (O_1776,N_29819,N_29190);
xnor UO_1777 (O_1777,N_29997,N_28565);
xor UO_1778 (O_1778,N_28415,N_29702);
nand UO_1779 (O_1779,N_28492,N_28502);
nor UO_1780 (O_1780,N_28686,N_29968);
xor UO_1781 (O_1781,N_28589,N_28791);
nor UO_1782 (O_1782,N_28642,N_28420);
nor UO_1783 (O_1783,N_28072,N_29394);
nand UO_1784 (O_1784,N_28237,N_29597);
nand UO_1785 (O_1785,N_29657,N_29481);
and UO_1786 (O_1786,N_28521,N_29451);
nand UO_1787 (O_1787,N_28702,N_29039);
and UO_1788 (O_1788,N_29209,N_29874);
and UO_1789 (O_1789,N_28123,N_29293);
and UO_1790 (O_1790,N_28188,N_29377);
and UO_1791 (O_1791,N_28993,N_28782);
or UO_1792 (O_1792,N_29506,N_28631);
nor UO_1793 (O_1793,N_29948,N_29944);
xor UO_1794 (O_1794,N_29131,N_28844);
or UO_1795 (O_1795,N_28869,N_28477);
and UO_1796 (O_1796,N_28340,N_29002);
or UO_1797 (O_1797,N_29944,N_28043);
xnor UO_1798 (O_1798,N_29878,N_29253);
or UO_1799 (O_1799,N_29183,N_29804);
nand UO_1800 (O_1800,N_29055,N_29159);
xnor UO_1801 (O_1801,N_28121,N_28271);
xor UO_1802 (O_1802,N_29102,N_28845);
xnor UO_1803 (O_1803,N_29935,N_28674);
nand UO_1804 (O_1804,N_28092,N_29847);
nand UO_1805 (O_1805,N_29829,N_29389);
nor UO_1806 (O_1806,N_28453,N_29607);
and UO_1807 (O_1807,N_28705,N_29236);
or UO_1808 (O_1808,N_29450,N_28718);
xnor UO_1809 (O_1809,N_28799,N_29820);
nand UO_1810 (O_1810,N_29860,N_29893);
nor UO_1811 (O_1811,N_28202,N_29114);
xnor UO_1812 (O_1812,N_28911,N_28492);
nand UO_1813 (O_1813,N_29040,N_29896);
xnor UO_1814 (O_1814,N_29261,N_29661);
or UO_1815 (O_1815,N_28777,N_28911);
nor UO_1816 (O_1816,N_28298,N_28609);
xor UO_1817 (O_1817,N_28181,N_29751);
xor UO_1818 (O_1818,N_28148,N_28960);
or UO_1819 (O_1819,N_28476,N_29832);
nor UO_1820 (O_1820,N_28095,N_29828);
nand UO_1821 (O_1821,N_29923,N_28409);
or UO_1822 (O_1822,N_29510,N_28644);
nand UO_1823 (O_1823,N_29459,N_28923);
and UO_1824 (O_1824,N_29104,N_29448);
nand UO_1825 (O_1825,N_29842,N_28677);
nor UO_1826 (O_1826,N_28032,N_28772);
or UO_1827 (O_1827,N_29446,N_29788);
and UO_1828 (O_1828,N_28579,N_29601);
nand UO_1829 (O_1829,N_28885,N_28079);
nand UO_1830 (O_1830,N_28100,N_28786);
and UO_1831 (O_1831,N_28162,N_29139);
nor UO_1832 (O_1832,N_28840,N_29300);
nand UO_1833 (O_1833,N_29570,N_29096);
nand UO_1834 (O_1834,N_29208,N_28617);
or UO_1835 (O_1835,N_29065,N_29094);
xnor UO_1836 (O_1836,N_28971,N_28543);
nor UO_1837 (O_1837,N_28090,N_28760);
xor UO_1838 (O_1838,N_28724,N_28733);
nor UO_1839 (O_1839,N_28662,N_29736);
nor UO_1840 (O_1840,N_29206,N_28068);
and UO_1841 (O_1841,N_29154,N_29203);
or UO_1842 (O_1842,N_28360,N_28548);
or UO_1843 (O_1843,N_28611,N_29117);
nand UO_1844 (O_1844,N_29912,N_28298);
or UO_1845 (O_1845,N_28077,N_29683);
or UO_1846 (O_1846,N_28008,N_29467);
nor UO_1847 (O_1847,N_29606,N_28897);
xnor UO_1848 (O_1848,N_29135,N_28595);
nand UO_1849 (O_1849,N_28289,N_29771);
or UO_1850 (O_1850,N_28974,N_29878);
and UO_1851 (O_1851,N_28177,N_29027);
or UO_1852 (O_1852,N_28789,N_28712);
nor UO_1853 (O_1853,N_29174,N_29874);
nand UO_1854 (O_1854,N_28413,N_28387);
or UO_1855 (O_1855,N_28709,N_29698);
nand UO_1856 (O_1856,N_29498,N_28586);
and UO_1857 (O_1857,N_29554,N_29092);
xor UO_1858 (O_1858,N_28845,N_28488);
nor UO_1859 (O_1859,N_28342,N_28628);
nor UO_1860 (O_1860,N_29435,N_29135);
xor UO_1861 (O_1861,N_28840,N_28997);
xnor UO_1862 (O_1862,N_28668,N_29176);
nor UO_1863 (O_1863,N_29093,N_29756);
or UO_1864 (O_1864,N_28140,N_28905);
nand UO_1865 (O_1865,N_28515,N_29488);
nor UO_1866 (O_1866,N_28480,N_28585);
or UO_1867 (O_1867,N_29428,N_29882);
nor UO_1868 (O_1868,N_29598,N_28771);
or UO_1869 (O_1869,N_29272,N_28974);
xor UO_1870 (O_1870,N_28247,N_28550);
nand UO_1871 (O_1871,N_28991,N_28984);
nand UO_1872 (O_1872,N_28528,N_29517);
nor UO_1873 (O_1873,N_29001,N_29381);
and UO_1874 (O_1874,N_28239,N_28102);
nor UO_1875 (O_1875,N_28387,N_29530);
and UO_1876 (O_1876,N_29513,N_28584);
xnor UO_1877 (O_1877,N_28558,N_28040);
nor UO_1878 (O_1878,N_29375,N_28993);
and UO_1879 (O_1879,N_29813,N_28080);
or UO_1880 (O_1880,N_29900,N_28771);
nor UO_1881 (O_1881,N_29166,N_28503);
nor UO_1882 (O_1882,N_29885,N_29868);
xor UO_1883 (O_1883,N_29020,N_29615);
and UO_1884 (O_1884,N_29673,N_29746);
or UO_1885 (O_1885,N_28931,N_29488);
xnor UO_1886 (O_1886,N_29678,N_29844);
nand UO_1887 (O_1887,N_28752,N_29731);
or UO_1888 (O_1888,N_28728,N_29402);
and UO_1889 (O_1889,N_29841,N_29925);
and UO_1890 (O_1890,N_29176,N_29728);
xnor UO_1891 (O_1891,N_29440,N_29431);
xnor UO_1892 (O_1892,N_29410,N_29826);
or UO_1893 (O_1893,N_29739,N_29117);
xor UO_1894 (O_1894,N_28436,N_29298);
or UO_1895 (O_1895,N_28925,N_29334);
xnor UO_1896 (O_1896,N_28059,N_28241);
xnor UO_1897 (O_1897,N_28584,N_29814);
and UO_1898 (O_1898,N_28616,N_28164);
and UO_1899 (O_1899,N_28732,N_29056);
nor UO_1900 (O_1900,N_28233,N_29781);
nand UO_1901 (O_1901,N_29346,N_29910);
nand UO_1902 (O_1902,N_28388,N_29312);
nor UO_1903 (O_1903,N_29987,N_28522);
xor UO_1904 (O_1904,N_28747,N_29224);
and UO_1905 (O_1905,N_29878,N_28807);
nor UO_1906 (O_1906,N_28843,N_28716);
or UO_1907 (O_1907,N_29768,N_28161);
xor UO_1908 (O_1908,N_29681,N_28528);
and UO_1909 (O_1909,N_29685,N_29973);
xor UO_1910 (O_1910,N_28335,N_29020);
or UO_1911 (O_1911,N_28137,N_29762);
and UO_1912 (O_1912,N_29804,N_28652);
or UO_1913 (O_1913,N_28417,N_29669);
nor UO_1914 (O_1914,N_29187,N_29749);
nor UO_1915 (O_1915,N_29262,N_29326);
xor UO_1916 (O_1916,N_28407,N_28161);
and UO_1917 (O_1917,N_28398,N_28993);
or UO_1918 (O_1918,N_29282,N_28205);
nor UO_1919 (O_1919,N_28141,N_28845);
and UO_1920 (O_1920,N_29315,N_28460);
nand UO_1921 (O_1921,N_29668,N_29879);
nor UO_1922 (O_1922,N_29720,N_29401);
or UO_1923 (O_1923,N_28494,N_28190);
xnor UO_1924 (O_1924,N_29056,N_28728);
xor UO_1925 (O_1925,N_28197,N_28582);
and UO_1926 (O_1926,N_29720,N_28711);
or UO_1927 (O_1927,N_28882,N_28762);
nand UO_1928 (O_1928,N_28410,N_29997);
xor UO_1929 (O_1929,N_28944,N_29063);
and UO_1930 (O_1930,N_28798,N_28852);
or UO_1931 (O_1931,N_29174,N_28583);
xnor UO_1932 (O_1932,N_29748,N_28556);
nor UO_1933 (O_1933,N_28299,N_29456);
nand UO_1934 (O_1934,N_29392,N_29462);
xor UO_1935 (O_1935,N_28099,N_28441);
nor UO_1936 (O_1936,N_28194,N_28023);
nand UO_1937 (O_1937,N_28022,N_28410);
or UO_1938 (O_1938,N_29904,N_29860);
or UO_1939 (O_1939,N_29016,N_29153);
or UO_1940 (O_1940,N_28421,N_29712);
and UO_1941 (O_1941,N_28506,N_28473);
and UO_1942 (O_1942,N_28877,N_28265);
nor UO_1943 (O_1943,N_29626,N_29861);
nand UO_1944 (O_1944,N_28482,N_29689);
or UO_1945 (O_1945,N_28803,N_29577);
xor UO_1946 (O_1946,N_29105,N_28924);
xnor UO_1947 (O_1947,N_28190,N_28285);
nand UO_1948 (O_1948,N_29463,N_28136);
and UO_1949 (O_1949,N_29509,N_28082);
and UO_1950 (O_1950,N_29469,N_29073);
xor UO_1951 (O_1951,N_28732,N_29425);
or UO_1952 (O_1952,N_28083,N_28868);
or UO_1953 (O_1953,N_29017,N_28407);
nor UO_1954 (O_1954,N_28475,N_29285);
and UO_1955 (O_1955,N_28070,N_29358);
nand UO_1956 (O_1956,N_28215,N_29152);
and UO_1957 (O_1957,N_28964,N_28811);
nor UO_1958 (O_1958,N_28291,N_28750);
and UO_1959 (O_1959,N_28754,N_29334);
nand UO_1960 (O_1960,N_28116,N_28098);
nor UO_1961 (O_1961,N_28409,N_29833);
nor UO_1962 (O_1962,N_29473,N_28045);
nand UO_1963 (O_1963,N_29047,N_29623);
nor UO_1964 (O_1964,N_28359,N_28866);
or UO_1965 (O_1965,N_29515,N_29134);
nand UO_1966 (O_1966,N_29005,N_29341);
xor UO_1967 (O_1967,N_29434,N_29734);
and UO_1968 (O_1968,N_29266,N_29286);
and UO_1969 (O_1969,N_28809,N_28838);
nor UO_1970 (O_1970,N_29550,N_29241);
or UO_1971 (O_1971,N_28801,N_29237);
nor UO_1972 (O_1972,N_29072,N_28098);
or UO_1973 (O_1973,N_29077,N_28588);
and UO_1974 (O_1974,N_29804,N_28940);
or UO_1975 (O_1975,N_29232,N_29112);
nor UO_1976 (O_1976,N_29390,N_29355);
xnor UO_1977 (O_1977,N_28371,N_28347);
xnor UO_1978 (O_1978,N_29110,N_28431);
or UO_1979 (O_1979,N_28720,N_29011);
nor UO_1980 (O_1980,N_29884,N_29630);
nor UO_1981 (O_1981,N_29873,N_29535);
and UO_1982 (O_1982,N_29692,N_28661);
nor UO_1983 (O_1983,N_28470,N_29910);
or UO_1984 (O_1984,N_28383,N_29496);
or UO_1985 (O_1985,N_29371,N_29539);
nor UO_1986 (O_1986,N_28044,N_28982);
nor UO_1987 (O_1987,N_28379,N_28479);
and UO_1988 (O_1988,N_29074,N_29463);
nor UO_1989 (O_1989,N_28775,N_28880);
xor UO_1990 (O_1990,N_28814,N_28854);
and UO_1991 (O_1991,N_28023,N_28490);
or UO_1992 (O_1992,N_28439,N_28143);
nor UO_1993 (O_1993,N_29638,N_28906);
nand UO_1994 (O_1994,N_29375,N_29029);
xnor UO_1995 (O_1995,N_29124,N_28821);
nand UO_1996 (O_1996,N_29128,N_28794);
xor UO_1997 (O_1997,N_28590,N_29149);
nor UO_1998 (O_1998,N_29979,N_29918);
nand UO_1999 (O_1999,N_28739,N_28367);
nor UO_2000 (O_2000,N_28608,N_28467);
and UO_2001 (O_2001,N_29709,N_29331);
nor UO_2002 (O_2002,N_28703,N_29172);
nand UO_2003 (O_2003,N_28935,N_29987);
xnor UO_2004 (O_2004,N_29665,N_29710);
xnor UO_2005 (O_2005,N_28411,N_29547);
xor UO_2006 (O_2006,N_29992,N_28615);
and UO_2007 (O_2007,N_28415,N_29725);
and UO_2008 (O_2008,N_28853,N_29994);
xor UO_2009 (O_2009,N_28969,N_29445);
nand UO_2010 (O_2010,N_28697,N_28982);
xnor UO_2011 (O_2011,N_29125,N_29457);
and UO_2012 (O_2012,N_29767,N_29340);
or UO_2013 (O_2013,N_28358,N_28837);
and UO_2014 (O_2014,N_28913,N_28091);
or UO_2015 (O_2015,N_29410,N_28900);
and UO_2016 (O_2016,N_29296,N_29083);
nand UO_2017 (O_2017,N_29537,N_28541);
nor UO_2018 (O_2018,N_29077,N_29488);
xnor UO_2019 (O_2019,N_28087,N_29384);
and UO_2020 (O_2020,N_29574,N_28082);
nor UO_2021 (O_2021,N_29368,N_29845);
nor UO_2022 (O_2022,N_29679,N_28149);
nand UO_2023 (O_2023,N_28681,N_28649);
xnor UO_2024 (O_2024,N_28984,N_29596);
nor UO_2025 (O_2025,N_29582,N_28616);
nand UO_2026 (O_2026,N_29330,N_29419);
or UO_2027 (O_2027,N_28309,N_29885);
nor UO_2028 (O_2028,N_28480,N_28500);
nand UO_2029 (O_2029,N_29395,N_28260);
nor UO_2030 (O_2030,N_29758,N_29740);
nor UO_2031 (O_2031,N_29776,N_28605);
and UO_2032 (O_2032,N_28954,N_28552);
and UO_2033 (O_2033,N_28953,N_29030);
xnor UO_2034 (O_2034,N_28340,N_29076);
nor UO_2035 (O_2035,N_29526,N_29278);
nor UO_2036 (O_2036,N_28008,N_28335);
or UO_2037 (O_2037,N_29974,N_29794);
and UO_2038 (O_2038,N_29124,N_28850);
nor UO_2039 (O_2039,N_28968,N_29781);
nand UO_2040 (O_2040,N_28157,N_29334);
or UO_2041 (O_2041,N_29896,N_28809);
xor UO_2042 (O_2042,N_28348,N_29164);
nor UO_2043 (O_2043,N_28892,N_28514);
nand UO_2044 (O_2044,N_29684,N_28121);
or UO_2045 (O_2045,N_29248,N_28275);
nor UO_2046 (O_2046,N_28872,N_28698);
nor UO_2047 (O_2047,N_29984,N_28829);
nor UO_2048 (O_2048,N_28029,N_28698);
and UO_2049 (O_2049,N_28073,N_29172);
nand UO_2050 (O_2050,N_28471,N_28361);
nand UO_2051 (O_2051,N_28615,N_29767);
nor UO_2052 (O_2052,N_28501,N_28554);
or UO_2053 (O_2053,N_28123,N_28501);
or UO_2054 (O_2054,N_28289,N_28707);
nand UO_2055 (O_2055,N_29649,N_29983);
or UO_2056 (O_2056,N_28683,N_29782);
nor UO_2057 (O_2057,N_28649,N_29585);
and UO_2058 (O_2058,N_29667,N_29484);
xnor UO_2059 (O_2059,N_28195,N_29061);
nor UO_2060 (O_2060,N_28621,N_28119);
and UO_2061 (O_2061,N_29569,N_28447);
xnor UO_2062 (O_2062,N_29193,N_28491);
nand UO_2063 (O_2063,N_28652,N_29715);
or UO_2064 (O_2064,N_29505,N_29986);
nor UO_2065 (O_2065,N_28820,N_29044);
xor UO_2066 (O_2066,N_28384,N_28732);
xnor UO_2067 (O_2067,N_29696,N_29489);
and UO_2068 (O_2068,N_28525,N_28041);
and UO_2069 (O_2069,N_28387,N_28191);
nor UO_2070 (O_2070,N_28553,N_28592);
xnor UO_2071 (O_2071,N_29712,N_29298);
and UO_2072 (O_2072,N_29209,N_29980);
or UO_2073 (O_2073,N_29099,N_28245);
nor UO_2074 (O_2074,N_29690,N_28776);
nand UO_2075 (O_2075,N_28552,N_29357);
nor UO_2076 (O_2076,N_28987,N_28297);
and UO_2077 (O_2077,N_29717,N_29881);
nor UO_2078 (O_2078,N_28572,N_28663);
nand UO_2079 (O_2079,N_29239,N_28247);
nand UO_2080 (O_2080,N_28580,N_29342);
or UO_2081 (O_2081,N_29291,N_29500);
xnor UO_2082 (O_2082,N_28409,N_28265);
nand UO_2083 (O_2083,N_28219,N_28400);
and UO_2084 (O_2084,N_29960,N_28924);
nor UO_2085 (O_2085,N_29821,N_28465);
nand UO_2086 (O_2086,N_28342,N_28172);
or UO_2087 (O_2087,N_28698,N_28975);
nor UO_2088 (O_2088,N_28157,N_28554);
nor UO_2089 (O_2089,N_29214,N_29308);
or UO_2090 (O_2090,N_29927,N_29040);
nand UO_2091 (O_2091,N_28548,N_29487);
xor UO_2092 (O_2092,N_29131,N_28968);
and UO_2093 (O_2093,N_28713,N_29177);
or UO_2094 (O_2094,N_28493,N_29268);
or UO_2095 (O_2095,N_29818,N_28537);
and UO_2096 (O_2096,N_29863,N_28185);
xor UO_2097 (O_2097,N_28764,N_28477);
xnor UO_2098 (O_2098,N_29061,N_29843);
nand UO_2099 (O_2099,N_28381,N_29908);
nor UO_2100 (O_2100,N_28692,N_29989);
or UO_2101 (O_2101,N_28738,N_29860);
xor UO_2102 (O_2102,N_29570,N_28187);
xnor UO_2103 (O_2103,N_28290,N_29026);
and UO_2104 (O_2104,N_29032,N_29844);
and UO_2105 (O_2105,N_28760,N_29768);
nor UO_2106 (O_2106,N_28643,N_29359);
or UO_2107 (O_2107,N_29363,N_28697);
and UO_2108 (O_2108,N_29803,N_29608);
nand UO_2109 (O_2109,N_29498,N_28889);
or UO_2110 (O_2110,N_29762,N_29520);
or UO_2111 (O_2111,N_29434,N_29036);
and UO_2112 (O_2112,N_28703,N_28193);
xor UO_2113 (O_2113,N_29861,N_29169);
and UO_2114 (O_2114,N_28981,N_29262);
and UO_2115 (O_2115,N_29738,N_29688);
nand UO_2116 (O_2116,N_28200,N_29589);
nand UO_2117 (O_2117,N_28170,N_28057);
and UO_2118 (O_2118,N_29725,N_28500);
or UO_2119 (O_2119,N_29031,N_29887);
and UO_2120 (O_2120,N_28187,N_28233);
and UO_2121 (O_2121,N_29382,N_29248);
nand UO_2122 (O_2122,N_29986,N_28438);
nor UO_2123 (O_2123,N_28741,N_29834);
nand UO_2124 (O_2124,N_28900,N_29161);
nand UO_2125 (O_2125,N_28186,N_29301);
nand UO_2126 (O_2126,N_29775,N_28746);
and UO_2127 (O_2127,N_28553,N_29994);
or UO_2128 (O_2128,N_29791,N_28330);
nand UO_2129 (O_2129,N_29723,N_28367);
nand UO_2130 (O_2130,N_29921,N_28192);
nor UO_2131 (O_2131,N_28372,N_29087);
and UO_2132 (O_2132,N_28708,N_28205);
nand UO_2133 (O_2133,N_28590,N_29560);
xnor UO_2134 (O_2134,N_28155,N_28749);
or UO_2135 (O_2135,N_29390,N_29557);
nand UO_2136 (O_2136,N_29874,N_29646);
and UO_2137 (O_2137,N_28751,N_28969);
nand UO_2138 (O_2138,N_28837,N_29114);
and UO_2139 (O_2139,N_29161,N_29915);
nor UO_2140 (O_2140,N_28236,N_28660);
xor UO_2141 (O_2141,N_28974,N_28738);
or UO_2142 (O_2142,N_29873,N_29042);
nor UO_2143 (O_2143,N_28141,N_29466);
nand UO_2144 (O_2144,N_29437,N_29455);
nand UO_2145 (O_2145,N_28015,N_28171);
xnor UO_2146 (O_2146,N_29874,N_29112);
or UO_2147 (O_2147,N_29016,N_28603);
or UO_2148 (O_2148,N_28549,N_29306);
or UO_2149 (O_2149,N_29382,N_29245);
xnor UO_2150 (O_2150,N_28322,N_29380);
or UO_2151 (O_2151,N_28187,N_29336);
xor UO_2152 (O_2152,N_28680,N_29580);
and UO_2153 (O_2153,N_28248,N_28307);
nor UO_2154 (O_2154,N_28902,N_28068);
or UO_2155 (O_2155,N_29008,N_29177);
and UO_2156 (O_2156,N_29696,N_28323);
xnor UO_2157 (O_2157,N_28999,N_28312);
nor UO_2158 (O_2158,N_28209,N_28352);
and UO_2159 (O_2159,N_29083,N_29659);
xor UO_2160 (O_2160,N_28734,N_28128);
nor UO_2161 (O_2161,N_28966,N_28448);
and UO_2162 (O_2162,N_29097,N_28724);
xnor UO_2163 (O_2163,N_29559,N_29177);
nand UO_2164 (O_2164,N_29224,N_28962);
nand UO_2165 (O_2165,N_29739,N_28010);
nor UO_2166 (O_2166,N_29913,N_29902);
or UO_2167 (O_2167,N_28895,N_29917);
and UO_2168 (O_2168,N_28076,N_29083);
nand UO_2169 (O_2169,N_28975,N_29354);
and UO_2170 (O_2170,N_28741,N_28426);
and UO_2171 (O_2171,N_29186,N_28115);
or UO_2172 (O_2172,N_29369,N_28279);
nand UO_2173 (O_2173,N_29841,N_29302);
nor UO_2174 (O_2174,N_29628,N_28279);
or UO_2175 (O_2175,N_29956,N_29972);
or UO_2176 (O_2176,N_28101,N_28686);
nand UO_2177 (O_2177,N_29091,N_28620);
xor UO_2178 (O_2178,N_28025,N_29031);
nor UO_2179 (O_2179,N_29061,N_28279);
nand UO_2180 (O_2180,N_28404,N_28945);
nand UO_2181 (O_2181,N_28721,N_28435);
nor UO_2182 (O_2182,N_28639,N_28050);
and UO_2183 (O_2183,N_28182,N_29299);
nand UO_2184 (O_2184,N_29150,N_29505);
and UO_2185 (O_2185,N_29794,N_29978);
nor UO_2186 (O_2186,N_29960,N_28989);
or UO_2187 (O_2187,N_29025,N_29301);
nor UO_2188 (O_2188,N_29973,N_29317);
nor UO_2189 (O_2189,N_29121,N_29975);
or UO_2190 (O_2190,N_28757,N_28765);
nor UO_2191 (O_2191,N_28109,N_28323);
and UO_2192 (O_2192,N_28221,N_29943);
or UO_2193 (O_2193,N_29854,N_28134);
xor UO_2194 (O_2194,N_29762,N_29279);
and UO_2195 (O_2195,N_28719,N_29133);
and UO_2196 (O_2196,N_29370,N_29907);
nor UO_2197 (O_2197,N_29159,N_29761);
nor UO_2198 (O_2198,N_29619,N_29409);
nand UO_2199 (O_2199,N_28960,N_28719);
nand UO_2200 (O_2200,N_29966,N_28471);
xnor UO_2201 (O_2201,N_28435,N_29294);
nor UO_2202 (O_2202,N_29731,N_29239);
xnor UO_2203 (O_2203,N_28007,N_28906);
xnor UO_2204 (O_2204,N_28908,N_29580);
and UO_2205 (O_2205,N_28086,N_29626);
and UO_2206 (O_2206,N_28689,N_29023);
and UO_2207 (O_2207,N_28211,N_28697);
xnor UO_2208 (O_2208,N_28037,N_29988);
nand UO_2209 (O_2209,N_29426,N_29115);
nand UO_2210 (O_2210,N_28501,N_29217);
or UO_2211 (O_2211,N_29920,N_28018);
nor UO_2212 (O_2212,N_29046,N_28810);
xnor UO_2213 (O_2213,N_28450,N_28418);
xor UO_2214 (O_2214,N_28955,N_28394);
and UO_2215 (O_2215,N_28987,N_29502);
and UO_2216 (O_2216,N_29967,N_28009);
nand UO_2217 (O_2217,N_28003,N_28698);
nand UO_2218 (O_2218,N_28420,N_28826);
nor UO_2219 (O_2219,N_28015,N_28090);
nor UO_2220 (O_2220,N_29261,N_28581);
and UO_2221 (O_2221,N_28774,N_29052);
xor UO_2222 (O_2222,N_28353,N_28307);
nor UO_2223 (O_2223,N_28735,N_28846);
nand UO_2224 (O_2224,N_29969,N_28378);
or UO_2225 (O_2225,N_28857,N_28115);
or UO_2226 (O_2226,N_29797,N_28505);
or UO_2227 (O_2227,N_29528,N_28501);
nor UO_2228 (O_2228,N_29203,N_28174);
nand UO_2229 (O_2229,N_28440,N_28222);
nor UO_2230 (O_2230,N_28315,N_28863);
or UO_2231 (O_2231,N_28802,N_29501);
xor UO_2232 (O_2232,N_29743,N_29638);
nand UO_2233 (O_2233,N_29044,N_28538);
and UO_2234 (O_2234,N_28283,N_28187);
or UO_2235 (O_2235,N_28763,N_28035);
nor UO_2236 (O_2236,N_28601,N_28520);
nor UO_2237 (O_2237,N_29794,N_28109);
and UO_2238 (O_2238,N_29257,N_29410);
or UO_2239 (O_2239,N_29902,N_28480);
and UO_2240 (O_2240,N_28653,N_28740);
nand UO_2241 (O_2241,N_28030,N_28548);
and UO_2242 (O_2242,N_28216,N_28581);
and UO_2243 (O_2243,N_29022,N_28425);
xor UO_2244 (O_2244,N_29921,N_29989);
and UO_2245 (O_2245,N_28810,N_28478);
nand UO_2246 (O_2246,N_28780,N_28450);
xnor UO_2247 (O_2247,N_29393,N_29617);
nand UO_2248 (O_2248,N_29368,N_28549);
or UO_2249 (O_2249,N_28493,N_29850);
nor UO_2250 (O_2250,N_28538,N_28743);
and UO_2251 (O_2251,N_28788,N_29447);
nand UO_2252 (O_2252,N_28149,N_29458);
or UO_2253 (O_2253,N_29174,N_28862);
nand UO_2254 (O_2254,N_29010,N_29155);
and UO_2255 (O_2255,N_29425,N_29267);
and UO_2256 (O_2256,N_29857,N_29193);
and UO_2257 (O_2257,N_29217,N_29348);
nor UO_2258 (O_2258,N_28672,N_28193);
or UO_2259 (O_2259,N_29004,N_28068);
and UO_2260 (O_2260,N_29687,N_29876);
xnor UO_2261 (O_2261,N_28986,N_28344);
nor UO_2262 (O_2262,N_28679,N_29690);
xnor UO_2263 (O_2263,N_29230,N_29820);
nand UO_2264 (O_2264,N_28044,N_28287);
nor UO_2265 (O_2265,N_28555,N_29089);
nand UO_2266 (O_2266,N_29342,N_28866);
nand UO_2267 (O_2267,N_29622,N_29418);
nor UO_2268 (O_2268,N_29269,N_28269);
and UO_2269 (O_2269,N_28044,N_29576);
xnor UO_2270 (O_2270,N_29365,N_28042);
and UO_2271 (O_2271,N_29885,N_28330);
and UO_2272 (O_2272,N_28539,N_28037);
or UO_2273 (O_2273,N_29359,N_28901);
or UO_2274 (O_2274,N_29254,N_28626);
xor UO_2275 (O_2275,N_28705,N_29981);
or UO_2276 (O_2276,N_29065,N_29325);
nand UO_2277 (O_2277,N_29811,N_29024);
or UO_2278 (O_2278,N_29353,N_28832);
or UO_2279 (O_2279,N_29460,N_28640);
nor UO_2280 (O_2280,N_29267,N_29334);
or UO_2281 (O_2281,N_29078,N_28605);
or UO_2282 (O_2282,N_28788,N_28389);
nor UO_2283 (O_2283,N_28955,N_28680);
and UO_2284 (O_2284,N_28249,N_28453);
nand UO_2285 (O_2285,N_29667,N_29338);
or UO_2286 (O_2286,N_29761,N_29835);
or UO_2287 (O_2287,N_29359,N_28347);
nand UO_2288 (O_2288,N_29222,N_28037);
and UO_2289 (O_2289,N_29101,N_29414);
or UO_2290 (O_2290,N_29812,N_28468);
nor UO_2291 (O_2291,N_29448,N_29582);
and UO_2292 (O_2292,N_29326,N_29193);
nand UO_2293 (O_2293,N_28692,N_29760);
xor UO_2294 (O_2294,N_29165,N_28429);
or UO_2295 (O_2295,N_29547,N_29659);
or UO_2296 (O_2296,N_29493,N_28575);
nor UO_2297 (O_2297,N_28756,N_28271);
or UO_2298 (O_2298,N_28589,N_29225);
nand UO_2299 (O_2299,N_29820,N_29816);
nor UO_2300 (O_2300,N_29004,N_28365);
nor UO_2301 (O_2301,N_29962,N_28199);
or UO_2302 (O_2302,N_28877,N_29295);
nor UO_2303 (O_2303,N_29847,N_28829);
nand UO_2304 (O_2304,N_29585,N_28466);
or UO_2305 (O_2305,N_29210,N_29231);
xor UO_2306 (O_2306,N_29388,N_28422);
and UO_2307 (O_2307,N_29370,N_29924);
or UO_2308 (O_2308,N_28358,N_29701);
or UO_2309 (O_2309,N_28564,N_28622);
nor UO_2310 (O_2310,N_28272,N_29514);
nand UO_2311 (O_2311,N_29888,N_28003);
xnor UO_2312 (O_2312,N_28781,N_29050);
or UO_2313 (O_2313,N_28497,N_28750);
and UO_2314 (O_2314,N_29104,N_28469);
and UO_2315 (O_2315,N_28985,N_29237);
nor UO_2316 (O_2316,N_28272,N_28803);
xnor UO_2317 (O_2317,N_29760,N_29939);
nor UO_2318 (O_2318,N_28986,N_28068);
nand UO_2319 (O_2319,N_29471,N_28164);
nor UO_2320 (O_2320,N_29321,N_28265);
nand UO_2321 (O_2321,N_29306,N_28483);
nor UO_2322 (O_2322,N_28639,N_29088);
xor UO_2323 (O_2323,N_28512,N_28945);
xnor UO_2324 (O_2324,N_29670,N_29820);
xor UO_2325 (O_2325,N_29213,N_28061);
nor UO_2326 (O_2326,N_29829,N_29185);
and UO_2327 (O_2327,N_28561,N_28821);
and UO_2328 (O_2328,N_29953,N_28789);
and UO_2329 (O_2329,N_28679,N_29719);
or UO_2330 (O_2330,N_29457,N_29197);
nand UO_2331 (O_2331,N_28189,N_28693);
nand UO_2332 (O_2332,N_29023,N_28759);
and UO_2333 (O_2333,N_28394,N_29401);
and UO_2334 (O_2334,N_29282,N_29564);
nand UO_2335 (O_2335,N_29279,N_28733);
and UO_2336 (O_2336,N_28666,N_29774);
nand UO_2337 (O_2337,N_28281,N_29642);
xor UO_2338 (O_2338,N_29120,N_28272);
xnor UO_2339 (O_2339,N_28231,N_29091);
and UO_2340 (O_2340,N_29187,N_29921);
nor UO_2341 (O_2341,N_28268,N_28304);
nand UO_2342 (O_2342,N_28577,N_29052);
nand UO_2343 (O_2343,N_28138,N_28088);
nand UO_2344 (O_2344,N_28297,N_29375);
nand UO_2345 (O_2345,N_29284,N_29298);
nand UO_2346 (O_2346,N_29061,N_29407);
nor UO_2347 (O_2347,N_29463,N_29175);
or UO_2348 (O_2348,N_29844,N_28120);
or UO_2349 (O_2349,N_29144,N_29410);
xnor UO_2350 (O_2350,N_29489,N_29558);
xor UO_2351 (O_2351,N_29270,N_28851);
xor UO_2352 (O_2352,N_29092,N_28290);
and UO_2353 (O_2353,N_29181,N_28742);
nand UO_2354 (O_2354,N_28114,N_28803);
nor UO_2355 (O_2355,N_29891,N_28227);
xnor UO_2356 (O_2356,N_28424,N_28641);
xor UO_2357 (O_2357,N_29871,N_28358);
nor UO_2358 (O_2358,N_28045,N_28756);
or UO_2359 (O_2359,N_28431,N_28224);
nor UO_2360 (O_2360,N_28473,N_29567);
nor UO_2361 (O_2361,N_29508,N_28080);
nand UO_2362 (O_2362,N_29889,N_29503);
nor UO_2363 (O_2363,N_29355,N_29456);
nand UO_2364 (O_2364,N_28593,N_29459);
xor UO_2365 (O_2365,N_29142,N_29667);
or UO_2366 (O_2366,N_28745,N_29584);
nand UO_2367 (O_2367,N_29392,N_29075);
nor UO_2368 (O_2368,N_28990,N_28252);
and UO_2369 (O_2369,N_29388,N_29696);
nor UO_2370 (O_2370,N_28179,N_29590);
nand UO_2371 (O_2371,N_29388,N_28731);
nand UO_2372 (O_2372,N_28954,N_28131);
or UO_2373 (O_2373,N_29345,N_29087);
nand UO_2374 (O_2374,N_29127,N_29330);
xnor UO_2375 (O_2375,N_28112,N_28009);
nor UO_2376 (O_2376,N_29696,N_28954);
xor UO_2377 (O_2377,N_28963,N_28005);
nand UO_2378 (O_2378,N_29019,N_28983);
or UO_2379 (O_2379,N_28881,N_29251);
nor UO_2380 (O_2380,N_28146,N_29662);
or UO_2381 (O_2381,N_28985,N_28961);
and UO_2382 (O_2382,N_28266,N_28288);
nand UO_2383 (O_2383,N_28192,N_28620);
and UO_2384 (O_2384,N_29947,N_29852);
nor UO_2385 (O_2385,N_29958,N_29723);
or UO_2386 (O_2386,N_28756,N_29132);
or UO_2387 (O_2387,N_29955,N_29264);
nand UO_2388 (O_2388,N_28752,N_28671);
nand UO_2389 (O_2389,N_28503,N_29398);
or UO_2390 (O_2390,N_28263,N_28910);
xor UO_2391 (O_2391,N_29735,N_28509);
xor UO_2392 (O_2392,N_29994,N_28496);
or UO_2393 (O_2393,N_28145,N_29734);
and UO_2394 (O_2394,N_28356,N_29961);
or UO_2395 (O_2395,N_28891,N_29237);
nand UO_2396 (O_2396,N_29678,N_29735);
xnor UO_2397 (O_2397,N_28588,N_29572);
xnor UO_2398 (O_2398,N_29397,N_29839);
xor UO_2399 (O_2399,N_29841,N_29629);
and UO_2400 (O_2400,N_28798,N_29423);
or UO_2401 (O_2401,N_29782,N_29272);
nor UO_2402 (O_2402,N_29840,N_28108);
or UO_2403 (O_2403,N_29704,N_28161);
nor UO_2404 (O_2404,N_29183,N_28479);
or UO_2405 (O_2405,N_29661,N_28182);
xor UO_2406 (O_2406,N_28788,N_28905);
and UO_2407 (O_2407,N_28821,N_29716);
xnor UO_2408 (O_2408,N_28290,N_29839);
and UO_2409 (O_2409,N_29492,N_28645);
and UO_2410 (O_2410,N_29327,N_28274);
xor UO_2411 (O_2411,N_29329,N_29133);
nor UO_2412 (O_2412,N_29119,N_28712);
xor UO_2413 (O_2413,N_28665,N_29980);
nand UO_2414 (O_2414,N_28508,N_28148);
and UO_2415 (O_2415,N_29738,N_28626);
nand UO_2416 (O_2416,N_28416,N_29466);
or UO_2417 (O_2417,N_29848,N_28307);
xor UO_2418 (O_2418,N_29681,N_29292);
xor UO_2419 (O_2419,N_29057,N_29595);
and UO_2420 (O_2420,N_28326,N_29413);
nand UO_2421 (O_2421,N_28364,N_29425);
nor UO_2422 (O_2422,N_29716,N_28645);
and UO_2423 (O_2423,N_28884,N_29837);
nor UO_2424 (O_2424,N_29022,N_29453);
nand UO_2425 (O_2425,N_29378,N_28635);
or UO_2426 (O_2426,N_28948,N_29702);
xnor UO_2427 (O_2427,N_29307,N_29117);
or UO_2428 (O_2428,N_28634,N_29103);
xor UO_2429 (O_2429,N_29590,N_29310);
nor UO_2430 (O_2430,N_28606,N_28088);
and UO_2431 (O_2431,N_28772,N_29049);
and UO_2432 (O_2432,N_28291,N_28582);
nand UO_2433 (O_2433,N_29050,N_29078);
nand UO_2434 (O_2434,N_28444,N_28484);
nor UO_2435 (O_2435,N_29874,N_29886);
xor UO_2436 (O_2436,N_28620,N_29554);
nor UO_2437 (O_2437,N_29502,N_28111);
xnor UO_2438 (O_2438,N_29793,N_28744);
nand UO_2439 (O_2439,N_28189,N_29959);
xnor UO_2440 (O_2440,N_28109,N_29296);
and UO_2441 (O_2441,N_29410,N_29313);
or UO_2442 (O_2442,N_29256,N_29452);
nor UO_2443 (O_2443,N_28621,N_28031);
xor UO_2444 (O_2444,N_29260,N_28081);
nand UO_2445 (O_2445,N_29318,N_28165);
nor UO_2446 (O_2446,N_28068,N_28703);
nand UO_2447 (O_2447,N_28037,N_29841);
nor UO_2448 (O_2448,N_29154,N_28745);
nor UO_2449 (O_2449,N_29565,N_28474);
nor UO_2450 (O_2450,N_28149,N_28926);
and UO_2451 (O_2451,N_28122,N_29208);
nor UO_2452 (O_2452,N_29820,N_28730);
or UO_2453 (O_2453,N_29683,N_29123);
nand UO_2454 (O_2454,N_28079,N_28444);
nand UO_2455 (O_2455,N_28162,N_28276);
and UO_2456 (O_2456,N_29075,N_28379);
nor UO_2457 (O_2457,N_29700,N_28225);
nor UO_2458 (O_2458,N_28518,N_28131);
nor UO_2459 (O_2459,N_29961,N_29535);
or UO_2460 (O_2460,N_28259,N_29839);
nand UO_2461 (O_2461,N_28135,N_28472);
or UO_2462 (O_2462,N_28704,N_29322);
xor UO_2463 (O_2463,N_29643,N_28226);
or UO_2464 (O_2464,N_29897,N_28154);
nand UO_2465 (O_2465,N_29264,N_28714);
nor UO_2466 (O_2466,N_29816,N_28694);
or UO_2467 (O_2467,N_28780,N_29156);
nor UO_2468 (O_2468,N_29590,N_29100);
or UO_2469 (O_2469,N_29559,N_29075);
nor UO_2470 (O_2470,N_29193,N_29899);
nand UO_2471 (O_2471,N_28775,N_28418);
and UO_2472 (O_2472,N_29001,N_29105);
nand UO_2473 (O_2473,N_29286,N_28820);
nand UO_2474 (O_2474,N_28375,N_28832);
xnor UO_2475 (O_2475,N_28684,N_29287);
or UO_2476 (O_2476,N_29163,N_28752);
and UO_2477 (O_2477,N_29062,N_29415);
and UO_2478 (O_2478,N_29866,N_28370);
nor UO_2479 (O_2479,N_29428,N_28268);
and UO_2480 (O_2480,N_29121,N_29412);
or UO_2481 (O_2481,N_29235,N_28761);
and UO_2482 (O_2482,N_29598,N_29369);
or UO_2483 (O_2483,N_29743,N_29616);
or UO_2484 (O_2484,N_28287,N_29829);
xor UO_2485 (O_2485,N_29022,N_28961);
or UO_2486 (O_2486,N_29645,N_28668);
nand UO_2487 (O_2487,N_29415,N_29224);
nor UO_2488 (O_2488,N_29054,N_29518);
or UO_2489 (O_2489,N_28390,N_29918);
nand UO_2490 (O_2490,N_29204,N_28871);
xor UO_2491 (O_2491,N_29554,N_28828);
nand UO_2492 (O_2492,N_28225,N_28640);
and UO_2493 (O_2493,N_29640,N_28019);
and UO_2494 (O_2494,N_29334,N_28063);
or UO_2495 (O_2495,N_28558,N_28786);
xor UO_2496 (O_2496,N_29045,N_28980);
or UO_2497 (O_2497,N_28044,N_28748);
nand UO_2498 (O_2498,N_29711,N_28329);
nor UO_2499 (O_2499,N_29652,N_29079);
or UO_2500 (O_2500,N_28849,N_29919);
and UO_2501 (O_2501,N_29375,N_29879);
xor UO_2502 (O_2502,N_28615,N_29034);
and UO_2503 (O_2503,N_28901,N_29987);
and UO_2504 (O_2504,N_28573,N_28804);
nor UO_2505 (O_2505,N_29881,N_29081);
nand UO_2506 (O_2506,N_29023,N_28116);
xor UO_2507 (O_2507,N_28674,N_28156);
nand UO_2508 (O_2508,N_29679,N_29488);
xor UO_2509 (O_2509,N_29798,N_28676);
nand UO_2510 (O_2510,N_29087,N_29546);
xor UO_2511 (O_2511,N_28744,N_29372);
or UO_2512 (O_2512,N_28252,N_29343);
xnor UO_2513 (O_2513,N_28349,N_28359);
and UO_2514 (O_2514,N_28129,N_28943);
nor UO_2515 (O_2515,N_29306,N_28984);
and UO_2516 (O_2516,N_28472,N_28609);
xnor UO_2517 (O_2517,N_29649,N_28305);
nand UO_2518 (O_2518,N_28483,N_29699);
xnor UO_2519 (O_2519,N_29752,N_28072);
or UO_2520 (O_2520,N_29191,N_28045);
or UO_2521 (O_2521,N_29434,N_29028);
nor UO_2522 (O_2522,N_29508,N_28473);
nor UO_2523 (O_2523,N_29477,N_28306);
xor UO_2524 (O_2524,N_29151,N_29067);
nor UO_2525 (O_2525,N_29676,N_28840);
and UO_2526 (O_2526,N_28725,N_29250);
nand UO_2527 (O_2527,N_29929,N_28454);
and UO_2528 (O_2528,N_29805,N_29611);
or UO_2529 (O_2529,N_29658,N_29981);
xnor UO_2530 (O_2530,N_29247,N_28021);
and UO_2531 (O_2531,N_28608,N_29408);
nor UO_2532 (O_2532,N_28160,N_28833);
nor UO_2533 (O_2533,N_29015,N_29297);
xor UO_2534 (O_2534,N_29494,N_28880);
or UO_2535 (O_2535,N_29568,N_28353);
xor UO_2536 (O_2536,N_29415,N_29969);
nor UO_2537 (O_2537,N_29681,N_28727);
and UO_2538 (O_2538,N_28571,N_28587);
xor UO_2539 (O_2539,N_28645,N_29835);
xnor UO_2540 (O_2540,N_28902,N_28836);
and UO_2541 (O_2541,N_29838,N_28602);
and UO_2542 (O_2542,N_28220,N_29343);
nand UO_2543 (O_2543,N_29215,N_29956);
nand UO_2544 (O_2544,N_29793,N_29409);
xor UO_2545 (O_2545,N_29000,N_29628);
nor UO_2546 (O_2546,N_28028,N_29224);
and UO_2547 (O_2547,N_29716,N_29075);
or UO_2548 (O_2548,N_28485,N_28414);
and UO_2549 (O_2549,N_28385,N_29211);
nor UO_2550 (O_2550,N_29743,N_29087);
and UO_2551 (O_2551,N_28122,N_28232);
nand UO_2552 (O_2552,N_29003,N_28469);
and UO_2553 (O_2553,N_29000,N_28501);
and UO_2554 (O_2554,N_28070,N_28560);
and UO_2555 (O_2555,N_29584,N_28646);
xnor UO_2556 (O_2556,N_29073,N_29925);
nor UO_2557 (O_2557,N_28399,N_29556);
or UO_2558 (O_2558,N_28227,N_28446);
or UO_2559 (O_2559,N_29786,N_29724);
nor UO_2560 (O_2560,N_29625,N_28253);
or UO_2561 (O_2561,N_29916,N_29817);
and UO_2562 (O_2562,N_29587,N_29510);
and UO_2563 (O_2563,N_28423,N_28791);
and UO_2564 (O_2564,N_28743,N_28732);
xor UO_2565 (O_2565,N_28744,N_29842);
or UO_2566 (O_2566,N_28830,N_28270);
nor UO_2567 (O_2567,N_28252,N_29919);
xnor UO_2568 (O_2568,N_28660,N_29443);
or UO_2569 (O_2569,N_28162,N_28653);
nor UO_2570 (O_2570,N_28713,N_28211);
and UO_2571 (O_2571,N_29389,N_29012);
and UO_2572 (O_2572,N_28316,N_28619);
and UO_2573 (O_2573,N_28079,N_29220);
or UO_2574 (O_2574,N_29408,N_29776);
nand UO_2575 (O_2575,N_28714,N_28553);
nor UO_2576 (O_2576,N_29492,N_29447);
nor UO_2577 (O_2577,N_28283,N_29734);
xor UO_2578 (O_2578,N_28673,N_29457);
xnor UO_2579 (O_2579,N_28685,N_29326);
and UO_2580 (O_2580,N_28033,N_28613);
or UO_2581 (O_2581,N_28449,N_29352);
nand UO_2582 (O_2582,N_28765,N_28024);
and UO_2583 (O_2583,N_28224,N_28844);
xnor UO_2584 (O_2584,N_28648,N_29746);
or UO_2585 (O_2585,N_28500,N_29785);
nand UO_2586 (O_2586,N_29485,N_28978);
xor UO_2587 (O_2587,N_29503,N_29901);
nand UO_2588 (O_2588,N_28026,N_28181);
nor UO_2589 (O_2589,N_29349,N_29191);
nand UO_2590 (O_2590,N_28840,N_29866);
and UO_2591 (O_2591,N_28974,N_29189);
and UO_2592 (O_2592,N_28978,N_28069);
xor UO_2593 (O_2593,N_29159,N_29852);
xor UO_2594 (O_2594,N_29280,N_29279);
or UO_2595 (O_2595,N_28336,N_29205);
or UO_2596 (O_2596,N_29619,N_28700);
or UO_2597 (O_2597,N_29741,N_29266);
or UO_2598 (O_2598,N_29586,N_29633);
nand UO_2599 (O_2599,N_29313,N_28636);
xor UO_2600 (O_2600,N_28601,N_29585);
xnor UO_2601 (O_2601,N_29773,N_28421);
and UO_2602 (O_2602,N_29789,N_28730);
and UO_2603 (O_2603,N_29562,N_28691);
or UO_2604 (O_2604,N_28559,N_29904);
xnor UO_2605 (O_2605,N_29789,N_29043);
or UO_2606 (O_2606,N_29175,N_28943);
and UO_2607 (O_2607,N_28950,N_28345);
nand UO_2608 (O_2608,N_29410,N_29342);
nand UO_2609 (O_2609,N_28262,N_28768);
nor UO_2610 (O_2610,N_29901,N_29436);
nor UO_2611 (O_2611,N_28945,N_29410);
nand UO_2612 (O_2612,N_28221,N_28176);
xor UO_2613 (O_2613,N_29152,N_29467);
xor UO_2614 (O_2614,N_28894,N_28454);
nand UO_2615 (O_2615,N_29666,N_29056);
nor UO_2616 (O_2616,N_28010,N_29834);
and UO_2617 (O_2617,N_29293,N_29332);
or UO_2618 (O_2618,N_29314,N_29886);
nand UO_2619 (O_2619,N_28845,N_28030);
and UO_2620 (O_2620,N_28528,N_29542);
and UO_2621 (O_2621,N_28372,N_28460);
xor UO_2622 (O_2622,N_29975,N_29503);
xnor UO_2623 (O_2623,N_28832,N_28494);
and UO_2624 (O_2624,N_29402,N_29094);
nor UO_2625 (O_2625,N_29719,N_29641);
xnor UO_2626 (O_2626,N_29751,N_29330);
and UO_2627 (O_2627,N_28240,N_29144);
or UO_2628 (O_2628,N_29297,N_29812);
nor UO_2629 (O_2629,N_28095,N_29142);
and UO_2630 (O_2630,N_28000,N_29171);
nand UO_2631 (O_2631,N_29278,N_28915);
nor UO_2632 (O_2632,N_28664,N_28833);
nor UO_2633 (O_2633,N_29801,N_28807);
xnor UO_2634 (O_2634,N_28247,N_29617);
nor UO_2635 (O_2635,N_29364,N_28783);
nand UO_2636 (O_2636,N_29972,N_28457);
xnor UO_2637 (O_2637,N_29465,N_29721);
and UO_2638 (O_2638,N_29414,N_28837);
nand UO_2639 (O_2639,N_28949,N_28654);
xnor UO_2640 (O_2640,N_29664,N_28131);
xor UO_2641 (O_2641,N_29353,N_29903);
xor UO_2642 (O_2642,N_28121,N_28849);
nor UO_2643 (O_2643,N_29662,N_29732);
or UO_2644 (O_2644,N_29305,N_29384);
nor UO_2645 (O_2645,N_28767,N_29265);
nand UO_2646 (O_2646,N_29775,N_28991);
nor UO_2647 (O_2647,N_29307,N_28476);
or UO_2648 (O_2648,N_28750,N_29118);
nand UO_2649 (O_2649,N_29531,N_29613);
or UO_2650 (O_2650,N_29759,N_29264);
nor UO_2651 (O_2651,N_28077,N_28116);
and UO_2652 (O_2652,N_28104,N_29026);
nor UO_2653 (O_2653,N_29331,N_29603);
xnor UO_2654 (O_2654,N_29620,N_29585);
xor UO_2655 (O_2655,N_29896,N_28233);
nand UO_2656 (O_2656,N_29900,N_28697);
and UO_2657 (O_2657,N_28555,N_28117);
or UO_2658 (O_2658,N_28441,N_28726);
nor UO_2659 (O_2659,N_29971,N_28696);
and UO_2660 (O_2660,N_29821,N_28280);
or UO_2661 (O_2661,N_28339,N_29848);
and UO_2662 (O_2662,N_29837,N_28443);
nand UO_2663 (O_2663,N_28344,N_28030);
nand UO_2664 (O_2664,N_29043,N_29884);
nand UO_2665 (O_2665,N_29265,N_28610);
and UO_2666 (O_2666,N_29385,N_28927);
or UO_2667 (O_2667,N_28802,N_29154);
and UO_2668 (O_2668,N_28391,N_29958);
xor UO_2669 (O_2669,N_29545,N_28853);
or UO_2670 (O_2670,N_28243,N_29999);
or UO_2671 (O_2671,N_29794,N_29201);
nor UO_2672 (O_2672,N_28513,N_28018);
or UO_2673 (O_2673,N_28925,N_28488);
and UO_2674 (O_2674,N_29504,N_28366);
nor UO_2675 (O_2675,N_28116,N_29816);
and UO_2676 (O_2676,N_29253,N_29929);
and UO_2677 (O_2677,N_29971,N_29466);
xnor UO_2678 (O_2678,N_29162,N_28690);
or UO_2679 (O_2679,N_28210,N_28953);
xnor UO_2680 (O_2680,N_28684,N_29254);
or UO_2681 (O_2681,N_29629,N_28349);
nand UO_2682 (O_2682,N_28499,N_29836);
xnor UO_2683 (O_2683,N_29468,N_28391);
nor UO_2684 (O_2684,N_28051,N_28027);
nand UO_2685 (O_2685,N_29660,N_29303);
or UO_2686 (O_2686,N_29136,N_28128);
or UO_2687 (O_2687,N_29986,N_28833);
xor UO_2688 (O_2688,N_29689,N_28205);
and UO_2689 (O_2689,N_28069,N_29363);
nand UO_2690 (O_2690,N_29977,N_29325);
nand UO_2691 (O_2691,N_28106,N_29335);
nand UO_2692 (O_2692,N_29188,N_28154);
nor UO_2693 (O_2693,N_28532,N_28843);
nor UO_2694 (O_2694,N_29181,N_28885);
nor UO_2695 (O_2695,N_28216,N_29193);
and UO_2696 (O_2696,N_28092,N_29811);
and UO_2697 (O_2697,N_29912,N_28684);
or UO_2698 (O_2698,N_28094,N_29920);
xnor UO_2699 (O_2699,N_28036,N_29779);
and UO_2700 (O_2700,N_29766,N_28423);
xor UO_2701 (O_2701,N_29417,N_29436);
xnor UO_2702 (O_2702,N_28894,N_28016);
nand UO_2703 (O_2703,N_29881,N_28915);
nand UO_2704 (O_2704,N_28861,N_28125);
nand UO_2705 (O_2705,N_28886,N_29132);
xnor UO_2706 (O_2706,N_29585,N_28367);
or UO_2707 (O_2707,N_28760,N_28211);
nor UO_2708 (O_2708,N_28069,N_28343);
or UO_2709 (O_2709,N_29240,N_29646);
xor UO_2710 (O_2710,N_29893,N_28416);
and UO_2711 (O_2711,N_29418,N_28761);
and UO_2712 (O_2712,N_29605,N_28911);
and UO_2713 (O_2713,N_29801,N_28422);
and UO_2714 (O_2714,N_29754,N_28569);
xor UO_2715 (O_2715,N_29356,N_29842);
nor UO_2716 (O_2716,N_29425,N_28354);
and UO_2717 (O_2717,N_28374,N_29766);
xnor UO_2718 (O_2718,N_29492,N_29893);
nor UO_2719 (O_2719,N_29288,N_28143);
or UO_2720 (O_2720,N_29106,N_29233);
nand UO_2721 (O_2721,N_29145,N_28203);
xor UO_2722 (O_2722,N_29002,N_28193);
nand UO_2723 (O_2723,N_28281,N_28922);
nor UO_2724 (O_2724,N_28111,N_28493);
or UO_2725 (O_2725,N_29901,N_29344);
and UO_2726 (O_2726,N_28232,N_29502);
nand UO_2727 (O_2727,N_28821,N_28092);
nor UO_2728 (O_2728,N_28024,N_28388);
or UO_2729 (O_2729,N_28945,N_29625);
nor UO_2730 (O_2730,N_29171,N_28169);
and UO_2731 (O_2731,N_28241,N_28626);
nor UO_2732 (O_2732,N_28860,N_29879);
xor UO_2733 (O_2733,N_29633,N_28347);
and UO_2734 (O_2734,N_28504,N_28897);
nor UO_2735 (O_2735,N_29240,N_28177);
nand UO_2736 (O_2736,N_29068,N_29330);
xnor UO_2737 (O_2737,N_29709,N_29815);
nand UO_2738 (O_2738,N_28099,N_29101);
xnor UO_2739 (O_2739,N_29011,N_28777);
xor UO_2740 (O_2740,N_29480,N_29675);
xnor UO_2741 (O_2741,N_28149,N_28643);
and UO_2742 (O_2742,N_28804,N_28586);
xnor UO_2743 (O_2743,N_29923,N_29614);
xnor UO_2744 (O_2744,N_28273,N_28173);
xor UO_2745 (O_2745,N_29312,N_29360);
nand UO_2746 (O_2746,N_29265,N_29938);
xnor UO_2747 (O_2747,N_29544,N_29336);
xor UO_2748 (O_2748,N_28880,N_29935);
nand UO_2749 (O_2749,N_29435,N_29902);
nor UO_2750 (O_2750,N_28819,N_28468);
nand UO_2751 (O_2751,N_28714,N_29321);
nand UO_2752 (O_2752,N_29572,N_29496);
and UO_2753 (O_2753,N_28626,N_28588);
or UO_2754 (O_2754,N_29254,N_29674);
xnor UO_2755 (O_2755,N_28017,N_28841);
nor UO_2756 (O_2756,N_29685,N_29607);
nand UO_2757 (O_2757,N_28356,N_28761);
and UO_2758 (O_2758,N_29206,N_29313);
and UO_2759 (O_2759,N_29348,N_29533);
nor UO_2760 (O_2760,N_29807,N_28156);
and UO_2761 (O_2761,N_28433,N_29464);
nand UO_2762 (O_2762,N_28430,N_28699);
xnor UO_2763 (O_2763,N_28049,N_29647);
and UO_2764 (O_2764,N_29561,N_28925);
nand UO_2765 (O_2765,N_28124,N_28431);
nor UO_2766 (O_2766,N_28554,N_29288);
nor UO_2767 (O_2767,N_28513,N_28765);
nand UO_2768 (O_2768,N_29118,N_29960);
nor UO_2769 (O_2769,N_29539,N_29490);
nand UO_2770 (O_2770,N_29269,N_28461);
xnor UO_2771 (O_2771,N_28853,N_28701);
xor UO_2772 (O_2772,N_28978,N_29709);
xor UO_2773 (O_2773,N_28178,N_28848);
and UO_2774 (O_2774,N_28919,N_28556);
and UO_2775 (O_2775,N_29401,N_28253);
nor UO_2776 (O_2776,N_29354,N_29770);
or UO_2777 (O_2777,N_28398,N_29622);
nor UO_2778 (O_2778,N_29124,N_28564);
or UO_2779 (O_2779,N_29494,N_28470);
nor UO_2780 (O_2780,N_28474,N_29916);
nand UO_2781 (O_2781,N_29171,N_28390);
xnor UO_2782 (O_2782,N_29027,N_28720);
xor UO_2783 (O_2783,N_29376,N_29149);
xnor UO_2784 (O_2784,N_29221,N_29772);
nor UO_2785 (O_2785,N_29289,N_29781);
or UO_2786 (O_2786,N_28017,N_28239);
nand UO_2787 (O_2787,N_29764,N_28949);
and UO_2788 (O_2788,N_29961,N_28114);
nor UO_2789 (O_2789,N_29521,N_29887);
nand UO_2790 (O_2790,N_28333,N_29159);
and UO_2791 (O_2791,N_28180,N_29842);
xor UO_2792 (O_2792,N_28710,N_28196);
nor UO_2793 (O_2793,N_29510,N_28377);
xor UO_2794 (O_2794,N_28599,N_29181);
nor UO_2795 (O_2795,N_29535,N_29393);
or UO_2796 (O_2796,N_28682,N_29990);
nor UO_2797 (O_2797,N_29485,N_29480);
nand UO_2798 (O_2798,N_28419,N_28681);
and UO_2799 (O_2799,N_29319,N_28495);
nor UO_2800 (O_2800,N_28336,N_29450);
and UO_2801 (O_2801,N_28176,N_29146);
xor UO_2802 (O_2802,N_28294,N_29151);
or UO_2803 (O_2803,N_28135,N_29816);
or UO_2804 (O_2804,N_28836,N_29167);
nor UO_2805 (O_2805,N_28488,N_28158);
nand UO_2806 (O_2806,N_28099,N_29240);
or UO_2807 (O_2807,N_28198,N_28743);
nor UO_2808 (O_2808,N_28534,N_28130);
or UO_2809 (O_2809,N_29125,N_29293);
and UO_2810 (O_2810,N_28234,N_28605);
and UO_2811 (O_2811,N_28956,N_29227);
nor UO_2812 (O_2812,N_29910,N_29831);
and UO_2813 (O_2813,N_29231,N_29767);
nand UO_2814 (O_2814,N_28549,N_28213);
xor UO_2815 (O_2815,N_28759,N_28966);
nand UO_2816 (O_2816,N_29017,N_29627);
nand UO_2817 (O_2817,N_29357,N_28837);
nand UO_2818 (O_2818,N_29717,N_29875);
nand UO_2819 (O_2819,N_29540,N_28284);
nor UO_2820 (O_2820,N_29399,N_28864);
xor UO_2821 (O_2821,N_28964,N_28528);
and UO_2822 (O_2822,N_28203,N_29473);
nand UO_2823 (O_2823,N_28453,N_28418);
xnor UO_2824 (O_2824,N_28988,N_28389);
nand UO_2825 (O_2825,N_29970,N_29101);
nand UO_2826 (O_2826,N_28293,N_29800);
nor UO_2827 (O_2827,N_28792,N_29017);
or UO_2828 (O_2828,N_29850,N_29244);
xnor UO_2829 (O_2829,N_28985,N_28210);
xor UO_2830 (O_2830,N_29205,N_29066);
or UO_2831 (O_2831,N_29132,N_28288);
nand UO_2832 (O_2832,N_28442,N_29631);
and UO_2833 (O_2833,N_28244,N_29433);
xor UO_2834 (O_2834,N_29370,N_28877);
xor UO_2835 (O_2835,N_28355,N_29524);
nand UO_2836 (O_2836,N_28831,N_28081);
and UO_2837 (O_2837,N_28227,N_29649);
xor UO_2838 (O_2838,N_29621,N_29996);
nor UO_2839 (O_2839,N_29976,N_29438);
xnor UO_2840 (O_2840,N_28121,N_29947);
or UO_2841 (O_2841,N_29384,N_29885);
and UO_2842 (O_2842,N_29741,N_28760);
and UO_2843 (O_2843,N_29442,N_28074);
nor UO_2844 (O_2844,N_29478,N_28772);
nand UO_2845 (O_2845,N_28033,N_28067);
xnor UO_2846 (O_2846,N_28059,N_29318);
nor UO_2847 (O_2847,N_28954,N_28264);
nand UO_2848 (O_2848,N_29344,N_28152);
nor UO_2849 (O_2849,N_29524,N_28624);
or UO_2850 (O_2850,N_28224,N_28019);
nand UO_2851 (O_2851,N_28593,N_29041);
or UO_2852 (O_2852,N_29213,N_29762);
or UO_2853 (O_2853,N_28748,N_29578);
xor UO_2854 (O_2854,N_29088,N_29064);
or UO_2855 (O_2855,N_29074,N_28541);
or UO_2856 (O_2856,N_29857,N_28944);
and UO_2857 (O_2857,N_28512,N_29777);
nand UO_2858 (O_2858,N_29720,N_28807);
or UO_2859 (O_2859,N_29110,N_29908);
nor UO_2860 (O_2860,N_28285,N_29166);
nand UO_2861 (O_2861,N_29775,N_29369);
nand UO_2862 (O_2862,N_29772,N_28948);
nand UO_2863 (O_2863,N_28830,N_28077);
nor UO_2864 (O_2864,N_28013,N_29198);
and UO_2865 (O_2865,N_28946,N_29898);
xnor UO_2866 (O_2866,N_29226,N_28718);
and UO_2867 (O_2867,N_28039,N_29893);
and UO_2868 (O_2868,N_29469,N_29642);
and UO_2869 (O_2869,N_29521,N_29767);
and UO_2870 (O_2870,N_28976,N_29526);
xnor UO_2871 (O_2871,N_29408,N_29273);
nor UO_2872 (O_2872,N_29519,N_29617);
xor UO_2873 (O_2873,N_29411,N_28649);
nor UO_2874 (O_2874,N_28252,N_28529);
xor UO_2875 (O_2875,N_28645,N_28782);
xnor UO_2876 (O_2876,N_29285,N_28658);
or UO_2877 (O_2877,N_28625,N_29211);
nor UO_2878 (O_2878,N_28451,N_29322);
or UO_2879 (O_2879,N_29558,N_29798);
nor UO_2880 (O_2880,N_29402,N_28651);
nor UO_2881 (O_2881,N_29421,N_29337);
or UO_2882 (O_2882,N_29223,N_28503);
nand UO_2883 (O_2883,N_28822,N_28671);
or UO_2884 (O_2884,N_29139,N_28294);
xor UO_2885 (O_2885,N_29575,N_29609);
xor UO_2886 (O_2886,N_28608,N_28771);
xnor UO_2887 (O_2887,N_28291,N_28530);
or UO_2888 (O_2888,N_28253,N_29281);
nor UO_2889 (O_2889,N_29778,N_29985);
or UO_2890 (O_2890,N_28957,N_29032);
or UO_2891 (O_2891,N_29573,N_29058);
nand UO_2892 (O_2892,N_28455,N_29454);
nand UO_2893 (O_2893,N_29907,N_28390);
or UO_2894 (O_2894,N_28763,N_29115);
and UO_2895 (O_2895,N_28439,N_29805);
or UO_2896 (O_2896,N_28706,N_28080);
nor UO_2897 (O_2897,N_29771,N_29629);
nand UO_2898 (O_2898,N_28662,N_28093);
xor UO_2899 (O_2899,N_29467,N_29186);
and UO_2900 (O_2900,N_28234,N_28875);
and UO_2901 (O_2901,N_29549,N_29563);
nor UO_2902 (O_2902,N_29346,N_28530);
xor UO_2903 (O_2903,N_28236,N_28707);
xor UO_2904 (O_2904,N_29346,N_29842);
xor UO_2905 (O_2905,N_29817,N_29679);
or UO_2906 (O_2906,N_28605,N_28439);
and UO_2907 (O_2907,N_29648,N_29505);
or UO_2908 (O_2908,N_28372,N_29173);
or UO_2909 (O_2909,N_28889,N_28595);
nand UO_2910 (O_2910,N_29219,N_29038);
xnor UO_2911 (O_2911,N_28890,N_28755);
nand UO_2912 (O_2912,N_29035,N_28830);
and UO_2913 (O_2913,N_28733,N_28723);
and UO_2914 (O_2914,N_29050,N_28425);
xnor UO_2915 (O_2915,N_28643,N_29453);
nand UO_2916 (O_2916,N_28878,N_29195);
xor UO_2917 (O_2917,N_29825,N_29551);
nor UO_2918 (O_2918,N_28682,N_28314);
nand UO_2919 (O_2919,N_29303,N_28016);
nor UO_2920 (O_2920,N_28400,N_28529);
or UO_2921 (O_2921,N_28845,N_28302);
xor UO_2922 (O_2922,N_28454,N_28986);
nand UO_2923 (O_2923,N_29170,N_29167);
and UO_2924 (O_2924,N_29026,N_29548);
nand UO_2925 (O_2925,N_29459,N_29886);
nand UO_2926 (O_2926,N_28233,N_28389);
xnor UO_2927 (O_2927,N_28824,N_29757);
xnor UO_2928 (O_2928,N_29538,N_29778);
or UO_2929 (O_2929,N_28175,N_28100);
xor UO_2930 (O_2930,N_28265,N_29096);
and UO_2931 (O_2931,N_28565,N_29932);
nand UO_2932 (O_2932,N_29150,N_28939);
xnor UO_2933 (O_2933,N_29923,N_29473);
xor UO_2934 (O_2934,N_29262,N_29230);
or UO_2935 (O_2935,N_29709,N_29587);
and UO_2936 (O_2936,N_29382,N_29342);
nor UO_2937 (O_2937,N_29686,N_29265);
or UO_2938 (O_2938,N_29681,N_29657);
nand UO_2939 (O_2939,N_28705,N_29232);
nand UO_2940 (O_2940,N_28743,N_29873);
nand UO_2941 (O_2941,N_28493,N_28277);
or UO_2942 (O_2942,N_28477,N_28407);
or UO_2943 (O_2943,N_29278,N_28579);
and UO_2944 (O_2944,N_28047,N_28851);
nand UO_2945 (O_2945,N_29067,N_28875);
xor UO_2946 (O_2946,N_29353,N_29897);
and UO_2947 (O_2947,N_29780,N_28714);
nand UO_2948 (O_2948,N_29347,N_29657);
or UO_2949 (O_2949,N_29162,N_29486);
nand UO_2950 (O_2950,N_29236,N_29411);
xnor UO_2951 (O_2951,N_28871,N_28498);
nor UO_2952 (O_2952,N_29731,N_29975);
xnor UO_2953 (O_2953,N_29411,N_29166);
nor UO_2954 (O_2954,N_28816,N_28930);
or UO_2955 (O_2955,N_29695,N_29557);
and UO_2956 (O_2956,N_29234,N_28232);
and UO_2957 (O_2957,N_29338,N_28131);
xnor UO_2958 (O_2958,N_28687,N_29844);
and UO_2959 (O_2959,N_28735,N_29719);
nand UO_2960 (O_2960,N_28867,N_28246);
and UO_2961 (O_2961,N_29644,N_28586);
xor UO_2962 (O_2962,N_28894,N_28677);
nor UO_2963 (O_2963,N_29533,N_28667);
nor UO_2964 (O_2964,N_29542,N_29985);
nand UO_2965 (O_2965,N_29597,N_29226);
or UO_2966 (O_2966,N_29931,N_28828);
nor UO_2967 (O_2967,N_29482,N_28042);
nor UO_2968 (O_2968,N_29912,N_28847);
and UO_2969 (O_2969,N_29483,N_29818);
or UO_2970 (O_2970,N_28453,N_28049);
or UO_2971 (O_2971,N_28669,N_29230);
nand UO_2972 (O_2972,N_28718,N_29962);
xnor UO_2973 (O_2973,N_29221,N_29479);
and UO_2974 (O_2974,N_28881,N_28976);
or UO_2975 (O_2975,N_29301,N_28563);
xnor UO_2976 (O_2976,N_28123,N_29075);
and UO_2977 (O_2977,N_28904,N_29185);
xor UO_2978 (O_2978,N_29394,N_28736);
nor UO_2979 (O_2979,N_28783,N_29410);
nand UO_2980 (O_2980,N_29151,N_29356);
and UO_2981 (O_2981,N_29178,N_28659);
xnor UO_2982 (O_2982,N_28636,N_29485);
nor UO_2983 (O_2983,N_29605,N_29154);
xnor UO_2984 (O_2984,N_28606,N_29466);
or UO_2985 (O_2985,N_29617,N_28873);
xor UO_2986 (O_2986,N_29394,N_28235);
xor UO_2987 (O_2987,N_28903,N_28310);
or UO_2988 (O_2988,N_29138,N_29787);
or UO_2989 (O_2989,N_28449,N_29581);
and UO_2990 (O_2990,N_28566,N_28181);
nand UO_2991 (O_2991,N_29344,N_28472);
and UO_2992 (O_2992,N_28051,N_29279);
xor UO_2993 (O_2993,N_28342,N_28422);
and UO_2994 (O_2994,N_29452,N_29315);
or UO_2995 (O_2995,N_29624,N_28057);
xnor UO_2996 (O_2996,N_29545,N_29503);
nor UO_2997 (O_2997,N_28740,N_28769);
nor UO_2998 (O_2998,N_28293,N_28030);
and UO_2999 (O_2999,N_28734,N_29696);
xnor UO_3000 (O_3000,N_29257,N_29222);
nand UO_3001 (O_3001,N_28106,N_28864);
xor UO_3002 (O_3002,N_29487,N_28064);
nor UO_3003 (O_3003,N_29362,N_29690);
xor UO_3004 (O_3004,N_29782,N_29301);
xnor UO_3005 (O_3005,N_29528,N_29222);
nor UO_3006 (O_3006,N_29585,N_29366);
or UO_3007 (O_3007,N_28032,N_28985);
and UO_3008 (O_3008,N_28581,N_28272);
or UO_3009 (O_3009,N_29009,N_29001);
and UO_3010 (O_3010,N_29250,N_29487);
or UO_3011 (O_3011,N_28097,N_28505);
or UO_3012 (O_3012,N_29847,N_29339);
nand UO_3013 (O_3013,N_28028,N_28935);
and UO_3014 (O_3014,N_28470,N_29721);
and UO_3015 (O_3015,N_28662,N_28713);
or UO_3016 (O_3016,N_29453,N_28405);
nand UO_3017 (O_3017,N_29412,N_28113);
and UO_3018 (O_3018,N_28699,N_29201);
and UO_3019 (O_3019,N_29621,N_28818);
nand UO_3020 (O_3020,N_29564,N_29649);
and UO_3021 (O_3021,N_28562,N_29363);
nor UO_3022 (O_3022,N_28717,N_28860);
and UO_3023 (O_3023,N_29517,N_28638);
xor UO_3024 (O_3024,N_28612,N_28686);
xor UO_3025 (O_3025,N_28033,N_28004);
xnor UO_3026 (O_3026,N_29383,N_28032);
nor UO_3027 (O_3027,N_28916,N_28879);
or UO_3028 (O_3028,N_29130,N_28185);
nand UO_3029 (O_3029,N_28864,N_28920);
and UO_3030 (O_3030,N_29914,N_29431);
nand UO_3031 (O_3031,N_29735,N_29760);
xnor UO_3032 (O_3032,N_29986,N_28413);
or UO_3033 (O_3033,N_29974,N_28404);
xor UO_3034 (O_3034,N_29218,N_28314);
nand UO_3035 (O_3035,N_28748,N_29299);
xor UO_3036 (O_3036,N_28581,N_29139);
and UO_3037 (O_3037,N_29879,N_28733);
and UO_3038 (O_3038,N_28100,N_29231);
or UO_3039 (O_3039,N_28441,N_28579);
xor UO_3040 (O_3040,N_29461,N_28296);
and UO_3041 (O_3041,N_29449,N_28151);
or UO_3042 (O_3042,N_28477,N_28492);
and UO_3043 (O_3043,N_28152,N_28394);
nand UO_3044 (O_3044,N_28983,N_28452);
xor UO_3045 (O_3045,N_29278,N_29791);
and UO_3046 (O_3046,N_28376,N_29695);
or UO_3047 (O_3047,N_29660,N_28109);
nand UO_3048 (O_3048,N_29736,N_29294);
or UO_3049 (O_3049,N_29771,N_28115);
nand UO_3050 (O_3050,N_29256,N_29968);
xnor UO_3051 (O_3051,N_29455,N_28962);
or UO_3052 (O_3052,N_29170,N_28391);
nor UO_3053 (O_3053,N_29195,N_29895);
xor UO_3054 (O_3054,N_29202,N_29090);
and UO_3055 (O_3055,N_28875,N_29177);
and UO_3056 (O_3056,N_29414,N_29410);
or UO_3057 (O_3057,N_29346,N_29548);
and UO_3058 (O_3058,N_29238,N_28353);
nand UO_3059 (O_3059,N_28416,N_28006);
nor UO_3060 (O_3060,N_29638,N_28664);
and UO_3061 (O_3061,N_29819,N_28649);
and UO_3062 (O_3062,N_28537,N_28368);
or UO_3063 (O_3063,N_29417,N_29175);
xor UO_3064 (O_3064,N_28133,N_29428);
nand UO_3065 (O_3065,N_29117,N_29823);
and UO_3066 (O_3066,N_29790,N_29911);
xnor UO_3067 (O_3067,N_29080,N_28929);
and UO_3068 (O_3068,N_29658,N_29970);
and UO_3069 (O_3069,N_29888,N_29380);
nand UO_3070 (O_3070,N_29322,N_28877);
or UO_3071 (O_3071,N_29946,N_28054);
and UO_3072 (O_3072,N_29760,N_29173);
nor UO_3073 (O_3073,N_28087,N_29640);
and UO_3074 (O_3074,N_28238,N_29506);
or UO_3075 (O_3075,N_28670,N_28383);
and UO_3076 (O_3076,N_28140,N_28715);
or UO_3077 (O_3077,N_29176,N_28701);
nor UO_3078 (O_3078,N_28179,N_29981);
nand UO_3079 (O_3079,N_28659,N_28591);
and UO_3080 (O_3080,N_29313,N_29159);
xor UO_3081 (O_3081,N_29685,N_28081);
xor UO_3082 (O_3082,N_29680,N_29830);
nor UO_3083 (O_3083,N_28036,N_29781);
xor UO_3084 (O_3084,N_29020,N_28308);
nand UO_3085 (O_3085,N_28627,N_29797);
nor UO_3086 (O_3086,N_29322,N_28485);
xor UO_3087 (O_3087,N_28466,N_29694);
or UO_3088 (O_3088,N_28600,N_29164);
or UO_3089 (O_3089,N_29275,N_29799);
or UO_3090 (O_3090,N_29176,N_28128);
nand UO_3091 (O_3091,N_29390,N_29520);
nor UO_3092 (O_3092,N_29036,N_28429);
nand UO_3093 (O_3093,N_28061,N_29336);
xnor UO_3094 (O_3094,N_29603,N_29812);
xor UO_3095 (O_3095,N_29775,N_29916);
nor UO_3096 (O_3096,N_28829,N_28658);
nand UO_3097 (O_3097,N_29956,N_29153);
or UO_3098 (O_3098,N_29053,N_29796);
nor UO_3099 (O_3099,N_28229,N_29168);
or UO_3100 (O_3100,N_28050,N_28115);
xor UO_3101 (O_3101,N_29145,N_28146);
xnor UO_3102 (O_3102,N_28540,N_28864);
and UO_3103 (O_3103,N_29405,N_28421);
nor UO_3104 (O_3104,N_29918,N_29811);
nor UO_3105 (O_3105,N_29537,N_28450);
nor UO_3106 (O_3106,N_28954,N_29024);
and UO_3107 (O_3107,N_29251,N_28678);
nand UO_3108 (O_3108,N_28017,N_28996);
or UO_3109 (O_3109,N_28385,N_28499);
nand UO_3110 (O_3110,N_28871,N_28966);
nor UO_3111 (O_3111,N_29302,N_29785);
nand UO_3112 (O_3112,N_28402,N_29426);
or UO_3113 (O_3113,N_29291,N_28424);
and UO_3114 (O_3114,N_28646,N_29585);
nand UO_3115 (O_3115,N_29825,N_28313);
nand UO_3116 (O_3116,N_29406,N_28222);
nand UO_3117 (O_3117,N_28916,N_28953);
or UO_3118 (O_3118,N_29578,N_29185);
nand UO_3119 (O_3119,N_29650,N_29288);
or UO_3120 (O_3120,N_29277,N_29580);
nor UO_3121 (O_3121,N_28934,N_29530);
nand UO_3122 (O_3122,N_28039,N_29527);
or UO_3123 (O_3123,N_28091,N_28101);
xor UO_3124 (O_3124,N_28167,N_28232);
nand UO_3125 (O_3125,N_29451,N_28706);
or UO_3126 (O_3126,N_28601,N_28990);
xor UO_3127 (O_3127,N_28373,N_28885);
and UO_3128 (O_3128,N_29713,N_29924);
and UO_3129 (O_3129,N_29976,N_29085);
and UO_3130 (O_3130,N_29511,N_28363);
nand UO_3131 (O_3131,N_29099,N_29175);
nor UO_3132 (O_3132,N_29937,N_29594);
nor UO_3133 (O_3133,N_28744,N_29911);
nor UO_3134 (O_3134,N_29770,N_28164);
and UO_3135 (O_3135,N_29608,N_29709);
nor UO_3136 (O_3136,N_28712,N_28689);
nand UO_3137 (O_3137,N_28545,N_29272);
or UO_3138 (O_3138,N_29465,N_29327);
and UO_3139 (O_3139,N_28821,N_29461);
and UO_3140 (O_3140,N_28151,N_28525);
and UO_3141 (O_3141,N_29251,N_28180);
or UO_3142 (O_3142,N_29019,N_28584);
nor UO_3143 (O_3143,N_28066,N_29403);
xor UO_3144 (O_3144,N_29684,N_29151);
nor UO_3145 (O_3145,N_29920,N_28642);
xnor UO_3146 (O_3146,N_29265,N_29194);
xnor UO_3147 (O_3147,N_29377,N_28736);
xnor UO_3148 (O_3148,N_28109,N_29846);
nand UO_3149 (O_3149,N_29616,N_28940);
nand UO_3150 (O_3150,N_28211,N_28429);
nor UO_3151 (O_3151,N_28596,N_28467);
nand UO_3152 (O_3152,N_28200,N_29380);
or UO_3153 (O_3153,N_28011,N_28982);
nor UO_3154 (O_3154,N_28968,N_28070);
nand UO_3155 (O_3155,N_28276,N_28539);
and UO_3156 (O_3156,N_29486,N_29370);
xnor UO_3157 (O_3157,N_28392,N_29709);
nor UO_3158 (O_3158,N_29605,N_28569);
nand UO_3159 (O_3159,N_29078,N_28695);
nor UO_3160 (O_3160,N_29360,N_28848);
and UO_3161 (O_3161,N_29905,N_28928);
or UO_3162 (O_3162,N_28235,N_29707);
nor UO_3163 (O_3163,N_29380,N_29163);
xor UO_3164 (O_3164,N_29202,N_28091);
xnor UO_3165 (O_3165,N_29361,N_28049);
nand UO_3166 (O_3166,N_28589,N_29642);
nor UO_3167 (O_3167,N_29704,N_28034);
nor UO_3168 (O_3168,N_29463,N_28247);
and UO_3169 (O_3169,N_28567,N_28077);
nand UO_3170 (O_3170,N_28289,N_29418);
nor UO_3171 (O_3171,N_29217,N_28402);
nor UO_3172 (O_3172,N_29845,N_29121);
nor UO_3173 (O_3173,N_28045,N_29659);
nand UO_3174 (O_3174,N_29109,N_29029);
xnor UO_3175 (O_3175,N_29066,N_29402);
or UO_3176 (O_3176,N_29227,N_29324);
and UO_3177 (O_3177,N_28854,N_28985);
or UO_3178 (O_3178,N_28847,N_29880);
or UO_3179 (O_3179,N_29783,N_29545);
xor UO_3180 (O_3180,N_29215,N_28656);
or UO_3181 (O_3181,N_28826,N_28750);
xnor UO_3182 (O_3182,N_29998,N_29018);
nand UO_3183 (O_3183,N_28031,N_29395);
and UO_3184 (O_3184,N_29554,N_28986);
nor UO_3185 (O_3185,N_29473,N_29652);
or UO_3186 (O_3186,N_28001,N_28590);
xnor UO_3187 (O_3187,N_29612,N_29063);
and UO_3188 (O_3188,N_28287,N_29686);
nor UO_3189 (O_3189,N_28773,N_28451);
xor UO_3190 (O_3190,N_29974,N_28064);
nand UO_3191 (O_3191,N_29803,N_29087);
or UO_3192 (O_3192,N_28548,N_28582);
and UO_3193 (O_3193,N_28119,N_29088);
nand UO_3194 (O_3194,N_29981,N_28645);
and UO_3195 (O_3195,N_28153,N_28546);
or UO_3196 (O_3196,N_29647,N_29720);
nand UO_3197 (O_3197,N_29359,N_28205);
nand UO_3198 (O_3198,N_28047,N_29409);
or UO_3199 (O_3199,N_29724,N_28178);
nor UO_3200 (O_3200,N_29675,N_28054);
and UO_3201 (O_3201,N_29820,N_28755);
nand UO_3202 (O_3202,N_29798,N_29286);
and UO_3203 (O_3203,N_28617,N_29511);
and UO_3204 (O_3204,N_28748,N_29074);
nor UO_3205 (O_3205,N_28299,N_28690);
or UO_3206 (O_3206,N_28940,N_28406);
or UO_3207 (O_3207,N_29254,N_28172);
and UO_3208 (O_3208,N_28437,N_29330);
xnor UO_3209 (O_3209,N_29313,N_29695);
xnor UO_3210 (O_3210,N_28800,N_29798);
and UO_3211 (O_3211,N_28848,N_29092);
nand UO_3212 (O_3212,N_28230,N_29923);
and UO_3213 (O_3213,N_29385,N_29170);
nand UO_3214 (O_3214,N_28441,N_28555);
nor UO_3215 (O_3215,N_28959,N_28820);
or UO_3216 (O_3216,N_29837,N_29775);
xor UO_3217 (O_3217,N_29142,N_28121);
nand UO_3218 (O_3218,N_28186,N_29780);
nand UO_3219 (O_3219,N_29476,N_29277);
xor UO_3220 (O_3220,N_29530,N_28888);
xnor UO_3221 (O_3221,N_28596,N_28992);
nor UO_3222 (O_3222,N_28763,N_29959);
xnor UO_3223 (O_3223,N_29403,N_28866);
nand UO_3224 (O_3224,N_28245,N_29908);
or UO_3225 (O_3225,N_28641,N_29094);
xnor UO_3226 (O_3226,N_29940,N_28690);
nand UO_3227 (O_3227,N_29744,N_28420);
or UO_3228 (O_3228,N_28345,N_29207);
and UO_3229 (O_3229,N_29746,N_29134);
nand UO_3230 (O_3230,N_28259,N_28338);
and UO_3231 (O_3231,N_29504,N_28891);
or UO_3232 (O_3232,N_28412,N_28387);
xor UO_3233 (O_3233,N_28236,N_29663);
and UO_3234 (O_3234,N_28807,N_28103);
and UO_3235 (O_3235,N_29063,N_29766);
nand UO_3236 (O_3236,N_28016,N_29076);
and UO_3237 (O_3237,N_28604,N_29044);
and UO_3238 (O_3238,N_28833,N_29194);
and UO_3239 (O_3239,N_29655,N_28516);
or UO_3240 (O_3240,N_28944,N_28263);
nand UO_3241 (O_3241,N_29840,N_29272);
and UO_3242 (O_3242,N_28047,N_29934);
or UO_3243 (O_3243,N_28281,N_29649);
and UO_3244 (O_3244,N_28302,N_28102);
and UO_3245 (O_3245,N_29807,N_28567);
and UO_3246 (O_3246,N_29051,N_29314);
xnor UO_3247 (O_3247,N_29214,N_28692);
nor UO_3248 (O_3248,N_29733,N_28166);
and UO_3249 (O_3249,N_29968,N_28724);
nor UO_3250 (O_3250,N_28480,N_29594);
nand UO_3251 (O_3251,N_29431,N_28786);
xnor UO_3252 (O_3252,N_28679,N_29640);
nor UO_3253 (O_3253,N_29773,N_29480);
xnor UO_3254 (O_3254,N_29500,N_28742);
or UO_3255 (O_3255,N_29353,N_29273);
xor UO_3256 (O_3256,N_28175,N_28634);
nor UO_3257 (O_3257,N_29288,N_29680);
or UO_3258 (O_3258,N_28139,N_28514);
nor UO_3259 (O_3259,N_28858,N_28004);
nor UO_3260 (O_3260,N_28324,N_29126);
nand UO_3261 (O_3261,N_29875,N_28386);
and UO_3262 (O_3262,N_28824,N_29053);
xor UO_3263 (O_3263,N_28598,N_29851);
nor UO_3264 (O_3264,N_28435,N_28128);
and UO_3265 (O_3265,N_29062,N_28077);
and UO_3266 (O_3266,N_29966,N_29585);
or UO_3267 (O_3267,N_29121,N_29628);
nand UO_3268 (O_3268,N_29784,N_29777);
nand UO_3269 (O_3269,N_28008,N_28277);
or UO_3270 (O_3270,N_29615,N_28591);
and UO_3271 (O_3271,N_28091,N_28036);
nor UO_3272 (O_3272,N_28370,N_29227);
xnor UO_3273 (O_3273,N_28909,N_28568);
and UO_3274 (O_3274,N_29478,N_28252);
nand UO_3275 (O_3275,N_29224,N_29683);
xnor UO_3276 (O_3276,N_28192,N_28905);
nor UO_3277 (O_3277,N_28209,N_29974);
nand UO_3278 (O_3278,N_28040,N_28436);
nor UO_3279 (O_3279,N_29980,N_29029);
and UO_3280 (O_3280,N_29290,N_28575);
nand UO_3281 (O_3281,N_29384,N_28082);
nand UO_3282 (O_3282,N_29862,N_29564);
and UO_3283 (O_3283,N_28052,N_28625);
and UO_3284 (O_3284,N_29287,N_28868);
nand UO_3285 (O_3285,N_28766,N_29727);
or UO_3286 (O_3286,N_29907,N_28683);
nand UO_3287 (O_3287,N_28099,N_28940);
xnor UO_3288 (O_3288,N_28245,N_28905);
and UO_3289 (O_3289,N_29330,N_28407);
and UO_3290 (O_3290,N_28120,N_28746);
nor UO_3291 (O_3291,N_29737,N_29831);
or UO_3292 (O_3292,N_28487,N_29948);
nor UO_3293 (O_3293,N_28065,N_28892);
and UO_3294 (O_3294,N_28600,N_28969);
or UO_3295 (O_3295,N_28138,N_28098);
nor UO_3296 (O_3296,N_28805,N_29639);
nor UO_3297 (O_3297,N_29948,N_29055);
nand UO_3298 (O_3298,N_29905,N_29429);
nor UO_3299 (O_3299,N_28480,N_28275);
or UO_3300 (O_3300,N_29594,N_28075);
nor UO_3301 (O_3301,N_28344,N_28868);
or UO_3302 (O_3302,N_28165,N_28911);
xor UO_3303 (O_3303,N_29942,N_29730);
and UO_3304 (O_3304,N_28435,N_29574);
nor UO_3305 (O_3305,N_28068,N_29105);
nor UO_3306 (O_3306,N_28872,N_29462);
nor UO_3307 (O_3307,N_29335,N_28432);
xor UO_3308 (O_3308,N_28839,N_28703);
and UO_3309 (O_3309,N_28337,N_28118);
or UO_3310 (O_3310,N_28983,N_29805);
nand UO_3311 (O_3311,N_28887,N_29670);
and UO_3312 (O_3312,N_28059,N_29496);
or UO_3313 (O_3313,N_29124,N_28041);
nor UO_3314 (O_3314,N_28910,N_29714);
and UO_3315 (O_3315,N_29861,N_29934);
nor UO_3316 (O_3316,N_28729,N_29220);
and UO_3317 (O_3317,N_29923,N_29095);
and UO_3318 (O_3318,N_29629,N_29528);
nand UO_3319 (O_3319,N_29302,N_28295);
and UO_3320 (O_3320,N_28978,N_28592);
and UO_3321 (O_3321,N_29566,N_28751);
and UO_3322 (O_3322,N_28992,N_29490);
nand UO_3323 (O_3323,N_28288,N_29354);
or UO_3324 (O_3324,N_28808,N_28977);
xor UO_3325 (O_3325,N_28444,N_29430);
nand UO_3326 (O_3326,N_29510,N_28448);
nand UO_3327 (O_3327,N_29854,N_28866);
and UO_3328 (O_3328,N_29183,N_28277);
nand UO_3329 (O_3329,N_28253,N_29055);
xnor UO_3330 (O_3330,N_29106,N_29876);
or UO_3331 (O_3331,N_28088,N_28690);
nor UO_3332 (O_3332,N_29605,N_29887);
and UO_3333 (O_3333,N_29568,N_29611);
or UO_3334 (O_3334,N_29920,N_29287);
and UO_3335 (O_3335,N_28247,N_29142);
or UO_3336 (O_3336,N_28175,N_28344);
xnor UO_3337 (O_3337,N_28730,N_29302);
xor UO_3338 (O_3338,N_28949,N_29747);
nor UO_3339 (O_3339,N_29821,N_28262);
or UO_3340 (O_3340,N_29284,N_28743);
or UO_3341 (O_3341,N_28938,N_29233);
and UO_3342 (O_3342,N_29885,N_29866);
or UO_3343 (O_3343,N_29263,N_28794);
or UO_3344 (O_3344,N_28295,N_29585);
xor UO_3345 (O_3345,N_29931,N_29483);
or UO_3346 (O_3346,N_29644,N_28528);
and UO_3347 (O_3347,N_28815,N_29225);
nor UO_3348 (O_3348,N_29286,N_28797);
or UO_3349 (O_3349,N_29854,N_28136);
nand UO_3350 (O_3350,N_29050,N_29646);
nor UO_3351 (O_3351,N_28966,N_28818);
or UO_3352 (O_3352,N_29004,N_28049);
and UO_3353 (O_3353,N_28357,N_28523);
nand UO_3354 (O_3354,N_29102,N_28892);
nand UO_3355 (O_3355,N_29581,N_28544);
or UO_3356 (O_3356,N_29719,N_29639);
or UO_3357 (O_3357,N_28387,N_28853);
and UO_3358 (O_3358,N_28246,N_29995);
nor UO_3359 (O_3359,N_28006,N_29156);
nor UO_3360 (O_3360,N_29589,N_28598);
nor UO_3361 (O_3361,N_28985,N_29311);
and UO_3362 (O_3362,N_29366,N_29175);
nand UO_3363 (O_3363,N_28710,N_29934);
or UO_3364 (O_3364,N_28001,N_28366);
xor UO_3365 (O_3365,N_29801,N_28887);
or UO_3366 (O_3366,N_28211,N_28305);
nand UO_3367 (O_3367,N_29055,N_28601);
and UO_3368 (O_3368,N_28847,N_29372);
and UO_3369 (O_3369,N_28666,N_28180);
xnor UO_3370 (O_3370,N_28029,N_28230);
nor UO_3371 (O_3371,N_29285,N_29077);
nor UO_3372 (O_3372,N_28048,N_28366);
xor UO_3373 (O_3373,N_28397,N_29916);
and UO_3374 (O_3374,N_28731,N_29021);
and UO_3375 (O_3375,N_28656,N_28795);
and UO_3376 (O_3376,N_28218,N_28338);
xor UO_3377 (O_3377,N_28533,N_28777);
or UO_3378 (O_3378,N_28477,N_29220);
or UO_3379 (O_3379,N_29158,N_28852);
nor UO_3380 (O_3380,N_29363,N_28232);
or UO_3381 (O_3381,N_28863,N_28103);
and UO_3382 (O_3382,N_29586,N_29159);
or UO_3383 (O_3383,N_28449,N_29657);
or UO_3384 (O_3384,N_28410,N_29138);
and UO_3385 (O_3385,N_28091,N_29342);
xnor UO_3386 (O_3386,N_28608,N_28057);
or UO_3387 (O_3387,N_28185,N_29559);
nor UO_3388 (O_3388,N_29866,N_28202);
or UO_3389 (O_3389,N_28236,N_29045);
nand UO_3390 (O_3390,N_28819,N_29733);
and UO_3391 (O_3391,N_29059,N_29039);
and UO_3392 (O_3392,N_29707,N_29167);
nand UO_3393 (O_3393,N_29067,N_28043);
or UO_3394 (O_3394,N_28984,N_29022);
or UO_3395 (O_3395,N_28218,N_29419);
xnor UO_3396 (O_3396,N_29913,N_29302);
or UO_3397 (O_3397,N_28229,N_29551);
nor UO_3398 (O_3398,N_29004,N_29841);
nor UO_3399 (O_3399,N_29632,N_29495);
xor UO_3400 (O_3400,N_28553,N_28382);
or UO_3401 (O_3401,N_29147,N_29862);
nand UO_3402 (O_3402,N_29920,N_29490);
and UO_3403 (O_3403,N_28913,N_28704);
xnor UO_3404 (O_3404,N_29868,N_29371);
nor UO_3405 (O_3405,N_28320,N_28625);
xor UO_3406 (O_3406,N_29327,N_29146);
xor UO_3407 (O_3407,N_29311,N_29629);
or UO_3408 (O_3408,N_28484,N_29815);
and UO_3409 (O_3409,N_29579,N_28274);
or UO_3410 (O_3410,N_28523,N_29557);
nand UO_3411 (O_3411,N_29239,N_28837);
or UO_3412 (O_3412,N_29668,N_28156);
nand UO_3413 (O_3413,N_29102,N_28210);
or UO_3414 (O_3414,N_29829,N_29586);
or UO_3415 (O_3415,N_29046,N_28016);
nor UO_3416 (O_3416,N_29558,N_28583);
or UO_3417 (O_3417,N_29973,N_28203);
nor UO_3418 (O_3418,N_28793,N_28135);
nand UO_3419 (O_3419,N_29439,N_29862);
xnor UO_3420 (O_3420,N_29491,N_29974);
xnor UO_3421 (O_3421,N_28191,N_28513);
or UO_3422 (O_3422,N_28023,N_29929);
xnor UO_3423 (O_3423,N_29003,N_29747);
and UO_3424 (O_3424,N_29347,N_28927);
or UO_3425 (O_3425,N_29987,N_28727);
and UO_3426 (O_3426,N_29201,N_28687);
nand UO_3427 (O_3427,N_29361,N_28072);
nand UO_3428 (O_3428,N_29293,N_29010);
nand UO_3429 (O_3429,N_28290,N_28841);
or UO_3430 (O_3430,N_29888,N_29436);
nand UO_3431 (O_3431,N_29163,N_28655);
and UO_3432 (O_3432,N_28000,N_29831);
or UO_3433 (O_3433,N_28210,N_29459);
and UO_3434 (O_3434,N_28548,N_28866);
nor UO_3435 (O_3435,N_29594,N_29020);
xor UO_3436 (O_3436,N_29660,N_29361);
and UO_3437 (O_3437,N_28695,N_28095);
and UO_3438 (O_3438,N_28653,N_28076);
or UO_3439 (O_3439,N_29818,N_28409);
and UO_3440 (O_3440,N_28855,N_28397);
xnor UO_3441 (O_3441,N_28302,N_28063);
or UO_3442 (O_3442,N_28561,N_28486);
xnor UO_3443 (O_3443,N_28763,N_28377);
nor UO_3444 (O_3444,N_28072,N_28119);
nor UO_3445 (O_3445,N_29343,N_28175);
nor UO_3446 (O_3446,N_29866,N_28829);
nor UO_3447 (O_3447,N_28072,N_28222);
or UO_3448 (O_3448,N_29117,N_28599);
nand UO_3449 (O_3449,N_29925,N_28950);
nand UO_3450 (O_3450,N_28798,N_29594);
or UO_3451 (O_3451,N_29910,N_28742);
nor UO_3452 (O_3452,N_29100,N_28948);
nor UO_3453 (O_3453,N_29124,N_28655);
xnor UO_3454 (O_3454,N_28837,N_29872);
or UO_3455 (O_3455,N_28371,N_28181);
nand UO_3456 (O_3456,N_29531,N_29803);
and UO_3457 (O_3457,N_28193,N_28521);
xnor UO_3458 (O_3458,N_29575,N_28476);
or UO_3459 (O_3459,N_28943,N_29560);
xor UO_3460 (O_3460,N_28823,N_28267);
or UO_3461 (O_3461,N_29860,N_28891);
xnor UO_3462 (O_3462,N_29842,N_29890);
xnor UO_3463 (O_3463,N_29969,N_29062);
and UO_3464 (O_3464,N_28800,N_29795);
nor UO_3465 (O_3465,N_29637,N_29620);
nand UO_3466 (O_3466,N_28240,N_29863);
and UO_3467 (O_3467,N_28766,N_29914);
nor UO_3468 (O_3468,N_28012,N_29146);
nor UO_3469 (O_3469,N_28738,N_28592);
nand UO_3470 (O_3470,N_29647,N_29027);
nand UO_3471 (O_3471,N_28300,N_29107);
or UO_3472 (O_3472,N_28755,N_29298);
nand UO_3473 (O_3473,N_29018,N_29914);
xor UO_3474 (O_3474,N_29223,N_28499);
nand UO_3475 (O_3475,N_28470,N_29613);
nand UO_3476 (O_3476,N_28651,N_29190);
nand UO_3477 (O_3477,N_28844,N_28862);
nand UO_3478 (O_3478,N_28161,N_29872);
nor UO_3479 (O_3479,N_29278,N_29012);
or UO_3480 (O_3480,N_28408,N_29379);
xnor UO_3481 (O_3481,N_28162,N_29702);
xnor UO_3482 (O_3482,N_28456,N_28752);
or UO_3483 (O_3483,N_29520,N_28464);
nor UO_3484 (O_3484,N_28885,N_29436);
nor UO_3485 (O_3485,N_28303,N_29652);
nand UO_3486 (O_3486,N_28994,N_28517);
nor UO_3487 (O_3487,N_29861,N_29849);
nand UO_3488 (O_3488,N_29324,N_29620);
nand UO_3489 (O_3489,N_28353,N_28399);
and UO_3490 (O_3490,N_28582,N_29931);
xor UO_3491 (O_3491,N_28879,N_28661);
and UO_3492 (O_3492,N_29573,N_28591);
or UO_3493 (O_3493,N_29971,N_28996);
xnor UO_3494 (O_3494,N_29711,N_28313);
xor UO_3495 (O_3495,N_28281,N_28546);
and UO_3496 (O_3496,N_29970,N_28992);
nor UO_3497 (O_3497,N_29419,N_29278);
or UO_3498 (O_3498,N_28281,N_28766);
or UO_3499 (O_3499,N_28101,N_28996);
endmodule