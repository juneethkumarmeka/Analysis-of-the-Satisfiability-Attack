module basic_500_3000_500_40_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_184,In_473);
nand U1 (N_1,In_108,In_393);
xor U2 (N_2,In_496,In_140);
nand U3 (N_3,In_495,In_361);
and U4 (N_4,In_106,In_251);
nor U5 (N_5,In_456,In_157);
nor U6 (N_6,In_176,In_490);
nand U7 (N_7,In_263,In_50);
or U8 (N_8,In_291,In_446);
or U9 (N_9,In_238,In_457);
and U10 (N_10,In_36,In_289);
and U11 (N_11,In_143,In_156);
xnor U12 (N_12,In_237,In_25);
and U13 (N_13,In_137,In_0);
xnor U14 (N_14,In_196,In_217);
nor U15 (N_15,In_380,In_312);
and U16 (N_16,In_61,In_135);
xor U17 (N_17,In_459,In_266);
xnor U18 (N_18,In_410,In_252);
and U19 (N_19,In_134,In_429);
or U20 (N_20,In_494,In_62);
xor U21 (N_21,In_353,In_453);
nand U22 (N_22,In_293,In_51);
nand U23 (N_23,In_439,In_345);
nor U24 (N_24,In_164,In_259);
or U25 (N_25,In_323,In_275);
or U26 (N_26,In_357,In_466);
and U27 (N_27,In_15,In_442);
or U28 (N_28,In_484,In_414);
xor U29 (N_29,In_138,In_209);
xnor U30 (N_30,In_16,In_454);
nor U31 (N_31,In_285,In_400);
xnor U32 (N_32,In_306,In_317);
xor U33 (N_33,In_445,In_94);
nor U34 (N_34,In_341,In_194);
nand U35 (N_35,In_347,In_120);
or U36 (N_36,In_255,In_449);
nor U37 (N_37,In_458,In_472);
or U38 (N_38,In_423,In_95);
xnor U39 (N_39,In_253,In_249);
nor U40 (N_40,In_428,In_364);
nand U41 (N_41,In_72,In_450);
nand U42 (N_42,In_272,In_425);
or U43 (N_43,In_235,In_435);
and U44 (N_44,In_205,In_152);
and U45 (N_45,In_204,In_60);
nor U46 (N_46,In_427,In_45);
xnor U47 (N_47,In_112,In_91);
nor U48 (N_48,In_100,In_127);
nand U49 (N_49,In_354,In_87);
and U50 (N_50,In_225,In_111);
xnor U51 (N_51,In_226,In_298);
xor U52 (N_52,In_296,In_227);
nand U53 (N_53,In_288,In_322);
nor U54 (N_54,In_367,In_417);
nand U55 (N_55,In_5,In_232);
nor U56 (N_56,In_114,In_228);
nor U57 (N_57,In_346,In_394);
and U58 (N_58,In_316,In_113);
and U59 (N_59,In_59,In_444);
xor U60 (N_60,In_131,In_158);
xor U61 (N_61,In_183,In_142);
nor U62 (N_62,In_460,In_250);
or U63 (N_63,In_186,In_40);
nand U64 (N_64,In_280,In_124);
or U65 (N_65,In_362,In_396);
or U66 (N_66,In_290,In_461);
or U67 (N_67,In_391,In_282);
nand U68 (N_68,In_213,In_177);
nand U69 (N_69,In_214,In_486);
xor U70 (N_70,In_485,In_30);
nand U71 (N_71,In_96,In_265);
xnor U72 (N_72,In_474,In_93);
nor U73 (N_73,In_21,In_154);
xnor U74 (N_74,In_125,In_413);
xor U75 (N_75,In_337,In_54);
nand U76 (N_76,N_32,In_27);
or U77 (N_77,In_167,N_30);
or U78 (N_78,In_338,In_198);
and U79 (N_79,In_271,In_151);
nand U80 (N_80,N_33,In_448);
xor U81 (N_81,N_31,In_348);
or U82 (N_82,In_351,In_58);
xor U83 (N_83,In_181,In_18);
and U84 (N_84,In_203,In_80);
nor U85 (N_85,In_32,In_97);
or U86 (N_86,In_144,In_231);
or U87 (N_87,In_133,In_452);
xor U88 (N_88,In_479,In_173);
nor U89 (N_89,In_355,In_487);
nand U90 (N_90,In_22,In_482);
xnor U91 (N_91,In_104,In_305);
and U92 (N_92,In_371,N_4);
or U93 (N_93,In_401,In_150);
xor U94 (N_94,In_169,In_79);
and U95 (N_95,In_23,In_294);
or U96 (N_96,In_76,In_276);
or U97 (N_97,N_46,In_162);
nor U98 (N_98,In_398,In_7);
and U99 (N_99,N_19,In_418);
and U100 (N_100,In_307,In_382);
xor U101 (N_101,In_246,In_116);
or U102 (N_102,N_61,In_287);
and U103 (N_103,In_292,In_369);
and U104 (N_104,In_360,N_0);
or U105 (N_105,In_363,In_122);
xnor U106 (N_106,In_223,In_78);
xnor U107 (N_107,N_62,In_202);
nand U108 (N_108,In_356,N_43);
xnor U109 (N_109,In_390,N_22);
and U110 (N_110,N_12,In_170);
xnor U111 (N_111,In_70,In_118);
or U112 (N_112,N_63,In_9);
nor U113 (N_113,In_119,In_310);
or U114 (N_114,N_47,N_18);
nor U115 (N_115,In_2,N_21);
or U116 (N_116,In_103,In_221);
nand U117 (N_117,N_64,In_53);
nand U118 (N_118,N_45,In_342);
and U119 (N_119,In_26,In_75);
nor U120 (N_120,In_77,In_208);
xnor U121 (N_121,In_86,In_408);
nor U122 (N_122,In_179,In_159);
xor U123 (N_123,In_303,In_437);
xnor U124 (N_124,In_480,N_70);
and U125 (N_125,In_281,In_180);
nand U126 (N_126,In_340,In_172);
nand U127 (N_127,In_300,In_239);
or U128 (N_128,In_405,In_318);
nor U129 (N_129,In_493,In_476);
and U130 (N_130,In_182,In_433);
xnor U131 (N_131,In_412,In_199);
and U132 (N_132,In_46,In_477);
xor U133 (N_133,N_23,In_229);
nor U134 (N_134,In_419,In_42);
nor U135 (N_135,In_234,In_14);
nand U136 (N_136,In_243,In_430);
or U137 (N_137,In_497,In_329);
nand U138 (N_138,In_222,In_483);
nor U139 (N_139,N_40,In_155);
or U140 (N_140,In_244,In_43);
xor U141 (N_141,N_13,N_24);
nand U142 (N_142,In_69,In_426);
and U143 (N_143,In_399,In_431);
or U144 (N_144,In_17,N_9);
nor U145 (N_145,In_161,In_163);
nor U146 (N_146,In_406,In_376);
xor U147 (N_147,In_19,In_185);
and U148 (N_148,In_421,In_37);
xor U149 (N_149,In_440,N_72);
and U150 (N_150,In_189,In_447);
nand U151 (N_151,In_270,In_311);
xor U152 (N_152,N_121,In_286);
or U153 (N_153,N_66,N_88);
and U154 (N_154,In_4,N_59);
and U155 (N_155,In_416,N_44);
nor U156 (N_156,N_11,N_16);
xor U157 (N_157,In_302,N_48);
xnor U158 (N_158,In_279,In_304);
nor U159 (N_159,In_105,In_402);
or U160 (N_160,In_471,N_110);
nor U161 (N_161,In_465,In_492);
and U162 (N_162,In_409,In_90);
or U163 (N_163,In_384,N_112);
or U164 (N_164,In_333,In_3);
nor U165 (N_165,In_381,N_130);
and U166 (N_166,In_57,N_39);
nor U167 (N_167,In_468,In_236);
nor U168 (N_168,In_88,In_278);
nand U169 (N_169,In_260,In_139);
or U170 (N_170,In_10,N_128);
and U171 (N_171,In_295,N_97);
nand U172 (N_172,In_191,In_257);
nor U173 (N_173,In_13,N_120);
nor U174 (N_174,In_136,In_462);
or U175 (N_175,In_219,N_139);
nand U176 (N_176,In_241,N_94);
nand U177 (N_177,N_50,N_73);
or U178 (N_178,N_3,N_106);
nand U179 (N_179,In_284,N_10);
nor U180 (N_180,N_101,In_377);
and U181 (N_181,In_478,In_123);
nor U182 (N_182,N_140,In_464);
or U183 (N_183,In_350,In_349);
and U184 (N_184,In_455,N_116);
or U185 (N_185,N_99,N_92);
xor U186 (N_186,In_85,In_370);
and U187 (N_187,In_110,In_212);
nand U188 (N_188,In_68,N_68);
or U189 (N_189,N_145,In_147);
and U190 (N_190,In_245,In_379);
nand U191 (N_191,N_25,N_76);
or U192 (N_192,In_24,In_215);
and U193 (N_193,In_321,N_6);
nor U194 (N_194,In_6,In_210);
nor U195 (N_195,N_29,N_2);
nor U196 (N_196,N_34,In_153);
nand U197 (N_197,In_301,In_368);
nor U198 (N_198,In_331,In_359);
xor U199 (N_199,In_463,In_207);
or U200 (N_200,In_488,N_91);
or U201 (N_201,In_499,In_89);
xnor U202 (N_202,In_82,In_395);
or U203 (N_203,In_262,N_102);
or U204 (N_204,In_192,N_80);
nor U205 (N_205,In_451,In_48);
or U206 (N_206,In_432,In_107);
or U207 (N_207,In_375,In_308);
nand U208 (N_208,N_105,N_118);
nand U209 (N_209,In_166,N_82);
nand U210 (N_210,In_274,In_28);
nand U211 (N_211,In_187,In_66);
or U212 (N_212,N_111,In_404);
xnor U213 (N_213,In_411,In_8);
nand U214 (N_214,In_470,In_240);
and U215 (N_215,In_128,In_130);
nor U216 (N_216,N_149,N_131);
nor U217 (N_217,N_83,N_85);
or U218 (N_218,N_37,N_28);
and U219 (N_219,In_247,In_267);
nor U220 (N_220,In_386,In_332);
nor U221 (N_221,In_160,In_39);
nand U222 (N_222,N_69,N_60);
or U223 (N_223,In_92,In_314);
xor U224 (N_224,In_268,In_63);
nand U225 (N_225,In_44,N_79);
nand U226 (N_226,N_36,In_126);
xor U227 (N_227,N_98,N_223);
xnor U228 (N_228,In_81,In_335);
nand U229 (N_229,In_220,N_202);
nor U230 (N_230,N_216,In_211);
nor U231 (N_231,In_12,N_123);
and U232 (N_232,N_188,N_218);
xor U233 (N_233,N_65,N_57);
nor U234 (N_234,N_208,In_197);
and U235 (N_235,N_194,In_101);
or U236 (N_236,N_191,In_269);
xor U237 (N_237,N_162,In_84);
and U238 (N_238,In_344,In_334);
nor U239 (N_239,In_174,N_56);
and U240 (N_240,N_221,N_200);
xor U241 (N_241,N_171,In_343);
nor U242 (N_242,In_374,N_164);
or U243 (N_243,In_438,N_178);
or U244 (N_244,N_143,In_20);
nor U245 (N_245,N_124,N_174);
nand U246 (N_246,N_169,In_168);
nand U247 (N_247,In_264,In_195);
nand U248 (N_248,In_149,In_98);
nand U249 (N_249,N_86,In_178);
nand U250 (N_250,N_129,N_206);
xor U251 (N_251,In_141,In_277);
and U252 (N_252,N_193,N_75);
xnor U253 (N_253,N_8,N_132);
and U254 (N_254,N_136,N_224);
xnor U255 (N_255,N_156,In_171);
or U256 (N_256,In_358,In_372);
nand U257 (N_257,N_209,N_210);
nor U258 (N_258,N_41,N_157);
and U259 (N_259,N_219,In_261);
nand U260 (N_260,N_93,N_152);
nor U261 (N_261,In_441,N_217);
nor U262 (N_262,In_224,N_58);
and U263 (N_263,N_212,In_145);
nor U264 (N_264,N_1,In_469);
xnor U265 (N_265,In_83,In_313);
nor U266 (N_266,N_142,N_182);
nor U267 (N_267,N_154,N_187);
and U268 (N_268,In_188,In_385);
xor U269 (N_269,In_216,N_213);
nand U270 (N_270,N_204,N_155);
nand U271 (N_271,N_5,N_192);
nand U272 (N_272,In_467,N_141);
xnor U273 (N_273,In_193,In_190);
nor U274 (N_274,In_248,N_179);
nor U275 (N_275,In_387,N_144);
and U276 (N_276,N_185,In_498);
xor U277 (N_277,In_422,N_220);
and U278 (N_278,N_148,N_189);
or U279 (N_279,N_53,N_205);
xor U280 (N_280,N_215,N_49);
and U281 (N_281,In_132,N_15);
and U282 (N_282,In_55,N_51);
nand U283 (N_283,N_67,In_242);
nor U284 (N_284,In_35,N_197);
xnor U285 (N_285,In_254,N_81);
nor U286 (N_286,N_89,In_129);
nand U287 (N_287,N_125,N_96);
nand U288 (N_288,N_180,In_99);
xor U289 (N_289,In_1,In_33);
xnor U290 (N_290,In_415,In_424);
nand U291 (N_291,N_17,N_104);
or U292 (N_292,In_383,In_339);
nand U293 (N_293,N_138,In_392);
nor U294 (N_294,N_20,N_151);
nand U295 (N_295,In_327,In_201);
and U296 (N_296,N_201,N_163);
nand U297 (N_297,N_84,N_168);
xnor U298 (N_298,In_71,In_299);
xnor U299 (N_299,N_107,N_195);
nand U300 (N_300,N_26,N_77);
nor U301 (N_301,N_260,In_38);
nor U302 (N_302,N_263,In_397);
and U303 (N_303,N_159,In_336);
and U304 (N_304,N_279,In_436);
nor U305 (N_305,In_256,N_74);
and U306 (N_306,N_183,N_114);
or U307 (N_307,N_266,N_250);
and U308 (N_308,In_320,N_113);
or U309 (N_309,N_255,In_491);
xor U310 (N_310,N_265,N_291);
nor U311 (N_311,N_115,In_315);
and U312 (N_312,N_172,In_73);
nand U313 (N_313,In_11,N_90);
xor U314 (N_314,In_330,In_273);
nor U315 (N_315,In_165,In_373);
nand U316 (N_316,N_242,N_160);
or U317 (N_317,N_87,N_277);
or U318 (N_318,In_175,In_67);
xnor U319 (N_319,N_167,N_283);
nand U320 (N_320,N_256,N_233);
xor U321 (N_321,N_273,In_146);
nand U322 (N_322,N_235,N_274);
xor U323 (N_323,N_137,In_109);
xor U324 (N_324,N_246,N_199);
nand U325 (N_325,N_231,In_200);
xor U326 (N_326,N_190,N_78);
or U327 (N_327,N_252,In_309);
xor U328 (N_328,In_49,N_281);
and U329 (N_329,N_292,In_297);
and U330 (N_330,N_103,In_407);
and U331 (N_331,N_122,N_14);
xor U332 (N_332,N_236,N_146);
or U333 (N_333,N_245,N_176);
or U334 (N_334,In_378,N_285);
or U335 (N_335,N_166,In_403);
nand U336 (N_336,N_153,N_158);
or U337 (N_337,N_177,N_109);
nor U338 (N_338,N_150,N_214);
nand U339 (N_339,In_52,In_31);
xnor U340 (N_340,N_243,N_95);
and U341 (N_341,N_267,N_55);
nand U342 (N_342,N_249,N_257);
xor U343 (N_343,In_481,N_133);
nand U344 (N_344,In_388,N_230);
xnor U345 (N_345,N_240,N_184);
or U346 (N_346,N_244,N_226);
and U347 (N_347,In_352,N_241);
and U348 (N_348,In_206,In_65);
xnor U349 (N_349,In_148,In_74);
or U350 (N_350,N_282,N_264);
nor U351 (N_351,N_181,In_230);
and U352 (N_352,N_299,N_254);
and U353 (N_353,In_47,In_258);
and U354 (N_354,In_389,N_54);
nand U355 (N_355,N_165,In_328);
or U356 (N_356,N_275,N_258);
xnor U357 (N_357,In_56,N_7);
nor U358 (N_358,N_211,In_117);
and U359 (N_359,In_41,In_443);
nand U360 (N_360,N_127,N_261);
or U361 (N_361,N_297,In_218);
and U362 (N_362,N_237,N_290);
or U363 (N_363,N_71,N_248);
nor U364 (N_364,In_121,N_287);
or U365 (N_365,N_251,N_289);
xnor U366 (N_366,N_284,N_253);
xnor U367 (N_367,N_295,N_203);
nand U368 (N_368,N_135,In_233);
xnor U369 (N_369,N_52,In_29);
nor U370 (N_370,In_102,N_298);
and U371 (N_371,N_207,N_126);
nand U372 (N_372,In_489,In_324);
and U373 (N_373,In_326,N_247);
nor U374 (N_374,In_34,In_115);
or U375 (N_375,N_350,N_301);
nand U376 (N_376,N_286,N_198);
or U377 (N_377,N_311,N_344);
nor U378 (N_378,N_370,N_359);
or U379 (N_379,N_368,N_331);
xor U380 (N_380,N_27,N_269);
nand U381 (N_381,N_304,N_315);
nand U382 (N_382,N_355,N_272);
and U383 (N_383,N_314,N_334);
and U384 (N_384,N_307,N_372);
nor U385 (N_385,N_371,N_300);
nand U386 (N_386,In_475,N_323);
xor U387 (N_387,N_318,N_108);
or U388 (N_388,N_280,N_225);
or U389 (N_389,N_321,N_336);
nor U390 (N_390,N_134,N_349);
and U391 (N_391,N_271,N_351);
and U392 (N_392,N_222,N_313);
or U393 (N_393,N_234,N_306);
nor U394 (N_394,N_262,N_329);
nor U395 (N_395,In_325,In_366);
nand U396 (N_396,N_325,N_347);
nand U397 (N_397,N_348,N_317);
or U398 (N_398,N_276,In_283);
xnor U399 (N_399,N_360,N_316);
nor U400 (N_400,N_322,N_38);
and U401 (N_401,N_353,N_305);
xnor U402 (N_402,N_337,N_228);
nor U403 (N_403,N_346,N_361);
or U404 (N_404,N_294,N_296);
or U405 (N_405,N_328,N_293);
xor U406 (N_406,N_100,N_342);
nor U407 (N_407,N_335,N_175);
xor U408 (N_408,N_268,N_365);
nor U409 (N_409,N_324,N_338);
nand U410 (N_410,N_330,N_367);
nor U411 (N_411,N_278,N_354);
xnor U412 (N_412,N_362,N_186);
nand U413 (N_413,N_333,N_227);
nand U414 (N_414,N_343,N_356);
xor U415 (N_415,In_64,N_173);
nor U416 (N_416,N_320,In_420);
xnor U417 (N_417,N_119,N_312);
nand U418 (N_418,N_147,N_341);
nand U419 (N_419,N_326,N_345);
and U420 (N_420,In_434,In_365);
or U421 (N_421,N_373,N_332);
xor U422 (N_422,In_319,N_364);
nand U423 (N_423,N_358,N_239);
nand U424 (N_424,N_259,N_232);
nand U425 (N_425,N_270,N_303);
xnor U426 (N_426,N_170,N_366);
xnor U427 (N_427,N_238,N_352);
nor U428 (N_428,N_340,N_310);
nand U429 (N_429,N_374,N_363);
xnor U430 (N_430,N_288,N_229);
nor U431 (N_431,N_369,N_42);
xor U432 (N_432,N_339,N_196);
and U433 (N_433,N_319,N_309);
and U434 (N_434,N_308,N_117);
xor U435 (N_435,N_161,N_357);
nand U436 (N_436,N_327,N_35);
nand U437 (N_437,N_302,N_276);
xor U438 (N_438,N_268,N_353);
nor U439 (N_439,N_309,N_294);
and U440 (N_440,N_234,N_339);
xnor U441 (N_441,N_339,N_349);
nor U442 (N_442,N_355,In_420);
and U443 (N_443,N_329,N_269);
and U444 (N_444,N_227,N_347);
nor U445 (N_445,N_280,N_198);
nand U446 (N_446,N_373,N_315);
nand U447 (N_447,N_366,N_334);
nand U448 (N_448,N_306,N_333);
nor U449 (N_449,N_352,N_278);
nand U450 (N_450,N_436,N_393);
nor U451 (N_451,N_378,N_432);
nor U452 (N_452,N_404,N_385);
nand U453 (N_453,N_396,N_403);
xnor U454 (N_454,N_415,N_388);
and U455 (N_455,N_375,N_442);
nand U456 (N_456,N_382,N_447);
nand U457 (N_457,N_410,N_377);
or U458 (N_458,N_427,N_376);
xor U459 (N_459,N_420,N_423);
or U460 (N_460,N_398,N_424);
and U461 (N_461,N_389,N_417);
nand U462 (N_462,N_414,N_387);
nor U463 (N_463,N_446,N_445);
xor U464 (N_464,N_433,N_448);
nor U465 (N_465,N_431,N_379);
or U466 (N_466,N_430,N_407);
nand U467 (N_467,N_399,N_419);
xor U468 (N_468,N_441,N_438);
nand U469 (N_469,N_402,N_406);
nand U470 (N_470,N_386,N_443);
or U471 (N_471,N_412,N_428);
nand U472 (N_472,N_392,N_444);
or U473 (N_473,N_437,N_405);
or U474 (N_474,N_426,N_384);
or U475 (N_475,N_413,N_418);
nand U476 (N_476,N_408,N_401);
nand U477 (N_477,N_429,N_395);
and U478 (N_478,N_397,N_391);
nor U479 (N_479,N_411,N_416);
nor U480 (N_480,N_421,N_390);
nand U481 (N_481,N_394,N_435);
and U482 (N_482,N_434,N_449);
nand U483 (N_483,N_381,N_400);
nand U484 (N_484,N_439,N_380);
and U485 (N_485,N_425,N_409);
nand U486 (N_486,N_422,N_383);
xor U487 (N_487,N_440,N_434);
and U488 (N_488,N_440,N_429);
nand U489 (N_489,N_416,N_428);
nor U490 (N_490,N_409,N_413);
nor U491 (N_491,N_387,N_443);
nand U492 (N_492,N_433,N_443);
nor U493 (N_493,N_378,N_442);
and U494 (N_494,N_402,N_423);
nand U495 (N_495,N_427,N_441);
xnor U496 (N_496,N_448,N_389);
xnor U497 (N_497,N_442,N_399);
nand U498 (N_498,N_427,N_375);
nor U499 (N_499,N_426,N_405);
or U500 (N_500,N_408,N_441);
xnor U501 (N_501,N_438,N_379);
nand U502 (N_502,N_386,N_408);
or U503 (N_503,N_405,N_429);
and U504 (N_504,N_434,N_386);
xor U505 (N_505,N_445,N_392);
xor U506 (N_506,N_429,N_403);
or U507 (N_507,N_436,N_386);
nor U508 (N_508,N_421,N_379);
nand U509 (N_509,N_387,N_386);
or U510 (N_510,N_449,N_412);
and U511 (N_511,N_394,N_418);
or U512 (N_512,N_433,N_375);
nor U513 (N_513,N_385,N_431);
xor U514 (N_514,N_378,N_390);
and U515 (N_515,N_445,N_380);
nand U516 (N_516,N_441,N_379);
nor U517 (N_517,N_392,N_383);
nor U518 (N_518,N_415,N_391);
xor U519 (N_519,N_391,N_425);
xnor U520 (N_520,N_382,N_406);
nand U521 (N_521,N_404,N_446);
and U522 (N_522,N_422,N_430);
nor U523 (N_523,N_423,N_376);
and U524 (N_524,N_436,N_413);
or U525 (N_525,N_465,N_503);
nor U526 (N_526,N_521,N_509);
and U527 (N_527,N_462,N_460);
or U528 (N_528,N_496,N_517);
xnor U529 (N_529,N_461,N_502);
or U530 (N_530,N_522,N_501);
nand U531 (N_531,N_471,N_512);
and U532 (N_532,N_472,N_475);
xnor U533 (N_533,N_494,N_464);
nand U534 (N_534,N_516,N_515);
or U535 (N_535,N_476,N_491);
and U536 (N_536,N_489,N_490);
nor U537 (N_537,N_524,N_520);
nand U538 (N_538,N_470,N_485);
and U539 (N_539,N_452,N_519);
or U540 (N_540,N_523,N_518);
xor U541 (N_541,N_459,N_480);
nand U542 (N_542,N_506,N_469);
nor U543 (N_543,N_510,N_453);
nand U544 (N_544,N_505,N_511);
nor U545 (N_545,N_495,N_498);
nor U546 (N_546,N_451,N_497);
and U547 (N_547,N_477,N_456);
xnor U548 (N_548,N_499,N_487);
nor U549 (N_549,N_468,N_514);
xor U550 (N_550,N_500,N_450);
xor U551 (N_551,N_458,N_488);
or U552 (N_552,N_504,N_513);
or U553 (N_553,N_467,N_479);
xor U554 (N_554,N_483,N_457);
nor U555 (N_555,N_508,N_492);
and U556 (N_556,N_507,N_486);
nand U557 (N_557,N_481,N_463);
xor U558 (N_558,N_455,N_466);
or U559 (N_559,N_454,N_473);
xnor U560 (N_560,N_482,N_474);
nand U561 (N_561,N_484,N_478);
nand U562 (N_562,N_493,N_520);
nor U563 (N_563,N_502,N_501);
nor U564 (N_564,N_473,N_485);
xnor U565 (N_565,N_486,N_495);
or U566 (N_566,N_512,N_503);
and U567 (N_567,N_450,N_463);
xnor U568 (N_568,N_492,N_459);
and U569 (N_569,N_475,N_506);
xor U570 (N_570,N_476,N_480);
nand U571 (N_571,N_477,N_523);
or U572 (N_572,N_503,N_452);
nor U573 (N_573,N_490,N_498);
nand U574 (N_574,N_473,N_523);
nand U575 (N_575,N_488,N_487);
nand U576 (N_576,N_523,N_495);
and U577 (N_577,N_462,N_486);
and U578 (N_578,N_509,N_478);
nand U579 (N_579,N_457,N_511);
nor U580 (N_580,N_474,N_487);
nor U581 (N_581,N_482,N_459);
and U582 (N_582,N_513,N_507);
nand U583 (N_583,N_470,N_468);
or U584 (N_584,N_450,N_464);
nor U585 (N_585,N_523,N_498);
xnor U586 (N_586,N_456,N_470);
nor U587 (N_587,N_515,N_484);
nor U588 (N_588,N_497,N_514);
nand U589 (N_589,N_461,N_456);
xor U590 (N_590,N_484,N_511);
xnor U591 (N_591,N_523,N_488);
or U592 (N_592,N_506,N_466);
and U593 (N_593,N_469,N_502);
nor U594 (N_594,N_524,N_465);
xor U595 (N_595,N_508,N_460);
or U596 (N_596,N_466,N_491);
nand U597 (N_597,N_460,N_484);
or U598 (N_598,N_510,N_454);
and U599 (N_599,N_473,N_513);
xor U600 (N_600,N_566,N_599);
nor U601 (N_601,N_588,N_563);
and U602 (N_602,N_589,N_597);
nor U603 (N_603,N_546,N_577);
or U604 (N_604,N_525,N_531);
xor U605 (N_605,N_526,N_534);
nor U606 (N_606,N_532,N_539);
nand U607 (N_607,N_568,N_576);
xor U608 (N_608,N_595,N_573);
or U609 (N_609,N_536,N_586);
xor U610 (N_610,N_564,N_541);
or U611 (N_611,N_584,N_572);
xor U612 (N_612,N_587,N_569);
nor U613 (N_613,N_561,N_593);
and U614 (N_614,N_560,N_571);
nand U615 (N_615,N_548,N_596);
or U616 (N_616,N_538,N_562);
nand U617 (N_617,N_552,N_580);
and U618 (N_618,N_542,N_598);
and U619 (N_619,N_529,N_579);
and U620 (N_620,N_575,N_545);
xnor U621 (N_621,N_582,N_549);
nand U622 (N_622,N_527,N_547);
nand U623 (N_623,N_581,N_550);
xor U624 (N_624,N_594,N_583);
and U625 (N_625,N_530,N_551);
nor U626 (N_626,N_565,N_553);
or U627 (N_627,N_555,N_590);
or U628 (N_628,N_544,N_528);
and U629 (N_629,N_574,N_558);
or U630 (N_630,N_554,N_570);
xor U631 (N_631,N_559,N_543);
xnor U632 (N_632,N_537,N_540);
and U633 (N_633,N_533,N_585);
and U634 (N_634,N_557,N_591);
xnor U635 (N_635,N_578,N_535);
or U636 (N_636,N_567,N_592);
xnor U637 (N_637,N_556,N_557);
xnor U638 (N_638,N_535,N_587);
or U639 (N_639,N_593,N_570);
and U640 (N_640,N_566,N_541);
nor U641 (N_641,N_555,N_584);
nor U642 (N_642,N_596,N_535);
xnor U643 (N_643,N_593,N_588);
and U644 (N_644,N_542,N_534);
nand U645 (N_645,N_549,N_585);
and U646 (N_646,N_557,N_535);
and U647 (N_647,N_549,N_572);
nor U648 (N_648,N_594,N_543);
nor U649 (N_649,N_587,N_529);
nand U650 (N_650,N_554,N_541);
nor U651 (N_651,N_550,N_554);
nor U652 (N_652,N_585,N_542);
nand U653 (N_653,N_564,N_596);
nand U654 (N_654,N_593,N_545);
xnor U655 (N_655,N_587,N_574);
nand U656 (N_656,N_545,N_594);
xnor U657 (N_657,N_598,N_551);
xor U658 (N_658,N_580,N_541);
nand U659 (N_659,N_529,N_527);
or U660 (N_660,N_565,N_589);
nand U661 (N_661,N_574,N_591);
nor U662 (N_662,N_598,N_569);
and U663 (N_663,N_576,N_529);
nand U664 (N_664,N_575,N_544);
nor U665 (N_665,N_546,N_529);
nor U666 (N_666,N_578,N_527);
nor U667 (N_667,N_537,N_562);
or U668 (N_668,N_584,N_545);
or U669 (N_669,N_577,N_527);
nor U670 (N_670,N_597,N_554);
nor U671 (N_671,N_534,N_590);
nor U672 (N_672,N_572,N_556);
nand U673 (N_673,N_541,N_593);
nor U674 (N_674,N_563,N_570);
xnor U675 (N_675,N_670,N_605);
xnor U676 (N_676,N_657,N_674);
nand U677 (N_677,N_604,N_628);
nand U678 (N_678,N_627,N_671);
and U679 (N_679,N_669,N_606);
or U680 (N_680,N_664,N_634);
nand U681 (N_681,N_631,N_646);
or U682 (N_682,N_614,N_641);
nor U683 (N_683,N_621,N_635);
and U684 (N_684,N_600,N_619);
nor U685 (N_685,N_611,N_650);
or U686 (N_686,N_618,N_644);
nand U687 (N_687,N_659,N_672);
nand U688 (N_688,N_653,N_610);
and U689 (N_689,N_602,N_633);
xnor U690 (N_690,N_662,N_630);
or U691 (N_691,N_638,N_656);
xnor U692 (N_692,N_617,N_660);
nor U693 (N_693,N_608,N_648);
or U694 (N_694,N_607,N_667);
or U695 (N_695,N_651,N_654);
nand U696 (N_696,N_626,N_640);
and U697 (N_697,N_645,N_622);
nand U698 (N_698,N_609,N_649);
xor U699 (N_699,N_668,N_652);
xnor U700 (N_700,N_665,N_663);
or U701 (N_701,N_658,N_673);
nor U702 (N_702,N_643,N_603);
nor U703 (N_703,N_615,N_639);
xor U704 (N_704,N_616,N_624);
xnor U705 (N_705,N_625,N_642);
nor U706 (N_706,N_636,N_637);
and U707 (N_707,N_612,N_661);
xor U708 (N_708,N_613,N_601);
xor U709 (N_709,N_666,N_647);
nand U710 (N_710,N_623,N_620);
and U711 (N_711,N_655,N_629);
nand U712 (N_712,N_632,N_634);
xnor U713 (N_713,N_659,N_607);
nand U714 (N_714,N_673,N_644);
or U715 (N_715,N_666,N_623);
nor U716 (N_716,N_603,N_607);
nand U717 (N_717,N_670,N_654);
xor U718 (N_718,N_657,N_670);
nor U719 (N_719,N_602,N_630);
or U720 (N_720,N_638,N_662);
nand U721 (N_721,N_617,N_673);
and U722 (N_722,N_618,N_610);
and U723 (N_723,N_607,N_621);
or U724 (N_724,N_612,N_629);
xnor U725 (N_725,N_625,N_665);
nand U726 (N_726,N_647,N_621);
or U727 (N_727,N_638,N_664);
and U728 (N_728,N_653,N_616);
nand U729 (N_729,N_637,N_625);
or U730 (N_730,N_613,N_671);
and U731 (N_731,N_625,N_628);
nand U732 (N_732,N_635,N_634);
or U733 (N_733,N_615,N_607);
nand U734 (N_734,N_620,N_669);
and U735 (N_735,N_648,N_620);
and U736 (N_736,N_665,N_611);
xnor U737 (N_737,N_639,N_650);
or U738 (N_738,N_653,N_646);
and U739 (N_739,N_673,N_668);
or U740 (N_740,N_645,N_601);
nor U741 (N_741,N_665,N_671);
and U742 (N_742,N_654,N_665);
and U743 (N_743,N_661,N_638);
or U744 (N_744,N_666,N_649);
xor U745 (N_745,N_621,N_672);
or U746 (N_746,N_646,N_602);
nand U747 (N_747,N_641,N_640);
or U748 (N_748,N_643,N_604);
nand U749 (N_749,N_642,N_648);
or U750 (N_750,N_684,N_707);
xor U751 (N_751,N_727,N_720);
xnor U752 (N_752,N_733,N_701);
or U753 (N_753,N_677,N_712);
nor U754 (N_754,N_688,N_722);
xnor U755 (N_755,N_681,N_747);
or U756 (N_756,N_695,N_725);
and U757 (N_757,N_749,N_743);
nor U758 (N_758,N_711,N_742);
or U759 (N_759,N_737,N_675);
xor U760 (N_760,N_696,N_689);
or U761 (N_761,N_724,N_736);
nand U762 (N_762,N_682,N_691);
xor U763 (N_763,N_683,N_690);
nand U764 (N_764,N_716,N_694);
nor U765 (N_765,N_686,N_700);
or U766 (N_766,N_735,N_745);
nand U767 (N_767,N_715,N_740);
or U768 (N_768,N_706,N_697);
and U769 (N_769,N_744,N_714);
xor U770 (N_770,N_704,N_676);
nor U771 (N_771,N_746,N_731);
and U772 (N_772,N_708,N_734);
or U773 (N_773,N_723,N_693);
nor U774 (N_774,N_728,N_719);
nor U775 (N_775,N_698,N_730);
and U776 (N_776,N_717,N_721);
xnor U777 (N_777,N_748,N_710);
nor U778 (N_778,N_726,N_718);
and U779 (N_779,N_687,N_680);
and U780 (N_780,N_685,N_738);
and U781 (N_781,N_692,N_699);
nor U782 (N_782,N_709,N_705);
nor U783 (N_783,N_732,N_713);
xnor U784 (N_784,N_703,N_741);
nor U785 (N_785,N_702,N_679);
nand U786 (N_786,N_678,N_739);
xor U787 (N_787,N_729,N_726);
and U788 (N_788,N_705,N_736);
or U789 (N_789,N_739,N_725);
xor U790 (N_790,N_706,N_731);
nand U791 (N_791,N_704,N_689);
nand U792 (N_792,N_746,N_702);
and U793 (N_793,N_706,N_736);
or U794 (N_794,N_690,N_700);
xor U795 (N_795,N_740,N_733);
nor U796 (N_796,N_731,N_728);
nand U797 (N_797,N_749,N_732);
nor U798 (N_798,N_734,N_677);
nor U799 (N_799,N_710,N_742);
nand U800 (N_800,N_746,N_690);
or U801 (N_801,N_688,N_712);
or U802 (N_802,N_728,N_696);
nor U803 (N_803,N_718,N_709);
nor U804 (N_804,N_705,N_679);
nand U805 (N_805,N_683,N_678);
xnor U806 (N_806,N_680,N_741);
xor U807 (N_807,N_694,N_711);
nand U808 (N_808,N_689,N_712);
nor U809 (N_809,N_711,N_734);
nand U810 (N_810,N_700,N_689);
or U811 (N_811,N_693,N_675);
and U812 (N_812,N_747,N_732);
xnor U813 (N_813,N_717,N_698);
nand U814 (N_814,N_723,N_683);
nand U815 (N_815,N_723,N_712);
nor U816 (N_816,N_749,N_697);
nand U817 (N_817,N_693,N_707);
nand U818 (N_818,N_723,N_717);
nand U819 (N_819,N_681,N_711);
nand U820 (N_820,N_677,N_686);
and U821 (N_821,N_676,N_723);
nor U822 (N_822,N_690,N_677);
and U823 (N_823,N_735,N_748);
and U824 (N_824,N_677,N_698);
nor U825 (N_825,N_758,N_819);
nor U826 (N_826,N_756,N_820);
and U827 (N_827,N_787,N_776);
xor U828 (N_828,N_777,N_818);
and U829 (N_829,N_788,N_750);
and U830 (N_830,N_773,N_764);
or U831 (N_831,N_803,N_769);
or U832 (N_832,N_763,N_784);
or U833 (N_833,N_779,N_772);
xnor U834 (N_834,N_800,N_766);
nand U835 (N_835,N_770,N_780);
xnor U836 (N_836,N_786,N_761);
nand U837 (N_837,N_822,N_809);
nor U838 (N_838,N_753,N_790);
or U839 (N_839,N_806,N_782);
and U840 (N_840,N_801,N_798);
or U841 (N_841,N_795,N_767);
xor U842 (N_842,N_816,N_775);
xnor U843 (N_843,N_759,N_783);
and U844 (N_844,N_796,N_824);
and U845 (N_845,N_794,N_814);
nand U846 (N_846,N_754,N_765);
and U847 (N_847,N_813,N_771);
or U848 (N_848,N_817,N_823);
nor U849 (N_849,N_810,N_811);
nand U850 (N_850,N_815,N_797);
and U851 (N_851,N_791,N_799);
nor U852 (N_852,N_778,N_762);
xnor U853 (N_853,N_760,N_812);
nand U854 (N_854,N_752,N_808);
nand U855 (N_855,N_807,N_751);
xnor U856 (N_856,N_802,N_757);
nor U857 (N_857,N_792,N_789);
nand U858 (N_858,N_821,N_755);
and U859 (N_859,N_768,N_804);
xor U860 (N_860,N_774,N_805);
or U861 (N_861,N_785,N_793);
nand U862 (N_862,N_781,N_815);
or U863 (N_863,N_765,N_801);
nor U864 (N_864,N_752,N_758);
xor U865 (N_865,N_761,N_800);
and U866 (N_866,N_817,N_752);
nor U867 (N_867,N_813,N_798);
and U868 (N_868,N_750,N_821);
and U869 (N_869,N_765,N_796);
nand U870 (N_870,N_815,N_808);
nand U871 (N_871,N_779,N_754);
nand U872 (N_872,N_760,N_754);
xnor U873 (N_873,N_785,N_757);
xnor U874 (N_874,N_795,N_760);
nand U875 (N_875,N_815,N_809);
and U876 (N_876,N_790,N_798);
and U877 (N_877,N_800,N_758);
nor U878 (N_878,N_765,N_752);
nor U879 (N_879,N_766,N_797);
xor U880 (N_880,N_764,N_770);
nand U881 (N_881,N_817,N_801);
nand U882 (N_882,N_780,N_814);
nor U883 (N_883,N_764,N_824);
xnor U884 (N_884,N_758,N_812);
nand U885 (N_885,N_787,N_810);
and U886 (N_886,N_819,N_755);
or U887 (N_887,N_789,N_754);
xor U888 (N_888,N_802,N_800);
nor U889 (N_889,N_756,N_750);
or U890 (N_890,N_812,N_774);
and U891 (N_891,N_768,N_772);
nand U892 (N_892,N_803,N_810);
xor U893 (N_893,N_790,N_810);
and U894 (N_894,N_810,N_821);
or U895 (N_895,N_763,N_801);
nand U896 (N_896,N_775,N_788);
or U897 (N_897,N_754,N_806);
and U898 (N_898,N_787,N_798);
or U899 (N_899,N_758,N_753);
nor U900 (N_900,N_892,N_868);
and U901 (N_901,N_840,N_854);
or U902 (N_902,N_860,N_852);
nand U903 (N_903,N_838,N_850);
or U904 (N_904,N_862,N_885);
nand U905 (N_905,N_878,N_863);
and U906 (N_906,N_886,N_865);
or U907 (N_907,N_893,N_842);
or U908 (N_908,N_889,N_887);
nand U909 (N_909,N_855,N_837);
and U910 (N_910,N_830,N_825);
or U911 (N_911,N_828,N_880);
or U912 (N_912,N_826,N_829);
nor U913 (N_913,N_890,N_899);
xor U914 (N_914,N_839,N_876);
xnor U915 (N_915,N_881,N_869);
and U916 (N_916,N_894,N_846);
or U917 (N_917,N_895,N_882);
xor U918 (N_918,N_832,N_861);
and U919 (N_919,N_836,N_867);
or U920 (N_920,N_898,N_859);
and U921 (N_921,N_874,N_831);
xnor U922 (N_922,N_872,N_848);
xor U923 (N_923,N_873,N_897);
xor U924 (N_924,N_845,N_843);
or U925 (N_925,N_877,N_834);
nor U926 (N_926,N_864,N_875);
or U927 (N_927,N_866,N_833);
nand U928 (N_928,N_883,N_891);
nand U929 (N_929,N_856,N_844);
nand U930 (N_930,N_888,N_857);
xor U931 (N_931,N_870,N_871);
xnor U932 (N_932,N_827,N_879);
and U933 (N_933,N_847,N_896);
xor U934 (N_934,N_851,N_858);
nor U935 (N_935,N_849,N_835);
or U936 (N_936,N_853,N_841);
and U937 (N_937,N_884,N_838);
nor U938 (N_938,N_888,N_881);
and U939 (N_939,N_870,N_841);
nand U940 (N_940,N_885,N_872);
xor U941 (N_941,N_891,N_898);
nand U942 (N_942,N_876,N_880);
xnor U943 (N_943,N_890,N_833);
and U944 (N_944,N_883,N_863);
and U945 (N_945,N_877,N_885);
or U946 (N_946,N_841,N_871);
nand U947 (N_947,N_869,N_888);
or U948 (N_948,N_893,N_848);
and U949 (N_949,N_835,N_880);
or U950 (N_950,N_864,N_857);
xnor U951 (N_951,N_899,N_861);
and U952 (N_952,N_892,N_872);
xor U953 (N_953,N_831,N_864);
or U954 (N_954,N_854,N_865);
or U955 (N_955,N_896,N_871);
and U956 (N_956,N_864,N_836);
and U957 (N_957,N_856,N_828);
or U958 (N_958,N_853,N_840);
nor U959 (N_959,N_859,N_886);
nand U960 (N_960,N_894,N_825);
nor U961 (N_961,N_840,N_845);
xor U962 (N_962,N_834,N_867);
and U963 (N_963,N_878,N_852);
nand U964 (N_964,N_892,N_827);
nor U965 (N_965,N_856,N_865);
nand U966 (N_966,N_889,N_879);
xor U967 (N_967,N_835,N_836);
or U968 (N_968,N_875,N_869);
or U969 (N_969,N_889,N_883);
or U970 (N_970,N_877,N_852);
or U971 (N_971,N_856,N_853);
nor U972 (N_972,N_827,N_847);
nand U973 (N_973,N_850,N_883);
nand U974 (N_974,N_895,N_849);
nand U975 (N_975,N_914,N_912);
and U976 (N_976,N_913,N_949);
and U977 (N_977,N_941,N_904);
or U978 (N_978,N_907,N_969);
and U979 (N_979,N_973,N_908);
xor U980 (N_980,N_910,N_944);
or U981 (N_981,N_936,N_964);
or U982 (N_982,N_924,N_929);
xnor U983 (N_983,N_923,N_947);
nor U984 (N_984,N_943,N_921);
or U985 (N_985,N_946,N_906);
xor U986 (N_986,N_959,N_958);
nor U987 (N_987,N_902,N_970);
and U988 (N_988,N_917,N_963);
nor U989 (N_989,N_920,N_905);
or U990 (N_990,N_931,N_953);
or U991 (N_991,N_915,N_942);
nor U992 (N_992,N_940,N_956);
or U993 (N_993,N_925,N_909);
xnor U994 (N_994,N_932,N_957);
and U995 (N_995,N_922,N_901);
xor U996 (N_996,N_954,N_927);
or U997 (N_997,N_974,N_926);
and U998 (N_998,N_948,N_919);
or U999 (N_999,N_968,N_952);
and U1000 (N_1000,N_967,N_955);
xor U1001 (N_1001,N_928,N_900);
nor U1002 (N_1002,N_935,N_962);
xor U1003 (N_1003,N_972,N_934);
or U1004 (N_1004,N_950,N_961);
nand U1005 (N_1005,N_960,N_933);
nand U1006 (N_1006,N_966,N_916);
xor U1007 (N_1007,N_939,N_911);
nor U1008 (N_1008,N_937,N_945);
xnor U1009 (N_1009,N_903,N_930);
nand U1010 (N_1010,N_938,N_918);
and U1011 (N_1011,N_951,N_965);
xor U1012 (N_1012,N_971,N_962);
and U1013 (N_1013,N_970,N_968);
nand U1014 (N_1014,N_901,N_914);
and U1015 (N_1015,N_900,N_957);
or U1016 (N_1016,N_905,N_950);
and U1017 (N_1017,N_916,N_973);
and U1018 (N_1018,N_903,N_952);
and U1019 (N_1019,N_905,N_957);
nor U1020 (N_1020,N_933,N_922);
or U1021 (N_1021,N_924,N_950);
xnor U1022 (N_1022,N_900,N_941);
nand U1023 (N_1023,N_924,N_914);
or U1024 (N_1024,N_960,N_925);
and U1025 (N_1025,N_914,N_932);
nor U1026 (N_1026,N_916,N_964);
xor U1027 (N_1027,N_903,N_973);
and U1028 (N_1028,N_931,N_961);
nand U1029 (N_1029,N_952,N_907);
xor U1030 (N_1030,N_906,N_912);
xnor U1031 (N_1031,N_903,N_901);
xnor U1032 (N_1032,N_951,N_946);
xnor U1033 (N_1033,N_966,N_908);
and U1034 (N_1034,N_970,N_955);
or U1035 (N_1035,N_952,N_925);
nor U1036 (N_1036,N_945,N_943);
xor U1037 (N_1037,N_947,N_922);
or U1038 (N_1038,N_904,N_928);
or U1039 (N_1039,N_927,N_909);
or U1040 (N_1040,N_932,N_904);
or U1041 (N_1041,N_904,N_954);
nand U1042 (N_1042,N_903,N_908);
xor U1043 (N_1043,N_909,N_951);
xor U1044 (N_1044,N_905,N_946);
nor U1045 (N_1045,N_949,N_943);
and U1046 (N_1046,N_955,N_912);
nor U1047 (N_1047,N_919,N_968);
nand U1048 (N_1048,N_957,N_961);
or U1049 (N_1049,N_972,N_909);
xnor U1050 (N_1050,N_1014,N_1040);
nor U1051 (N_1051,N_986,N_1018);
xnor U1052 (N_1052,N_1001,N_1041);
or U1053 (N_1053,N_1035,N_1002);
or U1054 (N_1054,N_1027,N_984);
xor U1055 (N_1055,N_1032,N_992);
nor U1056 (N_1056,N_977,N_988);
xnor U1057 (N_1057,N_1009,N_997);
or U1058 (N_1058,N_993,N_978);
nor U1059 (N_1059,N_1036,N_1024);
or U1060 (N_1060,N_1016,N_1042);
xnor U1061 (N_1061,N_1011,N_976);
nand U1062 (N_1062,N_975,N_1007);
and U1063 (N_1063,N_1022,N_985);
xnor U1064 (N_1064,N_1047,N_983);
xor U1065 (N_1065,N_1012,N_1017);
nand U1066 (N_1066,N_1030,N_1004);
nor U1067 (N_1067,N_1025,N_980);
xor U1068 (N_1068,N_1029,N_1023);
or U1069 (N_1069,N_1046,N_1021);
nand U1070 (N_1070,N_1026,N_987);
nor U1071 (N_1071,N_999,N_1033);
and U1072 (N_1072,N_1013,N_1031);
nor U1073 (N_1073,N_1039,N_1028);
or U1074 (N_1074,N_996,N_1020);
or U1075 (N_1075,N_1005,N_1019);
nor U1076 (N_1076,N_1015,N_991);
xnor U1077 (N_1077,N_990,N_1000);
nor U1078 (N_1078,N_1049,N_994);
and U1079 (N_1079,N_1008,N_1010);
xor U1080 (N_1080,N_982,N_1037);
xor U1081 (N_1081,N_1044,N_1003);
nand U1082 (N_1082,N_1034,N_1045);
or U1083 (N_1083,N_1006,N_1048);
nand U1084 (N_1084,N_1038,N_998);
or U1085 (N_1085,N_995,N_1043);
nor U1086 (N_1086,N_989,N_979);
nand U1087 (N_1087,N_981,N_1007);
or U1088 (N_1088,N_1012,N_990);
nor U1089 (N_1089,N_1002,N_1011);
xnor U1090 (N_1090,N_991,N_1027);
nand U1091 (N_1091,N_1011,N_1046);
xor U1092 (N_1092,N_995,N_996);
and U1093 (N_1093,N_1031,N_1009);
or U1094 (N_1094,N_1035,N_997);
nand U1095 (N_1095,N_1037,N_1049);
xor U1096 (N_1096,N_1044,N_1004);
or U1097 (N_1097,N_1026,N_984);
xnor U1098 (N_1098,N_1007,N_1034);
and U1099 (N_1099,N_990,N_978);
xnor U1100 (N_1100,N_1034,N_997);
and U1101 (N_1101,N_987,N_984);
or U1102 (N_1102,N_1028,N_1013);
nor U1103 (N_1103,N_1038,N_1037);
xor U1104 (N_1104,N_1034,N_1032);
nand U1105 (N_1105,N_990,N_1044);
nor U1106 (N_1106,N_1029,N_1015);
nor U1107 (N_1107,N_983,N_989);
and U1108 (N_1108,N_981,N_977);
and U1109 (N_1109,N_1023,N_1038);
nor U1110 (N_1110,N_977,N_1042);
or U1111 (N_1111,N_981,N_1004);
xnor U1112 (N_1112,N_1025,N_1023);
and U1113 (N_1113,N_996,N_1003);
nor U1114 (N_1114,N_1019,N_1046);
and U1115 (N_1115,N_986,N_1026);
and U1116 (N_1116,N_1026,N_1020);
nand U1117 (N_1117,N_1041,N_993);
nor U1118 (N_1118,N_976,N_1029);
xor U1119 (N_1119,N_1019,N_1018);
nor U1120 (N_1120,N_992,N_1005);
nor U1121 (N_1121,N_1023,N_984);
xor U1122 (N_1122,N_993,N_1048);
and U1123 (N_1123,N_1041,N_1030);
or U1124 (N_1124,N_1008,N_1020);
nand U1125 (N_1125,N_1061,N_1112);
nand U1126 (N_1126,N_1109,N_1121);
or U1127 (N_1127,N_1067,N_1094);
nand U1128 (N_1128,N_1091,N_1097);
nor U1129 (N_1129,N_1092,N_1056);
xor U1130 (N_1130,N_1096,N_1055);
and U1131 (N_1131,N_1059,N_1072);
xor U1132 (N_1132,N_1071,N_1050);
xor U1133 (N_1133,N_1074,N_1058);
or U1134 (N_1134,N_1060,N_1081);
and U1135 (N_1135,N_1117,N_1122);
nor U1136 (N_1136,N_1062,N_1107);
xnor U1137 (N_1137,N_1082,N_1080);
nand U1138 (N_1138,N_1084,N_1115);
nor U1139 (N_1139,N_1098,N_1053);
or U1140 (N_1140,N_1076,N_1085);
xor U1141 (N_1141,N_1095,N_1101);
nand U1142 (N_1142,N_1124,N_1075);
nand U1143 (N_1143,N_1100,N_1119);
or U1144 (N_1144,N_1078,N_1114);
or U1145 (N_1145,N_1123,N_1087);
or U1146 (N_1146,N_1073,N_1057);
nor U1147 (N_1147,N_1118,N_1054);
or U1148 (N_1148,N_1069,N_1063);
nand U1149 (N_1149,N_1093,N_1110);
or U1150 (N_1150,N_1083,N_1090);
nand U1151 (N_1151,N_1089,N_1104);
nand U1152 (N_1152,N_1065,N_1108);
nor U1153 (N_1153,N_1077,N_1111);
xnor U1154 (N_1154,N_1105,N_1052);
xnor U1155 (N_1155,N_1070,N_1099);
nor U1156 (N_1156,N_1079,N_1102);
or U1157 (N_1157,N_1086,N_1116);
xor U1158 (N_1158,N_1064,N_1088);
xnor U1159 (N_1159,N_1103,N_1051);
nor U1160 (N_1160,N_1106,N_1113);
nand U1161 (N_1161,N_1068,N_1066);
nor U1162 (N_1162,N_1120,N_1110);
and U1163 (N_1163,N_1094,N_1113);
or U1164 (N_1164,N_1094,N_1061);
and U1165 (N_1165,N_1106,N_1097);
nand U1166 (N_1166,N_1057,N_1112);
xor U1167 (N_1167,N_1080,N_1123);
and U1168 (N_1168,N_1072,N_1062);
xnor U1169 (N_1169,N_1114,N_1083);
xnor U1170 (N_1170,N_1052,N_1092);
and U1171 (N_1171,N_1109,N_1107);
xnor U1172 (N_1172,N_1102,N_1077);
and U1173 (N_1173,N_1061,N_1079);
and U1174 (N_1174,N_1102,N_1084);
nand U1175 (N_1175,N_1083,N_1112);
and U1176 (N_1176,N_1064,N_1107);
xnor U1177 (N_1177,N_1067,N_1050);
and U1178 (N_1178,N_1075,N_1076);
and U1179 (N_1179,N_1124,N_1106);
or U1180 (N_1180,N_1108,N_1097);
nand U1181 (N_1181,N_1082,N_1055);
xnor U1182 (N_1182,N_1082,N_1103);
and U1183 (N_1183,N_1110,N_1094);
or U1184 (N_1184,N_1117,N_1112);
or U1185 (N_1185,N_1050,N_1122);
or U1186 (N_1186,N_1092,N_1084);
nor U1187 (N_1187,N_1092,N_1074);
xor U1188 (N_1188,N_1117,N_1101);
or U1189 (N_1189,N_1057,N_1102);
nor U1190 (N_1190,N_1083,N_1086);
nand U1191 (N_1191,N_1098,N_1114);
and U1192 (N_1192,N_1100,N_1054);
or U1193 (N_1193,N_1050,N_1054);
nand U1194 (N_1194,N_1115,N_1089);
and U1195 (N_1195,N_1065,N_1116);
xor U1196 (N_1196,N_1078,N_1060);
or U1197 (N_1197,N_1121,N_1105);
nor U1198 (N_1198,N_1065,N_1099);
xnor U1199 (N_1199,N_1120,N_1088);
nor U1200 (N_1200,N_1180,N_1164);
and U1201 (N_1201,N_1140,N_1175);
or U1202 (N_1202,N_1126,N_1172);
and U1203 (N_1203,N_1149,N_1162);
nand U1204 (N_1204,N_1195,N_1135);
xnor U1205 (N_1205,N_1129,N_1196);
xnor U1206 (N_1206,N_1144,N_1194);
and U1207 (N_1207,N_1141,N_1167);
xor U1208 (N_1208,N_1134,N_1138);
nor U1209 (N_1209,N_1130,N_1145);
nor U1210 (N_1210,N_1127,N_1179);
and U1211 (N_1211,N_1166,N_1197);
xnor U1212 (N_1212,N_1173,N_1128);
nor U1213 (N_1213,N_1158,N_1131);
or U1214 (N_1214,N_1189,N_1160);
and U1215 (N_1215,N_1181,N_1155);
xnor U1216 (N_1216,N_1177,N_1168);
and U1217 (N_1217,N_1132,N_1146);
xor U1218 (N_1218,N_1186,N_1142);
nand U1219 (N_1219,N_1137,N_1191);
nor U1220 (N_1220,N_1185,N_1187);
nand U1221 (N_1221,N_1136,N_1154);
and U1222 (N_1222,N_1163,N_1171);
xnor U1223 (N_1223,N_1161,N_1139);
nor U1224 (N_1224,N_1157,N_1176);
nand U1225 (N_1225,N_1170,N_1184);
and U1226 (N_1226,N_1152,N_1159);
nor U1227 (N_1227,N_1143,N_1150);
nand U1228 (N_1228,N_1193,N_1183);
or U1229 (N_1229,N_1151,N_1125);
or U1230 (N_1230,N_1148,N_1188);
or U1231 (N_1231,N_1169,N_1153);
nand U1232 (N_1232,N_1133,N_1147);
nand U1233 (N_1233,N_1190,N_1182);
and U1234 (N_1234,N_1198,N_1156);
nand U1235 (N_1235,N_1174,N_1165);
or U1236 (N_1236,N_1199,N_1192);
xnor U1237 (N_1237,N_1178,N_1144);
xnor U1238 (N_1238,N_1198,N_1132);
xor U1239 (N_1239,N_1145,N_1176);
nand U1240 (N_1240,N_1131,N_1145);
nor U1241 (N_1241,N_1140,N_1173);
or U1242 (N_1242,N_1186,N_1158);
xor U1243 (N_1243,N_1159,N_1135);
xnor U1244 (N_1244,N_1147,N_1183);
nand U1245 (N_1245,N_1132,N_1190);
nand U1246 (N_1246,N_1183,N_1197);
or U1247 (N_1247,N_1186,N_1179);
xnor U1248 (N_1248,N_1199,N_1141);
nor U1249 (N_1249,N_1185,N_1174);
nor U1250 (N_1250,N_1196,N_1194);
and U1251 (N_1251,N_1172,N_1166);
xnor U1252 (N_1252,N_1180,N_1186);
or U1253 (N_1253,N_1178,N_1182);
xor U1254 (N_1254,N_1128,N_1164);
or U1255 (N_1255,N_1167,N_1188);
or U1256 (N_1256,N_1181,N_1154);
nor U1257 (N_1257,N_1128,N_1138);
nor U1258 (N_1258,N_1146,N_1193);
nand U1259 (N_1259,N_1145,N_1186);
and U1260 (N_1260,N_1151,N_1154);
xor U1261 (N_1261,N_1146,N_1195);
xnor U1262 (N_1262,N_1188,N_1156);
or U1263 (N_1263,N_1190,N_1191);
xnor U1264 (N_1264,N_1183,N_1132);
nor U1265 (N_1265,N_1186,N_1169);
or U1266 (N_1266,N_1170,N_1127);
or U1267 (N_1267,N_1175,N_1168);
and U1268 (N_1268,N_1172,N_1147);
nor U1269 (N_1269,N_1137,N_1171);
or U1270 (N_1270,N_1127,N_1169);
and U1271 (N_1271,N_1199,N_1152);
xor U1272 (N_1272,N_1196,N_1173);
and U1273 (N_1273,N_1194,N_1191);
and U1274 (N_1274,N_1167,N_1194);
or U1275 (N_1275,N_1240,N_1227);
and U1276 (N_1276,N_1244,N_1225);
xor U1277 (N_1277,N_1226,N_1241);
nand U1278 (N_1278,N_1247,N_1246);
nor U1279 (N_1279,N_1222,N_1210);
nor U1280 (N_1280,N_1209,N_1268);
and U1281 (N_1281,N_1250,N_1205);
nor U1282 (N_1282,N_1208,N_1274);
nor U1283 (N_1283,N_1239,N_1218);
nand U1284 (N_1284,N_1242,N_1215);
xor U1285 (N_1285,N_1223,N_1270);
nor U1286 (N_1286,N_1235,N_1273);
and U1287 (N_1287,N_1204,N_1252);
or U1288 (N_1288,N_1266,N_1200);
and U1289 (N_1289,N_1214,N_1253);
or U1290 (N_1290,N_1262,N_1257);
nor U1291 (N_1291,N_1249,N_1269);
xnor U1292 (N_1292,N_1264,N_1217);
xor U1293 (N_1293,N_1263,N_1231);
or U1294 (N_1294,N_1228,N_1202);
nand U1295 (N_1295,N_1206,N_1220);
nand U1296 (N_1296,N_1213,N_1233);
or U1297 (N_1297,N_1259,N_1261);
and U1298 (N_1298,N_1238,N_1251);
nand U1299 (N_1299,N_1256,N_1255);
nor U1300 (N_1300,N_1224,N_1237);
nor U1301 (N_1301,N_1272,N_1260);
nand U1302 (N_1302,N_1258,N_1211);
nand U1303 (N_1303,N_1229,N_1203);
nand U1304 (N_1304,N_1230,N_1243);
and U1305 (N_1305,N_1245,N_1248);
xnor U1306 (N_1306,N_1207,N_1271);
nand U1307 (N_1307,N_1221,N_1254);
or U1308 (N_1308,N_1216,N_1265);
or U1309 (N_1309,N_1236,N_1234);
and U1310 (N_1310,N_1212,N_1219);
xor U1311 (N_1311,N_1232,N_1267);
nand U1312 (N_1312,N_1201,N_1243);
and U1313 (N_1313,N_1207,N_1258);
nor U1314 (N_1314,N_1233,N_1260);
xnor U1315 (N_1315,N_1231,N_1219);
xnor U1316 (N_1316,N_1240,N_1234);
xor U1317 (N_1317,N_1269,N_1218);
xor U1318 (N_1318,N_1223,N_1263);
and U1319 (N_1319,N_1209,N_1240);
nor U1320 (N_1320,N_1260,N_1216);
xor U1321 (N_1321,N_1214,N_1256);
or U1322 (N_1322,N_1246,N_1241);
nand U1323 (N_1323,N_1216,N_1217);
nand U1324 (N_1324,N_1205,N_1265);
nor U1325 (N_1325,N_1267,N_1201);
and U1326 (N_1326,N_1258,N_1247);
xnor U1327 (N_1327,N_1212,N_1236);
nand U1328 (N_1328,N_1260,N_1226);
or U1329 (N_1329,N_1202,N_1233);
nor U1330 (N_1330,N_1218,N_1207);
or U1331 (N_1331,N_1239,N_1260);
xnor U1332 (N_1332,N_1224,N_1241);
xor U1333 (N_1333,N_1265,N_1236);
and U1334 (N_1334,N_1255,N_1236);
and U1335 (N_1335,N_1231,N_1223);
nor U1336 (N_1336,N_1222,N_1240);
or U1337 (N_1337,N_1261,N_1250);
nor U1338 (N_1338,N_1201,N_1270);
nor U1339 (N_1339,N_1250,N_1204);
nand U1340 (N_1340,N_1213,N_1209);
nor U1341 (N_1341,N_1260,N_1254);
xnor U1342 (N_1342,N_1240,N_1238);
xor U1343 (N_1343,N_1249,N_1229);
or U1344 (N_1344,N_1264,N_1228);
or U1345 (N_1345,N_1247,N_1234);
or U1346 (N_1346,N_1237,N_1212);
nor U1347 (N_1347,N_1244,N_1216);
nand U1348 (N_1348,N_1225,N_1229);
or U1349 (N_1349,N_1231,N_1234);
or U1350 (N_1350,N_1330,N_1317);
nor U1351 (N_1351,N_1285,N_1298);
nand U1352 (N_1352,N_1314,N_1294);
and U1353 (N_1353,N_1291,N_1299);
and U1354 (N_1354,N_1324,N_1303);
nand U1355 (N_1355,N_1290,N_1309);
and U1356 (N_1356,N_1307,N_1341);
and U1357 (N_1357,N_1284,N_1310);
and U1358 (N_1358,N_1321,N_1293);
and U1359 (N_1359,N_1275,N_1339);
nand U1360 (N_1360,N_1322,N_1302);
nor U1361 (N_1361,N_1287,N_1342);
nor U1362 (N_1362,N_1277,N_1311);
xor U1363 (N_1363,N_1347,N_1343);
xnor U1364 (N_1364,N_1279,N_1283);
nand U1365 (N_1365,N_1337,N_1282);
nand U1366 (N_1366,N_1316,N_1278);
nor U1367 (N_1367,N_1296,N_1335);
and U1368 (N_1368,N_1327,N_1280);
and U1369 (N_1369,N_1313,N_1292);
nor U1370 (N_1370,N_1295,N_1331);
nand U1371 (N_1371,N_1306,N_1346);
or U1372 (N_1372,N_1276,N_1315);
nor U1373 (N_1373,N_1328,N_1326);
and U1374 (N_1374,N_1301,N_1340);
and U1375 (N_1375,N_1286,N_1312);
xnor U1376 (N_1376,N_1305,N_1334);
or U1377 (N_1377,N_1338,N_1319);
nor U1378 (N_1378,N_1300,N_1333);
or U1379 (N_1379,N_1329,N_1323);
xnor U1380 (N_1380,N_1345,N_1332);
xor U1381 (N_1381,N_1289,N_1288);
and U1382 (N_1382,N_1297,N_1281);
nor U1383 (N_1383,N_1304,N_1344);
nor U1384 (N_1384,N_1318,N_1320);
nand U1385 (N_1385,N_1325,N_1348);
or U1386 (N_1386,N_1308,N_1336);
or U1387 (N_1387,N_1349,N_1328);
xnor U1388 (N_1388,N_1279,N_1296);
xor U1389 (N_1389,N_1329,N_1304);
and U1390 (N_1390,N_1325,N_1283);
and U1391 (N_1391,N_1279,N_1310);
xor U1392 (N_1392,N_1317,N_1340);
nor U1393 (N_1393,N_1277,N_1298);
or U1394 (N_1394,N_1280,N_1346);
and U1395 (N_1395,N_1318,N_1334);
nor U1396 (N_1396,N_1326,N_1298);
xnor U1397 (N_1397,N_1287,N_1308);
and U1398 (N_1398,N_1316,N_1304);
and U1399 (N_1399,N_1343,N_1334);
xor U1400 (N_1400,N_1291,N_1285);
xnor U1401 (N_1401,N_1277,N_1342);
and U1402 (N_1402,N_1288,N_1316);
and U1403 (N_1403,N_1276,N_1347);
or U1404 (N_1404,N_1335,N_1280);
nand U1405 (N_1405,N_1330,N_1343);
xnor U1406 (N_1406,N_1280,N_1347);
xor U1407 (N_1407,N_1347,N_1338);
nor U1408 (N_1408,N_1347,N_1293);
xor U1409 (N_1409,N_1303,N_1297);
xor U1410 (N_1410,N_1305,N_1310);
nor U1411 (N_1411,N_1276,N_1314);
nor U1412 (N_1412,N_1319,N_1285);
nor U1413 (N_1413,N_1300,N_1290);
xor U1414 (N_1414,N_1347,N_1345);
nand U1415 (N_1415,N_1302,N_1308);
xnor U1416 (N_1416,N_1342,N_1278);
and U1417 (N_1417,N_1279,N_1319);
xnor U1418 (N_1418,N_1278,N_1291);
nor U1419 (N_1419,N_1300,N_1299);
nor U1420 (N_1420,N_1331,N_1316);
xor U1421 (N_1421,N_1278,N_1310);
xor U1422 (N_1422,N_1308,N_1344);
nor U1423 (N_1423,N_1331,N_1300);
or U1424 (N_1424,N_1346,N_1304);
nand U1425 (N_1425,N_1414,N_1389);
or U1426 (N_1426,N_1364,N_1413);
xor U1427 (N_1427,N_1387,N_1400);
and U1428 (N_1428,N_1373,N_1422);
nor U1429 (N_1429,N_1369,N_1412);
nand U1430 (N_1430,N_1352,N_1381);
and U1431 (N_1431,N_1351,N_1410);
or U1432 (N_1432,N_1367,N_1376);
or U1433 (N_1433,N_1372,N_1393);
or U1434 (N_1434,N_1355,N_1365);
nand U1435 (N_1435,N_1380,N_1417);
or U1436 (N_1436,N_1406,N_1419);
xnor U1437 (N_1437,N_1392,N_1424);
or U1438 (N_1438,N_1363,N_1421);
or U1439 (N_1439,N_1362,N_1359);
and U1440 (N_1440,N_1388,N_1382);
xnor U1441 (N_1441,N_1350,N_1370);
and U1442 (N_1442,N_1383,N_1357);
and U1443 (N_1443,N_1407,N_1423);
or U1444 (N_1444,N_1408,N_1356);
nor U1445 (N_1445,N_1366,N_1399);
xnor U1446 (N_1446,N_1371,N_1416);
and U1447 (N_1447,N_1402,N_1404);
nor U1448 (N_1448,N_1354,N_1384);
nor U1449 (N_1449,N_1377,N_1397);
and U1450 (N_1450,N_1358,N_1403);
nand U1451 (N_1451,N_1418,N_1398);
or U1452 (N_1452,N_1386,N_1395);
or U1453 (N_1453,N_1409,N_1415);
xor U1454 (N_1454,N_1360,N_1390);
and U1455 (N_1455,N_1385,N_1368);
nand U1456 (N_1456,N_1391,N_1405);
or U1457 (N_1457,N_1394,N_1378);
nand U1458 (N_1458,N_1353,N_1361);
nand U1459 (N_1459,N_1420,N_1375);
xor U1460 (N_1460,N_1374,N_1379);
nand U1461 (N_1461,N_1396,N_1411);
nand U1462 (N_1462,N_1401,N_1359);
nor U1463 (N_1463,N_1422,N_1402);
nor U1464 (N_1464,N_1413,N_1411);
xor U1465 (N_1465,N_1352,N_1420);
or U1466 (N_1466,N_1419,N_1386);
or U1467 (N_1467,N_1416,N_1387);
nand U1468 (N_1468,N_1366,N_1371);
nand U1469 (N_1469,N_1396,N_1385);
and U1470 (N_1470,N_1383,N_1419);
or U1471 (N_1471,N_1398,N_1408);
nor U1472 (N_1472,N_1361,N_1383);
or U1473 (N_1473,N_1402,N_1355);
xor U1474 (N_1474,N_1386,N_1421);
and U1475 (N_1475,N_1373,N_1385);
or U1476 (N_1476,N_1424,N_1410);
or U1477 (N_1477,N_1397,N_1363);
or U1478 (N_1478,N_1369,N_1410);
xnor U1479 (N_1479,N_1401,N_1357);
and U1480 (N_1480,N_1372,N_1420);
nand U1481 (N_1481,N_1375,N_1374);
or U1482 (N_1482,N_1385,N_1369);
or U1483 (N_1483,N_1397,N_1351);
xnor U1484 (N_1484,N_1371,N_1410);
nor U1485 (N_1485,N_1362,N_1358);
and U1486 (N_1486,N_1414,N_1374);
nor U1487 (N_1487,N_1396,N_1360);
nor U1488 (N_1488,N_1389,N_1371);
nand U1489 (N_1489,N_1378,N_1363);
nor U1490 (N_1490,N_1376,N_1374);
and U1491 (N_1491,N_1423,N_1383);
or U1492 (N_1492,N_1394,N_1402);
nor U1493 (N_1493,N_1395,N_1356);
nor U1494 (N_1494,N_1381,N_1403);
or U1495 (N_1495,N_1415,N_1407);
nand U1496 (N_1496,N_1384,N_1365);
nand U1497 (N_1497,N_1372,N_1365);
xor U1498 (N_1498,N_1356,N_1386);
and U1499 (N_1499,N_1359,N_1352);
or U1500 (N_1500,N_1432,N_1467);
xnor U1501 (N_1501,N_1459,N_1473);
or U1502 (N_1502,N_1443,N_1426);
or U1503 (N_1503,N_1493,N_1430);
nand U1504 (N_1504,N_1450,N_1462);
nor U1505 (N_1505,N_1442,N_1435);
and U1506 (N_1506,N_1455,N_1497);
nand U1507 (N_1507,N_1492,N_1481);
nor U1508 (N_1508,N_1491,N_1496);
nor U1509 (N_1509,N_1431,N_1485);
nor U1510 (N_1510,N_1474,N_1427);
and U1511 (N_1511,N_1464,N_1495);
and U1512 (N_1512,N_1449,N_1444);
or U1513 (N_1513,N_1440,N_1483);
xor U1514 (N_1514,N_1461,N_1452);
nand U1515 (N_1515,N_1438,N_1482);
nand U1516 (N_1516,N_1479,N_1490);
nand U1517 (N_1517,N_1470,N_1439);
and U1518 (N_1518,N_1477,N_1499);
and U1519 (N_1519,N_1437,N_1475);
nand U1520 (N_1520,N_1447,N_1460);
xnor U1521 (N_1521,N_1458,N_1457);
xor U1522 (N_1522,N_1434,N_1466);
nand U1523 (N_1523,N_1468,N_1463);
nand U1524 (N_1524,N_1471,N_1480);
xnor U1525 (N_1525,N_1451,N_1433);
xor U1526 (N_1526,N_1428,N_1478);
xor U1527 (N_1527,N_1446,N_1489);
xnor U1528 (N_1528,N_1454,N_1445);
and U1529 (N_1529,N_1472,N_1476);
or U1530 (N_1530,N_1456,N_1487);
xor U1531 (N_1531,N_1448,N_1453);
nor U1532 (N_1532,N_1488,N_1425);
nand U1533 (N_1533,N_1441,N_1484);
xnor U1534 (N_1534,N_1498,N_1436);
or U1535 (N_1535,N_1494,N_1429);
and U1536 (N_1536,N_1469,N_1486);
or U1537 (N_1537,N_1465,N_1491);
nand U1538 (N_1538,N_1468,N_1460);
nor U1539 (N_1539,N_1477,N_1485);
and U1540 (N_1540,N_1494,N_1444);
or U1541 (N_1541,N_1437,N_1443);
xor U1542 (N_1542,N_1489,N_1431);
nand U1543 (N_1543,N_1454,N_1472);
or U1544 (N_1544,N_1475,N_1485);
xnor U1545 (N_1545,N_1495,N_1459);
or U1546 (N_1546,N_1459,N_1463);
nand U1547 (N_1547,N_1442,N_1449);
nor U1548 (N_1548,N_1445,N_1456);
or U1549 (N_1549,N_1468,N_1498);
and U1550 (N_1550,N_1483,N_1429);
nor U1551 (N_1551,N_1483,N_1427);
or U1552 (N_1552,N_1447,N_1480);
or U1553 (N_1553,N_1427,N_1460);
or U1554 (N_1554,N_1431,N_1497);
and U1555 (N_1555,N_1462,N_1435);
xnor U1556 (N_1556,N_1495,N_1436);
nand U1557 (N_1557,N_1444,N_1466);
and U1558 (N_1558,N_1497,N_1490);
xnor U1559 (N_1559,N_1454,N_1444);
and U1560 (N_1560,N_1451,N_1482);
nor U1561 (N_1561,N_1480,N_1493);
nand U1562 (N_1562,N_1478,N_1458);
and U1563 (N_1563,N_1467,N_1436);
xor U1564 (N_1564,N_1476,N_1492);
and U1565 (N_1565,N_1490,N_1429);
nand U1566 (N_1566,N_1442,N_1489);
and U1567 (N_1567,N_1461,N_1492);
or U1568 (N_1568,N_1428,N_1470);
xnor U1569 (N_1569,N_1427,N_1466);
and U1570 (N_1570,N_1446,N_1476);
nand U1571 (N_1571,N_1468,N_1454);
or U1572 (N_1572,N_1426,N_1466);
nor U1573 (N_1573,N_1467,N_1445);
nand U1574 (N_1574,N_1485,N_1498);
xor U1575 (N_1575,N_1573,N_1550);
xor U1576 (N_1576,N_1511,N_1565);
and U1577 (N_1577,N_1520,N_1508);
nand U1578 (N_1578,N_1566,N_1562);
nand U1579 (N_1579,N_1540,N_1500);
xor U1580 (N_1580,N_1564,N_1507);
nand U1581 (N_1581,N_1571,N_1522);
nand U1582 (N_1582,N_1574,N_1559);
nand U1583 (N_1583,N_1518,N_1521);
and U1584 (N_1584,N_1536,N_1557);
or U1585 (N_1585,N_1505,N_1553);
and U1586 (N_1586,N_1560,N_1572);
nand U1587 (N_1587,N_1541,N_1510);
and U1588 (N_1588,N_1561,N_1529);
nor U1589 (N_1589,N_1516,N_1525);
or U1590 (N_1590,N_1567,N_1558);
nor U1591 (N_1591,N_1502,N_1534);
or U1592 (N_1592,N_1530,N_1531);
nor U1593 (N_1593,N_1570,N_1547);
nand U1594 (N_1594,N_1535,N_1546);
and U1595 (N_1595,N_1503,N_1515);
and U1596 (N_1596,N_1528,N_1537);
and U1597 (N_1597,N_1506,N_1527);
nand U1598 (N_1598,N_1538,N_1556);
or U1599 (N_1599,N_1501,N_1568);
and U1600 (N_1600,N_1548,N_1549);
nor U1601 (N_1601,N_1554,N_1551);
and U1602 (N_1602,N_1544,N_1555);
nor U1603 (N_1603,N_1513,N_1509);
xnor U1604 (N_1604,N_1514,N_1545);
xor U1605 (N_1605,N_1512,N_1523);
or U1606 (N_1606,N_1532,N_1563);
nor U1607 (N_1607,N_1533,N_1552);
and U1608 (N_1608,N_1569,N_1519);
nor U1609 (N_1609,N_1542,N_1526);
or U1610 (N_1610,N_1543,N_1524);
nor U1611 (N_1611,N_1517,N_1539);
and U1612 (N_1612,N_1504,N_1526);
nor U1613 (N_1613,N_1528,N_1565);
and U1614 (N_1614,N_1531,N_1549);
xor U1615 (N_1615,N_1531,N_1545);
nor U1616 (N_1616,N_1545,N_1551);
xor U1617 (N_1617,N_1559,N_1541);
and U1618 (N_1618,N_1561,N_1563);
and U1619 (N_1619,N_1546,N_1521);
nor U1620 (N_1620,N_1513,N_1548);
and U1621 (N_1621,N_1508,N_1533);
nor U1622 (N_1622,N_1557,N_1529);
nand U1623 (N_1623,N_1501,N_1540);
xnor U1624 (N_1624,N_1513,N_1571);
nand U1625 (N_1625,N_1509,N_1528);
nor U1626 (N_1626,N_1532,N_1528);
nor U1627 (N_1627,N_1544,N_1515);
or U1628 (N_1628,N_1560,N_1515);
xnor U1629 (N_1629,N_1566,N_1559);
or U1630 (N_1630,N_1507,N_1544);
or U1631 (N_1631,N_1533,N_1521);
and U1632 (N_1632,N_1512,N_1528);
and U1633 (N_1633,N_1532,N_1543);
and U1634 (N_1634,N_1530,N_1552);
and U1635 (N_1635,N_1516,N_1532);
or U1636 (N_1636,N_1523,N_1552);
nor U1637 (N_1637,N_1511,N_1570);
nor U1638 (N_1638,N_1503,N_1544);
nand U1639 (N_1639,N_1551,N_1564);
or U1640 (N_1640,N_1539,N_1546);
xor U1641 (N_1641,N_1559,N_1572);
or U1642 (N_1642,N_1538,N_1533);
and U1643 (N_1643,N_1556,N_1533);
and U1644 (N_1644,N_1539,N_1520);
and U1645 (N_1645,N_1531,N_1507);
and U1646 (N_1646,N_1538,N_1530);
xnor U1647 (N_1647,N_1544,N_1522);
xor U1648 (N_1648,N_1505,N_1554);
and U1649 (N_1649,N_1544,N_1548);
and U1650 (N_1650,N_1612,N_1646);
xnor U1651 (N_1651,N_1649,N_1595);
or U1652 (N_1652,N_1637,N_1613);
and U1653 (N_1653,N_1580,N_1620);
and U1654 (N_1654,N_1586,N_1633);
nor U1655 (N_1655,N_1624,N_1594);
xor U1656 (N_1656,N_1575,N_1607);
and U1657 (N_1657,N_1577,N_1644);
xnor U1658 (N_1658,N_1626,N_1584);
xor U1659 (N_1659,N_1603,N_1629);
or U1660 (N_1660,N_1601,N_1632);
xor U1661 (N_1661,N_1581,N_1636);
or U1662 (N_1662,N_1605,N_1648);
or U1663 (N_1663,N_1588,N_1639);
and U1664 (N_1664,N_1641,N_1587);
nor U1665 (N_1665,N_1578,N_1596);
nand U1666 (N_1666,N_1614,N_1642);
nor U1667 (N_1667,N_1608,N_1582);
xnor U1668 (N_1668,N_1617,N_1635);
nor U1669 (N_1669,N_1597,N_1623);
xor U1670 (N_1670,N_1602,N_1627);
nand U1671 (N_1671,N_1600,N_1610);
xor U1672 (N_1672,N_1583,N_1579);
or U1673 (N_1673,N_1634,N_1593);
nand U1674 (N_1674,N_1609,N_1589);
nor U1675 (N_1675,N_1592,N_1604);
and U1676 (N_1676,N_1599,N_1606);
or U1677 (N_1677,N_1618,N_1619);
nor U1678 (N_1678,N_1640,N_1628);
nor U1679 (N_1679,N_1643,N_1576);
nand U1680 (N_1680,N_1616,N_1598);
xor U1681 (N_1681,N_1615,N_1621);
or U1682 (N_1682,N_1625,N_1631);
and U1683 (N_1683,N_1638,N_1622);
or U1684 (N_1684,N_1647,N_1590);
or U1685 (N_1685,N_1591,N_1611);
nor U1686 (N_1686,N_1645,N_1585);
xor U1687 (N_1687,N_1630,N_1621);
nor U1688 (N_1688,N_1648,N_1586);
nor U1689 (N_1689,N_1610,N_1609);
nand U1690 (N_1690,N_1648,N_1607);
nand U1691 (N_1691,N_1595,N_1606);
nand U1692 (N_1692,N_1635,N_1641);
xor U1693 (N_1693,N_1621,N_1632);
nor U1694 (N_1694,N_1646,N_1584);
nor U1695 (N_1695,N_1580,N_1612);
xnor U1696 (N_1696,N_1584,N_1577);
xnor U1697 (N_1697,N_1645,N_1641);
nor U1698 (N_1698,N_1583,N_1601);
xor U1699 (N_1699,N_1634,N_1622);
nand U1700 (N_1700,N_1625,N_1602);
or U1701 (N_1701,N_1595,N_1593);
nor U1702 (N_1702,N_1629,N_1590);
nor U1703 (N_1703,N_1633,N_1628);
xnor U1704 (N_1704,N_1590,N_1589);
nor U1705 (N_1705,N_1586,N_1593);
nor U1706 (N_1706,N_1586,N_1592);
and U1707 (N_1707,N_1619,N_1605);
nor U1708 (N_1708,N_1635,N_1578);
and U1709 (N_1709,N_1588,N_1583);
nor U1710 (N_1710,N_1628,N_1581);
xnor U1711 (N_1711,N_1609,N_1643);
nor U1712 (N_1712,N_1602,N_1632);
or U1713 (N_1713,N_1637,N_1642);
and U1714 (N_1714,N_1605,N_1585);
xnor U1715 (N_1715,N_1583,N_1593);
xor U1716 (N_1716,N_1593,N_1637);
nand U1717 (N_1717,N_1614,N_1593);
or U1718 (N_1718,N_1649,N_1633);
xor U1719 (N_1719,N_1615,N_1647);
xnor U1720 (N_1720,N_1628,N_1638);
nand U1721 (N_1721,N_1584,N_1640);
or U1722 (N_1722,N_1601,N_1589);
nor U1723 (N_1723,N_1625,N_1610);
nor U1724 (N_1724,N_1609,N_1601);
nand U1725 (N_1725,N_1658,N_1702);
nand U1726 (N_1726,N_1696,N_1720);
nor U1727 (N_1727,N_1690,N_1667);
and U1728 (N_1728,N_1695,N_1704);
nor U1729 (N_1729,N_1652,N_1677);
or U1730 (N_1730,N_1689,N_1723);
or U1731 (N_1731,N_1669,N_1706);
nand U1732 (N_1732,N_1709,N_1711);
nor U1733 (N_1733,N_1674,N_1694);
and U1734 (N_1734,N_1676,N_1680);
and U1735 (N_1735,N_1661,N_1666);
or U1736 (N_1736,N_1668,N_1697);
nor U1737 (N_1737,N_1700,N_1718);
and U1738 (N_1738,N_1651,N_1664);
xor U1739 (N_1739,N_1708,N_1698);
or U1740 (N_1740,N_1688,N_1654);
nor U1741 (N_1741,N_1692,N_1671);
nand U1742 (N_1742,N_1693,N_1660);
xnor U1743 (N_1743,N_1717,N_1707);
nand U1744 (N_1744,N_1679,N_1650);
or U1745 (N_1745,N_1653,N_1670);
xnor U1746 (N_1746,N_1710,N_1724);
nand U1747 (N_1747,N_1713,N_1673);
and U1748 (N_1748,N_1687,N_1683);
nand U1749 (N_1749,N_1715,N_1681);
and U1750 (N_1750,N_1656,N_1685);
and U1751 (N_1751,N_1712,N_1657);
xor U1752 (N_1752,N_1659,N_1678);
nor U1753 (N_1753,N_1686,N_1672);
nand U1754 (N_1754,N_1701,N_1662);
or U1755 (N_1755,N_1703,N_1699);
xor U1756 (N_1756,N_1684,N_1655);
nand U1757 (N_1757,N_1721,N_1705);
nand U1758 (N_1758,N_1663,N_1719);
xor U1759 (N_1759,N_1665,N_1714);
and U1760 (N_1760,N_1716,N_1722);
nand U1761 (N_1761,N_1675,N_1691);
xnor U1762 (N_1762,N_1682,N_1689);
or U1763 (N_1763,N_1674,N_1721);
nand U1764 (N_1764,N_1686,N_1660);
nor U1765 (N_1765,N_1652,N_1670);
xnor U1766 (N_1766,N_1717,N_1688);
nor U1767 (N_1767,N_1700,N_1693);
xnor U1768 (N_1768,N_1719,N_1724);
xnor U1769 (N_1769,N_1711,N_1707);
xnor U1770 (N_1770,N_1674,N_1711);
and U1771 (N_1771,N_1702,N_1679);
or U1772 (N_1772,N_1700,N_1698);
or U1773 (N_1773,N_1722,N_1676);
xnor U1774 (N_1774,N_1718,N_1694);
xor U1775 (N_1775,N_1659,N_1723);
or U1776 (N_1776,N_1683,N_1685);
nand U1777 (N_1777,N_1704,N_1698);
or U1778 (N_1778,N_1711,N_1719);
xnor U1779 (N_1779,N_1718,N_1714);
nor U1780 (N_1780,N_1678,N_1666);
xor U1781 (N_1781,N_1699,N_1701);
xor U1782 (N_1782,N_1696,N_1669);
xnor U1783 (N_1783,N_1703,N_1707);
and U1784 (N_1784,N_1683,N_1711);
nor U1785 (N_1785,N_1653,N_1682);
and U1786 (N_1786,N_1657,N_1659);
xnor U1787 (N_1787,N_1669,N_1675);
nor U1788 (N_1788,N_1652,N_1702);
xor U1789 (N_1789,N_1711,N_1682);
nor U1790 (N_1790,N_1658,N_1662);
nand U1791 (N_1791,N_1702,N_1723);
nor U1792 (N_1792,N_1681,N_1661);
nand U1793 (N_1793,N_1653,N_1680);
nand U1794 (N_1794,N_1663,N_1699);
xor U1795 (N_1795,N_1650,N_1685);
or U1796 (N_1796,N_1682,N_1710);
xor U1797 (N_1797,N_1667,N_1719);
and U1798 (N_1798,N_1687,N_1689);
xnor U1799 (N_1799,N_1663,N_1661);
xnor U1800 (N_1800,N_1782,N_1760);
nand U1801 (N_1801,N_1728,N_1750);
or U1802 (N_1802,N_1764,N_1795);
nand U1803 (N_1803,N_1729,N_1758);
and U1804 (N_1804,N_1786,N_1756);
nand U1805 (N_1805,N_1791,N_1743);
and U1806 (N_1806,N_1734,N_1772);
nor U1807 (N_1807,N_1735,N_1761);
nand U1808 (N_1808,N_1778,N_1773);
nor U1809 (N_1809,N_1789,N_1780);
or U1810 (N_1810,N_1794,N_1770);
nand U1811 (N_1811,N_1769,N_1781);
or U1812 (N_1812,N_1749,N_1744);
xnor U1813 (N_1813,N_1792,N_1788);
xnor U1814 (N_1814,N_1790,N_1741);
or U1815 (N_1815,N_1768,N_1774);
nor U1816 (N_1816,N_1751,N_1762);
or U1817 (N_1817,N_1745,N_1757);
or U1818 (N_1818,N_1731,N_1733);
and U1819 (N_1819,N_1763,N_1759);
nand U1820 (N_1820,N_1784,N_1775);
xor U1821 (N_1821,N_1736,N_1740);
and U1822 (N_1822,N_1730,N_1746);
xor U1823 (N_1823,N_1765,N_1752);
nor U1824 (N_1824,N_1799,N_1783);
nand U1825 (N_1825,N_1771,N_1726);
or U1826 (N_1826,N_1755,N_1747);
and U1827 (N_1827,N_1754,N_1797);
nor U1828 (N_1828,N_1738,N_1732);
nor U1829 (N_1829,N_1737,N_1796);
or U1830 (N_1830,N_1727,N_1787);
and U1831 (N_1831,N_1739,N_1785);
and U1832 (N_1832,N_1725,N_1776);
or U1833 (N_1833,N_1793,N_1767);
xor U1834 (N_1834,N_1777,N_1798);
nand U1835 (N_1835,N_1766,N_1748);
xor U1836 (N_1836,N_1779,N_1753);
nor U1837 (N_1837,N_1742,N_1751);
or U1838 (N_1838,N_1741,N_1746);
xnor U1839 (N_1839,N_1768,N_1795);
or U1840 (N_1840,N_1742,N_1790);
nor U1841 (N_1841,N_1786,N_1788);
or U1842 (N_1842,N_1725,N_1755);
and U1843 (N_1843,N_1739,N_1763);
xor U1844 (N_1844,N_1792,N_1740);
or U1845 (N_1845,N_1749,N_1731);
xor U1846 (N_1846,N_1734,N_1774);
and U1847 (N_1847,N_1785,N_1799);
nand U1848 (N_1848,N_1777,N_1772);
nand U1849 (N_1849,N_1799,N_1731);
nand U1850 (N_1850,N_1752,N_1756);
xnor U1851 (N_1851,N_1768,N_1781);
or U1852 (N_1852,N_1763,N_1769);
nand U1853 (N_1853,N_1796,N_1756);
and U1854 (N_1854,N_1730,N_1788);
xnor U1855 (N_1855,N_1777,N_1739);
nand U1856 (N_1856,N_1748,N_1774);
and U1857 (N_1857,N_1763,N_1789);
nor U1858 (N_1858,N_1752,N_1746);
xnor U1859 (N_1859,N_1783,N_1787);
nor U1860 (N_1860,N_1783,N_1734);
nand U1861 (N_1861,N_1748,N_1764);
xor U1862 (N_1862,N_1757,N_1746);
nor U1863 (N_1863,N_1783,N_1738);
nor U1864 (N_1864,N_1727,N_1743);
nand U1865 (N_1865,N_1755,N_1786);
nor U1866 (N_1866,N_1770,N_1732);
nand U1867 (N_1867,N_1797,N_1774);
or U1868 (N_1868,N_1782,N_1727);
nand U1869 (N_1869,N_1782,N_1791);
or U1870 (N_1870,N_1740,N_1757);
nor U1871 (N_1871,N_1767,N_1783);
xnor U1872 (N_1872,N_1783,N_1745);
and U1873 (N_1873,N_1745,N_1785);
or U1874 (N_1874,N_1790,N_1734);
and U1875 (N_1875,N_1827,N_1866);
nor U1876 (N_1876,N_1839,N_1804);
or U1877 (N_1877,N_1832,N_1823);
xnor U1878 (N_1878,N_1869,N_1801);
nor U1879 (N_1879,N_1857,N_1851);
nor U1880 (N_1880,N_1873,N_1860);
nand U1881 (N_1881,N_1816,N_1813);
or U1882 (N_1882,N_1824,N_1855);
xnor U1883 (N_1883,N_1803,N_1850);
and U1884 (N_1884,N_1829,N_1843);
nor U1885 (N_1885,N_1854,N_1830);
and U1886 (N_1886,N_1814,N_1806);
nor U1887 (N_1887,N_1809,N_1822);
nand U1888 (N_1888,N_1818,N_1858);
or U1889 (N_1889,N_1862,N_1871);
nand U1890 (N_1890,N_1874,N_1800);
xnor U1891 (N_1891,N_1828,N_1872);
xor U1892 (N_1892,N_1826,N_1825);
or U1893 (N_1893,N_1837,N_1810);
or U1894 (N_1894,N_1867,N_1838);
or U1895 (N_1895,N_1859,N_1841);
nor U1896 (N_1896,N_1836,N_1835);
or U1897 (N_1897,N_1847,N_1834);
xnor U1898 (N_1898,N_1852,N_1856);
nand U1899 (N_1899,N_1846,N_1808);
and U1900 (N_1900,N_1865,N_1807);
nor U1901 (N_1901,N_1820,N_1833);
or U1902 (N_1902,N_1848,N_1863);
or U1903 (N_1903,N_1868,N_1845);
and U1904 (N_1904,N_1831,N_1819);
and U1905 (N_1905,N_1849,N_1840);
or U1906 (N_1906,N_1870,N_1802);
nand U1907 (N_1907,N_1821,N_1815);
xnor U1908 (N_1908,N_1805,N_1812);
nand U1909 (N_1909,N_1842,N_1861);
and U1910 (N_1910,N_1864,N_1844);
xnor U1911 (N_1911,N_1853,N_1817);
nor U1912 (N_1912,N_1811,N_1872);
nand U1913 (N_1913,N_1821,N_1830);
and U1914 (N_1914,N_1827,N_1819);
and U1915 (N_1915,N_1805,N_1811);
xnor U1916 (N_1916,N_1853,N_1841);
or U1917 (N_1917,N_1847,N_1869);
and U1918 (N_1918,N_1849,N_1869);
nor U1919 (N_1919,N_1834,N_1801);
xnor U1920 (N_1920,N_1829,N_1834);
xor U1921 (N_1921,N_1861,N_1808);
nor U1922 (N_1922,N_1865,N_1838);
nand U1923 (N_1923,N_1806,N_1831);
nor U1924 (N_1924,N_1805,N_1826);
xnor U1925 (N_1925,N_1824,N_1856);
xnor U1926 (N_1926,N_1803,N_1802);
nand U1927 (N_1927,N_1825,N_1803);
or U1928 (N_1928,N_1849,N_1826);
xnor U1929 (N_1929,N_1863,N_1849);
nor U1930 (N_1930,N_1825,N_1859);
or U1931 (N_1931,N_1817,N_1850);
or U1932 (N_1932,N_1806,N_1853);
or U1933 (N_1933,N_1826,N_1807);
nand U1934 (N_1934,N_1848,N_1871);
and U1935 (N_1935,N_1804,N_1821);
or U1936 (N_1936,N_1824,N_1826);
or U1937 (N_1937,N_1857,N_1805);
and U1938 (N_1938,N_1802,N_1840);
or U1939 (N_1939,N_1842,N_1864);
nor U1940 (N_1940,N_1854,N_1807);
xnor U1941 (N_1941,N_1804,N_1807);
nand U1942 (N_1942,N_1869,N_1865);
nand U1943 (N_1943,N_1806,N_1866);
nand U1944 (N_1944,N_1833,N_1852);
nor U1945 (N_1945,N_1828,N_1870);
and U1946 (N_1946,N_1827,N_1822);
nand U1947 (N_1947,N_1850,N_1859);
nor U1948 (N_1948,N_1801,N_1866);
or U1949 (N_1949,N_1864,N_1814);
xnor U1950 (N_1950,N_1890,N_1896);
and U1951 (N_1951,N_1941,N_1948);
nor U1952 (N_1952,N_1921,N_1906);
xnor U1953 (N_1953,N_1909,N_1936);
or U1954 (N_1954,N_1884,N_1926);
nand U1955 (N_1955,N_1946,N_1939);
or U1956 (N_1956,N_1891,N_1893);
nor U1957 (N_1957,N_1930,N_1935);
nand U1958 (N_1958,N_1897,N_1875);
or U1959 (N_1959,N_1886,N_1882);
xor U1960 (N_1960,N_1892,N_1917);
nor U1961 (N_1961,N_1878,N_1915);
xor U1962 (N_1962,N_1889,N_1913);
and U1963 (N_1963,N_1880,N_1914);
xor U1964 (N_1964,N_1901,N_1883);
nand U1965 (N_1965,N_1931,N_1898);
nand U1966 (N_1966,N_1877,N_1944);
nor U1967 (N_1967,N_1942,N_1933);
xnor U1968 (N_1968,N_1919,N_1932);
and U1969 (N_1969,N_1900,N_1902);
nand U1970 (N_1970,N_1904,N_1949);
xor U1971 (N_1971,N_1940,N_1929);
or U1972 (N_1972,N_1905,N_1922);
nand U1973 (N_1973,N_1899,N_1907);
xor U1974 (N_1974,N_1887,N_1938);
or U1975 (N_1975,N_1895,N_1934);
xnor U1976 (N_1976,N_1920,N_1947);
and U1977 (N_1977,N_1894,N_1912);
and U1978 (N_1978,N_1923,N_1924);
and U1979 (N_1979,N_1888,N_1879);
nor U1980 (N_1980,N_1928,N_1945);
and U1981 (N_1981,N_1903,N_1916);
nand U1982 (N_1982,N_1943,N_1876);
nor U1983 (N_1983,N_1908,N_1918);
and U1984 (N_1984,N_1885,N_1881);
xnor U1985 (N_1985,N_1910,N_1911);
or U1986 (N_1986,N_1937,N_1925);
or U1987 (N_1987,N_1927,N_1890);
or U1988 (N_1988,N_1883,N_1899);
nor U1989 (N_1989,N_1875,N_1913);
xor U1990 (N_1990,N_1876,N_1883);
nand U1991 (N_1991,N_1891,N_1879);
nand U1992 (N_1992,N_1891,N_1880);
nor U1993 (N_1993,N_1883,N_1904);
nor U1994 (N_1994,N_1915,N_1917);
xnor U1995 (N_1995,N_1919,N_1891);
xnor U1996 (N_1996,N_1937,N_1949);
or U1997 (N_1997,N_1896,N_1894);
and U1998 (N_1998,N_1930,N_1903);
or U1999 (N_1999,N_1948,N_1883);
or U2000 (N_2000,N_1890,N_1911);
nand U2001 (N_2001,N_1912,N_1902);
nand U2002 (N_2002,N_1904,N_1942);
xor U2003 (N_2003,N_1899,N_1935);
nand U2004 (N_2004,N_1896,N_1933);
xor U2005 (N_2005,N_1909,N_1876);
and U2006 (N_2006,N_1901,N_1910);
xor U2007 (N_2007,N_1898,N_1896);
xnor U2008 (N_2008,N_1917,N_1931);
and U2009 (N_2009,N_1943,N_1889);
xnor U2010 (N_2010,N_1935,N_1902);
xnor U2011 (N_2011,N_1932,N_1907);
nand U2012 (N_2012,N_1898,N_1944);
nor U2013 (N_2013,N_1925,N_1916);
or U2014 (N_2014,N_1898,N_1877);
xor U2015 (N_2015,N_1916,N_1936);
xnor U2016 (N_2016,N_1933,N_1900);
or U2017 (N_2017,N_1881,N_1920);
nand U2018 (N_2018,N_1920,N_1902);
nand U2019 (N_2019,N_1944,N_1886);
nand U2020 (N_2020,N_1943,N_1883);
nand U2021 (N_2021,N_1945,N_1909);
xnor U2022 (N_2022,N_1913,N_1893);
and U2023 (N_2023,N_1934,N_1886);
nand U2024 (N_2024,N_1881,N_1890);
or U2025 (N_2025,N_1951,N_1996);
xnor U2026 (N_2026,N_1989,N_1966);
nand U2027 (N_2027,N_2017,N_1972);
or U2028 (N_2028,N_2007,N_1991);
or U2029 (N_2029,N_2008,N_1990);
and U2030 (N_2030,N_1988,N_1971);
nor U2031 (N_2031,N_1977,N_1955);
or U2032 (N_2032,N_2003,N_2020);
nand U2033 (N_2033,N_1998,N_1986);
nand U2034 (N_2034,N_1961,N_1994);
nand U2035 (N_2035,N_1992,N_1959);
nand U2036 (N_2036,N_1960,N_2018);
nand U2037 (N_2037,N_1987,N_1975);
nor U2038 (N_2038,N_1983,N_2024);
and U2039 (N_2039,N_1969,N_1993);
xor U2040 (N_2040,N_1997,N_2022);
xnor U2041 (N_2041,N_1973,N_1985);
or U2042 (N_2042,N_1967,N_1982);
and U2043 (N_2043,N_1965,N_1962);
nand U2044 (N_2044,N_1958,N_2010);
nand U2045 (N_2045,N_1957,N_1950);
or U2046 (N_2046,N_2014,N_2009);
xor U2047 (N_2047,N_1963,N_2021);
nor U2048 (N_2048,N_2001,N_2000);
or U2049 (N_2049,N_1974,N_1984);
nand U2050 (N_2050,N_1954,N_1995);
nand U2051 (N_2051,N_1953,N_2005);
nand U2052 (N_2052,N_1952,N_1999);
nor U2053 (N_2053,N_2016,N_1976);
nor U2054 (N_2054,N_2023,N_1980);
nand U2055 (N_2055,N_2019,N_2015);
xor U2056 (N_2056,N_1968,N_1981);
nor U2057 (N_2057,N_2013,N_2004);
or U2058 (N_2058,N_1978,N_2002);
nor U2059 (N_2059,N_2012,N_1979);
and U2060 (N_2060,N_1964,N_2011);
xor U2061 (N_2061,N_2006,N_1956);
xor U2062 (N_2062,N_1970,N_1962);
or U2063 (N_2063,N_2017,N_1954);
xor U2064 (N_2064,N_2003,N_1999);
xor U2065 (N_2065,N_1966,N_1996);
nand U2066 (N_2066,N_1965,N_1994);
nor U2067 (N_2067,N_1965,N_2013);
nand U2068 (N_2068,N_2011,N_2015);
nand U2069 (N_2069,N_1986,N_1989);
xnor U2070 (N_2070,N_1990,N_1980);
nor U2071 (N_2071,N_1980,N_1988);
xor U2072 (N_2072,N_2014,N_1973);
xor U2073 (N_2073,N_1991,N_1966);
or U2074 (N_2074,N_1953,N_2014);
nand U2075 (N_2075,N_1950,N_1979);
nor U2076 (N_2076,N_1952,N_2006);
nand U2077 (N_2077,N_1990,N_1965);
or U2078 (N_2078,N_1987,N_1960);
xor U2079 (N_2079,N_2011,N_2009);
nand U2080 (N_2080,N_2006,N_1974);
and U2081 (N_2081,N_2006,N_2024);
xnor U2082 (N_2082,N_1992,N_1960);
nor U2083 (N_2083,N_1972,N_2020);
or U2084 (N_2084,N_1966,N_2024);
or U2085 (N_2085,N_1952,N_1979);
xnor U2086 (N_2086,N_2024,N_1975);
or U2087 (N_2087,N_2017,N_2001);
xnor U2088 (N_2088,N_1988,N_1951);
xnor U2089 (N_2089,N_2021,N_1954);
nor U2090 (N_2090,N_1994,N_1960);
nor U2091 (N_2091,N_1992,N_1952);
nor U2092 (N_2092,N_1995,N_2005);
or U2093 (N_2093,N_1963,N_2011);
nand U2094 (N_2094,N_2001,N_1995);
and U2095 (N_2095,N_1990,N_1988);
xor U2096 (N_2096,N_2013,N_1998);
nor U2097 (N_2097,N_1987,N_2013);
xor U2098 (N_2098,N_1982,N_2022);
or U2099 (N_2099,N_2013,N_2019);
or U2100 (N_2100,N_2053,N_2096);
xor U2101 (N_2101,N_2078,N_2060);
and U2102 (N_2102,N_2047,N_2098);
nor U2103 (N_2103,N_2037,N_2055);
nand U2104 (N_2104,N_2065,N_2064);
xor U2105 (N_2105,N_2033,N_2049);
or U2106 (N_2106,N_2041,N_2044);
nor U2107 (N_2107,N_2029,N_2051);
or U2108 (N_2108,N_2067,N_2056);
or U2109 (N_2109,N_2089,N_2048);
nand U2110 (N_2110,N_2062,N_2081);
and U2111 (N_2111,N_2088,N_2076);
and U2112 (N_2112,N_2025,N_2063);
or U2113 (N_2113,N_2094,N_2027);
and U2114 (N_2114,N_2038,N_2045);
xor U2115 (N_2115,N_2034,N_2050);
nand U2116 (N_2116,N_2077,N_2040);
nor U2117 (N_2117,N_2087,N_2039);
nor U2118 (N_2118,N_2043,N_2071);
nand U2119 (N_2119,N_2035,N_2082);
or U2120 (N_2120,N_2046,N_2079);
and U2121 (N_2121,N_2099,N_2070);
nor U2122 (N_2122,N_2095,N_2073);
or U2123 (N_2123,N_2086,N_2092);
or U2124 (N_2124,N_2026,N_2042);
xor U2125 (N_2125,N_2097,N_2068);
xnor U2126 (N_2126,N_2090,N_2083);
nor U2127 (N_2127,N_2054,N_2061);
or U2128 (N_2128,N_2031,N_2058);
nand U2129 (N_2129,N_2059,N_2084);
and U2130 (N_2130,N_2066,N_2091);
nand U2131 (N_2131,N_2085,N_2032);
nand U2132 (N_2132,N_2036,N_2030);
and U2133 (N_2133,N_2069,N_2072);
nor U2134 (N_2134,N_2057,N_2080);
xnor U2135 (N_2135,N_2093,N_2028);
xor U2136 (N_2136,N_2075,N_2052);
nand U2137 (N_2137,N_2074,N_2080);
and U2138 (N_2138,N_2074,N_2094);
nand U2139 (N_2139,N_2047,N_2061);
nand U2140 (N_2140,N_2039,N_2071);
nor U2141 (N_2141,N_2075,N_2097);
nand U2142 (N_2142,N_2060,N_2068);
xor U2143 (N_2143,N_2048,N_2085);
and U2144 (N_2144,N_2031,N_2090);
or U2145 (N_2145,N_2091,N_2068);
nand U2146 (N_2146,N_2071,N_2098);
and U2147 (N_2147,N_2040,N_2085);
and U2148 (N_2148,N_2037,N_2031);
nand U2149 (N_2149,N_2026,N_2047);
and U2150 (N_2150,N_2031,N_2028);
and U2151 (N_2151,N_2061,N_2088);
nor U2152 (N_2152,N_2068,N_2083);
and U2153 (N_2153,N_2070,N_2071);
nand U2154 (N_2154,N_2094,N_2050);
nor U2155 (N_2155,N_2053,N_2074);
xnor U2156 (N_2156,N_2068,N_2087);
xnor U2157 (N_2157,N_2076,N_2097);
and U2158 (N_2158,N_2097,N_2030);
or U2159 (N_2159,N_2044,N_2063);
or U2160 (N_2160,N_2068,N_2040);
and U2161 (N_2161,N_2055,N_2081);
or U2162 (N_2162,N_2095,N_2099);
or U2163 (N_2163,N_2062,N_2078);
xor U2164 (N_2164,N_2042,N_2063);
nor U2165 (N_2165,N_2085,N_2025);
or U2166 (N_2166,N_2085,N_2030);
or U2167 (N_2167,N_2028,N_2030);
and U2168 (N_2168,N_2040,N_2056);
and U2169 (N_2169,N_2049,N_2063);
xor U2170 (N_2170,N_2028,N_2062);
xnor U2171 (N_2171,N_2048,N_2073);
xor U2172 (N_2172,N_2033,N_2079);
xnor U2173 (N_2173,N_2045,N_2028);
nor U2174 (N_2174,N_2066,N_2031);
nand U2175 (N_2175,N_2160,N_2107);
and U2176 (N_2176,N_2134,N_2115);
nor U2177 (N_2177,N_2123,N_2137);
nor U2178 (N_2178,N_2136,N_2120);
and U2179 (N_2179,N_2158,N_2147);
or U2180 (N_2180,N_2133,N_2174);
nor U2181 (N_2181,N_2172,N_2101);
xnor U2182 (N_2182,N_2148,N_2154);
xnor U2183 (N_2183,N_2152,N_2110);
or U2184 (N_2184,N_2143,N_2167);
xor U2185 (N_2185,N_2131,N_2135);
nand U2186 (N_2186,N_2125,N_2141);
and U2187 (N_2187,N_2103,N_2165);
xnor U2188 (N_2188,N_2171,N_2173);
nand U2189 (N_2189,N_2166,N_2170);
or U2190 (N_2190,N_2126,N_2128);
or U2191 (N_2191,N_2124,N_2109);
and U2192 (N_2192,N_2155,N_2100);
and U2193 (N_2193,N_2112,N_2168);
nor U2194 (N_2194,N_2104,N_2156);
and U2195 (N_2195,N_2138,N_2151);
or U2196 (N_2196,N_2102,N_2163);
xnor U2197 (N_2197,N_2108,N_2113);
and U2198 (N_2198,N_2116,N_2145);
nor U2199 (N_2199,N_2157,N_2106);
nand U2200 (N_2200,N_2139,N_2122);
and U2201 (N_2201,N_2162,N_2142);
and U2202 (N_2202,N_2117,N_2111);
xnor U2203 (N_2203,N_2130,N_2132);
and U2204 (N_2204,N_2129,N_2114);
and U2205 (N_2205,N_2149,N_2127);
nor U2206 (N_2206,N_2169,N_2150);
and U2207 (N_2207,N_2161,N_2146);
and U2208 (N_2208,N_2144,N_2159);
and U2209 (N_2209,N_2164,N_2118);
nor U2210 (N_2210,N_2119,N_2121);
nand U2211 (N_2211,N_2140,N_2153);
nor U2212 (N_2212,N_2105,N_2146);
nor U2213 (N_2213,N_2173,N_2141);
and U2214 (N_2214,N_2154,N_2157);
or U2215 (N_2215,N_2125,N_2171);
or U2216 (N_2216,N_2124,N_2101);
nand U2217 (N_2217,N_2140,N_2150);
nor U2218 (N_2218,N_2171,N_2135);
or U2219 (N_2219,N_2142,N_2123);
or U2220 (N_2220,N_2172,N_2133);
or U2221 (N_2221,N_2133,N_2102);
nand U2222 (N_2222,N_2168,N_2167);
and U2223 (N_2223,N_2149,N_2108);
nand U2224 (N_2224,N_2140,N_2128);
nor U2225 (N_2225,N_2161,N_2166);
or U2226 (N_2226,N_2132,N_2158);
or U2227 (N_2227,N_2147,N_2103);
xnor U2228 (N_2228,N_2151,N_2126);
xor U2229 (N_2229,N_2147,N_2128);
and U2230 (N_2230,N_2128,N_2103);
or U2231 (N_2231,N_2173,N_2118);
xnor U2232 (N_2232,N_2149,N_2169);
nor U2233 (N_2233,N_2150,N_2111);
nor U2234 (N_2234,N_2123,N_2152);
xnor U2235 (N_2235,N_2106,N_2142);
nor U2236 (N_2236,N_2167,N_2109);
nor U2237 (N_2237,N_2123,N_2112);
xor U2238 (N_2238,N_2169,N_2159);
and U2239 (N_2239,N_2163,N_2128);
xor U2240 (N_2240,N_2174,N_2144);
or U2241 (N_2241,N_2103,N_2119);
xnor U2242 (N_2242,N_2147,N_2146);
and U2243 (N_2243,N_2161,N_2130);
or U2244 (N_2244,N_2172,N_2116);
nor U2245 (N_2245,N_2171,N_2146);
or U2246 (N_2246,N_2103,N_2154);
xnor U2247 (N_2247,N_2139,N_2129);
nor U2248 (N_2248,N_2157,N_2104);
xor U2249 (N_2249,N_2174,N_2168);
nand U2250 (N_2250,N_2247,N_2206);
nor U2251 (N_2251,N_2198,N_2217);
nor U2252 (N_2252,N_2191,N_2235);
nand U2253 (N_2253,N_2200,N_2230);
nor U2254 (N_2254,N_2195,N_2240);
nand U2255 (N_2255,N_2189,N_2214);
and U2256 (N_2256,N_2221,N_2246);
nor U2257 (N_2257,N_2192,N_2176);
and U2258 (N_2258,N_2239,N_2218);
and U2259 (N_2259,N_2203,N_2222);
or U2260 (N_2260,N_2182,N_2234);
or U2261 (N_2261,N_2177,N_2197);
nand U2262 (N_2262,N_2181,N_2208);
or U2263 (N_2263,N_2201,N_2249);
nand U2264 (N_2264,N_2207,N_2187);
or U2265 (N_2265,N_2178,N_2224);
xor U2266 (N_2266,N_2216,N_2209);
nor U2267 (N_2267,N_2213,N_2244);
or U2268 (N_2268,N_2215,N_2236);
nand U2269 (N_2269,N_2185,N_2183);
or U2270 (N_2270,N_2180,N_2237);
or U2271 (N_2271,N_2229,N_2211);
xnor U2272 (N_2272,N_2232,N_2194);
nand U2273 (N_2273,N_2193,N_2202);
xor U2274 (N_2274,N_2199,N_2179);
or U2275 (N_2275,N_2205,N_2241);
and U2276 (N_2276,N_2243,N_2219);
or U2277 (N_2277,N_2242,N_2225);
or U2278 (N_2278,N_2175,N_2204);
or U2279 (N_2279,N_2212,N_2245);
xor U2280 (N_2280,N_2227,N_2186);
or U2281 (N_2281,N_2223,N_2228);
nand U2282 (N_2282,N_2238,N_2184);
nor U2283 (N_2283,N_2196,N_2210);
or U2284 (N_2284,N_2220,N_2190);
and U2285 (N_2285,N_2231,N_2248);
or U2286 (N_2286,N_2233,N_2226);
xnor U2287 (N_2287,N_2188,N_2179);
nor U2288 (N_2288,N_2235,N_2248);
xor U2289 (N_2289,N_2190,N_2191);
nor U2290 (N_2290,N_2198,N_2246);
nand U2291 (N_2291,N_2177,N_2205);
nor U2292 (N_2292,N_2232,N_2233);
and U2293 (N_2293,N_2198,N_2193);
and U2294 (N_2294,N_2218,N_2186);
nand U2295 (N_2295,N_2241,N_2178);
nor U2296 (N_2296,N_2234,N_2242);
and U2297 (N_2297,N_2189,N_2176);
and U2298 (N_2298,N_2210,N_2192);
nand U2299 (N_2299,N_2213,N_2188);
xor U2300 (N_2300,N_2191,N_2177);
xnor U2301 (N_2301,N_2222,N_2206);
and U2302 (N_2302,N_2184,N_2198);
or U2303 (N_2303,N_2211,N_2225);
or U2304 (N_2304,N_2194,N_2212);
nor U2305 (N_2305,N_2180,N_2176);
nor U2306 (N_2306,N_2235,N_2178);
nor U2307 (N_2307,N_2241,N_2189);
xor U2308 (N_2308,N_2197,N_2216);
and U2309 (N_2309,N_2234,N_2235);
or U2310 (N_2310,N_2207,N_2208);
and U2311 (N_2311,N_2248,N_2226);
or U2312 (N_2312,N_2202,N_2236);
or U2313 (N_2313,N_2202,N_2203);
nor U2314 (N_2314,N_2187,N_2218);
nor U2315 (N_2315,N_2243,N_2238);
and U2316 (N_2316,N_2241,N_2175);
or U2317 (N_2317,N_2205,N_2193);
and U2318 (N_2318,N_2211,N_2205);
nand U2319 (N_2319,N_2231,N_2234);
nand U2320 (N_2320,N_2209,N_2228);
and U2321 (N_2321,N_2193,N_2179);
and U2322 (N_2322,N_2206,N_2193);
nand U2323 (N_2323,N_2224,N_2226);
nand U2324 (N_2324,N_2245,N_2237);
or U2325 (N_2325,N_2268,N_2305);
nand U2326 (N_2326,N_2272,N_2323);
nor U2327 (N_2327,N_2308,N_2312);
or U2328 (N_2328,N_2321,N_2258);
nand U2329 (N_2329,N_2293,N_2299);
nand U2330 (N_2330,N_2252,N_2290);
and U2331 (N_2331,N_2263,N_2276);
nor U2332 (N_2332,N_2273,N_2298);
nor U2333 (N_2333,N_2288,N_2318);
nor U2334 (N_2334,N_2275,N_2316);
and U2335 (N_2335,N_2307,N_2253);
and U2336 (N_2336,N_2277,N_2314);
or U2337 (N_2337,N_2309,N_2281);
xnor U2338 (N_2338,N_2264,N_2267);
nand U2339 (N_2339,N_2301,N_2266);
xnor U2340 (N_2340,N_2296,N_2283);
or U2341 (N_2341,N_2262,N_2251);
and U2342 (N_2342,N_2285,N_2291);
xor U2343 (N_2343,N_2250,N_2287);
nand U2344 (N_2344,N_2292,N_2294);
or U2345 (N_2345,N_2297,N_2269);
or U2346 (N_2346,N_2303,N_2319);
nand U2347 (N_2347,N_2274,N_2256);
xor U2348 (N_2348,N_2320,N_2257);
and U2349 (N_2349,N_2300,N_2315);
or U2350 (N_2350,N_2295,N_2259);
nand U2351 (N_2351,N_2271,N_2313);
nor U2352 (N_2352,N_2311,N_2324);
nand U2353 (N_2353,N_2282,N_2284);
nand U2354 (N_2354,N_2270,N_2310);
nand U2355 (N_2355,N_2254,N_2265);
xor U2356 (N_2356,N_2279,N_2306);
and U2357 (N_2357,N_2302,N_2278);
nand U2358 (N_2358,N_2317,N_2255);
or U2359 (N_2359,N_2289,N_2304);
and U2360 (N_2360,N_2322,N_2260);
nor U2361 (N_2361,N_2286,N_2280);
and U2362 (N_2362,N_2261,N_2317);
and U2363 (N_2363,N_2294,N_2284);
nand U2364 (N_2364,N_2262,N_2290);
nand U2365 (N_2365,N_2269,N_2273);
and U2366 (N_2366,N_2270,N_2303);
and U2367 (N_2367,N_2308,N_2299);
nor U2368 (N_2368,N_2271,N_2316);
or U2369 (N_2369,N_2281,N_2290);
nor U2370 (N_2370,N_2252,N_2281);
xor U2371 (N_2371,N_2252,N_2322);
and U2372 (N_2372,N_2301,N_2285);
nor U2373 (N_2373,N_2311,N_2279);
xor U2374 (N_2374,N_2308,N_2251);
and U2375 (N_2375,N_2321,N_2251);
nand U2376 (N_2376,N_2286,N_2267);
or U2377 (N_2377,N_2302,N_2252);
or U2378 (N_2378,N_2265,N_2290);
nor U2379 (N_2379,N_2312,N_2257);
and U2380 (N_2380,N_2293,N_2284);
or U2381 (N_2381,N_2288,N_2291);
and U2382 (N_2382,N_2279,N_2307);
nor U2383 (N_2383,N_2267,N_2269);
or U2384 (N_2384,N_2268,N_2289);
nand U2385 (N_2385,N_2257,N_2300);
nor U2386 (N_2386,N_2265,N_2301);
or U2387 (N_2387,N_2306,N_2283);
xnor U2388 (N_2388,N_2252,N_2316);
or U2389 (N_2389,N_2301,N_2282);
xor U2390 (N_2390,N_2265,N_2323);
or U2391 (N_2391,N_2292,N_2267);
or U2392 (N_2392,N_2259,N_2264);
and U2393 (N_2393,N_2268,N_2285);
and U2394 (N_2394,N_2259,N_2293);
nand U2395 (N_2395,N_2283,N_2281);
nor U2396 (N_2396,N_2300,N_2265);
or U2397 (N_2397,N_2282,N_2274);
nand U2398 (N_2398,N_2260,N_2296);
xnor U2399 (N_2399,N_2284,N_2280);
xnor U2400 (N_2400,N_2382,N_2394);
nor U2401 (N_2401,N_2395,N_2381);
xnor U2402 (N_2402,N_2367,N_2327);
or U2403 (N_2403,N_2333,N_2376);
and U2404 (N_2404,N_2347,N_2391);
xor U2405 (N_2405,N_2358,N_2331);
nor U2406 (N_2406,N_2392,N_2325);
nor U2407 (N_2407,N_2326,N_2355);
and U2408 (N_2408,N_2328,N_2380);
xor U2409 (N_2409,N_2387,N_2332);
nand U2410 (N_2410,N_2372,N_2398);
nor U2411 (N_2411,N_2383,N_2384);
nand U2412 (N_2412,N_2349,N_2374);
and U2413 (N_2413,N_2359,N_2353);
nand U2414 (N_2414,N_2352,N_2345);
nand U2415 (N_2415,N_2385,N_2386);
and U2416 (N_2416,N_2341,N_2361);
xor U2417 (N_2417,N_2354,N_2368);
nor U2418 (N_2418,N_2390,N_2339);
or U2419 (N_2419,N_2343,N_2373);
or U2420 (N_2420,N_2337,N_2370);
nand U2421 (N_2421,N_2379,N_2336);
and U2422 (N_2422,N_2388,N_2362);
nor U2423 (N_2423,N_2365,N_2330);
nand U2424 (N_2424,N_2363,N_2356);
nor U2425 (N_2425,N_2360,N_2397);
xor U2426 (N_2426,N_2364,N_2340);
nor U2427 (N_2427,N_2357,N_2371);
or U2428 (N_2428,N_2346,N_2396);
and U2429 (N_2429,N_2348,N_2393);
nor U2430 (N_2430,N_2366,N_2389);
xor U2431 (N_2431,N_2378,N_2342);
or U2432 (N_2432,N_2350,N_2329);
and U2433 (N_2433,N_2399,N_2377);
nand U2434 (N_2434,N_2375,N_2351);
or U2435 (N_2435,N_2334,N_2369);
nor U2436 (N_2436,N_2344,N_2335);
nor U2437 (N_2437,N_2338,N_2391);
xor U2438 (N_2438,N_2357,N_2363);
xor U2439 (N_2439,N_2344,N_2382);
or U2440 (N_2440,N_2357,N_2374);
xor U2441 (N_2441,N_2336,N_2375);
and U2442 (N_2442,N_2328,N_2367);
and U2443 (N_2443,N_2354,N_2387);
or U2444 (N_2444,N_2345,N_2393);
and U2445 (N_2445,N_2365,N_2346);
nor U2446 (N_2446,N_2379,N_2399);
xor U2447 (N_2447,N_2359,N_2398);
xnor U2448 (N_2448,N_2377,N_2371);
nand U2449 (N_2449,N_2376,N_2355);
nor U2450 (N_2450,N_2335,N_2353);
xnor U2451 (N_2451,N_2330,N_2339);
nand U2452 (N_2452,N_2356,N_2382);
xor U2453 (N_2453,N_2351,N_2340);
and U2454 (N_2454,N_2337,N_2378);
nor U2455 (N_2455,N_2368,N_2344);
or U2456 (N_2456,N_2372,N_2333);
and U2457 (N_2457,N_2347,N_2350);
nand U2458 (N_2458,N_2327,N_2369);
xor U2459 (N_2459,N_2328,N_2396);
or U2460 (N_2460,N_2353,N_2390);
nor U2461 (N_2461,N_2398,N_2347);
or U2462 (N_2462,N_2379,N_2326);
or U2463 (N_2463,N_2384,N_2392);
or U2464 (N_2464,N_2327,N_2399);
xnor U2465 (N_2465,N_2337,N_2356);
and U2466 (N_2466,N_2374,N_2355);
nor U2467 (N_2467,N_2391,N_2328);
and U2468 (N_2468,N_2359,N_2349);
and U2469 (N_2469,N_2385,N_2369);
or U2470 (N_2470,N_2374,N_2373);
and U2471 (N_2471,N_2336,N_2398);
or U2472 (N_2472,N_2332,N_2347);
or U2473 (N_2473,N_2366,N_2347);
nand U2474 (N_2474,N_2359,N_2392);
or U2475 (N_2475,N_2463,N_2408);
nor U2476 (N_2476,N_2447,N_2459);
nor U2477 (N_2477,N_2427,N_2403);
nand U2478 (N_2478,N_2446,N_2467);
and U2479 (N_2479,N_2429,N_2416);
xnor U2480 (N_2480,N_2461,N_2462);
nand U2481 (N_2481,N_2425,N_2410);
nor U2482 (N_2482,N_2458,N_2434);
or U2483 (N_2483,N_2448,N_2472);
or U2484 (N_2484,N_2413,N_2424);
xnor U2485 (N_2485,N_2407,N_2473);
and U2486 (N_2486,N_2440,N_2449);
or U2487 (N_2487,N_2401,N_2450);
or U2488 (N_2488,N_2456,N_2460);
or U2489 (N_2489,N_2469,N_2468);
xnor U2490 (N_2490,N_2402,N_2406);
xnor U2491 (N_2491,N_2441,N_2474);
nor U2492 (N_2492,N_2444,N_2421);
and U2493 (N_2493,N_2404,N_2435);
and U2494 (N_2494,N_2465,N_2445);
xnor U2495 (N_2495,N_2418,N_2432);
nor U2496 (N_2496,N_2471,N_2420);
nor U2497 (N_2497,N_2431,N_2415);
and U2498 (N_2498,N_2442,N_2457);
nand U2499 (N_2499,N_2470,N_2439);
xor U2500 (N_2500,N_2422,N_2437);
xnor U2501 (N_2501,N_2433,N_2452);
nor U2502 (N_2502,N_2414,N_2453);
xor U2503 (N_2503,N_2411,N_2455);
nor U2504 (N_2504,N_2412,N_2409);
xnor U2505 (N_2505,N_2451,N_2417);
or U2506 (N_2506,N_2430,N_2405);
and U2507 (N_2507,N_2454,N_2423);
nand U2508 (N_2508,N_2443,N_2400);
or U2509 (N_2509,N_2436,N_2428);
nor U2510 (N_2510,N_2419,N_2438);
xor U2511 (N_2511,N_2426,N_2466);
nand U2512 (N_2512,N_2464,N_2412);
and U2513 (N_2513,N_2445,N_2410);
nand U2514 (N_2514,N_2422,N_2404);
xor U2515 (N_2515,N_2400,N_2473);
and U2516 (N_2516,N_2442,N_2459);
and U2517 (N_2517,N_2445,N_2471);
xor U2518 (N_2518,N_2474,N_2458);
nor U2519 (N_2519,N_2473,N_2455);
and U2520 (N_2520,N_2432,N_2404);
and U2521 (N_2521,N_2464,N_2465);
xnor U2522 (N_2522,N_2439,N_2446);
nand U2523 (N_2523,N_2450,N_2454);
or U2524 (N_2524,N_2450,N_2441);
xnor U2525 (N_2525,N_2439,N_2462);
xor U2526 (N_2526,N_2456,N_2455);
nor U2527 (N_2527,N_2473,N_2420);
and U2528 (N_2528,N_2405,N_2461);
nand U2529 (N_2529,N_2462,N_2402);
nand U2530 (N_2530,N_2422,N_2468);
and U2531 (N_2531,N_2405,N_2403);
or U2532 (N_2532,N_2465,N_2409);
or U2533 (N_2533,N_2422,N_2416);
or U2534 (N_2534,N_2428,N_2462);
and U2535 (N_2535,N_2416,N_2473);
and U2536 (N_2536,N_2456,N_2426);
xor U2537 (N_2537,N_2449,N_2461);
nand U2538 (N_2538,N_2421,N_2463);
nor U2539 (N_2539,N_2434,N_2423);
xor U2540 (N_2540,N_2425,N_2440);
and U2541 (N_2541,N_2428,N_2437);
xnor U2542 (N_2542,N_2465,N_2474);
and U2543 (N_2543,N_2443,N_2470);
nand U2544 (N_2544,N_2425,N_2402);
xnor U2545 (N_2545,N_2458,N_2442);
nand U2546 (N_2546,N_2452,N_2457);
or U2547 (N_2547,N_2455,N_2409);
xor U2548 (N_2548,N_2404,N_2453);
xnor U2549 (N_2549,N_2412,N_2415);
nand U2550 (N_2550,N_2540,N_2522);
or U2551 (N_2551,N_2491,N_2520);
or U2552 (N_2552,N_2490,N_2523);
nand U2553 (N_2553,N_2478,N_2497);
or U2554 (N_2554,N_2533,N_2546);
nor U2555 (N_2555,N_2531,N_2486);
nand U2556 (N_2556,N_2477,N_2510);
nand U2557 (N_2557,N_2492,N_2539);
xor U2558 (N_2558,N_2509,N_2541);
xnor U2559 (N_2559,N_2512,N_2537);
nor U2560 (N_2560,N_2521,N_2514);
nor U2561 (N_2561,N_2504,N_2544);
nor U2562 (N_2562,N_2515,N_2538);
or U2563 (N_2563,N_2495,N_2506);
and U2564 (N_2564,N_2547,N_2484);
and U2565 (N_2565,N_2487,N_2513);
xor U2566 (N_2566,N_2507,N_2517);
or U2567 (N_2567,N_2500,N_2488);
nor U2568 (N_2568,N_2516,N_2543);
or U2569 (N_2569,N_2524,N_2545);
nand U2570 (N_2570,N_2485,N_2528);
and U2571 (N_2571,N_2534,N_2505);
nand U2572 (N_2572,N_2493,N_2480);
xor U2573 (N_2573,N_2529,N_2535);
nor U2574 (N_2574,N_2525,N_2519);
nor U2575 (N_2575,N_2476,N_2502);
nor U2576 (N_2576,N_2503,N_2479);
and U2577 (N_2577,N_2489,N_2536);
nor U2578 (N_2578,N_2549,N_2501);
nand U2579 (N_2579,N_2494,N_2499);
nor U2580 (N_2580,N_2511,N_2482);
and U2581 (N_2581,N_2475,N_2481);
nand U2582 (N_2582,N_2508,N_2532);
nor U2583 (N_2583,N_2526,N_2542);
or U2584 (N_2584,N_2498,N_2527);
nand U2585 (N_2585,N_2483,N_2548);
nand U2586 (N_2586,N_2496,N_2518);
and U2587 (N_2587,N_2530,N_2525);
or U2588 (N_2588,N_2500,N_2516);
xnor U2589 (N_2589,N_2510,N_2512);
and U2590 (N_2590,N_2518,N_2520);
xor U2591 (N_2591,N_2498,N_2523);
or U2592 (N_2592,N_2515,N_2480);
nand U2593 (N_2593,N_2494,N_2544);
or U2594 (N_2594,N_2526,N_2497);
nand U2595 (N_2595,N_2506,N_2510);
or U2596 (N_2596,N_2483,N_2496);
xor U2597 (N_2597,N_2516,N_2508);
xor U2598 (N_2598,N_2536,N_2507);
nor U2599 (N_2599,N_2494,N_2525);
nor U2600 (N_2600,N_2516,N_2517);
or U2601 (N_2601,N_2539,N_2548);
nor U2602 (N_2602,N_2538,N_2478);
and U2603 (N_2603,N_2495,N_2479);
xnor U2604 (N_2604,N_2525,N_2524);
and U2605 (N_2605,N_2492,N_2528);
or U2606 (N_2606,N_2475,N_2492);
and U2607 (N_2607,N_2519,N_2500);
and U2608 (N_2608,N_2502,N_2534);
and U2609 (N_2609,N_2526,N_2544);
xnor U2610 (N_2610,N_2510,N_2496);
nor U2611 (N_2611,N_2503,N_2519);
nand U2612 (N_2612,N_2530,N_2542);
and U2613 (N_2613,N_2509,N_2502);
xnor U2614 (N_2614,N_2501,N_2512);
or U2615 (N_2615,N_2492,N_2477);
nand U2616 (N_2616,N_2495,N_2537);
xor U2617 (N_2617,N_2547,N_2496);
and U2618 (N_2618,N_2492,N_2493);
or U2619 (N_2619,N_2503,N_2533);
or U2620 (N_2620,N_2480,N_2523);
nand U2621 (N_2621,N_2535,N_2489);
nand U2622 (N_2622,N_2480,N_2487);
xnor U2623 (N_2623,N_2515,N_2528);
nor U2624 (N_2624,N_2481,N_2518);
or U2625 (N_2625,N_2583,N_2592);
or U2626 (N_2626,N_2607,N_2568);
nand U2627 (N_2627,N_2623,N_2553);
xnor U2628 (N_2628,N_2608,N_2579);
nand U2629 (N_2629,N_2560,N_2593);
xor U2630 (N_2630,N_2603,N_2591);
nor U2631 (N_2631,N_2580,N_2596);
nand U2632 (N_2632,N_2554,N_2588);
nand U2633 (N_2633,N_2597,N_2565);
or U2634 (N_2634,N_2599,N_2569);
and U2635 (N_2635,N_2563,N_2558);
and U2636 (N_2636,N_2616,N_2566);
nor U2637 (N_2637,N_2572,N_2550);
xnor U2638 (N_2638,N_2564,N_2556);
nand U2639 (N_2639,N_2587,N_2570);
xnor U2640 (N_2640,N_2606,N_2567);
nand U2641 (N_2641,N_2624,N_2590);
nand U2642 (N_2642,N_2552,N_2584);
or U2643 (N_2643,N_2600,N_2605);
and U2644 (N_2644,N_2609,N_2578);
and U2645 (N_2645,N_2586,N_2613);
nor U2646 (N_2646,N_2576,N_2612);
and U2647 (N_2647,N_2614,N_2601);
nand U2648 (N_2648,N_2557,N_2559);
and U2649 (N_2649,N_2575,N_2581);
and U2650 (N_2650,N_2622,N_2573);
xor U2651 (N_2651,N_2611,N_2602);
nor U2652 (N_2652,N_2619,N_2604);
or U2653 (N_2653,N_2562,N_2582);
nand U2654 (N_2654,N_2571,N_2551);
and U2655 (N_2655,N_2555,N_2589);
and U2656 (N_2656,N_2595,N_2617);
nand U2657 (N_2657,N_2620,N_2561);
or U2658 (N_2658,N_2610,N_2615);
and U2659 (N_2659,N_2574,N_2618);
nor U2660 (N_2660,N_2577,N_2621);
nand U2661 (N_2661,N_2594,N_2598);
nor U2662 (N_2662,N_2585,N_2575);
or U2663 (N_2663,N_2591,N_2553);
xor U2664 (N_2664,N_2603,N_2600);
nor U2665 (N_2665,N_2582,N_2615);
nand U2666 (N_2666,N_2618,N_2576);
or U2667 (N_2667,N_2566,N_2553);
and U2668 (N_2668,N_2612,N_2585);
nor U2669 (N_2669,N_2616,N_2619);
xor U2670 (N_2670,N_2589,N_2593);
xnor U2671 (N_2671,N_2563,N_2599);
nor U2672 (N_2672,N_2561,N_2556);
or U2673 (N_2673,N_2614,N_2604);
nand U2674 (N_2674,N_2569,N_2602);
nand U2675 (N_2675,N_2611,N_2567);
nand U2676 (N_2676,N_2586,N_2592);
xor U2677 (N_2677,N_2586,N_2582);
and U2678 (N_2678,N_2616,N_2599);
and U2679 (N_2679,N_2559,N_2589);
xnor U2680 (N_2680,N_2624,N_2605);
nand U2681 (N_2681,N_2582,N_2553);
nand U2682 (N_2682,N_2574,N_2551);
nand U2683 (N_2683,N_2572,N_2599);
and U2684 (N_2684,N_2558,N_2575);
and U2685 (N_2685,N_2605,N_2550);
or U2686 (N_2686,N_2616,N_2612);
and U2687 (N_2687,N_2624,N_2562);
nand U2688 (N_2688,N_2596,N_2599);
and U2689 (N_2689,N_2587,N_2556);
nor U2690 (N_2690,N_2554,N_2559);
or U2691 (N_2691,N_2584,N_2607);
xor U2692 (N_2692,N_2615,N_2572);
or U2693 (N_2693,N_2573,N_2569);
nand U2694 (N_2694,N_2564,N_2565);
xnor U2695 (N_2695,N_2609,N_2605);
nor U2696 (N_2696,N_2623,N_2581);
or U2697 (N_2697,N_2590,N_2564);
and U2698 (N_2698,N_2551,N_2623);
xor U2699 (N_2699,N_2573,N_2588);
and U2700 (N_2700,N_2679,N_2684);
nand U2701 (N_2701,N_2663,N_2668);
nor U2702 (N_2702,N_2625,N_2692);
nand U2703 (N_2703,N_2666,N_2658);
nor U2704 (N_2704,N_2657,N_2682);
nor U2705 (N_2705,N_2685,N_2687);
nor U2706 (N_2706,N_2676,N_2635);
xnor U2707 (N_2707,N_2675,N_2688);
xnor U2708 (N_2708,N_2695,N_2648);
nand U2709 (N_2709,N_2641,N_2698);
nand U2710 (N_2710,N_2645,N_2642);
nand U2711 (N_2711,N_2696,N_2671);
xor U2712 (N_2712,N_2652,N_2638);
or U2713 (N_2713,N_2636,N_2664);
nor U2714 (N_2714,N_2691,N_2689);
or U2715 (N_2715,N_2678,N_2697);
xor U2716 (N_2716,N_2660,N_2662);
nor U2717 (N_2717,N_2681,N_2665);
or U2718 (N_2718,N_2630,N_2653);
or U2719 (N_2719,N_2683,N_2654);
and U2720 (N_2720,N_2667,N_2644);
xnor U2721 (N_2721,N_2674,N_2647);
and U2722 (N_2722,N_2632,N_2661);
xor U2723 (N_2723,N_2656,N_2637);
and U2724 (N_2724,N_2650,N_2633);
nor U2725 (N_2725,N_2627,N_2694);
and U2726 (N_2726,N_2677,N_2651);
or U2727 (N_2727,N_2640,N_2672);
nor U2728 (N_2728,N_2631,N_2693);
nand U2729 (N_2729,N_2699,N_2659);
nor U2730 (N_2730,N_2649,N_2686);
nor U2731 (N_2731,N_2639,N_2634);
xor U2732 (N_2732,N_2680,N_2643);
or U2733 (N_2733,N_2655,N_2646);
and U2734 (N_2734,N_2670,N_2690);
nand U2735 (N_2735,N_2669,N_2673);
and U2736 (N_2736,N_2629,N_2626);
nor U2737 (N_2737,N_2628,N_2690);
or U2738 (N_2738,N_2633,N_2660);
xnor U2739 (N_2739,N_2643,N_2636);
or U2740 (N_2740,N_2692,N_2639);
or U2741 (N_2741,N_2678,N_2688);
xor U2742 (N_2742,N_2681,N_2685);
nor U2743 (N_2743,N_2650,N_2630);
or U2744 (N_2744,N_2670,N_2663);
nand U2745 (N_2745,N_2683,N_2627);
nand U2746 (N_2746,N_2650,N_2626);
xnor U2747 (N_2747,N_2666,N_2653);
and U2748 (N_2748,N_2689,N_2643);
nand U2749 (N_2749,N_2627,N_2635);
or U2750 (N_2750,N_2654,N_2666);
xnor U2751 (N_2751,N_2699,N_2686);
or U2752 (N_2752,N_2625,N_2693);
and U2753 (N_2753,N_2682,N_2694);
nor U2754 (N_2754,N_2669,N_2698);
xnor U2755 (N_2755,N_2666,N_2644);
nor U2756 (N_2756,N_2696,N_2673);
and U2757 (N_2757,N_2698,N_2629);
and U2758 (N_2758,N_2631,N_2688);
or U2759 (N_2759,N_2645,N_2691);
or U2760 (N_2760,N_2668,N_2677);
xor U2761 (N_2761,N_2695,N_2676);
nand U2762 (N_2762,N_2663,N_2654);
and U2763 (N_2763,N_2650,N_2662);
or U2764 (N_2764,N_2693,N_2646);
or U2765 (N_2765,N_2688,N_2661);
or U2766 (N_2766,N_2678,N_2651);
and U2767 (N_2767,N_2628,N_2669);
nand U2768 (N_2768,N_2646,N_2656);
nand U2769 (N_2769,N_2698,N_2633);
and U2770 (N_2770,N_2630,N_2628);
xor U2771 (N_2771,N_2666,N_2662);
xor U2772 (N_2772,N_2665,N_2698);
xor U2773 (N_2773,N_2681,N_2675);
xnor U2774 (N_2774,N_2637,N_2663);
and U2775 (N_2775,N_2740,N_2756);
xnor U2776 (N_2776,N_2726,N_2771);
xnor U2777 (N_2777,N_2750,N_2753);
or U2778 (N_2778,N_2734,N_2725);
nand U2779 (N_2779,N_2732,N_2737);
xnor U2780 (N_2780,N_2719,N_2754);
xor U2781 (N_2781,N_2745,N_2741);
nand U2782 (N_2782,N_2702,N_2724);
xnor U2783 (N_2783,N_2735,N_2765);
or U2784 (N_2784,N_2760,N_2711);
and U2785 (N_2785,N_2759,N_2723);
xor U2786 (N_2786,N_2703,N_2752);
or U2787 (N_2787,N_2769,N_2707);
xor U2788 (N_2788,N_2704,N_2717);
nand U2789 (N_2789,N_2772,N_2746);
nand U2790 (N_2790,N_2774,N_2710);
nor U2791 (N_2791,N_2716,N_2701);
nor U2792 (N_2792,N_2738,N_2705);
nor U2793 (N_2793,N_2763,N_2773);
xnor U2794 (N_2794,N_2721,N_2755);
nor U2795 (N_2795,N_2743,N_2764);
nand U2796 (N_2796,N_2714,N_2739);
nor U2797 (N_2797,N_2720,N_2748);
or U2798 (N_2798,N_2709,N_2713);
nor U2799 (N_2799,N_2728,N_2715);
nand U2800 (N_2800,N_2727,N_2731);
xnor U2801 (N_2801,N_2761,N_2722);
and U2802 (N_2802,N_2747,N_2736);
nor U2803 (N_2803,N_2749,N_2751);
or U2804 (N_2804,N_2708,N_2768);
xnor U2805 (N_2805,N_2770,N_2730);
nand U2806 (N_2806,N_2762,N_2766);
or U2807 (N_2807,N_2700,N_2742);
nor U2808 (N_2808,N_2712,N_2757);
nor U2809 (N_2809,N_2729,N_2733);
and U2810 (N_2810,N_2718,N_2706);
nand U2811 (N_2811,N_2767,N_2758);
and U2812 (N_2812,N_2744,N_2760);
xor U2813 (N_2813,N_2765,N_2720);
and U2814 (N_2814,N_2702,N_2723);
and U2815 (N_2815,N_2730,N_2766);
and U2816 (N_2816,N_2737,N_2702);
and U2817 (N_2817,N_2755,N_2752);
and U2818 (N_2818,N_2753,N_2720);
xnor U2819 (N_2819,N_2742,N_2753);
and U2820 (N_2820,N_2710,N_2715);
nor U2821 (N_2821,N_2710,N_2751);
nand U2822 (N_2822,N_2719,N_2710);
xnor U2823 (N_2823,N_2763,N_2727);
or U2824 (N_2824,N_2760,N_2725);
nor U2825 (N_2825,N_2732,N_2726);
and U2826 (N_2826,N_2749,N_2765);
nand U2827 (N_2827,N_2741,N_2759);
nor U2828 (N_2828,N_2760,N_2730);
xnor U2829 (N_2829,N_2719,N_2717);
nor U2830 (N_2830,N_2771,N_2765);
xor U2831 (N_2831,N_2751,N_2729);
xor U2832 (N_2832,N_2720,N_2702);
xor U2833 (N_2833,N_2746,N_2711);
or U2834 (N_2834,N_2722,N_2735);
nor U2835 (N_2835,N_2720,N_2727);
or U2836 (N_2836,N_2727,N_2735);
and U2837 (N_2837,N_2752,N_2758);
and U2838 (N_2838,N_2751,N_2742);
and U2839 (N_2839,N_2724,N_2725);
nor U2840 (N_2840,N_2765,N_2762);
nor U2841 (N_2841,N_2766,N_2738);
nor U2842 (N_2842,N_2735,N_2772);
and U2843 (N_2843,N_2736,N_2752);
xnor U2844 (N_2844,N_2773,N_2774);
xnor U2845 (N_2845,N_2749,N_2703);
or U2846 (N_2846,N_2752,N_2715);
and U2847 (N_2847,N_2745,N_2711);
xnor U2848 (N_2848,N_2767,N_2715);
nor U2849 (N_2849,N_2720,N_2728);
and U2850 (N_2850,N_2779,N_2809);
and U2851 (N_2851,N_2846,N_2844);
and U2852 (N_2852,N_2810,N_2806);
nand U2853 (N_2853,N_2789,N_2800);
nor U2854 (N_2854,N_2830,N_2781);
nor U2855 (N_2855,N_2802,N_2822);
xnor U2856 (N_2856,N_2834,N_2784);
or U2857 (N_2857,N_2796,N_2791);
and U2858 (N_2858,N_2795,N_2785);
or U2859 (N_2859,N_2821,N_2828);
and U2860 (N_2860,N_2788,N_2817);
xor U2861 (N_2861,N_2808,N_2835);
or U2862 (N_2862,N_2813,N_2783);
and U2863 (N_2863,N_2824,N_2838);
nand U2864 (N_2864,N_2807,N_2804);
xor U2865 (N_2865,N_2801,N_2820);
xor U2866 (N_2866,N_2840,N_2827);
nand U2867 (N_2867,N_2787,N_2793);
nand U2868 (N_2868,N_2776,N_2782);
nor U2869 (N_2869,N_2847,N_2797);
and U2870 (N_2870,N_2818,N_2836);
xor U2871 (N_2871,N_2805,N_2792);
xor U2872 (N_2872,N_2823,N_2837);
and U2873 (N_2873,N_2849,N_2842);
or U2874 (N_2874,N_2812,N_2794);
and U2875 (N_2875,N_2839,N_2829);
and U2876 (N_2876,N_2778,N_2832);
nor U2877 (N_2877,N_2841,N_2843);
nor U2878 (N_2878,N_2786,N_2819);
or U2879 (N_2879,N_2803,N_2775);
nor U2880 (N_2880,N_2848,N_2814);
and U2881 (N_2881,N_2815,N_2799);
nor U2882 (N_2882,N_2798,N_2831);
xor U2883 (N_2883,N_2811,N_2826);
nor U2884 (N_2884,N_2777,N_2816);
nor U2885 (N_2885,N_2833,N_2780);
and U2886 (N_2886,N_2825,N_2845);
xor U2887 (N_2887,N_2790,N_2831);
nand U2888 (N_2888,N_2822,N_2829);
nand U2889 (N_2889,N_2821,N_2793);
or U2890 (N_2890,N_2800,N_2819);
nor U2891 (N_2891,N_2836,N_2816);
nand U2892 (N_2892,N_2778,N_2801);
nor U2893 (N_2893,N_2822,N_2786);
nor U2894 (N_2894,N_2838,N_2804);
nor U2895 (N_2895,N_2798,N_2787);
nor U2896 (N_2896,N_2835,N_2789);
or U2897 (N_2897,N_2777,N_2791);
xor U2898 (N_2898,N_2801,N_2809);
and U2899 (N_2899,N_2838,N_2801);
nor U2900 (N_2900,N_2829,N_2778);
nor U2901 (N_2901,N_2834,N_2837);
nor U2902 (N_2902,N_2813,N_2841);
nand U2903 (N_2903,N_2805,N_2848);
nand U2904 (N_2904,N_2805,N_2784);
or U2905 (N_2905,N_2799,N_2840);
nand U2906 (N_2906,N_2780,N_2822);
xor U2907 (N_2907,N_2784,N_2833);
or U2908 (N_2908,N_2819,N_2803);
xor U2909 (N_2909,N_2844,N_2806);
or U2910 (N_2910,N_2787,N_2844);
and U2911 (N_2911,N_2779,N_2792);
xor U2912 (N_2912,N_2783,N_2845);
nor U2913 (N_2913,N_2820,N_2839);
nand U2914 (N_2914,N_2848,N_2842);
and U2915 (N_2915,N_2818,N_2809);
nand U2916 (N_2916,N_2842,N_2810);
or U2917 (N_2917,N_2785,N_2830);
nor U2918 (N_2918,N_2832,N_2795);
nand U2919 (N_2919,N_2838,N_2833);
or U2920 (N_2920,N_2809,N_2784);
or U2921 (N_2921,N_2814,N_2787);
nor U2922 (N_2922,N_2809,N_2847);
and U2923 (N_2923,N_2839,N_2778);
and U2924 (N_2924,N_2838,N_2780);
and U2925 (N_2925,N_2921,N_2857);
nand U2926 (N_2926,N_2909,N_2922);
and U2927 (N_2927,N_2856,N_2893);
or U2928 (N_2928,N_2883,N_2874);
nand U2929 (N_2929,N_2905,N_2903);
nor U2930 (N_2930,N_2898,N_2915);
and U2931 (N_2931,N_2855,N_2882);
nand U2932 (N_2932,N_2897,N_2864);
and U2933 (N_2933,N_2859,N_2850);
or U2934 (N_2934,N_2888,N_2891);
and U2935 (N_2935,N_2867,N_2881);
or U2936 (N_2936,N_2852,N_2853);
nand U2937 (N_2937,N_2912,N_2884);
nor U2938 (N_2938,N_2858,N_2911);
xor U2939 (N_2939,N_2873,N_2914);
or U2940 (N_2940,N_2923,N_2870);
xnor U2941 (N_2941,N_2904,N_2854);
and U2942 (N_2942,N_2916,N_2895);
nand U2943 (N_2943,N_2924,N_2868);
and U2944 (N_2944,N_2872,N_2863);
xnor U2945 (N_2945,N_2902,N_2918);
or U2946 (N_2946,N_2866,N_2878);
nand U2947 (N_2947,N_2900,N_2896);
and U2948 (N_2948,N_2890,N_2851);
and U2949 (N_2949,N_2869,N_2920);
nor U2950 (N_2950,N_2907,N_2879);
or U2951 (N_2951,N_2875,N_2901);
xor U2952 (N_2952,N_2892,N_2906);
xnor U2953 (N_2953,N_2876,N_2889);
or U2954 (N_2954,N_2871,N_2860);
nand U2955 (N_2955,N_2865,N_2886);
nand U2956 (N_2956,N_2861,N_2913);
nor U2957 (N_2957,N_2877,N_2894);
nor U2958 (N_2958,N_2910,N_2885);
or U2959 (N_2959,N_2887,N_2862);
and U2960 (N_2960,N_2917,N_2880);
nor U2961 (N_2961,N_2899,N_2919);
or U2962 (N_2962,N_2908,N_2892);
xor U2963 (N_2963,N_2892,N_2895);
xnor U2964 (N_2964,N_2888,N_2911);
or U2965 (N_2965,N_2883,N_2864);
or U2966 (N_2966,N_2864,N_2903);
and U2967 (N_2967,N_2892,N_2911);
nor U2968 (N_2968,N_2887,N_2850);
xnor U2969 (N_2969,N_2919,N_2920);
or U2970 (N_2970,N_2898,N_2872);
and U2971 (N_2971,N_2916,N_2906);
nor U2972 (N_2972,N_2910,N_2852);
nor U2973 (N_2973,N_2875,N_2899);
nor U2974 (N_2974,N_2873,N_2875);
or U2975 (N_2975,N_2869,N_2856);
and U2976 (N_2976,N_2910,N_2871);
nor U2977 (N_2977,N_2853,N_2867);
xnor U2978 (N_2978,N_2857,N_2887);
or U2979 (N_2979,N_2879,N_2904);
nand U2980 (N_2980,N_2855,N_2863);
and U2981 (N_2981,N_2867,N_2905);
or U2982 (N_2982,N_2879,N_2911);
nand U2983 (N_2983,N_2892,N_2918);
or U2984 (N_2984,N_2868,N_2908);
nand U2985 (N_2985,N_2920,N_2871);
nor U2986 (N_2986,N_2906,N_2851);
or U2987 (N_2987,N_2862,N_2875);
xor U2988 (N_2988,N_2903,N_2884);
xnor U2989 (N_2989,N_2923,N_2892);
and U2990 (N_2990,N_2888,N_2866);
or U2991 (N_2991,N_2881,N_2871);
or U2992 (N_2992,N_2906,N_2915);
xnor U2993 (N_2993,N_2911,N_2881);
and U2994 (N_2994,N_2924,N_2910);
nand U2995 (N_2995,N_2856,N_2909);
xnor U2996 (N_2996,N_2897,N_2875);
nor U2997 (N_2997,N_2864,N_2919);
nand U2998 (N_2998,N_2911,N_2917);
nor U2999 (N_2999,N_2854,N_2858);
nor UO_0 (O_0,N_2987,N_2990);
or UO_1 (O_1,N_2968,N_2936);
nor UO_2 (O_2,N_2945,N_2944);
nor UO_3 (O_3,N_2981,N_2982);
or UO_4 (O_4,N_2941,N_2980);
xor UO_5 (O_5,N_2985,N_2976);
or UO_6 (O_6,N_2940,N_2934);
nand UO_7 (O_7,N_2984,N_2973);
and UO_8 (O_8,N_2963,N_2933);
and UO_9 (O_9,N_2951,N_2932);
nand UO_10 (O_10,N_2986,N_2931);
nand UO_11 (O_11,N_2949,N_2966);
and UO_12 (O_12,N_2970,N_2978);
nand UO_13 (O_13,N_2955,N_2929);
xor UO_14 (O_14,N_2935,N_2959);
or UO_15 (O_15,N_2938,N_2926);
nor UO_16 (O_16,N_2954,N_2948);
nand UO_17 (O_17,N_2994,N_2977);
xnor UO_18 (O_18,N_2962,N_2939);
xor UO_19 (O_19,N_2956,N_2971);
nor UO_20 (O_20,N_2975,N_2988);
and UO_21 (O_21,N_2950,N_2965);
and UO_22 (O_22,N_2969,N_2958);
xor UO_23 (O_23,N_2952,N_2957);
or UO_24 (O_24,N_2996,N_2967);
and UO_25 (O_25,N_2997,N_2974);
nor UO_26 (O_26,N_2992,N_2991);
nand UO_27 (O_27,N_2961,N_2995);
and UO_28 (O_28,N_2930,N_2953);
nor UO_29 (O_29,N_2947,N_2943);
xnor UO_30 (O_30,N_2937,N_2972);
or UO_31 (O_31,N_2927,N_2993);
nand UO_32 (O_32,N_2989,N_2999);
and UO_33 (O_33,N_2964,N_2946);
or UO_34 (O_34,N_2979,N_2960);
nand UO_35 (O_35,N_2983,N_2928);
and UO_36 (O_36,N_2998,N_2942);
nand UO_37 (O_37,N_2925,N_2936);
and UO_38 (O_38,N_2975,N_2982);
or UO_39 (O_39,N_2926,N_2929);
xor UO_40 (O_40,N_2950,N_2939);
and UO_41 (O_41,N_2938,N_2970);
xor UO_42 (O_42,N_2928,N_2962);
and UO_43 (O_43,N_2979,N_2967);
nor UO_44 (O_44,N_2981,N_2954);
or UO_45 (O_45,N_2999,N_2969);
or UO_46 (O_46,N_2960,N_2942);
nor UO_47 (O_47,N_2960,N_2995);
nand UO_48 (O_48,N_2968,N_2987);
and UO_49 (O_49,N_2934,N_2965);
xor UO_50 (O_50,N_2965,N_2991);
nand UO_51 (O_51,N_2946,N_2985);
and UO_52 (O_52,N_2971,N_2936);
nand UO_53 (O_53,N_2969,N_2932);
nor UO_54 (O_54,N_2926,N_2997);
nor UO_55 (O_55,N_2980,N_2993);
or UO_56 (O_56,N_2988,N_2959);
and UO_57 (O_57,N_2991,N_2978);
or UO_58 (O_58,N_2934,N_2964);
nand UO_59 (O_59,N_2928,N_2926);
and UO_60 (O_60,N_2999,N_2932);
xnor UO_61 (O_61,N_2935,N_2974);
xor UO_62 (O_62,N_2928,N_2942);
xnor UO_63 (O_63,N_2979,N_2961);
and UO_64 (O_64,N_2999,N_2978);
nand UO_65 (O_65,N_2952,N_2987);
or UO_66 (O_66,N_2987,N_2960);
xor UO_67 (O_67,N_2967,N_2977);
and UO_68 (O_68,N_2944,N_2980);
xor UO_69 (O_69,N_2938,N_2986);
nand UO_70 (O_70,N_2972,N_2945);
and UO_71 (O_71,N_2929,N_2945);
and UO_72 (O_72,N_2981,N_2936);
or UO_73 (O_73,N_2944,N_2963);
nand UO_74 (O_74,N_2938,N_2952);
or UO_75 (O_75,N_2944,N_2928);
and UO_76 (O_76,N_2947,N_2983);
nand UO_77 (O_77,N_2985,N_2996);
and UO_78 (O_78,N_2960,N_2990);
or UO_79 (O_79,N_2926,N_2944);
xor UO_80 (O_80,N_2999,N_2972);
and UO_81 (O_81,N_2977,N_2943);
nand UO_82 (O_82,N_2980,N_2973);
xnor UO_83 (O_83,N_2929,N_2976);
or UO_84 (O_84,N_2937,N_2933);
nand UO_85 (O_85,N_2942,N_2956);
nor UO_86 (O_86,N_2962,N_2987);
xnor UO_87 (O_87,N_2950,N_2958);
and UO_88 (O_88,N_2954,N_2926);
xnor UO_89 (O_89,N_2934,N_2932);
xnor UO_90 (O_90,N_2944,N_2930);
and UO_91 (O_91,N_2956,N_2958);
or UO_92 (O_92,N_2927,N_2938);
nand UO_93 (O_93,N_2982,N_2959);
or UO_94 (O_94,N_2981,N_2987);
xnor UO_95 (O_95,N_2975,N_2956);
and UO_96 (O_96,N_2990,N_2936);
nor UO_97 (O_97,N_2965,N_2959);
xnor UO_98 (O_98,N_2974,N_2936);
nor UO_99 (O_99,N_2950,N_2925);
xor UO_100 (O_100,N_2927,N_2948);
and UO_101 (O_101,N_2934,N_2943);
or UO_102 (O_102,N_2955,N_2949);
or UO_103 (O_103,N_2928,N_2977);
or UO_104 (O_104,N_2943,N_2946);
or UO_105 (O_105,N_2963,N_2980);
nor UO_106 (O_106,N_2993,N_2960);
or UO_107 (O_107,N_2980,N_2962);
and UO_108 (O_108,N_2978,N_2926);
xnor UO_109 (O_109,N_2949,N_2984);
xor UO_110 (O_110,N_2952,N_2966);
nand UO_111 (O_111,N_2937,N_2968);
nor UO_112 (O_112,N_2926,N_2975);
xnor UO_113 (O_113,N_2942,N_2949);
nor UO_114 (O_114,N_2990,N_2946);
and UO_115 (O_115,N_2958,N_2954);
nor UO_116 (O_116,N_2976,N_2925);
nor UO_117 (O_117,N_2945,N_2994);
nand UO_118 (O_118,N_2981,N_2951);
nand UO_119 (O_119,N_2963,N_2964);
or UO_120 (O_120,N_2989,N_2982);
xor UO_121 (O_121,N_2947,N_2932);
or UO_122 (O_122,N_2942,N_2953);
nand UO_123 (O_123,N_2995,N_2943);
and UO_124 (O_124,N_2993,N_2995);
and UO_125 (O_125,N_2988,N_2931);
or UO_126 (O_126,N_2960,N_2989);
nor UO_127 (O_127,N_2963,N_2971);
xnor UO_128 (O_128,N_2995,N_2967);
or UO_129 (O_129,N_2996,N_2979);
nand UO_130 (O_130,N_2987,N_2991);
or UO_131 (O_131,N_2969,N_2962);
nand UO_132 (O_132,N_2996,N_2968);
and UO_133 (O_133,N_2954,N_2956);
xor UO_134 (O_134,N_2946,N_2997);
or UO_135 (O_135,N_2950,N_2974);
nand UO_136 (O_136,N_2956,N_2995);
nand UO_137 (O_137,N_2987,N_2978);
and UO_138 (O_138,N_2985,N_2990);
xor UO_139 (O_139,N_2992,N_2988);
and UO_140 (O_140,N_2967,N_2927);
xor UO_141 (O_141,N_2959,N_2976);
nor UO_142 (O_142,N_2942,N_2987);
nand UO_143 (O_143,N_2932,N_2949);
xnor UO_144 (O_144,N_2954,N_2985);
xor UO_145 (O_145,N_2933,N_2981);
nand UO_146 (O_146,N_2952,N_2954);
and UO_147 (O_147,N_2929,N_2994);
or UO_148 (O_148,N_2941,N_2948);
nor UO_149 (O_149,N_2975,N_2977);
or UO_150 (O_150,N_2936,N_2937);
nor UO_151 (O_151,N_2940,N_2947);
xor UO_152 (O_152,N_2955,N_2964);
or UO_153 (O_153,N_2956,N_2955);
nand UO_154 (O_154,N_2959,N_2932);
nor UO_155 (O_155,N_2978,N_2958);
or UO_156 (O_156,N_2954,N_2963);
nand UO_157 (O_157,N_2937,N_2966);
nor UO_158 (O_158,N_2931,N_2939);
nor UO_159 (O_159,N_2966,N_2929);
and UO_160 (O_160,N_2935,N_2927);
nor UO_161 (O_161,N_2981,N_2935);
nor UO_162 (O_162,N_2950,N_2996);
xor UO_163 (O_163,N_2968,N_2993);
or UO_164 (O_164,N_2935,N_2991);
nand UO_165 (O_165,N_2969,N_2972);
or UO_166 (O_166,N_2996,N_2977);
and UO_167 (O_167,N_2973,N_2931);
nand UO_168 (O_168,N_2967,N_2964);
nor UO_169 (O_169,N_2996,N_2931);
or UO_170 (O_170,N_2957,N_2981);
or UO_171 (O_171,N_2973,N_2925);
xnor UO_172 (O_172,N_2980,N_2943);
xor UO_173 (O_173,N_2981,N_2997);
xnor UO_174 (O_174,N_2976,N_2937);
nor UO_175 (O_175,N_2943,N_2963);
nand UO_176 (O_176,N_2932,N_2968);
or UO_177 (O_177,N_2934,N_2939);
and UO_178 (O_178,N_2967,N_2926);
and UO_179 (O_179,N_2987,N_2965);
and UO_180 (O_180,N_2986,N_2947);
and UO_181 (O_181,N_2974,N_2970);
and UO_182 (O_182,N_2994,N_2978);
xor UO_183 (O_183,N_2983,N_2926);
and UO_184 (O_184,N_2964,N_2995);
and UO_185 (O_185,N_2961,N_2970);
or UO_186 (O_186,N_2996,N_2980);
nor UO_187 (O_187,N_2965,N_2925);
nor UO_188 (O_188,N_2935,N_2979);
or UO_189 (O_189,N_2958,N_2942);
nand UO_190 (O_190,N_2969,N_2985);
xnor UO_191 (O_191,N_2944,N_2979);
or UO_192 (O_192,N_2989,N_2956);
and UO_193 (O_193,N_2937,N_2983);
or UO_194 (O_194,N_2961,N_2938);
nor UO_195 (O_195,N_2995,N_2945);
xnor UO_196 (O_196,N_2978,N_2950);
nor UO_197 (O_197,N_2951,N_2949);
xnor UO_198 (O_198,N_2947,N_2949);
or UO_199 (O_199,N_2930,N_2965);
and UO_200 (O_200,N_2942,N_2983);
nor UO_201 (O_201,N_2955,N_2954);
nand UO_202 (O_202,N_2955,N_2961);
nand UO_203 (O_203,N_2968,N_2965);
nand UO_204 (O_204,N_2961,N_2944);
nand UO_205 (O_205,N_2965,N_2960);
or UO_206 (O_206,N_2987,N_2959);
xor UO_207 (O_207,N_2993,N_2958);
and UO_208 (O_208,N_2960,N_2999);
nor UO_209 (O_209,N_2975,N_2966);
or UO_210 (O_210,N_2991,N_2931);
and UO_211 (O_211,N_2969,N_2944);
or UO_212 (O_212,N_2958,N_2936);
nor UO_213 (O_213,N_2947,N_2958);
nor UO_214 (O_214,N_2945,N_2942);
and UO_215 (O_215,N_2947,N_2938);
and UO_216 (O_216,N_2945,N_2975);
or UO_217 (O_217,N_2967,N_2987);
nand UO_218 (O_218,N_2956,N_2998);
nand UO_219 (O_219,N_2973,N_2975);
nand UO_220 (O_220,N_2946,N_2995);
and UO_221 (O_221,N_2992,N_2953);
or UO_222 (O_222,N_2928,N_2934);
and UO_223 (O_223,N_2946,N_2986);
nor UO_224 (O_224,N_2966,N_2994);
nor UO_225 (O_225,N_2981,N_2971);
and UO_226 (O_226,N_2927,N_2973);
nand UO_227 (O_227,N_2936,N_2934);
and UO_228 (O_228,N_2962,N_2991);
and UO_229 (O_229,N_2942,N_2935);
nand UO_230 (O_230,N_2974,N_2946);
and UO_231 (O_231,N_2986,N_2985);
nand UO_232 (O_232,N_2937,N_2975);
nor UO_233 (O_233,N_2969,N_2936);
and UO_234 (O_234,N_2961,N_2983);
and UO_235 (O_235,N_2991,N_2974);
nor UO_236 (O_236,N_2999,N_2925);
nor UO_237 (O_237,N_2993,N_2949);
nor UO_238 (O_238,N_2964,N_2966);
nand UO_239 (O_239,N_2983,N_2995);
and UO_240 (O_240,N_2960,N_2926);
and UO_241 (O_241,N_2975,N_2965);
or UO_242 (O_242,N_2958,N_2998);
xor UO_243 (O_243,N_2970,N_2962);
nand UO_244 (O_244,N_2933,N_2993);
xor UO_245 (O_245,N_2949,N_2953);
and UO_246 (O_246,N_2995,N_2969);
or UO_247 (O_247,N_2937,N_2979);
or UO_248 (O_248,N_2979,N_2957);
or UO_249 (O_249,N_2989,N_2977);
and UO_250 (O_250,N_2940,N_2928);
or UO_251 (O_251,N_2931,N_2948);
and UO_252 (O_252,N_2970,N_2972);
nor UO_253 (O_253,N_2957,N_2995);
or UO_254 (O_254,N_2974,N_2996);
xnor UO_255 (O_255,N_2941,N_2983);
or UO_256 (O_256,N_2946,N_2941);
or UO_257 (O_257,N_2926,N_2973);
and UO_258 (O_258,N_2985,N_2964);
xor UO_259 (O_259,N_2998,N_2948);
or UO_260 (O_260,N_2981,N_2967);
xor UO_261 (O_261,N_2994,N_2984);
nor UO_262 (O_262,N_2954,N_2987);
nand UO_263 (O_263,N_2974,N_2989);
and UO_264 (O_264,N_2994,N_2943);
nor UO_265 (O_265,N_2988,N_2937);
and UO_266 (O_266,N_2970,N_2994);
and UO_267 (O_267,N_2926,N_2989);
nand UO_268 (O_268,N_2948,N_2959);
nor UO_269 (O_269,N_2996,N_2962);
or UO_270 (O_270,N_2999,N_2957);
xnor UO_271 (O_271,N_2941,N_2944);
xnor UO_272 (O_272,N_2926,N_2980);
or UO_273 (O_273,N_2964,N_2974);
and UO_274 (O_274,N_2940,N_2981);
nor UO_275 (O_275,N_2977,N_2927);
or UO_276 (O_276,N_2937,N_2989);
or UO_277 (O_277,N_2954,N_2951);
and UO_278 (O_278,N_2960,N_2945);
and UO_279 (O_279,N_2928,N_2980);
or UO_280 (O_280,N_2933,N_2934);
or UO_281 (O_281,N_2951,N_2927);
nand UO_282 (O_282,N_2979,N_2973);
xnor UO_283 (O_283,N_2940,N_2980);
or UO_284 (O_284,N_2937,N_2934);
nand UO_285 (O_285,N_2944,N_2997);
xor UO_286 (O_286,N_2994,N_2975);
and UO_287 (O_287,N_2959,N_2967);
nand UO_288 (O_288,N_2958,N_2987);
nand UO_289 (O_289,N_2973,N_2992);
nor UO_290 (O_290,N_2953,N_2932);
nor UO_291 (O_291,N_2944,N_2936);
nor UO_292 (O_292,N_2943,N_2967);
nand UO_293 (O_293,N_2962,N_2936);
nand UO_294 (O_294,N_2982,N_2926);
and UO_295 (O_295,N_2977,N_2995);
and UO_296 (O_296,N_2986,N_2936);
xor UO_297 (O_297,N_2943,N_2982);
xor UO_298 (O_298,N_2967,N_2982);
nor UO_299 (O_299,N_2980,N_2932);
or UO_300 (O_300,N_2964,N_2962);
xnor UO_301 (O_301,N_2956,N_2957);
nor UO_302 (O_302,N_2932,N_2936);
nand UO_303 (O_303,N_2934,N_2955);
nor UO_304 (O_304,N_2974,N_2941);
xor UO_305 (O_305,N_2966,N_2996);
or UO_306 (O_306,N_2952,N_2985);
nand UO_307 (O_307,N_2989,N_2940);
xnor UO_308 (O_308,N_2943,N_2953);
xnor UO_309 (O_309,N_2985,N_2981);
or UO_310 (O_310,N_2994,N_2933);
and UO_311 (O_311,N_2972,N_2939);
or UO_312 (O_312,N_2975,N_2948);
nand UO_313 (O_313,N_2940,N_2979);
or UO_314 (O_314,N_2987,N_2996);
and UO_315 (O_315,N_2931,N_2949);
xnor UO_316 (O_316,N_2926,N_2966);
nor UO_317 (O_317,N_2998,N_2934);
xor UO_318 (O_318,N_2979,N_2992);
and UO_319 (O_319,N_2975,N_2978);
or UO_320 (O_320,N_2996,N_2963);
or UO_321 (O_321,N_2965,N_2935);
and UO_322 (O_322,N_2930,N_2933);
nand UO_323 (O_323,N_2995,N_2965);
nand UO_324 (O_324,N_2929,N_2960);
or UO_325 (O_325,N_2976,N_2942);
nor UO_326 (O_326,N_2926,N_2995);
xor UO_327 (O_327,N_2937,N_2965);
xnor UO_328 (O_328,N_2931,N_2954);
and UO_329 (O_329,N_2980,N_2985);
nor UO_330 (O_330,N_2976,N_2956);
xnor UO_331 (O_331,N_2997,N_2935);
or UO_332 (O_332,N_2971,N_2933);
or UO_333 (O_333,N_2928,N_2955);
or UO_334 (O_334,N_2951,N_2940);
xor UO_335 (O_335,N_2954,N_2976);
and UO_336 (O_336,N_2951,N_2935);
or UO_337 (O_337,N_2933,N_2945);
xor UO_338 (O_338,N_2984,N_2947);
nor UO_339 (O_339,N_2943,N_2926);
nor UO_340 (O_340,N_2993,N_2988);
or UO_341 (O_341,N_2976,N_2961);
nor UO_342 (O_342,N_2993,N_2967);
nand UO_343 (O_343,N_2964,N_2951);
xor UO_344 (O_344,N_2969,N_2930);
xor UO_345 (O_345,N_2979,N_2959);
nor UO_346 (O_346,N_2936,N_2938);
xnor UO_347 (O_347,N_2962,N_2955);
xor UO_348 (O_348,N_2993,N_2951);
and UO_349 (O_349,N_2977,N_2958);
and UO_350 (O_350,N_2977,N_2979);
nand UO_351 (O_351,N_2987,N_2936);
and UO_352 (O_352,N_2936,N_2953);
nand UO_353 (O_353,N_2935,N_2930);
nor UO_354 (O_354,N_2951,N_2955);
nand UO_355 (O_355,N_2962,N_2984);
nor UO_356 (O_356,N_2997,N_2940);
nand UO_357 (O_357,N_2930,N_2942);
nor UO_358 (O_358,N_2985,N_2947);
xnor UO_359 (O_359,N_2964,N_2988);
and UO_360 (O_360,N_2933,N_2986);
xor UO_361 (O_361,N_2941,N_2999);
nand UO_362 (O_362,N_2954,N_2947);
nor UO_363 (O_363,N_2932,N_2957);
nand UO_364 (O_364,N_2951,N_2968);
or UO_365 (O_365,N_2979,N_2958);
xnor UO_366 (O_366,N_2945,N_2934);
xnor UO_367 (O_367,N_2983,N_2956);
and UO_368 (O_368,N_2998,N_2954);
xnor UO_369 (O_369,N_2957,N_2997);
xnor UO_370 (O_370,N_2925,N_2985);
xor UO_371 (O_371,N_2991,N_2950);
nor UO_372 (O_372,N_2927,N_2995);
xor UO_373 (O_373,N_2956,N_2937);
and UO_374 (O_374,N_2963,N_2984);
nand UO_375 (O_375,N_2999,N_2965);
nor UO_376 (O_376,N_2982,N_2965);
nor UO_377 (O_377,N_2934,N_2974);
nor UO_378 (O_378,N_2952,N_2982);
xor UO_379 (O_379,N_2954,N_2928);
nand UO_380 (O_380,N_2962,N_2949);
nor UO_381 (O_381,N_2962,N_2979);
xor UO_382 (O_382,N_2928,N_2981);
or UO_383 (O_383,N_2950,N_2943);
xor UO_384 (O_384,N_2938,N_2940);
xor UO_385 (O_385,N_2973,N_2951);
xnor UO_386 (O_386,N_2999,N_2990);
and UO_387 (O_387,N_2963,N_2992);
and UO_388 (O_388,N_2958,N_2940);
and UO_389 (O_389,N_2926,N_2968);
and UO_390 (O_390,N_2995,N_2966);
nor UO_391 (O_391,N_2955,N_2959);
nand UO_392 (O_392,N_2929,N_2958);
xor UO_393 (O_393,N_2961,N_2925);
and UO_394 (O_394,N_2983,N_2959);
xor UO_395 (O_395,N_2932,N_2991);
and UO_396 (O_396,N_2985,N_2960);
nor UO_397 (O_397,N_2967,N_2945);
xnor UO_398 (O_398,N_2943,N_2944);
xor UO_399 (O_399,N_2972,N_2961);
and UO_400 (O_400,N_2994,N_2938);
nor UO_401 (O_401,N_2927,N_2947);
nand UO_402 (O_402,N_2977,N_2992);
or UO_403 (O_403,N_2970,N_2996);
xor UO_404 (O_404,N_2999,N_2963);
xor UO_405 (O_405,N_2955,N_2960);
and UO_406 (O_406,N_2975,N_2989);
and UO_407 (O_407,N_2982,N_2946);
xor UO_408 (O_408,N_2945,N_2980);
nand UO_409 (O_409,N_2964,N_2933);
xor UO_410 (O_410,N_2950,N_2989);
nand UO_411 (O_411,N_2996,N_2958);
and UO_412 (O_412,N_2944,N_2929);
and UO_413 (O_413,N_2942,N_2948);
nor UO_414 (O_414,N_2968,N_2959);
nand UO_415 (O_415,N_2949,N_2970);
and UO_416 (O_416,N_2964,N_2939);
or UO_417 (O_417,N_2974,N_2987);
nand UO_418 (O_418,N_2932,N_2986);
or UO_419 (O_419,N_2987,N_2989);
nor UO_420 (O_420,N_2991,N_2949);
and UO_421 (O_421,N_2925,N_2974);
nor UO_422 (O_422,N_2936,N_2973);
nor UO_423 (O_423,N_2938,N_2937);
and UO_424 (O_424,N_2946,N_2936);
xnor UO_425 (O_425,N_2992,N_2981);
or UO_426 (O_426,N_2973,N_2960);
nor UO_427 (O_427,N_2973,N_2988);
or UO_428 (O_428,N_2997,N_2978);
nor UO_429 (O_429,N_2978,N_2948);
nor UO_430 (O_430,N_2933,N_2996);
nor UO_431 (O_431,N_2938,N_2943);
and UO_432 (O_432,N_2972,N_2938);
or UO_433 (O_433,N_2993,N_2972);
and UO_434 (O_434,N_2990,N_2957);
nand UO_435 (O_435,N_2956,N_2952);
and UO_436 (O_436,N_2954,N_2959);
xor UO_437 (O_437,N_2960,N_2935);
xnor UO_438 (O_438,N_2993,N_2938);
nand UO_439 (O_439,N_2926,N_2979);
nand UO_440 (O_440,N_2971,N_2937);
or UO_441 (O_441,N_2925,N_2949);
nor UO_442 (O_442,N_2965,N_2949);
or UO_443 (O_443,N_2959,N_2998);
and UO_444 (O_444,N_2938,N_2982);
nand UO_445 (O_445,N_2976,N_2930);
nor UO_446 (O_446,N_2969,N_2937);
nand UO_447 (O_447,N_2970,N_2956);
or UO_448 (O_448,N_2960,N_2983);
or UO_449 (O_449,N_2990,N_2935);
or UO_450 (O_450,N_2969,N_2965);
nor UO_451 (O_451,N_2976,N_2993);
or UO_452 (O_452,N_2982,N_2972);
nor UO_453 (O_453,N_2984,N_2934);
and UO_454 (O_454,N_2980,N_2989);
nand UO_455 (O_455,N_2965,N_2953);
and UO_456 (O_456,N_2995,N_2988);
xor UO_457 (O_457,N_2934,N_2970);
xnor UO_458 (O_458,N_2944,N_2967);
xor UO_459 (O_459,N_2990,N_2998);
or UO_460 (O_460,N_2985,N_2962);
or UO_461 (O_461,N_2998,N_2999);
nand UO_462 (O_462,N_2948,N_2970);
xor UO_463 (O_463,N_2955,N_2977);
nand UO_464 (O_464,N_2926,N_2950);
or UO_465 (O_465,N_2989,N_2948);
or UO_466 (O_466,N_2978,N_2941);
and UO_467 (O_467,N_2995,N_2925);
nor UO_468 (O_468,N_2994,N_2926);
or UO_469 (O_469,N_2931,N_2983);
or UO_470 (O_470,N_2992,N_2999);
or UO_471 (O_471,N_2953,N_2951);
nand UO_472 (O_472,N_2989,N_2938);
or UO_473 (O_473,N_2961,N_2954);
or UO_474 (O_474,N_2999,N_2929);
nand UO_475 (O_475,N_2996,N_2940);
nand UO_476 (O_476,N_2927,N_2992);
nand UO_477 (O_477,N_2942,N_2925);
or UO_478 (O_478,N_2934,N_2999);
nand UO_479 (O_479,N_2939,N_2936);
or UO_480 (O_480,N_2992,N_2965);
xnor UO_481 (O_481,N_2991,N_2996);
and UO_482 (O_482,N_2955,N_2972);
nand UO_483 (O_483,N_2945,N_2935);
and UO_484 (O_484,N_2942,N_2932);
xnor UO_485 (O_485,N_2966,N_2932);
and UO_486 (O_486,N_2961,N_2971);
xor UO_487 (O_487,N_2945,N_2983);
nand UO_488 (O_488,N_2989,N_2979);
and UO_489 (O_489,N_2950,N_2951);
and UO_490 (O_490,N_2992,N_2957);
or UO_491 (O_491,N_2928,N_2931);
and UO_492 (O_492,N_2990,N_2983);
xnor UO_493 (O_493,N_2929,N_2989);
xor UO_494 (O_494,N_2996,N_2937);
nand UO_495 (O_495,N_2933,N_2970);
nand UO_496 (O_496,N_2945,N_2981);
xnor UO_497 (O_497,N_2969,N_2959);
and UO_498 (O_498,N_2974,N_2965);
nor UO_499 (O_499,N_2952,N_2935);
endmodule