module basic_750_5000_1000_2_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2502,N_2503,N_2504,N_2506,N_2508,N_2509,N_2510,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2530,N_2532,N_2534,N_2535,N_2537,N_2538,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2553,N_2554,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2566,N_2567,N_2568,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2592,N_2593,N_2594,N_2595,N_2596,N_2598,N_2599,N_2600,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2634,N_2635,N_2636,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2661,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2702,N_2703,N_2704,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2718,N_2719,N_2720,N_2721,N_2722,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2746,N_2747,N_2748,N_2749,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2768,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2783,N_2784,N_2785,N_2787,N_2790,N_2791,N_2792,N_2793,N_2794,N_2797,N_2798,N_2799,N_2801,N_2802,N_2804,N_2805,N_2806,N_2807,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2843,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2877,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2904,N_2905,N_2906,N_2907,N_2908,N_2910,N_2911,N_2912,N_2913,N_2914,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2925,N_2926,N_2928,N_2929,N_2930,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2947,N_2950,N_2951,N_2952,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2967,N_2968,N_2970,N_2971,N_2972,N_2973,N_2975,N_2976,N_2977,N_2979,N_2982,N_2984,N_2985,N_2986,N_2987,N_2988,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2997,N_2998,N_2999,N_3000,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3011,N_3012,N_3014,N_3015,N_3017,N_3018,N_3019,N_3022,N_3026,N_3028,N_3029,N_3032,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3047,N_3048,N_3051,N_3052,N_3053,N_3054,N_3056,N_3057,N_3058,N_3059,N_3061,N_3062,N_3064,N_3066,N_3067,N_3069,N_3071,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3083,N_3084,N_3085,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3102,N_3103,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3112,N_3113,N_3114,N_3115,N_3117,N_3118,N_3119,N_3120,N_3121,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3161,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3174,N_3175,N_3176,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3190,N_3191,N_3192,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3201,N_3203,N_3204,N_3205,N_3206,N_3208,N_3209,N_3210,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3223,N_3224,N_3225,N_3226,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3236,N_3237,N_3238,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3249,N_3250,N_3251,N_3252,N_3253,N_3255,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3264,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3296,N_3297,N_3298,N_3299,N_3300,N_3302,N_3304,N_3305,N_3307,N_3308,N_3309,N_3310,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3321,N_3323,N_3324,N_3325,N_3326,N_3328,N_3329,N_3330,N_3332,N_3334,N_3335,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3347,N_3348,N_3349,N_3350,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3361,N_3362,N_3363,N_3364,N_3366,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3380,N_3381,N_3383,N_3385,N_3387,N_3388,N_3389,N_3393,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3421,N_3422,N_3425,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3441,N_3442,N_3443,N_3444,N_3447,N_3449,N_3450,N_3451,N_3452,N_3454,N_3455,N_3456,N_3457,N_3458,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3469,N_3470,N_3472,N_3473,N_3474,N_3476,N_3478,N_3479,N_3480,N_3481,N_3483,N_3484,N_3486,N_3487,N_3488,N_3489,N_3490,N_3492,N_3495,N_3496,N_3497,N_3498,N_3500,N_3504,N_3505,N_3506,N_3507,N_3509,N_3510,N_3511,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3533,N_3534,N_3535,N_3536,N_3537,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3550,N_3551,N_3552,N_3553,N_3554,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3572,N_3573,N_3574,N_3575,N_3576,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3596,N_3597,N_3599,N_3600,N_3602,N_3603,N_3604,N_3605,N_3607,N_3608,N_3609,N_3610,N_3611,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3625,N_3626,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3661,N_3662,N_3663,N_3664,N_3666,N_3667,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3679,N_3681,N_3682,N_3683,N_3684,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3693,N_3694,N_3696,N_3697,N_3699,N_3700,N_3701,N_3702,N_3704,N_3705,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3727,N_3728,N_3729,N_3730,N_3731,N_3733,N_3735,N_3736,N_3737,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3749,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3759,N_3760,N_3761,N_3762,N_3764,N_3765,N_3767,N_3768,N_3769,N_3771,N_3772,N_3775,N_3776,N_3777,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3798,N_3799,N_3800,N_3801,N_3803,N_3805,N_3806,N_3807,N_3809,N_3811,N_3812,N_3813,N_3814,N_3817,N_3818,N_3820,N_3822,N_3823,N_3824,N_3825,N_3826,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3850,N_3851,N_3853,N_3854,N_3855,N_3856,N_3858,N_3860,N_3861,N_3863,N_3864,N_3865,N_3868,N_3870,N_3873,N_3874,N_3876,N_3877,N_3878,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3898,N_3899,N_3900,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3917,N_3918,N_3919,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3930,N_3931,N_3932,N_3933,N_3935,N_3937,N_3938,N_3939,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3957,N_3958,N_3959,N_3961,N_3962,N_3964,N_3965,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3974,N_3975,N_3976,N_3977,N_3978,N_3980,N_3981,N_3983,N_3985,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3998,N_3999,N_4000,N_4001,N_4005,N_4006,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4017,N_4018,N_4019,N_4020,N_4021,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4056,N_4057,N_4058,N_4059,N_4062,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4083,N_4085,N_4089,N_4091,N_4094,N_4095,N_4096,N_4097,N_4099,N_4101,N_4102,N_4104,N_4106,N_4107,N_4108,N_4111,N_4112,N_4113,N_4115,N_4116,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4128,N_4130,N_4131,N_4132,N_4133,N_4135,N_4136,N_4140,N_4142,N_4143,N_4144,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4216,N_4218,N_4219,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4236,N_4237,N_4240,N_4241,N_4242,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4297,N_4298,N_4300,N_4301,N_4302,N_4303,N_4304,N_4308,N_4309,N_4310,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4319,N_4321,N_4322,N_4325,N_4326,N_4327,N_4328,N_4329,N_4331,N_4333,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4355,N_4356,N_4357,N_4358,N_4359,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4369,N_4370,N_4371,N_4372,N_4373,N_4375,N_4376,N_4377,N_4378,N_4380,N_4381,N_4382,N_4383,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4401,N_4402,N_4404,N_4407,N_4408,N_4410,N_4412,N_4414,N_4416,N_4417,N_4418,N_4420,N_4421,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4430,N_4431,N_4434,N_4435,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4444,N_4445,N_4446,N_4447,N_4448,N_4451,N_4452,N_4453,N_4454,N_4455,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4473,N_4474,N_4476,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4505,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4519,N_4520,N_4521,N_4524,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4541,N_4542,N_4543,N_4545,N_4546,N_4547,N_4548,N_4549,N_4551,N_4552,N_4553,N_4555,N_4556,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4589,N_4590,N_4591,N_4592,N_4593,N_4595,N_4597,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4637,N_4638,N_4640,N_4641,N_4644,N_4645,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4681,N_4682,N_4683,N_4684,N_4686,N_4687,N_4690,N_4691,N_4692,N_4693,N_4695,N_4696,N_4697,N_4698,N_4699,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4714,N_4716,N_4717,N_4719,N_4720,N_4721,N_4722,N_4723,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4754,N_4755,N_4756,N_4759,N_4760,N_4762,N_4763,N_4764,N_4766,N_4767,N_4768,N_4770,N_4771,N_4774,N_4775,N_4776,N_4777,N_4778,N_4780,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4789,N_4790,N_4791,N_4792,N_4793,N_4795,N_4796,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4806,N_4807,N_4808,N_4810,N_4811,N_4813,N_4814,N_4816,N_4817,N_4818,N_4820,N_4823,N_4824,N_4826,N_4827,N_4828,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4841,N_4843,N_4844,N_4845,N_4847,N_4848,N_4849,N_4850,N_4851,N_4853,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4867,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4890,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4902,N_4903,N_4905,N_4909,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4934,N_4935,N_4936,N_4937,N_4938,N_4940,N_4941,N_4942,N_4943,N_4945,N_4946,N_4947,N_4948,N_4949,N_4952,N_4954,N_4956,N_4957,N_4958,N_4963,N_4964,N_4966,N_4967,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4978,N_4979,N_4980,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_255,In_299);
nand U1 (N_1,In_319,In_252);
nor U2 (N_2,In_73,In_179);
and U3 (N_3,In_532,In_12);
nor U4 (N_4,In_157,In_547);
xor U5 (N_5,In_449,In_355);
and U6 (N_6,In_172,In_257);
nand U7 (N_7,In_431,In_376);
xor U8 (N_8,In_639,In_698);
nand U9 (N_9,In_254,In_279);
or U10 (N_10,In_505,In_262);
xnor U11 (N_11,In_478,In_250);
and U12 (N_12,In_15,In_368);
and U13 (N_13,In_336,In_499);
nor U14 (N_14,In_328,In_79);
or U15 (N_15,In_161,In_354);
xor U16 (N_16,In_261,In_677);
or U17 (N_17,In_652,In_116);
or U18 (N_18,In_451,In_281);
or U19 (N_19,In_616,In_214);
nand U20 (N_20,In_468,In_231);
xnor U21 (N_21,In_174,In_62);
xnor U22 (N_22,In_373,In_703);
nand U23 (N_23,In_317,In_592);
xnor U24 (N_24,In_92,In_447);
nand U25 (N_25,In_171,In_503);
nor U26 (N_26,In_50,In_63);
nand U27 (N_27,In_168,In_207);
and U28 (N_28,In_393,In_372);
or U29 (N_29,In_697,In_264);
nand U30 (N_30,In_40,In_100);
xor U31 (N_31,In_342,In_506);
xor U32 (N_32,In_126,In_102);
or U33 (N_33,In_464,In_632);
or U34 (N_34,In_270,In_98);
nand U35 (N_35,In_541,In_184);
xnor U36 (N_36,In_334,In_351);
or U37 (N_37,In_203,In_398);
and U38 (N_38,In_635,In_143);
and U39 (N_39,In_327,In_346);
or U40 (N_40,In_21,In_687);
xnor U41 (N_41,In_491,In_2);
and U42 (N_42,In_484,In_735);
and U43 (N_43,In_104,In_52);
and U44 (N_44,In_717,In_719);
nor U45 (N_45,In_511,In_278);
xnor U46 (N_46,In_650,In_529);
and U47 (N_47,In_572,In_238);
or U48 (N_48,In_326,In_227);
nor U49 (N_49,In_366,In_187);
nand U50 (N_50,In_221,In_256);
and U51 (N_51,In_260,In_438);
nand U52 (N_52,In_331,In_378);
nor U53 (N_53,In_708,In_25);
or U54 (N_54,In_646,In_681);
nor U55 (N_55,In_230,In_425);
nand U56 (N_56,In_688,In_672);
xnor U57 (N_57,In_640,In_686);
or U58 (N_58,In_661,In_212);
nor U59 (N_59,In_525,In_399);
nor U60 (N_60,In_141,In_200);
xor U61 (N_61,In_655,In_169);
or U62 (N_62,In_713,In_285);
nor U63 (N_63,In_300,In_27);
nand U64 (N_64,In_690,In_313);
nand U65 (N_65,In_612,In_87);
and U66 (N_66,In_287,In_587);
nand U67 (N_67,In_24,In_213);
xor U68 (N_68,In_195,In_452);
or U69 (N_69,In_266,In_105);
or U70 (N_70,In_177,In_35);
xnor U71 (N_71,In_404,In_392);
nand U72 (N_72,In_429,In_275);
xor U73 (N_73,In_704,In_527);
or U74 (N_74,In_208,In_526);
or U75 (N_75,In_34,In_144);
and U76 (N_76,In_185,In_94);
nor U77 (N_77,In_479,In_340);
and U78 (N_78,In_454,In_14);
nand U79 (N_79,In_442,In_173);
or U80 (N_80,In_736,In_394);
or U81 (N_81,In_155,In_246);
xnor U82 (N_82,In_515,In_546);
nor U83 (N_83,In_306,In_647);
nand U84 (N_84,In_241,In_406);
xnor U85 (N_85,In_217,In_630);
and U86 (N_86,In_65,In_348);
xor U87 (N_87,In_95,In_47);
and U88 (N_88,In_699,In_358);
nor U89 (N_89,In_339,In_320);
and U90 (N_90,In_443,In_568);
xor U91 (N_91,In_705,In_83);
and U92 (N_92,In_508,In_20);
xnor U93 (N_93,In_183,In_710);
nor U94 (N_94,In_298,In_408);
or U95 (N_95,In_69,In_232);
or U96 (N_96,In_223,In_82);
xor U97 (N_97,In_78,In_510);
nor U98 (N_98,In_46,In_163);
xor U99 (N_99,In_165,In_108);
xnor U100 (N_100,In_124,In_607);
or U101 (N_101,In_471,In_553);
or U102 (N_102,In_741,In_676);
nor U103 (N_103,In_42,In_347);
nand U104 (N_104,In_90,In_110);
nor U105 (N_105,In_463,In_193);
xnor U106 (N_106,In_170,In_590);
or U107 (N_107,In_536,In_577);
nand U108 (N_108,In_582,In_718);
or U109 (N_109,In_53,In_413);
xnor U110 (N_110,In_588,In_18);
or U111 (N_111,In_96,In_473);
nor U112 (N_112,In_625,In_29);
nor U113 (N_113,In_337,In_322);
xnor U114 (N_114,In_109,In_222);
nand U115 (N_115,In_733,In_528);
xnor U116 (N_116,In_595,In_216);
or U117 (N_117,In_742,In_335);
nor U118 (N_118,In_234,In_701);
xnor U119 (N_119,In_269,In_516);
and U120 (N_120,In_706,In_305);
nor U121 (N_121,In_501,In_122);
or U122 (N_122,In_312,In_498);
or U123 (N_123,In_416,In_16);
and U124 (N_124,In_395,In_537);
and U125 (N_125,In_1,In_660);
xor U126 (N_126,In_74,In_307);
nor U127 (N_127,In_680,In_389);
or U128 (N_128,In_80,In_417);
nor U129 (N_129,In_68,In_75);
xor U130 (N_130,In_602,In_103);
nor U131 (N_131,In_59,In_477);
or U132 (N_132,In_411,In_301);
xnor U133 (N_133,In_39,In_286);
xor U134 (N_134,In_675,In_695);
or U135 (N_135,In_436,In_684);
or U136 (N_136,In_485,In_437);
or U137 (N_137,In_175,In_722);
nor U138 (N_138,In_600,In_581);
nor U139 (N_139,In_380,In_707);
nand U140 (N_140,In_666,In_518);
or U141 (N_141,In_629,In_237);
or U142 (N_142,In_749,In_455);
xor U143 (N_143,In_397,In_245);
xor U144 (N_144,In_199,In_127);
xor U145 (N_145,In_106,In_148);
nor U146 (N_146,In_93,In_130);
or U147 (N_147,In_194,In_494);
and U148 (N_148,In_283,In_166);
nand U149 (N_149,In_633,In_272);
nand U150 (N_150,In_186,In_382);
nor U151 (N_151,In_44,In_435);
or U152 (N_152,In_86,In_303);
nand U153 (N_153,In_598,In_349);
nor U154 (N_154,In_641,In_315);
nand U155 (N_155,In_152,In_353);
nor U156 (N_156,In_357,In_49);
xor U157 (N_157,In_739,In_330);
nor U158 (N_158,In_290,In_81);
nand U159 (N_159,In_259,In_524);
nand U160 (N_160,In_206,In_424);
or U161 (N_161,In_663,In_111);
nor U162 (N_162,In_651,In_534);
or U163 (N_163,In_211,In_115);
nor U164 (N_164,In_388,In_570);
and U165 (N_165,In_282,In_198);
nor U166 (N_166,In_428,In_530);
nand U167 (N_167,In_539,In_11);
nand U168 (N_168,In_609,In_365);
and U169 (N_169,In_673,In_377);
nand U170 (N_170,In_421,In_731);
nor U171 (N_171,In_268,In_402);
nand U172 (N_172,In_386,In_407);
or U173 (N_173,In_531,In_734);
nand U174 (N_174,In_26,In_369);
nor U175 (N_175,In_434,In_744);
xor U176 (N_176,In_176,In_670);
nor U177 (N_177,In_644,In_72);
nor U178 (N_178,In_637,In_575);
or U179 (N_179,In_132,In_167);
and U180 (N_180,In_419,In_329);
or U181 (N_181,In_310,In_64);
nand U182 (N_182,In_461,In_0);
nor U183 (N_183,In_201,In_113);
xnor U184 (N_184,In_476,In_679);
and U185 (N_185,In_32,In_37);
or U186 (N_186,In_469,In_38);
nor U187 (N_187,In_239,In_542);
nand U188 (N_188,In_138,In_274);
nand U189 (N_189,In_444,In_22);
xnor U190 (N_190,In_601,In_296);
nand U191 (N_191,In_263,In_89);
and U192 (N_192,In_638,In_385);
or U193 (N_193,In_658,In_605);
or U194 (N_194,In_117,In_209);
nor U195 (N_195,In_521,In_215);
nand U196 (N_196,In_360,In_613);
xor U197 (N_197,In_375,In_668);
nand U198 (N_198,In_645,In_604);
xor U199 (N_199,In_314,In_573);
and U200 (N_200,In_456,In_128);
nor U201 (N_201,In_308,In_709);
or U202 (N_202,In_235,In_316);
nor U203 (N_203,In_147,In_101);
nor U204 (N_204,In_164,In_17);
or U205 (N_205,In_715,In_747);
or U206 (N_206,In_657,In_420);
nand U207 (N_207,In_487,In_669);
or U208 (N_208,In_664,In_77);
or U209 (N_209,In_384,In_76);
or U210 (N_210,In_691,In_125);
and U211 (N_211,In_273,In_13);
nor U212 (N_212,In_696,In_370);
xor U213 (N_213,In_31,In_61);
or U214 (N_214,In_129,In_154);
nand U215 (N_215,In_514,In_359);
or U216 (N_216,In_569,In_114);
and U217 (N_217,In_57,In_190);
nand U218 (N_218,In_615,In_544);
and U219 (N_219,In_674,In_390);
nand U220 (N_220,In_692,In_276);
or U221 (N_221,In_379,In_121);
nor U222 (N_222,In_492,In_160);
nand U223 (N_223,In_627,In_567);
nor U224 (N_224,In_247,In_689);
xor U225 (N_225,In_162,In_220);
or U226 (N_226,In_445,In_594);
nor U227 (N_227,In_711,In_383);
or U228 (N_228,In_659,In_396);
nand U229 (N_229,In_146,In_586);
xor U230 (N_230,In_362,In_648);
nor U231 (N_231,In_562,In_432);
and U232 (N_232,In_563,In_345);
and U233 (N_233,In_422,In_457);
and U234 (N_234,In_520,In_311);
or U235 (N_235,In_367,In_597);
nor U236 (N_236,In_665,In_728);
and U237 (N_237,In_448,In_504);
and U238 (N_238,In_682,In_671);
or U239 (N_239,In_374,In_19);
xor U240 (N_240,In_325,In_656);
nor U241 (N_241,In_636,In_410);
xor U242 (N_242,In_294,In_423);
nand U243 (N_243,In_611,In_140);
xor U244 (N_244,In_551,In_361);
nand U245 (N_245,In_191,In_667);
nor U246 (N_246,In_277,In_589);
xnor U247 (N_247,In_614,In_500);
xnor U248 (N_248,In_540,In_565);
xor U249 (N_249,In_149,In_721);
nand U250 (N_250,In_248,In_210);
nor U251 (N_251,In_723,In_558);
nand U252 (N_252,In_585,In_700);
nor U253 (N_253,In_371,In_48);
or U254 (N_254,In_617,In_694);
or U255 (N_255,In_30,In_550);
xor U256 (N_256,In_579,In_566);
nor U257 (N_257,In_97,In_134);
nor U258 (N_258,In_189,In_137);
xor U259 (N_259,In_318,In_88);
xor U260 (N_260,In_490,In_578);
nor U261 (N_261,In_242,In_466);
nand U262 (N_262,In_10,In_634);
nor U263 (N_263,In_60,In_71);
nand U264 (N_264,In_7,In_352);
or U265 (N_265,In_488,In_297);
nand U266 (N_266,In_120,In_8);
and U267 (N_267,In_150,In_497);
nand U268 (N_268,In_462,In_626);
or U269 (N_269,In_430,In_561);
nand U270 (N_270,In_649,In_350);
or U271 (N_271,In_653,In_538);
nor U272 (N_272,In_243,In_182);
and U273 (N_273,In_219,In_267);
nor U274 (N_274,In_738,In_743);
nor U275 (N_275,In_284,In_493);
xor U276 (N_276,In_470,In_543);
or U277 (N_277,In_439,In_433);
or U278 (N_278,In_574,In_55);
nor U279 (N_279,In_412,In_599);
nor U280 (N_280,In_486,In_344);
xnor U281 (N_281,In_745,In_584);
nand U282 (N_282,In_643,In_323);
nand U283 (N_283,In_84,In_99);
and U284 (N_284,In_249,In_475);
and U285 (N_285,In_218,In_460);
nor U286 (N_286,In_321,In_85);
or U287 (N_287,In_4,In_554);
or U288 (N_288,In_3,In_123);
and U289 (N_289,In_180,In_603);
or U290 (N_290,In_642,In_156);
nor U291 (N_291,In_291,In_740);
nor U292 (N_292,In_236,In_480);
nor U293 (N_293,In_446,In_414);
xor U294 (N_294,In_387,In_181);
and U295 (N_295,In_729,In_610);
and U296 (N_296,In_324,In_43);
nor U297 (N_297,In_440,In_233);
nand U298 (N_298,In_304,In_560);
nand U299 (N_299,In_712,In_409);
nor U300 (N_300,In_107,In_228);
nor U301 (N_301,In_482,In_522);
nand U302 (N_302,In_622,In_564);
nor U303 (N_303,In_606,In_67);
and U304 (N_304,In_158,In_621);
and U305 (N_305,In_224,In_662);
xnor U306 (N_306,In_118,In_244);
or U307 (N_307,In_474,In_205);
or U308 (N_308,In_293,In_131);
or U309 (N_309,In_748,In_58);
nor U310 (N_310,In_202,In_702);
nand U311 (N_311,In_136,In_557);
nor U312 (N_312,In_683,In_608);
nor U313 (N_313,In_288,In_280);
and U314 (N_314,In_495,In_596);
nand U315 (N_315,In_545,In_555);
or U316 (N_316,In_467,In_618);
nand U317 (N_317,In_289,In_502);
and U318 (N_318,In_41,In_583);
and U319 (N_319,In_401,In_591);
nor U320 (N_320,In_552,In_513);
and U321 (N_321,In_619,In_251);
or U322 (N_322,In_453,In_620);
nor U323 (N_323,In_54,In_341);
xnor U324 (N_324,In_654,In_441);
and U325 (N_325,In_559,In_28);
and U326 (N_326,In_204,In_746);
xor U327 (N_327,In_693,In_727);
nand U328 (N_328,In_523,In_403);
and U329 (N_329,In_391,In_631);
nor U330 (N_330,In_405,In_225);
or U331 (N_331,In_509,In_678);
nor U332 (N_332,In_139,In_623);
nand U333 (N_333,In_253,In_685);
nand U334 (N_334,In_483,In_549);
xnor U335 (N_335,In_178,In_418);
nand U336 (N_336,In_400,In_548);
nand U337 (N_337,In_119,In_512);
and U338 (N_338,In_624,In_427);
nor U339 (N_339,In_295,In_338);
or U340 (N_340,In_472,In_56);
nor U341 (N_341,In_197,In_450);
nor U342 (N_342,In_302,In_240);
xor U343 (N_343,In_23,In_732);
and U344 (N_344,In_45,In_151);
and U345 (N_345,In_133,In_737);
nand U346 (N_346,In_70,In_142);
nand U347 (N_347,In_724,In_265);
and U348 (N_348,In_343,In_33);
or U349 (N_349,In_6,In_714);
or U350 (N_350,In_145,In_309);
nand U351 (N_351,In_153,In_333);
xor U352 (N_352,In_135,In_519);
nor U353 (N_353,In_258,In_271);
and U354 (N_354,In_112,In_364);
and U355 (N_355,In_51,In_229);
and U356 (N_356,In_576,In_363);
and U357 (N_357,In_517,In_580);
nor U358 (N_358,In_628,In_91);
nor U359 (N_359,In_36,In_226);
nor U360 (N_360,In_9,In_459);
xnor U361 (N_361,In_188,In_5);
nor U362 (N_362,In_465,In_571);
nand U363 (N_363,In_720,In_292);
and U364 (N_364,In_725,In_66);
and U365 (N_365,In_192,In_159);
or U366 (N_366,In_533,In_726);
nand U367 (N_367,In_481,In_496);
nand U368 (N_368,In_458,In_730);
xor U369 (N_369,In_426,In_556);
nand U370 (N_370,In_507,In_332);
nand U371 (N_371,In_196,In_415);
nor U372 (N_372,In_356,In_593);
xnor U373 (N_373,In_716,In_489);
nand U374 (N_374,In_381,In_535);
and U375 (N_375,In_733,In_715);
and U376 (N_376,In_715,In_486);
and U377 (N_377,In_230,In_545);
or U378 (N_378,In_559,In_549);
xor U379 (N_379,In_163,In_547);
nor U380 (N_380,In_76,In_29);
or U381 (N_381,In_495,In_164);
xnor U382 (N_382,In_229,In_727);
nand U383 (N_383,In_103,In_593);
or U384 (N_384,In_663,In_91);
nand U385 (N_385,In_23,In_36);
nor U386 (N_386,In_68,In_453);
nor U387 (N_387,In_150,In_675);
and U388 (N_388,In_325,In_725);
or U389 (N_389,In_76,In_207);
and U390 (N_390,In_303,In_197);
and U391 (N_391,In_320,In_672);
nor U392 (N_392,In_503,In_404);
nand U393 (N_393,In_530,In_90);
nor U394 (N_394,In_208,In_44);
xnor U395 (N_395,In_608,In_56);
xnor U396 (N_396,In_660,In_68);
or U397 (N_397,In_13,In_416);
xnor U398 (N_398,In_44,In_441);
and U399 (N_399,In_210,In_4);
and U400 (N_400,In_668,In_35);
nor U401 (N_401,In_735,In_443);
xor U402 (N_402,In_233,In_615);
nor U403 (N_403,In_103,In_611);
nor U404 (N_404,In_198,In_69);
nor U405 (N_405,In_26,In_351);
nor U406 (N_406,In_630,In_385);
nor U407 (N_407,In_405,In_75);
and U408 (N_408,In_78,In_625);
nor U409 (N_409,In_168,In_219);
or U410 (N_410,In_123,In_649);
nand U411 (N_411,In_145,In_124);
nor U412 (N_412,In_316,In_365);
xnor U413 (N_413,In_291,In_121);
nor U414 (N_414,In_369,In_487);
nor U415 (N_415,In_608,In_567);
xor U416 (N_416,In_43,In_672);
xor U417 (N_417,In_104,In_277);
and U418 (N_418,In_262,In_280);
or U419 (N_419,In_644,In_546);
xor U420 (N_420,In_577,In_552);
nand U421 (N_421,In_595,In_122);
xor U422 (N_422,In_738,In_631);
xor U423 (N_423,In_698,In_202);
nand U424 (N_424,In_249,In_383);
nor U425 (N_425,In_248,In_140);
and U426 (N_426,In_626,In_644);
nand U427 (N_427,In_12,In_722);
xor U428 (N_428,In_244,In_645);
nand U429 (N_429,In_473,In_101);
nand U430 (N_430,In_240,In_724);
xnor U431 (N_431,In_480,In_37);
nor U432 (N_432,In_446,In_626);
or U433 (N_433,In_598,In_723);
or U434 (N_434,In_430,In_658);
nand U435 (N_435,In_345,In_349);
or U436 (N_436,In_523,In_673);
nand U437 (N_437,In_648,In_592);
or U438 (N_438,In_509,In_423);
or U439 (N_439,In_166,In_194);
nor U440 (N_440,In_729,In_375);
or U441 (N_441,In_587,In_557);
nor U442 (N_442,In_366,In_499);
nand U443 (N_443,In_184,In_256);
and U444 (N_444,In_113,In_548);
nor U445 (N_445,In_354,In_725);
or U446 (N_446,In_203,In_214);
and U447 (N_447,In_189,In_541);
nor U448 (N_448,In_131,In_357);
and U449 (N_449,In_189,In_37);
nor U450 (N_450,In_467,In_605);
nand U451 (N_451,In_365,In_430);
nor U452 (N_452,In_489,In_448);
xor U453 (N_453,In_69,In_725);
xnor U454 (N_454,In_87,In_245);
and U455 (N_455,In_164,In_694);
nand U456 (N_456,In_128,In_313);
and U457 (N_457,In_606,In_131);
xor U458 (N_458,In_684,In_726);
xor U459 (N_459,In_743,In_679);
xnor U460 (N_460,In_450,In_368);
or U461 (N_461,In_340,In_588);
and U462 (N_462,In_584,In_386);
nand U463 (N_463,In_65,In_591);
nor U464 (N_464,In_729,In_146);
nor U465 (N_465,In_317,In_160);
nand U466 (N_466,In_221,In_192);
and U467 (N_467,In_81,In_555);
xnor U468 (N_468,In_316,In_67);
or U469 (N_469,In_545,In_17);
nor U470 (N_470,In_262,In_650);
xnor U471 (N_471,In_316,In_32);
and U472 (N_472,In_50,In_683);
nand U473 (N_473,In_312,In_7);
xnor U474 (N_474,In_69,In_255);
xnor U475 (N_475,In_99,In_55);
nor U476 (N_476,In_528,In_137);
or U477 (N_477,In_536,In_603);
and U478 (N_478,In_534,In_476);
nor U479 (N_479,In_68,In_733);
nand U480 (N_480,In_603,In_346);
xnor U481 (N_481,In_423,In_395);
or U482 (N_482,In_686,In_167);
nor U483 (N_483,In_610,In_398);
or U484 (N_484,In_665,In_597);
xor U485 (N_485,In_186,In_372);
or U486 (N_486,In_113,In_151);
nor U487 (N_487,In_20,In_314);
and U488 (N_488,In_375,In_517);
nand U489 (N_489,In_416,In_46);
xnor U490 (N_490,In_462,In_103);
xnor U491 (N_491,In_499,In_265);
nor U492 (N_492,In_92,In_14);
xnor U493 (N_493,In_557,In_717);
xor U494 (N_494,In_80,In_503);
or U495 (N_495,In_296,In_548);
xnor U496 (N_496,In_500,In_737);
nand U497 (N_497,In_587,In_210);
nor U498 (N_498,In_467,In_470);
or U499 (N_499,In_9,In_34);
and U500 (N_500,In_558,In_76);
or U501 (N_501,In_445,In_578);
or U502 (N_502,In_740,In_76);
nor U503 (N_503,In_694,In_387);
nand U504 (N_504,In_511,In_383);
and U505 (N_505,In_503,In_610);
and U506 (N_506,In_109,In_664);
nand U507 (N_507,In_211,In_677);
xor U508 (N_508,In_208,In_475);
and U509 (N_509,In_290,In_480);
and U510 (N_510,In_139,In_663);
nand U511 (N_511,In_368,In_183);
nand U512 (N_512,In_688,In_469);
nor U513 (N_513,In_564,In_243);
nand U514 (N_514,In_741,In_683);
nand U515 (N_515,In_279,In_709);
xnor U516 (N_516,In_183,In_448);
nand U517 (N_517,In_94,In_644);
nand U518 (N_518,In_188,In_442);
and U519 (N_519,In_491,In_243);
xnor U520 (N_520,In_564,In_62);
nor U521 (N_521,In_105,In_698);
or U522 (N_522,In_446,In_665);
xnor U523 (N_523,In_140,In_552);
nor U524 (N_524,In_422,In_112);
or U525 (N_525,In_742,In_508);
and U526 (N_526,In_476,In_309);
nor U527 (N_527,In_518,In_235);
nand U528 (N_528,In_291,In_69);
nor U529 (N_529,In_541,In_249);
nor U530 (N_530,In_535,In_132);
nand U531 (N_531,In_215,In_301);
nor U532 (N_532,In_272,In_210);
nand U533 (N_533,In_593,In_491);
or U534 (N_534,In_588,In_551);
or U535 (N_535,In_380,In_326);
and U536 (N_536,In_559,In_564);
nor U537 (N_537,In_379,In_330);
and U538 (N_538,In_469,In_7);
nand U539 (N_539,In_6,In_244);
nand U540 (N_540,In_221,In_642);
and U541 (N_541,In_632,In_327);
xnor U542 (N_542,In_381,In_148);
and U543 (N_543,In_360,In_280);
nand U544 (N_544,In_168,In_56);
and U545 (N_545,In_597,In_648);
nand U546 (N_546,In_191,In_283);
xor U547 (N_547,In_202,In_333);
xor U548 (N_548,In_2,In_235);
xor U549 (N_549,In_279,In_147);
and U550 (N_550,In_629,In_231);
or U551 (N_551,In_330,In_9);
and U552 (N_552,In_154,In_628);
nand U553 (N_553,In_286,In_743);
xnor U554 (N_554,In_663,In_616);
xnor U555 (N_555,In_435,In_205);
nor U556 (N_556,In_121,In_734);
nor U557 (N_557,In_452,In_596);
or U558 (N_558,In_113,In_380);
xnor U559 (N_559,In_665,In_179);
and U560 (N_560,In_75,In_515);
nand U561 (N_561,In_63,In_212);
or U562 (N_562,In_483,In_387);
or U563 (N_563,In_427,In_663);
or U564 (N_564,In_460,In_135);
xor U565 (N_565,In_26,In_86);
nor U566 (N_566,In_725,In_462);
nor U567 (N_567,In_642,In_195);
nand U568 (N_568,In_518,In_505);
xor U569 (N_569,In_467,In_571);
or U570 (N_570,In_266,In_132);
nor U571 (N_571,In_445,In_387);
xnor U572 (N_572,In_534,In_263);
or U573 (N_573,In_577,In_617);
xnor U574 (N_574,In_340,In_24);
or U575 (N_575,In_351,In_21);
nor U576 (N_576,In_504,In_136);
xnor U577 (N_577,In_512,In_680);
or U578 (N_578,In_595,In_55);
nor U579 (N_579,In_236,In_54);
xnor U580 (N_580,In_642,In_125);
and U581 (N_581,In_397,In_489);
and U582 (N_582,In_452,In_255);
xnor U583 (N_583,In_413,In_234);
nand U584 (N_584,In_18,In_95);
nor U585 (N_585,In_607,In_623);
and U586 (N_586,In_620,In_484);
and U587 (N_587,In_400,In_131);
and U588 (N_588,In_615,In_644);
nand U589 (N_589,In_606,In_665);
and U590 (N_590,In_293,In_499);
nor U591 (N_591,In_362,In_450);
nand U592 (N_592,In_523,In_109);
nor U593 (N_593,In_581,In_322);
or U594 (N_594,In_656,In_283);
or U595 (N_595,In_126,In_165);
nor U596 (N_596,In_494,In_537);
or U597 (N_597,In_748,In_384);
xor U598 (N_598,In_700,In_239);
or U599 (N_599,In_417,In_515);
xnor U600 (N_600,In_62,In_623);
nor U601 (N_601,In_649,In_291);
xor U602 (N_602,In_416,In_142);
and U603 (N_603,In_654,In_130);
nor U604 (N_604,In_738,In_127);
xnor U605 (N_605,In_393,In_674);
xnor U606 (N_606,In_73,In_392);
xor U607 (N_607,In_331,In_613);
nor U608 (N_608,In_1,In_480);
nor U609 (N_609,In_61,In_607);
or U610 (N_610,In_451,In_208);
nand U611 (N_611,In_188,In_401);
nand U612 (N_612,In_235,In_181);
or U613 (N_613,In_533,In_312);
and U614 (N_614,In_137,In_75);
and U615 (N_615,In_177,In_420);
or U616 (N_616,In_42,In_304);
or U617 (N_617,In_368,In_145);
nand U618 (N_618,In_570,In_655);
or U619 (N_619,In_249,In_24);
nand U620 (N_620,In_551,In_311);
nor U621 (N_621,In_200,In_671);
nand U622 (N_622,In_701,In_16);
nand U623 (N_623,In_593,In_735);
xor U624 (N_624,In_195,In_187);
nor U625 (N_625,In_498,In_149);
or U626 (N_626,In_124,In_47);
xnor U627 (N_627,In_70,In_276);
and U628 (N_628,In_569,In_393);
xnor U629 (N_629,In_682,In_186);
or U630 (N_630,In_550,In_349);
and U631 (N_631,In_379,In_90);
and U632 (N_632,In_565,In_510);
nor U633 (N_633,In_736,In_601);
xnor U634 (N_634,In_40,In_447);
nor U635 (N_635,In_203,In_424);
or U636 (N_636,In_555,In_653);
and U637 (N_637,In_116,In_344);
nand U638 (N_638,In_611,In_626);
nor U639 (N_639,In_350,In_380);
or U640 (N_640,In_652,In_602);
or U641 (N_641,In_104,In_424);
nand U642 (N_642,In_336,In_2);
nand U643 (N_643,In_419,In_367);
xor U644 (N_644,In_512,In_691);
xnor U645 (N_645,In_623,In_693);
and U646 (N_646,In_208,In_747);
and U647 (N_647,In_250,In_499);
and U648 (N_648,In_513,In_253);
nand U649 (N_649,In_565,In_459);
nand U650 (N_650,In_314,In_256);
and U651 (N_651,In_123,In_224);
or U652 (N_652,In_458,In_242);
nor U653 (N_653,In_189,In_481);
or U654 (N_654,In_212,In_520);
nor U655 (N_655,In_289,In_653);
xnor U656 (N_656,In_553,In_519);
nor U657 (N_657,In_119,In_536);
nand U658 (N_658,In_264,In_571);
xnor U659 (N_659,In_60,In_697);
and U660 (N_660,In_705,In_261);
and U661 (N_661,In_595,In_584);
or U662 (N_662,In_691,In_597);
nand U663 (N_663,In_68,In_29);
nor U664 (N_664,In_378,In_116);
and U665 (N_665,In_112,In_159);
and U666 (N_666,In_499,In_37);
or U667 (N_667,In_230,In_702);
nor U668 (N_668,In_208,In_352);
nor U669 (N_669,In_363,In_416);
xnor U670 (N_670,In_673,In_422);
and U671 (N_671,In_134,In_14);
nand U672 (N_672,In_282,In_101);
xor U673 (N_673,In_349,In_735);
nor U674 (N_674,In_227,In_343);
or U675 (N_675,In_254,In_298);
nand U676 (N_676,In_40,In_18);
xnor U677 (N_677,In_233,In_396);
nor U678 (N_678,In_299,In_31);
nor U679 (N_679,In_153,In_226);
nor U680 (N_680,In_528,In_676);
xor U681 (N_681,In_440,In_162);
or U682 (N_682,In_324,In_624);
and U683 (N_683,In_640,In_225);
and U684 (N_684,In_105,In_404);
xor U685 (N_685,In_235,In_697);
nor U686 (N_686,In_56,In_505);
or U687 (N_687,In_400,In_156);
xor U688 (N_688,In_132,In_571);
nand U689 (N_689,In_285,In_75);
nand U690 (N_690,In_652,In_495);
or U691 (N_691,In_272,In_303);
or U692 (N_692,In_408,In_403);
nand U693 (N_693,In_340,In_229);
and U694 (N_694,In_289,In_273);
and U695 (N_695,In_392,In_239);
nor U696 (N_696,In_654,In_574);
or U697 (N_697,In_269,In_47);
or U698 (N_698,In_735,In_599);
or U699 (N_699,In_32,In_723);
nand U700 (N_700,In_105,In_132);
nor U701 (N_701,In_530,In_649);
nor U702 (N_702,In_355,In_387);
xor U703 (N_703,In_29,In_386);
and U704 (N_704,In_319,In_123);
nor U705 (N_705,In_263,In_434);
nand U706 (N_706,In_435,In_1);
and U707 (N_707,In_156,In_676);
and U708 (N_708,In_478,In_168);
xnor U709 (N_709,In_317,In_620);
xnor U710 (N_710,In_147,In_439);
xor U711 (N_711,In_289,In_703);
nor U712 (N_712,In_690,In_414);
and U713 (N_713,In_560,In_528);
xnor U714 (N_714,In_287,In_525);
and U715 (N_715,In_528,In_31);
nand U716 (N_716,In_490,In_106);
or U717 (N_717,In_192,In_176);
and U718 (N_718,In_716,In_125);
xnor U719 (N_719,In_589,In_668);
and U720 (N_720,In_710,In_261);
or U721 (N_721,In_206,In_145);
nand U722 (N_722,In_432,In_565);
or U723 (N_723,In_540,In_2);
nand U724 (N_724,In_513,In_582);
nand U725 (N_725,In_552,In_586);
xor U726 (N_726,In_171,In_42);
and U727 (N_727,In_411,In_740);
and U728 (N_728,In_527,In_415);
nand U729 (N_729,In_434,In_129);
nand U730 (N_730,In_676,In_335);
or U731 (N_731,In_343,In_239);
or U732 (N_732,In_579,In_692);
and U733 (N_733,In_76,In_736);
nor U734 (N_734,In_127,In_708);
nand U735 (N_735,In_638,In_733);
xnor U736 (N_736,In_596,In_559);
or U737 (N_737,In_41,In_303);
xor U738 (N_738,In_625,In_487);
xnor U739 (N_739,In_686,In_285);
nor U740 (N_740,In_726,In_667);
nor U741 (N_741,In_304,In_615);
and U742 (N_742,In_407,In_343);
xor U743 (N_743,In_650,In_169);
and U744 (N_744,In_109,In_267);
xnor U745 (N_745,In_691,In_290);
xnor U746 (N_746,In_671,In_289);
nor U747 (N_747,In_448,In_594);
xor U748 (N_748,In_40,In_562);
and U749 (N_749,In_60,In_276);
nand U750 (N_750,In_398,In_89);
xnor U751 (N_751,In_205,In_110);
xnor U752 (N_752,In_730,In_474);
or U753 (N_753,In_27,In_105);
nor U754 (N_754,In_169,In_337);
or U755 (N_755,In_15,In_599);
or U756 (N_756,In_665,In_660);
xnor U757 (N_757,In_358,In_102);
nor U758 (N_758,In_353,In_626);
nor U759 (N_759,In_121,In_672);
xnor U760 (N_760,In_438,In_28);
or U761 (N_761,In_416,In_494);
nand U762 (N_762,In_208,In_581);
nand U763 (N_763,In_170,In_520);
and U764 (N_764,In_624,In_470);
nand U765 (N_765,In_160,In_72);
xor U766 (N_766,In_280,In_196);
or U767 (N_767,In_707,In_122);
or U768 (N_768,In_115,In_739);
nor U769 (N_769,In_377,In_221);
or U770 (N_770,In_708,In_419);
xnor U771 (N_771,In_54,In_423);
xnor U772 (N_772,In_321,In_255);
or U773 (N_773,In_511,In_644);
or U774 (N_774,In_630,In_613);
nor U775 (N_775,In_210,In_722);
xnor U776 (N_776,In_418,In_75);
nor U777 (N_777,In_383,In_76);
xor U778 (N_778,In_352,In_694);
and U779 (N_779,In_26,In_681);
xnor U780 (N_780,In_634,In_630);
xnor U781 (N_781,In_692,In_508);
xnor U782 (N_782,In_411,In_305);
nor U783 (N_783,In_646,In_115);
or U784 (N_784,In_360,In_744);
xnor U785 (N_785,In_398,In_513);
or U786 (N_786,In_684,In_27);
and U787 (N_787,In_525,In_91);
nor U788 (N_788,In_405,In_192);
nand U789 (N_789,In_253,In_322);
nor U790 (N_790,In_693,In_671);
xor U791 (N_791,In_118,In_258);
nand U792 (N_792,In_380,In_643);
nor U793 (N_793,In_102,In_656);
xnor U794 (N_794,In_304,In_484);
nor U795 (N_795,In_219,In_212);
xnor U796 (N_796,In_328,In_329);
xnor U797 (N_797,In_145,In_477);
and U798 (N_798,In_260,In_161);
and U799 (N_799,In_299,In_21);
nand U800 (N_800,In_61,In_656);
nor U801 (N_801,In_116,In_62);
and U802 (N_802,In_257,In_380);
or U803 (N_803,In_269,In_578);
or U804 (N_804,In_218,In_149);
and U805 (N_805,In_33,In_631);
nand U806 (N_806,In_31,In_186);
or U807 (N_807,In_66,In_520);
nor U808 (N_808,In_448,In_289);
and U809 (N_809,In_163,In_420);
and U810 (N_810,In_423,In_118);
xor U811 (N_811,In_269,In_353);
nor U812 (N_812,In_54,In_576);
or U813 (N_813,In_214,In_166);
or U814 (N_814,In_139,In_592);
xor U815 (N_815,In_310,In_593);
nand U816 (N_816,In_117,In_641);
xor U817 (N_817,In_455,In_516);
and U818 (N_818,In_682,In_453);
xnor U819 (N_819,In_5,In_74);
and U820 (N_820,In_398,In_10);
and U821 (N_821,In_200,In_729);
or U822 (N_822,In_406,In_455);
and U823 (N_823,In_536,In_198);
nand U824 (N_824,In_454,In_349);
xnor U825 (N_825,In_461,In_280);
nand U826 (N_826,In_149,In_111);
or U827 (N_827,In_79,In_296);
or U828 (N_828,In_24,In_182);
xnor U829 (N_829,In_676,In_179);
nand U830 (N_830,In_481,In_27);
or U831 (N_831,In_7,In_577);
nand U832 (N_832,In_276,In_49);
xor U833 (N_833,In_571,In_331);
and U834 (N_834,In_720,In_237);
or U835 (N_835,In_43,In_518);
xor U836 (N_836,In_44,In_581);
and U837 (N_837,In_572,In_514);
or U838 (N_838,In_416,In_193);
or U839 (N_839,In_530,In_484);
or U840 (N_840,In_416,In_589);
nand U841 (N_841,In_393,In_433);
nor U842 (N_842,In_105,In_397);
nor U843 (N_843,In_529,In_227);
nand U844 (N_844,In_349,In_117);
and U845 (N_845,In_76,In_748);
xor U846 (N_846,In_535,In_530);
nor U847 (N_847,In_720,In_489);
and U848 (N_848,In_223,In_416);
or U849 (N_849,In_456,In_534);
xor U850 (N_850,In_486,In_451);
nor U851 (N_851,In_315,In_98);
nor U852 (N_852,In_393,In_118);
nand U853 (N_853,In_707,In_490);
or U854 (N_854,In_308,In_543);
nor U855 (N_855,In_464,In_85);
xnor U856 (N_856,In_730,In_414);
nand U857 (N_857,In_243,In_90);
nand U858 (N_858,In_696,In_441);
and U859 (N_859,In_667,In_584);
or U860 (N_860,In_568,In_46);
and U861 (N_861,In_549,In_260);
and U862 (N_862,In_415,In_252);
xor U863 (N_863,In_671,In_198);
or U864 (N_864,In_395,In_514);
nand U865 (N_865,In_292,In_5);
xor U866 (N_866,In_479,In_384);
xor U867 (N_867,In_302,In_490);
nor U868 (N_868,In_699,In_199);
or U869 (N_869,In_107,In_84);
nand U870 (N_870,In_258,In_247);
and U871 (N_871,In_78,In_366);
and U872 (N_872,In_545,In_232);
nand U873 (N_873,In_721,In_749);
nand U874 (N_874,In_173,In_605);
and U875 (N_875,In_211,In_630);
and U876 (N_876,In_291,In_11);
or U877 (N_877,In_224,In_370);
nand U878 (N_878,In_514,In_643);
nor U879 (N_879,In_440,In_114);
xnor U880 (N_880,In_541,In_455);
xnor U881 (N_881,In_748,In_455);
xor U882 (N_882,In_240,In_353);
nor U883 (N_883,In_375,In_726);
nand U884 (N_884,In_147,In_186);
and U885 (N_885,In_68,In_333);
and U886 (N_886,In_201,In_154);
or U887 (N_887,In_186,In_79);
xor U888 (N_888,In_213,In_575);
or U889 (N_889,In_539,In_309);
or U890 (N_890,In_396,In_142);
nor U891 (N_891,In_601,In_632);
or U892 (N_892,In_603,In_145);
xor U893 (N_893,In_21,In_25);
and U894 (N_894,In_117,In_549);
or U895 (N_895,In_534,In_652);
and U896 (N_896,In_160,In_491);
nor U897 (N_897,In_213,In_216);
nor U898 (N_898,In_726,In_24);
or U899 (N_899,In_238,In_288);
nand U900 (N_900,In_18,In_459);
xor U901 (N_901,In_661,In_693);
nand U902 (N_902,In_77,In_55);
and U903 (N_903,In_462,In_749);
xnor U904 (N_904,In_62,In_13);
xnor U905 (N_905,In_365,In_195);
nand U906 (N_906,In_730,In_40);
nand U907 (N_907,In_449,In_575);
or U908 (N_908,In_435,In_300);
nand U909 (N_909,In_712,In_57);
and U910 (N_910,In_651,In_602);
nand U911 (N_911,In_128,In_206);
xnor U912 (N_912,In_265,In_385);
nand U913 (N_913,In_590,In_259);
or U914 (N_914,In_113,In_594);
or U915 (N_915,In_79,In_646);
or U916 (N_916,In_596,In_502);
or U917 (N_917,In_704,In_646);
nor U918 (N_918,In_185,In_548);
and U919 (N_919,In_220,In_659);
and U920 (N_920,In_71,In_362);
nor U921 (N_921,In_82,In_600);
and U922 (N_922,In_142,In_181);
or U923 (N_923,In_667,In_102);
nand U924 (N_924,In_299,In_150);
or U925 (N_925,In_648,In_497);
nand U926 (N_926,In_633,In_700);
and U927 (N_927,In_494,In_356);
or U928 (N_928,In_680,In_8);
nor U929 (N_929,In_465,In_484);
nand U930 (N_930,In_2,In_735);
nor U931 (N_931,In_193,In_513);
nor U932 (N_932,In_344,In_164);
or U933 (N_933,In_388,In_227);
nand U934 (N_934,In_382,In_655);
nor U935 (N_935,In_271,In_584);
nand U936 (N_936,In_239,In_559);
or U937 (N_937,In_154,In_225);
xor U938 (N_938,In_315,In_94);
and U939 (N_939,In_188,In_296);
nand U940 (N_940,In_649,In_729);
or U941 (N_941,In_465,In_449);
or U942 (N_942,In_282,In_249);
xnor U943 (N_943,In_234,In_124);
nand U944 (N_944,In_507,In_42);
xor U945 (N_945,In_361,In_347);
and U946 (N_946,In_200,In_429);
nor U947 (N_947,In_355,In_197);
or U948 (N_948,In_209,In_423);
xor U949 (N_949,In_696,In_327);
xnor U950 (N_950,In_96,In_633);
xor U951 (N_951,In_20,In_571);
or U952 (N_952,In_416,In_154);
nor U953 (N_953,In_413,In_3);
nand U954 (N_954,In_460,In_215);
nor U955 (N_955,In_556,In_577);
xnor U956 (N_956,In_159,In_58);
xor U957 (N_957,In_363,In_580);
xnor U958 (N_958,In_577,In_379);
or U959 (N_959,In_422,In_530);
and U960 (N_960,In_337,In_551);
nor U961 (N_961,In_496,In_295);
or U962 (N_962,In_500,In_322);
or U963 (N_963,In_534,In_452);
xnor U964 (N_964,In_665,In_326);
xor U965 (N_965,In_3,In_227);
or U966 (N_966,In_398,In_579);
nand U967 (N_967,In_694,In_651);
or U968 (N_968,In_630,In_56);
nand U969 (N_969,In_548,In_734);
and U970 (N_970,In_364,In_318);
xnor U971 (N_971,In_459,In_82);
nor U972 (N_972,In_314,In_126);
or U973 (N_973,In_402,In_3);
nor U974 (N_974,In_299,In_189);
or U975 (N_975,In_681,In_388);
nor U976 (N_976,In_476,In_615);
and U977 (N_977,In_511,In_115);
xnor U978 (N_978,In_381,In_332);
nor U979 (N_979,In_71,In_659);
and U980 (N_980,In_628,In_525);
or U981 (N_981,In_540,In_312);
and U982 (N_982,In_61,In_539);
xor U983 (N_983,In_470,In_474);
xor U984 (N_984,In_426,In_146);
and U985 (N_985,In_232,In_88);
nand U986 (N_986,In_220,In_561);
xnor U987 (N_987,In_729,In_533);
xnor U988 (N_988,In_374,In_320);
and U989 (N_989,In_483,In_472);
and U990 (N_990,In_560,In_202);
and U991 (N_991,In_215,In_633);
xnor U992 (N_992,In_75,In_725);
or U993 (N_993,In_556,In_525);
or U994 (N_994,In_267,In_365);
and U995 (N_995,In_249,In_447);
xor U996 (N_996,In_714,In_177);
nor U997 (N_997,In_548,In_746);
xor U998 (N_998,In_284,In_603);
and U999 (N_999,In_420,In_207);
and U1000 (N_1000,In_307,In_722);
xor U1001 (N_1001,In_702,In_643);
nor U1002 (N_1002,In_206,In_688);
xnor U1003 (N_1003,In_125,In_24);
xor U1004 (N_1004,In_326,In_519);
and U1005 (N_1005,In_696,In_500);
xnor U1006 (N_1006,In_26,In_40);
and U1007 (N_1007,In_684,In_708);
xor U1008 (N_1008,In_718,In_478);
nor U1009 (N_1009,In_91,In_371);
nand U1010 (N_1010,In_138,In_186);
or U1011 (N_1011,In_357,In_140);
nor U1012 (N_1012,In_487,In_520);
xnor U1013 (N_1013,In_157,In_431);
xor U1014 (N_1014,In_579,In_520);
nand U1015 (N_1015,In_115,In_168);
xnor U1016 (N_1016,In_24,In_185);
nand U1017 (N_1017,In_385,In_614);
nand U1018 (N_1018,In_165,In_247);
nand U1019 (N_1019,In_299,In_30);
nor U1020 (N_1020,In_585,In_265);
and U1021 (N_1021,In_264,In_259);
and U1022 (N_1022,In_500,In_387);
xnor U1023 (N_1023,In_332,In_410);
nor U1024 (N_1024,In_390,In_384);
or U1025 (N_1025,In_729,In_199);
nor U1026 (N_1026,In_651,In_428);
and U1027 (N_1027,In_260,In_453);
nand U1028 (N_1028,In_184,In_115);
and U1029 (N_1029,In_691,In_277);
and U1030 (N_1030,In_20,In_541);
nand U1031 (N_1031,In_409,In_522);
nor U1032 (N_1032,In_334,In_77);
nand U1033 (N_1033,In_496,In_8);
or U1034 (N_1034,In_463,In_206);
xnor U1035 (N_1035,In_27,In_597);
and U1036 (N_1036,In_530,In_209);
nand U1037 (N_1037,In_25,In_517);
or U1038 (N_1038,In_306,In_441);
nor U1039 (N_1039,In_595,In_226);
or U1040 (N_1040,In_532,In_451);
nor U1041 (N_1041,In_345,In_489);
nand U1042 (N_1042,In_143,In_475);
and U1043 (N_1043,In_64,In_554);
or U1044 (N_1044,In_387,In_185);
nand U1045 (N_1045,In_748,In_580);
or U1046 (N_1046,In_270,In_306);
and U1047 (N_1047,In_642,In_235);
nand U1048 (N_1048,In_553,In_325);
nand U1049 (N_1049,In_635,In_64);
xnor U1050 (N_1050,In_576,In_528);
and U1051 (N_1051,In_305,In_568);
nor U1052 (N_1052,In_271,In_561);
and U1053 (N_1053,In_527,In_47);
nor U1054 (N_1054,In_55,In_238);
nand U1055 (N_1055,In_0,In_317);
and U1056 (N_1056,In_169,In_525);
nand U1057 (N_1057,In_69,In_302);
xor U1058 (N_1058,In_118,In_602);
xor U1059 (N_1059,In_606,In_745);
xnor U1060 (N_1060,In_545,In_650);
nand U1061 (N_1061,In_476,In_300);
and U1062 (N_1062,In_182,In_731);
and U1063 (N_1063,In_269,In_581);
xnor U1064 (N_1064,In_479,In_239);
nor U1065 (N_1065,In_614,In_395);
nand U1066 (N_1066,In_261,In_35);
xnor U1067 (N_1067,In_182,In_308);
and U1068 (N_1068,In_662,In_737);
xnor U1069 (N_1069,In_693,In_740);
or U1070 (N_1070,In_526,In_438);
nor U1071 (N_1071,In_552,In_515);
and U1072 (N_1072,In_475,In_95);
nand U1073 (N_1073,In_124,In_59);
xor U1074 (N_1074,In_233,In_494);
nor U1075 (N_1075,In_449,In_189);
or U1076 (N_1076,In_312,In_667);
nand U1077 (N_1077,In_307,In_389);
xnor U1078 (N_1078,In_279,In_156);
or U1079 (N_1079,In_329,In_636);
nand U1080 (N_1080,In_538,In_691);
nand U1081 (N_1081,In_546,In_86);
nand U1082 (N_1082,In_201,In_381);
nand U1083 (N_1083,In_35,In_699);
and U1084 (N_1084,In_389,In_334);
or U1085 (N_1085,In_223,In_710);
xor U1086 (N_1086,In_522,In_518);
nor U1087 (N_1087,In_492,In_725);
or U1088 (N_1088,In_198,In_138);
and U1089 (N_1089,In_302,In_26);
nand U1090 (N_1090,In_517,In_48);
xor U1091 (N_1091,In_554,In_563);
and U1092 (N_1092,In_713,In_608);
nor U1093 (N_1093,In_562,In_130);
nor U1094 (N_1094,In_637,In_742);
xnor U1095 (N_1095,In_520,In_659);
xnor U1096 (N_1096,In_410,In_623);
nor U1097 (N_1097,In_723,In_97);
or U1098 (N_1098,In_506,In_624);
xor U1099 (N_1099,In_614,In_468);
and U1100 (N_1100,In_493,In_11);
nand U1101 (N_1101,In_67,In_65);
and U1102 (N_1102,In_87,In_262);
and U1103 (N_1103,In_402,In_224);
or U1104 (N_1104,In_367,In_578);
nand U1105 (N_1105,In_238,In_365);
nor U1106 (N_1106,In_624,In_328);
nor U1107 (N_1107,In_698,In_498);
nand U1108 (N_1108,In_36,In_372);
and U1109 (N_1109,In_493,In_208);
xnor U1110 (N_1110,In_47,In_670);
and U1111 (N_1111,In_204,In_448);
xor U1112 (N_1112,In_455,In_153);
xnor U1113 (N_1113,In_743,In_88);
nand U1114 (N_1114,In_52,In_638);
or U1115 (N_1115,In_3,In_102);
xor U1116 (N_1116,In_679,In_624);
nand U1117 (N_1117,In_58,In_203);
or U1118 (N_1118,In_237,In_254);
nand U1119 (N_1119,In_338,In_356);
and U1120 (N_1120,In_329,In_709);
xor U1121 (N_1121,In_134,In_576);
or U1122 (N_1122,In_484,In_140);
or U1123 (N_1123,In_129,In_225);
nand U1124 (N_1124,In_257,In_602);
xnor U1125 (N_1125,In_613,In_654);
xnor U1126 (N_1126,In_160,In_715);
nor U1127 (N_1127,In_388,In_547);
nand U1128 (N_1128,In_52,In_413);
xnor U1129 (N_1129,In_549,In_320);
or U1130 (N_1130,In_627,In_25);
or U1131 (N_1131,In_345,In_140);
nand U1132 (N_1132,In_138,In_407);
or U1133 (N_1133,In_94,In_85);
and U1134 (N_1134,In_739,In_655);
nand U1135 (N_1135,In_138,In_454);
or U1136 (N_1136,In_309,In_408);
nor U1137 (N_1137,In_268,In_11);
nor U1138 (N_1138,In_228,In_439);
or U1139 (N_1139,In_524,In_403);
xnor U1140 (N_1140,In_476,In_106);
or U1141 (N_1141,In_149,In_549);
nor U1142 (N_1142,In_647,In_493);
nand U1143 (N_1143,In_522,In_649);
or U1144 (N_1144,In_320,In_738);
xnor U1145 (N_1145,In_74,In_201);
and U1146 (N_1146,In_554,In_666);
and U1147 (N_1147,In_137,In_725);
nand U1148 (N_1148,In_69,In_33);
and U1149 (N_1149,In_564,In_555);
xnor U1150 (N_1150,In_442,In_742);
nand U1151 (N_1151,In_247,In_720);
nand U1152 (N_1152,In_697,In_414);
xor U1153 (N_1153,In_335,In_127);
nand U1154 (N_1154,In_487,In_7);
nor U1155 (N_1155,In_314,In_53);
or U1156 (N_1156,In_374,In_17);
and U1157 (N_1157,In_169,In_54);
and U1158 (N_1158,In_339,In_688);
nor U1159 (N_1159,In_227,In_729);
nand U1160 (N_1160,In_188,In_63);
nand U1161 (N_1161,In_29,In_683);
xor U1162 (N_1162,In_611,In_590);
xnor U1163 (N_1163,In_710,In_501);
xor U1164 (N_1164,In_590,In_451);
nand U1165 (N_1165,In_350,In_46);
nand U1166 (N_1166,In_649,In_423);
or U1167 (N_1167,In_735,In_75);
xnor U1168 (N_1168,In_368,In_27);
nand U1169 (N_1169,In_683,In_706);
nand U1170 (N_1170,In_599,In_721);
nand U1171 (N_1171,In_146,In_733);
nor U1172 (N_1172,In_634,In_160);
nor U1173 (N_1173,In_526,In_512);
or U1174 (N_1174,In_227,In_177);
nand U1175 (N_1175,In_600,In_319);
and U1176 (N_1176,In_109,In_275);
and U1177 (N_1177,In_273,In_295);
and U1178 (N_1178,In_577,In_220);
xnor U1179 (N_1179,In_58,In_527);
nor U1180 (N_1180,In_579,In_616);
xnor U1181 (N_1181,In_26,In_652);
xnor U1182 (N_1182,In_596,In_363);
nand U1183 (N_1183,In_399,In_62);
nand U1184 (N_1184,In_709,In_86);
and U1185 (N_1185,In_81,In_409);
or U1186 (N_1186,In_543,In_547);
nor U1187 (N_1187,In_172,In_605);
or U1188 (N_1188,In_641,In_209);
nor U1189 (N_1189,In_187,In_227);
nor U1190 (N_1190,In_36,In_313);
or U1191 (N_1191,In_567,In_521);
nand U1192 (N_1192,In_125,In_478);
xor U1193 (N_1193,In_723,In_72);
or U1194 (N_1194,In_19,In_49);
xor U1195 (N_1195,In_383,In_70);
nand U1196 (N_1196,In_683,In_256);
and U1197 (N_1197,In_174,In_409);
nor U1198 (N_1198,In_734,In_361);
or U1199 (N_1199,In_259,In_95);
nand U1200 (N_1200,In_213,In_594);
nand U1201 (N_1201,In_530,In_235);
xor U1202 (N_1202,In_232,In_105);
xor U1203 (N_1203,In_5,In_654);
nor U1204 (N_1204,In_682,In_734);
nor U1205 (N_1205,In_155,In_551);
nor U1206 (N_1206,In_399,In_379);
and U1207 (N_1207,In_588,In_488);
nand U1208 (N_1208,In_297,In_73);
xor U1209 (N_1209,In_153,In_444);
xnor U1210 (N_1210,In_441,In_12);
nand U1211 (N_1211,In_65,In_190);
xnor U1212 (N_1212,In_257,In_41);
and U1213 (N_1213,In_148,In_430);
nor U1214 (N_1214,In_137,In_191);
nor U1215 (N_1215,In_721,In_355);
or U1216 (N_1216,In_365,In_258);
nor U1217 (N_1217,In_625,In_443);
nor U1218 (N_1218,In_365,In_544);
nor U1219 (N_1219,In_529,In_308);
xnor U1220 (N_1220,In_189,In_441);
and U1221 (N_1221,In_54,In_147);
nor U1222 (N_1222,In_489,In_561);
and U1223 (N_1223,In_326,In_749);
or U1224 (N_1224,In_180,In_746);
xnor U1225 (N_1225,In_260,In_293);
xor U1226 (N_1226,In_362,In_637);
or U1227 (N_1227,In_572,In_617);
xor U1228 (N_1228,In_516,In_63);
or U1229 (N_1229,In_379,In_283);
and U1230 (N_1230,In_22,In_285);
or U1231 (N_1231,In_685,In_202);
or U1232 (N_1232,In_459,In_238);
or U1233 (N_1233,In_568,In_44);
or U1234 (N_1234,In_447,In_452);
xor U1235 (N_1235,In_392,In_573);
and U1236 (N_1236,In_701,In_139);
and U1237 (N_1237,In_65,In_266);
nor U1238 (N_1238,In_148,In_205);
and U1239 (N_1239,In_92,In_30);
nor U1240 (N_1240,In_645,In_494);
and U1241 (N_1241,In_459,In_686);
and U1242 (N_1242,In_277,In_161);
nor U1243 (N_1243,In_700,In_561);
and U1244 (N_1244,In_377,In_680);
xnor U1245 (N_1245,In_146,In_39);
nor U1246 (N_1246,In_262,In_606);
nor U1247 (N_1247,In_554,In_235);
xor U1248 (N_1248,In_601,In_94);
and U1249 (N_1249,In_421,In_274);
nand U1250 (N_1250,In_121,In_48);
xnor U1251 (N_1251,In_677,In_680);
nor U1252 (N_1252,In_696,In_7);
nor U1253 (N_1253,In_144,In_220);
nor U1254 (N_1254,In_403,In_529);
or U1255 (N_1255,In_319,In_363);
xor U1256 (N_1256,In_185,In_573);
nor U1257 (N_1257,In_109,In_119);
nand U1258 (N_1258,In_714,In_311);
xnor U1259 (N_1259,In_349,In_55);
nor U1260 (N_1260,In_202,In_111);
or U1261 (N_1261,In_258,In_472);
and U1262 (N_1262,In_360,In_666);
or U1263 (N_1263,In_325,In_68);
nor U1264 (N_1264,In_259,In_458);
and U1265 (N_1265,In_677,In_391);
nand U1266 (N_1266,In_452,In_94);
or U1267 (N_1267,In_524,In_7);
nand U1268 (N_1268,In_463,In_159);
nand U1269 (N_1269,In_239,In_641);
nor U1270 (N_1270,In_682,In_197);
nand U1271 (N_1271,In_436,In_474);
and U1272 (N_1272,In_628,In_617);
xor U1273 (N_1273,In_328,In_585);
nand U1274 (N_1274,In_625,In_490);
and U1275 (N_1275,In_704,In_113);
or U1276 (N_1276,In_193,In_595);
or U1277 (N_1277,In_406,In_618);
and U1278 (N_1278,In_283,In_582);
and U1279 (N_1279,In_134,In_32);
nand U1280 (N_1280,In_242,In_238);
xor U1281 (N_1281,In_455,In_53);
or U1282 (N_1282,In_169,In_460);
nor U1283 (N_1283,In_60,In_262);
xnor U1284 (N_1284,In_128,In_572);
and U1285 (N_1285,In_440,In_286);
or U1286 (N_1286,In_259,In_685);
xnor U1287 (N_1287,In_296,In_546);
and U1288 (N_1288,In_651,In_388);
and U1289 (N_1289,In_534,In_528);
and U1290 (N_1290,In_237,In_22);
or U1291 (N_1291,In_257,In_181);
or U1292 (N_1292,In_185,In_732);
nand U1293 (N_1293,In_317,In_26);
nand U1294 (N_1294,In_149,In_596);
or U1295 (N_1295,In_523,In_160);
or U1296 (N_1296,In_390,In_258);
and U1297 (N_1297,In_492,In_546);
or U1298 (N_1298,In_339,In_744);
and U1299 (N_1299,In_579,In_488);
nor U1300 (N_1300,In_655,In_231);
xor U1301 (N_1301,In_83,In_267);
or U1302 (N_1302,In_675,In_411);
nand U1303 (N_1303,In_327,In_124);
xor U1304 (N_1304,In_387,In_563);
and U1305 (N_1305,In_647,In_225);
or U1306 (N_1306,In_415,In_580);
and U1307 (N_1307,In_420,In_521);
nor U1308 (N_1308,In_678,In_478);
or U1309 (N_1309,In_253,In_155);
nand U1310 (N_1310,In_397,In_372);
nor U1311 (N_1311,In_196,In_37);
or U1312 (N_1312,In_235,In_585);
nand U1313 (N_1313,In_375,In_730);
nor U1314 (N_1314,In_528,In_431);
and U1315 (N_1315,In_543,In_82);
or U1316 (N_1316,In_488,In_85);
and U1317 (N_1317,In_128,In_607);
nor U1318 (N_1318,In_474,In_266);
nor U1319 (N_1319,In_296,In_520);
nor U1320 (N_1320,In_581,In_704);
nor U1321 (N_1321,In_228,In_188);
xnor U1322 (N_1322,In_499,In_221);
nor U1323 (N_1323,In_144,In_101);
xnor U1324 (N_1324,In_155,In_477);
nand U1325 (N_1325,In_724,In_517);
and U1326 (N_1326,In_708,In_7);
xnor U1327 (N_1327,In_536,In_100);
nor U1328 (N_1328,In_40,In_459);
and U1329 (N_1329,In_360,In_652);
xnor U1330 (N_1330,In_176,In_715);
xor U1331 (N_1331,In_6,In_224);
xor U1332 (N_1332,In_691,In_8);
nand U1333 (N_1333,In_24,In_277);
and U1334 (N_1334,In_103,In_537);
nor U1335 (N_1335,In_177,In_97);
and U1336 (N_1336,In_397,In_119);
nand U1337 (N_1337,In_600,In_211);
nor U1338 (N_1338,In_443,In_218);
xnor U1339 (N_1339,In_652,In_660);
nor U1340 (N_1340,In_368,In_455);
and U1341 (N_1341,In_254,In_336);
or U1342 (N_1342,In_26,In_542);
or U1343 (N_1343,In_139,In_137);
and U1344 (N_1344,In_258,In_90);
or U1345 (N_1345,In_2,In_102);
nor U1346 (N_1346,In_155,In_360);
xnor U1347 (N_1347,In_730,In_285);
or U1348 (N_1348,In_30,In_366);
nand U1349 (N_1349,In_258,In_716);
xnor U1350 (N_1350,In_397,In_308);
and U1351 (N_1351,In_625,In_261);
xor U1352 (N_1352,In_77,In_449);
xor U1353 (N_1353,In_384,In_598);
and U1354 (N_1354,In_682,In_570);
xnor U1355 (N_1355,In_721,In_625);
nor U1356 (N_1356,In_315,In_680);
and U1357 (N_1357,In_661,In_544);
xor U1358 (N_1358,In_397,In_326);
xor U1359 (N_1359,In_59,In_87);
nand U1360 (N_1360,In_263,In_258);
or U1361 (N_1361,In_324,In_200);
or U1362 (N_1362,In_663,In_408);
and U1363 (N_1363,In_641,In_394);
nand U1364 (N_1364,In_267,In_78);
xnor U1365 (N_1365,In_622,In_223);
nor U1366 (N_1366,In_268,In_113);
or U1367 (N_1367,In_416,In_68);
nand U1368 (N_1368,In_472,In_599);
nor U1369 (N_1369,In_185,In_441);
nand U1370 (N_1370,In_71,In_651);
and U1371 (N_1371,In_91,In_147);
nand U1372 (N_1372,In_32,In_395);
xnor U1373 (N_1373,In_570,In_692);
nor U1374 (N_1374,In_483,In_590);
nor U1375 (N_1375,In_443,In_395);
and U1376 (N_1376,In_190,In_466);
nor U1377 (N_1377,In_319,In_514);
or U1378 (N_1378,In_547,In_586);
and U1379 (N_1379,In_97,In_376);
nor U1380 (N_1380,In_578,In_225);
xor U1381 (N_1381,In_65,In_69);
and U1382 (N_1382,In_732,In_388);
nand U1383 (N_1383,In_227,In_178);
nor U1384 (N_1384,In_80,In_23);
nand U1385 (N_1385,In_688,In_515);
xor U1386 (N_1386,In_22,In_473);
and U1387 (N_1387,In_274,In_222);
or U1388 (N_1388,In_190,In_214);
nor U1389 (N_1389,In_281,In_682);
nor U1390 (N_1390,In_149,In_410);
nand U1391 (N_1391,In_180,In_331);
xnor U1392 (N_1392,In_711,In_420);
or U1393 (N_1393,In_97,In_327);
nor U1394 (N_1394,In_657,In_592);
and U1395 (N_1395,In_445,In_571);
and U1396 (N_1396,In_324,In_269);
nor U1397 (N_1397,In_111,In_467);
xor U1398 (N_1398,In_206,In_654);
nor U1399 (N_1399,In_81,In_122);
xor U1400 (N_1400,In_476,In_26);
xor U1401 (N_1401,In_153,In_181);
nor U1402 (N_1402,In_628,In_658);
nand U1403 (N_1403,In_564,In_130);
nand U1404 (N_1404,In_118,In_199);
xnor U1405 (N_1405,In_547,In_260);
and U1406 (N_1406,In_114,In_8);
xnor U1407 (N_1407,In_552,In_517);
nor U1408 (N_1408,In_146,In_161);
nor U1409 (N_1409,In_500,In_299);
nand U1410 (N_1410,In_225,In_747);
nor U1411 (N_1411,In_288,In_378);
and U1412 (N_1412,In_602,In_698);
xor U1413 (N_1413,In_313,In_334);
xnor U1414 (N_1414,In_443,In_656);
and U1415 (N_1415,In_688,In_432);
nor U1416 (N_1416,In_599,In_78);
nand U1417 (N_1417,In_508,In_734);
xor U1418 (N_1418,In_454,In_190);
nand U1419 (N_1419,In_83,In_573);
or U1420 (N_1420,In_515,In_652);
and U1421 (N_1421,In_524,In_743);
nand U1422 (N_1422,In_673,In_568);
xnor U1423 (N_1423,In_631,In_665);
and U1424 (N_1424,In_77,In_9);
nand U1425 (N_1425,In_271,In_424);
and U1426 (N_1426,In_196,In_666);
and U1427 (N_1427,In_348,In_554);
nand U1428 (N_1428,In_536,In_159);
xnor U1429 (N_1429,In_561,In_11);
nor U1430 (N_1430,In_583,In_616);
xnor U1431 (N_1431,In_598,In_339);
or U1432 (N_1432,In_253,In_275);
or U1433 (N_1433,In_667,In_585);
and U1434 (N_1434,In_606,In_452);
nand U1435 (N_1435,In_697,In_66);
and U1436 (N_1436,In_668,In_715);
or U1437 (N_1437,In_594,In_677);
xor U1438 (N_1438,In_121,In_189);
and U1439 (N_1439,In_743,In_694);
nand U1440 (N_1440,In_723,In_136);
and U1441 (N_1441,In_247,In_743);
and U1442 (N_1442,In_112,In_99);
or U1443 (N_1443,In_403,In_509);
or U1444 (N_1444,In_206,In_429);
xnor U1445 (N_1445,In_185,In_486);
or U1446 (N_1446,In_330,In_332);
and U1447 (N_1447,In_468,In_195);
or U1448 (N_1448,In_245,In_588);
nand U1449 (N_1449,In_729,In_405);
xor U1450 (N_1450,In_582,In_238);
and U1451 (N_1451,In_132,In_9);
nand U1452 (N_1452,In_238,In_631);
xor U1453 (N_1453,In_712,In_374);
nor U1454 (N_1454,In_556,In_357);
nor U1455 (N_1455,In_639,In_688);
xnor U1456 (N_1456,In_674,In_449);
and U1457 (N_1457,In_377,In_233);
nor U1458 (N_1458,In_235,In_96);
and U1459 (N_1459,In_232,In_399);
xor U1460 (N_1460,In_612,In_2);
and U1461 (N_1461,In_257,In_710);
xnor U1462 (N_1462,In_519,In_170);
and U1463 (N_1463,In_257,In_653);
and U1464 (N_1464,In_441,In_112);
and U1465 (N_1465,In_713,In_609);
nor U1466 (N_1466,In_127,In_401);
or U1467 (N_1467,In_150,In_692);
and U1468 (N_1468,In_398,In_638);
nor U1469 (N_1469,In_620,In_75);
nand U1470 (N_1470,In_623,In_532);
or U1471 (N_1471,In_449,In_269);
nand U1472 (N_1472,In_234,In_122);
nand U1473 (N_1473,In_2,In_166);
nor U1474 (N_1474,In_550,In_677);
or U1475 (N_1475,In_309,In_602);
and U1476 (N_1476,In_290,In_253);
xor U1477 (N_1477,In_748,In_199);
nand U1478 (N_1478,In_48,In_208);
and U1479 (N_1479,In_200,In_92);
and U1480 (N_1480,In_556,In_495);
nor U1481 (N_1481,In_314,In_396);
or U1482 (N_1482,In_568,In_328);
xor U1483 (N_1483,In_715,In_675);
and U1484 (N_1484,In_14,In_404);
nand U1485 (N_1485,In_519,In_165);
or U1486 (N_1486,In_552,In_519);
nor U1487 (N_1487,In_299,In_195);
xnor U1488 (N_1488,In_628,In_673);
nand U1489 (N_1489,In_267,In_392);
or U1490 (N_1490,In_373,In_35);
and U1491 (N_1491,In_318,In_67);
or U1492 (N_1492,In_380,In_31);
and U1493 (N_1493,In_45,In_538);
or U1494 (N_1494,In_511,In_604);
nand U1495 (N_1495,In_91,In_197);
and U1496 (N_1496,In_382,In_61);
nor U1497 (N_1497,In_251,In_563);
and U1498 (N_1498,In_605,In_440);
or U1499 (N_1499,In_39,In_74);
nor U1500 (N_1500,In_46,In_122);
and U1501 (N_1501,In_170,In_555);
xor U1502 (N_1502,In_724,In_161);
nor U1503 (N_1503,In_673,In_48);
nor U1504 (N_1504,In_693,In_147);
xor U1505 (N_1505,In_410,In_312);
nor U1506 (N_1506,In_513,In_293);
and U1507 (N_1507,In_625,In_371);
nand U1508 (N_1508,In_310,In_286);
and U1509 (N_1509,In_285,In_53);
and U1510 (N_1510,In_524,In_157);
and U1511 (N_1511,In_653,In_706);
or U1512 (N_1512,In_481,In_325);
xnor U1513 (N_1513,In_494,In_729);
nor U1514 (N_1514,In_20,In_538);
and U1515 (N_1515,In_590,In_561);
xnor U1516 (N_1516,In_146,In_93);
nor U1517 (N_1517,In_673,In_326);
and U1518 (N_1518,In_257,In_637);
nor U1519 (N_1519,In_100,In_431);
xnor U1520 (N_1520,In_661,In_378);
nor U1521 (N_1521,In_371,In_6);
nand U1522 (N_1522,In_126,In_675);
and U1523 (N_1523,In_10,In_489);
xnor U1524 (N_1524,In_639,In_186);
xor U1525 (N_1525,In_597,In_524);
xor U1526 (N_1526,In_643,In_330);
nand U1527 (N_1527,In_127,In_439);
xor U1528 (N_1528,In_372,In_82);
or U1529 (N_1529,In_449,In_217);
and U1530 (N_1530,In_41,In_668);
xnor U1531 (N_1531,In_447,In_24);
and U1532 (N_1532,In_477,In_505);
and U1533 (N_1533,In_610,In_175);
or U1534 (N_1534,In_462,In_646);
nand U1535 (N_1535,In_279,In_375);
nand U1536 (N_1536,In_646,In_147);
xor U1537 (N_1537,In_558,In_404);
nor U1538 (N_1538,In_375,In_457);
nor U1539 (N_1539,In_78,In_363);
and U1540 (N_1540,In_21,In_180);
xor U1541 (N_1541,In_230,In_10);
xnor U1542 (N_1542,In_726,In_527);
or U1543 (N_1543,In_331,In_722);
xnor U1544 (N_1544,In_205,In_545);
xor U1545 (N_1545,In_737,In_511);
nor U1546 (N_1546,In_658,In_348);
nor U1547 (N_1547,In_564,In_474);
nor U1548 (N_1548,In_297,In_119);
or U1549 (N_1549,In_32,In_285);
nor U1550 (N_1550,In_650,In_363);
xnor U1551 (N_1551,In_706,In_45);
and U1552 (N_1552,In_226,In_667);
xor U1553 (N_1553,In_652,In_220);
nor U1554 (N_1554,In_341,In_524);
xor U1555 (N_1555,In_303,In_386);
nand U1556 (N_1556,In_433,In_457);
xor U1557 (N_1557,In_371,In_283);
and U1558 (N_1558,In_541,In_311);
xor U1559 (N_1559,In_156,In_320);
or U1560 (N_1560,In_537,In_635);
and U1561 (N_1561,In_183,In_591);
xor U1562 (N_1562,In_197,In_490);
and U1563 (N_1563,In_511,In_324);
and U1564 (N_1564,In_690,In_328);
xor U1565 (N_1565,In_107,In_718);
xor U1566 (N_1566,In_675,In_574);
nand U1567 (N_1567,In_182,In_19);
or U1568 (N_1568,In_322,In_693);
xor U1569 (N_1569,In_559,In_380);
nand U1570 (N_1570,In_464,In_613);
or U1571 (N_1571,In_20,In_380);
and U1572 (N_1572,In_677,In_393);
xnor U1573 (N_1573,In_407,In_414);
nor U1574 (N_1574,In_688,In_459);
and U1575 (N_1575,In_255,In_118);
nand U1576 (N_1576,In_82,In_48);
and U1577 (N_1577,In_271,In_506);
and U1578 (N_1578,In_463,In_57);
or U1579 (N_1579,In_570,In_362);
xnor U1580 (N_1580,In_108,In_738);
and U1581 (N_1581,In_532,In_402);
xor U1582 (N_1582,In_403,In_466);
nor U1583 (N_1583,In_573,In_67);
or U1584 (N_1584,In_331,In_553);
and U1585 (N_1585,In_246,In_14);
or U1586 (N_1586,In_175,In_477);
nor U1587 (N_1587,In_499,In_98);
nand U1588 (N_1588,In_2,In_28);
nor U1589 (N_1589,In_240,In_565);
or U1590 (N_1590,In_72,In_460);
and U1591 (N_1591,In_727,In_101);
or U1592 (N_1592,In_46,In_100);
xor U1593 (N_1593,In_657,In_275);
or U1594 (N_1594,In_456,In_77);
or U1595 (N_1595,In_84,In_354);
or U1596 (N_1596,In_667,In_282);
nor U1597 (N_1597,In_277,In_310);
and U1598 (N_1598,In_47,In_644);
xor U1599 (N_1599,In_254,In_377);
and U1600 (N_1600,In_157,In_707);
or U1601 (N_1601,In_8,In_70);
xnor U1602 (N_1602,In_522,In_285);
nor U1603 (N_1603,In_718,In_96);
and U1604 (N_1604,In_251,In_105);
xnor U1605 (N_1605,In_568,In_653);
or U1606 (N_1606,In_318,In_521);
xnor U1607 (N_1607,In_602,In_270);
xor U1608 (N_1608,In_747,In_88);
or U1609 (N_1609,In_283,In_545);
and U1610 (N_1610,In_476,In_685);
xor U1611 (N_1611,In_591,In_132);
and U1612 (N_1612,In_251,In_647);
nor U1613 (N_1613,In_6,In_628);
xor U1614 (N_1614,In_76,In_46);
or U1615 (N_1615,In_635,In_550);
nand U1616 (N_1616,In_614,In_732);
nor U1617 (N_1617,In_206,In_263);
and U1618 (N_1618,In_737,In_391);
xor U1619 (N_1619,In_667,In_422);
or U1620 (N_1620,In_524,In_295);
xor U1621 (N_1621,In_212,In_321);
nor U1622 (N_1622,In_333,In_6);
nor U1623 (N_1623,In_312,In_135);
and U1624 (N_1624,In_27,In_530);
xnor U1625 (N_1625,In_210,In_361);
xnor U1626 (N_1626,In_580,In_210);
or U1627 (N_1627,In_491,In_295);
nor U1628 (N_1628,In_635,In_532);
nor U1629 (N_1629,In_509,In_320);
and U1630 (N_1630,In_151,In_342);
nand U1631 (N_1631,In_441,In_232);
and U1632 (N_1632,In_433,In_297);
or U1633 (N_1633,In_596,In_540);
nor U1634 (N_1634,In_690,In_654);
nand U1635 (N_1635,In_561,In_407);
or U1636 (N_1636,In_145,In_356);
and U1637 (N_1637,In_465,In_662);
and U1638 (N_1638,In_438,In_573);
xor U1639 (N_1639,In_605,In_291);
nand U1640 (N_1640,In_586,In_388);
and U1641 (N_1641,In_319,In_420);
xor U1642 (N_1642,In_318,In_655);
and U1643 (N_1643,In_178,In_295);
and U1644 (N_1644,In_257,In_728);
and U1645 (N_1645,In_406,In_705);
and U1646 (N_1646,In_126,In_471);
nand U1647 (N_1647,In_370,In_385);
nor U1648 (N_1648,In_181,In_195);
and U1649 (N_1649,In_212,In_651);
nand U1650 (N_1650,In_476,In_338);
and U1651 (N_1651,In_160,In_152);
and U1652 (N_1652,In_472,In_208);
and U1653 (N_1653,In_408,In_125);
nor U1654 (N_1654,In_140,In_8);
or U1655 (N_1655,In_748,In_629);
xnor U1656 (N_1656,In_571,In_185);
and U1657 (N_1657,In_397,In_157);
nor U1658 (N_1658,In_738,In_485);
nor U1659 (N_1659,In_633,In_622);
or U1660 (N_1660,In_528,In_321);
and U1661 (N_1661,In_482,In_418);
and U1662 (N_1662,In_584,In_141);
and U1663 (N_1663,In_379,In_503);
xor U1664 (N_1664,In_108,In_242);
and U1665 (N_1665,In_194,In_409);
nor U1666 (N_1666,In_603,In_424);
nor U1667 (N_1667,In_144,In_103);
xnor U1668 (N_1668,In_646,In_469);
and U1669 (N_1669,In_69,In_614);
xor U1670 (N_1670,In_337,In_314);
xor U1671 (N_1671,In_17,In_85);
and U1672 (N_1672,In_124,In_459);
or U1673 (N_1673,In_496,In_249);
and U1674 (N_1674,In_725,In_306);
nor U1675 (N_1675,In_369,In_122);
nand U1676 (N_1676,In_353,In_363);
nor U1677 (N_1677,In_428,In_391);
or U1678 (N_1678,In_252,In_369);
or U1679 (N_1679,In_6,In_433);
nor U1680 (N_1680,In_90,In_628);
xnor U1681 (N_1681,In_221,In_565);
or U1682 (N_1682,In_595,In_728);
and U1683 (N_1683,In_438,In_311);
or U1684 (N_1684,In_599,In_42);
or U1685 (N_1685,In_242,In_737);
nand U1686 (N_1686,In_385,In_313);
nand U1687 (N_1687,In_635,In_614);
nand U1688 (N_1688,In_272,In_680);
xor U1689 (N_1689,In_637,In_45);
nand U1690 (N_1690,In_60,In_558);
nor U1691 (N_1691,In_630,In_139);
or U1692 (N_1692,In_104,In_8);
or U1693 (N_1693,In_82,In_210);
xnor U1694 (N_1694,In_201,In_229);
xor U1695 (N_1695,In_224,In_721);
and U1696 (N_1696,In_122,In_712);
and U1697 (N_1697,In_170,In_231);
nand U1698 (N_1698,In_164,In_311);
xnor U1699 (N_1699,In_652,In_385);
nand U1700 (N_1700,In_357,In_420);
or U1701 (N_1701,In_426,In_127);
xor U1702 (N_1702,In_521,In_115);
or U1703 (N_1703,In_220,In_137);
nand U1704 (N_1704,In_458,In_569);
or U1705 (N_1705,In_424,In_358);
and U1706 (N_1706,In_723,In_298);
or U1707 (N_1707,In_669,In_458);
nor U1708 (N_1708,In_742,In_513);
xor U1709 (N_1709,In_311,In_306);
nor U1710 (N_1710,In_605,In_649);
xnor U1711 (N_1711,In_383,In_721);
and U1712 (N_1712,In_545,In_673);
or U1713 (N_1713,In_542,In_741);
or U1714 (N_1714,In_533,In_426);
nor U1715 (N_1715,In_563,In_242);
nor U1716 (N_1716,In_547,In_493);
or U1717 (N_1717,In_417,In_291);
nand U1718 (N_1718,In_544,In_322);
nand U1719 (N_1719,In_634,In_416);
nor U1720 (N_1720,In_705,In_348);
xnor U1721 (N_1721,In_675,In_367);
nor U1722 (N_1722,In_563,In_428);
nor U1723 (N_1723,In_538,In_562);
nand U1724 (N_1724,In_170,In_508);
or U1725 (N_1725,In_76,In_40);
or U1726 (N_1726,In_347,In_443);
xnor U1727 (N_1727,In_110,In_140);
nand U1728 (N_1728,In_616,In_546);
and U1729 (N_1729,In_726,In_153);
nand U1730 (N_1730,In_72,In_432);
or U1731 (N_1731,In_270,In_597);
xor U1732 (N_1732,In_183,In_586);
nand U1733 (N_1733,In_192,In_87);
nor U1734 (N_1734,In_115,In_603);
xor U1735 (N_1735,In_702,In_191);
or U1736 (N_1736,In_228,In_747);
and U1737 (N_1737,In_523,In_387);
nor U1738 (N_1738,In_691,In_207);
xor U1739 (N_1739,In_599,In_492);
nor U1740 (N_1740,In_247,In_112);
and U1741 (N_1741,In_683,In_392);
or U1742 (N_1742,In_561,In_295);
and U1743 (N_1743,In_102,In_433);
nor U1744 (N_1744,In_427,In_612);
and U1745 (N_1745,In_297,In_447);
xnor U1746 (N_1746,In_582,In_441);
xnor U1747 (N_1747,In_406,In_537);
xor U1748 (N_1748,In_623,In_29);
and U1749 (N_1749,In_352,In_613);
xnor U1750 (N_1750,In_564,In_495);
nor U1751 (N_1751,In_427,In_340);
or U1752 (N_1752,In_103,In_358);
or U1753 (N_1753,In_102,In_692);
or U1754 (N_1754,In_514,In_475);
nand U1755 (N_1755,In_562,In_627);
xnor U1756 (N_1756,In_509,In_237);
nand U1757 (N_1757,In_112,In_639);
xor U1758 (N_1758,In_451,In_36);
and U1759 (N_1759,In_1,In_425);
nor U1760 (N_1760,In_244,In_482);
xnor U1761 (N_1761,In_373,In_362);
xnor U1762 (N_1762,In_93,In_518);
xor U1763 (N_1763,In_639,In_396);
nand U1764 (N_1764,In_395,In_446);
and U1765 (N_1765,In_702,In_15);
nor U1766 (N_1766,In_339,In_72);
or U1767 (N_1767,In_618,In_209);
nor U1768 (N_1768,In_262,In_351);
or U1769 (N_1769,In_608,In_404);
and U1770 (N_1770,In_351,In_578);
xnor U1771 (N_1771,In_253,In_307);
xor U1772 (N_1772,In_544,In_30);
nand U1773 (N_1773,In_468,In_336);
and U1774 (N_1774,In_642,In_27);
nor U1775 (N_1775,In_420,In_299);
and U1776 (N_1776,In_423,In_717);
or U1777 (N_1777,In_419,In_506);
xnor U1778 (N_1778,In_511,In_696);
nand U1779 (N_1779,In_484,In_420);
and U1780 (N_1780,In_97,In_434);
or U1781 (N_1781,In_487,In_462);
xor U1782 (N_1782,In_27,In_327);
or U1783 (N_1783,In_248,In_327);
or U1784 (N_1784,In_133,In_543);
nor U1785 (N_1785,In_537,In_453);
nor U1786 (N_1786,In_272,In_87);
nor U1787 (N_1787,In_374,In_629);
or U1788 (N_1788,In_143,In_274);
or U1789 (N_1789,In_720,In_735);
nand U1790 (N_1790,In_89,In_691);
nor U1791 (N_1791,In_88,In_457);
nand U1792 (N_1792,In_673,In_610);
nor U1793 (N_1793,In_17,In_236);
xnor U1794 (N_1794,In_611,In_121);
and U1795 (N_1795,In_736,In_398);
nor U1796 (N_1796,In_433,In_564);
or U1797 (N_1797,In_196,In_258);
and U1798 (N_1798,In_445,In_78);
or U1799 (N_1799,In_9,In_300);
and U1800 (N_1800,In_726,In_379);
nor U1801 (N_1801,In_613,In_484);
nor U1802 (N_1802,In_263,In_729);
nor U1803 (N_1803,In_647,In_236);
and U1804 (N_1804,In_654,In_447);
nor U1805 (N_1805,In_599,In_279);
and U1806 (N_1806,In_149,In_234);
xor U1807 (N_1807,In_423,In_243);
and U1808 (N_1808,In_263,In_128);
or U1809 (N_1809,In_514,In_637);
nor U1810 (N_1810,In_168,In_541);
nand U1811 (N_1811,In_96,In_28);
or U1812 (N_1812,In_601,In_332);
nor U1813 (N_1813,In_507,In_172);
or U1814 (N_1814,In_523,In_571);
nand U1815 (N_1815,In_138,In_524);
or U1816 (N_1816,In_641,In_111);
nand U1817 (N_1817,In_67,In_561);
or U1818 (N_1818,In_281,In_626);
xor U1819 (N_1819,In_219,In_3);
nor U1820 (N_1820,In_671,In_484);
xnor U1821 (N_1821,In_725,In_588);
xnor U1822 (N_1822,In_195,In_332);
nand U1823 (N_1823,In_203,In_527);
nand U1824 (N_1824,In_513,In_334);
and U1825 (N_1825,In_718,In_409);
nand U1826 (N_1826,In_303,In_166);
and U1827 (N_1827,In_689,In_299);
or U1828 (N_1828,In_215,In_416);
or U1829 (N_1829,In_652,In_384);
xor U1830 (N_1830,In_655,In_441);
nor U1831 (N_1831,In_124,In_696);
xnor U1832 (N_1832,In_235,In_198);
xnor U1833 (N_1833,In_444,In_517);
and U1834 (N_1834,In_185,In_270);
nand U1835 (N_1835,In_89,In_207);
nand U1836 (N_1836,In_108,In_392);
and U1837 (N_1837,In_453,In_493);
nand U1838 (N_1838,In_578,In_468);
and U1839 (N_1839,In_330,In_498);
and U1840 (N_1840,In_385,In_687);
nand U1841 (N_1841,In_740,In_228);
nand U1842 (N_1842,In_461,In_514);
nand U1843 (N_1843,In_247,In_496);
nor U1844 (N_1844,In_713,In_522);
or U1845 (N_1845,In_369,In_4);
nand U1846 (N_1846,In_275,In_472);
or U1847 (N_1847,In_88,In_728);
nor U1848 (N_1848,In_566,In_265);
nand U1849 (N_1849,In_497,In_532);
nand U1850 (N_1850,In_565,In_515);
or U1851 (N_1851,In_630,In_9);
nand U1852 (N_1852,In_27,In_567);
nor U1853 (N_1853,In_552,In_384);
or U1854 (N_1854,In_29,In_277);
xor U1855 (N_1855,In_369,In_91);
xor U1856 (N_1856,In_232,In_470);
nor U1857 (N_1857,In_80,In_156);
nor U1858 (N_1858,In_419,In_634);
xor U1859 (N_1859,In_174,In_218);
nand U1860 (N_1860,In_371,In_275);
and U1861 (N_1861,In_257,In_7);
nand U1862 (N_1862,In_527,In_744);
nor U1863 (N_1863,In_232,In_461);
nor U1864 (N_1864,In_501,In_289);
xnor U1865 (N_1865,In_635,In_427);
and U1866 (N_1866,In_539,In_676);
or U1867 (N_1867,In_165,In_439);
xor U1868 (N_1868,In_578,In_27);
nand U1869 (N_1869,In_352,In_440);
nand U1870 (N_1870,In_191,In_293);
nor U1871 (N_1871,In_653,In_240);
and U1872 (N_1872,In_476,In_403);
xor U1873 (N_1873,In_561,In_165);
xor U1874 (N_1874,In_122,In_116);
nor U1875 (N_1875,In_149,In_148);
nand U1876 (N_1876,In_364,In_56);
or U1877 (N_1877,In_572,In_186);
nand U1878 (N_1878,In_35,In_160);
nor U1879 (N_1879,In_0,In_566);
or U1880 (N_1880,In_693,In_368);
and U1881 (N_1881,In_153,In_514);
nor U1882 (N_1882,In_102,In_86);
and U1883 (N_1883,In_12,In_525);
nor U1884 (N_1884,In_500,In_543);
or U1885 (N_1885,In_165,In_20);
nor U1886 (N_1886,In_594,In_1);
and U1887 (N_1887,In_580,In_109);
nor U1888 (N_1888,In_136,In_486);
or U1889 (N_1889,In_576,In_642);
nor U1890 (N_1890,In_343,In_422);
nand U1891 (N_1891,In_175,In_9);
xnor U1892 (N_1892,In_632,In_74);
xor U1893 (N_1893,In_628,In_0);
or U1894 (N_1894,In_539,In_660);
and U1895 (N_1895,In_150,In_589);
or U1896 (N_1896,In_124,In_743);
and U1897 (N_1897,In_404,In_368);
xnor U1898 (N_1898,In_378,In_420);
or U1899 (N_1899,In_677,In_662);
nor U1900 (N_1900,In_136,In_445);
or U1901 (N_1901,In_683,In_346);
and U1902 (N_1902,In_445,In_391);
xnor U1903 (N_1903,In_731,In_74);
nand U1904 (N_1904,In_425,In_636);
nand U1905 (N_1905,In_301,In_645);
or U1906 (N_1906,In_50,In_188);
xor U1907 (N_1907,In_494,In_153);
xnor U1908 (N_1908,In_353,In_339);
xor U1909 (N_1909,In_250,In_233);
nand U1910 (N_1910,In_427,In_211);
nand U1911 (N_1911,In_52,In_507);
nor U1912 (N_1912,In_195,In_127);
nand U1913 (N_1913,In_432,In_728);
nand U1914 (N_1914,In_24,In_115);
nand U1915 (N_1915,In_282,In_541);
nand U1916 (N_1916,In_725,In_616);
nor U1917 (N_1917,In_307,In_35);
nand U1918 (N_1918,In_311,In_123);
or U1919 (N_1919,In_454,In_738);
nand U1920 (N_1920,In_538,In_213);
nand U1921 (N_1921,In_527,In_205);
xor U1922 (N_1922,In_665,In_306);
or U1923 (N_1923,In_300,In_646);
nand U1924 (N_1924,In_535,In_312);
and U1925 (N_1925,In_138,In_476);
nand U1926 (N_1926,In_404,In_398);
nand U1927 (N_1927,In_336,In_109);
nor U1928 (N_1928,In_526,In_485);
nand U1929 (N_1929,In_366,In_211);
and U1930 (N_1930,In_392,In_559);
nand U1931 (N_1931,In_244,In_372);
nor U1932 (N_1932,In_17,In_740);
nor U1933 (N_1933,In_505,In_359);
nand U1934 (N_1934,In_75,In_460);
and U1935 (N_1935,In_518,In_229);
xnor U1936 (N_1936,In_654,In_34);
nand U1937 (N_1937,In_15,In_346);
or U1938 (N_1938,In_389,In_41);
nor U1939 (N_1939,In_134,In_556);
or U1940 (N_1940,In_593,In_479);
and U1941 (N_1941,In_268,In_222);
nor U1942 (N_1942,In_497,In_707);
nand U1943 (N_1943,In_607,In_344);
nand U1944 (N_1944,In_47,In_700);
nor U1945 (N_1945,In_610,In_481);
nand U1946 (N_1946,In_87,In_33);
nor U1947 (N_1947,In_339,In_507);
nand U1948 (N_1948,In_467,In_116);
nor U1949 (N_1949,In_76,In_16);
or U1950 (N_1950,In_301,In_673);
nor U1951 (N_1951,In_541,In_130);
or U1952 (N_1952,In_601,In_65);
and U1953 (N_1953,In_207,In_329);
or U1954 (N_1954,In_430,In_6);
nor U1955 (N_1955,In_51,In_177);
or U1956 (N_1956,In_583,In_64);
and U1957 (N_1957,In_426,In_558);
and U1958 (N_1958,In_741,In_185);
nor U1959 (N_1959,In_222,In_438);
xor U1960 (N_1960,In_605,In_311);
nand U1961 (N_1961,In_102,In_744);
xor U1962 (N_1962,In_312,In_497);
and U1963 (N_1963,In_347,In_591);
nand U1964 (N_1964,In_534,In_150);
xor U1965 (N_1965,In_381,In_223);
or U1966 (N_1966,In_144,In_93);
and U1967 (N_1967,In_476,In_711);
xor U1968 (N_1968,In_314,In_27);
nor U1969 (N_1969,In_629,In_505);
xnor U1970 (N_1970,In_712,In_219);
or U1971 (N_1971,In_145,In_300);
xor U1972 (N_1972,In_249,In_369);
nor U1973 (N_1973,In_172,In_228);
nor U1974 (N_1974,In_511,In_568);
or U1975 (N_1975,In_594,In_687);
and U1976 (N_1976,In_362,In_180);
nand U1977 (N_1977,In_95,In_682);
nor U1978 (N_1978,In_540,In_413);
xor U1979 (N_1979,In_503,In_40);
and U1980 (N_1980,In_271,In_306);
xnor U1981 (N_1981,In_512,In_105);
and U1982 (N_1982,In_97,In_159);
nor U1983 (N_1983,In_137,In_718);
or U1984 (N_1984,In_705,In_100);
nor U1985 (N_1985,In_710,In_417);
or U1986 (N_1986,In_225,In_660);
xor U1987 (N_1987,In_57,In_611);
and U1988 (N_1988,In_12,In_162);
nor U1989 (N_1989,In_668,In_365);
or U1990 (N_1990,In_50,In_320);
and U1991 (N_1991,In_156,In_327);
nand U1992 (N_1992,In_345,In_458);
and U1993 (N_1993,In_205,In_712);
nand U1994 (N_1994,In_552,In_666);
nor U1995 (N_1995,In_691,In_224);
xor U1996 (N_1996,In_156,In_203);
nand U1997 (N_1997,In_533,In_537);
or U1998 (N_1998,In_288,In_496);
and U1999 (N_1999,In_200,In_569);
or U2000 (N_2000,In_389,In_625);
nor U2001 (N_2001,In_749,In_649);
nand U2002 (N_2002,In_423,In_556);
nand U2003 (N_2003,In_494,In_521);
or U2004 (N_2004,In_406,In_274);
xor U2005 (N_2005,In_585,In_670);
nor U2006 (N_2006,In_701,In_596);
nor U2007 (N_2007,In_68,In_16);
xor U2008 (N_2008,In_541,In_453);
nor U2009 (N_2009,In_240,In_5);
nand U2010 (N_2010,In_556,In_720);
xnor U2011 (N_2011,In_639,In_602);
or U2012 (N_2012,In_245,In_138);
or U2013 (N_2013,In_404,In_498);
nor U2014 (N_2014,In_351,In_292);
xor U2015 (N_2015,In_355,In_598);
and U2016 (N_2016,In_337,In_133);
xnor U2017 (N_2017,In_482,In_383);
xor U2018 (N_2018,In_677,In_131);
nand U2019 (N_2019,In_645,In_272);
nand U2020 (N_2020,In_349,In_270);
nand U2021 (N_2021,In_526,In_359);
or U2022 (N_2022,In_183,In_317);
nor U2023 (N_2023,In_253,In_151);
or U2024 (N_2024,In_136,In_731);
xnor U2025 (N_2025,In_474,In_61);
or U2026 (N_2026,In_621,In_672);
and U2027 (N_2027,In_502,In_249);
nor U2028 (N_2028,In_414,In_392);
or U2029 (N_2029,In_553,In_54);
and U2030 (N_2030,In_593,In_270);
xor U2031 (N_2031,In_582,In_428);
xnor U2032 (N_2032,In_349,In_372);
xor U2033 (N_2033,In_254,In_242);
or U2034 (N_2034,In_66,In_274);
or U2035 (N_2035,In_672,In_533);
nor U2036 (N_2036,In_645,In_136);
nor U2037 (N_2037,In_626,In_275);
nand U2038 (N_2038,In_241,In_631);
or U2039 (N_2039,In_164,In_706);
nor U2040 (N_2040,In_447,In_539);
nor U2041 (N_2041,In_515,In_388);
xor U2042 (N_2042,In_421,In_595);
xnor U2043 (N_2043,In_17,In_509);
or U2044 (N_2044,In_256,In_258);
or U2045 (N_2045,In_588,In_249);
xnor U2046 (N_2046,In_83,In_257);
and U2047 (N_2047,In_326,In_22);
nand U2048 (N_2048,In_302,In_96);
or U2049 (N_2049,In_80,In_711);
xnor U2050 (N_2050,In_327,In_729);
or U2051 (N_2051,In_469,In_471);
nor U2052 (N_2052,In_364,In_663);
or U2053 (N_2053,In_90,In_170);
or U2054 (N_2054,In_419,In_74);
xor U2055 (N_2055,In_398,In_479);
nor U2056 (N_2056,In_630,In_144);
nand U2057 (N_2057,In_633,In_730);
or U2058 (N_2058,In_488,In_37);
nor U2059 (N_2059,In_270,In_376);
or U2060 (N_2060,In_59,In_465);
nor U2061 (N_2061,In_655,In_219);
xnor U2062 (N_2062,In_407,In_628);
nand U2063 (N_2063,In_244,In_544);
xnor U2064 (N_2064,In_253,In_241);
xor U2065 (N_2065,In_447,In_274);
and U2066 (N_2066,In_162,In_712);
nand U2067 (N_2067,In_688,In_187);
nor U2068 (N_2068,In_496,In_283);
or U2069 (N_2069,In_630,In_39);
nor U2070 (N_2070,In_235,In_299);
or U2071 (N_2071,In_374,In_513);
or U2072 (N_2072,In_595,In_59);
nand U2073 (N_2073,In_180,In_508);
nand U2074 (N_2074,In_635,In_286);
xnor U2075 (N_2075,In_412,In_582);
nand U2076 (N_2076,In_481,In_32);
and U2077 (N_2077,In_736,In_173);
and U2078 (N_2078,In_749,In_182);
or U2079 (N_2079,In_157,In_512);
and U2080 (N_2080,In_464,In_584);
nand U2081 (N_2081,In_586,In_595);
nor U2082 (N_2082,In_74,In_231);
or U2083 (N_2083,In_603,In_691);
nor U2084 (N_2084,In_392,In_312);
xnor U2085 (N_2085,In_744,In_516);
and U2086 (N_2086,In_114,In_496);
nand U2087 (N_2087,In_388,In_8);
or U2088 (N_2088,In_89,In_16);
nand U2089 (N_2089,In_587,In_666);
or U2090 (N_2090,In_55,In_715);
nand U2091 (N_2091,In_253,In_575);
nor U2092 (N_2092,In_85,In_266);
xnor U2093 (N_2093,In_56,In_678);
and U2094 (N_2094,In_473,In_248);
xor U2095 (N_2095,In_98,In_569);
or U2096 (N_2096,In_564,In_477);
or U2097 (N_2097,In_222,In_367);
or U2098 (N_2098,In_127,In_261);
or U2099 (N_2099,In_642,In_505);
or U2100 (N_2100,In_160,In_512);
nor U2101 (N_2101,In_374,In_151);
xor U2102 (N_2102,In_221,In_643);
nor U2103 (N_2103,In_349,In_563);
or U2104 (N_2104,In_188,In_747);
xor U2105 (N_2105,In_379,In_223);
nor U2106 (N_2106,In_383,In_648);
nand U2107 (N_2107,In_359,In_239);
xnor U2108 (N_2108,In_307,In_164);
nor U2109 (N_2109,In_501,In_278);
nor U2110 (N_2110,In_159,In_166);
or U2111 (N_2111,In_336,In_669);
or U2112 (N_2112,In_552,In_408);
and U2113 (N_2113,In_616,In_129);
xor U2114 (N_2114,In_48,In_143);
and U2115 (N_2115,In_59,In_420);
nand U2116 (N_2116,In_408,In_255);
nand U2117 (N_2117,In_350,In_377);
nor U2118 (N_2118,In_638,In_78);
nor U2119 (N_2119,In_107,In_747);
nand U2120 (N_2120,In_284,In_511);
nor U2121 (N_2121,In_54,In_186);
or U2122 (N_2122,In_498,In_414);
nand U2123 (N_2123,In_16,In_133);
nand U2124 (N_2124,In_198,In_449);
nor U2125 (N_2125,In_572,In_95);
nand U2126 (N_2126,In_669,In_151);
and U2127 (N_2127,In_476,In_688);
nor U2128 (N_2128,In_40,In_337);
xnor U2129 (N_2129,In_449,In_584);
or U2130 (N_2130,In_182,In_682);
nand U2131 (N_2131,In_409,In_568);
or U2132 (N_2132,In_172,In_311);
nor U2133 (N_2133,In_88,In_179);
and U2134 (N_2134,In_367,In_227);
nor U2135 (N_2135,In_134,In_255);
or U2136 (N_2136,In_2,In_214);
or U2137 (N_2137,In_305,In_285);
nand U2138 (N_2138,In_454,In_468);
or U2139 (N_2139,In_152,In_665);
and U2140 (N_2140,In_200,In_407);
xnor U2141 (N_2141,In_224,In_487);
and U2142 (N_2142,In_195,In_388);
nor U2143 (N_2143,In_445,In_507);
or U2144 (N_2144,In_56,In_642);
nand U2145 (N_2145,In_169,In_588);
xnor U2146 (N_2146,In_217,In_592);
and U2147 (N_2147,In_25,In_604);
nand U2148 (N_2148,In_199,In_37);
nand U2149 (N_2149,In_83,In_178);
nand U2150 (N_2150,In_46,In_580);
nand U2151 (N_2151,In_421,In_139);
or U2152 (N_2152,In_611,In_122);
nand U2153 (N_2153,In_569,In_476);
xor U2154 (N_2154,In_743,In_248);
nor U2155 (N_2155,In_209,In_464);
and U2156 (N_2156,In_654,In_29);
xor U2157 (N_2157,In_293,In_689);
xnor U2158 (N_2158,In_25,In_649);
nand U2159 (N_2159,In_546,In_653);
or U2160 (N_2160,In_126,In_517);
and U2161 (N_2161,In_17,In_13);
xnor U2162 (N_2162,In_724,In_640);
xnor U2163 (N_2163,In_538,In_164);
or U2164 (N_2164,In_33,In_599);
and U2165 (N_2165,In_68,In_433);
and U2166 (N_2166,In_150,In_630);
nor U2167 (N_2167,In_627,In_102);
nor U2168 (N_2168,In_6,In_62);
xnor U2169 (N_2169,In_602,In_50);
nor U2170 (N_2170,In_267,In_670);
nor U2171 (N_2171,In_423,In_171);
xor U2172 (N_2172,In_193,In_657);
or U2173 (N_2173,In_2,In_548);
nor U2174 (N_2174,In_480,In_238);
nand U2175 (N_2175,In_482,In_330);
and U2176 (N_2176,In_95,In_481);
nand U2177 (N_2177,In_563,In_40);
nand U2178 (N_2178,In_670,In_452);
or U2179 (N_2179,In_459,In_705);
nand U2180 (N_2180,In_646,In_327);
xor U2181 (N_2181,In_650,In_70);
and U2182 (N_2182,In_705,In_394);
xnor U2183 (N_2183,In_61,In_501);
nand U2184 (N_2184,In_279,In_522);
or U2185 (N_2185,In_477,In_651);
xor U2186 (N_2186,In_631,In_444);
nor U2187 (N_2187,In_252,In_307);
nor U2188 (N_2188,In_191,In_603);
nand U2189 (N_2189,In_166,In_134);
and U2190 (N_2190,In_521,In_638);
or U2191 (N_2191,In_427,In_471);
nor U2192 (N_2192,In_152,In_362);
nand U2193 (N_2193,In_400,In_515);
nand U2194 (N_2194,In_361,In_641);
or U2195 (N_2195,In_24,In_159);
xor U2196 (N_2196,In_71,In_333);
xor U2197 (N_2197,In_703,In_592);
or U2198 (N_2198,In_672,In_554);
and U2199 (N_2199,In_599,In_747);
or U2200 (N_2200,In_474,In_68);
and U2201 (N_2201,In_430,In_700);
and U2202 (N_2202,In_84,In_26);
and U2203 (N_2203,In_130,In_718);
nand U2204 (N_2204,In_500,In_700);
xnor U2205 (N_2205,In_267,In_563);
nor U2206 (N_2206,In_72,In_685);
xnor U2207 (N_2207,In_207,In_366);
nand U2208 (N_2208,In_167,In_604);
nand U2209 (N_2209,In_171,In_476);
nor U2210 (N_2210,In_259,In_641);
or U2211 (N_2211,In_61,In_48);
and U2212 (N_2212,In_518,In_364);
or U2213 (N_2213,In_144,In_664);
nor U2214 (N_2214,In_613,In_688);
xnor U2215 (N_2215,In_460,In_749);
nand U2216 (N_2216,In_337,In_341);
or U2217 (N_2217,In_139,In_278);
xor U2218 (N_2218,In_536,In_504);
nor U2219 (N_2219,In_106,In_423);
and U2220 (N_2220,In_615,In_738);
nand U2221 (N_2221,In_288,In_598);
and U2222 (N_2222,In_259,In_410);
or U2223 (N_2223,In_633,In_477);
and U2224 (N_2224,In_16,In_403);
nor U2225 (N_2225,In_155,In_407);
and U2226 (N_2226,In_249,In_435);
nor U2227 (N_2227,In_115,In_448);
nor U2228 (N_2228,In_542,In_187);
nor U2229 (N_2229,In_168,In_110);
or U2230 (N_2230,In_278,In_328);
xnor U2231 (N_2231,In_243,In_102);
xor U2232 (N_2232,In_561,In_58);
nand U2233 (N_2233,In_269,In_105);
and U2234 (N_2234,In_243,In_327);
nand U2235 (N_2235,In_237,In_285);
or U2236 (N_2236,In_168,In_383);
xor U2237 (N_2237,In_541,In_526);
nand U2238 (N_2238,In_68,In_418);
nor U2239 (N_2239,In_180,In_120);
nand U2240 (N_2240,In_18,In_583);
nor U2241 (N_2241,In_667,In_633);
and U2242 (N_2242,In_155,In_455);
nor U2243 (N_2243,In_461,In_742);
xor U2244 (N_2244,In_237,In_321);
nor U2245 (N_2245,In_330,In_510);
or U2246 (N_2246,In_134,In_473);
xor U2247 (N_2247,In_308,In_502);
nand U2248 (N_2248,In_736,In_159);
or U2249 (N_2249,In_576,In_653);
nor U2250 (N_2250,In_657,In_263);
nor U2251 (N_2251,In_129,In_744);
nor U2252 (N_2252,In_196,In_141);
and U2253 (N_2253,In_72,In_466);
or U2254 (N_2254,In_241,In_498);
and U2255 (N_2255,In_725,In_648);
xor U2256 (N_2256,In_382,In_352);
or U2257 (N_2257,In_171,In_571);
nor U2258 (N_2258,In_99,In_195);
xnor U2259 (N_2259,In_66,In_148);
nor U2260 (N_2260,In_363,In_138);
nand U2261 (N_2261,In_676,In_460);
nor U2262 (N_2262,In_455,In_16);
xnor U2263 (N_2263,In_118,In_682);
nand U2264 (N_2264,In_710,In_717);
or U2265 (N_2265,In_232,In_155);
and U2266 (N_2266,In_171,In_666);
or U2267 (N_2267,In_154,In_580);
nand U2268 (N_2268,In_498,In_451);
or U2269 (N_2269,In_382,In_457);
nor U2270 (N_2270,In_7,In_599);
or U2271 (N_2271,In_319,In_198);
xnor U2272 (N_2272,In_683,In_134);
nor U2273 (N_2273,In_43,In_653);
nand U2274 (N_2274,In_267,In_543);
or U2275 (N_2275,In_463,In_529);
xor U2276 (N_2276,In_314,In_180);
nor U2277 (N_2277,In_16,In_603);
nor U2278 (N_2278,In_277,In_42);
nand U2279 (N_2279,In_541,In_331);
nand U2280 (N_2280,In_719,In_64);
or U2281 (N_2281,In_73,In_656);
xnor U2282 (N_2282,In_93,In_369);
nor U2283 (N_2283,In_600,In_497);
and U2284 (N_2284,In_680,In_587);
nor U2285 (N_2285,In_588,In_351);
nor U2286 (N_2286,In_112,In_432);
and U2287 (N_2287,In_552,In_584);
nor U2288 (N_2288,In_10,In_142);
nand U2289 (N_2289,In_549,In_474);
nor U2290 (N_2290,In_385,In_634);
nor U2291 (N_2291,In_525,In_146);
nand U2292 (N_2292,In_317,In_245);
nor U2293 (N_2293,In_29,In_71);
xnor U2294 (N_2294,In_277,In_218);
nand U2295 (N_2295,In_201,In_159);
nand U2296 (N_2296,In_531,In_719);
nand U2297 (N_2297,In_363,In_559);
xor U2298 (N_2298,In_570,In_444);
or U2299 (N_2299,In_282,In_85);
nor U2300 (N_2300,In_397,In_598);
xor U2301 (N_2301,In_689,In_684);
nor U2302 (N_2302,In_203,In_512);
nand U2303 (N_2303,In_546,In_161);
nor U2304 (N_2304,In_62,In_400);
nor U2305 (N_2305,In_616,In_141);
xnor U2306 (N_2306,In_400,In_433);
nand U2307 (N_2307,In_77,In_110);
nand U2308 (N_2308,In_570,In_207);
nor U2309 (N_2309,In_462,In_4);
and U2310 (N_2310,In_622,In_567);
or U2311 (N_2311,In_680,In_184);
nor U2312 (N_2312,In_510,In_718);
and U2313 (N_2313,In_507,In_658);
and U2314 (N_2314,In_543,In_227);
nor U2315 (N_2315,In_15,In_319);
nor U2316 (N_2316,In_408,In_470);
xnor U2317 (N_2317,In_739,In_292);
xnor U2318 (N_2318,In_611,In_549);
or U2319 (N_2319,In_49,In_387);
xnor U2320 (N_2320,In_240,In_341);
xor U2321 (N_2321,In_493,In_477);
xnor U2322 (N_2322,In_466,In_171);
and U2323 (N_2323,In_339,In_578);
and U2324 (N_2324,In_413,In_325);
or U2325 (N_2325,In_96,In_482);
nand U2326 (N_2326,In_440,In_410);
nand U2327 (N_2327,In_453,In_504);
xnor U2328 (N_2328,In_578,In_251);
nand U2329 (N_2329,In_582,In_629);
nor U2330 (N_2330,In_197,In_254);
or U2331 (N_2331,In_269,In_219);
xor U2332 (N_2332,In_294,In_23);
or U2333 (N_2333,In_688,In_275);
and U2334 (N_2334,In_631,In_255);
xnor U2335 (N_2335,In_326,In_727);
xor U2336 (N_2336,In_711,In_604);
xor U2337 (N_2337,In_494,In_459);
xor U2338 (N_2338,In_486,In_641);
xor U2339 (N_2339,In_573,In_151);
and U2340 (N_2340,In_607,In_64);
nand U2341 (N_2341,In_370,In_413);
xnor U2342 (N_2342,In_130,In_435);
nor U2343 (N_2343,In_278,In_354);
nor U2344 (N_2344,In_248,In_612);
xor U2345 (N_2345,In_232,In_636);
or U2346 (N_2346,In_212,In_230);
nor U2347 (N_2347,In_191,In_275);
and U2348 (N_2348,In_735,In_245);
nor U2349 (N_2349,In_483,In_318);
nor U2350 (N_2350,In_50,In_303);
nand U2351 (N_2351,In_720,In_29);
or U2352 (N_2352,In_666,In_339);
nand U2353 (N_2353,In_346,In_338);
and U2354 (N_2354,In_106,In_718);
nand U2355 (N_2355,In_366,In_697);
and U2356 (N_2356,In_26,In_583);
nor U2357 (N_2357,In_363,In_83);
nand U2358 (N_2358,In_659,In_722);
nor U2359 (N_2359,In_708,In_516);
xnor U2360 (N_2360,In_192,In_52);
xnor U2361 (N_2361,In_414,In_317);
xor U2362 (N_2362,In_21,In_563);
xor U2363 (N_2363,In_120,In_128);
or U2364 (N_2364,In_94,In_272);
and U2365 (N_2365,In_472,In_482);
and U2366 (N_2366,In_72,In_239);
nor U2367 (N_2367,In_429,In_539);
or U2368 (N_2368,In_376,In_501);
nor U2369 (N_2369,In_53,In_559);
nor U2370 (N_2370,In_241,In_464);
and U2371 (N_2371,In_215,In_548);
or U2372 (N_2372,In_312,In_501);
xor U2373 (N_2373,In_269,In_436);
nand U2374 (N_2374,In_157,In_196);
xor U2375 (N_2375,In_459,In_588);
nand U2376 (N_2376,In_389,In_287);
xnor U2377 (N_2377,In_743,In_688);
nand U2378 (N_2378,In_23,In_60);
nor U2379 (N_2379,In_474,In_590);
nand U2380 (N_2380,In_447,In_598);
and U2381 (N_2381,In_143,In_577);
nor U2382 (N_2382,In_272,In_240);
nand U2383 (N_2383,In_739,In_73);
nand U2384 (N_2384,In_358,In_427);
or U2385 (N_2385,In_518,In_194);
nand U2386 (N_2386,In_49,In_79);
nand U2387 (N_2387,In_111,In_359);
nand U2388 (N_2388,In_235,In_462);
nand U2389 (N_2389,In_359,In_738);
or U2390 (N_2390,In_566,In_24);
and U2391 (N_2391,In_480,In_440);
and U2392 (N_2392,In_252,In_385);
or U2393 (N_2393,In_420,In_348);
and U2394 (N_2394,In_628,In_491);
xor U2395 (N_2395,In_232,In_707);
nand U2396 (N_2396,In_25,In_59);
xor U2397 (N_2397,In_260,In_384);
or U2398 (N_2398,In_509,In_234);
or U2399 (N_2399,In_609,In_367);
nor U2400 (N_2400,In_434,In_416);
nand U2401 (N_2401,In_225,In_81);
and U2402 (N_2402,In_681,In_271);
nand U2403 (N_2403,In_268,In_697);
xnor U2404 (N_2404,In_709,In_595);
or U2405 (N_2405,In_475,In_156);
and U2406 (N_2406,In_671,In_568);
xor U2407 (N_2407,In_504,In_514);
nand U2408 (N_2408,In_133,In_396);
nand U2409 (N_2409,In_405,In_607);
and U2410 (N_2410,In_699,In_593);
and U2411 (N_2411,In_602,In_633);
nand U2412 (N_2412,In_240,In_34);
nand U2413 (N_2413,In_642,In_174);
xnor U2414 (N_2414,In_200,In_182);
and U2415 (N_2415,In_414,In_157);
and U2416 (N_2416,In_178,In_483);
or U2417 (N_2417,In_203,In_75);
nor U2418 (N_2418,In_397,In_620);
or U2419 (N_2419,In_408,In_488);
or U2420 (N_2420,In_117,In_52);
nor U2421 (N_2421,In_325,In_582);
and U2422 (N_2422,In_407,In_430);
xor U2423 (N_2423,In_105,In_529);
or U2424 (N_2424,In_94,In_530);
and U2425 (N_2425,In_85,In_445);
and U2426 (N_2426,In_425,In_148);
xnor U2427 (N_2427,In_701,In_263);
xnor U2428 (N_2428,In_179,In_651);
nand U2429 (N_2429,In_530,In_747);
xnor U2430 (N_2430,In_657,In_426);
nor U2431 (N_2431,In_67,In_605);
or U2432 (N_2432,In_73,In_692);
or U2433 (N_2433,In_356,In_91);
and U2434 (N_2434,In_494,In_622);
and U2435 (N_2435,In_9,In_320);
nand U2436 (N_2436,In_508,In_302);
or U2437 (N_2437,In_276,In_726);
xor U2438 (N_2438,In_119,In_29);
xnor U2439 (N_2439,In_531,In_291);
xor U2440 (N_2440,In_521,In_75);
nand U2441 (N_2441,In_540,In_19);
or U2442 (N_2442,In_61,In_411);
and U2443 (N_2443,In_694,In_216);
or U2444 (N_2444,In_231,In_166);
xor U2445 (N_2445,In_390,In_552);
nand U2446 (N_2446,In_358,In_716);
nand U2447 (N_2447,In_382,In_357);
or U2448 (N_2448,In_636,In_422);
nor U2449 (N_2449,In_710,In_591);
and U2450 (N_2450,In_197,In_359);
or U2451 (N_2451,In_361,In_218);
and U2452 (N_2452,In_115,In_367);
or U2453 (N_2453,In_345,In_225);
or U2454 (N_2454,In_617,In_63);
nor U2455 (N_2455,In_506,In_437);
and U2456 (N_2456,In_605,In_78);
nand U2457 (N_2457,In_560,In_415);
or U2458 (N_2458,In_207,In_644);
and U2459 (N_2459,In_458,In_682);
xnor U2460 (N_2460,In_622,In_524);
and U2461 (N_2461,In_213,In_677);
or U2462 (N_2462,In_295,In_201);
or U2463 (N_2463,In_702,In_32);
nand U2464 (N_2464,In_464,In_731);
xnor U2465 (N_2465,In_615,In_468);
and U2466 (N_2466,In_439,In_593);
nand U2467 (N_2467,In_566,In_86);
xor U2468 (N_2468,In_686,In_254);
and U2469 (N_2469,In_638,In_305);
nor U2470 (N_2470,In_379,In_397);
nand U2471 (N_2471,In_499,In_636);
nand U2472 (N_2472,In_540,In_118);
xnor U2473 (N_2473,In_674,In_86);
nor U2474 (N_2474,In_363,In_58);
nand U2475 (N_2475,In_529,In_663);
nand U2476 (N_2476,In_92,In_573);
xnor U2477 (N_2477,In_112,In_401);
or U2478 (N_2478,In_740,In_512);
xor U2479 (N_2479,In_9,In_476);
and U2480 (N_2480,In_552,In_704);
or U2481 (N_2481,In_674,In_535);
nand U2482 (N_2482,In_445,In_115);
nand U2483 (N_2483,In_190,In_716);
xor U2484 (N_2484,In_278,In_214);
nor U2485 (N_2485,In_632,In_287);
or U2486 (N_2486,In_186,In_635);
nand U2487 (N_2487,In_339,In_319);
nand U2488 (N_2488,In_653,In_668);
and U2489 (N_2489,In_197,In_652);
nor U2490 (N_2490,In_615,In_192);
nor U2491 (N_2491,In_373,In_622);
or U2492 (N_2492,In_434,In_600);
and U2493 (N_2493,In_170,In_98);
xnor U2494 (N_2494,In_724,In_257);
nor U2495 (N_2495,In_435,In_5);
or U2496 (N_2496,In_485,In_299);
xor U2497 (N_2497,In_585,In_738);
or U2498 (N_2498,In_708,In_699);
nand U2499 (N_2499,In_424,In_488);
nor U2500 (N_2500,N_2047,N_446);
nand U2501 (N_2501,N_1497,N_2350);
and U2502 (N_2502,N_321,N_1926);
or U2503 (N_2503,N_449,N_137);
nand U2504 (N_2504,N_2346,N_2131);
nor U2505 (N_2505,N_2101,N_1632);
xnor U2506 (N_2506,N_1611,N_1571);
and U2507 (N_2507,N_2467,N_582);
xor U2508 (N_2508,N_2174,N_2414);
nor U2509 (N_2509,N_564,N_1620);
nor U2510 (N_2510,N_574,N_2291);
or U2511 (N_2511,N_103,N_828);
and U2512 (N_2512,N_2354,N_1508);
xor U2513 (N_2513,N_1826,N_2442);
and U2514 (N_2514,N_1799,N_1474);
nand U2515 (N_2515,N_1405,N_577);
or U2516 (N_2516,N_2033,N_36);
nor U2517 (N_2517,N_1201,N_1433);
nor U2518 (N_2518,N_1931,N_1911);
and U2519 (N_2519,N_28,N_482);
xor U2520 (N_2520,N_204,N_179);
and U2521 (N_2521,N_1297,N_300);
nand U2522 (N_2522,N_2483,N_1473);
or U2523 (N_2523,N_1424,N_205);
xor U2524 (N_2524,N_1537,N_202);
nand U2525 (N_2525,N_1205,N_1998);
and U2526 (N_2526,N_2477,N_73);
and U2527 (N_2527,N_241,N_1524);
nand U2528 (N_2528,N_1130,N_2024);
or U2529 (N_2529,N_1533,N_1888);
or U2530 (N_2530,N_2040,N_1189);
xnor U2531 (N_2531,N_439,N_2066);
and U2532 (N_2532,N_2378,N_2320);
or U2533 (N_2533,N_2492,N_2085);
xnor U2534 (N_2534,N_166,N_399);
nand U2535 (N_2535,N_1725,N_2470);
nor U2536 (N_2536,N_852,N_1574);
xor U2537 (N_2537,N_401,N_333);
nor U2538 (N_2538,N_55,N_1085);
xnor U2539 (N_2539,N_939,N_1621);
or U2540 (N_2540,N_1939,N_432);
xor U2541 (N_2541,N_1949,N_301);
nor U2542 (N_2542,N_686,N_1882);
nor U2543 (N_2543,N_102,N_614);
xor U2544 (N_2544,N_834,N_724);
nor U2545 (N_2545,N_2261,N_1715);
nand U2546 (N_2546,N_1785,N_1486);
xor U2547 (N_2547,N_912,N_226);
xor U2548 (N_2548,N_1338,N_1285);
nand U2549 (N_2549,N_810,N_1220);
and U2550 (N_2550,N_525,N_1208);
xnor U2551 (N_2551,N_144,N_1019);
nor U2552 (N_2552,N_452,N_1359);
and U2553 (N_2553,N_1634,N_1562);
or U2554 (N_2554,N_502,N_111);
and U2555 (N_2555,N_1090,N_2459);
and U2556 (N_2556,N_937,N_917);
or U2557 (N_2557,N_1616,N_1464);
and U2558 (N_2558,N_1197,N_892);
nand U2559 (N_2559,N_200,N_165);
nand U2560 (N_2560,N_1141,N_113);
xnor U2561 (N_2561,N_1292,N_485);
nor U2562 (N_2562,N_781,N_1552);
or U2563 (N_2563,N_745,N_1892);
nand U2564 (N_2564,N_1328,N_2155);
xor U2565 (N_2565,N_1767,N_907);
nand U2566 (N_2566,N_1116,N_1749);
or U2567 (N_2567,N_1569,N_529);
xor U2568 (N_2568,N_651,N_732);
or U2569 (N_2569,N_1315,N_2218);
xnor U2570 (N_2570,N_1195,N_1123);
and U2571 (N_2571,N_1327,N_2349);
nor U2572 (N_2572,N_2400,N_203);
nor U2573 (N_2573,N_1352,N_1403);
nor U2574 (N_2574,N_1243,N_623);
or U2575 (N_2575,N_801,N_265);
nand U2576 (N_2576,N_1301,N_63);
xor U2577 (N_2577,N_1042,N_692);
nand U2578 (N_2578,N_1371,N_1385);
nand U2579 (N_2579,N_34,N_1692);
nand U2580 (N_2580,N_1717,N_1002);
nand U2581 (N_2581,N_2173,N_2123);
xnor U2582 (N_2582,N_2335,N_326);
or U2583 (N_2583,N_469,N_1505);
nor U2584 (N_2584,N_555,N_1481);
nor U2585 (N_2585,N_1412,N_2021);
or U2586 (N_2586,N_531,N_1860);
and U2587 (N_2587,N_327,N_925);
or U2588 (N_2588,N_1649,N_2413);
and U2589 (N_2589,N_899,N_2267);
xnor U2590 (N_2590,N_415,N_296);
nor U2591 (N_2591,N_2433,N_2284);
xor U2592 (N_2592,N_764,N_713);
nand U2593 (N_2593,N_1365,N_1993);
xnor U2594 (N_2594,N_230,N_51);
nor U2595 (N_2595,N_2468,N_1868);
nand U2596 (N_2596,N_1284,N_1314);
or U2597 (N_2597,N_1770,N_1542);
nor U2598 (N_2598,N_381,N_1659);
nor U2599 (N_2599,N_755,N_2336);
nand U2600 (N_2600,N_1759,N_1748);
or U2601 (N_2601,N_1335,N_1206);
xnor U2602 (N_2602,N_107,N_257);
xnor U2603 (N_2603,N_1721,N_1483);
xor U2604 (N_2604,N_1633,N_843);
xnor U2605 (N_2605,N_1999,N_1408);
nor U2606 (N_2606,N_2077,N_1270);
or U2607 (N_2607,N_526,N_1738);
and U2608 (N_2608,N_661,N_1257);
or U2609 (N_2609,N_122,N_1758);
nor U2610 (N_2610,N_978,N_1752);
nand U2611 (N_2611,N_58,N_911);
xor U2612 (N_2612,N_310,N_313);
xnor U2613 (N_2613,N_2403,N_1191);
or U2614 (N_2614,N_920,N_94);
xnor U2615 (N_2615,N_2427,N_2264);
or U2616 (N_2616,N_2089,N_1991);
nor U2617 (N_2617,N_1641,N_342);
nor U2618 (N_2618,N_1716,N_2493);
xnor U2619 (N_2619,N_998,N_80);
xor U2620 (N_2620,N_463,N_735);
xor U2621 (N_2621,N_744,N_2053);
xnor U2622 (N_2622,N_2387,N_1112);
nand U2623 (N_2623,N_1094,N_220);
nor U2624 (N_2624,N_969,N_2120);
nor U2625 (N_2625,N_2306,N_2265);
and U2626 (N_2626,N_2460,N_979);
xor U2627 (N_2627,N_626,N_2049);
and U2628 (N_2628,N_2048,N_2154);
nor U2629 (N_2629,N_796,N_856);
xor U2630 (N_2630,N_1828,N_2418);
and U2631 (N_2631,N_1095,N_832);
nand U2632 (N_2632,N_649,N_2344);
nor U2633 (N_2633,N_1955,N_1531);
and U2634 (N_2634,N_1513,N_219);
or U2635 (N_2635,N_589,N_1591);
xor U2636 (N_2636,N_2422,N_1152);
and U2637 (N_2637,N_69,N_1582);
nor U2638 (N_2638,N_2011,N_1200);
and U2639 (N_2639,N_628,N_535);
or U2640 (N_2640,N_168,N_1107);
nand U2641 (N_2641,N_1318,N_728);
or U2642 (N_2642,N_1751,N_1614);
or U2643 (N_2643,N_259,N_444);
and U2644 (N_2644,N_1444,N_503);
nand U2645 (N_2645,N_1033,N_2094);
xor U2646 (N_2646,N_1625,N_586);
or U2647 (N_2647,N_403,N_492);
nor U2648 (N_2648,N_1765,N_1650);
or U2649 (N_2649,N_588,N_981);
or U2650 (N_2650,N_2328,N_490);
xnor U2651 (N_2651,N_1103,N_541);
or U2652 (N_2652,N_1264,N_1006);
nor U2653 (N_2653,N_935,N_619);
and U2654 (N_2654,N_2305,N_2162);
xnor U2655 (N_2655,N_930,N_962);
and U2656 (N_2656,N_1983,N_769);
and U2657 (N_2657,N_1645,N_1904);
and U2658 (N_2658,N_593,N_557);
nand U2659 (N_2659,N_1730,N_1276);
and U2660 (N_2660,N_1629,N_1982);
and U2661 (N_2661,N_1272,N_1972);
xnor U2662 (N_2662,N_364,N_1399);
xnor U2663 (N_2663,N_288,N_1579);
and U2664 (N_2664,N_1581,N_2103);
nor U2665 (N_2665,N_1875,N_295);
xnor U2666 (N_2666,N_1583,N_1646);
nor U2667 (N_2667,N_1083,N_1710);
xnor U2668 (N_2668,N_835,N_2038);
nand U2669 (N_2669,N_388,N_2319);
and U2670 (N_2670,N_297,N_1994);
nor U2671 (N_2671,N_1363,N_706);
xor U2672 (N_2672,N_1409,N_1989);
nor U2673 (N_2673,N_1111,N_990);
and U2674 (N_2674,N_79,N_1138);
xnor U2675 (N_2675,N_615,N_1812);
nand U2676 (N_2676,N_105,N_1122);
xnor U2677 (N_2677,N_2022,N_2213);
or U2678 (N_2678,N_2435,N_668);
or U2679 (N_2679,N_491,N_1852);
and U2680 (N_2680,N_783,N_1572);
or U2681 (N_2681,N_215,N_1708);
nor U2682 (N_2682,N_1615,N_12);
nor U2683 (N_2683,N_1032,N_1743);
nand U2684 (N_2684,N_1238,N_2452);
nor U2685 (N_2685,N_2163,N_1558);
nor U2686 (N_2686,N_815,N_1557);
nand U2687 (N_2687,N_2314,N_678);
xnor U2688 (N_2688,N_1973,N_1745);
nand U2689 (N_2689,N_1452,N_2420);
nand U2690 (N_2690,N_2484,N_59);
nand U2691 (N_2691,N_440,N_521);
nand U2692 (N_2692,N_127,N_149);
nand U2693 (N_2693,N_948,N_1737);
or U2694 (N_2694,N_19,N_1736);
xor U2695 (N_2695,N_352,N_1437);
xnor U2696 (N_2696,N_1332,N_464);
nand U2697 (N_2697,N_554,N_468);
and U2698 (N_2698,N_919,N_1522);
nor U2699 (N_2699,N_1011,N_763);
or U2700 (N_2700,N_2296,N_1000);
xor U2701 (N_2701,N_1054,N_1115);
or U2702 (N_2702,N_1550,N_2379);
and U2703 (N_2703,N_1833,N_747);
nand U2704 (N_2704,N_2090,N_2072);
xor U2705 (N_2705,N_2116,N_2496);
and U2706 (N_2706,N_174,N_697);
and U2707 (N_2707,N_1469,N_2451);
xor U2708 (N_2708,N_1246,N_1990);
xor U2709 (N_2709,N_1119,N_229);
nand U2710 (N_2710,N_734,N_2200);
nand U2711 (N_2711,N_1043,N_2027);
nor U2712 (N_2712,N_1209,N_986);
or U2713 (N_2713,N_2251,N_943);
xor U2714 (N_2714,N_1515,N_1089);
nand U2715 (N_2715,N_2061,N_556);
and U2716 (N_2716,N_110,N_1357);
nor U2717 (N_2717,N_2316,N_888);
and U2718 (N_2718,N_1252,N_2143);
or U2719 (N_2719,N_942,N_594);
and U2720 (N_2720,N_1733,N_1075);
and U2721 (N_2721,N_1961,N_306);
or U2722 (N_2722,N_29,N_737);
xor U2723 (N_2723,N_1434,N_2210);
nor U2724 (N_2724,N_2,N_1499);
xor U2725 (N_2725,N_605,N_632);
and U2726 (N_2726,N_2494,N_1925);
nand U2727 (N_2727,N_1213,N_654);
nor U2728 (N_2728,N_1202,N_1128);
nor U2729 (N_2729,N_1394,N_926);
nor U2730 (N_2730,N_2015,N_775);
or U2731 (N_2731,N_96,N_1559);
and U2732 (N_2732,N_2398,N_170);
or U2733 (N_2733,N_128,N_209);
and U2734 (N_2734,N_198,N_1139);
xor U2735 (N_2735,N_1420,N_1347);
xor U2736 (N_2736,N_1647,N_273);
or U2737 (N_2737,N_477,N_1462);
and U2738 (N_2738,N_2421,N_2463);
xnor U2739 (N_2739,N_308,N_2455);
and U2740 (N_2740,N_361,N_1341);
or U2741 (N_2741,N_1300,N_182);
and U2742 (N_2742,N_2003,N_1761);
xnor U2743 (N_2743,N_777,N_650);
xnor U2744 (N_2744,N_1881,N_372);
and U2745 (N_2745,N_1204,N_1847);
nor U2746 (N_2746,N_1110,N_599);
and U2747 (N_2747,N_252,N_853);
nor U2748 (N_2748,N_573,N_980);
nor U2749 (N_2749,N_1471,N_1068);
or U2750 (N_2750,N_1150,N_1077);
nand U2751 (N_2751,N_2487,N_1482);
nor U2752 (N_2752,N_1305,N_516);
xor U2753 (N_2753,N_2209,N_1064);
nand U2754 (N_2754,N_1968,N_1664);
nand U2755 (N_2755,N_2023,N_1373);
nand U2756 (N_2756,N_1066,N_946);
nor U2757 (N_2757,N_2287,N_509);
nand U2758 (N_2758,N_1149,N_1142);
xnor U2759 (N_2759,N_1082,N_2255);
and U2760 (N_2760,N_2223,N_237);
or U2761 (N_2761,N_1447,N_889);
or U2762 (N_2762,N_1311,N_1350);
xnor U2763 (N_2763,N_2249,N_1601);
nor U2764 (N_2764,N_1884,N_1084);
nor U2765 (N_2765,N_1281,N_1376);
xnor U2766 (N_2766,N_2067,N_999);
or U2767 (N_2767,N_2371,N_2203);
nor U2768 (N_2768,N_1263,N_913);
or U2769 (N_2769,N_1308,N_1895);
and U2770 (N_2770,N_1954,N_2068);
or U2771 (N_2771,N_1519,N_2397);
nor U2772 (N_2772,N_2097,N_303);
xnor U2773 (N_2773,N_1151,N_1596);
nand U2774 (N_2774,N_1548,N_2221);
nand U2775 (N_2775,N_253,N_1182);
nor U2776 (N_2776,N_157,N_695);
or U2777 (N_2777,N_595,N_2177);
xnor U2778 (N_2778,N_1857,N_1807);
nor U2779 (N_2779,N_1223,N_279);
nand U2780 (N_2780,N_1231,N_2180);
xor U2781 (N_2781,N_1889,N_2104);
or U2782 (N_2782,N_1342,N_2004);
xnor U2783 (N_2783,N_772,N_1689);
nand U2784 (N_2784,N_27,N_790);
or U2785 (N_2785,N_679,N_936);
nand U2786 (N_2786,N_1040,N_450);
nor U2787 (N_2787,N_151,N_667);
or U2788 (N_2788,N_1836,N_474);
and U2789 (N_2789,N_65,N_2332);
and U2790 (N_2790,N_208,N_848);
nor U2791 (N_2791,N_720,N_424);
and U2792 (N_2792,N_660,N_1101);
and U2793 (N_2793,N_2222,N_2217);
and U2794 (N_2794,N_498,N_1127);
and U2795 (N_2795,N_2357,N_2124);
nor U2796 (N_2796,N_1188,N_2119);
and U2797 (N_2797,N_785,N_1436);
nand U2798 (N_2798,N_2432,N_1277);
and U2799 (N_2799,N_1878,N_1796);
and U2800 (N_2800,N_1156,N_1161);
nand U2801 (N_2801,N_2241,N_1912);
nor U2802 (N_2802,N_367,N_1458);
nand U2803 (N_2803,N_1502,N_1406);
nand U2804 (N_2804,N_1766,N_505);
or U2805 (N_2805,N_567,N_1735);
nor U2806 (N_2806,N_275,N_2031);
or U2807 (N_2807,N_1919,N_85);
or U2808 (N_2808,N_1283,N_1791);
or U2809 (N_2809,N_2252,N_414);
and U2810 (N_2810,N_419,N_560);
nor U2811 (N_2811,N_371,N_2363);
nand U2812 (N_2812,N_1454,N_2254);
nor U2813 (N_2813,N_1226,N_1996);
or U2814 (N_2814,N_687,N_579);
xor U2815 (N_2815,N_315,N_2245);
nor U2816 (N_2816,N_1254,N_1544);
and U2817 (N_2817,N_1768,N_2340);
nand U2818 (N_2818,N_2130,N_1459);
or U2819 (N_2819,N_1563,N_150);
nand U2820 (N_2820,N_1538,N_1099);
nor U2821 (N_2821,N_1224,N_609);
nor U2822 (N_2822,N_2157,N_2288);
and U2823 (N_2823,N_2204,N_1597);
nand U2824 (N_2824,N_1456,N_17);
and U2825 (N_2825,N_1913,N_991);
nand U2826 (N_2826,N_532,N_2189);
and U2827 (N_2827,N_375,N_647);
or U2828 (N_2828,N_607,N_236);
xnor U2829 (N_2829,N_696,N_376);
or U2830 (N_2830,N_2273,N_400);
nor U2831 (N_2831,N_2194,N_126);
nand U2832 (N_2832,N_2497,N_119);
nor U2833 (N_2833,N_1718,N_365);
or U2834 (N_2834,N_1975,N_1561);
and U2835 (N_2835,N_2449,N_304);
or U2836 (N_2836,N_2491,N_1594);
nor U2837 (N_2837,N_355,N_756);
nand U2838 (N_2838,N_88,N_89);
xor U2839 (N_2839,N_1903,N_1387);
or U2840 (N_2840,N_1916,N_1534);
nor U2841 (N_2841,N_2293,N_1414);
xor U2842 (N_2842,N_1484,N_1753);
nand U2843 (N_2843,N_1494,N_2342);
nor U2844 (N_2844,N_539,N_2201);
or U2845 (N_2845,N_1247,N_959);
nor U2846 (N_2846,N_1811,N_2257);
or U2847 (N_2847,N_1593,N_1957);
or U2848 (N_2848,N_1027,N_1815);
and U2849 (N_2849,N_771,N_2495);
nand U2850 (N_2850,N_1974,N_1724);
xor U2851 (N_2851,N_1838,N_1215);
and U2852 (N_2852,N_2458,N_1590);
nand U2853 (N_2853,N_495,N_759);
nand U2854 (N_2854,N_1653,N_1180);
and U2855 (N_2855,N_1349,N_245);
xor U2856 (N_2856,N_878,N_1845);
or U2857 (N_2857,N_1120,N_901);
nor U2858 (N_2858,N_49,N_1817);
xnor U2859 (N_2859,N_322,N_1539);
nand U2860 (N_2860,N_1404,N_54);
and U2861 (N_2861,N_1603,N_2469);
nand U2862 (N_2862,N_1290,N_791);
nand U2863 (N_2863,N_773,N_116);
nand U2864 (N_2864,N_1477,N_709);
nand U2865 (N_2865,N_373,N_2039);
xor U2866 (N_2866,N_787,N_604);
and U2867 (N_2867,N_2198,N_2450);
xor U2868 (N_2868,N_1942,N_1900);
xor U2869 (N_2869,N_1523,N_1905);
and U2870 (N_2870,N_461,N_1763);
nor U2871 (N_2871,N_2016,N_2114);
nand U2872 (N_2872,N_786,N_625);
nand U2873 (N_2873,N_722,N_638);
nor U2874 (N_2874,N_181,N_121);
nand U2875 (N_2875,N_2220,N_2171);
and U2876 (N_2876,N_1867,N_445);
nor U2877 (N_2877,N_486,N_2205);
nor U2878 (N_2878,N_243,N_1741);
nand U2879 (N_2879,N_1945,N_1163);
or U2880 (N_2880,N_2149,N_1048);
or U2881 (N_2881,N_891,N_2348);
nand U2882 (N_2882,N_738,N_575);
xnor U2883 (N_2883,N_1422,N_1685);
nor U2884 (N_2884,N_1822,N_1367);
and U2885 (N_2885,N_378,N_680);
and U2886 (N_2886,N_808,N_460);
or U2887 (N_2887,N_863,N_1179);
xnor U2888 (N_2888,N_2429,N_954);
nor U2889 (N_2889,N_778,N_223);
nand U2890 (N_2890,N_1344,N_363);
or U2891 (N_2891,N_1691,N_553);
nor U2892 (N_2892,N_2165,N_1545);
nand U2893 (N_2893,N_1829,N_2055);
xnor U2894 (N_2894,N_819,N_1160);
and U2895 (N_2895,N_2148,N_14);
nand U2896 (N_2896,N_2071,N_1728);
or U2897 (N_2897,N_1410,N_694);
nor U2898 (N_2898,N_1104,N_698);
and U2899 (N_2899,N_26,N_903);
xor U2900 (N_2900,N_578,N_1253);
nand U2901 (N_2901,N_864,N_1901);
and U2902 (N_2902,N_1891,N_809);
xor U2903 (N_2903,N_914,N_2034);
xnor U2904 (N_2904,N_2044,N_186);
xor U2905 (N_2905,N_812,N_2376);
and U2906 (N_2906,N_2014,N_2275);
nand U2907 (N_2907,N_830,N_1713);
or U2908 (N_2908,N_1712,N_101);
and U2909 (N_2909,N_2358,N_643);
xnor U2910 (N_2910,N_641,N_2401);
or U2911 (N_2911,N_1637,N_2286);
or U2912 (N_2912,N_2445,N_916);
and U2913 (N_2913,N_187,N_451);
or U2914 (N_2914,N_1937,N_1416);
or U2915 (N_2915,N_1525,N_2444);
or U2916 (N_2916,N_141,N_779);
nor U2917 (N_2917,N_1389,N_2112);
nand U2918 (N_2918,N_1662,N_231);
xor U2919 (N_2919,N_2285,N_1747);
nor U2920 (N_2920,N_2109,N_571);
nand U2921 (N_2921,N_1964,N_1532);
and U2922 (N_2922,N_2002,N_479);
and U2923 (N_2923,N_2471,N_2018);
xor U2924 (N_2924,N_2443,N_387);
xnor U2925 (N_2925,N_627,N_1962);
nor U2926 (N_2926,N_992,N_1057);
or U2927 (N_2927,N_1941,N_489);
nor U2928 (N_2928,N_1566,N_1880);
xnor U2929 (N_2929,N_1175,N_1856);
or U2930 (N_2930,N_309,N_768);
or U2931 (N_2931,N_824,N_1952);
nor U2932 (N_2932,N_854,N_1677);
or U2933 (N_2933,N_25,N_496);
or U2934 (N_2934,N_2425,N_82);
nand U2935 (N_2935,N_542,N_1805);
nor U2936 (N_2936,N_2141,N_2482);
nand U2937 (N_2937,N_1475,N_271);
or U2938 (N_2938,N_2416,N_816);
nor U2939 (N_2939,N_1227,N_330);
and U2940 (N_2940,N_2246,N_1176);
xnor U2941 (N_2941,N_433,N_736);
nand U2942 (N_2942,N_869,N_2297);
or U2943 (N_2943,N_1310,N_1449);
xnor U2944 (N_2944,N_434,N_860);
nand U2945 (N_2945,N_2446,N_1701);
nor U2946 (N_2946,N_2384,N_2440);
nor U2947 (N_2947,N_1652,N_480);
and U2948 (N_2948,N_454,N_865);
nor U2949 (N_2949,N_92,N_339);
xor U2950 (N_2950,N_481,N_793);
and U2951 (N_2951,N_1045,N_1682);
xnor U2952 (N_2952,N_1794,N_1148);
nor U2953 (N_2953,N_1560,N_533);
nand U2954 (N_2954,N_1488,N_1832);
nand U2955 (N_2955,N_1627,N_246);
and U2956 (N_2956,N_1038,N_2448);
nand U2957 (N_2957,N_1930,N_2391);
and U2958 (N_2958,N_1814,N_955);
nand U2959 (N_2959,N_1024,N_971);
xor U2960 (N_2960,N_527,N_610);
nand U2961 (N_2961,N_2152,N_247);
and U2962 (N_2962,N_2351,N_2490);
nor U2963 (N_2963,N_117,N_1825);
nand U2964 (N_2964,N_194,N_1663);
nand U2965 (N_2965,N_1154,N_37);
nand U2966 (N_2966,N_634,N_1478);
nor U2967 (N_2967,N_248,N_318);
nor U2968 (N_2968,N_1907,N_30);
xor U2969 (N_2969,N_1987,N_1036);
or U2970 (N_2970,N_983,N_1551);
nor U2971 (N_2971,N_2447,N_875);
xor U2972 (N_2972,N_1965,N_2231);
nor U2973 (N_2973,N_1896,N_1096);
or U2974 (N_2974,N_839,N_358);
xor U2975 (N_2975,N_1178,N_2475);
nand U2976 (N_2976,N_1927,N_1118);
nand U2977 (N_2977,N_576,N_154);
xor U2978 (N_2978,N_346,N_893);
xor U2979 (N_2979,N_859,N_263);
or U2980 (N_2980,N_621,N_319);
and U2981 (N_2981,N_699,N_1869);
or U2982 (N_2982,N_172,N_580);
nand U2983 (N_2983,N_2050,N_214);
nor U2984 (N_2984,N_918,N_1296);
or U2985 (N_2985,N_1804,N_1169);
nor U2986 (N_2986,N_193,N_2480);
or U2987 (N_2987,N_2106,N_1898);
xor U2988 (N_2988,N_2125,N_497);
and U2989 (N_2989,N_293,N_1657);
nand U2990 (N_2990,N_2408,N_360);
xnor U2991 (N_2991,N_2183,N_1210);
xnor U2992 (N_2992,N_1014,N_951);
xor U2993 (N_2993,N_1088,N_1321);
or U2994 (N_2994,N_169,N_5);
nand U2995 (N_2995,N_1286,N_289);
nand U2996 (N_2996,N_2405,N_540);
xnor U2997 (N_2997,N_1719,N_162);
xor U2998 (N_2998,N_1021,N_2309);
and U2999 (N_2999,N_2105,N_2290);
xor U3000 (N_3000,N_2374,N_1131);
nand U3001 (N_3001,N_1186,N_2035);
and U3002 (N_3002,N_2431,N_2282);
and U3003 (N_3003,N_2486,N_1280);
nand U3004 (N_3004,N_2054,N_565);
and U3005 (N_3005,N_792,N_842);
or U3006 (N_3006,N_871,N_1626);
or U3007 (N_3007,N_671,N_453);
xor U3008 (N_3008,N_2247,N_2084);
and U3009 (N_3009,N_1121,N_1739);
nor U3010 (N_3010,N_1065,N_2234);
and U3011 (N_3011,N_1678,N_1319);
or U3012 (N_3012,N_644,N_1383);
nor U3013 (N_3013,N_201,N_290);
or U3014 (N_3014,N_1181,N_2235);
nand U3015 (N_3015,N_675,N_645);
nor U3016 (N_3016,N_1050,N_2059);
xor U3017 (N_3017,N_255,N_590);
xor U3018 (N_3018,N_897,N_749);
xnor U3019 (N_3019,N_1438,N_125);
and U3020 (N_3020,N_266,N_1177);
nor U3021 (N_3021,N_2188,N_40);
nor U3022 (N_3022,N_1810,N_1316);
or U3023 (N_3023,N_1849,N_1451);
or U3024 (N_3024,N_1808,N_1470);
nand U3025 (N_3025,N_1669,N_1585);
nor U3026 (N_3026,N_1556,N_592);
xor U3027 (N_3027,N_2179,N_1086);
nor U3028 (N_3028,N_1102,N_1700);
or U3029 (N_3029,N_2229,N_630);
and U3030 (N_3030,N_639,N_390);
nor U3031 (N_3031,N_46,N_254);
nor U3032 (N_3032,N_928,N_1442);
xnor U3033 (N_3033,N_1015,N_2301);
or U3034 (N_3034,N_408,N_1547);
nor U3035 (N_3035,N_807,N_1702);
or U3036 (N_3036,N_997,N_2409);
and U3037 (N_3037,N_499,N_1846);
xnor U3038 (N_3038,N_1506,N_2383);
xnor U3039 (N_3039,N_591,N_423);
xor U3040 (N_3040,N_118,N_761);
or U3041 (N_3041,N_1417,N_2372);
nand U3042 (N_3042,N_183,N_844);
or U3043 (N_3043,N_1429,N_1543);
xnor U3044 (N_3044,N_338,N_572);
nand U3045 (N_3045,N_1588,N_351);
nor U3046 (N_3046,N_1516,N_191);
xor U3047 (N_3047,N_2184,N_2407);
nor U3048 (N_3048,N_323,N_1369);
nor U3049 (N_3049,N_1168,N_2100);
xor U3050 (N_3050,N_2274,N_2268);
and U3051 (N_3051,N_1235,N_530);
xnor U3052 (N_3052,N_1498,N_1823);
nor U3053 (N_3053,N_1136,N_1997);
or U3054 (N_3054,N_748,N_862);
nor U3055 (N_3055,N_316,N_510);
nor U3056 (N_3056,N_447,N_1278);
and U3057 (N_3057,N_2041,N_1874);
nand U3058 (N_3058,N_845,N_1190);
nor U3059 (N_3059,N_190,N_826);
or U3060 (N_3060,N_1782,N_2207);
or U3061 (N_3061,N_120,N_2216);
nor U3062 (N_3062,N_39,N_1091);
and U3063 (N_3063,N_2377,N_292);
and U3064 (N_3064,N_550,N_2300);
or U3065 (N_3065,N_988,N_2347);
nand U3066 (N_3066,N_2412,N_1520);
and U3067 (N_3067,N_384,N_473);
xor U3068 (N_3068,N_1025,N_1443);
xnor U3069 (N_3069,N_1688,N_2005);
nand U3070 (N_3070,N_410,N_83);
or U3071 (N_3071,N_2426,N_1871);
nor U3072 (N_3072,N_833,N_416);
nand U3073 (N_3073,N_1779,N_488);
nor U3074 (N_3074,N_298,N_350);
and U3075 (N_3075,N_1549,N_2258);
nor U3076 (N_3076,N_2091,N_2338);
nor U3077 (N_3077,N_391,N_1801);
xor U3078 (N_3078,N_1671,N_109);
xnor U3079 (N_3079,N_87,N_1613);
xor U3080 (N_3080,N_1966,N_2390);
xor U3081 (N_3081,N_472,N_2199);
or U3082 (N_3082,N_1140,N_2352);
nand U3083 (N_3083,N_1375,N_383);
nor U3084 (N_3084,N_264,N_1518);
and U3085 (N_3085,N_837,N_1013);
nand U3086 (N_3086,N_1052,N_283);
nor U3087 (N_3087,N_721,N_2240);
and U3088 (N_3088,N_754,N_377);
nor U3089 (N_3089,N_940,N_885);
xor U3090 (N_3090,N_1978,N_739);
or U3091 (N_3091,N_278,N_258);
xor U3092 (N_3092,N_921,N_558);
xor U3093 (N_3093,N_965,N_1267);
and U3094 (N_3094,N_138,N_1595);
xnor U3095 (N_3095,N_1078,N_20);
nor U3096 (N_3096,N_1893,N_2312);
nor U3097 (N_3097,N_269,N_537);
nand U3098 (N_3098,N_2190,N_393);
or U3099 (N_3099,N_1521,N_1468);
and U3100 (N_3100,N_232,N_1126);
and U3101 (N_3101,N_683,N_1325);
nand U3102 (N_3102,N_2488,N_1312);
xor U3103 (N_3103,N_933,N_1890);
or U3104 (N_3104,N_2259,N_1500);
and U3105 (N_3105,N_343,N_846);
or U3106 (N_3106,N_890,N_345);
or U3107 (N_3107,N_1665,N_2065);
and U3108 (N_3108,N_2058,N_616);
nor U3109 (N_3109,N_710,N_1797);
nor U3110 (N_3110,N_1028,N_2156);
and U3111 (N_3111,N_836,N_2239);
xnor U3112 (N_3112,N_2232,N_442);
or U3113 (N_3113,N_953,N_1294);
nor U3114 (N_3114,N_915,N_1658);
or U3115 (N_3115,N_1017,N_1419);
and U3116 (N_3116,N_723,N_1764);
nor U3117 (N_3117,N_484,N_244);
or U3118 (N_3118,N_1222,N_2253);
nand U3119 (N_3119,N_2279,N_1586);
xnor U3120 (N_3120,N_2113,N_476);
nor U3121 (N_3121,N_2437,N_7);
nor U3122 (N_3122,N_1988,N_1395);
xor U3123 (N_3123,N_16,N_905);
or U3124 (N_3124,N_2263,N_1565);
nand U3125 (N_3125,N_1654,N_507);
nor U3126 (N_3126,N_142,N_1362);
nor U3127 (N_3127,N_2327,N_1309);
or U3128 (N_3128,N_1514,N_1711);
nor U3129 (N_3129,N_2434,N_506);
xnor U3130 (N_3130,N_536,N_1604);
nor U3131 (N_3131,N_1249,N_430);
xnor U3132 (N_3132,N_2070,N_2032);
nor U3133 (N_3133,N_1124,N_2233);
nor U3134 (N_3134,N_1298,N_1165);
xor U3135 (N_3135,N_1287,N_294);
and U3136 (N_3136,N_299,N_167);
or U3137 (N_3137,N_1479,N_711);
nor U3138 (N_3138,N_789,N_906);
nand U3139 (N_3139,N_163,N_898);
or U3140 (N_3140,N_2472,N_780);
nand U3141 (N_3141,N_873,N_2419);
nor U3142 (N_3142,N_944,N_1029);
nand U3143 (N_3143,N_2395,N_544);
nor U3144 (N_3144,N_1809,N_1504);
or U3145 (N_3145,N_1773,N_1378);
nand U3146 (N_3146,N_1800,N_794);
xnor U3147 (N_3147,N_2410,N_2186);
nand U3148 (N_3148,N_685,N_196);
xnor U3149 (N_3149,N_2260,N_847);
or U3150 (N_3150,N_1125,N_874);
nand U3151 (N_3151,N_2359,N_1034);
nor U3152 (N_3152,N_1173,N_1306);
nand U3153 (N_3153,N_2008,N_1783);
nor U3154 (N_3154,N_2176,N_33);
or U3155 (N_3155,N_1750,N_1839);
nor U3156 (N_3156,N_690,N_585);
or U3157 (N_3157,N_385,N_1777);
or U3158 (N_3158,N_185,N_2168);
or U3159 (N_3159,N_534,N_64);
nor U3160 (N_3160,N_189,N_1827);
and U3161 (N_3161,N_284,N_1170);
or U3162 (N_3162,N_129,N_1053);
xor U3163 (N_3163,N_1164,N_2080);
nand U3164 (N_3164,N_2313,N_867);
nor U3165 (N_3165,N_1007,N_2441);
nor U3166 (N_3166,N_97,N_282);
nor U3167 (N_3167,N_1740,N_887);
and U3168 (N_3168,N_1303,N_1265);
or U3169 (N_3169,N_581,N_569);
nand U3170 (N_3170,N_1245,N_1693);
and U3171 (N_3171,N_1114,N_311);
or U3172 (N_3172,N_2028,N_331);
nand U3173 (N_3173,N_1806,N_1944);
nand U3174 (N_3174,N_2380,N_985);
xor U3175 (N_3175,N_561,N_934);
or U3176 (N_3176,N_850,N_2402);
xnor U3177 (N_3177,N_9,N_731);
nand U3178 (N_3178,N_1517,N_970);
nand U3179 (N_3179,N_1269,N_470);
and U3180 (N_3180,N_188,N_409);
or U3181 (N_3181,N_2436,N_455);
or U3182 (N_3182,N_2182,N_1628);
nand U3183 (N_3183,N_1167,N_1606);
and U3184 (N_3184,N_956,N_1695);
xor U3185 (N_3185,N_199,N_1567);
and U3186 (N_3186,N_814,N_601);
and U3187 (N_3187,N_1106,N_975);
nor U3188 (N_3188,N_1386,N_1947);
or U3189 (N_3189,N_600,N_1275);
xnor U3190 (N_3190,N_822,N_217);
or U3191 (N_3191,N_653,N_994);
and U3192 (N_3192,N_2191,N_274);
and U3193 (N_3193,N_1729,N_2108);
nand U3194 (N_3194,N_1971,N_2136);
xor U3195 (N_3195,N_1492,N_302);
and U3196 (N_3196,N_2013,N_2345);
and U3197 (N_3197,N_2062,N_1853);
and U3198 (N_3198,N_1776,N_2056);
nor U3199 (N_3199,N_2262,N_2063);
or U3200 (N_3200,N_1948,N_396);
xor U3201 (N_3201,N_18,N_1351);
xnor U3202 (N_3202,N_1720,N_967);
xnor U3203 (N_3203,N_2046,N_1324);
and U3204 (N_3204,N_1157,N_684);
nand U3205 (N_3205,N_1346,N_1023);
or U3206 (N_3206,N_1233,N_2289);
and U3207 (N_3207,N_2096,N_2388);
xor U3208 (N_3208,N_1986,N_1495);
xor U3209 (N_3209,N_2330,N_72);
and U3210 (N_3210,N_1570,N_272);
xnor U3211 (N_3211,N_2310,N_2158);
nand U3212 (N_3212,N_158,N_1323);
and U3213 (N_3213,N_2098,N_672);
nand U3214 (N_3214,N_1599,N_1490);
nor U3215 (N_3215,N_1788,N_973);
and U3216 (N_3216,N_471,N_406);
xor U3217 (N_3217,N_1251,N_770);
nor U3218 (N_3218,N_1918,N_2298);
nand U3219 (N_3219,N_374,N_1946);
nand U3220 (N_3220,N_285,N_640);
nor U3221 (N_3221,N_2036,N_1824);
nor U3222 (N_3222,N_1676,N_2224);
xor U3223 (N_3223,N_2474,N_693);
xnor U3224 (N_3224,N_1915,N_178);
and U3225 (N_3225,N_1906,N_598);
xnor U3226 (N_3226,N_1374,N_851);
and U3227 (N_3227,N_1413,N_238);
nor U3228 (N_3228,N_1589,N_1360);
nand U3229 (N_3229,N_1756,N_1274);
or U3230 (N_3230,N_1016,N_1917);
nor U3231 (N_3231,N_84,N_75);
nor U3232 (N_3232,N_2006,N_1929);
nor U3233 (N_3233,N_106,N_669);
and U3234 (N_3234,N_379,N_1153);
xnor U3235 (N_3235,N_2466,N_1059);
nor U3236 (N_3236,N_160,N_2043);
nand U3237 (N_3237,N_38,N_2118);
nand U3238 (N_3238,N_1307,N_543);
and U3239 (N_3239,N_2160,N_613);
xor U3240 (N_3240,N_1607,N_1232);
nor U3241 (N_3241,N_1831,N_2454);
xnor U3242 (N_3242,N_658,N_2007);
nand U3243 (N_3243,N_1392,N_932);
nand U3244 (N_3244,N_1787,N_317);
nand U3245 (N_3245,N_2331,N_1980);
nor U3246 (N_3246,N_77,N_344);
or U3247 (N_3247,N_1802,N_1820);
or U3248 (N_3248,N_466,N_61);
nand U3249 (N_3249,N_249,N_348);
and U3250 (N_3250,N_803,N_240);
nor U3251 (N_3251,N_947,N_465);
nor U3252 (N_3252,N_1618,N_799);
or U3253 (N_3253,N_1910,N_587);
or U3254 (N_3254,N_1976,N_2227);
nor U3255 (N_3255,N_462,N_211);
nor U3256 (N_3256,N_1651,N_562);
and U3257 (N_3257,N_1850,N_1183);
nand U3258 (N_3258,N_2457,N_457);
xor U3259 (N_3259,N_2140,N_1580);
and U3260 (N_3260,N_1631,N_1732);
xor U3261 (N_3261,N_1031,N_1273);
or U3262 (N_3262,N_2465,N_71);
xnor U3263 (N_3263,N_1792,N_3);
nor U3264 (N_3264,N_1639,N_1295);
nor U3265 (N_3265,N_1198,N_821);
xnor U3266 (N_3266,N_931,N_523);
xor U3267 (N_3267,N_2009,N_817);
nor U3268 (N_3268,N_1780,N_1171);
or U3269 (N_3269,N_133,N_602);
and U3270 (N_3270,N_1840,N_927);
nand U3271 (N_3271,N_1771,N_982);
xor U3272 (N_3272,N_287,N_60);
nand U3273 (N_3273,N_1062,N_441);
and U3274 (N_3274,N_877,N_1536);
nor U3275 (N_3275,N_312,N_1885);
or U3276 (N_3276,N_1921,N_1466);
xor U3277 (N_3277,N_90,N_2146);
nor U3278 (N_3278,N_886,N_281);
nand U3279 (N_3279,N_1667,N_957);
xor U3280 (N_3280,N_1147,N_132);
and U3281 (N_3281,N_1018,N_1854);
nand U3282 (N_3282,N_546,N_1240);
or U3283 (N_3283,N_362,N_1446);
and U3284 (N_3284,N_1746,N_806);
nor U3285 (N_3285,N_1366,N_2181);
nand U3286 (N_3286,N_1070,N_2476);
or U3287 (N_3287,N_413,N_2020);
nand U3288 (N_3288,N_2326,N_538);
nand U3289 (N_3289,N_1211,N_114);
or U3290 (N_3290,N_67,N_1834);
and U3291 (N_3291,N_788,N_2276);
nand U3292 (N_3292,N_782,N_1940);
xor U3293 (N_3293,N_740,N_1960);
nand U3294 (N_3294,N_1679,N_702);
or U3295 (N_3295,N_1400,N_68);
and U3296 (N_3296,N_2439,N_2499);
nand U3297 (N_3297,N_329,N_1899);
xor U3298 (N_3298,N_235,N_1953);
or U3299 (N_3299,N_501,N_1714);
nand U3300 (N_3300,N_2462,N_1546);
nand U3301 (N_3301,N_1218,N_412);
nand U3302 (N_3302,N_99,N_425);
and U3303 (N_3303,N_2117,N_829);
or U3304 (N_3304,N_2308,N_23);
xnor U3305 (N_3305,N_1398,N_1058);
nor U3306 (N_3306,N_2317,N_1005);
xnor U3307 (N_3307,N_1221,N_1174);
nor U3308 (N_3308,N_147,N_1592);
nor U3309 (N_3309,N_192,N_2172);
nand U3310 (N_3310,N_2366,N_336);
nand U3311 (N_3311,N_1302,N_929);
and U3312 (N_3312,N_1145,N_1865);
xor U3313 (N_3313,N_2369,N_66);
and U3314 (N_3314,N_2430,N_805);
and U3315 (N_3315,N_1977,N_1705);
or U3316 (N_3316,N_353,N_504);
nand U3317 (N_3317,N_280,N_335);
or U3318 (N_3318,N_1760,N_1476);
xnor U3319 (N_3319,N_2236,N_548);
or U3320 (N_3320,N_270,N_145);
and U3321 (N_3321,N_2001,N_1635);
xor U3322 (N_3322,N_2396,N_2461);
nor U3323 (N_3323,N_950,N_1784);
nor U3324 (N_3324,N_622,N_2370);
and U3325 (N_3325,N_1605,N_1541);
xnor U3326 (N_3326,N_1393,N_8);
and U3327 (N_3327,N_148,N_2211);
or U3328 (N_3328,N_210,N_1041);
xor U3329 (N_3329,N_1969,N_1821);
and U3330 (N_3330,N_2244,N_422);
xnor U3331 (N_3331,N_2088,N_478);
nor U3332 (N_3332,N_1528,N_1781);
and U3333 (N_3333,N_1754,N_880);
and U3334 (N_3334,N_1073,N_1087);
nand U3335 (N_3335,N_566,N_2248);
nor U3336 (N_3336,N_514,N_1061);
or U3337 (N_3337,N_974,N_2150);
and U3338 (N_3338,N_1199,N_517);
nor U3339 (N_3339,N_1841,N_528);
nor U3340 (N_3340,N_2375,N_1576);
or U3341 (N_3341,N_508,N_1587);
nand U3342 (N_3342,N_2074,N_2115);
nor U3343 (N_3343,N_421,N_2277);
xnor U3344 (N_3344,N_1461,N_314);
and U3345 (N_3345,N_1722,N_2322);
nand U3346 (N_3346,N_2318,N_883);
and U3347 (N_3347,N_563,N_139);
or U3348 (N_3348,N_2323,N_767);
and U3349 (N_3349,N_2237,N_631);
and U3350 (N_3350,N_1619,N_1855);
nand U3351 (N_3351,N_443,N_2266);
xnor U3352 (N_3352,N_881,N_674);
nor U3353 (N_3353,N_2242,N_909);
and U3354 (N_3354,N_1922,N_2367);
nor U3355 (N_3355,N_584,N_1624);
xor U3356 (N_3356,N_1870,N_1744);
and U3357 (N_3357,N_320,N_2362);
nor U3358 (N_3358,N_617,N_458);
xor U3359 (N_3359,N_228,N_977);
nor U3360 (N_3360,N_1909,N_1908);
or U3361 (N_3361,N_612,N_1577);
nor U3362 (N_3362,N_757,N_2438);
or U3363 (N_3363,N_1440,N_1859);
nor U3364 (N_3364,N_741,N_648);
xnor U3365 (N_3365,N_2075,N_603);
xor U3366 (N_3366,N_305,N_1706);
and U3367 (N_3367,N_1877,N_1);
nor U3368 (N_3368,N_2060,N_2399);
and U3369 (N_3369,N_752,N_2473);
nor U3370 (N_3370,N_712,N_1463);
nor U3371 (N_3371,N_993,N_718);
and U3372 (N_3372,N_1196,N_2368);
nand U3373 (N_3373,N_682,N_1397);
and U3374 (N_3374,N_123,N_1155);
and U3375 (N_3375,N_1686,N_1135);
or U3376 (N_3376,N_1010,N_984);
nand U3377 (N_3377,N_1241,N_1568);
and U3378 (N_3378,N_1472,N_1039);
xor U3379 (N_3379,N_515,N_784);
nand U3380 (N_3380,N_2133,N_104);
or U3381 (N_3381,N_715,N_2381);
nand U3382 (N_3382,N_407,N_774);
nor U3383 (N_3383,N_1230,N_1370);
or U3384 (N_3384,N_841,N_1079);
nand U3385 (N_3385,N_872,N_1936);
xnor U3386 (N_3386,N_2321,N_1648);
xnor U3387 (N_3387,N_1959,N_286);
nor U3388 (N_3388,N_437,N_2164);
or U3389 (N_3389,N_1289,N_2464);
and U3390 (N_3390,N_620,N_224);
xor U3391 (N_3391,N_884,N_966);
and U3392 (N_3392,N_1842,N_216);
and U3393 (N_3393,N_689,N_2373);
and U3394 (N_3394,N_1453,N_261);
xor U3395 (N_3395,N_2147,N_2353);
or U3396 (N_3396,N_1670,N_1610);
xnor U3397 (N_3397,N_2037,N_10);
xor U3398 (N_3398,N_95,N_239);
nand U3399 (N_3399,N_798,N_2029);
nor U3400 (N_3400,N_2159,N_1602);
nor U3401 (N_3401,N_2064,N_1288);
or U3402 (N_3402,N_1984,N_307);
nand U3403 (N_3403,N_44,N_742);
xnor U3404 (N_3404,N_1709,N_2196);
nor U3405 (N_3405,N_0,N_2000);
or U3406 (N_3406,N_1009,N_2069);
nor U3407 (N_3407,N_2132,N_958);
nand U3408 (N_3408,N_2382,N_159);
xor U3409 (N_3409,N_2456,N_100);
or U3410 (N_3410,N_1934,N_1234);
nand U3411 (N_3411,N_547,N_276);
nand U3412 (N_3412,N_1203,N_135);
or U3413 (N_3413,N_11,N_2197);
nand U3414 (N_3414,N_1844,N_1259);
nor U3415 (N_3415,N_2386,N_1584);
and U3416 (N_3416,N_727,N_765);
xor U3417 (N_3417,N_429,N_1109);
or U3418 (N_3418,N_825,N_1225);
xor U3419 (N_3419,N_1675,N_1866);
and U3420 (N_3420,N_758,N_389);
nor U3421 (N_3421,N_1162,N_91);
xnor U3422 (N_3422,N_428,N_2052);
or U3423 (N_3423,N_130,N_1330);
and U3424 (N_3424,N_426,N_1600);
or U3425 (N_3425,N_1622,N_1343);
or U3426 (N_3426,N_153,N_268);
nand U3427 (N_3427,N_606,N_2256);
and U3428 (N_3428,N_2178,N_1320);
and U3429 (N_3429,N_1428,N_2453);
nor U3430 (N_3430,N_112,N_2030);
xnor U3431 (N_3431,N_1266,N_1643);
and U3432 (N_3432,N_52,N_776);
and U3433 (N_3433,N_1661,N_448);
nor U3434 (N_3434,N_1450,N_1851);
and U3435 (N_3435,N_1432,N_53);
nand U3436 (N_3436,N_1248,N_729);
nand U3437 (N_3437,N_212,N_2339);
nor U3438 (N_3438,N_2294,N_583);
nand U3439 (N_3439,N_1100,N_2214);
nor U3440 (N_3440,N_840,N_2355);
xnor U3441 (N_3441,N_2083,N_93);
nand U3442 (N_3442,N_676,N_1803);
nand U3443 (N_3443,N_227,N_1935);
nand U3444 (N_3444,N_2012,N_2481);
and U3445 (N_3445,N_1044,N_2281);
xnor U3446 (N_3446,N_184,N_2226);
or U3447 (N_3447,N_1361,N_1455);
and U3448 (N_3448,N_1133,N_633);
nand U3449 (N_3449,N_1356,N_2406);
or U3450 (N_3450,N_746,N_334);
or U3451 (N_3451,N_941,N_1690);
xor U3452 (N_3452,N_32,N_511);
or U3453 (N_3453,N_1396,N_716);
nor U3454 (N_3454,N_750,N_500);
xnor U3455 (N_3455,N_177,N_519);
and U3456 (N_3456,N_820,N_493);
nand U3457 (N_3457,N_963,N_1345);
nand U3458 (N_3458,N_838,N_2175);
and U3459 (N_3459,N_2169,N_1216);
xor U3460 (N_3460,N_1049,N_70);
and U3461 (N_3461,N_1026,N_1790);
and U3462 (N_3462,N_762,N_1887);
or U3463 (N_3463,N_2139,N_1425);
nor U3464 (N_3464,N_1146,N_1046);
or U3465 (N_3465,N_1037,N_24);
nor U3466 (N_3466,N_1022,N_1507);
nand U3467 (N_3467,N_357,N_1260);
xnor U3468 (N_3468,N_642,N_1774);
xnor U3469 (N_3469,N_2137,N_1426);
xor U3470 (N_3470,N_2167,N_520);
nor U3471 (N_3471,N_707,N_902);
or U3472 (N_3472,N_1268,N_2333);
or U3473 (N_3473,N_1813,N_4);
xnor U3474 (N_3474,N_124,N_1876);
or U3475 (N_3475,N_666,N_1666);
and U3476 (N_3476,N_57,N_1640);
xor U3477 (N_3477,N_1819,N_1407);
xnor U3478 (N_3478,N_1681,N_1069);
xnor U3479 (N_3479,N_663,N_596);
xnor U3480 (N_3480,N_743,N_277);
or U3481 (N_3481,N_207,N_1158);
xor U3482 (N_3482,N_559,N_146);
nor U3483 (N_3483,N_1623,N_1554);
xor U3484 (N_3484,N_487,N_1501);
xor U3485 (N_3485,N_152,N_1193);
nor U3486 (N_3486,N_197,N_260);
nor U3487 (N_3487,N_250,N_76);
nor U3488 (N_3488,N_1928,N_618);
nand U3489 (N_3489,N_1527,N_952);
nor U3490 (N_3490,N_1883,N_726);
xor U3491 (N_3491,N_857,N_1421);
nor U3492 (N_3492,N_22,N_1228);
xor U3493 (N_3493,N_1423,N_2192);
nor U3494 (N_3494,N_513,N_1992);
or U3495 (N_3495,N_418,N_2138);
and U3496 (N_3496,N_156,N_904);
nor U3497 (N_3497,N_438,N_1638);
or U3498 (N_3498,N_140,N_1430);
and U3499 (N_3499,N_21,N_1818);
and U3500 (N_3500,N_368,N_218);
or U3501 (N_3501,N_2126,N_1415);
xnor U3502 (N_3502,N_2082,N_50);
nand U3503 (N_3503,N_1734,N_2269);
nor U3504 (N_3504,N_1239,N_1435);
or U3505 (N_3505,N_1642,N_1097);
and U3506 (N_3506,N_1920,N_910);
or U3507 (N_3507,N_1256,N_1795);
nor U3508 (N_3508,N_161,N_2343);
xor U3509 (N_3509,N_459,N_938);
nor U3510 (N_3510,N_1742,N_1786);
nand U3511 (N_3511,N_143,N_1313);
nand U3512 (N_3512,N_1493,N_131);
or U3513 (N_3513,N_2428,N_2212);
nor U3514 (N_3514,N_2498,N_15);
nor U3515 (N_3515,N_483,N_394);
and U3516 (N_3516,N_47,N_1933);
or U3517 (N_3517,N_1258,N_369);
and U3518 (N_3518,N_1143,N_1755);
or U3519 (N_3519,N_976,N_1334);
xnor U3520 (N_3520,N_1512,N_1098);
xor U3521 (N_3521,N_908,N_2272);
xor U3522 (N_3522,N_417,N_435);
and U3523 (N_3523,N_134,N_1914);
nand U3524 (N_3524,N_1879,N_405);
and U3525 (N_3525,N_1339,N_961);
nor U3526 (N_3526,N_1465,N_1612);
and U3527 (N_3527,N_2485,N_1093);
and U3528 (N_3528,N_2417,N_518);
nand U3529 (N_3529,N_1336,N_813);
or U3530 (N_3530,N_811,N_1485);
nand U3531 (N_3531,N_1229,N_1353);
nand U3532 (N_3532,N_2389,N_171);
or U3533 (N_3533,N_1329,N_1575);
nor U3534 (N_3534,N_597,N_233);
nand U3535 (N_3535,N_41,N_2042);
nand U3536 (N_3536,N_45,N_1074);
nand U3537 (N_3537,N_1237,N_1535);
nand U3538 (N_3538,N_552,N_1630);
xor U3539 (N_3539,N_1250,N_1873);
and U3540 (N_3540,N_882,N_2076);
nand U3541 (N_3541,N_549,N_1698);
xor U3542 (N_3542,N_673,N_2225);
or U3543 (N_3543,N_1056,N_855);
xor U3544 (N_3544,N_1951,N_251);
nand U3545 (N_3545,N_1457,N_1159);
and U3546 (N_3546,N_1391,N_2128);
and U3547 (N_3547,N_427,N_1503);
nor U3548 (N_3548,N_1731,N_1020);
nor U3549 (N_3549,N_2479,N_900);
and U3550 (N_3550,N_1236,N_717);
nand U3551 (N_3551,N_1282,N_380);
and U3552 (N_3552,N_2292,N_924);
or U3553 (N_3553,N_688,N_213);
or U3554 (N_3554,N_823,N_2193);
and U3555 (N_3555,N_221,N_1924);
xnor U3556 (N_3556,N_751,N_2202);
nor U3557 (N_3557,N_923,N_395);
and U3558 (N_3558,N_2051,N_512);
nor U3559 (N_3559,N_1789,N_1337);
nand U3560 (N_3560,N_714,N_1368);
xnor U3561 (N_3561,N_551,N_56);
nor U3562 (N_3562,N_2111,N_2102);
nor U3563 (N_3563,N_1055,N_1003);
and U3564 (N_3564,N_2356,N_662);
or U3565 (N_3565,N_341,N_1331);
and U3566 (N_3566,N_356,N_1704);
xnor U3567 (N_3567,N_1956,N_922);
nand U3568 (N_3568,N_436,N_646);
xnor U3569 (N_3569,N_1411,N_2385);
nand U3570 (N_3570,N_1105,N_1381);
and U3571 (N_3571,N_234,N_831);
xor U3572 (N_3572,N_1798,N_1364);
xnor U3573 (N_3573,N_467,N_1441);
or U3574 (N_3574,N_2107,N_629);
xnor U3575 (N_3575,N_2329,N_86);
or U3576 (N_3576,N_704,N_291);
xnor U3577 (N_3577,N_2081,N_1480);
nand U3578 (N_3578,N_2415,N_411);
nand U3579 (N_3579,N_1897,N_1769);
or U3580 (N_3580,N_173,N_1491);
or U3581 (N_3581,N_949,N_1144);
xor U3582 (N_3582,N_1355,N_703);
xor U3583 (N_3583,N_2280,N_420);
nor U3584 (N_3584,N_337,N_2478);
or U3585 (N_3585,N_2334,N_989);
and U3586 (N_3586,N_818,N_2127);
nand U3587 (N_3587,N_1835,N_895);
nand U3588 (N_3588,N_1207,N_522);
xnor U3589 (N_3589,N_1384,N_2078);
or U3590 (N_3590,N_1445,N_1979);
xor U3591 (N_3591,N_1609,N_402);
nand U3592 (N_3592,N_2134,N_1326);
xor U3593 (N_3593,N_1340,N_1967);
nand U3594 (N_3594,N_960,N_1660);
xnor U3595 (N_3595,N_1872,N_968);
xnor U3596 (N_3596,N_652,N_1757);
xor U3597 (N_3597,N_1684,N_1510);
and U3598 (N_3598,N_655,N_681);
or U3599 (N_3599,N_996,N_2283);
nand U3600 (N_3600,N_2299,N_1886);
xnor U3601 (N_3601,N_2219,N_849);
nor U3602 (N_3602,N_366,N_78);
nor U3603 (N_3603,N_635,N_802);
nand U3604 (N_3604,N_262,N_1063);
nand U3605 (N_3605,N_31,N_108);
xor U3606 (N_3606,N_1932,N_2142);
and U3607 (N_3607,N_1071,N_2144);
nand U3608 (N_3608,N_324,N_1943);
nor U3609 (N_3609,N_1793,N_656);
xor U3610 (N_3610,N_1864,N_74);
nand U3611 (N_3611,N_2270,N_2243);
nor U3612 (N_3612,N_1699,N_1697);
and U3613 (N_3613,N_1816,N_636);
and U3614 (N_3614,N_1214,N_2215);
nand U3615 (N_3615,N_1862,N_1489);
or U3616 (N_3616,N_206,N_2166);
or U3617 (N_3617,N_659,N_1051);
or U3618 (N_3618,N_2364,N_2057);
nand U3619 (N_3619,N_42,N_1081);
nor U3620 (N_3620,N_155,N_1187);
and U3621 (N_3621,N_1772,N_1418);
nor U3622 (N_3622,N_1656,N_858);
xnor U3623 (N_3623,N_1509,N_1192);
nand U3624 (N_3624,N_2361,N_242);
nand U3625 (N_3625,N_2019,N_115);
xnor U3626 (N_3626,N_876,N_797);
or U3627 (N_3627,N_1322,N_1372);
or U3628 (N_3628,N_2135,N_1317);
nand U3629 (N_3629,N_1072,N_987);
and U3630 (N_3630,N_2278,N_225);
and U3631 (N_3631,N_1134,N_2325);
or U3632 (N_3632,N_392,N_2271);
nand U3633 (N_3633,N_136,N_800);
and U3634 (N_3634,N_1726,N_1680);
nor U3635 (N_3635,N_972,N_894);
xor U3636 (N_3636,N_753,N_35);
nor U3637 (N_3637,N_1902,N_2206);
and U3638 (N_3638,N_1271,N_2161);
and U3639 (N_3639,N_1837,N_2025);
xor U3640 (N_3640,N_1448,N_670);
or U3641 (N_3641,N_1578,N_175);
xor U3642 (N_3642,N_2295,N_1598);
or U3643 (N_3643,N_2304,N_1348);
xnor U3644 (N_3644,N_475,N_1067);
or U3645 (N_3645,N_2121,N_2324);
or U3646 (N_3646,N_1861,N_2093);
and U3647 (N_3647,N_1950,N_1380);
nand U3648 (N_3648,N_180,N_1467);
nor U3649 (N_3649,N_2151,N_1291);
xnor U3650 (N_3650,N_1217,N_1608);
xnor U3651 (N_3651,N_1004,N_397);
nor U3652 (N_3652,N_705,N_1299);
nand U3653 (N_3653,N_1553,N_1030);
nor U3654 (N_3654,N_2337,N_456);
xnor U3655 (N_3655,N_657,N_81);
or U3656 (N_3656,N_730,N_164);
xor U3657 (N_3657,N_325,N_1212);
and U3658 (N_3658,N_6,N_1617);
and U3659 (N_3659,N_608,N_1108);
and U3660 (N_3660,N_1530,N_677);
nand U3661 (N_3661,N_1382,N_370);
and U3662 (N_3662,N_664,N_1762);
nor U3663 (N_3663,N_398,N_1117);
xor U3664 (N_3664,N_1255,N_386);
or U3665 (N_3665,N_1460,N_1843);
nor U3666 (N_3666,N_2303,N_2110);
nand U3667 (N_3667,N_1775,N_1555);
nand U3668 (N_3668,N_725,N_1511);
nor U3669 (N_3669,N_2238,N_2404);
xor U3670 (N_3670,N_340,N_2087);
or U3671 (N_3671,N_1092,N_1008);
nor U3672 (N_3672,N_2086,N_1894);
xnor U3673 (N_3673,N_1923,N_1129);
or U3674 (N_3674,N_568,N_804);
nor U3675 (N_3675,N_1970,N_2073);
and U3676 (N_3676,N_62,N_1858);
nand U3677 (N_3677,N_1242,N_1402);
xor U3678 (N_3678,N_2311,N_870);
and U3679 (N_3679,N_2411,N_1703);
nor U3680 (N_3680,N_1995,N_328);
nor U3681 (N_3681,N_1985,N_2010);
nand U3682 (N_3682,N_1655,N_43);
xor U3683 (N_3683,N_349,N_665);
nand U3684 (N_3684,N_1401,N_1707);
xor U3685 (N_3685,N_1674,N_2185);
and U3686 (N_3686,N_2250,N_868);
nand U3687 (N_3687,N_2145,N_1526);
or U3688 (N_3688,N_2394,N_2392);
nand U3689 (N_3689,N_176,N_2423);
xnor U3690 (N_3690,N_524,N_1830);
nor U3691 (N_3691,N_2195,N_719);
nand U3692 (N_3692,N_1529,N_98);
xnor U3693 (N_3693,N_2230,N_1293);
and U3694 (N_3694,N_1848,N_2026);
or U3695 (N_3695,N_2153,N_1938);
and U3696 (N_3696,N_2170,N_1573);
xor U3697 (N_3697,N_1863,N_1358);
nor U3698 (N_3698,N_2228,N_1113);
xor U3699 (N_3699,N_2045,N_1137);
xor U3700 (N_3700,N_222,N_13);
xor U3701 (N_3701,N_1439,N_1047);
or U3702 (N_3702,N_1388,N_2489);
and U3703 (N_3703,N_359,N_1012);
nand U3704 (N_3704,N_1184,N_1727);
nand U3705 (N_3705,N_2122,N_760);
nor U3706 (N_3706,N_195,N_1132);
nand U3707 (N_3707,N_1958,N_1668);
nand U3708 (N_3708,N_896,N_2393);
nor U3709 (N_3709,N_879,N_611);
xnor U3710 (N_3710,N_1564,N_1333);
nand U3711 (N_3711,N_1060,N_866);
nand U3712 (N_3712,N_1487,N_2208);
or U3713 (N_3713,N_2302,N_701);
xor U3714 (N_3714,N_1687,N_1778);
nand U3715 (N_3715,N_2095,N_1672);
and U3716 (N_3716,N_1694,N_1194);
xnor U3717 (N_3717,N_1279,N_708);
or U3718 (N_3718,N_964,N_700);
and U3719 (N_3719,N_1696,N_354);
and U3720 (N_3720,N_1166,N_1683);
nand U3721 (N_3721,N_570,N_1540);
xor U3722 (N_3722,N_1076,N_2341);
xnor U3723 (N_3723,N_733,N_1354);
xor U3724 (N_3724,N_2307,N_545);
or U3725 (N_3725,N_431,N_795);
nand U3726 (N_3726,N_1080,N_1185);
nor U3727 (N_3727,N_332,N_267);
nand U3728 (N_3728,N_1219,N_2017);
xnor U3729 (N_3729,N_1035,N_1963);
or U3730 (N_3730,N_2187,N_637);
or U3731 (N_3731,N_347,N_404);
nand U3732 (N_3732,N_2079,N_1496);
nor U3733 (N_3733,N_1673,N_1261);
or U3734 (N_3734,N_2360,N_691);
and U3735 (N_3735,N_1644,N_1636);
nor U3736 (N_3736,N_382,N_1001);
nor U3737 (N_3737,N_945,N_2099);
nor U3738 (N_3738,N_766,N_827);
or U3739 (N_3739,N_1172,N_1244);
nand U3740 (N_3740,N_256,N_1723);
and U3741 (N_3741,N_2424,N_861);
and U3742 (N_3742,N_2315,N_494);
xor U3743 (N_3743,N_2092,N_2129);
or U3744 (N_3744,N_1427,N_1377);
and U3745 (N_3745,N_1304,N_995);
nand U3746 (N_3746,N_2365,N_624);
or U3747 (N_3747,N_1390,N_1262);
nand U3748 (N_3748,N_48,N_1379);
nor U3749 (N_3749,N_1981,N_1431);
or U3750 (N_3750,N_1542,N_2479);
nand U3751 (N_3751,N_1563,N_113);
or U3752 (N_3752,N_407,N_198);
or U3753 (N_3753,N_370,N_376);
nand U3754 (N_3754,N_823,N_2296);
xor U3755 (N_3755,N_261,N_1983);
xor U3756 (N_3756,N_1090,N_1614);
xor U3757 (N_3757,N_1515,N_2463);
or U3758 (N_3758,N_3,N_2462);
or U3759 (N_3759,N_1450,N_1922);
or U3760 (N_3760,N_111,N_515);
nand U3761 (N_3761,N_2213,N_2240);
xnor U3762 (N_3762,N_1267,N_2109);
and U3763 (N_3763,N_1833,N_1904);
xor U3764 (N_3764,N_1392,N_641);
and U3765 (N_3765,N_2026,N_688);
and U3766 (N_3766,N_924,N_1624);
xor U3767 (N_3767,N_808,N_505);
and U3768 (N_3768,N_9,N_1840);
nor U3769 (N_3769,N_1067,N_856);
nand U3770 (N_3770,N_682,N_58);
nand U3771 (N_3771,N_1667,N_23);
nor U3772 (N_3772,N_1845,N_2155);
or U3773 (N_3773,N_1318,N_2036);
nor U3774 (N_3774,N_1029,N_2436);
or U3775 (N_3775,N_2154,N_1002);
nand U3776 (N_3776,N_2288,N_594);
or U3777 (N_3777,N_37,N_576);
xnor U3778 (N_3778,N_2261,N_633);
xnor U3779 (N_3779,N_183,N_1404);
nor U3780 (N_3780,N_1907,N_174);
or U3781 (N_3781,N_623,N_1511);
nor U3782 (N_3782,N_833,N_1252);
nand U3783 (N_3783,N_1115,N_21);
or U3784 (N_3784,N_2102,N_1985);
or U3785 (N_3785,N_1545,N_1960);
and U3786 (N_3786,N_1521,N_1151);
and U3787 (N_3787,N_1230,N_729);
and U3788 (N_3788,N_2205,N_1922);
and U3789 (N_3789,N_462,N_825);
xnor U3790 (N_3790,N_789,N_672);
nor U3791 (N_3791,N_1328,N_1443);
nor U3792 (N_3792,N_1490,N_1779);
xnor U3793 (N_3793,N_1182,N_1261);
or U3794 (N_3794,N_1554,N_1117);
or U3795 (N_3795,N_1795,N_1570);
and U3796 (N_3796,N_565,N_501);
nor U3797 (N_3797,N_2218,N_449);
xor U3798 (N_3798,N_2469,N_2262);
xor U3799 (N_3799,N_551,N_479);
or U3800 (N_3800,N_576,N_1072);
nor U3801 (N_3801,N_9,N_413);
or U3802 (N_3802,N_342,N_2349);
or U3803 (N_3803,N_2424,N_549);
nand U3804 (N_3804,N_1394,N_1516);
xnor U3805 (N_3805,N_419,N_1413);
xor U3806 (N_3806,N_832,N_774);
or U3807 (N_3807,N_791,N_880);
or U3808 (N_3808,N_156,N_1077);
or U3809 (N_3809,N_207,N_521);
and U3810 (N_3810,N_2444,N_693);
and U3811 (N_3811,N_155,N_996);
nand U3812 (N_3812,N_1086,N_93);
nor U3813 (N_3813,N_2337,N_888);
and U3814 (N_3814,N_1443,N_855);
nor U3815 (N_3815,N_1906,N_1467);
xor U3816 (N_3816,N_971,N_586);
nor U3817 (N_3817,N_1391,N_1245);
nor U3818 (N_3818,N_1747,N_2253);
and U3819 (N_3819,N_795,N_2492);
or U3820 (N_3820,N_2235,N_939);
nor U3821 (N_3821,N_1187,N_2297);
nor U3822 (N_3822,N_2461,N_469);
xor U3823 (N_3823,N_2070,N_780);
or U3824 (N_3824,N_391,N_512);
xor U3825 (N_3825,N_2239,N_2133);
and U3826 (N_3826,N_2087,N_2209);
or U3827 (N_3827,N_1847,N_306);
nor U3828 (N_3828,N_1571,N_498);
nor U3829 (N_3829,N_792,N_2440);
nor U3830 (N_3830,N_1847,N_1346);
nor U3831 (N_3831,N_352,N_1819);
or U3832 (N_3832,N_2253,N_2428);
nor U3833 (N_3833,N_1936,N_1840);
xor U3834 (N_3834,N_1838,N_1169);
xnor U3835 (N_3835,N_1885,N_1948);
and U3836 (N_3836,N_2430,N_1671);
or U3837 (N_3837,N_1757,N_1713);
or U3838 (N_3838,N_115,N_998);
xor U3839 (N_3839,N_1762,N_1040);
xnor U3840 (N_3840,N_1902,N_1654);
xor U3841 (N_3841,N_1102,N_1336);
and U3842 (N_3842,N_1893,N_1483);
or U3843 (N_3843,N_358,N_2094);
and U3844 (N_3844,N_162,N_1515);
or U3845 (N_3845,N_1787,N_856);
and U3846 (N_3846,N_2169,N_2034);
or U3847 (N_3847,N_1242,N_734);
nand U3848 (N_3848,N_404,N_1430);
nor U3849 (N_3849,N_1475,N_1085);
and U3850 (N_3850,N_2443,N_1422);
xor U3851 (N_3851,N_140,N_583);
nand U3852 (N_3852,N_101,N_850);
nor U3853 (N_3853,N_2484,N_1843);
or U3854 (N_3854,N_1177,N_1383);
nor U3855 (N_3855,N_904,N_2078);
nand U3856 (N_3856,N_1156,N_2078);
nor U3857 (N_3857,N_649,N_1006);
nand U3858 (N_3858,N_1084,N_56);
xnor U3859 (N_3859,N_1953,N_1260);
or U3860 (N_3860,N_871,N_779);
or U3861 (N_3861,N_1518,N_2390);
or U3862 (N_3862,N_1927,N_822);
nand U3863 (N_3863,N_1817,N_113);
and U3864 (N_3864,N_2233,N_2064);
xnor U3865 (N_3865,N_629,N_746);
xor U3866 (N_3866,N_2181,N_397);
or U3867 (N_3867,N_2278,N_1698);
and U3868 (N_3868,N_1281,N_270);
nand U3869 (N_3869,N_63,N_2375);
and U3870 (N_3870,N_1433,N_1474);
xnor U3871 (N_3871,N_1449,N_1030);
or U3872 (N_3872,N_499,N_1419);
and U3873 (N_3873,N_2459,N_1284);
and U3874 (N_3874,N_1912,N_1565);
nand U3875 (N_3875,N_591,N_467);
or U3876 (N_3876,N_2442,N_1803);
nor U3877 (N_3877,N_2459,N_11);
xor U3878 (N_3878,N_1700,N_619);
or U3879 (N_3879,N_1959,N_1362);
nand U3880 (N_3880,N_375,N_1392);
nor U3881 (N_3881,N_1689,N_121);
nor U3882 (N_3882,N_2361,N_685);
xnor U3883 (N_3883,N_55,N_1650);
nor U3884 (N_3884,N_1576,N_1820);
xnor U3885 (N_3885,N_1895,N_955);
and U3886 (N_3886,N_771,N_119);
xnor U3887 (N_3887,N_1145,N_609);
or U3888 (N_3888,N_372,N_806);
nor U3889 (N_3889,N_1878,N_926);
and U3890 (N_3890,N_109,N_229);
nand U3891 (N_3891,N_1310,N_2462);
nand U3892 (N_3892,N_2015,N_1260);
and U3893 (N_3893,N_987,N_75);
nand U3894 (N_3894,N_859,N_356);
and U3895 (N_3895,N_793,N_1483);
xor U3896 (N_3896,N_85,N_1196);
or U3897 (N_3897,N_24,N_360);
nor U3898 (N_3898,N_1263,N_397);
or U3899 (N_3899,N_1854,N_534);
nor U3900 (N_3900,N_2364,N_1346);
and U3901 (N_3901,N_105,N_1175);
and U3902 (N_3902,N_1407,N_896);
xor U3903 (N_3903,N_2472,N_972);
nand U3904 (N_3904,N_1048,N_1956);
xnor U3905 (N_3905,N_1876,N_1751);
or U3906 (N_3906,N_1339,N_1098);
or U3907 (N_3907,N_64,N_1961);
xor U3908 (N_3908,N_338,N_2140);
nor U3909 (N_3909,N_426,N_207);
nor U3910 (N_3910,N_593,N_1879);
nor U3911 (N_3911,N_2021,N_198);
nor U3912 (N_3912,N_335,N_321);
or U3913 (N_3913,N_171,N_433);
xnor U3914 (N_3914,N_2032,N_1473);
nand U3915 (N_3915,N_1516,N_956);
nand U3916 (N_3916,N_2222,N_2037);
xor U3917 (N_3917,N_60,N_1253);
nor U3918 (N_3918,N_1971,N_1815);
nand U3919 (N_3919,N_1951,N_1985);
and U3920 (N_3920,N_224,N_2269);
or U3921 (N_3921,N_2273,N_1913);
or U3922 (N_3922,N_2434,N_482);
nor U3923 (N_3923,N_1070,N_2490);
or U3924 (N_3924,N_1706,N_730);
and U3925 (N_3925,N_1929,N_562);
nand U3926 (N_3926,N_2409,N_2065);
and U3927 (N_3927,N_1859,N_2055);
xnor U3928 (N_3928,N_110,N_552);
nand U3929 (N_3929,N_1549,N_1443);
or U3930 (N_3930,N_300,N_1723);
nand U3931 (N_3931,N_851,N_610);
nand U3932 (N_3932,N_2419,N_2165);
and U3933 (N_3933,N_2482,N_55);
xnor U3934 (N_3934,N_319,N_2203);
or U3935 (N_3935,N_538,N_2418);
and U3936 (N_3936,N_244,N_1970);
nand U3937 (N_3937,N_1028,N_2448);
or U3938 (N_3938,N_544,N_1373);
xor U3939 (N_3939,N_1369,N_1204);
or U3940 (N_3940,N_484,N_2154);
nor U3941 (N_3941,N_347,N_1633);
or U3942 (N_3942,N_1141,N_325);
or U3943 (N_3943,N_2262,N_1129);
nor U3944 (N_3944,N_2302,N_1110);
nand U3945 (N_3945,N_829,N_1985);
and U3946 (N_3946,N_822,N_82);
nand U3947 (N_3947,N_1049,N_1678);
xnor U3948 (N_3948,N_518,N_1485);
xnor U3949 (N_3949,N_642,N_1919);
xor U3950 (N_3950,N_2085,N_206);
nor U3951 (N_3951,N_2330,N_1294);
or U3952 (N_3952,N_649,N_1216);
nor U3953 (N_3953,N_2130,N_329);
nor U3954 (N_3954,N_2245,N_663);
xnor U3955 (N_3955,N_1538,N_2199);
nor U3956 (N_3956,N_1180,N_57);
and U3957 (N_3957,N_1088,N_664);
xnor U3958 (N_3958,N_2364,N_1265);
and U3959 (N_3959,N_2028,N_2236);
nor U3960 (N_3960,N_940,N_253);
nand U3961 (N_3961,N_560,N_2267);
nand U3962 (N_3962,N_2426,N_1287);
or U3963 (N_3963,N_407,N_1684);
or U3964 (N_3964,N_2151,N_1188);
xor U3965 (N_3965,N_835,N_1556);
or U3966 (N_3966,N_191,N_168);
nor U3967 (N_3967,N_2010,N_1474);
nor U3968 (N_3968,N_909,N_1592);
nand U3969 (N_3969,N_217,N_131);
or U3970 (N_3970,N_1315,N_234);
nor U3971 (N_3971,N_2457,N_1835);
nor U3972 (N_3972,N_2141,N_872);
nor U3973 (N_3973,N_272,N_827);
nor U3974 (N_3974,N_826,N_29);
nor U3975 (N_3975,N_1698,N_1232);
and U3976 (N_3976,N_960,N_1598);
xnor U3977 (N_3977,N_1138,N_1753);
xnor U3978 (N_3978,N_1412,N_1046);
xnor U3979 (N_3979,N_2067,N_684);
xnor U3980 (N_3980,N_2075,N_2031);
nor U3981 (N_3981,N_2045,N_793);
and U3982 (N_3982,N_749,N_1385);
xor U3983 (N_3983,N_1380,N_2440);
xor U3984 (N_3984,N_204,N_2202);
or U3985 (N_3985,N_866,N_1383);
nor U3986 (N_3986,N_2381,N_527);
and U3987 (N_3987,N_308,N_2410);
nor U3988 (N_3988,N_625,N_387);
and U3989 (N_3989,N_1935,N_2281);
or U3990 (N_3990,N_1000,N_1251);
nand U3991 (N_3991,N_1409,N_43);
and U3992 (N_3992,N_1288,N_418);
nand U3993 (N_3993,N_1695,N_1200);
and U3994 (N_3994,N_252,N_1827);
nand U3995 (N_3995,N_412,N_280);
and U3996 (N_3996,N_482,N_1490);
xnor U3997 (N_3997,N_1459,N_2189);
xor U3998 (N_3998,N_1815,N_391);
and U3999 (N_3999,N_1069,N_555);
nand U4000 (N_4000,N_546,N_687);
nor U4001 (N_4001,N_490,N_1115);
xor U4002 (N_4002,N_2363,N_790);
or U4003 (N_4003,N_866,N_1056);
nor U4004 (N_4004,N_2460,N_2223);
nor U4005 (N_4005,N_1831,N_1926);
and U4006 (N_4006,N_2461,N_1565);
nand U4007 (N_4007,N_1769,N_1872);
or U4008 (N_4008,N_558,N_298);
nand U4009 (N_4009,N_2257,N_1151);
nand U4010 (N_4010,N_932,N_137);
nand U4011 (N_4011,N_354,N_776);
nor U4012 (N_4012,N_110,N_667);
xor U4013 (N_4013,N_1675,N_441);
nor U4014 (N_4014,N_620,N_1883);
nand U4015 (N_4015,N_78,N_2019);
nor U4016 (N_4016,N_203,N_1102);
xor U4017 (N_4017,N_644,N_844);
nand U4018 (N_4018,N_115,N_1107);
nand U4019 (N_4019,N_417,N_2274);
nand U4020 (N_4020,N_867,N_896);
nor U4021 (N_4021,N_622,N_1406);
xnor U4022 (N_4022,N_1031,N_269);
xnor U4023 (N_4023,N_1649,N_254);
and U4024 (N_4024,N_1945,N_1670);
nor U4025 (N_4025,N_2267,N_2229);
and U4026 (N_4026,N_1927,N_1245);
nand U4027 (N_4027,N_1234,N_959);
nor U4028 (N_4028,N_1487,N_1949);
xor U4029 (N_4029,N_72,N_158);
and U4030 (N_4030,N_2152,N_706);
nor U4031 (N_4031,N_2269,N_613);
and U4032 (N_4032,N_1435,N_769);
nor U4033 (N_4033,N_1976,N_1593);
or U4034 (N_4034,N_779,N_1828);
nor U4035 (N_4035,N_2256,N_913);
and U4036 (N_4036,N_1457,N_1391);
xnor U4037 (N_4037,N_859,N_1306);
nand U4038 (N_4038,N_1088,N_1135);
xor U4039 (N_4039,N_429,N_2162);
or U4040 (N_4040,N_1995,N_355);
or U4041 (N_4041,N_215,N_1075);
xor U4042 (N_4042,N_2490,N_2454);
or U4043 (N_4043,N_1961,N_1732);
nand U4044 (N_4044,N_318,N_128);
or U4045 (N_4045,N_2075,N_2067);
nor U4046 (N_4046,N_385,N_602);
nor U4047 (N_4047,N_1289,N_2357);
and U4048 (N_4048,N_2400,N_2085);
nor U4049 (N_4049,N_1265,N_2156);
or U4050 (N_4050,N_2474,N_1952);
and U4051 (N_4051,N_2441,N_2308);
xnor U4052 (N_4052,N_966,N_743);
nand U4053 (N_4053,N_653,N_676);
or U4054 (N_4054,N_1644,N_1756);
and U4055 (N_4055,N_832,N_798);
xor U4056 (N_4056,N_2490,N_496);
and U4057 (N_4057,N_952,N_85);
or U4058 (N_4058,N_699,N_2092);
xor U4059 (N_4059,N_2094,N_1976);
nand U4060 (N_4060,N_324,N_800);
or U4061 (N_4061,N_1848,N_1854);
xnor U4062 (N_4062,N_390,N_2030);
nor U4063 (N_4063,N_2433,N_1069);
or U4064 (N_4064,N_2106,N_2049);
nor U4065 (N_4065,N_1853,N_2232);
nand U4066 (N_4066,N_1216,N_2437);
or U4067 (N_4067,N_762,N_2140);
nor U4068 (N_4068,N_1710,N_1898);
and U4069 (N_4069,N_949,N_29);
or U4070 (N_4070,N_1786,N_2409);
or U4071 (N_4071,N_1403,N_179);
nand U4072 (N_4072,N_22,N_2345);
xnor U4073 (N_4073,N_107,N_1806);
nor U4074 (N_4074,N_1374,N_2028);
nor U4075 (N_4075,N_1699,N_1929);
xor U4076 (N_4076,N_1138,N_1624);
nand U4077 (N_4077,N_1803,N_2178);
nor U4078 (N_4078,N_2499,N_921);
or U4079 (N_4079,N_1715,N_1296);
or U4080 (N_4080,N_582,N_2068);
nand U4081 (N_4081,N_1349,N_1212);
or U4082 (N_4082,N_309,N_1236);
nor U4083 (N_4083,N_1769,N_726);
xnor U4084 (N_4084,N_1339,N_1947);
nand U4085 (N_4085,N_117,N_1246);
nor U4086 (N_4086,N_2042,N_2339);
or U4087 (N_4087,N_1681,N_118);
xor U4088 (N_4088,N_384,N_590);
nand U4089 (N_4089,N_1522,N_1165);
or U4090 (N_4090,N_2052,N_574);
nor U4091 (N_4091,N_1301,N_1862);
or U4092 (N_4092,N_162,N_1168);
nand U4093 (N_4093,N_317,N_2249);
nor U4094 (N_4094,N_1722,N_2414);
or U4095 (N_4095,N_1935,N_1250);
and U4096 (N_4096,N_994,N_1513);
xor U4097 (N_4097,N_1981,N_2199);
and U4098 (N_4098,N_1384,N_1164);
nand U4099 (N_4099,N_673,N_1195);
and U4100 (N_4100,N_695,N_5);
nor U4101 (N_4101,N_2203,N_2257);
nor U4102 (N_4102,N_1281,N_10);
xnor U4103 (N_4103,N_1118,N_1676);
xor U4104 (N_4104,N_2066,N_2362);
nand U4105 (N_4105,N_1685,N_2307);
nand U4106 (N_4106,N_2451,N_911);
or U4107 (N_4107,N_1581,N_835);
xor U4108 (N_4108,N_75,N_403);
nor U4109 (N_4109,N_1633,N_748);
xnor U4110 (N_4110,N_1873,N_2064);
xnor U4111 (N_4111,N_1304,N_2200);
xor U4112 (N_4112,N_1540,N_51);
nand U4113 (N_4113,N_410,N_1059);
and U4114 (N_4114,N_280,N_1387);
nor U4115 (N_4115,N_673,N_1446);
or U4116 (N_4116,N_1237,N_672);
xor U4117 (N_4117,N_2195,N_716);
nand U4118 (N_4118,N_2090,N_1684);
nand U4119 (N_4119,N_699,N_1898);
nor U4120 (N_4120,N_800,N_342);
nand U4121 (N_4121,N_1474,N_597);
and U4122 (N_4122,N_1575,N_2487);
nor U4123 (N_4123,N_843,N_1375);
xnor U4124 (N_4124,N_2392,N_1947);
xnor U4125 (N_4125,N_836,N_685);
nand U4126 (N_4126,N_50,N_972);
nand U4127 (N_4127,N_1074,N_319);
xor U4128 (N_4128,N_1934,N_1259);
nand U4129 (N_4129,N_1567,N_2384);
nor U4130 (N_4130,N_1675,N_2351);
xor U4131 (N_4131,N_2421,N_1355);
xor U4132 (N_4132,N_1705,N_1479);
and U4133 (N_4133,N_2016,N_542);
xnor U4134 (N_4134,N_1921,N_1692);
xor U4135 (N_4135,N_407,N_2341);
or U4136 (N_4136,N_18,N_1776);
and U4137 (N_4137,N_1429,N_224);
and U4138 (N_4138,N_2041,N_26);
nor U4139 (N_4139,N_1788,N_2162);
and U4140 (N_4140,N_1491,N_1376);
nand U4141 (N_4141,N_2041,N_488);
xor U4142 (N_4142,N_774,N_770);
or U4143 (N_4143,N_1778,N_1811);
or U4144 (N_4144,N_1624,N_2488);
xor U4145 (N_4145,N_2111,N_433);
and U4146 (N_4146,N_497,N_2483);
or U4147 (N_4147,N_1146,N_695);
xor U4148 (N_4148,N_2422,N_1659);
and U4149 (N_4149,N_303,N_568);
nor U4150 (N_4150,N_255,N_1805);
nor U4151 (N_4151,N_1792,N_1295);
xnor U4152 (N_4152,N_404,N_298);
or U4153 (N_4153,N_731,N_1187);
nand U4154 (N_4154,N_176,N_1206);
and U4155 (N_4155,N_2307,N_1440);
xor U4156 (N_4156,N_1603,N_1481);
xor U4157 (N_4157,N_910,N_1348);
nor U4158 (N_4158,N_2051,N_1942);
or U4159 (N_4159,N_1216,N_2248);
nor U4160 (N_4160,N_2084,N_1551);
nor U4161 (N_4161,N_880,N_2122);
nand U4162 (N_4162,N_631,N_790);
xor U4163 (N_4163,N_1715,N_98);
nand U4164 (N_4164,N_2438,N_1362);
nand U4165 (N_4165,N_2025,N_1153);
xnor U4166 (N_4166,N_30,N_1);
or U4167 (N_4167,N_1872,N_571);
nand U4168 (N_4168,N_1762,N_1572);
and U4169 (N_4169,N_1946,N_1160);
xnor U4170 (N_4170,N_2406,N_1231);
nand U4171 (N_4171,N_112,N_1369);
nor U4172 (N_4172,N_280,N_534);
nand U4173 (N_4173,N_2173,N_2108);
nor U4174 (N_4174,N_1735,N_309);
nor U4175 (N_4175,N_1013,N_1397);
xnor U4176 (N_4176,N_426,N_735);
and U4177 (N_4177,N_721,N_1779);
or U4178 (N_4178,N_1758,N_1450);
nand U4179 (N_4179,N_2124,N_1467);
and U4180 (N_4180,N_1035,N_521);
nand U4181 (N_4181,N_531,N_2308);
xor U4182 (N_4182,N_1905,N_1954);
nand U4183 (N_4183,N_567,N_2347);
and U4184 (N_4184,N_1747,N_348);
xor U4185 (N_4185,N_2229,N_1844);
nor U4186 (N_4186,N_444,N_1461);
nor U4187 (N_4187,N_1222,N_2182);
and U4188 (N_4188,N_106,N_416);
xnor U4189 (N_4189,N_2000,N_2192);
and U4190 (N_4190,N_1540,N_2036);
xnor U4191 (N_4191,N_5,N_841);
nor U4192 (N_4192,N_429,N_297);
xnor U4193 (N_4193,N_1539,N_170);
xnor U4194 (N_4194,N_518,N_1207);
nor U4195 (N_4195,N_1101,N_1444);
or U4196 (N_4196,N_497,N_638);
nor U4197 (N_4197,N_2410,N_318);
and U4198 (N_4198,N_2457,N_1702);
nand U4199 (N_4199,N_447,N_1122);
or U4200 (N_4200,N_2189,N_2147);
and U4201 (N_4201,N_1535,N_445);
and U4202 (N_4202,N_2123,N_2411);
or U4203 (N_4203,N_1515,N_2090);
or U4204 (N_4204,N_2094,N_234);
or U4205 (N_4205,N_2176,N_2293);
xnor U4206 (N_4206,N_1686,N_1049);
nand U4207 (N_4207,N_832,N_2493);
or U4208 (N_4208,N_1826,N_1107);
xor U4209 (N_4209,N_1533,N_651);
and U4210 (N_4210,N_1035,N_1961);
xnor U4211 (N_4211,N_437,N_1658);
xnor U4212 (N_4212,N_175,N_2469);
nand U4213 (N_4213,N_360,N_903);
nor U4214 (N_4214,N_756,N_1523);
and U4215 (N_4215,N_2193,N_97);
and U4216 (N_4216,N_349,N_1488);
nor U4217 (N_4217,N_2260,N_1454);
nor U4218 (N_4218,N_251,N_2043);
and U4219 (N_4219,N_1931,N_1001);
and U4220 (N_4220,N_1805,N_183);
or U4221 (N_4221,N_1506,N_1414);
nor U4222 (N_4222,N_586,N_362);
and U4223 (N_4223,N_500,N_828);
xnor U4224 (N_4224,N_2463,N_997);
xnor U4225 (N_4225,N_1299,N_1366);
nand U4226 (N_4226,N_2277,N_23);
and U4227 (N_4227,N_141,N_2496);
nor U4228 (N_4228,N_122,N_1015);
nor U4229 (N_4229,N_2428,N_1016);
nand U4230 (N_4230,N_146,N_2457);
and U4231 (N_4231,N_1282,N_1907);
nand U4232 (N_4232,N_951,N_2420);
and U4233 (N_4233,N_1877,N_160);
or U4234 (N_4234,N_707,N_654);
or U4235 (N_4235,N_647,N_2262);
nor U4236 (N_4236,N_1724,N_431);
and U4237 (N_4237,N_1017,N_2460);
nor U4238 (N_4238,N_390,N_1443);
and U4239 (N_4239,N_2279,N_308);
or U4240 (N_4240,N_521,N_614);
and U4241 (N_4241,N_777,N_681);
nand U4242 (N_4242,N_2439,N_128);
or U4243 (N_4243,N_1272,N_385);
or U4244 (N_4244,N_214,N_1958);
nand U4245 (N_4245,N_2243,N_2391);
xor U4246 (N_4246,N_1898,N_484);
nor U4247 (N_4247,N_1185,N_2264);
nand U4248 (N_4248,N_2388,N_2140);
xor U4249 (N_4249,N_2163,N_2239);
xnor U4250 (N_4250,N_1692,N_2018);
and U4251 (N_4251,N_1957,N_1035);
xnor U4252 (N_4252,N_929,N_1460);
or U4253 (N_4253,N_1955,N_902);
xor U4254 (N_4254,N_513,N_2411);
nor U4255 (N_4255,N_2471,N_795);
or U4256 (N_4256,N_1857,N_1436);
nor U4257 (N_4257,N_774,N_1086);
nand U4258 (N_4258,N_1459,N_1433);
nor U4259 (N_4259,N_1480,N_1645);
xnor U4260 (N_4260,N_1240,N_1794);
nand U4261 (N_4261,N_647,N_1871);
nand U4262 (N_4262,N_1294,N_1367);
or U4263 (N_4263,N_1579,N_159);
xor U4264 (N_4264,N_1686,N_664);
xnor U4265 (N_4265,N_1264,N_1424);
or U4266 (N_4266,N_1780,N_184);
nor U4267 (N_4267,N_350,N_1292);
nor U4268 (N_4268,N_793,N_498);
and U4269 (N_4269,N_310,N_164);
nand U4270 (N_4270,N_1004,N_1309);
nand U4271 (N_4271,N_2192,N_2498);
nand U4272 (N_4272,N_2276,N_997);
or U4273 (N_4273,N_1486,N_2218);
xnor U4274 (N_4274,N_1480,N_1433);
and U4275 (N_4275,N_1495,N_1515);
xor U4276 (N_4276,N_598,N_574);
nor U4277 (N_4277,N_1537,N_1251);
nor U4278 (N_4278,N_2121,N_1143);
nand U4279 (N_4279,N_634,N_1628);
xor U4280 (N_4280,N_1090,N_876);
xor U4281 (N_4281,N_2231,N_543);
xor U4282 (N_4282,N_2128,N_95);
nor U4283 (N_4283,N_1648,N_2046);
nor U4284 (N_4284,N_1090,N_805);
nor U4285 (N_4285,N_1221,N_862);
and U4286 (N_4286,N_458,N_1482);
and U4287 (N_4287,N_882,N_517);
xor U4288 (N_4288,N_1264,N_98);
nand U4289 (N_4289,N_504,N_1090);
nor U4290 (N_4290,N_1492,N_801);
nand U4291 (N_4291,N_2173,N_1863);
and U4292 (N_4292,N_502,N_1526);
or U4293 (N_4293,N_1619,N_14);
and U4294 (N_4294,N_438,N_1933);
and U4295 (N_4295,N_1968,N_231);
nor U4296 (N_4296,N_1706,N_1436);
xor U4297 (N_4297,N_2466,N_1325);
nand U4298 (N_4298,N_929,N_1218);
nor U4299 (N_4299,N_758,N_945);
nand U4300 (N_4300,N_1859,N_489);
and U4301 (N_4301,N_294,N_2187);
nand U4302 (N_4302,N_180,N_1593);
nand U4303 (N_4303,N_1312,N_140);
or U4304 (N_4304,N_112,N_629);
nand U4305 (N_4305,N_1322,N_1641);
nor U4306 (N_4306,N_787,N_1456);
or U4307 (N_4307,N_213,N_2313);
or U4308 (N_4308,N_267,N_540);
nand U4309 (N_4309,N_2034,N_1360);
or U4310 (N_4310,N_585,N_2097);
nand U4311 (N_4311,N_1781,N_818);
nor U4312 (N_4312,N_684,N_2011);
nand U4313 (N_4313,N_2341,N_817);
xor U4314 (N_4314,N_115,N_2087);
or U4315 (N_4315,N_1724,N_1759);
and U4316 (N_4316,N_767,N_1052);
nand U4317 (N_4317,N_628,N_82);
xnor U4318 (N_4318,N_142,N_1670);
or U4319 (N_4319,N_691,N_628);
nor U4320 (N_4320,N_105,N_1517);
or U4321 (N_4321,N_821,N_1802);
and U4322 (N_4322,N_544,N_2037);
xnor U4323 (N_4323,N_640,N_1243);
xnor U4324 (N_4324,N_324,N_957);
xnor U4325 (N_4325,N_2435,N_1623);
and U4326 (N_4326,N_1152,N_343);
nor U4327 (N_4327,N_652,N_1930);
and U4328 (N_4328,N_535,N_1108);
or U4329 (N_4329,N_1694,N_111);
xnor U4330 (N_4330,N_447,N_2139);
nand U4331 (N_4331,N_1124,N_1807);
nand U4332 (N_4332,N_1905,N_1756);
nor U4333 (N_4333,N_1981,N_195);
nor U4334 (N_4334,N_129,N_1741);
nand U4335 (N_4335,N_424,N_2205);
nor U4336 (N_4336,N_1999,N_1225);
and U4337 (N_4337,N_2069,N_2137);
nor U4338 (N_4338,N_1996,N_909);
and U4339 (N_4339,N_1667,N_861);
or U4340 (N_4340,N_1547,N_2181);
and U4341 (N_4341,N_1829,N_1373);
nor U4342 (N_4342,N_2052,N_1100);
nor U4343 (N_4343,N_812,N_325);
or U4344 (N_4344,N_148,N_177);
or U4345 (N_4345,N_278,N_1272);
or U4346 (N_4346,N_192,N_1797);
xor U4347 (N_4347,N_2170,N_347);
or U4348 (N_4348,N_51,N_1595);
xnor U4349 (N_4349,N_1562,N_92);
or U4350 (N_4350,N_1299,N_51);
or U4351 (N_4351,N_954,N_1574);
or U4352 (N_4352,N_422,N_2456);
nand U4353 (N_4353,N_357,N_2410);
and U4354 (N_4354,N_557,N_266);
nor U4355 (N_4355,N_1809,N_1040);
and U4356 (N_4356,N_429,N_544);
nor U4357 (N_4357,N_1051,N_1478);
nor U4358 (N_4358,N_2350,N_1193);
nor U4359 (N_4359,N_1441,N_1249);
nor U4360 (N_4360,N_1609,N_1639);
nor U4361 (N_4361,N_480,N_1558);
nand U4362 (N_4362,N_2326,N_935);
nor U4363 (N_4363,N_11,N_2072);
and U4364 (N_4364,N_2143,N_2473);
or U4365 (N_4365,N_284,N_478);
or U4366 (N_4366,N_1744,N_657);
or U4367 (N_4367,N_488,N_561);
xor U4368 (N_4368,N_1427,N_1649);
nand U4369 (N_4369,N_2340,N_179);
and U4370 (N_4370,N_2458,N_1073);
or U4371 (N_4371,N_380,N_452);
or U4372 (N_4372,N_2370,N_362);
xor U4373 (N_4373,N_1556,N_900);
nor U4374 (N_4374,N_610,N_1060);
xnor U4375 (N_4375,N_1559,N_2418);
and U4376 (N_4376,N_1578,N_1603);
nor U4377 (N_4377,N_146,N_2267);
nor U4378 (N_4378,N_825,N_2026);
xnor U4379 (N_4379,N_2202,N_1582);
nand U4380 (N_4380,N_1480,N_2076);
or U4381 (N_4381,N_325,N_666);
nor U4382 (N_4382,N_2360,N_2444);
nand U4383 (N_4383,N_2302,N_771);
or U4384 (N_4384,N_1842,N_118);
and U4385 (N_4385,N_2083,N_283);
nor U4386 (N_4386,N_362,N_519);
or U4387 (N_4387,N_1466,N_2440);
xor U4388 (N_4388,N_1585,N_1000);
nor U4389 (N_4389,N_2343,N_2375);
xnor U4390 (N_4390,N_1212,N_766);
and U4391 (N_4391,N_368,N_1921);
xnor U4392 (N_4392,N_1411,N_2328);
or U4393 (N_4393,N_1171,N_7);
nand U4394 (N_4394,N_2116,N_1007);
xnor U4395 (N_4395,N_1860,N_1400);
xor U4396 (N_4396,N_775,N_951);
or U4397 (N_4397,N_1240,N_1265);
xnor U4398 (N_4398,N_1960,N_1955);
nor U4399 (N_4399,N_467,N_464);
and U4400 (N_4400,N_973,N_1158);
nor U4401 (N_4401,N_2299,N_2039);
nor U4402 (N_4402,N_1484,N_1816);
nor U4403 (N_4403,N_1583,N_1985);
xor U4404 (N_4404,N_811,N_1991);
xnor U4405 (N_4405,N_999,N_702);
or U4406 (N_4406,N_1139,N_1097);
nor U4407 (N_4407,N_1001,N_972);
and U4408 (N_4408,N_1843,N_409);
or U4409 (N_4409,N_86,N_414);
and U4410 (N_4410,N_2371,N_1638);
nor U4411 (N_4411,N_64,N_1914);
or U4412 (N_4412,N_701,N_153);
and U4413 (N_4413,N_1419,N_405);
or U4414 (N_4414,N_13,N_1634);
and U4415 (N_4415,N_807,N_551);
nand U4416 (N_4416,N_125,N_1542);
xor U4417 (N_4417,N_929,N_414);
xnor U4418 (N_4418,N_390,N_1782);
and U4419 (N_4419,N_2204,N_943);
xnor U4420 (N_4420,N_2026,N_1642);
nor U4421 (N_4421,N_395,N_439);
nand U4422 (N_4422,N_525,N_1935);
and U4423 (N_4423,N_173,N_1528);
nor U4424 (N_4424,N_2437,N_1036);
nand U4425 (N_4425,N_50,N_2484);
xor U4426 (N_4426,N_2269,N_2472);
or U4427 (N_4427,N_2206,N_1405);
and U4428 (N_4428,N_740,N_1044);
and U4429 (N_4429,N_599,N_2433);
nor U4430 (N_4430,N_1357,N_2301);
xnor U4431 (N_4431,N_1913,N_72);
nor U4432 (N_4432,N_1651,N_1462);
xnor U4433 (N_4433,N_1417,N_2450);
or U4434 (N_4434,N_605,N_1579);
or U4435 (N_4435,N_1890,N_901);
and U4436 (N_4436,N_1837,N_462);
nand U4437 (N_4437,N_1030,N_564);
and U4438 (N_4438,N_133,N_130);
nand U4439 (N_4439,N_1291,N_1305);
xnor U4440 (N_4440,N_1039,N_405);
or U4441 (N_4441,N_19,N_1313);
and U4442 (N_4442,N_256,N_1516);
nand U4443 (N_4443,N_666,N_155);
nand U4444 (N_4444,N_1529,N_1927);
or U4445 (N_4445,N_728,N_1587);
and U4446 (N_4446,N_1493,N_1174);
nor U4447 (N_4447,N_74,N_1566);
nor U4448 (N_4448,N_142,N_398);
or U4449 (N_4449,N_374,N_884);
xor U4450 (N_4450,N_941,N_1978);
xor U4451 (N_4451,N_1237,N_795);
nand U4452 (N_4452,N_2462,N_752);
nand U4453 (N_4453,N_219,N_842);
or U4454 (N_4454,N_1174,N_1714);
and U4455 (N_4455,N_595,N_2319);
xor U4456 (N_4456,N_1304,N_2486);
nand U4457 (N_4457,N_1768,N_1270);
xor U4458 (N_4458,N_1545,N_2026);
nand U4459 (N_4459,N_1544,N_1213);
nor U4460 (N_4460,N_256,N_1636);
nand U4461 (N_4461,N_1973,N_1989);
and U4462 (N_4462,N_1734,N_386);
nor U4463 (N_4463,N_304,N_491);
nor U4464 (N_4464,N_1029,N_996);
and U4465 (N_4465,N_2064,N_1703);
nand U4466 (N_4466,N_1762,N_973);
or U4467 (N_4467,N_1092,N_954);
nor U4468 (N_4468,N_1532,N_2345);
xor U4469 (N_4469,N_167,N_2004);
or U4470 (N_4470,N_1755,N_1612);
and U4471 (N_4471,N_2134,N_1365);
and U4472 (N_4472,N_1568,N_2403);
xnor U4473 (N_4473,N_1204,N_1249);
and U4474 (N_4474,N_521,N_1796);
nor U4475 (N_4475,N_900,N_1115);
and U4476 (N_4476,N_2105,N_922);
nor U4477 (N_4477,N_1757,N_1957);
nand U4478 (N_4478,N_1865,N_169);
xnor U4479 (N_4479,N_651,N_1168);
nor U4480 (N_4480,N_2225,N_1282);
nand U4481 (N_4481,N_82,N_269);
and U4482 (N_4482,N_2232,N_299);
and U4483 (N_4483,N_218,N_970);
nand U4484 (N_4484,N_1071,N_2271);
xnor U4485 (N_4485,N_639,N_1628);
and U4486 (N_4486,N_1461,N_2301);
nor U4487 (N_4487,N_2360,N_538);
and U4488 (N_4488,N_705,N_1);
xnor U4489 (N_4489,N_1907,N_156);
xnor U4490 (N_4490,N_913,N_481);
xnor U4491 (N_4491,N_1121,N_114);
nand U4492 (N_4492,N_2148,N_1432);
xor U4493 (N_4493,N_91,N_884);
xnor U4494 (N_4494,N_338,N_1761);
xor U4495 (N_4495,N_835,N_549);
xor U4496 (N_4496,N_2054,N_2034);
and U4497 (N_4497,N_2349,N_2267);
nor U4498 (N_4498,N_1669,N_1072);
nand U4499 (N_4499,N_2296,N_522);
nor U4500 (N_4500,N_1039,N_1633);
or U4501 (N_4501,N_1565,N_1228);
xor U4502 (N_4502,N_2175,N_293);
nand U4503 (N_4503,N_407,N_929);
or U4504 (N_4504,N_1362,N_1942);
xnor U4505 (N_4505,N_1724,N_190);
nor U4506 (N_4506,N_1056,N_1101);
and U4507 (N_4507,N_1185,N_1186);
and U4508 (N_4508,N_1754,N_1082);
nor U4509 (N_4509,N_1767,N_1231);
xor U4510 (N_4510,N_1495,N_333);
and U4511 (N_4511,N_2376,N_180);
or U4512 (N_4512,N_174,N_1228);
or U4513 (N_4513,N_1822,N_402);
xnor U4514 (N_4514,N_555,N_416);
nand U4515 (N_4515,N_2082,N_1409);
or U4516 (N_4516,N_880,N_923);
nand U4517 (N_4517,N_2413,N_1751);
and U4518 (N_4518,N_2466,N_292);
nand U4519 (N_4519,N_275,N_393);
and U4520 (N_4520,N_1338,N_1897);
nor U4521 (N_4521,N_982,N_816);
and U4522 (N_4522,N_1813,N_1881);
or U4523 (N_4523,N_2457,N_698);
and U4524 (N_4524,N_1305,N_2148);
and U4525 (N_4525,N_1918,N_200);
nand U4526 (N_4526,N_923,N_668);
or U4527 (N_4527,N_1764,N_297);
or U4528 (N_4528,N_1155,N_2089);
xnor U4529 (N_4529,N_553,N_447);
or U4530 (N_4530,N_2035,N_1795);
nor U4531 (N_4531,N_1453,N_736);
and U4532 (N_4532,N_645,N_402);
nor U4533 (N_4533,N_628,N_2066);
or U4534 (N_4534,N_878,N_1122);
nor U4535 (N_4535,N_1036,N_856);
xor U4536 (N_4536,N_1476,N_1271);
nand U4537 (N_4537,N_2373,N_307);
xnor U4538 (N_4538,N_128,N_2282);
or U4539 (N_4539,N_264,N_2039);
and U4540 (N_4540,N_897,N_1988);
nand U4541 (N_4541,N_2499,N_580);
nand U4542 (N_4542,N_1277,N_537);
nor U4543 (N_4543,N_2223,N_2194);
or U4544 (N_4544,N_2309,N_1077);
and U4545 (N_4545,N_1501,N_1268);
nor U4546 (N_4546,N_1271,N_1714);
nand U4547 (N_4547,N_1387,N_297);
xnor U4548 (N_4548,N_1410,N_1619);
or U4549 (N_4549,N_1883,N_307);
and U4550 (N_4550,N_460,N_1051);
nand U4551 (N_4551,N_794,N_1803);
nand U4552 (N_4552,N_757,N_2035);
nor U4553 (N_4553,N_274,N_670);
xor U4554 (N_4554,N_1943,N_2328);
and U4555 (N_4555,N_1805,N_629);
nor U4556 (N_4556,N_1376,N_242);
nand U4557 (N_4557,N_1688,N_2028);
and U4558 (N_4558,N_309,N_471);
nor U4559 (N_4559,N_1085,N_1270);
or U4560 (N_4560,N_2074,N_132);
nand U4561 (N_4561,N_1610,N_159);
nor U4562 (N_4562,N_1202,N_1539);
xor U4563 (N_4563,N_985,N_1487);
and U4564 (N_4564,N_1696,N_1142);
nor U4565 (N_4565,N_656,N_23);
or U4566 (N_4566,N_192,N_1252);
or U4567 (N_4567,N_953,N_848);
xor U4568 (N_4568,N_173,N_1295);
xnor U4569 (N_4569,N_166,N_1427);
nor U4570 (N_4570,N_885,N_1510);
or U4571 (N_4571,N_1533,N_2080);
nor U4572 (N_4572,N_1728,N_2087);
and U4573 (N_4573,N_1659,N_1071);
and U4574 (N_4574,N_2453,N_2046);
or U4575 (N_4575,N_164,N_1578);
xor U4576 (N_4576,N_1111,N_861);
nor U4577 (N_4577,N_2163,N_193);
nand U4578 (N_4578,N_1660,N_571);
nor U4579 (N_4579,N_1692,N_1254);
and U4580 (N_4580,N_2331,N_681);
nand U4581 (N_4581,N_310,N_1203);
or U4582 (N_4582,N_925,N_765);
nor U4583 (N_4583,N_597,N_1498);
nand U4584 (N_4584,N_1369,N_78);
or U4585 (N_4585,N_211,N_2035);
nand U4586 (N_4586,N_2299,N_1902);
and U4587 (N_4587,N_564,N_2184);
nand U4588 (N_4588,N_909,N_188);
and U4589 (N_4589,N_1555,N_371);
nor U4590 (N_4590,N_962,N_386);
and U4591 (N_4591,N_102,N_522);
xnor U4592 (N_4592,N_2097,N_409);
and U4593 (N_4593,N_613,N_1360);
nand U4594 (N_4594,N_2101,N_284);
nand U4595 (N_4595,N_555,N_1627);
xor U4596 (N_4596,N_1546,N_1466);
and U4597 (N_4597,N_1990,N_1040);
or U4598 (N_4598,N_813,N_2041);
nand U4599 (N_4599,N_775,N_1849);
nor U4600 (N_4600,N_1816,N_23);
and U4601 (N_4601,N_243,N_396);
nor U4602 (N_4602,N_1429,N_879);
xor U4603 (N_4603,N_1822,N_1313);
and U4604 (N_4604,N_2248,N_12);
nand U4605 (N_4605,N_1011,N_1196);
xnor U4606 (N_4606,N_1179,N_1043);
and U4607 (N_4607,N_2008,N_1548);
or U4608 (N_4608,N_610,N_2098);
or U4609 (N_4609,N_1115,N_2442);
nor U4610 (N_4610,N_1380,N_1395);
nand U4611 (N_4611,N_2243,N_77);
nand U4612 (N_4612,N_2138,N_611);
or U4613 (N_4613,N_1943,N_1743);
xnor U4614 (N_4614,N_828,N_1541);
or U4615 (N_4615,N_1604,N_777);
and U4616 (N_4616,N_1163,N_1481);
and U4617 (N_4617,N_1347,N_1934);
and U4618 (N_4618,N_2148,N_1375);
and U4619 (N_4619,N_715,N_2184);
and U4620 (N_4620,N_2138,N_2445);
and U4621 (N_4621,N_1213,N_2133);
nor U4622 (N_4622,N_2220,N_711);
or U4623 (N_4623,N_766,N_1707);
and U4624 (N_4624,N_2134,N_912);
and U4625 (N_4625,N_35,N_30);
nand U4626 (N_4626,N_583,N_81);
or U4627 (N_4627,N_1937,N_1672);
and U4628 (N_4628,N_509,N_1375);
nor U4629 (N_4629,N_1924,N_1498);
and U4630 (N_4630,N_1789,N_329);
nor U4631 (N_4631,N_2448,N_305);
nand U4632 (N_4632,N_2235,N_1713);
nand U4633 (N_4633,N_596,N_1116);
nand U4634 (N_4634,N_763,N_251);
xor U4635 (N_4635,N_674,N_6);
and U4636 (N_4636,N_2169,N_2245);
nor U4637 (N_4637,N_1444,N_108);
or U4638 (N_4638,N_249,N_455);
nand U4639 (N_4639,N_194,N_1794);
nand U4640 (N_4640,N_348,N_939);
nand U4641 (N_4641,N_2268,N_222);
xor U4642 (N_4642,N_1748,N_1223);
nor U4643 (N_4643,N_888,N_382);
nand U4644 (N_4644,N_2135,N_332);
or U4645 (N_4645,N_549,N_111);
nand U4646 (N_4646,N_92,N_2479);
or U4647 (N_4647,N_724,N_1649);
xnor U4648 (N_4648,N_105,N_576);
nor U4649 (N_4649,N_2206,N_841);
nand U4650 (N_4650,N_2155,N_273);
and U4651 (N_4651,N_1581,N_546);
and U4652 (N_4652,N_2382,N_301);
nand U4653 (N_4653,N_1253,N_853);
or U4654 (N_4654,N_1898,N_2226);
nand U4655 (N_4655,N_563,N_582);
nand U4656 (N_4656,N_615,N_1865);
or U4657 (N_4657,N_2480,N_316);
xor U4658 (N_4658,N_369,N_1312);
nor U4659 (N_4659,N_2348,N_1199);
or U4660 (N_4660,N_1340,N_691);
and U4661 (N_4661,N_1995,N_82);
or U4662 (N_4662,N_216,N_1523);
nor U4663 (N_4663,N_1261,N_2257);
or U4664 (N_4664,N_58,N_1926);
nand U4665 (N_4665,N_1580,N_1696);
nor U4666 (N_4666,N_215,N_1356);
xnor U4667 (N_4667,N_147,N_2238);
nand U4668 (N_4668,N_907,N_2471);
and U4669 (N_4669,N_444,N_172);
or U4670 (N_4670,N_1787,N_1674);
or U4671 (N_4671,N_1111,N_1713);
nand U4672 (N_4672,N_47,N_1143);
nor U4673 (N_4673,N_1344,N_630);
nor U4674 (N_4674,N_1671,N_472);
and U4675 (N_4675,N_1338,N_1564);
and U4676 (N_4676,N_2434,N_719);
xnor U4677 (N_4677,N_1530,N_1870);
or U4678 (N_4678,N_284,N_427);
nor U4679 (N_4679,N_1572,N_1677);
and U4680 (N_4680,N_213,N_1925);
xnor U4681 (N_4681,N_943,N_2032);
and U4682 (N_4682,N_1153,N_1740);
nand U4683 (N_4683,N_2282,N_1295);
and U4684 (N_4684,N_2309,N_231);
nand U4685 (N_4685,N_1116,N_1499);
and U4686 (N_4686,N_827,N_1600);
nand U4687 (N_4687,N_1741,N_760);
nand U4688 (N_4688,N_1275,N_255);
nand U4689 (N_4689,N_297,N_1311);
nor U4690 (N_4690,N_846,N_824);
nor U4691 (N_4691,N_1098,N_2314);
xnor U4692 (N_4692,N_2067,N_171);
and U4693 (N_4693,N_1230,N_2312);
or U4694 (N_4694,N_1771,N_1514);
xnor U4695 (N_4695,N_876,N_2067);
nor U4696 (N_4696,N_101,N_1778);
nor U4697 (N_4697,N_1506,N_393);
xor U4698 (N_4698,N_645,N_2499);
nand U4699 (N_4699,N_634,N_740);
nor U4700 (N_4700,N_121,N_1133);
nand U4701 (N_4701,N_327,N_1038);
nor U4702 (N_4702,N_266,N_146);
xor U4703 (N_4703,N_2189,N_1300);
and U4704 (N_4704,N_2423,N_300);
or U4705 (N_4705,N_2029,N_257);
and U4706 (N_4706,N_880,N_969);
or U4707 (N_4707,N_532,N_1283);
xor U4708 (N_4708,N_2442,N_1118);
or U4709 (N_4709,N_2170,N_1075);
xor U4710 (N_4710,N_252,N_341);
nand U4711 (N_4711,N_189,N_1762);
nand U4712 (N_4712,N_1863,N_3);
or U4713 (N_4713,N_1619,N_1393);
nand U4714 (N_4714,N_864,N_1005);
and U4715 (N_4715,N_298,N_1726);
and U4716 (N_4716,N_463,N_1077);
xnor U4717 (N_4717,N_2338,N_335);
nor U4718 (N_4718,N_420,N_828);
nor U4719 (N_4719,N_763,N_25);
and U4720 (N_4720,N_232,N_56);
or U4721 (N_4721,N_2316,N_718);
or U4722 (N_4722,N_669,N_2403);
and U4723 (N_4723,N_1191,N_2300);
and U4724 (N_4724,N_651,N_945);
nand U4725 (N_4725,N_1220,N_2467);
nand U4726 (N_4726,N_1171,N_1221);
and U4727 (N_4727,N_604,N_543);
and U4728 (N_4728,N_1844,N_274);
nand U4729 (N_4729,N_352,N_103);
and U4730 (N_4730,N_1213,N_389);
and U4731 (N_4731,N_153,N_1642);
nor U4732 (N_4732,N_407,N_2281);
or U4733 (N_4733,N_1979,N_939);
and U4734 (N_4734,N_731,N_1527);
xnor U4735 (N_4735,N_1249,N_490);
xnor U4736 (N_4736,N_1445,N_1888);
nor U4737 (N_4737,N_541,N_2477);
nor U4738 (N_4738,N_40,N_2297);
nor U4739 (N_4739,N_2437,N_1955);
and U4740 (N_4740,N_1558,N_622);
xor U4741 (N_4741,N_1497,N_1935);
or U4742 (N_4742,N_326,N_1861);
or U4743 (N_4743,N_483,N_835);
nand U4744 (N_4744,N_2352,N_1901);
and U4745 (N_4745,N_1719,N_726);
or U4746 (N_4746,N_1041,N_1107);
or U4747 (N_4747,N_921,N_444);
xor U4748 (N_4748,N_1464,N_1337);
nor U4749 (N_4749,N_2027,N_1429);
xnor U4750 (N_4750,N_2178,N_837);
xnor U4751 (N_4751,N_607,N_119);
nor U4752 (N_4752,N_1549,N_862);
xnor U4753 (N_4753,N_1185,N_890);
nand U4754 (N_4754,N_2152,N_1325);
or U4755 (N_4755,N_777,N_2305);
nand U4756 (N_4756,N_2474,N_1837);
or U4757 (N_4757,N_662,N_649);
or U4758 (N_4758,N_486,N_1415);
or U4759 (N_4759,N_362,N_445);
and U4760 (N_4760,N_323,N_426);
or U4761 (N_4761,N_46,N_757);
nand U4762 (N_4762,N_1293,N_2465);
nand U4763 (N_4763,N_245,N_306);
and U4764 (N_4764,N_900,N_254);
nor U4765 (N_4765,N_1534,N_2419);
nor U4766 (N_4766,N_1241,N_50);
nor U4767 (N_4767,N_1457,N_1224);
nor U4768 (N_4768,N_1345,N_140);
xor U4769 (N_4769,N_1651,N_618);
xnor U4770 (N_4770,N_2030,N_495);
nor U4771 (N_4771,N_2334,N_416);
and U4772 (N_4772,N_1384,N_43);
and U4773 (N_4773,N_1535,N_407);
nand U4774 (N_4774,N_806,N_730);
nand U4775 (N_4775,N_2322,N_307);
or U4776 (N_4776,N_1173,N_2139);
nor U4777 (N_4777,N_502,N_2330);
and U4778 (N_4778,N_818,N_773);
nor U4779 (N_4779,N_2212,N_1584);
and U4780 (N_4780,N_1769,N_874);
nor U4781 (N_4781,N_462,N_1987);
and U4782 (N_4782,N_13,N_1308);
xor U4783 (N_4783,N_1765,N_911);
nand U4784 (N_4784,N_510,N_519);
and U4785 (N_4785,N_1617,N_319);
xor U4786 (N_4786,N_1676,N_493);
nor U4787 (N_4787,N_2215,N_1572);
nor U4788 (N_4788,N_1414,N_2467);
nor U4789 (N_4789,N_2421,N_1274);
and U4790 (N_4790,N_1049,N_904);
xnor U4791 (N_4791,N_1177,N_796);
xnor U4792 (N_4792,N_1683,N_309);
nand U4793 (N_4793,N_186,N_2199);
nand U4794 (N_4794,N_1853,N_56);
nand U4795 (N_4795,N_1918,N_1528);
and U4796 (N_4796,N_741,N_1512);
nand U4797 (N_4797,N_2272,N_1002);
nand U4798 (N_4798,N_2416,N_192);
or U4799 (N_4799,N_753,N_2415);
nand U4800 (N_4800,N_80,N_183);
nor U4801 (N_4801,N_479,N_723);
and U4802 (N_4802,N_1830,N_548);
and U4803 (N_4803,N_1747,N_1603);
or U4804 (N_4804,N_1899,N_1589);
nand U4805 (N_4805,N_2174,N_86);
nand U4806 (N_4806,N_322,N_20);
xnor U4807 (N_4807,N_45,N_450);
nor U4808 (N_4808,N_1389,N_1682);
or U4809 (N_4809,N_2322,N_516);
nor U4810 (N_4810,N_1377,N_235);
nor U4811 (N_4811,N_1671,N_593);
nand U4812 (N_4812,N_2285,N_589);
nor U4813 (N_4813,N_1255,N_551);
nor U4814 (N_4814,N_442,N_2466);
or U4815 (N_4815,N_2240,N_594);
and U4816 (N_4816,N_655,N_1430);
and U4817 (N_4817,N_1826,N_1447);
or U4818 (N_4818,N_1066,N_839);
xor U4819 (N_4819,N_1385,N_418);
nand U4820 (N_4820,N_985,N_1744);
and U4821 (N_4821,N_67,N_839);
nor U4822 (N_4822,N_1620,N_1288);
nor U4823 (N_4823,N_1465,N_1933);
xnor U4824 (N_4824,N_1334,N_230);
nand U4825 (N_4825,N_456,N_1743);
nor U4826 (N_4826,N_70,N_1466);
nor U4827 (N_4827,N_1142,N_1329);
nor U4828 (N_4828,N_1981,N_1419);
and U4829 (N_4829,N_970,N_676);
nor U4830 (N_4830,N_1324,N_980);
and U4831 (N_4831,N_1152,N_945);
xnor U4832 (N_4832,N_1513,N_1282);
nor U4833 (N_4833,N_1410,N_798);
nand U4834 (N_4834,N_1066,N_1982);
nand U4835 (N_4835,N_2094,N_254);
nand U4836 (N_4836,N_385,N_327);
xnor U4837 (N_4837,N_1237,N_1276);
nor U4838 (N_4838,N_894,N_185);
nor U4839 (N_4839,N_49,N_1244);
or U4840 (N_4840,N_2168,N_1398);
nand U4841 (N_4841,N_633,N_1235);
nand U4842 (N_4842,N_458,N_1287);
xnor U4843 (N_4843,N_540,N_1068);
nand U4844 (N_4844,N_1968,N_1164);
xor U4845 (N_4845,N_297,N_1080);
nand U4846 (N_4846,N_493,N_31);
xnor U4847 (N_4847,N_2495,N_1318);
or U4848 (N_4848,N_1305,N_1203);
nor U4849 (N_4849,N_1566,N_423);
or U4850 (N_4850,N_193,N_1903);
and U4851 (N_4851,N_1124,N_804);
nand U4852 (N_4852,N_1620,N_1284);
nor U4853 (N_4853,N_312,N_1740);
nand U4854 (N_4854,N_966,N_672);
or U4855 (N_4855,N_2495,N_2015);
xnor U4856 (N_4856,N_2136,N_1300);
nand U4857 (N_4857,N_1480,N_2183);
and U4858 (N_4858,N_213,N_1297);
or U4859 (N_4859,N_1121,N_446);
and U4860 (N_4860,N_1442,N_2376);
nand U4861 (N_4861,N_323,N_1862);
nand U4862 (N_4862,N_718,N_879);
nor U4863 (N_4863,N_1352,N_2218);
and U4864 (N_4864,N_1603,N_957);
nor U4865 (N_4865,N_720,N_2116);
nand U4866 (N_4866,N_1562,N_817);
nor U4867 (N_4867,N_1779,N_1403);
or U4868 (N_4868,N_1846,N_598);
or U4869 (N_4869,N_1795,N_1375);
xor U4870 (N_4870,N_1711,N_1923);
xnor U4871 (N_4871,N_755,N_2209);
or U4872 (N_4872,N_186,N_771);
nor U4873 (N_4873,N_273,N_2338);
nand U4874 (N_4874,N_2482,N_1557);
nand U4875 (N_4875,N_67,N_2028);
xnor U4876 (N_4876,N_531,N_580);
xor U4877 (N_4877,N_2446,N_2376);
and U4878 (N_4878,N_2457,N_1534);
nor U4879 (N_4879,N_157,N_37);
xnor U4880 (N_4880,N_1296,N_1837);
nand U4881 (N_4881,N_2024,N_471);
nand U4882 (N_4882,N_671,N_1088);
or U4883 (N_4883,N_1906,N_705);
xnor U4884 (N_4884,N_1551,N_1632);
or U4885 (N_4885,N_1580,N_1024);
nor U4886 (N_4886,N_390,N_1119);
nand U4887 (N_4887,N_1632,N_83);
nand U4888 (N_4888,N_288,N_1576);
and U4889 (N_4889,N_2053,N_1297);
or U4890 (N_4890,N_548,N_1631);
nand U4891 (N_4891,N_758,N_1409);
or U4892 (N_4892,N_1409,N_1999);
nand U4893 (N_4893,N_1653,N_208);
nor U4894 (N_4894,N_1178,N_2403);
xor U4895 (N_4895,N_256,N_2348);
and U4896 (N_4896,N_992,N_1156);
nor U4897 (N_4897,N_2190,N_1582);
nor U4898 (N_4898,N_736,N_775);
nand U4899 (N_4899,N_213,N_2108);
xor U4900 (N_4900,N_1642,N_1244);
xor U4901 (N_4901,N_2180,N_902);
or U4902 (N_4902,N_1874,N_456);
nor U4903 (N_4903,N_1994,N_2011);
and U4904 (N_4904,N_149,N_779);
and U4905 (N_4905,N_1886,N_1558);
xnor U4906 (N_4906,N_2039,N_263);
xnor U4907 (N_4907,N_2153,N_220);
xnor U4908 (N_4908,N_1939,N_420);
xnor U4909 (N_4909,N_478,N_1326);
nand U4910 (N_4910,N_2157,N_2338);
or U4911 (N_4911,N_2172,N_1524);
xnor U4912 (N_4912,N_795,N_984);
nand U4913 (N_4913,N_649,N_1936);
xor U4914 (N_4914,N_449,N_1886);
nand U4915 (N_4915,N_1899,N_545);
nand U4916 (N_4916,N_2069,N_565);
or U4917 (N_4917,N_910,N_782);
or U4918 (N_4918,N_836,N_863);
and U4919 (N_4919,N_304,N_1226);
or U4920 (N_4920,N_1949,N_1453);
and U4921 (N_4921,N_132,N_296);
nor U4922 (N_4922,N_1352,N_1720);
xnor U4923 (N_4923,N_2285,N_1464);
xor U4924 (N_4924,N_1362,N_711);
xnor U4925 (N_4925,N_1402,N_1091);
or U4926 (N_4926,N_951,N_901);
nand U4927 (N_4927,N_1247,N_1090);
or U4928 (N_4928,N_351,N_1792);
or U4929 (N_4929,N_1055,N_1536);
xor U4930 (N_4930,N_1386,N_1959);
nor U4931 (N_4931,N_1519,N_92);
and U4932 (N_4932,N_2498,N_553);
and U4933 (N_4933,N_1340,N_579);
and U4934 (N_4934,N_497,N_2009);
and U4935 (N_4935,N_1940,N_1292);
nand U4936 (N_4936,N_1185,N_1912);
and U4937 (N_4937,N_638,N_631);
nor U4938 (N_4938,N_2316,N_2419);
nand U4939 (N_4939,N_1212,N_2292);
and U4940 (N_4940,N_34,N_407);
xor U4941 (N_4941,N_1740,N_926);
or U4942 (N_4942,N_1867,N_2198);
nor U4943 (N_4943,N_2096,N_569);
nor U4944 (N_4944,N_413,N_2274);
xnor U4945 (N_4945,N_1295,N_508);
nor U4946 (N_4946,N_2335,N_685);
and U4947 (N_4947,N_1033,N_2449);
or U4948 (N_4948,N_1910,N_1707);
xor U4949 (N_4949,N_366,N_826);
or U4950 (N_4950,N_1347,N_1135);
or U4951 (N_4951,N_75,N_679);
nand U4952 (N_4952,N_744,N_90);
or U4953 (N_4953,N_1081,N_0);
nand U4954 (N_4954,N_1309,N_1097);
nor U4955 (N_4955,N_1852,N_240);
nor U4956 (N_4956,N_2023,N_565);
or U4957 (N_4957,N_643,N_802);
or U4958 (N_4958,N_1121,N_1967);
nand U4959 (N_4959,N_385,N_1165);
nor U4960 (N_4960,N_677,N_355);
or U4961 (N_4961,N_992,N_314);
or U4962 (N_4962,N_1909,N_651);
or U4963 (N_4963,N_1431,N_1022);
nor U4964 (N_4964,N_1108,N_2186);
or U4965 (N_4965,N_745,N_2392);
nor U4966 (N_4966,N_1958,N_2370);
or U4967 (N_4967,N_2493,N_217);
or U4968 (N_4968,N_1585,N_1357);
or U4969 (N_4969,N_278,N_522);
or U4970 (N_4970,N_412,N_1420);
xor U4971 (N_4971,N_856,N_1261);
and U4972 (N_4972,N_1862,N_2355);
nor U4973 (N_4973,N_1357,N_902);
xor U4974 (N_4974,N_655,N_2031);
nor U4975 (N_4975,N_506,N_1107);
nor U4976 (N_4976,N_327,N_2470);
and U4977 (N_4977,N_674,N_2130);
nor U4978 (N_4978,N_1177,N_2027);
and U4979 (N_4979,N_306,N_2385);
xor U4980 (N_4980,N_2287,N_891);
and U4981 (N_4981,N_490,N_385);
nor U4982 (N_4982,N_2444,N_1500);
nor U4983 (N_4983,N_1418,N_803);
nor U4984 (N_4984,N_256,N_1780);
or U4985 (N_4985,N_1902,N_126);
and U4986 (N_4986,N_1432,N_139);
nor U4987 (N_4987,N_2246,N_1046);
and U4988 (N_4988,N_2111,N_1333);
nor U4989 (N_4989,N_1274,N_1000);
or U4990 (N_4990,N_851,N_1005);
or U4991 (N_4991,N_2037,N_146);
and U4992 (N_4992,N_352,N_479);
nand U4993 (N_4993,N_2031,N_391);
nand U4994 (N_4994,N_928,N_531);
or U4995 (N_4995,N_2118,N_450);
and U4996 (N_4996,N_2462,N_352);
and U4997 (N_4997,N_60,N_2234);
and U4998 (N_4998,N_2253,N_413);
or U4999 (N_4999,N_1823,N_2344);
nor UO_0 (O_0,N_2736,N_4461);
xor UO_1 (O_1,N_3483,N_3028);
xor UO_2 (O_2,N_3125,N_4101);
xor UO_3 (O_3,N_3961,N_3620);
or UO_4 (O_4,N_3965,N_4372);
or UO_5 (O_5,N_3628,N_4645);
xor UO_6 (O_6,N_4219,N_3410);
nand UO_7 (O_7,N_3309,N_3438);
or UO_8 (O_8,N_3109,N_2880);
or UO_9 (O_9,N_4562,N_2990);
and UO_10 (O_10,N_4592,N_3909);
or UO_11 (O_11,N_3541,N_3416);
and UO_12 (O_12,N_4530,N_4678);
nor UO_13 (O_13,N_4572,N_2920);
or UO_14 (O_14,N_3161,N_2961);
or UO_15 (O_15,N_3845,N_3566);
xnor UO_16 (O_16,N_4875,N_4115);
or UO_17 (O_17,N_3281,N_4470);
or UO_18 (O_18,N_3949,N_3128);
or UO_19 (O_19,N_4513,N_2659);
nand UO_20 (O_20,N_3137,N_3230);
or UO_21 (O_21,N_4610,N_3334);
and UO_22 (O_22,N_3231,N_3238);
nand UO_23 (O_23,N_4792,N_3343);
nor UO_24 (O_24,N_3964,N_3015);
nand UO_25 (O_25,N_4494,N_4350);
and UO_26 (O_26,N_4847,N_3602);
xor UO_27 (O_27,N_3618,N_3720);
nand UO_28 (O_28,N_3185,N_3837);
nor UO_29 (O_29,N_3728,N_4223);
nor UO_30 (O_30,N_4813,N_4741);
and UO_31 (O_31,N_4553,N_2682);
nand UO_32 (O_32,N_4573,N_3619);
xnor UO_33 (O_33,N_4417,N_4708);
xor UO_34 (O_34,N_4776,N_3561);
nand UO_35 (O_35,N_2928,N_4008);
and UO_36 (O_36,N_4510,N_3919);
or UO_37 (O_37,N_2885,N_4966);
nor UO_38 (O_38,N_3203,N_3385);
nor UO_39 (O_39,N_2515,N_4180);
xor UO_40 (O_40,N_4000,N_4696);
or UO_41 (O_41,N_4782,N_4785);
or UO_42 (O_42,N_3900,N_2790);
nor UO_43 (O_43,N_4770,N_4612);
xnor UO_44 (O_44,N_4184,N_3951);
xnor UO_45 (O_45,N_3682,N_4984);
nand UO_46 (O_46,N_3372,N_3145);
nand UO_47 (O_47,N_4172,N_4340);
nand UO_48 (O_48,N_2672,N_2673);
or UO_49 (O_49,N_3567,N_4013);
nor UO_50 (O_50,N_4070,N_3332);
xnor UO_51 (O_51,N_2611,N_2729);
xor UO_52 (O_52,N_2509,N_2860);
and UO_53 (O_53,N_4760,N_3724);
or UO_54 (O_54,N_2817,N_3974);
and UO_55 (O_55,N_4896,N_4982);
xnor UO_56 (O_56,N_4291,N_3224);
nand UO_57 (O_57,N_3119,N_3898);
and UO_58 (O_58,N_3051,N_3430);
and UO_59 (O_59,N_3252,N_4439);
and UO_60 (O_60,N_4900,N_3812);
nand UO_61 (O_61,N_4668,N_2958);
xnor UO_62 (O_62,N_3314,N_3476);
nor UO_63 (O_63,N_2999,N_3464);
nand UO_64 (O_64,N_4622,N_4698);
and UO_65 (O_65,N_2839,N_2896);
or UO_66 (O_66,N_3253,N_2779);
nor UO_67 (O_67,N_3838,N_4416);
nor UO_68 (O_68,N_4282,N_2665);
and UO_69 (O_69,N_2976,N_4485);
and UO_70 (O_70,N_2607,N_3368);
nor UO_71 (O_71,N_4048,N_3342);
nand UO_72 (O_72,N_4570,N_3489);
nand UO_73 (O_73,N_3765,N_3569);
nand UO_74 (O_74,N_3383,N_4615);
nand UO_75 (O_75,N_4499,N_2760);
and UO_76 (O_76,N_2545,N_3591);
or UO_77 (O_77,N_2900,N_3741);
and UO_78 (O_78,N_4867,N_2874);
nand UO_79 (O_79,N_4186,N_2612);
or UO_80 (O_80,N_3081,N_4835);
xor UO_81 (O_81,N_2588,N_4182);
or UO_82 (O_82,N_4444,N_3304);
nand UO_83 (O_83,N_4561,N_2934);
nor UO_84 (O_84,N_4203,N_4860);
xnor UO_85 (O_85,N_3413,N_2604);
and UO_86 (O_86,N_4756,N_4791);
and UO_87 (O_87,N_4558,N_3208);
xor UO_88 (O_88,N_4322,N_3434);
or UO_89 (O_89,N_2828,N_3110);
nand UO_90 (O_90,N_3731,N_3318);
nor UO_91 (O_91,N_4659,N_3112);
and UO_92 (O_92,N_2582,N_2763);
and UO_93 (O_93,N_4932,N_3752);
nand UO_94 (O_94,N_3221,N_3933);
xnor UO_95 (O_95,N_3364,N_4763);
and UO_96 (O_96,N_3590,N_3597);
nor UO_97 (O_97,N_3335,N_2734);
or UO_98 (O_98,N_3158,N_2911);
and UO_99 (O_99,N_3860,N_3380);
nor UO_100 (O_100,N_4672,N_4166);
nand UO_101 (O_101,N_2596,N_2957);
or UO_102 (O_102,N_4920,N_4464);
xor UO_103 (O_103,N_3691,N_3709);
nand UO_104 (O_104,N_4113,N_3574);
and UO_105 (O_105,N_3213,N_3504);
nor UO_106 (O_106,N_3348,N_2730);
nor UO_107 (O_107,N_3576,N_4451);
nand UO_108 (O_108,N_3705,N_4980);
or UO_109 (O_109,N_4517,N_3874);
nand UO_110 (O_110,N_4635,N_3942);
nor UO_111 (O_111,N_3911,N_4975);
nor UO_112 (O_112,N_2791,N_4853);
and UO_113 (O_113,N_2831,N_3772);
nor UO_114 (O_114,N_4625,N_3825);
nand UO_115 (O_115,N_4483,N_4035);
nor UO_116 (O_116,N_3465,N_4057);
xnor UO_117 (O_117,N_3747,N_4814);
nand UO_118 (O_118,N_3407,N_4560);
nor UO_119 (O_119,N_3722,N_4885);
xnor UO_120 (O_120,N_4097,N_2873);
or UO_121 (O_121,N_3578,N_3302);
nor UO_122 (O_122,N_3182,N_3516);
xnor UO_123 (O_123,N_3120,N_4978);
and UO_124 (O_124,N_2575,N_3408);
nand UO_125 (O_125,N_4440,N_4268);
nand UO_126 (O_126,N_3626,N_3074);
or UO_127 (O_127,N_3847,N_2866);
nand UO_128 (O_128,N_4640,N_4378);
xnor UO_129 (O_129,N_3894,N_4569);
nor UO_130 (O_130,N_4839,N_3868);
nor UO_131 (O_131,N_4010,N_3928);
and UO_132 (O_132,N_3036,N_4810);
and UO_133 (O_133,N_3131,N_3950);
xnor UO_134 (O_134,N_4638,N_2884);
and UO_135 (O_135,N_4589,N_2576);
nor UO_136 (O_136,N_3688,N_4380);
and UO_137 (O_137,N_4170,N_4431);
or UO_138 (O_138,N_4759,N_2642);
xor UO_139 (O_139,N_3150,N_3506);
and UO_140 (O_140,N_3684,N_4206);
nor UO_141 (O_141,N_4263,N_4582);
nor UO_142 (O_142,N_2719,N_3910);
nor UO_143 (O_143,N_3733,N_2706);
nor UO_144 (O_144,N_2955,N_2773);
xnor UO_145 (O_145,N_4945,N_3249);
and UO_146 (O_146,N_4376,N_2586);
nor UO_147 (O_147,N_3514,N_2688);
xnor UO_148 (O_148,N_3736,N_3536);
or UO_149 (O_149,N_4029,N_3777);
or UO_150 (O_150,N_4241,N_4546);
nor UO_151 (O_151,N_2959,N_3114);
or UO_152 (O_152,N_2947,N_4079);
and UO_153 (O_153,N_3633,N_4691);
or UO_154 (O_154,N_4019,N_3908);
nand UO_155 (O_155,N_4096,N_3169);
nor UO_156 (O_156,N_3534,N_4873);
xor UO_157 (O_157,N_4408,N_3607);
xnor UO_158 (O_158,N_3431,N_3533);
xor UO_159 (O_159,N_4762,N_2666);
and UO_160 (O_160,N_4744,N_2806);
xor UO_161 (O_161,N_3641,N_3844);
nor UO_162 (O_162,N_3505,N_3895);
nor UO_163 (O_163,N_4627,N_4928);
nand UO_164 (O_164,N_4005,N_3258);
xnor UO_165 (O_165,N_3658,N_2544);
or UO_166 (O_166,N_3210,N_3518);
and UO_167 (O_167,N_3850,N_4397);
and UO_168 (O_168,N_4298,N_4872);
nand UO_169 (O_169,N_3796,N_4686);
or UO_170 (O_170,N_2762,N_4534);
nand UO_171 (O_171,N_2618,N_4652);
and UO_172 (O_172,N_4418,N_4921);
or UO_173 (O_173,N_4617,N_3341);
xnor UO_174 (O_174,N_3694,N_4430);
nand UO_175 (O_175,N_3425,N_4196);
nand UO_176 (O_176,N_4198,N_2766);
xor UO_177 (O_177,N_3756,N_4447);
xnor UO_178 (O_178,N_3593,N_4309);
or UO_179 (O_179,N_4877,N_3681);
or UO_180 (O_180,N_4212,N_3059);
and UO_181 (O_181,N_4199,N_4717);
xnor UO_182 (O_182,N_2695,N_2549);
nand UO_183 (O_183,N_3347,N_3645);
and UO_184 (O_184,N_4207,N_3463);
and UO_185 (O_185,N_2756,N_3156);
nor UO_186 (O_186,N_2548,N_3117);
or UO_187 (O_187,N_3157,N_4112);
xor UO_188 (O_188,N_4099,N_3427);
nor UO_189 (O_189,N_3537,N_4861);
and UO_190 (O_190,N_2712,N_4169);
and UO_191 (O_191,N_3599,N_4269);
and UO_192 (O_192,N_2615,N_2914);
nand UO_193 (O_193,N_2853,N_3631);
or UO_194 (O_194,N_4834,N_3798);
nand UO_195 (O_195,N_2675,N_2621);
nand UO_196 (O_196,N_3194,N_4362);
or UO_197 (O_197,N_2707,N_3274);
and UO_198 (O_198,N_4064,N_2902);
nor UO_199 (O_199,N_3746,N_4068);
nand UO_200 (O_200,N_4665,N_3472);
nor UO_201 (O_201,N_2669,N_2534);
xor UO_202 (O_202,N_4290,N_4209);
xor UO_203 (O_203,N_3075,N_3244);
nand UO_204 (O_204,N_4168,N_4826);
or UO_205 (O_205,N_3057,N_4364);
xor UO_206 (O_206,N_2811,N_4520);
and UO_207 (O_207,N_4663,N_2975);
nand UO_208 (O_208,N_4069,N_4969);
and UO_209 (O_209,N_2567,N_4548);
nor UO_210 (O_210,N_2563,N_4247);
xnor UO_211 (O_211,N_4748,N_4383);
xnor UO_212 (O_212,N_4690,N_2517);
or UO_213 (O_213,N_2585,N_3762);
nor UO_214 (O_214,N_3927,N_2605);
or UO_215 (O_215,N_3735,N_4001);
xnor UO_216 (O_216,N_3629,N_4993);
xnor UO_217 (O_217,N_4527,N_2812);
and UO_218 (O_218,N_2737,N_2747);
or UO_219 (O_219,N_3642,N_2561);
xnor UO_220 (O_220,N_3455,N_3932);
and UO_221 (O_221,N_3976,N_4590);
nor UO_222 (O_222,N_3307,N_3826);
and UO_223 (O_223,N_2973,N_3967);
nor UO_224 (O_224,N_4915,N_2614);
or UO_225 (O_225,N_4695,N_3888);
and UO_226 (O_226,N_3099,N_4874);
or UO_227 (O_227,N_4404,N_3497);
nor UO_228 (O_228,N_4012,N_3362);
or UO_229 (O_229,N_4858,N_3917);
nor UO_230 (O_230,N_4751,N_4230);
nor UO_231 (O_231,N_2858,N_3127);
or UO_232 (O_232,N_4058,N_4133);
and UO_233 (O_233,N_4675,N_4111);
and UO_234 (O_234,N_3757,N_3700);
nand UO_235 (O_235,N_3575,N_2506);
or UO_236 (O_236,N_4466,N_4987);
nand UO_237 (O_237,N_4943,N_4796);
nand UO_238 (O_238,N_4654,N_4754);
and UO_239 (O_239,N_4339,N_3291);
or UO_240 (O_240,N_3292,N_2599);
nor UO_241 (O_241,N_3418,N_4793);
nor UO_242 (O_242,N_2513,N_4947);
or UO_243 (O_243,N_2821,N_3811);
and UO_244 (O_244,N_3164,N_3530);
and UO_245 (O_245,N_3241,N_3889);
xor UO_246 (O_246,N_3393,N_2690);
nand UO_247 (O_247,N_3205,N_3921);
or UO_248 (O_248,N_3470,N_3012);
nand UO_249 (O_249,N_3179,N_4934);
and UO_250 (O_250,N_2882,N_3284);
or UO_251 (O_251,N_4865,N_3638);
xnor UO_252 (O_252,N_3554,N_2661);
or UO_253 (O_253,N_4514,N_4492);
or UO_254 (O_254,N_4882,N_4018);
xor UO_255 (O_255,N_2716,N_4964);
xnor UO_256 (O_256,N_3596,N_2984);
or UO_257 (O_257,N_2648,N_3474);
nand UO_258 (O_258,N_2699,N_3201);
xor UO_259 (O_259,N_4401,N_4563);
or UO_260 (O_260,N_2512,N_4999);
and UO_261 (O_261,N_3317,N_4123);
nand UO_262 (O_262,N_4116,N_4733);
and UO_263 (O_263,N_3613,N_4491);
xnor UO_264 (O_264,N_4072,N_4160);
or UO_265 (O_265,N_3795,N_3938);
nor UO_266 (O_266,N_4041,N_4997);
nor UO_267 (O_267,N_2653,N_3035);
and UO_268 (O_268,N_3761,N_3995);
nor UO_269 (O_269,N_2935,N_4030);
and UO_270 (O_270,N_3106,N_3269);
xor UO_271 (O_271,N_4532,N_3990);
or UO_272 (O_272,N_3863,N_4077);
nor UO_273 (O_273,N_3622,N_2819);
or UO_274 (O_274,N_4065,N_3085);
or UO_275 (O_275,N_2713,N_3310);
and UO_276 (O_276,N_3495,N_3674);
nor UO_277 (O_277,N_2657,N_3262);
nor UO_278 (O_278,N_4666,N_3297);
and UO_279 (O_279,N_2643,N_2748);
and UO_280 (O_280,N_3625,N_2504);
nor UO_281 (O_281,N_3551,N_4375);
or UO_282 (O_282,N_3704,N_4434);
or UO_283 (O_283,N_3487,N_2967);
nand UO_284 (O_284,N_3047,N_4356);
nor UO_285 (O_285,N_3861,N_3880);
nor UO_286 (O_286,N_3417,N_2754);
and UO_287 (O_287,N_3998,N_2970);
nand UO_288 (O_288,N_3939,N_2619);
nand UO_289 (O_289,N_3359,N_3149);
or UO_290 (O_290,N_2587,N_3115);
nor UO_291 (O_291,N_4670,N_2540);
nor UO_292 (O_292,N_4593,N_4124);
and UO_293 (O_293,N_4887,N_2630);
and UO_294 (O_294,N_2617,N_4849);
xor UO_295 (O_295,N_4130,N_3764);
and UO_296 (O_296,N_3415,N_4869);
and UO_297 (O_297,N_4927,N_2805);
xor UO_298 (O_298,N_3824,N_4803);
nor UO_299 (O_299,N_3184,N_3153);
nand UO_300 (O_300,N_2963,N_4528);
nor UO_301 (O_301,N_2733,N_2936);
or UO_302 (O_302,N_3617,N_4720);
nor UO_303 (O_303,N_2829,N_3839);
nor UO_304 (O_304,N_3776,N_3683);
nand UO_305 (O_305,N_2950,N_3461);
nand UO_306 (O_306,N_2650,N_3039);
xor UO_307 (O_307,N_2820,N_4074);
xor UO_308 (O_308,N_3133,N_4623);
xnor UO_309 (O_309,N_2854,N_4524);
and UO_310 (O_310,N_2658,N_3353);
or UO_311 (O_311,N_3801,N_3147);
xnor UO_312 (O_312,N_3245,N_2939);
and UO_313 (O_313,N_4727,N_4614);
nor UO_314 (O_314,N_3955,N_4076);
and UO_315 (O_315,N_3199,N_2606);
nand UO_316 (O_316,N_2759,N_4600);
nand UO_317 (O_317,N_4787,N_4837);
nand UO_318 (O_318,N_3215,N_2571);
or UO_319 (O_319,N_3229,N_3174);
and UO_320 (O_320,N_4963,N_4579);
or UO_321 (O_321,N_3283,N_4511);
xor UO_322 (O_322,N_4581,N_2671);
or UO_323 (O_323,N_2778,N_4738);
nor UO_324 (O_324,N_4293,N_2785);
xnor UO_325 (O_325,N_4798,N_4938);
nand UO_326 (O_326,N_3978,N_4507);
xor UO_327 (O_327,N_3711,N_2646);
xor UO_328 (O_328,N_4722,N_2813);
or UO_329 (O_329,N_3640,N_3496);
and UO_330 (O_330,N_3676,N_4246);
or UO_331 (O_331,N_4618,N_4661);
xor UO_332 (O_332,N_4693,N_3702);
nand UO_333 (O_333,N_3975,N_4551);
and UO_334 (O_334,N_3293,N_3195);
and UO_335 (O_335,N_3753,N_3124);
xor UO_336 (O_336,N_3319,N_4190);
or UO_337 (O_337,N_3443,N_4034);
xnor UO_338 (O_338,N_4038,N_3977);
xnor UO_339 (O_339,N_3480,N_3401);
nor UO_340 (O_340,N_4174,N_2772);
or UO_341 (O_341,N_2502,N_3255);
and UO_342 (O_342,N_2992,N_2865);
nand UO_343 (O_343,N_4047,N_4505);
xnor UO_344 (O_344,N_3616,N_4841);
and UO_345 (O_345,N_2768,N_2523);
xnor UO_346 (O_346,N_4862,N_2678);
xnor UO_347 (O_347,N_4484,N_4025);
or UO_348 (O_348,N_3377,N_3467);
and UO_349 (O_349,N_2944,N_3488);
xor UO_350 (O_350,N_4648,N_2893);
nand UO_351 (O_351,N_3126,N_3315);
nor UO_352 (O_352,N_3373,N_2765);
or UO_353 (O_353,N_3357,N_4660);
or UO_354 (O_354,N_2855,N_4347);
and UO_355 (O_355,N_3907,N_4619);
xor UO_356 (O_356,N_3903,N_2824);
and UO_357 (O_357,N_3077,N_3345);
or UO_358 (O_358,N_3649,N_3029);
nand UO_359 (O_359,N_4800,N_4537);
xor UO_360 (O_360,N_4024,N_4128);
and UO_361 (O_361,N_3079,N_3429);
or UO_362 (O_362,N_3584,N_4363);
and UO_363 (O_363,N_2834,N_3018);
nor UO_364 (O_364,N_3287,N_3264);
and UO_365 (O_365,N_3924,N_3484);
xnor UO_366 (O_366,N_3831,N_3271);
nor UO_367 (O_367,N_3183,N_2644);
nand UO_368 (O_368,N_4566,N_3941);
and UO_369 (O_369,N_3098,N_2538);
or UO_370 (O_370,N_2830,N_2696);
and UO_371 (O_371,N_3188,N_4059);
and UO_372 (O_372,N_3931,N_2832);
nor UO_373 (O_373,N_3775,N_4843);
nor UO_374 (O_374,N_3568,N_3991);
xnor UO_375 (O_375,N_4148,N_4119);
nor UO_376 (O_376,N_2647,N_3813);
or UO_377 (O_377,N_4580,N_3587);
nand UO_378 (O_378,N_2508,N_3759);
and UO_379 (O_379,N_2543,N_2693);
nor UO_380 (O_380,N_3686,N_4300);
nand UO_381 (O_381,N_4163,N_3089);
and UO_382 (O_382,N_2845,N_4385);
xnor UO_383 (O_383,N_2583,N_3611);
nor UO_384 (O_384,N_4147,N_4929);
and UO_385 (O_385,N_3651,N_3044);
and UO_386 (O_386,N_4996,N_2573);
or UO_387 (O_387,N_4159,N_4441);
nand UO_388 (O_388,N_3447,N_3376);
and UO_389 (O_389,N_3526,N_3737);
nand UO_390 (O_390,N_4348,N_3522);
xor UO_391 (O_391,N_3833,N_3486);
or UO_392 (O_392,N_4836,N_2901);
nand UO_393 (O_393,N_4667,N_2616);
nor UO_394 (O_394,N_3904,N_3088);
nor UO_395 (O_395,N_3080,N_3523);
nand UO_396 (O_396,N_3954,N_3771);
and UO_397 (O_397,N_4739,N_3206);
and UO_398 (O_398,N_4726,N_3621);
nor UO_399 (O_399,N_4585,N_2720);
xor UO_400 (O_400,N_3404,N_2985);
nand UO_401 (O_401,N_2952,N_3717);
nand UO_402 (O_402,N_3247,N_3548);
and UO_403 (O_403,N_4899,N_3993);
or UO_404 (O_404,N_4280,N_3460);
and UO_405 (O_405,N_4630,N_4395);
xor UO_406 (O_406,N_4091,N_3652);
nor UO_407 (O_407,N_3915,N_3040);
or UO_408 (O_408,N_4479,N_2589);
xnor UO_409 (O_409,N_4699,N_4925);
nor UO_410 (O_410,N_4205,N_3469);
xnor UO_411 (O_411,N_3782,N_2771);
or UO_412 (O_412,N_4767,N_4750);
and UO_413 (O_413,N_4543,N_4731);
xnor UO_414 (O_414,N_3450,N_4656);
nand UO_415 (O_415,N_2519,N_4676);
nand UO_416 (O_416,N_4080,N_2770);
nor UO_417 (O_417,N_3041,N_3084);
or UO_418 (O_418,N_4231,N_2681);
or UO_419 (O_419,N_3968,N_3251);
or UO_420 (O_420,N_3002,N_4480);
or UO_421 (O_421,N_4784,N_2557);
and UO_422 (O_422,N_4644,N_3398);
xor UO_423 (O_423,N_2722,N_4807);
or UO_424 (O_424,N_3354,N_3246);
and UO_425 (O_425,N_2809,N_4818);
xnor UO_426 (O_426,N_4802,N_3946);
or UO_427 (O_427,N_3048,N_4154);
nor UO_428 (O_428,N_4574,N_4185);
nand UO_429 (O_429,N_2835,N_2631);
nor UO_430 (O_430,N_4601,N_4463);
nor UO_431 (O_431,N_2739,N_4467);
and UO_432 (O_432,N_4095,N_4200);
nand UO_433 (O_433,N_4294,N_4914);
nand UO_434 (O_434,N_4248,N_3767);
or UO_435 (O_435,N_3062,N_3893);
nand UO_436 (O_436,N_4712,N_2546);
and UO_437 (O_437,N_3865,N_3187);
nand UO_438 (O_438,N_3056,N_4728);
xnor UO_439 (O_439,N_4301,N_4325);
nand UO_440 (O_440,N_4786,N_3073);
and UO_441 (O_441,N_4271,N_4711);
or UO_442 (O_442,N_4455,N_2925);
xor UO_443 (O_443,N_4565,N_4051);
and UO_444 (O_444,N_3725,N_2764);
or UO_445 (O_445,N_4349,N_4545);
or UO_446 (O_446,N_4542,N_4649);
nand UO_447 (O_447,N_2535,N_4308);
or UO_448 (O_448,N_4893,N_3139);
nor UO_449 (O_449,N_3037,N_3672);
or UO_450 (O_450,N_2687,N_3097);
nand UO_451 (O_451,N_3788,N_3799);
nand UO_452 (O_452,N_2641,N_3152);
nand UO_453 (O_453,N_2941,N_4732);
and UO_454 (O_454,N_2943,N_3326);
and UO_455 (O_455,N_4193,N_4224);
xnor UO_456 (O_456,N_4040,N_2592);
xnor UO_457 (O_457,N_4924,N_4682);
or UO_458 (O_458,N_4341,N_4237);
nor UO_459 (O_459,N_4028,N_3118);
nand UO_460 (O_460,N_3378,N_4314);
xnor UO_461 (O_461,N_4388,N_3592);
xor UO_462 (O_462,N_4578,N_4303);
xnor UO_463 (O_463,N_4150,N_3583);
nand UO_464 (O_464,N_4135,N_3632);
nor UO_465 (O_465,N_3462,N_2718);
and UO_466 (O_466,N_4707,N_4435);
nand UO_467 (O_467,N_4442,N_4912);
nor UO_468 (O_468,N_4469,N_4336);
or UO_469 (O_469,N_4216,N_4764);
and UO_470 (O_470,N_3481,N_4871);
nor UO_471 (O_471,N_4357,N_2871);
and UO_472 (O_472,N_4257,N_3096);
xnor UO_473 (O_473,N_2993,N_4603);
or UO_474 (O_474,N_4624,N_3280);
nor UO_475 (O_475,N_4178,N_3608);
xor UO_476 (O_476,N_3543,N_4344);
or UO_477 (O_477,N_4496,N_4998);
and UO_478 (O_478,N_3699,N_4226);
or UO_479 (O_479,N_2741,N_4536);
nor UO_480 (O_480,N_3170,N_2632);
nand UO_481 (O_481,N_3656,N_4254);
nand UO_482 (O_482,N_3891,N_4859);
nor UO_483 (O_483,N_4173,N_4394);
xnor UO_484 (O_484,N_3324,N_3276);
and UO_485 (O_485,N_2908,N_3884);
or UO_486 (O_486,N_4233,N_2578);
nor UO_487 (O_487,N_4549,N_3906);
xnor UO_488 (O_488,N_3814,N_3713);
nor UO_489 (O_489,N_4342,N_2856);
xor UO_490 (O_490,N_4351,N_4118);
and UO_491 (O_491,N_2807,N_2776);
or UO_492 (O_492,N_4983,N_3662);
or UO_493 (O_493,N_2680,N_3361);
nand UO_494 (O_494,N_3218,N_3832);
nor UO_495 (O_495,N_3542,N_2704);
or UO_496 (O_496,N_3854,N_4721);
nor UO_497 (O_497,N_4778,N_3563);
nand UO_498 (O_498,N_4897,N_3389);
and UO_499 (O_499,N_3167,N_2794);
and UO_500 (O_500,N_4252,N_4369);
xor UO_501 (O_501,N_2684,N_3178);
xor UO_502 (O_502,N_2982,N_4027);
xnor UO_503 (O_503,N_3953,N_2995);
or UO_504 (O_504,N_2574,N_3744);
and UO_505 (O_505,N_4541,N_4986);
nand UO_506 (O_506,N_2691,N_4253);
nand UO_507 (O_507,N_3142,N_4211);
and UO_508 (O_508,N_3003,N_2887);
nand UO_509 (O_509,N_3267,N_4042);
and UO_510 (O_510,N_2727,N_3479);
xor UO_511 (O_511,N_2715,N_4521);
xnor UO_512 (O_512,N_4423,N_4976);
nand UO_513 (O_513,N_2654,N_4462);
xnor UO_514 (O_514,N_3313,N_2801);
xor UO_515 (O_515,N_4677,N_4045);
nand UO_516 (O_516,N_2977,N_3789);
nand UO_517 (O_517,N_4629,N_3107);
or UO_518 (O_518,N_3585,N_3358);
xnor UO_519 (O_519,N_4037,N_4856);
nand UO_520 (O_520,N_3433,N_4371);
nand UO_521 (O_521,N_4884,N_3790);
xnor UO_522 (O_522,N_4650,N_3196);
and UO_523 (O_523,N_2742,N_4365);
nor UO_524 (O_524,N_4850,N_3134);
xnor UO_525 (O_525,N_3442,N_2938);
xnor UO_526 (O_526,N_4108,N_4031);
nor UO_527 (O_527,N_3755,N_3026);
nand UO_528 (O_528,N_4420,N_4954);
and UO_529 (O_529,N_2862,N_3233);
nor UO_530 (O_530,N_3610,N_4425);
nor UO_531 (O_531,N_3654,N_3912);
and UO_532 (O_532,N_4709,N_2721);
xnor UO_533 (O_533,N_2851,N_3586);
nor UO_534 (O_534,N_3687,N_4801);
or UO_535 (O_535,N_2676,N_4512);
nand UO_536 (O_536,N_4081,N_4774);
nor UO_537 (O_537,N_3971,N_4575);
nor UO_538 (O_538,N_4244,N_2668);
or UO_539 (O_539,N_4876,N_3272);
xnor UO_540 (O_540,N_4674,N_3395);
nand UO_541 (O_541,N_4152,N_4164);
nor UO_542 (O_542,N_2655,N_4453);
xor UO_543 (O_543,N_3983,N_3219);
or UO_544 (O_544,N_3856,N_3873);
nand UO_545 (O_545,N_3492,N_4533);
or UO_546 (O_546,N_4273,N_3999);
xor UO_547 (O_547,N_3996,N_3557);
or UO_548 (O_548,N_2677,N_2960);
or UO_549 (O_549,N_4225,N_4359);
and UO_550 (O_550,N_3154,N_4156);
or UO_551 (O_551,N_2988,N_3240);
and UO_552 (O_552,N_3667,N_3298);
nand UO_553 (O_553,N_2883,N_4473);
xnor UO_554 (O_554,N_4844,N_2781);
or UO_555 (O_555,N_2994,N_2881);
xnor UO_556 (O_556,N_4465,N_4310);
nand UO_557 (O_557,N_3288,N_4187);
xor UO_558 (O_558,N_3511,N_4555);
nand UO_559 (O_559,N_2686,N_2746);
nand UO_560 (O_560,N_4795,N_3300);
nand UO_561 (O_561,N_4790,N_3769);
nor UO_562 (O_562,N_3043,N_4468);
or UO_563 (O_563,N_4501,N_4783);
and UO_564 (O_564,N_3337,N_4519);
nand UO_565 (O_565,N_3604,N_4265);
nor UO_566 (O_566,N_3022,N_2971);
or UO_567 (O_567,N_3019,N_3582);
xor UO_568 (O_568,N_3052,N_3260);
or UO_569 (O_569,N_3817,N_3560);
or UO_570 (O_570,N_3108,N_3718);
nand UO_571 (O_571,N_2635,N_3513);
nand UO_572 (O_572,N_3094,N_2841);
nor UO_573 (O_573,N_3540,N_4179);
and UO_574 (O_574,N_3855,N_4552);
xor UO_575 (O_575,N_4234,N_4020);
and UO_576 (O_576,N_3405,N_3980);
nor UO_577 (O_577,N_2702,N_4806);
nand UO_578 (O_578,N_3008,N_4845);
nor UO_579 (O_579,N_3005,N_4278);
nand UO_580 (O_580,N_2634,N_3989);
nand UO_581 (O_581,N_2731,N_3957);
and UO_582 (O_582,N_4681,N_4974);
nor UO_583 (O_583,N_3212,N_2510);
xor UO_584 (O_584,N_4122,N_3565);
and UO_585 (O_585,N_2628,N_2590);
nor UO_586 (O_586,N_4973,N_3851);
nor UO_587 (O_587,N_2892,N_3650);
xnor UO_588 (O_588,N_4410,N_4358);
xnor UO_589 (O_589,N_3308,N_3539);
nand UO_590 (O_590,N_2863,N_4684);
xor UO_591 (O_591,N_2799,N_4387);
and UO_592 (O_592,N_2838,N_4633);
or UO_593 (O_593,N_3930,N_4078);
nand UO_594 (O_594,N_4229,N_3572);
xnor UO_595 (O_595,N_2933,N_3305);
or UO_596 (O_596,N_2907,N_3432);
or UO_597 (O_597,N_4281,N_4611);
nand UO_598 (O_598,N_4424,N_3806);
nor UO_599 (O_599,N_4402,N_4476);
xnor UO_600 (O_600,N_3171,N_3054);
nand UO_601 (O_601,N_4905,N_4327);
xnor UO_602 (O_602,N_4609,N_2572);
or UO_603 (O_603,N_4489,N_2753);
xor UO_604 (O_604,N_3509,N_4390);
or UO_605 (O_605,N_3981,N_3794);
nor UO_606 (O_606,N_3714,N_4328);
and UO_607 (O_607,N_3666,N_4941);
or UO_608 (O_608,N_2921,N_3388);
or UO_609 (O_609,N_2525,N_2916);
and UO_610 (O_610,N_4857,N_4498);
xor UO_611 (O_611,N_4106,N_2537);
xnor UO_612 (O_612,N_3296,N_4295);
nand UO_613 (O_613,N_3696,N_2584);
nor UO_614 (O_614,N_3780,N_2726);
and UO_615 (O_615,N_3935,N_3138);
xnor UO_616 (O_616,N_3076,N_4583);
and UO_617 (O_617,N_3328,N_2526);
nor UO_618 (O_618,N_3087,N_4755);
or UO_619 (O_619,N_3061,N_2986);
and UO_620 (O_620,N_4958,N_4531);
or UO_621 (O_621,N_4256,N_3719);
nor UO_622 (O_622,N_4333,N_4808);
nor UO_623 (O_623,N_4370,N_3234);
and UO_624 (O_624,N_3397,N_4036);
or UO_625 (O_625,N_2674,N_3792);
or UO_626 (O_626,N_3690,N_4535);
nor UO_627 (O_627,N_4804,N_4437);
or UO_628 (O_628,N_3414,N_4714);
or UO_629 (O_629,N_2700,N_4426);
xor UO_630 (O_630,N_4547,N_3290);
nor UO_631 (O_631,N_4706,N_3456);
xnor UO_632 (O_632,N_3890,N_2735);
xnor UO_633 (O_633,N_4276,N_3473);
and UO_634 (O_634,N_4317,N_4710);
xor UO_635 (O_635,N_2728,N_2848);
xnor UO_636 (O_636,N_4742,N_3129);
or UO_637 (O_637,N_3102,N_2919);
nor UO_638 (O_638,N_2979,N_3647);
or UO_639 (O_639,N_2656,N_3925);
nor UO_640 (O_640,N_3615,N_4326);
or UO_641 (O_641,N_3006,N_4673);
and UO_642 (O_642,N_2725,N_3521);
and UO_643 (O_643,N_3066,N_2598);
and UO_644 (O_644,N_3751,N_4937);
or UO_645 (O_645,N_3176,N_4302);
nor UO_646 (O_646,N_3994,N_2593);
and UO_647 (O_647,N_3243,N_3071);
xor UO_648 (O_648,N_3403,N_2698);
xor UO_649 (O_649,N_4641,N_4502);
xor UO_650 (O_650,N_4260,N_3146);
nor UO_651 (O_651,N_2749,N_4508);
nand UO_652 (O_652,N_2956,N_3236);
nand UO_653 (O_653,N_3653,N_2836);
nor UO_654 (O_654,N_4454,N_4799);
xor UO_655 (O_655,N_3175,N_2872);
nor UO_656 (O_656,N_2798,N_3943);
nand UO_657 (O_657,N_4120,N_4272);
and UO_658 (O_658,N_3552,N_3242);
nor UO_659 (O_659,N_4242,N_2804);
nor UO_660 (O_660,N_3623,N_4460);
or UO_661 (O_661,N_4620,N_3121);
or UO_662 (O_662,N_4428,N_2703);
or UO_663 (O_663,N_2527,N_4971);
nand UO_664 (O_664,N_4823,N_3250);
nand UO_665 (O_665,N_3130,N_3452);
nand UO_666 (O_666,N_3697,N_3273);
xor UO_667 (O_667,N_2926,N_4863);
and UO_668 (O_668,N_2837,N_2899);
or UO_669 (O_669,N_4669,N_4811);
nor UO_670 (O_670,N_4880,N_3329);
nor UO_671 (O_671,N_2683,N_4851);
nand UO_672 (O_672,N_2627,N_4382);
and UO_673 (O_673,N_2922,N_3870);
nand UO_674 (O_674,N_4655,N_3655);
nand UO_675 (O_675,N_3441,N_4107);
or UO_676 (O_676,N_4149,N_3701);
and UO_677 (O_677,N_4175,N_3214);
nand UO_678 (O_678,N_4985,N_4970);
xnor UO_679 (O_679,N_4194,N_4275);
xnor UO_680 (O_680,N_4734,N_2625);
nor UO_681 (O_681,N_3458,N_3286);
or UO_682 (O_682,N_3350,N_3009);
nor UO_683 (O_683,N_3078,N_2710);
or UO_684 (O_684,N_4771,N_4155);
or UO_685 (O_685,N_4923,N_3330);
or UO_686 (O_686,N_3449,N_4634);
and UO_687 (O_687,N_3321,N_4942);
xnor UO_688 (O_688,N_2917,N_3105);
nor UO_689 (O_689,N_4398,N_4197);
or UO_690 (O_690,N_3661,N_3500);
and UO_691 (O_691,N_2889,N_3198);
xnor UO_692 (O_692,N_4261,N_4956);
or UO_693 (O_693,N_3589,N_4052);
nand UO_694 (O_694,N_2823,N_4604);
xnor UO_695 (O_695,N_4775,N_3926);
nor UO_696 (O_696,N_3457,N_3637);
and UO_697 (O_697,N_4011,N_2553);
and UO_698 (O_698,N_2991,N_3843);
nand UO_699 (O_699,N_4637,N_4591);
xor UO_700 (O_700,N_3729,N_4373);
xnor UO_701 (O_701,N_4855,N_4789);
or UO_702 (O_702,N_3220,N_3708);
and UO_703 (O_703,N_2784,N_4222);
xnor UO_704 (O_704,N_4056,N_3818);
or UO_705 (O_705,N_2554,N_4481);
or UO_706 (O_706,N_4073,N_3093);
xnor UO_707 (O_707,N_4192,N_3340);
nor UO_708 (O_708,N_3168,N_2929);
nor UO_709 (O_709,N_4564,N_2859);
nor UO_710 (O_710,N_3546,N_3266);
nand UO_711 (O_711,N_3899,N_4161);
nand UO_712 (O_712,N_3103,N_3344);
and UO_713 (O_713,N_2711,N_4516);
nor UO_714 (O_714,N_4393,N_3922);
nor UO_715 (O_715,N_2564,N_3325);
or UO_716 (O_716,N_3886,N_2913);
or UO_717 (O_717,N_4820,N_4201);
nand UO_718 (O_718,N_4895,N_4730);
and UO_719 (O_719,N_4021,N_4664);
nor UO_720 (O_720,N_4331,N_3525);
and UO_721 (O_721,N_4827,N_3835);
nor UO_722 (O_722,N_3947,N_2558);
nand UO_723 (O_723,N_2503,N_4838);
nor UO_724 (O_724,N_3659,N_2843);
or UO_725 (O_725,N_3282,N_3809);
or UO_726 (O_726,N_4448,N_4458);
xnor UO_727 (O_727,N_4493,N_2743);
nand UO_728 (O_728,N_2581,N_2775);
and UO_729 (O_729,N_3435,N_2861);
nand UO_730 (O_730,N_4704,N_3186);
or UO_731 (O_731,N_2997,N_3677);
and UO_732 (O_732,N_2751,N_3689);
and UO_733 (O_733,N_4816,N_2708);
and UO_734 (O_734,N_4459,N_4421);
xor UO_735 (O_735,N_4407,N_4144);
and UO_736 (O_736,N_3603,N_3498);
xnor UO_737 (O_737,N_2595,N_2602);
and UO_738 (O_738,N_4062,N_4102);
xnor UO_739 (O_739,N_3132,N_2777);
nor UO_740 (O_740,N_2651,N_3881);
nand UO_741 (O_741,N_3237,N_3864);
and UO_742 (O_742,N_2550,N_2802);
xor UO_743 (O_743,N_3339,N_3069);
nor UO_744 (O_744,N_4104,N_3535);
and UO_745 (O_745,N_3820,N_2904);
nor UO_746 (O_746,N_2608,N_3952);
nand UO_747 (O_747,N_3805,N_2709);
xor UO_748 (O_748,N_3630,N_3092);
nand UO_749 (O_749,N_4270,N_4881);
nor UO_750 (O_750,N_2877,N_3400);
nand UO_751 (O_751,N_2639,N_2697);
nor UO_752 (O_752,N_4452,N_4486);
nor UO_753 (O_753,N_3779,N_3517);
xnor UO_754 (O_754,N_4017,N_3370);
xor UO_755 (O_755,N_3017,N_3594);
and UO_756 (O_756,N_2629,N_3913);
or UO_757 (O_757,N_2664,N_4414);
nand UO_758 (O_758,N_3723,N_2528);
and UO_759 (O_759,N_3992,N_4571);
nand UO_760 (O_760,N_3545,N_3369);
xor UO_761 (O_761,N_3163,N_2568);
xnor UO_762 (O_762,N_3090,N_4935);
nand UO_763 (O_763,N_4692,N_3958);
xor UO_764 (O_764,N_3972,N_2679);
or UO_765 (O_765,N_3573,N_2609);
nor UO_766 (O_766,N_4745,N_4361);
xor UO_767 (O_767,N_4264,N_4329);
or UO_768 (O_768,N_4949,N_3091);
xor UO_769 (O_769,N_3004,N_2894);
and UO_770 (O_770,N_4245,N_3834);
or UO_771 (O_771,N_4288,N_3100);
xor UO_772 (O_772,N_3693,N_4736);
and UO_773 (O_773,N_3648,N_4026);
xnor UO_774 (O_774,N_4046,N_2783);
and UO_775 (O_775,N_4482,N_3643);
and UO_776 (O_776,N_4386,N_4250);
or UO_777 (O_777,N_2833,N_3375);
or UO_778 (O_778,N_3712,N_4729);
and UO_779 (O_779,N_3204,N_4979);
xor UO_780 (O_780,N_4653,N_4355);
or UO_781 (O_781,N_4766,N_4377);
or UO_782 (O_782,N_2761,N_3278);
xnor UO_783 (O_783,N_3466,N_3371);
nor UO_784 (O_784,N_3225,N_2744);
or UO_785 (O_785,N_3387,N_2827);
nand UO_786 (O_786,N_4142,N_3673);
nor UO_787 (O_787,N_4824,N_4315);
nand UO_788 (O_788,N_2918,N_2815);
nand UO_789 (O_789,N_4286,N_4181);
nor UO_790 (O_790,N_3679,N_3294);
nand UO_791 (O_791,N_3356,N_3064);
xnor UO_792 (O_792,N_3644,N_3490);
nor UO_793 (O_793,N_4445,N_3223);
or UO_794 (O_794,N_2514,N_4768);
and UO_795 (O_795,N_2910,N_2930);
and UO_796 (O_796,N_4616,N_3646);
and UO_797 (O_797,N_2816,N_4381);
nor UO_798 (O_798,N_3259,N_4719);
nor UO_799 (O_799,N_3451,N_3349);
and UO_800 (O_800,N_3083,N_2937);
nand UO_801 (O_801,N_3478,N_3406);
or UO_802 (O_802,N_3366,N_3787);
or UO_803 (O_803,N_4353,N_3740);
nand UO_804 (O_804,N_3636,N_4083);
and UO_805 (O_805,N_3095,N_3053);
nor UO_806 (O_806,N_2810,N_4438);
nor UO_807 (O_807,N_3058,N_3559);
or UO_808 (O_808,N_4162,N_3885);
nand UO_809 (O_809,N_4671,N_3876);
and UO_810 (O_810,N_2846,N_3745);
and UO_811 (O_811,N_2867,N_2886);
and UO_812 (O_812,N_2875,N_2951);
nor UO_813 (O_813,N_4687,N_4221);
xnor UO_814 (O_814,N_4171,N_2864);
xor UO_815 (O_815,N_2972,N_4886);
xnor UO_816 (O_816,N_4258,N_2962);
and UO_817 (O_817,N_3600,N_2620);
and UO_818 (O_818,N_2524,N_3363);
nand UO_819 (O_819,N_4140,N_3760);
or UO_820 (O_820,N_3166,N_2520);
nor UO_821 (O_821,N_4992,N_4683);
nor UO_822 (O_822,N_3730,N_4204);
nand UO_823 (O_823,N_3011,N_2826);
and UO_824 (O_824,N_3710,N_4828);
or UO_825 (O_825,N_4183,N_3671);
or UO_826 (O_826,N_4957,N_4946);
and UO_827 (O_827,N_2822,N_4832);
nor UO_828 (O_828,N_4883,N_3419);
nor UO_829 (O_829,N_2792,N_2912);
xnor UO_830 (O_830,N_3609,N_4657);
and UO_831 (O_831,N_3437,N_4607);
xor UO_832 (O_832,N_2752,N_3454);
xnor UO_833 (O_833,N_3190,N_4478);
and UO_834 (O_834,N_2906,N_4006);
xor UO_835 (O_835,N_3743,N_4337);
and UO_836 (O_836,N_2521,N_4890);
and UO_837 (O_837,N_4267,N_4497);
nand UO_838 (O_838,N_4747,N_3123);
nor UO_839 (O_839,N_3657,N_2888);
nor UO_840 (O_840,N_4312,N_4490);
nand UO_841 (O_841,N_3905,N_3807);
or UO_842 (O_842,N_3721,N_4909);
nand UO_843 (O_843,N_4167,N_4189);
nand UO_844 (O_844,N_4227,N_4777);
nor UO_845 (O_845,N_4725,N_2694);
and UO_846 (O_846,N_3882,N_4240);
nor UO_847 (O_847,N_2998,N_2638);
nand UO_848 (O_848,N_3042,N_2940);
nor UO_849 (O_849,N_3836,N_3959);
nor UO_850 (O_850,N_3140,N_4251);
and UO_851 (O_851,N_4471,N_4132);
or UO_852 (O_852,N_4723,N_4515);
or UO_853 (O_853,N_3969,N_3507);
xnor UO_854 (O_854,N_4931,N_2560);
xnor UO_855 (O_855,N_3923,N_3793);
nor UO_856 (O_856,N_3544,N_2755);
or UO_857 (O_857,N_2965,N_4389);
nand UO_858 (O_858,N_2740,N_3768);
xor UO_859 (O_859,N_4903,N_2964);
xnor UO_860 (O_860,N_2898,N_2840);
or UO_861 (O_861,N_2667,N_4319);
or UO_862 (O_862,N_3355,N_3520);
nand UO_863 (O_863,N_4679,N_3217);
and UO_864 (O_864,N_4697,N_3409);
or UO_865 (O_865,N_4043,N_3842);
xnor UO_866 (O_866,N_3316,N_4831);
nand UO_867 (O_867,N_3948,N_3944);
or UO_868 (O_868,N_3180,N_3529);
nor UO_869 (O_869,N_4427,N_3141);
or UO_870 (O_870,N_4538,N_4995);
or UO_871 (O_871,N_4879,N_4917);
or UO_872 (O_872,N_4870,N_4143);
xor UO_873 (O_873,N_3553,N_3268);
nor UO_874 (O_874,N_2774,N_4151);
xor UO_875 (O_875,N_3670,N_4737);
xor UO_876 (O_876,N_2532,N_3783);
xor UO_877 (O_877,N_4749,N_3299);
nor UO_878 (O_878,N_2566,N_4283);
nor UO_879 (O_879,N_4658,N_2547);
nand UO_880 (O_880,N_2932,N_3945);
nor UO_881 (O_881,N_2954,N_3634);
and UO_882 (O_882,N_4989,N_4321);
xor UO_883 (O_883,N_4817,N_3038);
and UO_884 (O_884,N_3270,N_4366);
and UO_885 (O_885,N_3192,N_4304);
nand UO_886 (O_886,N_2849,N_3510);
and UO_887 (O_887,N_3853,N_3428);
or UO_888 (O_888,N_3985,N_2577);
and UO_889 (O_889,N_4584,N_4049);
and UO_890 (O_890,N_3918,N_4346);
nor UO_891 (O_891,N_4157,N_4587);
nor UO_892 (O_892,N_4367,N_2559);
and UO_893 (O_893,N_3754,N_4279);
nor UO_894 (O_894,N_3791,N_2518);
and UO_895 (O_895,N_4930,N_4833);
and UO_896 (O_896,N_4972,N_3892);
nand UO_897 (O_897,N_3519,N_4632);
nor UO_898 (O_898,N_3781,N_3113);
nand UO_899 (O_899,N_3675,N_3338);
and UO_900 (O_900,N_4509,N_3605);
and UO_901 (O_901,N_4352,N_3396);
and UO_902 (O_902,N_2787,N_2689);
nor UO_903 (O_903,N_3550,N_4894);
or UO_904 (O_904,N_3896,N_2692);
and UO_905 (O_905,N_4188,N_4597);
nor UO_906 (O_906,N_3257,N_4743);
and UO_907 (O_907,N_3275,N_3527);
or UO_908 (O_908,N_3562,N_3785);
nand UO_909 (O_909,N_3846,N_2542);
nand UO_910 (O_910,N_3742,N_2895);
xnor UO_911 (O_911,N_3444,N_3439);
xor UO_912 (O_912,N_4412,N_4094);
nor UO_913 (O_913,N_2818,N_4131);
or UO_914 (O_914,N_4297,N_3878);
xor UO_915 (O_915,N_3822,N_3381);
xnor UO_916 (O_916,N_4121,N_2640);
nor UO_917 (O_917,N_2850,N_3564);
nand UO_918 (O_918,N_4396,N_2714);
or UO_919 (O_919,N_4146,N_4153);
and UO_920 (O_920,N_4948,N_4529);
and UO_921 (O_921,N_2594,N_3515);
xnor UO_922 (O_922,N_2869,N_4628);
nand UO_923 (O_923,N_3191,N_4285);
nor UO_924 (O_924,N_3614,N_3727);
nor UO_925 (O_925,N_3014,N_4399);
or UO_926 (O_926,N_4039,N_4236);
nor UO_927 (O_927,N_4940,N_4391);
nand UO_928 (O_928,N_4136,N_4345);
xnor UO_929 (O_929,N_4495,N_4705);
nand UO_930 (O_930,N_3962,N_3749);
nor UO_931 (O_931,N_4602,N_4988);
and UO_932 (O_932,N_4892,N_3374);
nor UO_933 (O_933,N_3528,N_4266);
or UO_934 (O_934,N_3181,N_4446);
and UO_935 (O_935,N_3830,N_3558);
nor UO_936 (O_936,N_2987,N_2793);
xor UO_937 (O_937,N_3289,N_4919);
and UO_938 (O_938,N_3828,N_2551);
or UO_939 (O_939,N_4338,N_4292);
nand UO_940 (O_940,N_3877,N_2600);
and UO_941 (O_941,N_3067,N_2610);
nand UO_942 (O_942,N_2968,N_3172);
nand UO_943 (O_943,N_3399,N_3800);
or UO_944 (O_944,N_4089,N_4313);
nand UO_945 (O_945,N_2541,N_3914);
xor UO_946 (O_946,N_2530,N_4559);
and UO_947 (O_947,N_4210,N_4274);
and UO_948 (O_948,N_3635,N_3209);
xnor UO_949 (O_949,N_4075,N_2556);
nand UO_950 (O_950,N_3000,N_4567);
nor UO_951 (O_951,N_3829,N_4898);
nand UO_952 (O_952,N_3261,N_4916);
or UO_953 (O_953,N_4289,N_3883);
xor UO_954 (O_954,N_4716,N_4066);
xnor UO_955 (O_955,N_2945,N_4259);
or UO_956 (O_956,N_3135,N_2897);
nor UO_957 (O_957,N_4878,N_4232);
nor UO_958 (O_958,N_2780,N_2636);
or UO_959 (O_959,N_4913,N_4208);
and UO_960 (O_960,N_4556,N_4500);
nand UO_961 (O_961,N_3581,N_3216);
nor UO_962 (O_962,N_4848,N_2522);
or UO_963 (O_963,N_2622,N_4085);
and UO_964 (O_964,N_3155,N_4752);
or UO_965 (O_965,N_4994,N_3422);
nor UO_966 (O_966,N_4586,N_2626);
nand UO_967 (O_967,N_4936,N_3547);
nor UO_968 (O_968,N_2870,N_4631);
and UO_969 (O_969,N_2663,N_3007);
or UO_970 (O_970,N_4218,N_4991);
nand UO_971 (O_971,N_4032,N_2905);
or UO_972 (O_972,N_3970,N_3226);
xor UO_973 (O_973,N_4474,N_3148);
nor UO_974 (O_974,N_3663,N_2797);
nand UO_975 (O_975,N_4249,N_3045);
nor UO_976 (O_976,N_4050,N_4922);
xor UO_977 (O_977,N_3784,N_2562);
and UO_978 (O_978,N_4568,N_3803);
and UO_979 (O_979,N_4621,N_4392);
nor UO_980 (O_980,N_4952,N_3323);
or UO_981 (O_981,N_2814,N_3144);
and UO_982 (O_982,N_2847,N_4651);
xnor UO_983 (O_983,N_3858,N_2942);
and UO_984 (O_984,N_4316,N_3580);
nand UO_985 (O_985,N_2649,N_2852);
or UO_986 (O_986,N_2603,N_2516);
or UO_987 (O_987,N_3436,N_4902);
and UO_988 (O_988,N_4195,N_4595);
xor UO_989 (O_989,N_3579,N_3823);
and UO_990 (O_990,N_3032,N_4780);
nand UO_991 (O_991,N_3197,N_3279);
xnor UO_992 (O_992,N_4599,N_4067);
or UO_993 (O_993,N_4926,N_4608);
nand UO_994 (O_994,N_3937,N_2879);
xor UO_995 (O_995,N_2732,N_3165);
nand UO_996 (O_996,N_4864,N_3421);
or UO_997 (O_997,N_4967,N_4740);
nor UO_998 (O_998,N_3664,N_3232);
nand UO_999 (O_999,N_4009,N_4287);
endmodule