module basic_3000_30000_3500_60_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_1375,In_1289);
xor U1 (N_1,In_2863,In_2998);
nand U2 (N_2,In_1319,In_2686);
or U3 (N_3,In_2518,In_2890);
xnor U4 (N_4,In_1839,In_393);
and U5 (N_5,In_1421,In_2960);
or U6 (N_6,In_2549,In_1000);
nand U7 (N_7,In_1649,In_2205);
nand U8 (N_8,In_2075,In_2544);
nand U9 (N_9,In_1064,In_1489);
nor U10 (N_10,In_104,In_506);
xor U11 (N_11,In_1197,In_127);
xor U12 (N_12,In_1951,In_232);
nor U13 (N_13,In_842,In_2651);
nor U14 (N_14,In_1745,In_2555);
or U15 (N_15,In_229,In_2839);
nor U16 (N_16,In_2985,In_1184);
and U17 (N_17,In_977,In_1730);
nand U18 (N_18,In_1211,In_1809);
nor U19 (N_19,In_1129,In_1728);
and U20 (N_20,In_2577,In_1876);
nor U21 (N_21,In_1294,In_844);
or U22 (N_22,In_2941,In_1066);
nand U23 (N_23,In_338,In_279);
nor U24 (N_24,In_2114,In_1552);
nand U25 (N_25,In_418,In_2212);
xor U26 (N_26,In_1468,In_649);
and U27 (N_27,In_2855,In_1061);
xnor U28 (N_28,In_353,In_1367);
and U29 (N_29,In_133,In_1723);
and U30 (N_30,In_165,In_845);
nand U31 (N_31,In_493,In_1223);
and U32 (N_32,In_2608,In_2828);
nor U33 (N_33,In_864,In_171);
and U34 (N_34,In_18,In_996);
nor U35 (N_35,In_1877,In_2167);
nor U36 (N_36,In_1984,In_2439);
nor U37 (N_37,In_2929,In_1970);
or U38 (N_38,In_1398,In_2055);
or U39 (N_39,In_868,In_93);
nand U40 (N_40,In_2599,In_26);
or U41 (N_41,In_488,In_1466);
and U42 (N_42,In_566,In_1547);
or U43 (N_43,In_2705,In_2742);
xor U44 (N_44,In_863,In_1896);
nor U45 (N_45,In_2028,In_1588);
xor U46 (N_46,In_2311,In_2783);
xor U47 (N_47,In_1964,In_1739);
and U48 (N_48,In_752,In_434);
nand U49 (N_49,In_2229,In_2852);
nand U50 (N_50,In_1352,In_101);
nand U51 (N_51,In_2942,In_2163);
and U52 (N_52,In_2967,In_430);
and U53 (N_53,In_2209,In_2709);
or U54 (N_54,In_2217,In_1677);
nor U55 (N_55,In_777,In_2889);
or U56 (N_56,In_1264,In_1540);
and U57 (N_57,In_2735,In_2513);
and U58 (N_58,In_2168,In_1406);
nand U59 (N_59,In_2778,In_399);
nor U60 (N_60,In_385,In_143);
nand U61 (N_61,In_732,In_391);
or U62 (N_62,In_745,In_439);
nor U63 (N_63,In_861,In_1616);
and U64 (N_64,In_283,In_541);
or U65 (N_65,In_90,In_627);
nor U66 (N_66,In_2943,In_1630);
and U67 (N_67,In_2566,In_1541);
or U68 (N_68,In_900,In_1621);
nor U69 (N_69,In_1538,In_873);
and U70 (N_70,In_2265,In_1667);
or U71 (N_71,In_1336,In_2085);
or U72 (N_72,In_1027,In_2860);
xnor U73 (N_73,In_1408,In_2576);
nor U74 (N_74,In_605,In_125);
nand U75 (N_75,In_1762,In_1248);
or U76 (N_76,In_2791,In_2614);
nor U77 (N_77,In_2550,In_619);
nor U78 (N_78,In_1875,In_1034);
or U79 (N_79,In_1228,In_1057);
nand U80 (N_80,In_2830,In_2479);
nand U81 (N_81,In_699,In_950);
and U82 (N_82,In_1535,In_982);
xnor U83 (N_83,In_961,In_1956);
xor U84 (N_84,In_1861,In_1308);
xor U85 (N_85,In_1437,In_2635);
xor U86 (N_86,In_2861,In_675);
nor U87 (N_87,In_1593,In_1442);
nand U88 (N_88,In_1212,In_1788);
and U89 (N_89,In_2474,In_162);
nor U90 (N_90,In_78,In_1718);
nand U91 (N_91,In_20,In_598);
and U92 (N_92,In_1881,In_2428);
and U93 (N_93,In_436,In_645);
nand U94 (N_94,In_2922,In_718);
nand U95 (N_95,In_289,In_1756);
nor U96 (N_96,In_755,In_2134);
and U97 (N_97,In_342,In_68);
nor U98 (N_98,In_967,In_2844);
or U99 (N_99,In_1700,In_2722);
nand U100 (N_100,In_1536,In_2988);
nand U101 (N_101,In_2367,In_2082);
or U102 (N_102,In_888,In_2720);
or U103 (N_103,In_145,In_875);
or U104 (N_104,In_2460,In_813);
nor U105 (N_105,In_2096,In_2851);
nor U106 (N_106,In_2763,In_1270);
xor U107 (N_107,In_651,In_2416);
or U108 (N_108,In_193,In_1794);
or U109 (N_109,In_526,In_15);
nor U110 (N_110,In_1586,In_2369);
nor U111 (N_111,In_1744,In_1166);
nor U112 (N_112,In_612,In_2071);
or U113 (N_113,In_543,In_1163);
nand U114 (N_114,In_2769,In_572);
nand U115 (N_115,In_2107,In_77);
nand U116 (N_116,In_511,In_1574);
xor U117 (N_117,In_2165,In_218);
nand U118 (N_118,In_1065,In_759);
and U119 (N_119,In_510,In_2485);
nand U120 (N_120,In_1385,In_2595);
nor U121 (N_121,In_2939,In_2658);
and U122 (N_122,In_2891,In_2013);
xnor U123 (N_123,In_444,In_1594);
nand U124 (N_124,In_2468,In_464);
or U125 (N_125,In_1342,In_1925);
or U126 (N_126,In_2154,In_797);
xnor U127 (N_127,In_764,In_979);
nor U128 (N_128,In_2208,In_452);
nand U129 (N_129,In_2568,In_1642);
nor U130 (N_130,In_2809,In_374);
or U131 (N_131,In_692,In_2696);
nor U132 (N_132,In_2878,In_2029);
or U133 (N_133,In_2237,In_637);
and U134 (N_134,In_1396,In_582);
nor U135 (N_135,In_2521,In_1268);
and U136 (N_136,In_2562,In_2571);
nand U137 (N_137,In_1172,In_858);
or U138 (N_138,In_1190,In_2068);
nand U139 (N_139,In_1662,In_2616);
xnor U140 (N_140,In_589,In_1518);
xor U141 (N_141,In_742,In_2321);
nor U142 (N_142,In_1329,In_2898);
nand U143 (N_143,In_1904,In_1988);
or U144 (N_144,In_336,In_81);
and U145 (N_145,In_50,In_1345);
or U146 (N_146,In_1845,In_639);
nor U147 (N_147,In_988,In_2829);
nand U148 (N_148,In_1765,In_1313);
xnor U149 (N_149,In_2282,In_297);
and U150 (N_150,In_1397,In_275);
xnor U151 (N_151,In_2279,In_1331);
nand U152 (N_152,In_2359,In_1237);
nor U153 (N_153,In_1678,In_787);
nor U154 (N_154,In_384,In_2415);
and U155 (N_155,In_517,In_515);
xnor U156 (N_156,In_2842,In_1917);
nor U157 (N_157,In_1058,In_1423);
nand U158 (N_158,In_243,In_725);
nor U159 (N_159,In_154,In_1224);
nor U160 (N_160,In_267,In_1870);
nor U161 (N_161,In_539,In_2190);
nand U162 (N_162,In_2181,In_2919);
nand U163 (N_163,In_1637,In_375);
and U164 (N_164,In_206,In_335);
nand U165 (N_165,In_2100,In_502);
and U166 (N_166,In_103,In_2470);
xor U167 (N_167,In_377,In_547);
or U168 (N_168,In_2031,In_1450);
and U169 (N_169,In_367,In_1288);
nand U170 (N_170,In_1400,In_1589);
and U171 (N_171,In_2370,In_705);
nand U172 (N_172,In_1068,In_2400);
nand U173 (N_173,In_2419,In_2600);
or U174 (N_174,In_2565,In_1692);
and U175 (N_175,In_2663,In_2202);
nand U176 (N_176,In_2040,In_1561);
or U177 (N_177,In_1451,In_422);
and U178 (N_178,In_1123,In_597);
and U179 (N_179,In_2827,In_521);
xnor U180 (N_180,In_1985,In_1822);
nor U181 (N_181,In_2307,In_1360);
and U182 (N_182,In_1100,In_720);
nand U183 (N_183,In_2533,In_579);
or U184 (N_184,In_1405,In_794);
nor U185 (N_185,In_1118,In_2270);
and U186 (N_186,In_1186,In_499);
xor U187 (N_187,In_792,In_2526);
nor U188 (N_188,In_1003,In_671);
and U189 (N_189,In_2802,In_1370);
nand U190 (N_190,In_1250,In_1439);
nor U191 (N_191,In_1980,In_2131);
nor U192 (N_192,In_230,In_2816);
nor U193 (N_193,In_1269,In_2932);
nor U194 (N_194,In_2540,In_2634);
nand U195 (N_195,In_169,In_2669);
nor U196 (N_196,In_1151,In_288);
nor U197 (N_197,In_226,In_2308);
nand U198 (N_198,In_333,In_501);
xnor U199 (N_199,In_886,In_1074);
nand U200 (N_200,In_721,In_1112);
xor U201 (N_201,In_14,In_100);
and U202 (N_202,In_558,In_1417);
xor U203 (N_203,In_1435,In_1615);
xnor U204 (N_204,In_10,In_459);
or U205 (N_205,In_1191,In_944);
nand U206 (N_206,In_2818,In_733);
xor U207 (N_207,In_1915,In_1539);
xnor U208 (N_208,In_144,In_2671);
or U209 (N_209,In_1585,In_487);
nor U210 (N_210,In_1444,In_2335);
or U211 (N_211,In_2664,In_1038);
and U212 (N_212,In_321,In_1015);
or U213 (N_213,In_2430,In_2053);
xnor U214 (N_214,In_2143,In_544);
or U215 (N_215,In_1998,In_1841);
nand U216 (N_216,In_743,In_1524);
and U217 (N_217,In_161,In_29);
nor U218 (N_218,In_1598,In_1638);
nor U219 (N_219,In_2707,In_2593);
nor U220 (N_220,In_1858,In_41);
nor U221 (N_221,In_601,In_296);
and U222 (N_222,In_298,In_1202);
nor U223 (N_223,In_2341,In_2346);
nand U224 (N_224,In_1001,In_657);
nand U225 (N_225,In_241,In_327);
nand U226 (N_226,In_2976,In_24);
nor U227 (N_227,In_851,In_2999);
xor U228 (N_228,In_1819,In_2272);
and U229 (N_229,In_766,In_223);
nand U230 (N_230,In_1651,In_2358);
nand U231 (N_231,In_2963,In_1495);
or U232 (N_232,In_2498,In_409);
and U233 (N_233,In_1101,In_2353);
or U234 (N_234,In_2807,In_1654);
nand U235 (N_235,In_2743,In_984);
nand U236 (N_236,In_2567,In_2357);
nor U237 (N_237,In_1275,In_1646);
or U238 (N_238,In_2453,In_1492);
xor U239 (N_239,In_2095,In_398);
xor U240 (N_240,In_1415,In_1154);
and U241 (N_241,In_1147,In_52);
xnor U242 (N_242,In_1726,In_912);
nand U243 (N_243,In_1207,In_1577);
nor U244 (N_244,In_121,In_271);
nor U245 (N_245,In_465,In_1244);
xor U246 (N_246,In_2937,In_2427);
and U247 (N_247,In_795,In_287);
and U248 (N_248,In_1773,In_2866);
xnor U249 (N_249,In_999,In_1880);
nand U250 (N_250,In_2139,In_2136);
or U251 (N_251,In_1363,In_2711);
and U252 (N_252,In_2340,In_1559);
nor U253 (N_253,In_2684,In_669);
xnor U254 (N_254,In_830,In_1835);
nor U255 (N_255,In_63,In_1470);
and U256 (N_256,In_1155,In_2384);
and U257 (N_257,In_2968,In_2284);
or U258 (N_258,In_553,In_542);
and U259 (N_259,In_1935,In_257);
xnor U260 (N_260,In_954,In_1712);
or U261 (N_261,In_2613,In_1084);
and U262 (N_262,In_1284,In_1920);
nor U263 (N_263,In_1316,In_835);
and U264 (N_264,In_1124,In_74);
and U265 (N_265,In_1203,In_307);
nand U266 (N_266,In_1204,In_1368);
nand U267 (N_267,In_1227,In_2322);
nand U268 (N_268,In_148,In_202);
or U269 (N_269,In_2491,In_753);
nor U270 (N_270,In_2219,In_2982);
nor U271 (N_271,In_435,In_951);
or U272 (N_272,In_805,In_1087);
and U273 (N_273,In_681,In_2009);
or U274 (N_274,In_1812,In_1401);
or U275 (N_275,In_2820,In_56);
xnor U276 (N_276,In_1431,In_2318);
or U277 (N_277,In_152,In_2724);
or U278 (N_278,In_2621,In_891);
nor U279 (N_279,In_2821,In_768);
or U280 (N_280,In_2245,In_856);
nor U281 (N_281,In_1688,In_463);
nand U282 (N_282,In_1633,In_1195);
nand U283 (N_283,In_334,In_2620);
xor U284 (N_284,In_1340,In_118);
nand U285 (N_285,In_1919,In_2670);
nand U286 (N_286,In_183,In_368);
or U287 (N_287,In_1945,In_2728);
nand U288 (N_288,In_2377,In_1814);
xnor U289 (N_289,In_505,In_2563);
and U290 (N_290,In_1735,In_1175);
and U291 (N_291,In_27,In_1500);
xnor U292 (N_292,In_1694,In_2733);
or U293 (N_293,In_449,In_884);
nand U294 (N_294,In_1210,In_952);
or U295 (N_295,In_1683,In_475);
or U296 (N_296,In_936,In_1800);
or U297 (N_297,In_1792,In_396);
nand U298 (N_298,In_744,In_2276);
xnor U299 (N_299,In_620,In_2961);
nand U300 (N_300,In_2597,In_848);
xor U301 (N_301,In_1140,In_1302);
and U302 (N_302,In_2730,In_840);
nand U303 (N_303,In_2652,In_2520);
and U304 (N_304,In_1452,In_2630);
xor U305 (N_305,In_280,In_673);
nand U306 (N_306,In_47,In_1252);
nand U307 (N_307,In_1384,In_802);
or U308 (N_308,In_909,In_926);
xor U309 (N_309,In_2674,In_723);
nand U310 (N_310,In_528,In_2257);
or U311 (N_311,In_1868,In_200);
and U312 (N_312,In_1987,In_432);
and U313 (N_313,In_1837,In_2347);
xor U314 (N_314,In_235,In_306);
and U315 (N_315,In_453,In_2266);
nor U316 (N_316,In_933,In_691);
nand U317 (N_317,In_1967,In_551);
nand U318 (N_318,In_2192,In_2708);
nand U319 (N_319,In_1299,In_2868);
and U320 (N_320,In_2339,In_2066);
and U321 (N_321,In_2099,In_2056);
nand U322 (N_322,In_484,In_2184);
and U323 (N_323,In_832,In_2456);
or U324 (N_324,In_2622,In_2719);
nor U325 (N_325,In_259,In_2657);
or U326 (N_326,In_1453,In_934);
xnor U327 (N_327,In_1560,In_1565);
nand U328 (N_328,In_1963,In_2414);
or U329 (N_329,In_316,In_1961);
or U330 (N_330,In_1042,In_2232);
xor U331 (N_331,In_2280,In_438);
nor U332 (N_332,In_1440,In_914);
and U333 (N_333,In_1070,In_2200);
nand U334 (N_334,In_1067,In_1648);
nor U335 (N_335,In_1848,In_88);
nor U336 (N_336,In_2538,In_650);
and U337 (N_337,In_1986,In_877);
xnor U338 (N_338,In_2499,In_1901);
and U339 (N_339,In_2602,In_548);
xor U340 (N_340,In_2754,In_2090);
xor U341 (N_341,In_2574,In_1395);
nor U342 (N_342,In_2945,In_734);
or U343 (N_343,In_2310,In_2086);
and U344 (N_344,In_2413,In_379);
xor U345 (N_345,In_80,In_1887);
nand U346 (N_346,In_2559,In_34);
nand U347 (N_347,In_910,In_1149);
nor U348 (N_348,In_390,In_2036);
and U349 (N_349,In_993,In_1626);
or U350 (N_350,In_904,In_1425);
and U351 (N_351,In_2203,In_395);
nand U352 (N_352,In_824,In_1078);
and U353 (N_353,In_414,In_2121);
or U354 (N_354,In_853,In_1239);
and U355 (N_355,In_1750,In_1566);
and U356 (N_356,In_1516,In_2870);
or U357 (N_357,In_2104,In_735);
nand U358 (N_358,In_1690,In_323);
or U359 (N_359,In_325,In_2843);
nor U360 (N_360,In_2760,In_878);
or U361 (N_361,In_2966,In_1357);
and U362 (N_362,In_689,In_789);
or U363 (N_363,In_146,In_217);
and U364 (N_364,In_1092,In_326);
nor U365 (N_365,In_437,In_1113);
and U366 (N_366,In_804,In_1706);
nor U367 (N_367,In_416,In_1869);
or U368 (N_368,In_277,In_2238);
nor U369 (N_369,In_1245,In_2546);
and U370 (N_370,In_507,In_2759);
xor U371 (N_371,In_1791,In_1082);
xor U372 (N_372,In_2695,In_1131);
xnor U373 (N_373,In_2410,In_1663);
nor U374 (N_374,In_1389,In_2133);
nor U375 (N_375,In_2481,In_1238);
nand U376 (N_376,In_2417,In_2834);
nor U377 (N_377,In_1139,In_773);
and U378 (N_378,In_1517,In_928);
or U379 (N_379,In_2320,In_1668);
or U380 (N_380,In_2281,In_2477);
nor U381 (N_381,In_1206,In_2761);
xnor U382 (N_382,In_917,In_2046);
and U383 (N_383,In_750,In_1691);
nand U384 (N_384,In_1088,In_172);
xor U385 (N_385,In_1590,In_1213);
xnor U386 (N_386,In_1684,In_2041);
and U387 (N_387,In_893,In_1254);
nor U388 (N_388,In_1031,In_2352);
and U389 (N_389,In_1995,In_343);
and U390 (N_390,In_2330,In_2247);
and U391 (N_391,In_1366,In_1196);
or U392 (N_392,In_2469,In_1624);
or U393 (N_393,In_722,In_22);
and U394 (N_394,In_1862,In_867);
or U395 (N_395,In_1009,In_1811);
or U396 (N_396,In_1183,In_383);
nand U397 (N_397,In_2749,In_2348);
or U398 (N_398,In_1827,In_916);
or U399 (N_399,In_1337,In_485);
or U400 (N_400,In_1596,In_2689);
nand U401 (N_401,In_1893,In_1362);
xor U402 (N_402,In_738,In_1682);
nor U403 (N_403,In_1815,In_2893);
and U404 (N_404,In_1643,In_780);
nor U405 (N_405,In_1923,In_2779);
or U406 (N_406,In_788,In_1382);
and U407 (N_407,In_2530,In_2242);
and U408 (N_408,In_2476,In_320);
nand U409 (N_409,In_739,In_220);
and U410 (N_410,In_362,In_2458);
or U411 (N_411,In_2064,In_117);
nor U412 (N_412,In_555,In_2291);
or U413 (N_413,In_339,In_1023);
nand U414 (N_414,In_2497,In_1371);
xor U415 (N_415,In_1666,In_2198);
and U416 (N_416,In_2706,In_953);
or U417 (N_417,In_2610,In_622);
xor U418 (N_418,In_2534,In_407);
or U419 (N_419,In_1493,In_2261);
or U420 (N_420,In_1906,In_1836);
nand U421 (N_421,In_1388,In_1619);
or U422 (N_422,In_532,In_2931);
nor U423 (N_423,In_1059,In_2473);
nand U424 (N_424,In_2901,In_2007);
and U425 (N_425,In_299,In_2011);
nand U426 (N_426,In_549,In_380);
xnor U427 (N_427,In_2024,In_2336);
or U428 (N_428,In_33,In_1287);
xor U429 (N_429,In_106,In_2973);
nand U430 (N_430,In_209,In_315);
nand U431 (N_431,In_2248,In_670);
or U432 (N_432,In_779,In_2044);
xor U433 (N_433,In_301,In_2455);
or U434 (N_434,In_2145,In_216);
nand U435 (N_435,In_84,In_823);
xor U436 (N_436,In_2611,In_2153);
nor U437 (N_437,In_468,In_2063);
xor U438 (N_438,In_2687,In_603);
or U439 (N_439,In_791,In_67);
or U440 (N_440,In_2106,In_621);
or U441 (N_441,In_329,In_2793);
xnor U442 (N_442,In_490,In_43);
xnor U443 (N_443,In_445,In_2659);
xor U444 (N_444,In_1569,In_2723);
and U445 (N_445,In_1958,In_2034);
nor U446 (N_446,In_1364,In_2527);
xor U447 (N_447,In_2426,In_1699);
nor U448 (N_448,In_1514,In_2636);
xnor U449 (N_449,In_2487,In_331);
xnor U450 (N_450,In_686,In_2289);
xnor U451 (N_451,In_625,In_2691);
or U452 (N_452,In_978,In_1576);
nand U453 (N_453,In_1855,In_2846);
xnor U454 (N_454,In_131,In_1424);
and U455 (N_455,In_1128,In_2558);
and U456 (N_456,In_577,In_786);
nor U457 (N_457,In_2298,In_1013);
nor U458 (N_458,In_2297,In_630);
nor U459 (N_459,In_1532,In_2074);
or U460 (N_460,In_923,In_2685);
nand U461 (N_461,In_1449,In_1927);
nor U462 (N_462,In_1079,In_2319);
nand U463 (N_463,In_882,In_516);
xor U464 (N_464,In_483,In_330);
nor U465 (N_465,In_1977,In_1290);
and U466 (N_466,In_1286,In_73);
and U467 (N_467,In_1892,In_2449);
xnor U468 (N_468,In_1736,In_1158);
nor U469 (N_469,In_2531,In_807);
xnor U470 (N_470,In_2551,In_1170);
xor U471 (N_471,In_2598,In_2510);
nor U472 (N_472,In_378,In_1929);
xnor U473 (N_473,In_1673,In_1355);
or U474 (N_474,In_2792,In_633);
and U475 (N_475,In_609,In_1020);
xnor U476 (N_476,In_1969,In_2152);
xor U477 (N_477,In_1146,In_1161);
and U478 (N_478,In_2758,In_1789);
xnor U479 (N_479,In_1,In_1055);
or U480 (N_480,In_2101,In_214);
nor U481 (N_481,In_1679,In_2629);
xnor U482 (N_482,In_1912,In_70);
nor U483 (N_483,In_682,In_666);
nand U484 (N_484,In_2949,In_1698);
nand U485 (N_485,In_546,In_401);
nor U486 (N_486,In_491,In_1035);
or U487 (N_487,In_568,In_2446);
nor U488 (N_488,In_2093,In_1181);
or U489 (N_489,In_1114,In_1446);
nor U490 (N_490,In_1693,In_246);
or U491 (N_491,In_1454,In_2971);
or U492 (N_492,In_290,In_1509);
nor U493 (N_493,In_1888,In_40);
or U494 (N_494,In_2983,In_2331);
or U495 (N_495,In_1942,In_2483);
or U496 (N_496,In_168,In_2268);
or U497 (N_497,In_76,In_1982);
nor U498 (N_498,In_871,In_1098);
nor U499 (N_499,In_1077,In_2808);
nor U500 (N_500,In_1222,In_32);
xnor U501 (N_501,In_1781,In_221);
nor U502 (N_502,In_2928,N_348);
xor U503 (N_503,In_2172,In_13);
xor U504 (N_504,In_2363,N_477);
xnor U505 (N_505,N_83,In_1826);
and U506 (N_506,In_1132,In_1188);
nor U507 (N_507,In_1377,In_1860);
or U508 (N_508,In_1932,In_1506);
xor U509 (N_509,In_1475,In_212);
and U510 (N_510,In_898,In_1661);
nand U511 (N_511,N_207,In_1808);
xor U512 (N_512,In_2327,In_119);
xor U513 (N_513,In_2964,In_61);
nor U514 (N_514,In_2383,In_676);
nor U515 (N_515,N_495,N_183);
xnor U516 (N_516,In_994,In_1613);
or U517 (N_517,In_2869,N_111);
nand U518 (N_518,In_1708,In_1898);
nand U519 (N_519,In_1966,In_890);
nand U520 (N_520,In_997,In_1665);
nand U521 (N_521,In_2376,In_1832);
or U522 (N_522,In_341,In_31);
nor U523 (N_523,In_476,In_854);
and U524 (N_524,In_458,In_2586);
and U525 (N_525,N_74,In_1640);
nor U526 (N_526,In_2718,In_939);
nor U527 (N_527,N_96,In_2437);
nand U528 (N_528,In_1926,In_2201);
nor U529 (N_529,N_438,In_1233);
nor U530 (N_530,In_2523,In_2117);
and U531 (N_531,In_2269,N_140);
nand U532 (N_532,N_409,In_942);
and U533 (N_533,In_160,N_213);
nor U534 (N_534,In_2740,In_2698);
nand U535 (N_535,In_932,N_441);
or U536 (N_536,In_796,In_1199);
or U537 (N_537,N_122,In_1740);
nor U538 (N_538,In_358,In_1004);
or U539 (N_539,In_2161,In_1310);
xor U540 (N_540,In_2258,N_159);
xor U541 (N_541,In_1217,In_346);
xor U542 (N_542,In_876,In_1419);
or U543 (N_543,In_1685,In_2374);
and U544 (N_544,In_2697,N_374);
nand U545 (N_545,N_360,In_429);
xnor U546 (N_546,In_2033,In_2182);
nor U547 (N_547,In_1962,In_1187);
nand U548 (N_548,N_497,In_1867);
or U549 (N_549,In_1469,N_186);
xnor U550 (N_550,In_606,In_2155);
xor U551 (N_551,In_664,In_1404);
xor U552 (N_552,N_234,In_1938);
nand U553 (N_553,In_2118,In_2507);
or U554 (N_554,In_489,In_1722);
nor U555 (N_555,In_2681,N_80);
nor U556 (N_556,In_1622,In_2881);
or U557 (N_557,N_193,N_117);
and U558 (N_558,In_1137,In_1564);
nor U559 (N_559,N_101,N_340);
nor U560 (N_560,In_2059,N_126);
or U561 (N_561,In_128,N_197);
xor U562 (N_562,N_440,N_65);
nor U563 (N_563,In_5,In_1656);
nor U564 (N_564,In_1544,In_2906);
nor U565 (N_565,In_8,In_1521);
nor U566 (N_566,In_674,In_1655);
and U567 (N_567,N_142,In_638);
and U568 (N_568,In_2867,In_2061);
nand U569 (N_569,In_2008,N_162);
xnor U570 (N_570,In_2344,In_1391);
or U571 (N_571,In_964,In_2097);
nand U572 (N_572,In_2825,In_317);
nand U573 (N_573,In_1768,In_1960);
xnor U574 (N_574,In_1556,In_1177);
or U575 (N_575,In_1767,In_1871);
nor U576 (N_576,In_2950,In_958);
or U577 (N_577,In_1018,In_584);
nand U578 (N_578,In_576,In_2433);
nand U579 (N_579,In_2704,In_931);
or U580 (N_580,In_2240,In_1089);
xnor U581 (N_581,In_965,N_342);
xnor U582 (N_582,N_323,In_701);
or U583 (N_583,In_1806,N_23);
and U584 (N_584,In_2638,In_197);
and U585 (N_585,In_1028,In_2677);
and U586 (N_586,N_308,In_811);
nor U587 (N_587,In_2235,In_2129);
xnor U588 (N_588,In_1631,In_1751);
nor U589 (N_589,In_2603,In_302);
and U590 (N_590,In_2128,N_398);
nor U591 (N_591,In_1763,In_2986);
or U592 (N_592,In_1924,In_1978);
nor U593 (N_593,In_2646,In_2349);
and U594 (N_594,In_83,In_2772);
or U595 (N_595,In_1026,N_408);
and U596 (N_596,In_1063,In_2582);
or U597 (N_597,In_2196,In_749);
or U598 (N_598,In_2978,In_902);
nor U599 (N_599,In_611,In_1676);
or U600 (N_600,In_1192,In_2037);
nor U601 (N_601,In_28,In_2462);
and U602 (N_602,In_2076,In_264);
or U603 (N_603,N_132,In_1081);
or U604 (N_604,In_2912,In_2023);
xor U605 (N_605,In_1039,In_837);
or U606 (N_606,In_2552,In_1818);
or U607 (N_607,In_956,N_450);
and U608 (N_608,In_2004,N_62);
or U609 (N_609,In_1443,In_2020);
and U610 (N_610,In_1142,In_2872);
and U611 (N_611,In_973,In_1324);
nand U612 (N_612,In_1753,N_384);
nand U613 (N_613,In_2899,N_76);
nor U614 (N_614,In_269,In_266);
and U615 (N_615,N_357,In_2399);
and U616 (N_616,In_1025,In_1278);
or U617 (N_617,N_198,In_1358);
xnor U618 (N_618,N_93,N_371);
nand U619 (N_619,In_2262,In_2786);
nand U620 (N_620,In_870,In_2805);
nor U621 (N_621,N_402,In_1178);
xnor U622 (N_622,In_1432,In_2070);
or U623 (N_623,In_2286,In_2832);
nand U624 (N_624,N_325,In_714);
or U625 (N_625,In_518,In_1810);
xnor U626 (N_626,In_373,In_1347);
xnor U627 (N_627,In_312,N_410);
and U628 (N_628,In_1006,In_21);
or U629 (N_629,In_1772,In_1526);
xor U630 (N_630,N_149,In_2224);
and U631 (N_631,N_88,N_57);
nor U632 (N_632,In_2012,N_429);
nor U633 (N_633,In_455,In_1946);
or U634 (N_634,In_251,N_187);
and U635 (N_635,In_588,In_2984);
and U636 (N_636,N_237,In_2690);
nor U637 (N_637,In_1711,In_1407);
nand U638 (N_638,In_1570,In_49);
nor U639 (N_639,N_486,In_1482);
and U640 (N_640,In_1721,In_1992);
nor U641 (N_641,In_2637,In_737);
xnor U642 (N_642,In_2946,In_2528);
and U643 (N_643,In_1053,In_2000);
and U644 (N_644,In_2025,In_2725);
xor U645 (N_645,In_2493,In_1729);
nor U646 (N_646,In_205,In_2785);
xor U647 (N_647,In_1847,In_1629);
xor U648 (N_648,In_921,In_359);
and U649 (N_649,In_126,In_2837);
nand U650 (N_650,In_1136,N_121);
nand U651 (N_651,In_1842,In_2333);
or U652 (N_652,In_762,N_457);
nand U653 (N_653,In_207,In_2423);
nor U654 (N_654,In_39,In_2102);
xnor U655 (N_655,In_2343,N_393);
xor U656 (N_656,In_1165,N_152);
nor U657 (N_657,In_201,In_182);
nand U658 (N_658,In_252,N_12);
nand U659 (N_659,In_1458,In_2222);
xor U660 (N_660,In_313,N_480);
xor U661 (N_661,N_86,N_157);
xor U662 (N_662,In_188,In_1109);
xnor U663 (N_663,In_2178,In_2073);
or U664 (N_664,In_1834,In_2264);
xor U665 (N_665,In_2524,In_2157);
or U666 (N_666,In_1528,In_2246);
and U667 (N_667,In_2612,N_87);
or U668 (N_668,N_32,In_2226);
xor U669 (N_669,In_2680,In_852);
nand U670 (N_670,In_2103,In_874);
nand U671 (N_671,In_688,In_2892);
or U672 (N_672,In_1701,In_2158);
or U673 (N_673,In_1083,N_469);
nand U674 (N_674,In_529,In_1515);
or U675 (N_675,In_2757,In_2702);
nor U676 (N_676,In_285,N_481);
nor U677 (N_677,N_353,In_406);
xnor U678 (N_678,In_2615,In_204);
and U679 (N_679,In_195,In_2173);
nand U680 (N_680,In_2796,N_386);
and U681 (N_681,In_1386,In_1882);
or U682 (N_682,In_2241,In_2512);
or U683 (N_683,In_114,N_196);
and U684 (N_684,In_175,In_2098);
nand U685 (N_685,In_1909,In_2450);
xor U686 (N_686,In_710,N_29);
and U687 (N_687,In_1402,N_456);
nand U688 (N_688,In_255,In_783);
nor U689 (N_689,N_82,In_2529);
and U690 (N_690,In_1277,In_2804);
nor U691 (N_691,In_2016,In_618);
and U692 (N_692,In_1303,In_2768);
and U693 (N_693,N_130,In_801);
nand U694 (N_694,In_2210,In_2864);
xnor U695 (N_695,In_2463,In_2385);
nor U696 (N_696,In_2436,In_1266);
nand U697 (N_697,In_2688,In_2151);
or U698 (N_698,In_514,In_178);
nor U699 (N_699,In_1030,In_2645);
xor U700 (N_700,N_246,In_817);
and U701 (N_701,In_69,In_1831);
or U702 (N_702,In_2541,In_2030);
nand U703 (N_703,In_2570,In_1497);
and U704 (N_704,In_1587,In_1143);
nor U705 (N_705,In_2032,In_137);
or U706 (N_706,In_2954,In_1785);
nand U707 (N_707,In_2432,In_1669);
and U708 (N_708,N_219,In_1758);
nor U709 (N_709,In_2492,N_223);
or U710 (N_710,In_1805,In_2448);
nand U711 (N_711,In_2909,In_1734);
xnor U712 (N_712,N_272,In_23);
nand U713 (N_713,In_1392,In_706);
nand U714 (N_714,N_364,In_2144);
and U715 (N_715,In_2371,In_411);
xor U716 (N_716,N_466,N_331);
nand U717 (N_717,In_2716,In_2774);
nor U718 (N_718,In_1297,In_1890);
nand U719 (N_719,In_1749,In_1863);
xnor U720 (N_720,N_199,In_906);
nor U721 (N_721,N_14,In_1445);
or U722 (N_722,N_40,In_2536);
nand U723 (N_723,In_369,N_230);
nor U724 (N_724,In_2390,In_730);
nor U725 (N_725,In_2926,In_1949);
nor U726 (N_726,In_2147,In_2712);
and U727 (N_727,In_2915,In_2278);
nor U728 (N_728,In_1096,In_519);
xnor U729 (N_729,In_278,In_2486);
or U730 (N_730,In_1607,N_359);
or U731 (N_731,N_205,N_228);
xnor U732 (N_732,N_73,In_456);
xnor U733 (N_733,In_2781,N_137);
and U734 (N_734,In_0,N_401);
nor U735 (N_735,In_2596,In_159);
nor U736 (N_736,N_379,In_1874);
nand U737 (N_737,In_1766,In_2840);
and U738 (N_738,In_319,In_943);
nand U739 (N_739,In_1420,N_69);
xnor U740 (N_740,In_1879,In_929);
and U741 (N_741,N_107,In_2607);
and U742 (N_742,In_1635,In_1955);
or U743 (N_743,In_2290,In_2109);
nor U744 (N_744,In_2296,N_350);
nor U745 (N_745,In_1002,In_693);
or U746 (N_746,In_1801,In_2752);
and U747 (N_747,In_1457,N_283);
nor U748 (N_748,In_1777,In_2407);
xnor U749 (N_749,In_615,In_370);
nand U750 (N_750,In_1491,N_204);
nand U751 (N_751,In_2233,In_1567);
nand U752 (N_752,In_1309,In_2267);
xnor U753 (N_753,In_1720,N_321);
and U754 (N_754,In_1104,In_1376);
nand U755 (N_755,In_1850,In_2216);
nor U756 (N_756,In_2256,In_2655);
nand U757 (N_757,In_1438,In_1135);
nand U758 (N_758,In_2628,In_1681);
or U759 (N_759,In_2606,In_962);
xor U760 (N_760,In_1944,In_520);
or U761 (N_761,In_2252,In_256);
nor U762 (N_762,In_2115,In_1430);
or U763 (N_763,In_477,In_644);
xor U764 (N_764,In_1216,In_2162);
xnor U765 (N_765,In_2452,N_376);
nor U766 (N_766,In_304,In_1017);
and U767 (N_767,In_635,In_1764);
nor U768 (N_768,In_1918,N_280);
nor U769 (N_769,N_239,In_2488);
xor U770 (N_770,In_2250,In_1325);
or U771 (N_771,In_1144,In_2411);
and U772 (N_772,In_613,In_2179);
xnor U773 (N_773,In_1557,In_2831);
xnor U774 (N_774,In_2515,In_2625);
xor U775 (N_775,In_729,In_2903);
and U776 (N_776,N_492,In_2975);
nor U777 (N_777,N_42,In_1612);
or U778 (N_778,N_344,N_349);
nor U779 (N_779,In_174,In_949);
and U780 (N_780,In_975,In_1383);
xnor U781 (N_781,In_2260,In_60);
and U782 (N_782,In_1703,In_2848);
nor U783 (N_783,In_1205,N_263);
nor U784 (N_784,In_908,In_1816);
or U785 (N_785,In_150,In_2213);
nand U786 (N_786,In_1296,In_1553);
nor U787 (N_787,In_1354,In_36);
nor U788 (N_788,N_59,In_16);
nor U789 (N_789,In_1525,In_2305);
or U790 (N_790,In_1189,In_276);
nand U791 (N_791,In_2744,In_616);
xor U792 (N_792,N_46,N_78);
xnor U793 (N_793,In_983,In_2314);
or U794 (N_794,In_2273,In_1582);
or U795 (N_795,In_1226,In_2519);
xor U796 (N_796,In_2682,In_1111);
nand U797 (N_797,In_86,In_2236);
xnor U798 (N_798,In_2500,In_2002);
nand U799 (N_799,In_210,In_2884);
nor U800 (N_800,N_339,N_124);
or U801 (N_801,In_2021,In_97);
or U802 (N_802,In_680,In_1122);
or U803 (N_803,In_1043,In_249);
and U804 (N_804,N_209,N_295);
and U805 (N_805,In_1770,In_402);
nand U806 (N_806,In_1527,In_2366);
and U807 (N_807,N_229,N_278);
or U808 (N_808,In_107,In_1859);
or U809 (N_809,In_2288,In_1973);
or U810 (N_810,In_678,In_968);
or U811 (N_811,In_1546,In_1878);
or U812 (N_812,In_2745,In_1033);
or U813 (N_813,In_2299,In_2936);
nor U814 (N_814,N_244,In_1687);
nor U815 (N_815,In_736,In_1012);
xnor U816 (N_816,In_345,In_397);
or U817 (N_817,In_969,In_1428);
xor U818 (N_818,In_442,In_1381);
and U819 (N_819,In_865,In_2047);
nor U820 (N_820,In_1710,In_1314);
nand U821 (N_821,N_118,In_587);
nor U822 (N_822,In_1864,N_143);
and U823 (N_823,In_859,N_166);
and U824 (N_824,In_2244,In_897);
nor U825 (N_825,In_1090,N_439);
nor U826 (N_826,In_2777,In_1322);
nand U827 (N_827,In_2583,N_221);
xor U828 (N_828,In_537,N_432);
and U829 (N_829,In_2124,In_1821);
and U830 (N_830,In_446,In_2283);
xor U831 (N_831,N_375,In_1436);
nand U832 (N_832,In_1804,In_305);
nor U833 (N_833,In_1116,In_1073);
or U834 (N_834,In_1091,In_1477);
and U835 (N_835,N_358,In_1323);
xnor U836 (N_836,N_154,In_2925);
and U837 (N_837,In_2727,In_2721);
nand U838 (N_838,In_1697,In_2459);
nand U839 (N_839,In_1085,N_225);
or U840 (N_840,In_1032,N_395);
xor U841 (N_841,In_1260,In_2243);
nand U842 (N_842,In_2382,In_1120);
nor U843 (N_843,In_2656,In_1441);
nor U844 (N_844,In_1545,In_311);
nand U845 (N_845,In_147,In_1093);
xnor U846 (N_846,In_1707,N_474);
or U847 (N_847,In_992,In_2771);
and U848 (N_848,N_227,In_552);
xor U849 (N_849,In_2907,In_268);
and U850 (N_850,In_2970,In_1220);
xor U851 (N_851,In_1976,N_110);
and U852 (N_852,In_559,N_214);
or U853 (N_853,In_1076,In_561);
and U854 (N_854,In_2185,In_2293);
nor U855 (N_855,In_440,In_2923);
nor U856 (N_856,In_2365,In_1046);
and U857 (N_857,In_2356,In_55);
or U858 (N_858,In_1513,In_1737);
nand U859 (N_859,N_471,In_919);
or U860 (N_860,In_1276,In_2396);
and U861 (N_861,In_646,In_2123);
and U862 (N_862,In_99,In_2871);
or U863 (N_863,In_2902,In_1298);
nand U864 (N_864,In_1846,In_141);
and U865 (N_865,In_2231,In_2164);
or U866 (N_866,In_727,In_2974);
xor U867 (N_867,In_2644,In_1505);
nor U868 (N_868,In_2381,N_328);
nor U869 (N_869,In_2301,In_1119);
or U870 (N_870,In_746,In_545);
or U871 (N_871,In_1072,In_2700);
nand U872 (N_872,In_108,In_1787);
nand U873 (N_873,In_2126,In_273);
nor U874 (N_874,In_2197,In_660);
and U875 (N_875,In_2556,N_265);
xor U876 (N_876,In_533,N_460);
nand U877 (N_877,In_1473,In_648);
or U878 (N_878,N_498,N_160);
xnor U879 (N_879,In_2955,In_2886);
or U880 (N_880,In_828,In_158);
xnor U881 (N_881,N_282,In_1328);
nand U882 (N_882,In_907,In_1994);
or U883 (N_883,In_2876,In_1680);
xnor U884 (N_884,In_1422,In_2188);
nor U885 (N_885,In_1267,In_53);
or U886 (N_886,In_1071,In_2368);
nor U887 (N_887,In_1103,In_1380);
xor U888 (N_888,In_1455,N_355);
xor U889 (N_889,In_392,In_318);
or U890 (N_890,In_704,In_1752);
nand U891 (N_891,In_1069,In_1644);
nor U892 (N_892,In_1599,In_348);
nor U893 (N_893,In_1833,In_781);
nor U894 (N_894,In_2113,N_377);
xnor U895 (N_895,In_474,In_643);
nand U896 (N_896,In_2443,In_2391);
or U897 (N_897,In_2873,In_2776);
and U898 (N_898,In_2362,In_2478);
nor U899 (N_899,In_531,In_1242);
and U900 (N_900,N_195,In_525);
nand U901 (N_901,In_2150,N_341);
nand U902 (N_902,In_2585,In_607);
and U903 (N_903,In_2865,In_2501);
xor U904 (N_904,N_92,N_165);
xnor U905 (N_905,In_690,In_1786);
and U906 (N_906,In_1549,In_1844);
xor U907 (N_907,In_1583,In_1427);
and U908 (N_908,In_1157,In_386);
nand U909 (N_909,In_1461,N_22);
and U910 (N_910,In_1746,N_269);
or U911 (N_911,In_1261,N_161);
nor U912 (N_912,In_1885,In_156);
nand U913 (N_913,N_28,In_189);
xor U914 (N_914,In_1410,In_508);
nor U915 (N_915,In_2859,In_793);
nand U916 (N_916,In_2398,In_2532);
and U917 (N_917,In_2174,N_472);
xnor U918 (N_918,N_430,N_414);
and U919 (N_919,In_2263,In_2350);
and U920 (N_920,N_425,In_129);
or U921 (N_921,In_2951,In_2590);
or U922 (N_922,N_458,In_2801);
and U923 (N_923,In_1611,In_2762);
and U924 (N_924,In_1472,In_2993);
and U925 (N_925,In_1097,In_244);
nand U926 (N_926,In_2274,In_1253);
nand U927 (N_927,N_312,In_798);
xor U928 (N_928,In_2300,In_1727);
xor U929 (N_929,In_2442,N_15);
xor U930 (N_930,In_1849,N_258);
nor U931 (N_931,In_1597,In_179);
and U932 (N_932,In_937,In_857);
or U933 (N_933,In_2522,In_2019);
or U934 (N_934,In_981,In_2896);
and U935 (N_935,In_1198,In_1164);
or U936 (N_936,In_1460,In_2739);
xnor U937 (N_937,In_2717,In_1232);
or U938 (N_938,In_866,In_2253);
nand U939 (N_939,In_96,In_1465);
nand U940 (N_940,N_394,In_724);
or U941 (N_941,In_2018,N_288);
and U942 (N_942,In_2475,N_268);
or U943 (N_943,N_257,N_97);
nand U944 (N_944,In_1501,N_172);
nand U945 (N_945,In_659,In_1080);
and U946 (N_946,N_254,In_2189);
nand U947 (N_947,N_277,In_540);
or U948 (N_948,N_365,N_61);
xor U949 (N_949,In_2767,In_2466);
nand U950 (N_950,N_48,In_486);
xor U951 (N_951,In_534,In_441);
and U952 (N_952,In_142,In_260);
nand U953 (N_953,In_2050,In_2920);
or U954 (N_954,In_2511,N_109);
and U955 (N_955,In_2042,In_1214);
and U956 (N_956,In_2736,In_2991);
and U957 (N_957,In_426,N_184);
and U958 (N_958,In_2325,N_153);
and U959 (N_959,N_419,In_1099);
xor U960 (N_960,N_286,In_337);
xnor U961 (N_961,In_110,In_941);
or U962 (N_962,N_302,In_57);
xor U963 (N_963,In_2457,N_178);
nand U964 (N_964,In_1803,In_2806);
xor U965 (N_965,In_2713,In_1280);
xor U966 (N_966,In_2654,N_405);
nand U967 (N_967,In_600,In_903);
nor U968 (N_968,In_1579,N_293);
nor U969 (N_969,In_2302,In_2895);
xor U970 (N_970,N_335,In_2678);
or U971 (N_971,In_2054,N_235);
nand U972 (N_972,In_702,In_272);
nor U973 (N_973,In_924,In_1660);
and U974 (N_974,In_2441,In_2088);
nand U975 (N_975,In_2387,In_1884);
and U976 (N_976,In_1823,In_2017);
or U977 (N_977,In_989,In_683);
xor U978 (N_978,In_896,N_403);
and U979 (N_979,In_1941,In_415);
or U980 (N_980,N_188,In_1393);
xnor U981 (N_981,In_2914,In_2026);
nand U982 (N_982,In_524,In_1107);
xnor U983 (N_983,In_2089,In_166);
nand U984 (N_984,In_122,In_990);
xor U985 (N_985,In_1338,In_111);
and U986 (N_986,In_2092,In_1044);
nor U987 (N_987,In_945,In_2666);
nor U988 (N_988,In_1056,In_2447);
xor U989 (N_989,In_2303,In_1838);
and U990 (N_990,In_1990,In_1784);
and U991 (N_991,In_1047,In_136);
or U992 (N_992,N_191,In_12);
and U993 (N_993,In_462,In_2693);
nor U994 (N_994,In_1409,In_2962);
and U995 (N_995,In_1153,In_2027);
and U996 (N_996,In_2561,In_428);
nor U997 (N_997,In_194,In_1695);
and U998 (N_998,N_361,In_2138);
or U999 (N_999,In_2176,In_2835);
nor U1000 (N_1000,N_804,In_2480);
xor U1001 (N_1001,N_763,In_451);
and U1002 (N_1002,N_488,In_102);
xor U1003 (N_1003,N_973,N_138);
and U1004 (N_1004,N_544,In_2604);
nand U1005 (N_1005,In_286,N_827);
or U1006 (N_1006,N_600,N_318);
xnor U1007 (N_1007,N_959,In_1705);
and U1008 (N_1008,In_2039,In_2632);
xnor U1009 (N_1009,In_2180,In_2171);
and U1010 (N_1010,In_1824,In_696);
nor U1011 (N_1011,In_2668,N_559);
nor U1012 (N_1012,In_829,In_2627);
or U1013 (N_1013,N_853,In_1776);
nor U1014 (N_1014,N_686,N_796);
xnor U1015 (N_1015,In_1341,N_289);
or U1016 (N_1016,In_2641,N_850);
nor U1017 (N_1017,In_2800,N_974);
nor U1018 (N_1018,N_433,N_108);
nand U1019 (N_1019,In_2956,In_716);
nand U1020 (N_1020,In_1330,In_2401);
nand U1021 (N_1021,N_803,N_764);
xor U1022 (N_1022,N_612,In_423);
and U1023 (N_1023,In_2006,N_666);
nor U1024 (N_1024,N_176,N_524);
or U1025 (N_1025,N_327,N_554);
nor U1026 (N_1026,N_884,N_636);
nand U1027 (N_1027,N_928,N_580);
nor U1028 (N_1028,N_505,N_482);
nor U1029 (N_1029,In_184,In_45);
and U1030 (N_1030,In_728,In_1372);
xnor U1031 (N_1031,In_2003,N_816);
and U1032 (N_1032,N_533,In_862);
nor U1033 (N_1033,In_134,N_383);
and U1034 (N_1034,N_232,N_839);
nor U1035 (N_1035,In_1709,In_2661);
xor U1036 (N_1036,In_2675,In_1487);
nor U1037 (N_1037,N_951,In_227);
nand U1038 (N_1038,In_1914,N_728);
xnor U1039 (N_1039,In_1152,In_1019);
and U1040 (N_1040,N_427,In_186);
nor U1041 (N_1041,N_872,In_800);
and U1042 (N_1042,In_2897,In_215);
and U1043 (N_1043,N_210,In_623);
or U1044 (N_1044,In_889,N_91);
nand U1045 (N_1045,N_864,N_445);
nand U1046 (N_1046,In_2833,In_1265);
and U1047 (N_1047,In_784,In_1105);
or U1048 (N_1048,N_942,In_2764);
xor U1049 (N_1049,N_813,In_2810);
and U1050 (N_1050,N_876,N_593);
xnor U1051 (N_1051,N_780,N_496);
or U1052 (N_1052,N_512,In_1334);
xnor U1053 (N_1053,In_687,N_743);
and U1054 (N_1054,N_597,N_865);
nand U1055 (N_1055,N_236,N_628);
or U1056 (N_1056,N_880,In_2924);
nor U1057 (N_1057,In_1671,In_2022);
nor U1058 (N_1058,In_2653,In_2077);
nand U1059 (N_1059,In_1790,In_1664);
nor U1060 (N_1060,In_1581,In_2662);
nor U1061 (N_1061,In_1156,In_2108);
nand U1062 (N_1062,N_506,In_1448);
nor U1063 (N_1063,In_957,In_282);
nor U1064 (N_1064,In_1169,In_665);
xor U1065 (N_1065,In_1236,In_1485);
nor U1066 (N_1066,In_708,In_2094);
or U1067 (N_1067,In_1498,In_1348);
nor U1068 (N_1068,In_2354,N_464);
nand U1069 (N_1069,In_270,N_182);
or U1070 (N_1070,N_950,N_452);
nand U1071 (N_1071,In_2797,In_2683);
nor U1072 (N_1072,N_777,In_2251);
nand U1073 (N_1073,N_285,In_1639);
and U1074 (N_1074,In_140,In_652);
nand U1075 (N_1075,In_663,In_1502);
or U1076 (N_1076,In_1933,N_55);
nand U1077 (N_1077,In_2588,In_599);
or U1078 (N_1078,In_2207,N_72);
or U1079 (N_1079,N_787,In_1173);
nand U1080 (N_1080,In_2292,In_1641);
nand U1081 (N_1081,N_25,In_120);
nor U1082 (N_1082,In_1954,In_2930);
xnor U1083 (N_1083,In_899,N_64);
xor U1084 (N_1084,N_317,N_737);
or U1085 (N_1085,In_420,N_33);
and U1086 (N_1086,In_2545,N_446);
nand U1087 (N_1087,In_496,N_535);
and U1088 (N_1088,In_946,N_851);
nor U1089 (N_1089,N_961,In_1563);
xnor U1090 (N_1090,In_1094,In_2631);
nor U1091 (N_1091,N_841,In_2879);
nor U1092 (N_1092,N_627,N_650);
or U1093 (N_1093,N_795,In_1614);
nor U1094 (N_1094,In_2894,In_2773);
nor U1095 (N_1095,N_49,N_490);
nand U1096 (N_1096,In_155,In_535);
and U1097 (N_1097,N_382,N_461);
or U1098 (N_1098,N_212,N_943);
nand U1099 (N_1099,In_1530,In_253);
or U1100 (N_1100,In_7,N_776);
nor U1101 (N_1101,In_2496,In_192);
xnor U1102 (N_1102,N_882,N_447);
nor U1103 (N_1103,N_731,N_870);
or U1104 (N_1104,In_1040,N_908);
xor U1105 (N_1105,N_329,In_1036);
nor U1106 (N_1106,In_2748,In_1462);
nor U1107 (N_1107,In_2045,N_769);
xnor U1108 (N_1108,In_2782,In_2746);
xor U1109 (N_1109,N_774,In_1426);
xor U1110 (N_1110,N_833,N_681);
xnor U1111 (N_1111,In_573,N_805);
nor U1112 (N_1112,N_575,In_894);
xor U1113 (N_1113,In_1295,In_59);
or U1114 (N_1114,N_760,N_745);
xnor U1115 (N_1115,N_248,N_4);
xor U1116 (N_1116,In_448,N_563);
or U1117 (N_1117,In_470,In_1608);
xor U1118 (N_1118,In_2787,N_333);
xor U1119 (N_1119,In_2204,N_698);
nand U1120 (N_1120,In_1062,N_832);
or U1121 (N_1121,N_296,In_2454);
nand U1122 (N_1122,N_638,In_2862);
and U1123 (N_1123,In_261,In_62);
and U1124 (N_1124,N_685,N_381);
or U1125 (N_1125,In_1636,In_247);
nand U1126 (N_1126,In_1418,N_955);
nand U1127 (N_1127,N_68,N_242);
nand U1128 (N_1128,N_459,In_2514);
and U1129 (N_1129,In_1182,In_2360);
nor U1130 (N_1130,In_2058,In_109);
or U1131 (N_1131,N_556,In_2215);
xor U1132 (N_1132,In_2166,N_292);
and U1133 (N_1133,In_1595,N_949);
or U1134 (N_1134,In_71,In_1279);
and U1135 (N_1135,N_977,N_674);
and U1136 (N_1136,N_799,In_847);
nand U1137 (N_1137,In_2617,In_1160);
and U1138 (N_1138,In_382,In_987);
xor U1139 (N_1139,In_1550,In_2490);
nor U1140 (N_1140,N_699,In_356);
nand U1141 (N_1141,N_792,N_794);
nand U1142 (N_1142,N_798,In_656);
nand U1143 (N_1143,In_1555,In_151);
or U1144 (N_1144,In_1374,N_418);
nor U1145 (N_1145,In_846,In_940);
nor U1146 (N_1146,In_2921,N_704);
xnor U1147 (N_1147,In_1403,N_347);
or U1148 (N_1148,N_608,In_1731);
nor U1149 (N_1149,In_190,N_967);
nand U1150 (N_1150,N_661,In_46);
or U1151 (N_1151,In_1051,N_276);
and U1152 (N_1152,In_1974,In_1931);
xnor U1153 (N_1153,In_347,In_2537);
nor U1154 (N_1154,N_590,N_979);
or U1155 (N_1155,In_2815,In_30);
nand U1156 (N_1156,In_2494,In_827);
xor U1157 (N_1157,In_770,In_2506);
and U1158 (N_1158,In_1714,N_75);
nand U1159 (N_1159,N_818,In_697);
or U1160 (N_1160,N_105,N_702);
and U1161 (N_1161,N_915,In_2259);
nand U1162 (N_1162,In_1484,In_849);
or U1163 (N_1163,N_255,In_629);
nor U1164 (N_1164,In_709,In_447);
nand U1165 (N_1165,In_2803,In_424);
xnor U1166 (N_1166,In_575,N_500);
xnor U1167 (N_1167,In_1657,In_2351);
or U1168 (N_1168,N_66,In_2277);
xnor U1169 (N_1169,N_513,N_709);
nor U1170 (N_1170,N_782,In_2295);
and U1171 (N_1171,In_2619,N_985);
or U1172 (N_1172,In_885,N_747);
or U1173 (N_1173,In_2811,In_1603);
nor U1174 (N_1174,In_1048,In_608);
nor U1175 (N_1175,N_356,N_483);
nor U1176 (N_1176,In_35,N_680);
and U1177 (N_1177,N_536,N_718);
and U1178 (N_1178,N_588,In_550);
xnor U1179 (N_1179,In_1899,In_2429);
and U1180 (N_1180,In_831,N_494);
and U1181 (N_1181,N_582,N_643);
nor U1182 (N_1182,In_631,In_1971);
and U1183 (N_1183,In_2910,In_1174);
nor U1184 (N_1184,In_1940,N_523);
xnor U1185 (N_1185,N_502,In_1476);
xor U1186 (N_1186,In_2814,In_1208);
nand U1187 (N_1187,In_2195,N_220);
or U1188 (N_1188,In_2364,In_1604);
or U1189 (N_1189,In_1724,In_2091);
xnor U1190 (N_1190,N_3,N_633);
xor U1191 (N_1191,N_368,N_808);
xor U1192 (N_1192,N_883,In_494);
and U1193 (N_1193,In_1447,In_2467);
nand U1194 (N_1194,In_115,N_920);
nor U1195 (N_1195,N_203,N_290);
nor U1196 (N_1196,In_2908,N_442);
xor U1197 (N_1197,N_946,In_2214);
xor U1198 (N_1198,N_812,N_270);
nor U1199 (N_1199,N_304,In_387);
xnor U1200 (N_1200,In_1797,N_271);
nor U1201 (N_1201,In_1333,In_79);
or U1202 (N_1202,N_617,N_13);
xor U1203 (N_1203,N_960,In_349);
nand U1204 (N_1204,In_2422,In_1628);
nor U1205 (N_1205,In_960,N_622);
or U1206 (N_1206,N_904,N_262);
or U1207 (N_1207,In_703,In_748);
xor U1208 (N_1208,N_528,N_5);
or U1209 (N_1209,N_820,In_825);
nand U1210 (N_1210,N_81,In_1005);
or U1211 (N_1211,In_11,N_913);
nand U1212 (N_1212,In_2795,In_1895);
xor U1213 (N_1213,In_2392,N_930);
xor U1214 (N_1214,N_781,In_1022);
xor U1215 (N_1215,In_2580,In_350);
and U1216 (N_1216,In_472,In_985);
and U1217 (N_1217,N_8,N_119);
nand U1218 (N_1218,In_1620,N_931);
nand U1219 (N_1219,N_875,N_266);
or U1220 (N_1220,N_697,In_2035);
and U1221 (N_1221,In_157,N_420);
nand U1222 (N_1222,In_1512,In_726);
xor U1223 (N_1223,N_243,In_460);
xnor U1224 (N_1224,N_957,In_1271);
nor U1225 (N_1225,N_530,N_874);
nand U1226 (N_1226,In_2324,In_821);
nand U1227 (N_1227,In_2838,N_250);
nand U1228 (N_1228,In_1474,In_2183);
nor U1229 (N_1229,In_2249,N_260);
or U1230 (N_1230,N_390,N_707);
and U1231 (N_1231,In_1490,N_41);
and U1232 (N_1232,N_990,N_560);
or U1233 (N_1233,N_89,N_733);
nand U1234 (N_1234,N_937,In_2633);
nand U1235 (N_1235,N_969,In_2065);
nand U1236 (N_1236,In_1851,N_552);
or U1237 (N_1237,In_431,In_196);
nand U1238 (N_1238,In_292,N_95);
xnor U1239 (N_1239,N_367,N_542);
or U1240 (N_1240,N_37,In_1856);
and U1241 (N_1241,N_684,In_105);
or U1242 (N_1242,In_677,In_2673);
or U1243 (N_1243,In_1774,N_863);
nand U1244 (N_1244,N_303,In_1702);
and U1245 (N_1245,N_972,N_726);
and U1246 (N_1246,N_896,In_2067);
xor U1247 (N_1247,In_2332,N_10);
or U1248 (N_1248,N_315,In_1981);
or U1249 (N_1249,In_1897,In_87);
nor U1250 (N_1250,In_782,N_899);
nand U1251 (N_1251,N_877,In_1519);
xnor U1252 (N_1252,In_523,In_1133);
nor U1253 (N_1253,In_2425,N_256);
nor U1254 (N_1254,N_476,In_2465);
or U1255 (N_1255,In_180,In_911);
nand U1256 (N_1256,N_712,In_164);
nand U1257 (N_1257,N_35,N_706);
nand U1258 (N_1258,In_2798,In_586);
nor U1259 (N_1259,In_711,In_1843);
and U1260 (N_1260,N_635,N_840);
and U1261 (N_1261,In_772,In_1130);
nand U1262 (N_1262,In_258,In_112);
nand U1263 (N_1263,In_641,N_2);
nor U1264 (N_1264,N_922,N_789);
or U1265 (N_1265,In_1075,In_92);
nand U1266 (N_1266,N_507,N_842);
and U1267 (N_1267,In_1999,In_2794);
and U1268 (N_1268,In_1820,N_744);
xor U1269 (N_1269,In_185,N_676);
nor U1270 (N_1270,N_735,N_539);
nor U1271 (N_1271,N_802,In_1601);
and U1272 (N_1272,N_611,N_670);
xor U1273 (N_1273,N_591,N_895);
xnor U1274 (N_1274,N_294,In_583);
xor U1275 (N_1275,In_1321,N_655);
nand U1276 (N_1276,N_759,In_461);
nand U1277 (N_1277,In_879,N_604);
or U1278 (N_1278,In_58,N_595);
or U1279 (N_1279,N_573,N_598);
xnor U1280 (N_1280,N_44,In_684);
or U1281 (N_1281,In_2948,N_652);
nand U1282 (N_1282,In_2747,In_1258);
nand U1283 (N_1283,In_1907,In_64);
nor U1284 (N_1284,In_294,N_669);
or U1285 (N_1285,In_1231,In_211);
nor U1286 (N_1286,In_662,In_2193);
and U1287 (N_1287,In_2584,In_1145);
or U1288 (N_1288,N_547,N_868);
and U1289 (N_1289,N_846,N_836);
or U1290 (N_1290,In_816,N_800);
and U1291 (N_1291,In_562,In_2788);
xnor U1292 (N_1292,In_2304,In_1218);
nand U1293 (N_1293,In_2726,N_151);
nand U1294 (N_1294,In_2618,N_99);
nand U1295 (N_1295,N_996,In_913);
nand U1296 (N_1296,In_1281,In_2699);
or U1297 (N_1297,In_2591,N_692);
or U1298 (N_1298,In_1503,N_281);
nor U1299 (N_1299,N_775,N_284);
and U1300 (N_1300,In_1813,In_427);
and U1301 (N_1301,In_72,N_694);
xnor U1302 (N_1302,N_103,In_2355);
and U1303 (N_1303,In_570,In_1050);
nand U1304 (N_1304,In_37,In_986);
and U1305 (N_1305,In_585,In_2345);
nand U1306 (N_1306,N_114,In_1240);
or U1307 (N_1307,In_2461,N_311);
nand U1308 (N_1308,In_2,N_190);
nand U1309 (N_1309,In_1891,In_959);
and U1310 (N_1310,In_1311,In_760);
nor U1311 (N_1311,In_1416,N_847);
nand U1312 (N_1312,In_1285,In_2125);
and U1313 (N_1313,N_941,N_648);
nor U1314 (N_1314,N_437,In_2175);
and U1315 (N_1315,In_740,N_583);
nor U1316 (N_1316,In_839,In_203);
or U1317 (N_1317,In_1910,In_130);
or U1318 (N_1318,In_1394,In_2081);
nor U1319 (N_1319,N_202,In_1024);
nor U1320 (N_1320,N_806,In_2737);
nor U1321 (N_1321,In_2186,N_826);
and U1322 (N_1322,In_2715,In_1201);
xnor U1323 (N_1323,In_765,In_2057);
nor U1324 (N_1324,In_1900,In_1991);
or U1325 (N_1325,In_324,In_265);
and U1326 (N_1326,In_228,N_939);
or U1327 (N_1327,In_1817,In_234);
nand U1328 (N_1328,In_450,N_411);
or U1329 (N_1329,In_2397,In_2445);
xor U1330 (N_1330,In_2194,In_1488);
nand U1331 (N_1331,In_1429,In_1760);
or U1332 (N_1332,N_18,N_729);
xnor U1333 (N_1333,In_1373,In_1645);
or U1334 (N_1334,N_324,N_790);
nor U1335 (N_1335,N_332,In_2640);
and U1336 (N_1336,N_654,N_918);
nor U1337 (N_1337,In_479,In_363);
nand U1338 (N_1338,N_566,N_917);
and U1339 (N_1339,N_565,In_2313);
nor U1340 (N_1340,N_938,N_786);
or U1341 (N_1341,In_2918,N_784);
nor U1342 (N_1342,N_468,N_215);
xnor U1343 (N_1343,N_910,N_435);
xnor U1344 (N_1344,N_940,In_1796);
and U1345 (N_1345,N_678,In_2160);
nor U1346 (N_1346,In_2421,In_2140);
nand U1347 (N_1347,In_1743,N_298);
and U1348 (N_1348,In_2069,In_2882);
nor U1349 (N_1349,In_1937,In_2306);
and U1350 (N_1350,N_634,In_2756);
xnor U1351 (N_1351,In_1306,In_1399);
xor U1352 (N_1352,N_319,In_66);
nand U1353 (N_1353,In_2223,In_2412);
or U1354 (N_1354,In_976,N_703);
or U1355 (N_1355,In_1948,In_17);
nand U1356 (N_1356,In_421,N_463);
or U1357 (N_1357,In_138,N_965);
nor U1358 (N_1358,In_1571,In_248);
or U1359 (N_1359,In_883,In_153);
nor U1360 (N_1360,N_642,In_1483);
xor U1361 (N_1361,N_21,N_185);
or U1362 (N_1362,In_284,In_1670);
and U1363 (N_1363,N_300,In_478);
and U1364 (N_1364,In_1041,N_343);
nand U1365 (N_1365,In_1713,In_2969);
nand U1366 (N_1366,In_245,In_2220);
and U1367 (N_1367,In_719,In_2790);
or U1368 (N_1368,N_935,In_1471);
and U1369 (N_1369,In_1168,N_881);
nand U1370 (N_1370,In_1305,In_1496);
and U1371 (N_1371,N_336,In_2234);
or U1372 (N_1372,N_519,In_2789);
and U1373 (N_1373,In_176,In_1037);
and U1374 (N_1374,In_1274,In_991);
or U1375 (N_1375,N_671,N_690);
and U1376 (N_1376,In_2589,In_2979);
xnor U1377 (N_1377,N_609,N_587);
and U1378 (N_1378,In_790,N_129);
or U1379 (N_1379,N_785,N_467);
nor U1380 (N_1380,N_56,In_1529);
nand U1381 (N_1381,In_880,In_578);
or U1382 (N_1382,N_102,In_1049);
nand U1383 (N_1383,N_879,N_128);
xor U1384 (N_1384,In_1176,N_51);
or U1385 (N_1385,N_952,N_106);
xor U1386 (N_1386,N_462,In_2547);
xnor U1387 (N_1387,N_663,In_820);
xnor U1388 (N_1388,N_17,In_2911);
or U1389 (N_1389,In_2409,In_636);
and U1390 (N_1390,In_1568,In_355);
or U1391 (N_1391,In_497,In_1854);
nor U1392 (N_1392,In_872,N_660);
and U1393 (N_1393,N_695,N_948);
nor U1394 (N_1394,In_574,N_742);
xnor U1395 (N_1395,N_451,N_520);
xnor U1396 (N_1396,N_993,N_120);
nor U1397 (N_1397,In_1957,In_181);
nand U1398 (N_1398,N_163,In_2995);
and U1399 (N_1399,In_2120,N_619);
nand U1400 (N_1400,In_1659,In_2958);
and U1401 (N_1401,In_2388,In_208);
or U1402 (N_1402,N_825,In_1747);
xor U1403 (N_1403,In_836,In_2435);
nor U1404 (N_1404,N_810,N_779);
nor U1405 (N_1405,N_645,In_1572);
nand U1406 (N_1406,N_174,In_2660);
nor U1407 (N_1407,N_814,N_987);
and U1408 (N_1408,N_892,N_388);
xor U1409 (N_1409,In_473,N_180);
and U1410 (N_1410,In_2947,In_2072);
xnor U1411 (N_1411,N_123,N_407);
or U1412 (N_1412,In_2642,N_52);
and U1413 (N_1413,N_578,N_629);
nor U1414 (N_1414,N_857,In_974);
xor U1415 (N_1415,In_843,In_2944);
nand U1416 (N_1416,In_2812,N_834);
or U1417 (N_1417,In_2078,In_1167);
and U1418 (N_1418,N_576,In_1249);
nand U1419 (N_1419,In_1349,N_501);
xor U1420 (N_1420,N_926,In_1434);
or U1421 (N_1421,N_249,In_2609);
or U1422 (N_1422,In_1141,In_2957);
or U1423 (N_1423,N_94,N_936);
and U1424 (N_1424,N_54,N_337);
nand U1425 (N_1425,In_2361,N_475);
xor U1426 (N_1426,In_1481,N_104);
and U1427 (N_1427,In_2887,In_2334);
xor U1428 (N_1428,In_1543,In_388);
xnor U1429 (N_1429,N_537,In_1365);
nor U1430 (N_1430,N_738,In_2750);
or U1431 (N_1431,N_351,In_509);
and U1432 (N_1432,N_646,In_624);
and U1433 (N_1433,In_1761,In_2572);
xor U1434 (N_1434,N_772,In_308);
nor U1435 (N_1435,N_701,In_1715);
nor U1436 (N_1436,In_2010,N_756);
and U1437 (N_1437,In_1959,In_1825);
xnor U1438 (N_1438,In_2885,In_1351);
nand U1439 (N_1439,N_444,N_6);
or U1440 (N_1440,N_168,N_38);
and U1441 (N_1441,N_473,N_264);
xnor U1442 (N_1442,In_322,N_201);
nor U1443 (N_1443,In_2953,N_891);
xor U1444 (N_1444,N_326,N_724);
xor U1445 (N_1445,In_254,In_1257);
nand U1446 (N_1446,In_2933,In_814);
nor U1447 (N_1447,N_529,In_2516);
and U1448 (N_1448,In_198,In_1996);
and U1449 (N_1449,In_1617,In_2375);
and U1450 (N_1450,In_2710,In_1262);
nand U1451 (N_1451,N_231,In_2509);
or U1452 (N_1452,In_167,In_1798);
and U1453 (N_1453,N_181,N_297);
xor U1454 (N_1454,In_1356,In_2775);
nor U1455 (N_1455,In_1716,In_403);
nand U1456 (N_1456,N_139,N_9);
or U1457 (N_1457,In_778,In_947);
and U1458 (N_1458,N_887,N_252);
nand U1459 (N_1459,In_2573,In_1675);
xnor U1460 (N_1460,In_225,In_2996);
nand U1461 (N_1461,In_2731,N_60);
xnor U1462 (N_1462,N_391,N_569);
xor U1463 (N_1463,In_1326,In_1263);
nor U1464 (N_1464,N_24,In_1387);
or U1465 (N_1465,N_396,In_1997);
or U1466 (N_1466,N_531,N_200);
xor U1467 (N_1467,N_416,N_131);
nor U1468 (N_1468,N_534,In_922);
and U1469 (N_1469,In_1780,In_1127);
and U1470 (N_1470,N_888,N_912);
and U1471 (N_1471,In_1095,N_354);
or U1472 (N_1472,N_553,N_797);
xnor U1473 (N_1473,In_1029,In_2539);
nor U1474 (N_1474,N_783,N_434);
nor U1475 (N_1475,In_469,N_599);
or U1476 (N_1476,In_1578,In_1255);
nand U1477 (N_1477,N_36,N_171);
or U1478 (N_1478,N_761,N_150);
nor U1479 (N_1479,In_2001,N_392);
nand U1480 (N_1480,In_2505,N_549);
xnor U1481 (N_1481,In_2199,In_513);
nand U1482 (N_1482,N_830,In_1606);
nand U1483 (N_1483,N_992,In_1674);
xnor U1484 (N_1484,In_563,N_426);
and U1485 (N_1485,N_594,In_901);
xnor U1486 (N_1486,N_871,In_1014);
xor U1487 (N_1487,N_510,In_594);
nor U1488 (N_1488,In_2934,N_71);
and U1489 (N_1489,In_1908,In_2904);
nand U1490 (N_1490,In_425,N_758);
or U1491 (N_1491,In_1121,In_6);
and U1492 (N_1492,N_767,In_1795);
and U1493 (N_1493,N_30,N_484);
and U1494 (N_1494,In_2822,N_241);
nor U1495 (N_1495,In_2959,In_963);
or U1496 (N_1496,In_1251,In_295);
and U1497 (N_1497,N_240,In_1548);
nor U1498 (N_1498,N_963,In_556);
nand U1499 (N_1499,In_2503,N_508);
xnor U1500 (N_1500,In_2913,In_38);
and U1501 (N_1501,N_1341,N_1244);
and U1502 (N_1502,N_1069,In_328);
xor U1503 (N_1503,In_2015,N_134);
and U1504 (N_1504,N_1183,In_1108);
and U1505 (N_1505,N_1430,N_144);
nor U1506 (N_1506,In_51,N_889);
nor U1507 (N_1507,N_1120,N_1235);
xor U1508 (N_1508,N_791,In_1312);
nand U1509 (N_1509,N_1106,N_1463);
xor U1510 (N_1510,N_1493,In_262);
and U1511 (N_1511,In_2770,N_1008);
xor U1512 (N_1512,In_1783,N_449);
nand U1513 (N_1513,In_2271,N_1323);
and U1514 (N_1514,In_1209,N_251);
or U1515 (N_1515,In_593,In_2127);
or U1516 (N_1516,In_1930,N_601);
or U1517 (N_1517,In_1979,In_695);
and U1518 (N_1518,N_869,N_1266);
or U1519 (N_1519,In_1463,N_1389);
or U1520 (N_1520,N_1337,N_521);
or U1521 (N_1521,In_2994,In_747);
xor U1522 (N_1522,In_2857,In_361);
nand U1523 (N_1523,N_765,In_2380);
nor U1524 (N_1524,N_141,N_148);
nand U1525 (N_1525,In_685,N_1422);
xor U1526 (N_1526,N_1275,N_736);
nor U1527 (N_1527,In_2420,In_1241);
or U1528 (N_1528,N_750,In_2285);
and U1529 (N_1529,In_2495,In_2799);
nor U1530 (N_1530,In_1562,In_1291);
and U1531 (N_1531,N_1078,In_1782);
or U1532 (N_1532,N_175,N_412);
xnor U1533 (N_1533,In_1993,N_1237);
xnor U1534 (N_1534,N_548,In_1179);
xnor U1535 (N_1535,In_1634,N_561);
nor U1536 (N_1536,In_647,In_376);
and U1537 (N_1537,N_1420,N_1233);
nand U1538 (N_1538,N_1461,In_2122);
xnor U1539 (N_1539,In_2111,N_664);
xor U1540 (N_1540,In_2378,In_1953);
or U1541 (N_1541,N_424,In_1989);
nand U1542 (N_1542,N_1425,N_603);
xnor U1543 (N_1543,N_1017,In_1110);
xnor U1544 (N_1544,In_1339,In_838);
and U1545 (N_1545,In_1802,N_1052);
or U1546 (N_1546,N_43,In_2992);
xor U1547 (N_1547,In_132,N_1381);
or U1548 (N_1548,N_1234,In_1008);
xnor U1549 (N_1549,In_2753,N_267);
nand U1550 (N_1550,N_1188,In_2845);
and U1551 (N_1551,In_1283,In_419);
or U1552 (N_1552,In_925,N_1159);
and U1553 (N_1553,N_1496,N_1334);
or U1554 (N_1554,In_2905,In_2440);
nand U1555 (N_1555,N_1391,N_1312);
and U1556 (N_1556,In_2484,N_1343);
xnor U1557 (N_1557,In_1866,In_2560);
or U1558 (N_1558,In_372,In_527);
nand U1559 (N_1559,N_934,N_532);
and U1560 (N_1560,In_1799,N_1190);
xor U1561 (N_1561,N_1221,N_1442);
or U1562 (N_1562,N_1260,N_1129);
and U1563 (N_1563,N_1113,N_1415);
nor U1564 (N_1564,N_665,N_1387);
and U1565 (N_1565,N_1492,In_2525);
or U1566 (N_1566,In_1194,In_1793);
nand U1567 (N_1567,In_239,N_1224);
nand U1568 (N_1568,N_1448,N_499);
and U1569 (N_1569,N_1038,In_2766);
nand U1570 (N_1570,N_721,N_316);
or U1571 (N_1571,In_2471,N_1390);
xnor U1572 (N_1572,In_1456,N_858);
nand U1573 (N_1573,In_1738,N_1451);
nor U1574 (N_1574,N_218,N_793);
xor U1575 (N_1575,N_1025,In_1125);
and U1576 (N_1576,N_1388,N_1024);
xnor U1577 (N_1577,N_305,In_763);
nand U1578 (N_1578,N_1377,N_616);
nor U1579 (N_1579,N_1403,In_187);
nor U1580 (N_1580,In_1769,N_373);
xnor U1581 (N_1581,N_672,In_2393);
nor U1582 (N_1582,N_606,N_980);
nor U1583 (N_1583,N_338,N_700);
nand U1584 (N_1584,N_551,In_2858);
or U1585 (N_1585,In_834,N_307);
nand U1586 (N_1586,N_1278,In_2275);
xor U1587 (N_1587,N_1319,N_1400);
nor U1588 (N_1588,N_164,N_831);
or U1589 (N_1589,In_1717,In_640);
xnor U1590 (N_1590,N_1444,N_1321);
xor U1591 (N_1591,N_1404,N_1373);
and U1592 (N_1592,N_757,In_826);
nand U1593 (N_1593,In_1459,N_1112);
and U1594 (N_1594,N_644,In_2817);
nor U1595 (N_1595,N_522,N_1070);
or U1596 (N_1596,N_1262,N_1481);
or U1597 (N_1597,N_727,In_2987);
or U1598 (N_1598,N_1124,N_1003);
nand U1599 (N_1599,N_862,In_1235);
nand U1600 (N_1600,N_807,In_2594);
xnor U1601 (N_1601,N_886,In_1317);
nand U1602 (N_1602,N_705,N_1097);
xnor U1603 (N_1603,N_1392,N_1145);
or U1604 (N_1604,N_1140,In_2156);
and U1605 (N_1605,N_1454,N_146);
and U1606 (N_1606,In_1054,N_156);
xnor U1607 (N_1607,N_1366,In_2980);
and U1608 (N_1608,In_642,In_1272);
nand U1609 (N_1609,In_48,N_567);
and U1610 (N_1610,N_1335,N_1193);
or U1611 (N_1611,N_788,In_2149);
xor U1612 (N_1612,N_1417,N_1280);
or U1613 (N_1613,N_1349,N_385);
and U1614 (N_1614,N_478,In_1134);
or U1615 (N_1615,In_1936,N_287);
xnor U1616 (N_1616,N_1303,In_2819);
xor U1617 (N_1617,In_512,N_1258);
nand U1618 (N_1618,N_746,In_139);
and U1619 (N_1619,In_1467,N_667);
nor U1620 (N_1620,N_809,N_1028);
nor U1621 (N_1621,N_1402,N_1302);
nand U1622 (N_1622,In_1511,N_1315);
xor U1623 (N_1623,N_725,N_1307);
xor U1624 (N_1624,N_1022,N_247);
or U1625 (N_1625,In_310,N_1111);
xor U1626 (N_1626,N_584,In_2418);
nor U1627 (N_1627,N_1206,N_1095);
or U1628 (N_1628,In_1010,N_1134);
or U1629 (N_1629,In_2639,N_1379);
nor U1630 (N_1630,In_998,In_1520);
nand U1631 (N_1631,N_404,In_1234);
nor U1632 (N_1632,N_179,N_995);
or U1633 (N_1633,In_498,N_1288);
nor U1634 (N_1634,N_1185,In_2049);
and U1635 (N_1635,N_1384,N_1346);
and U1636 (N_1636,N_852,In_1828);
nor U1637 (N_1637,In_2874,N_1220);
or U1638 (N_1638,In_2938,N_1245);
xor U1639 (N_1639,N_1181,N_878);
xor U1640 (N_1640,N_1453,N_454);
nand U1641 (N_1641,In_1741,N_1027);
and U1642 (N_1642,N_579,In_1609);
nand U1643 (N_1643,In_1650,N_662);
xnor U1644 (N_1644,In_1647,N_299);
nor U1645 (N_1645,In_408,N_222);
nand U1646 (N_1646,In_1301,N_614);
and U1647 (N_1647,N_1071,In_2408);
nor U1648 (N_1648,In_567,N_1178);
xor U1649 (N_1649,N_632,N_504);
or U1650 (N_1650,N_1058,N_1225);
nand U1651 (N_1651,In_2228,N_1248);
xnor U1652 (N_1652,N_1317,In_1943);
and U1653 (N_1653,In_2323,In_1185);
xnor U1654 (N_1654,N_1094,In_1558);
or U1655 (N_1655,N_1273,N_1470);
or U1656 (N_1656,In_98,N_1174);
nand U1657 (N_1657,In_236,In_1686);
or U1658 (N_1658,N_1267,N_1127);
nand U1659 (N_1659,N_1229,N_1401);
nand U1660 (N_1660,N_301,In_2326);
nor U1661 (N_1661,N_314,N_415);
nor U1662 (N_1662,N_417,N_1158);
nor U1663 (N_1663,In_2569,N_1155);
nor U1664 (N_1664,In_2315,N_194);
xor U1665 (N_1665,In_2972,In_466);
nand U1666 (N_1666,In_1531,N_1460);
nor U1667 (N_1667,N_916,In_2403);
xor U1668 (N_1668,N_956,N_525);
and U1669 (N_1669,N_1016,In_966);
and U1670 (N_1670,In_1346,In_604);
and U1671 (N_1671,N_493,In_413);
and U1672 (N_1672,N_1416,N_1298);
or U1673 (N_1673,In_667,N_1170);
or U1674 (N_1674,N_708,N_905);
nand U1675 (N_1675,N_274,In_2038);
nor U1676 (N_1676,In_213,N_866);
or U1677 (N_1677,N_1318,In_351);
nand U1678 (N_1678,N_516,In_2649);
xor U1679 (N_1679,N_1059,In_2557);
nand U1680 (N_1680,N_1057,In_1433);
nor U1681 (N_1681,In_1754,N_116);
xor U1682 (N_1682,N_1133,In_2587);
or U1683 (N_1683,N_766,N_1438);
nor U1684 (N_1684,In_2043,N_997);
or U1685 (N_1685,In_1554,N_637);
nand U1686 (N_1686,In_94,In_1117);
nor U1687 (N_1687,In_1504,In_672);
and U1688 (N_1688,N_526,N_1359);
xnor U1689 (N_1689,In_2780,In_536);
xnor U1690 (N_1690,N_1385,In_1928);
nand U1691 (N_1691,N_1396,N_1327);
nor U1692 (N_1692,In_538,N_423);
nor U1693 (N_1693,N_63,N_1279);
nand U1694 (N_1694,N_1072,In_371);
or U1695 (N_1695,N_749,N_1010);
or U1696 (N_1696,N_620,In_1632);
nand U1697 (N_1697,N_79,N_914);
nor U1698 (N_1698,In_2601,N_1305);
or U1699 (N_1699,N_740,In_522);
and U1700 (N_1700,In_2105,N_1365);
nor U1701 (N_1701,N_1247,In_1771);
and U1702 (N_1702,N_602,In_565);
xor U1703 (N_1703,N_1223,N_1434);
xnor U1704 (N_1704,In_332,In_700);
nor U1705 (N_1705,In_628,N_1109);
xnor U1706 (N_1706,N_1399,N_683);
nor U1707 (N_1707,N_1217,N_1314);
nand U1708 (N_1708,In_2981,N_1421);
nand U1709 (N_1709,In_3,N_1007);
nand U1710 (N_1710,In_123,In_1379);
nor U1711 (N_1711,In_314,N_596);
and U1712 (N_1712,N_1261,N_309);
nand U1713 (N_1713,N_1255,In_1115);
and U1714 (N_1714,In_774,N_1458);
nand U1715 (N_1715,N_1311,N_574);
or U1716 (N_1716,N_924,In_1507);
nor U1717 (N_1717,In_2553,N_70);
or U1718 (N_1718,N_1167,In_1369);
xor U1719 (N_1719,N_1287,In_812);
xnor U1720 (N_1720,In_1575,In_242);
nor U1721 (N_1721,In_410,N_1354);
xor U1722 (N_1722,In_626,In_818);
or U1723 (N_1723,N_1293,N_1483);
nor U1724 (N_1724,N_541,N_413);
and U1725 (N_1725,N_1427,N_835);
or U1726 (N_1726,N_253,N_1424);
or U1727 (N_1727,N_1215,In_19);
xnor U1728 (N_1728,N_158,In_364);
or U1729 (N_1729,In_1413,In_2935);
or U1730 (N_1730,N_543,In_2965);
and U1731 (N_1731,N_1414,N_1466);
xnor U1732 (N_1732,N_1253,N_1032);
and U1733 (N_1733,N_1485,In_2338);
xnor U1734 (N_1734,N_897,N_1256);
nor U1735 (N_1735,In_1229,N_1393);
nand U1736 (N_1736,In_1618,N_989);
or U1737 (N_1737,N_313,In_707);
xor U1738 (N_1738,In_2751,N_564);
and U1739 (N_1739,N_659,N_907);
xor U1740 (N_1740,N_346,In_850);
and U1741 (N_1741,In_2062,N_1482);
and U1742 (N_1742,N_1202,In_2856);
and U1743 (N_1743,N_1019,N_1428);
nor U1744 (N_1744,In_357,N_734);
and U1745 (N_1745,In_2130,N_489);
or U1746 (N_1746,N_0,In_1508);
and U1747 (N_1747,N_1447,N_487);
and U1748 (N_1748,N_1316,N_233);
or U1749 (N_1749,In_381,N_125);
and U1750 (N_1750,N_1103,In_1725);
or U1751 (N_1751,In_530,N_1081);
or U1752 (N_1752,N_550,N_1117);
and U1753 (N_1753,N_631,N_1395);
and U1754 (N_1754,In_2679,In_2434);
nor U1755 (N_1755,N_933,In_443);
nor U1756 (N_1756,In_860,In_1150);
and U1757 (N_1757,In_1021,N_1410);
xnor U1758 (N_1758,In_2317,N_1394);
and U1759 (N_1759,In_2826,In_892);
nand U1760 (N_1760,In_785,In_1719);
and U1761 (N_1761,In_240,In_2701);
nand U1762 (N_1762,N_275,In_2014);
and U1763 (N_1763,N_778,N_1358);
and U1764 (N_1764,N_748,N_1462);
nor U1765 (N_1765,N_925,In_1872);
or U1766 (N_1766,N_1222,N_1201);
or U1767 (N_1767,In_1016,In_806);
nand U1768 (N_1768,N_1161,N_1355);
xor U1769 (N_1769,In_955,N_964);
nor U1770 (N_1770,N_1240,In_309);
or U1771 (N_1771,In_971,In_1045);
nand U1772 (N_1772,N_958,In_300);
nor U1773 (N_1773,N_192,In_1748);
xor U1774 (N_1774,In_340,In_2142);
xor U1775 (N_1775,In_454,N_848);
and U1776 (N_1776,N_1118,N_679);
xor U1777 (N_1777,N_1306,In_654);
nand U1778 (N_1778,N_968,N_1236);
or U1779 (N_1779,N_719,In_1602);
nor U1780 (N_1780,N_1207,In_365);
xnor U1781 (N_1781,N_647,In_75);
nor U1782 (N_1782,In_1921,N_715);
or U1783 (N_1783,N_453,N_1491);
xor U1784 (N_1784,N_1338,In_810);
nor U1785 (N_1785,In_1106,In_2535);
xnor U1786 (N_1786,In_2623,N_1435);
and U1787 (N_1787,N_722,In_191);
and U1788 (N_1788,N_1264,In_2389);
xnor U1789 (N_1789,N_1409,N_1465);
and U1790 (N_1790,N_1271,N_1116);
xor U1791 (N_1791,N_741,N_1270);
or U1792 (N_1792,In_2119,In_679);
nor U1793 (N_1793,N_1363,N_1342);
and U1794 (N_1794,N_1163,In_2438);
xor U1795 (N_1795,N_1246,N_673);
nand U1796 (N_1796,N_621,N_983);
nor U1797 (N_1797,N_586,In_2135);
nand U1798 (N_1798,In_2755,N_615);
nor U1799 (N_1799,N_1214,In_457);
nor U1800 (N_1800,In_170,In_2952);
nor U1801 (N_1801,N_1325,N_517);
or U1802 (N_1802,In_2402,N_1494);
xor U1803 (N_1803,N_397,N_1144);
and U1804 (N_1804,In_2060,N_859);
or U1805 (N_1805,N_1412,N_651);
nor U1806 (N_1806,N_653,N_546);
xor U1807 (N_1807,In_1610,N_562);
and U1808 (N_1808,In_1148,N_1080);
nor U1809 (N_1809,N_1367,In_1865);
xor U1810 (N_1810,N_224,N_649);
or U1811 (N_1811,N_1064,N_1160);
or U1812 (N_1812,In_2841,In_2472);
and U1813 (N_1813,In_581,N_921);
nor U1814 (N_1814,N_1476,In_2703);
nor U1815 (N_1815,In_2824,N_1005);
or U1816 (N_1816,In_2316,N_720);
or U1817 (N_1817,N_739,N_1066);
xor U1818 (N_1818,N_693,N_1289);
nor U1819 (N_1819,In_731,In_1162);
xnor U1820 (N_1820,In_2051,N_978);
xnor U1821 (N_1821,N_1353,In_1011);
and U1822 (N_1822,N_1099,N_1093);
and U1823 (N_1823,N_291,In_808);
nand U1824 (N_1824,In_905,N_363);
and U1825 (N_1825,N_362,In_9);
and U1826 (N_1826,N_259,In_799);
or U1827 (N_1827,N_399,In_1627);
and U1828 (N_1828,N_1068,In_2543);
nand U1829 (N_1829,N_1176,N_1296);
and U1830 (N_1830,N_372,N_1);
nand U1831 (N_1831,N_986,In_1779);
xor U1832 (N_1832,N_998,N_823);
or U1833 (N_1833,In_2579,N_1308);
nor U1834 (N_1834,In_2694,N_1169);
xnor U1835 (N_1835,N_1397,In_1412);
or U1836 (N_1836,N_610,N_713);
nand U1837 (N_1837,In_715,N_927);
and U1838 (N_1838,N_717,N_822);
and U1839 (N_1839,In_1343,N_1031);
nor U1840 (N_1840,In_2554,N_1443);
nor U1841 (N_1841,In_2227,In_2990);
xnor U1842 (N_1842,N_1281,N_1446);
nand U1843 (N_1843,In_124,In_1542);
and U1844 (N_1844,N_135,In_389);
or U1845 (N_1845,In_2451,N_1243);
nor U1846 (N_1846,In_1102,N_1209);
nor U1847 (N_1847,N_389,N_1002);
or U1848 (N_1848,N_1004,N_1360);
or U1849 (N_1849,N_689,In_2676);
and U1850 (N_1850,N_136,In_1479);
xor U1851 (N_1851,In_1390,In_2148);
or U1852 (N_1852,In_1573,In_281);
or U1853 (N_1853,In_2312,In_1903);
or U1854 (N_1854,N_238,In_554);
and U1855 (N_1855,In_815,N_436);
and U1856 (N_1856,N_1055,In_2672);
nor U1857 (N_1857,N_1218,In_2230);
nor U1858 (N_1858,In_1658,In_2626);
and U1859 (N_1859,In_417,N_1063);
nand U1860 (N_1860,N_45,In_2784);
nor U1861 (N_1861,In_2255,In_1414);
xnor U1862 (N_1862,N_443,In_930);
and U1863 (N_1863,In_433,In_757);
and U1864 (N_1864,In_1950,N_954);
nor U1865 (N_1865,In_95,In_2080);
xor U1866 (N_1866,N_169,N_1431);
and U1867 (N_1867,In_590,N_320);
xor U1868 (N_1868,N_1230,N_1175);
nor U1869 (N_1869,N_592,In_1335);
and U1870 (N_1870,N_1432,N_1285);
or U1871 (N_1871,N_752,N_1423);
xnor U1872 (N_1872,N_1339,N_1457);
nor U1873 (N_1873,N_1232,In_2548);
nand U1874 (N_1874,N_829,N_1128);
and U1875 (N_1875,In_2379,N_1054);
or U1876 (N_1876,In_1652,N_1282);
and U1877 (N_1877,N_817,In_2386);
nor U1878 (N_1878,N_1131,N_1468);
nor U1879 (N_1879,In_352,In_2084);
nor U1880 (N_1880,In_2575,N_47);
xor U1881 (N_1881,In_303,N_1021);
nand U1882 (N_1882,In_222,N_1336);
and U1883 (N_1883,N_1408,N_1418);
nor U1884 (N_1884,N_768,N_1108);
or U1885 (N_1885,In_2592,N_1090);
xor U1886 (N_1886,In_2329,N_1020);
xor U1887 (N_1887,In_238,In_2132);
xor U1888 (N_1888,N_1172,N_1369);
or U1889 (N_1889,N_1291,N_1182);
xor U1890 (N_1890,N_1376,In_1523);
and U1891 (N_1891,N_1030,N_1228);
or U1892 (N_1892,N_1123,In_1778);
or U1893 (N_1893,N_815,N_723);
and U1894 (N_1894,N_1370,In_394);
xor U1895 (N_1895,In_1830,N_1371);
xor U1896 (N_1896,N_1173,N_1204);
xnor U1897 (N_1897,In_1600,N_1301);
xor U1898 (N_1898,N_470,N_1075);
and U1899 (N_1899,In_2342,N_1047);
nor U1900 (N_1900,In_1965,In_655);
nor U1901 (N_1901,N_929,N_557);
or U1902 (N_1902,N_837,N_1456);
or U1903 (N_1903,N_900,In_1464);
nor U1904 (N_1904,N_1356,N_1251);
nor U1905 (N_1905,N_975,In_291);
nor U1906 (N_1906,N_1061,In_2650);
and U1907 (N_1907,N_1138,In_2287);
or U1908 (N_1908,In_2648,N_1125);
or U1909 (N_1909,In_2504,N_1141);
or U1910 (N_1910,N_1089,N_873);
and U1911 (N_1911,N_273,N_906);
or U1912 (N_1912,In_65,In_25);
or U1913 (N_1913,N_1091,In_400);
nor U1914 (N_1914,N_1110,N_801);
nor U1915 (N_1915,N_1014,In_972);
nor U1916 (N_1916,In_354,N_1276);
nor U1917 (N_1917,N_1179,N_90);
or U1918 (N_1918,In_653,In_855);
and U1919 (N_1919,N_730,N_639);
nor U1920 (N_1920,In_1889,N_1135);
and U1921 (N_1921,N_1479,N_1362);
and U1922 (N_1922,N_555,N_1073);
and U1923 (N_1923,In_1361,In_1221);
nand U1924 (N_1924,In_1533,N_1489);
and U1925 (N_1925,In_614,N_1051);
nor U1926 (N_1926,In_591,N_1357);
or U1927 (N_1927,N_1187,N_1330);
nor U1928 (N_1928,N_844,N_1227);
or U1929 (N_1929,N_1473,In_2431);
xnor U1930 (N_1930,In_2116,N_898);
and U1931 (N_1931,In_1852,N_1477);
nor U1932 (N_1932,In_712,N_1211);
and U1933 (N_1933,N_558,In_741);
and U1934 (N_1934,N_20,In_938);
xor U1935 (N_1935,In_1807,N_485);
xor U1936 (N_1936,N_39,N_1252);
or U1937 (N_1937,N_981,N_626);
xnor U1938 (N_1938,N_687,In_1052);
nand U1939 (N_1939,In_1060,In_595);
nor U1940 (N_1940,N_1368,N_545);
or U1941 (N_1941,N_538,N_1084);
xor U1942 (N_1942,N_465,In_2853);
xor U1943 (N_1943,In_113,In_1359);
and U1944 (N_1944,In_1934,N_991);
or U1945 (N_1945,In_1215,N_819);
or U1946 (N_1946,In_504,In_771);
or U1947 (N_1947,In_564,N_824);
xnor U1948 (N_1948,N_1150,In_1983);
and U1949 (N_1949,N_155,N_1274);
and U1950 (N_1950,In_809,N_984);
or U1951 (N_1951,In_980,N_1340);
or U1952 (N_1952,N_1151,N_53);
nor U1953 (N_1953,In_116,N_1241);
or U1954 (N_1954,In_970,In_1625);
xor U1955 (N_1955,N_1411,N_1198);
nor U1956 (N_1956,N_1085,In_149);
nor U1957 (N_1957,In_492,In_1672);
nor U1958 (N_1958,N_1433,In_42);
or U1959 (N_1959,In_2294,N_1041);
nand U1960 (N_1960,N_773,In_1086);
or U1961 (N_1961,N_261,N_527);
xor U1962 (N_1962,N_1361,In_91);
nor U1963 (N_1963,N_1137,In_634);
nand U1964 (N_1964,In_1293,In_1256);
nor U1965 (N_1965,N_1320,In_2424);
nor U1966 (N_1966,N_1352,N_1044);
and U1967 (N_1967,In_1534,N_589);
xor U1968 (N_1968,In_344,N_245);
or U1969 (N_1969,In_2900,In_2170);
and U1970 (N_1970,In_2917,In_1225);
or U1971 (N_1971,N_167,N_226);
nor U1972 (N_1972,In_694,N_901);
or U1973 (N_1973,N_1046,In_1353);
nand U1974 (N_1974,N_1105,N_115);
and U1975 (N_1975,In_1704,N_1498);
xor U1976 (N_1976,In_1732,N_378);
and U1977 (N_1977,In_713,N_1486);
nand U1978 (N_1978,In_1230,In_482);
or U1979 (N_1979,N_1249,In_602);
nand U1980 (N_1980,N_514,N_67);
nand U1981 (N_1981,In_803,N_345);
nand U1982 (N_1982,In_2738,In_173);
nand U1983 (N_1983,In_2581,In_2254);
and U1984 (N_1984,N_431,In_2823);
and U1985 (N_1985,In_2875,N_422);
xor U1986 (N_1986,N_113,N_380);
nor U1987 (N_1987,In_250,N_860);
or U1988 (N_1988,In_2880,N_1497);
xnor U1989 (N_1989,In_610,In_2489);
and U1990 (N_1990,In_2159,N_518);
xor U1991 (N_1991,In_698,In_2206);
nand U1992 (N_1992,In_2372,In_927);
nand U1993 (N_1993,N_1350,In_263);
nor U1994 (N_1994,In_841,N_1042);
and U1995 (N_1995,In_1307,N_613);
or U1996 (N_1996,N_206,N_1100);
nor U1997 (N_1997,N_369,N_1043);
nor U1998 (N_1998,N_902,N_127);
or U1999 (N_1999,N_1012,In_1537);
nand U2000 (N_2000,N_1561,N_1351);
or U2001 (N_2001,N_1231,N_1901);
and U2002 (N_2002,In_274,N_1753);
xnor U2003 (N_2003,N_1592,N_1849);
nand U2004 (N_2004,N_1326,N_751);
or U2005 (N_2005,In_1300,N_1982);
or U2006 (N_2006,In_2221,N_1991);
or U2007 (N_2007,N_1048,N_1717);
nor U2008 (N_2008,In_2836,N_1999);
and U2009 (N_2009,In_1857,In_366);
or U2010 (N_2010,N_1205,N_1283);
nor U2011 (N_2011,In_1840,N_691);
nor U2012 (N_2012,N_1521,N_1907);
nand U2013 (N_2013,N_98,In_596);
nor U2014 (N_2014,N_1795,N_1671);
and U2015 (N_2015,In_918,N_1798);
and U2016 (N_2016,N_1761,N_1310);
or U2017 (N_2017,N_1953,In_2187);
or U2018 (N_2018,N_1933,N_1923);
nand U2019 (N_2019,N_682,N_1049);
and U2020 (N_2020,N_1559,N_1634);
xnor U2021 (N_2021,N_1941,N_1037);
nand U2022 (N_2022,N_1852,In_1913);
and U2023 (N_2023,N_1869,N_1934);
or U2024 (N_2024,N_1194,N_1695);
nand U2025 (N_2025,N_1006,N_1572);
xnor U2026 (N_2026,N_1730,N_1896);
xnor U2027 (N_2027,N_856,N_607);
nor U2028 (N_2028,N_1723,N_1897);
xnor U2029 (N_2029,N_828,In_500);
or U2030 (N_2030,N_1612,In_2169);
or U2031 (N_2031,N_1513,N_1807);
and U2032 (N_2032,In_1883,N_1725);
nand U2033 (N_2033,N_1467,In_1886);
and U2034 (N_2034,N_1908,N_1503);
nor U2035 (N_2035,In_2079,N_1579);
and U2036 (N_2036,N_1653,N_1894);
or U2037 (N_2037,N_1752,N_1805);
nor U2038 (N_2038,In_1171,N_1599);
or U2039 (N_2039,N_1670,N_1578);
nand U2040 (N_2040,N_911,N_1587);
nor U2041 (N_2041,N_1804,N_1487);
xor U2042 (N_2042,N_1567,N_1566);
or U2043 (N_2043,N_1917,N_1874);
nor U2044 (N_2044,N_1573,N_1687);
xnor U2045 (N_2045,In_2647,In_1350);
and U2046 (N_2046,In_1689,N_1644);
and U2047 (N_2047,N_1856,In_1853);
and U2048 (N_2048,N_1978,N_1906);
nand U2049 (N_2049,N_1146,N_503);
or U2050 (N_2050,N_1833,N_511);
nor U2051 (N_2051,In_1551,N_1819);
and U2052 (N_2052,N_1732,N_1976);
or U2053 (N_2053,N_1782,In_2813);
xnor U2054 (N_2054,In_1259,N_1386);
nand U2055 (N_2055,N_1657,N_1556);
and U2056 (N_2056,N_1268,In_2916);
and U2057 (N_2057,In_2729,N_1879);
nand U2058 (N_2058,N_1911,N_1775);
or U2059 (N_2059,N_945,In_560);
xnor U2060 (N_2060,In_1486,N_1977);
xor U2061 (N_2061,N_1574,N_1726);
or U2062 (N_2062,N_1951,N_771);
and U2063 (N_2063,N_1452,In_1522);
nor U2064 (N_2064,N_1083,N_1669);
nor U2065 (N_2065,N_581,In_2218);
nor U2066 (N_2066,In_1378,N_1506);
xnor U2067 (N_2067,N_1629,N_1382);
and U2068 (N_2068,In_85,N_1813);
and U2069 (N_2069,N_1778,N_1846);
nand U2070 (N_2070,N_1546,N_1347);
and U2071 (N_2071,In_1411,N_1745);
or U2072 (N_2072,In_1922,N_1710);
and U2073 (N_2073,N_1992,N_1810);
nor U2074 (N_2074,N_571,N_1668);
nor U2075 (N_2075,In_1126,N_1664);
and U2076 (N_2076,N_1372,N_1968);
and U2077 (N_2077,N_944,In_881);
and U2078 (N_2078,N_1680,N_1216);
xor U2079 (N_2079,N_1889,In_2177);
xnor U2080 (N_2080,In_412,N_1995);
xor U2081 (N_2081,N_1966,N_1171);
nor U2082 (N_2082,N_1300,N_1297);
nor U2083 (N_2083,N_1250,N_1294);
and U2084 (N_2084,In_1916,In_2732);
or U2085 (N_2085,N_1104,N_1742);
nor U2086 (N_2086,N_1863,In_1584);
xnor U2087 (N_2087,N_1769,N_1963);
or U2088 (N_2088,N_100,N_1983);
nand U2089 (N_2089,N_1490,N_1591);
xnor U2090 (N_2090,N_1760,In_1247);
and U2091 (N_2091,In_1193,N_1550);
and U2092 (N_2092,N_1520,N_1949);
nor U2093 (N_2093,N_1945,N_1984);
nor U2094 (N_2094,N_1830,N_1484);
nor U2095 (N_2095,N_1437,In_1911);
xor U2096 (N_2096,N_1082,N_1646);
xor U2097 (N_2097,N_1974,N_1877);
and U2098 (N_2098,N_1847,N_1796);
nand U2099 (N_2099,N_1586,N_1762);
nand U2100 (N_2100,N_1809,N_208);
nand U2101 (N_2101,N_1565,N_1815);
or U2102 (N_2102,N_1715,N_1783);
and U2103 (N_2103,N_1239,N_1617);
and U2104 (N_2104,N_1821,N_1625);
nand U2105 (N_2105,N_1806,N_1696);
and U2106 (N_2106,In_1755,N_1607);
and U2107 (N_2107,N_1737,N_387);
and U2108 (N_2108,N_1867,N_1870);
nor U2109 (N_2109,N_1195,N_1866);
xor U2110 (N_2110,N_855,In_471);
nand U2111 (N_2111,N_1773,In_2847);
xor U2112 (N_2112,N_540,N_1584);
xor U2113 (N_2113,N_1603,N_1900);
or U2114 (N_2114,N_1943,N_625);
and U2115 (N_2115,N_1802,N_1839);
xnor U2116 (N_2116,N_1551,N_334);
xnor U2117 (N_2117,In_1902,N_1748);
nand U2118 (N_2118,In_1243,N_1980);
and U2119 (N_2119,N_1528,In_1968);
nand U2120 (N_2120,N_710,N_716);
xnor U2121 (N_2121,N_1855,N_675);
or U2122 (N_2122,In_2854,N_1946);
nand U2123 (N_2123,N_84,N_1053);
and U2124 (N_2124,N_1534,N_1034);
and U2125 (N_2125,In_2404,In_1138);
nor U2126 (N_2126,N_34,In_2508);
nor U2127 (N_2127,N_1872,N_641);
or U2128 (N_2128,In_1478,N_1259);
and U2129 (N_2129,N_1101,N_1009);
and U2130 (N_2130,N_1700,In_754);
xnor U2131 (N_2131,N_400,N_1708);
or U2132 (N_2132,N_1691,N_893);
nor U2133 (N_2133,N_1588,N_838);
nand U2134 (N_2134,N_1970,N_953);
nand U2135 (N_2135,N_455,N_1153);
nor U2136 (N_2136,N_932,N_1292);
xor U2137 (N_2137,N_1596,N_1547);
or U2138 (N_2138,N_1419,In_1292);
nor U2139 (N_2139,N_1767,N_1562);
and U2140 (N_2140,N_1962,N_1450);
and U2141 (N_2141,N_58,In_569);
nand U2142 (N_2142,N_370,In_1696);
xnor U2143 (N_2143,N_50,N_1601);
or U2144 (N_2144,N_1474,N_1157);
and U2145 (N_2145,N_1107,N_1590);
nand U2146 (N_2146,N_1557,N_1640);
nand U2147 (N_2147,In_2083,N_1598);
nand U2148 (N_2148,N_1823,N_1000);
nor U2149 (N_2149,N_1790,In_467);
nand U2150 (N_2150,N_1985,N_1887);
and U2151 (N_2151,N_982,In_717);
or U2152 (N_2152,In_2373,N_1875);
or U2153 (N_2153,N_1641,N_1013);
nor U2154 (N_2154,N_1208,N_1820);
and U2155 (N_2155,N_1750,N_1618);
and U2156 (N_2156,N_1472,N_1927);
and U2157 (N_2157,N_1189,N_1543);
nor U2158 (N_2158,N_1121,In_758);
nand U2159 (N_2159,N_630,In_2191);
or U2160 (N_2160,N_211,N_890);
nand U2161 (N_2161,N_1238,N_1878);
nand U2162 (N_2162,N_1841,N_1880);
xor U2163 (N_2163,In_1320,N_310);
or U2164 (N_2164,N_1619,N_7);
and U2165 (N_2165,N_1589,N_1794);
or U2166 (N_2166,N_570,N_1130);
or U2167 (N_2167,N_1254,N_1940);
and U2168 (N_2168,N_1862,N_1803);
nor U2169 (N_2169,N_1666,N_568);
nor U2170 (N_2170,N_1743,In_1873);
or U2171 (N_2171,In_1282,In_2564);
nor U2172 (N_2172,N_1060,N_1515);
nand U2173 (N_2173,N_1720,N_173);
or U2174 (N_2174,N_1577,N_1098);
and U2175 (N_2175,N_19,N_1533);
nand U2176 (N_2176,N_1937,N_1865);
nand U2177 (N_2177,N_849,N_1831);
or U2178 (N_2178,N_1624,N_1413);
nand U2179 (N_2179,In_935,N_1164);
or U2180 (N_2180,N_1564,In_1733);
xnor U2181 (N_2181,N_509,N_1526);
and U2182 (N_2182,In_2502,In_2052);
xor U2183 (N_2183,N_1536,N_1333);
xor U2184 (N_2184,N_1848,In_2542);
nand U2185 (N_2185,N_1439,N_1738);
or U2186 (N_2186,N_1699,N_1784);
nand U2187 (N_2187,N_1295,In_54);
xnor U2188 (N_2188,N_711,N_1015);
xnor U2189 (N_2189,N_1686,In_2765);
nand U2190 (N_2190,N_1604,In_2394);
and U2191 (N_2191,N_1544,N_1665);
xnor U2192 (N_2192,N_1651,N_1147);
xor U2193 (N_2193,N_754,N_1132);
or U2194 (N_2194,N_1593,N_1994);
nand U2195 (N_2195,In_2997,N_1480);
xnor U2196 (N_2196,N_1729,N_1744);
xor U2197 (N_2197,N_1751,In_775);
nand U2198 (N_2198,In_1742,N_1772);
nor U2199 (N_2199,N_1514,In_89);
and U2200 (N_2200,N_1018,N_1344);
and U2201 (N_2201,N_1639,N_1517);
nand U2202 (N_2202,N_1661,N_1495);
xor U2203 (N_2203,N_1585,N_1518);
and U2204 (N_2204,N_1570,N_657);
nor U2205 (N_2205,N_1967,N_1902);
xor U2206 (N_2206,N_1861,N_1662);
xor U2207 (N_2207,In_4,N_762);
and U2208 (N_2208,N_133,N_1029);
or U2209 (N_2209,N_1859,N_1724);
nand U2210 (N_2210,N_330,In_2989);
nor U2211 (N_2211,In_1775,N_1505);
nor U2212 (N_2212,N_1426,N_1727);
and U2213 (N_2213,N_947,N_1212);
xor U2214 (N_2214,N_1986,N_1678);
nand U2215 (N_2215,In_1623,N_1965);
nand U2216 (N_2216,N_1582,N_1119);
xnor U2217 (N_2217,N_1913,N_572);
xnor U2218 (N_2218,N_1184,N_1840);
and U2219 (N_2219,N_1191,N_1697);
nand U2220 (N_2220,N_962,N_1667);
or U2221 (N_2221,N_1675,N_1154);
xnor U2222 (N_2222,In_948,N_1930);
nor U2223 (N_2223,N_1960,N_1660);
nor U2224 (N_2224,N_1455,N_1226);
or U2225 (N_2225,N_1793,N_1922);
and U2226 (N_2226,N_1685,N_1200);
xor U2227 (N_2227,N_1380,N_845);
nand U2228 (N_2228,N_1011,N_515);
and U2229 (N_2229,N_1449,N_1265);
and U2230 (N_2230,N_1735,N_1290);
nor U2231 (N_2231,N_1904,N_885);
nand U2232 (N_2232,N_1719,N_1749);
and U2233 (N_2233,N_1755,N_1873);
nand U2234 (N_2234,In_360,In_2406);
nor U2235 (N_2235,In_571,N_1885);
xnor U2236 (N_2236,N_1786,N_1523);
nand U2237 (N_2237,N_1890,N_1638);
nand U2238 (N_2238,N_1529,N_1502);
nor U2239 (N_2239,N_1812,In_1580);
xor U2240 (N_2240,N_1429,N_1508);
nor U2241 (N_2241,N_1219,N_1633);
and U2242 (N_2242,N_1971,N_1835);
xnor U2243 (N_2243,N_1555,N_1575);
xor U2244 (N_2244,N_1808,N_1628);
and U2245 (N_2245,N_1522,N_1711);
nand U2246 (N_2246,N_1964,N_1162);
or U2247 (N_2247,N_1510,N_1035);
xnor U2248 (N_2248,N_1854,In_2146);
xnor U2249 (N_2249,N_1001,N_1535);
xnor U2250 (N_2250,N_1791,In_82);
xor U2251 (N_2251,N_1597,N_145);
nor U2252 (N_2252,N_1771,In_769);
nor U2253 (N_2253,N_1989,In_224);
xnor U2254 (N_2254,N_1757,N_1939);
nor U2255 (N_2255,In_2239,N_1581);
or U2256 (N_2256,N_1088,In_293);
or U2257 (N_2257,N_1956,N_1549);
or U2258 (N_2258,N_1407,In_592);
xnor U2259 (N_2259,N_1348,N_755);
or U2260 (N_2260,N_1816,N_1284);
nor U2261 (N_2261,N_1756,N_1524);
and U2262 (N_2262,N_1655,N_1822);
xnor U2263 (N_2263,N_1837,In_2977);
nor U2264 (N_2264,N_1186,N_1857);
nand U2265 (N_2265,N_1876,N_867);
xor U2266 (N_2266,In_617,In_2734);
xnor U2267 (N_2267,In_2048,N_406);
nand U2268 (N_2268,N_1548,In_915);
and U2269 (N_2269,N_1152,In_2112);
nand U2270 (N_2270,In_2464,N_1036);
or U2271 (N_2271,N_1077,N_1690);
nand U2272 (N_2272,N_1914,N_1608);
nor U2273 (N_2273,N_1716,N_1683);
nor U2274 (N_2274,N_1610,N_1688);
and U2275 (N_2275,N_1383,N_1919);
nand U2276 (N_2276,N_1658,N_1684);
nor U2277 (N_2277,N_1682,In_2578);
and U2278 (N_2278,N_1309,N_1636);
or U2279 (N_2279,N_732,In_1510);
nand U2280 (N_2280,N_1979,N_491);
and U2281 (N_2281,N_1033,N_1627);
nor U2282 (N_2282,N_1705,N_1703);
nand U2283 (N_2283,N_1026,N_1817);
or U2284 (N_2284,N_1987,In_761);
xnor U2285 (N_2285,N_1728,In_1653);
and U2286 (N_2286,N_1958,In_1605);
nor U2287 (N_2287,In_2405,N_366);
nor U2288 (N_2288,N_1328,N_1650);
nor U2289 (N_2289,In_1759,N_909);
and U2290 (N_2290,N_753,N_1993);
or U2291 (N_2291,N_1560,N_1398);
xor U2292 (N_2292,N_1950,N_1779);
or U2293 (N_2293,In_2888,N_1663);
or U2294 (N_2294,N_1196,N_1527);
nand U2295 (N_2295,N_1788,In_756);
and U2296 (N_2296,N_1834,N_1681);
or U2297 (N_2297,N_1539,N_854);
or U2298 (N_2298,N_1948,N_1269);
nand U2299 (N_2299,N_1115,N_999);
xnor U2300 (N_2300,N_189,N_1471);
nor U2301 (N_2301,N_27,In_895);
xor U2302 (N_2302,N_1918,N_1286);
nand U2303 (N_2303,N_147,N_1166);
or U2304 (N_2304,In_1200,N_1928);
or U2305 (N_2305,N_1643,In_668);
and U2306 (N_2306,N_1500,N_1858);
or U2307 (N_2307,N_1747,N_1192);
and U2308 (N_2308,N_1884,N_1997);
or U2309 (N_2309,N_1954,N_85);
and U2310 (N_2310,In_2225,N_1540);
nand U2311 (N_2311,N_1079,N_1910);
or U2312 (N_2312,N_1893,In_480);
nor U2313 (N_2313,N_1512,N_1067);
nor U2314 (N_2314,N_1272,N_1768);
nor U2315 (N_2315,N_1996,N_1924);
nand U2316 (N_2316,N_1507,N_1076);
and U2317 (N_2317,N_1114,N_1647);
xor U2318 (N_2318,N_1595,N_1792);
xor U2319 (N_2319,N_1800,N_1766);
nor U2320 (N_2320,In_503,N_1955);
nand U2321 (N_2321,In_1947,N_1645);
or U2322 (N_2322,N_1611,N_919);
nor U2323 (N_2323,N_1741,N_1552);
nand U2324 (N_2324,N_1441,N_1197);
or U2325 (N_2325,N_1516,In_2395);
or U2326 (N_2326,N_1649,In_2087);
nor U2327 (N_2327,In_920,N_216);
and U2328 (N_2328,N_1142,N_1499);
xnor U2329 (N_2329,N_1780,In_822);
xor U2330 (N_2330,N_1542,In_557);
xor U2331 (N_2331,N_1713,N_479);
and U2332 (N_2332,N_1673,N_1621);
or U2333 (N_2333,N_1436,In_819);
nand U2334 (N_2334,N_1765,N_1942);
or U2335 (N_2335,N_1818,N_1733);
and U2336 (N_2336,N_1136,N_1039);
nor U2337 (N_2337,In_2309,N_1797);
xnor U2338 (N_2338,N_1938,N_770);
or U2339 (N_2339,N_1758,N_1538);
and U2340 (N_2340,N_1701,In_2667);
and U2341 (N_2341,N_1969,N_1981);
or U2342 (N_2342,N_1801,N_1040);
or U2343 (N_2343,In_163,N_322);
nor U2344 (N_2344,N_1836,In_661);
or U2345 (N_2345,N_1475,N_170);
nor U2346 (N_2346,In_2517,N_1777);
nand U2347 (N_2347,N_1926,N_1213);
xnor U2348 (N_2348,N_658,In_2005);
xnor U2349 (N_2349,N_1537,In_1952);
or U2350 (N_2350,N_1746,N_1576);
or U2351 (N_2351,In_404,In_887);
nor U2352 (N_2352,N_1895,N_677);
xnor U2353 (N_2353,N_1322,N_1092);
xnor U2354 (N_2354,N_1065,N_1883);
or U2355 (N_2355,N_577,N_1563);
xor U2356 (N_2356,N_1990,In_1273);
nand U2357 (N_2357,N_656,N_1864);
xor U2358 (N_2358,N_1459,N_1853);
xnor U2359 (N_2359,N_1102,In_2211);
nor U2360 (N_2360,N_1925,N_988);
xnor U2361 (N_2361,N_1959,N_605);
xnor U2362 (N_2362,N_1139,N_1706);
xor U2363 (N_2363,N_1722,N_11);
and U2364 (N_2364,N_1957,N_1909);
nand U2365 (N_2365,In_1304,N_1935);
or U2366 (N_2366,In_580,N_1530);
nor U2367 (N_2367,N_1961,In_2883);
xor U2368 (N_2368,N_1210,In_776);
nand U2369 (N_2369,N_1676,In_44);
nand U2370 (N_2370,N_1405,N_696);
xnor U2371 (N_2371,In_995,N_1860);
nand U2372 (N_2372,N_971,N_1143);
nand U2373 (N_2373,In_1591,N_306);
nor U2374 (N_2374,In_1499,In_1246);
xor U2375 (N_2375,N_1631,N_1659);
nand U2376 (N_2376,N_668,N_1406);
nor U2377 (N_2377,N_1799,In_219);
xor U2378 (N_2378,N_1126,N_1886);
or U2379 (N_2379,N_1672,N_1693);
nand U2380 (N_2380,N_1828,N_1609);
nand U2381 (N_2381,N_1714,N_1652);
or U2382 (N_2382,N_1656,In_231);
nor U2383 (N_2383,N_1844,N_1998);
nand U2384 (N_2384,In_405,In_1939);
xor U2385 (N_2385,N_1811,In_2337);
xor U2386 (N_2386,N_1605,N_1731);
nand U2387 (N_2387,N_1571,N_1898);
and U2388 (N_2388,N_1947,N_16);
and U2389 (N_2389,N_77,N_1882);
nand U2390 (N_2390,N_279,In_2741);
nand U2391 (N_2391,N_1613,In_833);
or U2392 (N_2392,N_1637,N_1975);
nor U2393 (N_2393,N_1622,N_1242);
nand U2394 (N_2394,N_714,N_1988);
nand U2395 (N_2395,N_1850,N_1888);
xnor U2396 (N_2396,In_199,N_1785);
xnor U2397 (N_2397,N_1600,N_618);
xnor U2398 (N_2398,N_1827,In_2940);
nor U2399 (N_2399,N_1824,In_2849);
nor U2400 (N_2400,N_177,In_2444);
or U2401 (N_2401,N_1632,In_2927);
and U2402 (N_2402,In_2714,N_1096);
nand U2403 (N_2403,N_1606,N_217);
nand U2404 (N_2404,N_1654,N_1718);
nand U2405 (N_2405,N_1826,N_1842);
xor U2406 (N_2406,In_1327,N_1694);
xor U2407 (N_2407,In_2141,N_1916);
and U2408 (N_2408,In_237,N_428);
or U2409 (N_2409,N_1871,N_976);
and U2410 (N_2410,N_1329,N_811);
nand U2411 (N_2411,N_1944,N_1263);
nand U2412 (N_2412,N_1554,N_1378);
xnor U2413 (N_2413,In_869,In_632);
xor U2414 (N_2414,N_1177,N_1478);
nand U2415 (N_2415,N_1829,In_2328);
or U2416 (N_2416,N_1912,N_1440);
and U2417 (N_2417,N_1759,In_1344);
or U2418 (N_2418,N_1375,N_1838);
or U2419 (N_2419,N_1148,N_1932);
nand U2420 (N_2420,N_1774,N_1648);
nor U2421 (N_2421,In_1219,N_1331);
nand U2422 (N_2422,In_2850,N_1734);
and U2423 (N_2423,In_2605,N_1062);
xor U2424 (N_2424,N_1509,N_1023);
xnor U2425 (N_2425,N_1525,N_1704);
nor U2426 (N_2426,N_1677,N_1374);
and U2427 (N_2427,N_1532,N_1531);
nand U2428 (N_2428,N_1787,In_1894);
or U2429 (N_2429,N_1776,N_1891);
xor U2430 (N_2430,N_1168,N_1074);
nand U2431 (N_2431,In_1332,N_421);
nor U2432 (N_2432,N_1332,N_966);
nand U2433 (N_2433,N_1199,N_1568);
nor U2434 (N_2434,N_1045,N_585);
nand U2435 (N_2435,N_1615,N_1936);
or U2436 (N_2436,N_1920,N_1511);
nor U2437 (N_2437,In_2624,In_2110);
and U2438 (N_2438,N_1345,N_970);
xnor U2439 (N_2439,N_1501,N_1594);
xor U2440 (N_2440,N_1868,N_26);
xnor U2441 (N_2441,In_177,N_1635);
and U2442 (N_2442,N_994,N_1277);
nand U2443 (N_2443,N_1709,N_1721);
or U2444 (N_2444,N_1915,N_923);
nor U2445 (N_2445,N_1623,N_1832);
and U2446 (N_2446,N_1679,In_1318);
xnor U2447 (N_2447,N_1469,In_1592);
and U2448 (N_2448,N_1364,In_1315);
xnor U2449 (N_2449,N_1086,N_1973);
nor U2450 (N_2450,N_1614,N_861);
or U2451 (N_2451,N_1707,N_1257);
xnor U2452 (N_2452,N_1905,N_1764);
or U2453 (N_2453,N_894,N_1580);
or U2454 (N_2454,N_1304,N_1087);
and U2455 (N_2455,In_1180,N_1692);
or U2456 (N_2456,N_1602,In_1494);
and U2457 (N_2457,N_1892,N_1781);
nor U2458 (N_2458,In_1975,N_1770);
or U2459 (N_2459,N_1626,N_1620);
nor U2460 (N_2460,In_495,In_481);
nor U2461 (N_2461,N_1642,N_623);
nand U2462 (N_2462,N_1881,N_1931);
nand U2463 (N_2463,N_1583,N_1324);
nor U2464 (N_2464,In_1480,In_1757);
or U2465 (N_2465,N_624,In_751);
nand U2466 (N_2466,N_1299,N_1165);
nand U2467 (N_2467,N_1843,N_1921);
xor U2468 (N_2468,N_1972,N_1553);
and U2469 (N_2469,N_1952,N_1814);
or U2470 (N_2470,N_1689,N_1630);
nor U2471 (N_2471,In_233,In_2877);
nand U2472 (N_2472,N_1313,N_1569);
and U2473 (N_2473,N_1056,N_1851);
and U2474 (N_2474,N_1464,N_1050);
nor U2475 (N_2475,In_2665,N_1180);
nand U2476 (N_2476,N_1698,In_1905);
or U2477 (N_2477,N_1519,In_1007);
xor U2478 (N_2478,N_1203,N_688);
xor U2479 (N_2479,N_1754,N_1156);
or U2480 (N_2480,N_1541,N_112);
and U2481 (N_2481,N_1702,N_1845);
nand U2482 (N_2482,In_658,In_2482);
nor U2483 (N_2483,N_1545,In_1829);
nand U2484 (N_2484,N_1488,N_448);
and U2485 (N_2485,N_1763,N_1558);
nand U2486 (N_2486,N_903,In_2137);
nor U2487 (N_2487,In_2643,N_1739);
or U2488 (N_2488,N_31,N_1899);
nand U2489 (N_2489,In_1972,In_767);
nand U2490 (N_2490,N_1789,N_640);
nor U2491 (N_2491,N_843,N_1712);
and U2492 (N_2492,N_1903,N_1674);
or U2493 (N_2493,N_1149,N_1616);
nor U2494 (N_2494,N_1825,N_1736);
nand U2495 (N_2495,N_352,N_1445);
nor U2496 (N_2496,N_821,N_1740);
xnor U2497 (N_2497,In_135,In_1159);
nor U2498 (N_2498,N_1122,N_1929);
nand U2499 (N_2499,N_1504,In_2692);
or U2500 (N_2500,N_2410,N_2343);
xnor U2501 (N_2501,N_2001,N_2095);
nor U2502 (N_2502,N_2327,N_2121);
nor U2503 (N_2503,N_2429,N_2240);
and U2504 (N_2504,N_2292,N_2259);
xor U2505 (N_2505,N_2146,N_2243);
xor U2506 (N_2506,N_2149,N_2481);
nand U2507 (N_2507,N_2123,N_2318);
or U2508 (N_2508,N_2031,N_2023);
nor U2509 (N_2509,N_2353,N_2345);
and U2510 (N_2510,N_2004,N_2443);
and U2511 (N_2511,N_2043,N_2349);
nand U2512 (N_2512,N_2332,N_2080);
or U2513 (N_2513,N_2423,N_2256);
or U2514 (N_2514,N_2272,N_2113);
nand U2515 (N_2515,N_2270,N_2066);
or U2516 (N_2516,N_2276,N_2331);
xor U2517 (N_2517,N_2226,N_2457);
nand U2518 (N_2518,N_2394,N_2025);
and U2519 (N_2519,N_2225,N_2147);
xor U2520 (N_2520,N_2328,N_2300);
and U2521 (N_2521,N_2083,N_2290);
or U2522 (N_2522,N_2315,N_2101);
nor U2523 (N_2523,N_2164,N_2071);
nand U2524 (N_2524,N_2373,N_2430);
and U2525 (N_2525,N_2491,N_2335);
nor U2526 (N_2526,N_2236,N_2428);
nand U2527 (N_2527,N_2417,N_2143);
and U2528 (N_2528,N_2406,N_2026);
nor U2529 (N_2529,N_2037,N_2237);
or U2530 (N_2530,N_2049,N_2145);
or U2531 (N_2531,N_2057,N_2397);
xor U2532 (N_2532,N_2062,N_2171);
nand U2533 (N_2533,N_2364,N_2486);
and U2534 (N_2534,N_2210,N_2303);
nand U2535 (N_2535,N_2483,N_2393);
nand U2536 (N_2536,N_2021,N_2378);
nor U2537 (N_2537,N_2196,N_2116);
xnor U2538 (N_2538,N_2405,N_2374);
and U2539 (N_2539,N_2260,N_2007);
or U2540 (N_2540,N_2231,N_2494);
and U2541 (N_2541,N_2176,N_2006);
and U2542 (N_2542,N_2120,N_2469);
nand U2543 (N_2543,N_2161,N_2306);
and U2544 (N_2544,N_2202,N_2163);
and U2545 (N_2545,N_2440,N_2117);
or U2546 (N_2546,N_2126,N_2453);
or U2547 (N_2547,N_2365,N_2449);
nand U2548 (N_2548,N_2319,N_2036);
nand U2549 (N_2549,N_2358,N_2132);
nand U2550 (N_2550,N_2380,N_2056);
xnor U2551 (N_2551,N_2351,N_2361);
xnor U2552 (N_2552,N_2170,N_2400);
and U2553 (N_2553,N_2368,N_2076);
xnor U2554 (N_2554,N_2341,N_2371);
nor U2555 (N_2555,N_2392,N_2114);
nor U2556 (N_2556,N_2468,N_2325);
and U2557 (N_2557,N_2246,N_2254);
xnor U2558 (N_2558,N_2340,N_2388);
or U2559 (N_2559,N_2191,N_2017);
or U2560 (N_2560,N_2496,N_2234);
or U2561 (N_2561,N_2168,N_2263);
or U2562 (N_2562,N_2019,N_2297);
nand U2563 (N_2563,N_2250,N_2182);
or U2564 (N_2564,N_2252,N_2474);
nand U2565 (N_2565,N_2151,N_2442);
or U2566 (N_2566,N_2248,N_2134);
nor U2567 (N_2567,N_2310,N_2424);
nand U2568 (N_2568,N_2222,N_2142);
xor U2569 (N_2569,N_2369,N_2399);
nor U2570 (N_2570,N_2301,N_2154);
nor U2571 (N_2571,N_2375,N_2452);
nand U2572 (N_2572,N_2081,N_2199);
nor U2573 (N_2573,N_2412,N_2352);
xnor U2574 (N_2574,N_2213,N_2065);
nor U2575 (N_2575,N_2419,N_2032);
xnor U2576 (N_2576,N_2158,N_2459);
or U2577 (N_2577,N_2135,N_2063);
xnor U2578 (N_2578,N_2175,N_2466);
nor U2579 (N_2579,N_2401,N_2233);
and U2580 (N_2580,N_2268,N_2011);
or U2581 (N_2581,N_2067,N_2133);
nand U2582 (N_2582,N_2311,N_2125);
nand U2583 (N_2583,N_2185,N_2489);
and U2584 (N_2584,N_2344,N_2472);
and U2585 (N_2585,N_2389,N_2497);
or U2586 (N_2586,N_2055,N_2077);
or U2587 (N_2587,N_2153,N_2040);
xnor U2588 (N_2588,N_2109,N_2090);
nand U2589 (N_2589,N_2304,N_2041);
nor U2590 (N_2590,N_2159,N_2262);
xnor U2591 (N_2591,N_2299,N_2277);
xnor U2592 (N_2592,N_2008,N_2316);
nand U2593 (N_2593,N_2033,N_2293);
nand U2594 (N_2594,N_2314,N_2321);
or U2595 (N_2595,N_2356,N_2039);
nand U2596 (N_2596,N_2330,N_2470);
and U2597 (N_2597,N_2326,N_2172);
or U2598 (N_2598,N_2035,N_2278);
or U2599 (N_2599,N_2433,N_2279);
or U2600 (N_2600,N_2460,N_2238);
xor U2601 (N_2601,N_2432,N_2102);
nor U2602 (N_2602,N_2415,N_2169);
or U2603 (N_2603,N_2018,N_2088);
nand U2604 (N_2604,N_2408,N_2436);
or U2605 (N_2605,N_2187,N_2287);
and U2606 (N_2606,N_2334,N_2059);
and U2607 (N_2607,N_2028,N_2354);
xor U2608 (N_2608,N_2480,N_2091);
or U2609 (N_2609,N_2228,N_2178);
nor U2610 (N_2610,N_2136,N_2195);
and U2611 (N_2611,N_2112,N_2479);
and U2612 (N_2612,N_2414,N_2317);
nor U2613 (N_2613,N_2336,N_2087);
xor U2614 (N_2614,N_2488,N_2167);
nand U2615 (N_2615,N_2082,N_2044);
xor U2616 (N_2616,N_2291,N_2129);
and U2617 (N_2617,N_2014,N_2431);
or U2618 (N_2618,N_2402,N_2329);
or U2619 (N_2619,N_2435,N_2390);
xor U2620 (N_2620,N_2387,N_2070);
and U2621 (N_2621,N_2339,N_2338);
and U2622 (N_2622,N_2425,N_2286);
nand U2623 (N_2623,N_2212,N_2103);
nor U2624 (N_2624,N_2219,N_2235);
and U2625 (N_2625,N_2376,N_2485);
nor U2626 (N_2626,N_2060,N_2174);
or U2627 (N_2627,N_2477,N_2285);
or U2628 (N_2628,N_2024,N_2094);
nand U2629 (N_2629,N_2015,N_2463);
xor U2630 (N_2630,N_2258,N_2451);
and U2631 (N_2631,N_2438,N_2005);
nor U2632 (N_2632,N_2128,N_2002);
nand U2633 (N_2633,N_2323,N_2131);
xor U2634 (N_2634,N_2089,N_2478);
nand U2635 (N_2635,N_2458,N_2162);
or U2636 (N_2636,N_2052,N_2072);
or U2637 (N_2637,N_2189,N_2296);
nand U2638 (N_2638,N_2229,N_2421);
xor U2639 (N_2639,N_2152,N_2079);
nand U2640 (N_2640,N_2230,N_2075);
nor U2641 (N_2641,N_2267,N_2064);
or U2642 (N_2642,N_2156,N_2192);
and U2643 (N_2643,N_2115,N_2359);
or U2644 (N_2644,N_2122,N_2398);
and U2645 (N_2645,N_2096,N_2367);
nand U2646 (N_2646,N_2241,N_2097);
nand U2647 (N_2647,N_2216,N_2180);
and U2648 (N_2648,N_2073,N_2404);
or U2649 (N_2649,N_2000,N_2181);
or U2650 (N_2650,N_2355,N_2061);
xnor U2651 (N_2651,N_2038,N_2141);
xor U2652 (N_2652,N_2224,N_2119);
nand U2653 (N_2653,N_2194,N_2160);
or U2654 (N_2654,N_2068,N_2223);
or U2655 (N_2655,N_2207,N_2475);
nor U2656 (N_2656,N_2030,N_2016);
and U2657 (N_2657,N_2420,N_2211);
nand U2658 (N_2658,N_2370,N_2499);
and U2659 (N_2659,N_2034,N_2385);
and U2660 (N_2660,N_2053,N_2454);
nand U2661 (N_2661,N_2245,N_2188);
or U2662 (N_2662,N_2092,N_2084);
nand U2663 (N_2663,N_2003,N_2273);
nand U2664 (N_2664,N_2281,N_2221);
nand U2665 (N_2665,N_2027,N_2382);
or U2666 (N_2666,N_2009,N_2283);
xor U2667 (N_2667,N_2029,N_2298);
nand U2668 (N_2668,N_2455,N_2322);
nand U2669 (N_2669,N_2437,N_2342);
and U2670 (N_2670,N_2434,N_2013);
xnor U2671 (N_2671,N_2379,N_2179);
and U2672 (N_2672,N_2461,N_2183);
nand U2673 (N_2673,N_2372,N_2232);
nand U2674 (N_2674,N_2208,N_2280);
nand U2675 (N_2675,N_2193,N_2465);
and U2676 (N_2676,N_2289,N_2138);
and U2677 (N_2677,N_2209,N_2155);
nand U2678 (N_2678,N_2139,N_2493);
xnor U2679 (N_2679,N_2418,N_2020);
nor U2680 (N_2680,N_2074,N_2242);
and U2681 (N_2681,N_2140,N_2487);
xor U2682 (N_2682,N_2190,N_2107);
nand U2683 (N_2683,N_2058,N_2106);
nor U2684 (N_2684,N_2462,N_2274);
and U2685 (N_2685,N_2492,N_2100);
nand U2686 (N_2686,N_2022,N_2383);
and U2687 (N_2687,N_2409,N_2490);
and U2688 (N_2688,N_2403,N_2085);
nor U2689 (N_2689,N_2220,N_2456);
nor U2690 (N_2690,N_2484,N_2377);
nor U2691 (N_2691,N_2148,N_2214);
xnor U2692 (N_2692,N_2395,N_2294);
nor U2693 (N_2693,N_2047,N_2086);
or U2694 (N_2694,N_2426,N_2203);
and U2695 (N_2695,N_2166,N_2108);
nand U2696 (N_2696,N_2444,N_2307);
and U2697 (N_2697,N_2205,N_2105);
or U2698 (N_2698,N_2467,N_2337);
or U2699 (N_2699,N_2320,N_2157);
and U2700 (N_2700,N_2045,N_2261);
nand U2701 (N_2701,N_2251,N_2144);
xor U2702 (N_2702,N_2305,N_2098);
or U2703 (N_2703,N_2165,N_2284);
xnor U2704 (N_2704,N_2275,N_2093);
or U2705 (N_2705,N_2295,N_2054);
nor U2706 (N_2706,N_2288,N_2150);
xnor U2707 (N_2707,N_2333,N_2416);
and U2708 (N_2708,N_2204,N_2244);
and U2709 (N_2709,N_2111,N_2201);
nand U2710 (N_2710,N_2069,N_2313);
and U2711 (N_2711,N_2264,N_2445);
xor U2712 (N_2712,N_2366,N_2448);
nand U2713 (N_2713,N_2206,N_2441);
nand U2714 (N_2714,N_2363,N_2124);
and U2715 (N_2715,N_2396,N_2422);
nand U2716 (N_2716,N_2099,N_2253);
nand U2717 (N_2717,N_2266,N_2347);
or U2718 (N_2718,N_2200,N_2217);
or U2719 (N_2719,N_2498,N_2257);
or U2720 (N_2720,N_2476,N_2177);
nand U2721 (N_2721,N_2350,N_2186);
nor U2722 (N_2722,N_2473,N_2249);
nand U2723 (N_2723,N_2197,N_2184);
nor U2724 (N_2724,N_2471,N_2269);
or U2725 (N_2725,N_2384,N_2427);
xor U2726 (N_2726,N_2271,N_2042);
and U2727 (N_2727,N_2446,N_2309);
nand U2728 (N_2728,N_2215,N_2198);
nor U2729 (N_2729,N_2447,N_2247);
and U2730 (N_2730,N_2130,N_2104);
nor U2731 (N_2731,N_2407,N_2348);
nand U2732 (N_2732,N_2239,N_2110);
or U2733 (N_2733,N_2346,N_2360);
xor U2734 (N_2734,N_2439,N_2413);
xor U2735 (N_2735,N_2312,N_2218);
nor U2736 (N_2736,N_2051,N_2450);
or U2737 (N_2737,N_2464,N_2381);
nand U2738 (N_2738,N_2127,N_2227);
or U2739 (N_2739,N_2173,N_2050);
xnor U2740 (N_2740,N_2411,N_2482);
xor U2741 (N_2741,N_2137,N_2048);
nand U2742 (N_2742,N_2495,N_2357);
or U2743 (N_2743,N_2391,N_2118);
nor U2744 (N_2744,N_2386,N_2046);
nor U2745 (N_2745,N_2324,N_2078);
nand U2746 (N_2746,N_2308,N_2362);
xnor U2747 (N_2747,N_2282,N_2302);
xnor U2748 (N_2748,N_2012,N_2265);
nand U2749 (N_2749,N_2255,N_2010);
and U2750 (N_2750,N_2084,N_2362);
and U2751 (N_2751,N_2390,N_2044);
xor U2752 (N_2752,N_2237,N_2248);
nand U2753 (N_2753,N_2400,N_2135);
or U2754 (N_2754,N_2045,N_2429);
and U2755 (N_2755,N_2300,N_2354);
xor U2756 (N_2756,N_2239,N_2259);
or U2757 (N_2757,N_2056,N_2333);
and U2758 (N_2758,N_2297,N_2396);
and U2759 (N_2759,N_2091,N_2326);
nand U2760 (N_2760,N_2027,N_2214);
nor U2761 (N_2761,N_2235,N_2091);
xor U2762 (N_2762,N_2015,N_2323);
xor U2763 (N_2763,N_2448,N_2153);
nor U2764 (N_2764,N_2326,N_2103);
nand U2765 (N_2765,N_2426,N_2278);
xnor U2766 (N_2766,N_2301,N_2027);
nor U2767 (N_2767,N_2432,N_2064);
nand U2768 (N_2768,N_2281,N_2026);
xnor U2769 (N_2769,N_2275,N_2261);
and U2770 (N_2770,N_2104,N_2276);
nand U2771 (N_2771,N_2143,N_2079);
nor U2772 (N_2772,N_2153,N_2401);
or U2773 (N_2773,N_2187,N_2141);
and U2774 (N_2774,N_2323,N_2218);
nor U2775 (N_2775,N_2318,N_2319);
nor U2776 (N_2776,N_2479,N_2178);
nor U2777 (N_2777,N_2345,N_2299);
nor U2778 (N_2778,N_2116,N_2232);
nor U2779 (N_2779,N_2230,N_2199);
or U2780 (N_2780,N_2091,N_2029);
and U2781 (N_2781,N_2129,N_2397);
and U2782 (N_2782,N_2317,N_2293);
xor U2783 (N_2783,N_2230,N_2071);
or U2784 (N_2784,N_2431,N_2386);
nor U2785 (N_2785,N_2292,N_2070);
and U2786 (N_2786,N_2470,N_2351);
and U2787 (N_2787,N_2366,N_2486);
nor U2788 (N_2788,N_2422,N_2420);
nand U2789 (N_2789,N_2334,N_2268);
or U2790 (N_2790,N_2061,N_2284);
and U2791 (N_2791,N_2100,N_2289);
nand U2792 (N_2792,N_2130,N_2242);
or U2793 (N_2793,N_2337,N_2330);
nor U2794 (N_2794,N_2070,N_2121);
or U2795 (N_2795,N_2028,N_2007);
and U2796 (N_2796,N_2305,N_2140);
or U2797 (N_2797,N_2304,N_2084);
or U2798 (N_2798,N_2050,N_2047);
and U2799 (N_2799,N_2132,N_2313);
nand U2800 (N_2800,N_2209,N_2437);
or U2801 (N_2801,N_2435,N_2279);
nand U2802 (N_2802,N_2349,N_2114);
xnor U2803 (N_2803,N_2366,N_2218);
nand U2804 (N_2804,N_2400,N_2257);
xor U2805 (N_2805,N_2118,N_2119);
or U2806 (N_2806,N_2259,N_2258);
or U2807 (N_2807,N_2156,N_2260);
nor U2808 (N_2808,N_2100,N_2183);
nand U2809 (N_2809,N_2003,N_2022);
and U2810 (N_2810,N_2082,N_2010);
xnor U2811 (N_2811,N_2264,N_2475);
xor U2812 (N_2812,N_2057,N_2322);
nor U2813 (N_2813,N_2322,N_2442);
nor U2814 (N_2814,N_2247,N_2227);
and U2815 (N_2815,N_2079,N_2442);
xnor U2816 (N_2816,N_2072,N_2431);
nor U2817 (N_2817,N_2488,N_2412);
xnor U2818 (N_2818,N_2147,N_2217);
xor U2819 (N_2819,N_2008,N_2423);
nand U2820 (N_2820,N_2228,N_2149);
and U2821 (N_2821,N_2480,N_2056);
and U2822 (N_2822,N_2481,N_2282);
nor U2823 (N_2823,N_2374,N_2093);
or U2824 (N_2824,N_2271,N_2173);
and U2825 (N_2825,N_2163,N_2295);
or U2826 (N_2826,N_2091,N_2110);
and U2827 (N_2827,N_2320,N_2041);
nand U2828 (N_2828,N_2234,N_2095);
and U2829 (N_2829,N_2261,N_2271);
xnor U2830 (N_2830,N_2471,N_2294);
or U2831 (N_2831,N_2380,N_2412);
nor U2832 (N_2832,N_2480,N_2403);
or U2833 (N_2833,N_2399,N_2323);
nand U2834 (N_2834,N_2384,N_2198);
xnor U2835 (N_2835,N_2032,N_2340);
nand U2836 (N_2836,N_2098,N_2378);
or U2837 (N_2837,N_2393,N_2353);
and U2838 (N_2838,N_2295,N_2097);
nor U2839 (N_2839,N_2162,N_2405);
and U2840 (N_2840,N_2425,N_2071);
and U2841 (N_2841,N_2317,N_2320);
nor U2842 (N_2842,N_2320,N_2295);
nor U2843 (N_2843,N_2245,N_2033);
nand U2844 (N_2844,N_2024,N_2406);
nand U2845 (N_2845,N_2047,N_2436);
and U2846 (N_2846,N_2379,N_2284);
nand U2847 (N_2847,N_2474,N_2065);
and U2848 (N_2848,N_2409,N_2069);
and U2849 (N_2849,N_2243,N_2296);
and U2850 (N_2850,N_2231,N_2480);
and U2851 (N_2851,N_2230,N_2233);
or U2852 (N_2852,N_2181,N_2450);
or U2853 (N_2853,N_2010,N_2042);
xnor U2854 (N_2854,N_2105,N_2132);
nor U2855 (N_2855,N_2386,N_2250);
and U2856 (N_2856,N_2090,N_2348);
nand U2857 (N_2857,N_2196,N_2050);
nor U2858 (N_2858,N_2118,N_2360);
nor U2859 (N_2859,N_2312,N_2253);
or U2860 (N_2860,N_2283,N_2394);
and U2861 (N_2861,N_2373,N_2066);
or U2862 (N_2862,N_2246,N_2043);
xnor U2863 (N_2863,N_2426,N_2464);
xnor U2864 (N_2864,N_2029,N_2219);
and U2865 (N_2865,N_2382,N_2085);
and U2866 (N_2866,N_2466,N_2396);
nand U2867 (N_2867,N_2032,N_2456);
xor U2868 (N_2868,N_2155,N_2140);
and U2869 (N_2869,N_2481,N_2463);
or U2870 (N_2870,N_2402,N_2068);
xnor U2871 (N_2871,N_2244,N_2274);
and U2872 (N_2872,N_2149,N_2169);
xnor U2873 (N_2873,N_2083,N_2306);
or U2874 (N_2874,N_2118,N_2043);
and U2875 (N_2875,N_2188,N_2337);
nand U2876 (N_2876,N_2125,N_2277);
or U2877 (N_2877,N_2493,N_2067);
xor U2878 (N_2878,N_2020,N_2361);
or U2879 (N_2879,N_2494,N_2411);
xor U2880 (N_2880,N_2305,N_2422);
xnor U2881 (N_2881,N_2179,N_2232);
xor U2882 (N_2882,N_2296,N_2410);
nor U2883 (N_2883,N_2284,N_2447);
nor U2884 (N_2884,N_2057,N_2078);
or U2885 (N_2885,N_2129,N_2446);
xor U2886 (N_2886,N_2367,N_2170);
nor U2887 (N_2887,N_2398,N_2428);
xor U2888 (N_2888,N_2472,N_2337);
nor U2889 (N_2889,N_2096,N_2083);
xnor U2890 (N_2890,N_2289,N_2066);
nand U2891 (N_2891,N_2362,N_2201);
xor U2892 (N_2892,N_2033,N_2333);
nor U2893 (N_2893,N_2381,N_2066);
xor U2894 (N_2894,N_2396,N_2314);
xnor U2895 (N_2895,N_2373,N_2268);
nand U2896 (N_2896,N_2280,N_2454);
nor U2897 (N_2897,N_2328,N_2255);
nand U2898 (N_2898,N_2275,N_2360);
or U2899 (N_2899,N_2333,N_2419);
nand U2900 (N_2900,N_2473,N_2170);
nor U2901 (N_2901,N_2244,N_2495);
nor U2902 (N_2902,N_2454,N_2078);
xnor U2903 (N_2903,N_2352,N_2357);
nand U2904 (N_2904,N_2249,N_2222);
nor U2905 (N_2905,N_2165,N_2464);
nor U2906 (N_2906,N_2265,N_2291);
and U2907 (N_2907,N_2475,N_2431);
xor U2908 (N_2908,N_2182,N_2197);
xor U2909 (N_2909,N_2358,N_2454);
nand U2910 (N_2910,N_2315,N_2221);
xor U2911 (N_2911,N_2144,N_2451);
nor U2912 (N_2912,N_2407,N_2310);
nor U2913 (N_2913,N_2020,N_2005);
xnor U2914 (N_2914,N_2120,N_2410);
or U2915 (N_2915,N_2141,N_2265);
nor U2916 (N_2916,N_2137,N_2196);
nand U2917 (N_2917,N_2399,N_2222);
nand U2918 (N_2918,N_2070,N_2490);
or U2919 (N_2919,N_2319,N_2487);
and U2920 (N_2920,N_2174,N_2048);
or U2921 (N_2921,N_2311,N_2455);
and U2922 (N_2922,N_2150,N_2181);
nor U2923 (N_2923,N_2205,N_2371);
nand U2924 (N_2924,N_2433,N_2072);
nand U2925 (N_2925,N_2287,N_2156);
nor U2926 (N_2926,N_2056,N_2120);
xor U2927 (N_2927,N_2279,N_2247);
nand U2928 (N_2928,N_2001,N_2100);
or U2929 (N_2929,N_2011,N_2280);
and U2930 (N_2930,N_2298,N_2038);
xnor U2931 (N_2931,N_2342,N_2419);
xnor U2932 (N_2932,N_2339,N_2180);
nor U2933 (N_2933,N_2145,N_2401);
xnor U2934 (N_2934,N_2091,N_2186);
xor U2935 (N_2935,N_2402,N_2303);
or U2936 (N_2936,N_2056,N_2409);
xnor U2937 (N_2937,N_2395,N_2108);
and U2938 (N_2938,N_2227,N_2238);
or U2939 (N_2939,N_2312,N_2411);
xor U2940 (N_2940,N_2200,N_2382);
xnor U2941 (N_2941,N_2468,N_2462);
and U2942 (N_2942,N_2420,N_2403);
or U2943 (N_2943,N_2269,N_2315);
nor U2944 (N_2944,N_2131,N_2000);
nor U2945 (N_2945,N_2004,N_2338);
and U2946 (N_2946,N_2238,N_2360);
nor U2947 (N_2947,N_2248,N_2238);
xnor U2948 (N_2948,N_2358,N_2260);
or U2949 (N_2949,N_2367,N_2198);
and U2950 (N_2950,N_2122,N_2366);
or U2951 (N_2951,N_2097,N_2322);
nand U2952 (N_2952,N_2380,N_2300);
nor U2953 (N_2953,N_2353,N_2492);
or U2954 (N_2954,N_2221,N_2179);
and U2955 (N_2955,N_2048,N_2464);
xor U2956 (N_2956,N_2224,N_2352);
or U2957 (N_2957,N_2106,N_2212);
nor U2958 (N_2958,N_2351,N_2112);
nor U2959 (N_2959,N_2422,N_2272);
nor U2960 (N_2960,N_2039,N_2226);
nor U2961 (N_2961,N_2184,N_2401);
or U2962 (N_2962,N_2064,N_2494);
xor U2963 (N_2963,N_2444,N_2151);
nand U2964 (N_2964,N_2114,N_2030);
and U2965 (N_2965,N_2421,N_2458);
and U2966 (N_2966,N_2383,N_2177);
xor U2967 (N_2967,N_2031,N_2140);
or U2968 (N_2968,N_2003,N_2101);
nor U2969 (N_2969,N_2240,N_2467);
xor U2970 (N_2970,N_2354,N_2454);
nor U2971 (N_2971,N_2268,N_2031);
nand U2972 (N_2972,N_2208,N_2414);
nor U2973 (N_2973,N_2454,N_2047);
and U2974 (N_2974,N_2391,N_2124);
xnor U2975 (N_2975,N_2254,N_2080);
nand U2976 (N_2976,N_2390,N_2170);
and U2977 (N_2977,N_2180,N_2014);
and U2978 (N_2978,N_2239,N_2490);
xor U2979 (N_2979,N_2371,N_2296);
nor U2980 (N_2980,N_2168,N_2320);
and U2981 (N_2981,N_2003,N_2270);
or U2982 (N_2982,N_2275,N_2084);
nand U2983 (N_2983,N_2201,N_2447);
xor U2984 (N_2984,N_2334,N_2208);
nand U2985 (N_2985,N_2180,N_2206);
and U2986 (N_2986,N_2341,N_2349);
nor U2987 (N_2987,N_2092,N_2160);
and U2988 (N_2988,N_2204,N_2340);
nand U2989 (N_2989,N_2434,N_2052);
nand U2990 (N_2990,N_2097,N_2173);
nand U2991 (N_2991,N_2075,N_2416);
nor U2992 (N_2992,N_2180,N_2119);
xor U2993 (N_2993,N_2411,N_2377);
or U2994 (N_2994,N_2323,N_2280);
nor U2995 (N_2995,N_2260,N_2235);
and U2996 (N_2996,N_2000,N_2388);
and U2997 (N_2997,N_2187,N_2258);
and U2998 (N_2998,N_2256,N_2284);
xor U2999 (N_2999,N_2277,N_2021);
nor U3000 (N_3000,N_2545,N_2890);
nand U3001 (N_3001,N_2956,N_2945);
and U3002 (N_3002,N_2584,N_2693);
xor U3003 (N_3003,N_2643,N_2874);
xnor U3004 (N_3004,N_2975,N_2656);
nor U3005 (N_3005,N_2638,N_2875);
nor U3006 (N_3006,N_2591,N_2520);
and U3007 (N_3007,N_2926,N_2561);
or U3008 (N_3008,N_2614,N_2585);
xor U3009 (N_3009,N_2665,N_2774);
xor U3010 (N_3010,N_2634,N_2647);
and U3011 (N_3011,N_2941,N_2501);
nor U3012 (N_3012,N_2703,N_2842);
nor U3013 (N_3013,N_2780,N_2531);
and U3014 (N_3014,N_2611,N_2723);
xor U3015 (N_3015,N_2893,N_2543);
or U3016 (N_3016,N_2789,N_2912);
nand U3017 (N_3017,N_2848,N_2982);
and U3018 (N_3018,N_2580,N_2546);
nor U3019 (N_3019,N_2675,N_2880);
nor U3020 (N_3020,N_2720,N_2903);
xor U3021 (N_3021,N_2544,N_2939);
or U3022 (N_3022,N_2637,N_2564);
xnor U3023 (N_3023,N_2557,N_2819);
or U3024 (N_3024,N_2562,N_2700);
xor U3025 (N_3025,N_2777,N_2914);
xor U3026 (N_3026,N_2521,N_2855);
nor U3027 (N_3027,N_2683,N_2917);
xnor U3028 (N_3028,N_2600,N_2595);
nor U3029 (N_3029,N_2786,N_2663);
xor U3030 (N_3030,N_2862,N_2826);
nand U3031 (N_3031,N_2995,N_2886);
nor U3032 (N_3032,N_2962,N_2761);
and U3033 (N_3033,N_2568,N_2757);
or U3034 (N_3034,N_2778,N_2714);
xor U3035 (N_3035,N_2971,N_2835);
xor U3036 (N_3036,N_2759,N_2541);
or U3037 (N_3037,N_2905,N_2690);
and U3038 (N_3038,N_2642,N_2922);
xor U3039 (N_3039,N_2705,N_2594);
nand U3040 (N_3040,N_2813,N_2678);
or U3041 (N_3041,N_2692,N_2709);
nand U3042 (N_3042,N_2861,N_2624);
and U3043 (N_3043,N_2571,N_2728);
or U3044 (N_3044,N_2770,N_2756);
and U3045 (N_3045,N_2574,N_2873);
nor U3046 (N_3046,N_2716,N_2741);
and U3047 (N_3047,N_2876,N_2581);
xor U3048 (N_3048,N_2653,N_2506);
and U3049 (N_3049,N_2850,N_2816);
nand U3050 (N_3050,N_2689,N_2844);
or U3051 (N_3051,N_2871,N_2762);
nor U3052 (N_3052,N_2864,N_2978);
nor U3053 (N_3053,N_2996,N_2824);
or U3054 (N_3054,N_2619,N_2805);
and U3055 (N_3055,N_2821,N_2935);
and U3056 (N_3056,N_2740,N_2773);
nor U3057 (N_3057,N_2578,N_2815);
or U3058 (N_3058,N_2660,N_2645);
nand U3059 (N_3059,N_2948,N_2934);
nand U3060 (N_3060,N_2860,N_2888);
xor U3061 (N_3061,N_2615,N_2901);
or U3062 (N_3062,N_2500,N_2526);
nand U3063 (N_3063,N_2516,N_2814);
or U3064 (N_3064,N_2721,N_2603);
and U3065 (N_3065,N_2785,N_2572);
nor U3066 (N_3066,N_2522,N_2735);
and U3067 (N_3067,N_2902,N_2950);
nor U3068 (N_3068,N_2984,N_2547);
and U3069 (N_3069,N_2836,N_2953);
or U3070 (N_3070,N_2588,N_2837);
xnor U3071 (N_3071,N_2599,N_2664);
or U3072 (N_3072,N_2587,N_2839);
xnor U3073 (N_3073,N_2527,N_2609);
or U3074 (N_3074,N_2993,N_2617);
and U3075 (N_3075,N_2523,N_2991);
xnor U3076 (N_3076,N_2717,N_2753);
nand U3077 (N_3077,N_2992,N_2936);
xnor U3078 (N_3078,N_2712,N_2845);
and U3079 (N_3079,N_2630,N_2507);
and U3080 (N_3080,N_2877,N_2811);
and U3081 (N_3081,N_2517,N_2820);
xnor U3082 (N_3082,N_2928,N_2998);
and U3083 (N_3083,N_2997,N_2818);
xnor U3084 (N_3084,N_2649,N_2970);
or U3085 (N_3085,N_2552,N_2966);
xnor U3086 (N_3086,N_2627,N_2560);
xnor U3087 (N_3087,N_2754,N_2648);
nor U3088 (N_3088,N_2865,N_2921);
and U3089 (N_3089,N_2597,N_2592);
nor U3090 (N_3090,N_2632,N_2658);
nor U3091 (N_3091,N_2904,N_2909);
nor U3092 (N_3092,N_2726,N_2608);
or U3093 (N_3093,N_2622,N_2682);
nor U3094 (N_3094,N_2535,N_2673);
and U3095 (N_3095,N_2884,N_2528);
and U3096 (N_3096,N_2881,N_2687);
nand U3097 (N_3097,N_2937,N_2787);
or U3098 (N_3098,N_2979,N_2791);
or U3099 (N_3099,N_2671,N_2987);
and U3100 (N_3100,N_2822,N_2504);
nand U3101 (N_3101,N_2707,N_2736);
and U3102 (N_3102,N_2929,N_2532);
nor U3103 (N_3103,N_2503,N_2825);
and U3104 (N_3104,N_2722,N_2573);
nor U3105 (N_3105,N_2974,N_2679);
xnor U3106 (N_3106,N_2932,N_2764);
nand U3107 (N_3107,N_2925,N_2512);
nand U3108 (N_3108,N_2633,N_2755);
nand U3109 (N_3109,N_2563,N_2897);
and U3110 (N_3110,N_2924,N_2866);
xnor U3111 (N_3111,N_2843,N_2605);
xnor U3112 (N_3112,N_2575,N_2559);
or U3113 (N_3113,N_2746,N_2999);
xor U3114 (N_3114,N_2807,N_2894);
or U3115 (N_3115,N_2960,N_2976);
nor U3116 (N_3116,N_2856,N_2616);
nand U3117 (N_3117,N_2907,N_2550);
nand U3118 (N_3118,N_2601,N_2688);
or U3119 (N_3119,N_2988,N_2567);
or U3120 (N_3120,N_2666,N_2579);
xnor U3121 (N_3121,N_2704,N_2919);
nand U3122 (N_3122,N_2795,N_2829);
nand U3123 (N_3123,N_2667,N_2920);
xnor U3124 (N_3124,N_2607,N_2885);
or U3125 (N_3125,N_2593,N_2708);
and U3126 (N_3126,N_2725,N_2784);
or U3127 (N_3127,N_2576,N_2849);
nor U3128 (N_3128,N_2697,N_2834);
and U3129 (N_3129,N_2792,N_2539);
xnor U3130 (N_3130,N_2662,N_2951);
nand U3131 (N_3131,N_2681,N_2803);
nand U3132 (N_3132,N_2906,N_2900);
and U3133 (N_3133,N_2765,N_2955);
xnor U3134 (N_3134,N_2577,N_2731);
xor U3135 (N_3135,N_2968,N_2859);
nand U3136 (N_3136,N_2801,N_2628);
nor U3137 (N_3137,N_2646,N_2680);
and U3138 (N_3138,N_2706,N_2651);
nand U3139 (N_3139,N_2832,N_2878);
and U3140 (N_3140,N_2827,N_2779);
and U3141 (N_3141,N_2732,N_2661);
or U3142 (N_3142,N_2613,N_2916);
xnor U3143 (N_3143,N_2769,N_2911);
xor U3144 (N_3144,N_2655,N_2640);
xor U3145 (N_3145,N_2794,N_2879);
and U3146 (N_3146,N_2699,N_2959);
xor U3147 (N_3147,N_2954,N_2729);
xor U3148 (N_3148,N_2691,N_2763);
xnor U3149 (N_3149,N_2684,N_2542);
nor U3150 (N_3150,N_2898,N_2808);
and U3151 (N_3151,N_2851,N_2551);
xor U3152 (N_3152,N_2915,N_2533);
or U3153 (N_3153,N_2830,N_2793);
and U3154 (N_3154,N_2589,N_2771);
nor U3155 (N_3155,N_2798,N_2782);
and U3156 (N_3156,N_2685,N_2641);
nor U3157 (N_3157,N_2980,N_2812);
xnor U3158 (N_3158,N_2872,N_2739);
nand U3159 (N_3159,N_2969,N_2621);
or U3160 (N_3160,N_2702,N_2990);
nand U3161 (N_3161,N_2511,N_2940);
nand U3162 (N_3162,N_2797,N_2644);
or U3163 (N_3163,N_2854,N_2538);
xor U3164 (N_3164,N_2891,N_2910);
or U3165 (N_3165,N_2841,N_2513);
xnor U3166 (N_3166,N_2636,N_2867);
xnor U3167 (N_3167,N_2887,N_2927);
xor U3168 (N_3168,N_2515,N_2745);
nand U3169 (N_3169,N_2788,N_2781);
nor U3170 (N_3170,N_2670,N_2566);
xnor U3171 (N_3171,N_2549,N_2514);
and U3172 (N_3172,N_2847,N_2870);
or U3173 (N_3173,N_2558,N_2519);
nand U3174 (N_3174,N_2809,N_2677);
or U3175 (N_3175,N_2749,N_2751);
nand U3176 (N_3176,N_2967,N_2652);
xnor U3177 (N_3177,N_2596,N_2548);
and U3178 (N_3178,N_2711,N_2852);
and U3179 (N_3179,N_2623,N_2570);
nor U3180 (N_3180,N_2650,N_2895);
and U3181 (N_3181,N_2973,N_2947);
or U3182 (N_3182,N_2530,N_2804);
nand U3183 (N_3183,N_2767,N_2738);
nand U3184 (N_3184,N_2858,N_2776);
nand U3185 (N_3185,N_2529,N_2734);
and U3186 (N_3186,N_2853,N_2744);
nand U3187 (N_3187,N_2802,N_2718);
and U3188 (N_3188,N_2840,N_2620);
or U3189 (N_3189,N_2701,N_2719);
nand U3190 (N_3190,N_2817,N_2657);
and U3191 (N_3191,N_2989,N_2534);
nor U3192 (N_3192,N_2509,N_2882);
xor U3193 (N_3193,N_2654,N_2508);
xnor U3194 (N_3194,N_2946,N_2583);
nor U3195 (N_3195,N_2696,N_2750);
or U3196 (N_3196,N_2833,N_2913);
and U3197 (N_3197,N_2554,N_2944);
nor U3198 (N_3198,N_2505,N_2669);
and U3199 (N_3199,N_2889,N_2510);
nand U3200 (N_3200,N_2724,N_2635);
xnor U3201 (N_3201,N_2659,N_2598);
nor U3202 (N_3202,N_2604,N_2612);
and U3203 (N_3203,N_2863,N_2977);
nor U3204 (N_3204,N_2730,N_2676);
nor U3205 (N_3205,N_2629,N_2896);
or U3206 (N_3206,N_2602,N_2930);
nand U3207 (N_3207,N_2626,N_2772);
nand U3208 (N_3208,N_2958,N_2672);
xor U3209 (N_3209,N_2715,N_2828);
xor U3210 (N_3210,N_2983,N_2565);
nand U3211 (N_3211,N_2868,N_2892);
and U3212 (N_3212,N_2752,N_2965);
and U3213 (N_3213,N_2838,N_2727);
and U3214 (N_3214,N_2748,N_2790);
or U3215 (N_3215,N_2800,N_2899);
nor U3216 (N_3216,N_2710,N_2957);
and U3217 (N_3217,N_2985,N_2606);
nand U3218 (N_3218,N_2768,N_2569);
and U3219 (N_3219,N_2775,N_2918);
or U3220 (N_3220,N_2986,N_2625);
xnor U3221 (N_3221,N_2810,N_2733);
or U3222 (N_3222,N_2869,N_2799);
xnor U3223 (N_3223,N_2536,N_2923);
xor U3224 (N_3224,N_2938,N_2668);
and U3225 (N_3225,N_2883,N_2555);
or U3226 (N_3226,N_2796,N_2972);
or U3227 (N_3227,N_2952,N_2524);
xor U3228 (N_3228,N_2943,N_2525);
nor U3229 (N_3229,N_2846,N_2553);
nand U3230 (N_3230,N_2518,N_2823);
or U3231 (N_3231,N_2760,N_2618);
and U3232 (N_3232,N_2582,N_2806);
nand U3233 (N_3233,N_2737,N_2766);
or U3234 (N_3234,N_2747,N_2961);
nor U3235 (N_3235,N_2502,N_2942);
and U3236 (N_3236,N_2674,N_2686);
nor U3237 (N_3237,N_2908,N_2857);
xnor U3238 (N_3238,N_2639,N_2590);
or U3239 (N_3239,N_2933,N_2994);
nor U3240 (N_3240,N_2694,N_2981);
or U3241 (N_3241,N_2695,N_2783);
nand U3242 (N_3242,N_2556,N_2610);
nand U3243 (N_3243,N_2540,N_2537);
nand U3244 (N_3244,N_2743,N_2964);
and U3245 (N_3245,N_2758,N_2713);
and U3246 (N_3246,N_2742,N_2931);
xor U3247 (N_3247,N_2586,N_2949);
xor U3248 (N_3248,N_2831,N_2698);
nor U3249 (N_3249,N_2631,N_2963);
and U3250 (N_3250,N_2709,N_2779);
xor U3251 (N_3251,N_2500,N_2795);
xor U3252 (N_3252,N_2892,N_2664);
or U3253 (N_3253,N_2849,N_2565);
or U3254 (N_3254,N_2751,N_2738);
nor U3255 (N_3255,N_2684,N_2613);
and U3256 (N_3256,N_2621,N_2576);
or U3257 (N_3257,N_2513,N_2554);
nor U3258 (N_3258,N_2552,N_2921);
nand U3259 (N_3259,N_2816,N_2596);
or U3260 (N_3260,N_2627,N_2566);
or U3261 (N_3261,N_2772,N_2767);
or U3262 (N_3262,N_2913,N_2557);
xor U3263 (N_3263,N_2574,N_2585);
xor U3264 (N_3264,N_2811,N_2585);
xor U3265 (N_3265,N_2769,N_2577);
nor U3266 (N_3266,N_2537,N_2998);
xnor U3267 (N_3267,N_2903,N_2872);
xnor U3268 (N_3268,N_2504,N_2870);
or U3269 (N_3269,N_2506,N_2996);
or U3270 (N_3270,N_2881,N_2609);
and U3271 (N_3271,N_2859,N_2815);
nor U3272 (N_3272,N_2877,N_2552);
xnor U3273 (N_3273,N_2633,N_2636);
or U3274 (N_3274,N_2813,N_2857);
and U3275 (N_3275,N_2970,N_2531);
xor U3276 (N_3276,N_2617,N_2730);
nor U3277 (N_3277,N_2543,N_2671);
xor U3278 (N_3278,N_2735,N_2646);
nand U3279 (N_3279,N_2855,N_2718);
and U3280 (N_3280,N_2958,N_2553);
nor U3281 (N_3281,N_2802,N_2902);
nand U3282 (N_3282,N_2632,N_2822);
nand U3283 (N_3283,N_2852,N_2818);
xnor U3284 (N_3284,N_2810,N_2821);
and U3285 (N_3285,N_2881,N_2936);
xnor U3286 (N_3286,N_2760,N_2985);
and U3287 (N_3287,N_2620,N_2855);
and U3288 (N_3288,N_2946,N_2939);
nor U3289 (N_3289,N_2650,N_2921);
and U3290 (N_3290,N_2599,N_2572);
nor U3291 (N_3291,N_2536,N_2769);
nand U3292 (N_3292,N_2615,N_2666);
nor U3293 (N_3293,N_2596,N_2868);
xor U3294 (N_3294,N_2720,N_2901);
nor U3295 (N_3295,N_2759,N_2932);
and U3296 (N_3296,N_2710,N_2956);
nand U3297 (N_3297,N_2700,N_2640);
nand U3298 (N_3298,N_2903,N_2937);
nor U3299 (N_3299,N_2787,N_2708);
nand U3300 (N_3300,N_2645,N_2940);
nand U3301 (N_3301,N_2744,N_2795);
nand U3302 (N_3302,N_2831,N_2856);
or U3303 (N_3303,N_2633,N_2681);
xor U3304 (N_3304,N_2958,N_2704);
nand U3305 (N_3305,N_2881,N_2920);
or U3306 (N_3306,N_2519,N_2684);
xor U3307 (N_3307,N_2947,N_2897);
xnor U3308 (N_3308,N_2886,N_2981);
or U3309 (N_3309,N_2730,N_2665);
nand U3310 (N_3310,N_2570,N_2976);
or U3311 (N_3311,N_2996,N_2852);
or U3312 (N_3312,N_2595,N_2515);
or U3313 (N_3313,N_2926,N_2782);
and U3314 (N_3314,N_2677,N_2527);
nor U3315 (N_3315,N_2889,N_2925);
or U3316 (N_3316,N_2954,N_2565);
or U3317 (N_3317,N_2771,N_2651);
or U3318 (N_3318,N_2715,N_2800);
xnor U3319 (N_3319,N_2582,N_2525);
or U3320 (N_3320,N_2679,N_2837);
nand U3321 (N_3321,N_2593,N_2508);
and U3322 (N_3322,N_2543,N_2875);
xnor U3323 (N_3323,N_2846,N_2829);
nand U3324 (N_3324,N_2894,N_2564);
nand U3325 (N_3325,N_2846,N_2876);
xnor U3326 (N_3326,N_2734,N_2595);
nor U3327 (N_3327,N_2675,N_2627);
and U3328 (N_3328,N_2727,N_2935);
xor U3329 (N_3329,N_2724,N_2977);
nor U3330 (N_3330,N_2537,N_2832);
and U3331 (N_3331,N_2858,N_2576);
nand U3332 (N_3332,N_2908,N_2656);
nor U3333 (N_3333,N_2543,N_2582);
and U3334 (N_3334,N_2900,N_2568);
xnor U3335 (N_3335,N_2535,N_2894);
xor U3336 (N_3336,N_2706,N_2551);
and U3337 (N_3337,N_2735,N_2795);
xor U3338 (N_3338,N_2562,N_2667);
nor U3339 (N_3339,N_2526,N_2586);
and U3340 (N_3340,N_2789,N_2796);
or U3341 (N_3341,N_2800,N_2815);
nand U3342 (N_3342,N_2687,N_2974);
and U3343 (N_3343,N_2944,N_2655);
nor U3344 (N_3344,N_2861,N_2695);
nor U3345 (N_3345,N_2597,N_2512);
or U3346 (N_3346,N_2615,N_2543);
nor U3347 (N_3347,N_2881,N_2536);
nor U3348 (N_3348,N_2701,N_2843);
nand U3349 (N_3349,N_2536,N_2518);
or U3350 (N_3350,N_2925,N_2775);
or U3351 (N_3351,N_2970,N_2519);
or U3352 (N_3352,N_2680,N_2700);
nand U3353 (N_3353,N_2926,N_2581);
nor U3354 (N_3354,N_2511,N_2623);
nand U3355 (N_3355,N_2885,N_2706);
nand U3356 (N_3356,N_2603,N_2955);
and U3357 (N_3357,N_2701,N_2769);
and U3358 (N_3358,N_2785,N_2772);
xor U3359 (N_3359,N_2734,N_2611);
nand U3360 (N_3360,N_2948,N_2505);
nor U3361 (N_3361,N_2992,N_2973);
and U3362 (N_3362,N_2593,N_2626);
nand U3363 (N_3363,N_2584,N_2995);
nand U3364 (N_3364,N_2636,N_2918);
nand U3365 (N_3365,N_2819,N_2675);
nand U3366 (N_3366,N_2950,N_2541);
xor U3367 (N_3367,N_2537,N_2796);
xnor U3368 (N_3368,N_2669,N_2732);
or U3369 (N_3369,N_2762,N_2739);
and U3370 (N_3370,N_2914,N_2920);
or U3371 (N_3371,N_2735,N_2680);
or U3372 (N_3372,N_2890,N_2769);
nor U3373 (N_3373,N_2979,N_2658);
xnor U3374 (N_3374,N_2890,N_2843);
nor U3375 (N_3375,N_2755,N_2866);
nand U3376 (N_3376,N_2833,N_2623);
xor U3377 (N_3377,N_2891,N_2923);
xnor U3378 (N_3378,N_2639,N_2886);
xnor U3379 (N_3379,N_2856,N_2590);
nand U3380 (N_3380,N_2645,N_2630);
and U3381 (N_3381,N_2963,N_2854);
and U3382 (N_3382,N_2679,N_2993);
xor U3383 (N_3383,N_2537,N_2689);
nand U3384 (N_3384,N_2614,N_2920);
xor U3385 (N_3385,N_2945,N_2576);
nand U3386 (N_3386,N_2665,N_2793);
nand U3387 (N_3387,N_2887,N_2708);
and U3388 (N_3388,N_2674,N_2949);
or U3389 (N_3389,N_2871,N_2944);
or U3390 (N_3390,N_2546,N_2916);
nand U3391 (N_3391,N_2680,N_2811);
nand U3392 (N_3392,N_2748,N_2888);
nand U3393 (N_3393,N_2791,N_2544);
or U3394 (N_3394,N_2807,N_2869);
nor U3395 (N_3395,N_2694,N_2774);
and U3396 (N_3396,N_2883,N_2867);
nor U3397 (N_3397,N_2999,N_2630);
xor U3398 (N_3398,N_2958,N_2526);
or U3399 (N_3399,N_2610,N_2548);
nand U3400 (N_3400,N_2797,N_2578);
xor U3401 (N_3401,N_2525,N_2593);
nand U3402 (N_3402,N_2725,N_2917);
nand U3403 (N_3403,N_2514,N_2873);
nand U3404 (N_3404,N_2695,N_2655);
xnor U3405 (N_3405,N_2763,N_2695);
or U3406 (N_3406,N_2833,N_2590);
nand U3407 (N_3407,N_2638,N_2937);
nand U3408 (N_3408,N_2901,N_2674);
xnor U3409 (N_3409,N_2581,N_2533);
and U3410 (N_3410,N_2673,N_2956);
xnor U3411 (N_3411,N_2642,N_2777);
nand U3412 (N_3412,N_2828,N_2688);
nor U3413 (N_3413,N_2929,N_2629);
nor U3414 (N_3414,N_2708,N_2577);
nor U3415 (N_3415,N_2969,N_2780);
or U3416 (N_3416,N_2835,N_2912);
nand U3417 (N_3417,N_2857,N_2986);
nor U3418 (N_3418,N_2808,N_2628);
xnor U3419 (N_3419,N_2746,N_2757);
and U3420 (N_3420,N_2553,N_2991);
nor U3421 (N_3421,N_2606,N_2672);
and U3422 (N_3422,N_2857,N_2764);
and U3423 (N_3423,N_2974,N_2806);
or U3424 (N_3424,N_2932,N_2781);
or U3425 (N_3425,N_2658,N_2807);
and U3426 (N_3426,N_2593,N_2669);
nand U3427 (N_3427,N_2716,N_2897);
xnor U3428 (N_3428,N_2748,N_2995);
nor U3429 (N_3429,N_2594,N_2685);
or U3430 (N_3430,N_2851,N_2918);
nand U3431 (N_3431,N_2578,N_2604);
nand U3432 (N_3432,N_2770,N_2607);
nand U3433 (N_3433,N_2743,N_2582);
nor U3434 (N_3434,N_2883,N_2780);
nand U3435 (N_3435,N_2599,N_2792);
xor U3436 (N_3436,N_2957,N_2700);
nor U3437 (N_3437,N_2836,N_2630);
xor U3438 (N_3438,N_2903,N_2718);
or U3439 (N_3439,N_2808,N_2812);
and U3440 (N_3440,N_2618,N_2541);
and U3441 (N_3441,N_2731,N_2959);
nor U3442 (N_3442,N_2565,N_2908);
or U3443 (N_3443,N_2558,N_2707);
xnor U3444 (N_3444,N_2785,N_2589);
xnor U3445 (N_3445,N_2530,N_2987);
or U3446 (N_3446,N_2918,N_2797);
xor U3447 (N_3447,N_2968,N_2692);
xor U3448 (N_3448,N_2987,N_2890);
xor U3449 (N_3449,N_2956,N_2662);
or U3450 (N_3450,N_2812,N_2964);
or U3451 (N_3451,N_2921,N_2711);
or U3452 (N_3452,N_2849,N_2667);
nor U3453 (N_3453,N_2879,N_2986);
xor U3454 (N_3454,N_2678,N_2731);
nor U3455 (N_3455,N_2605,N_2997);
or U3456 (N_3456,N_2764,N_2713);
nand U3457 (N_3457,N_2855,N_2843);
or U3458 (N_3458,N_2913,N_2837);
or U3459 (N_3459,N_2988,N_2571);
and U3460 (N_3460,N_2648,N_2798);
and U3461 (N_3461,N_2720,N_2588);
and U3462 (N_3462,N_2511,N_2580);
nand U3463 (N_3463,N_2835,N_2904);
xnor U3464 (N_3464,N_2506,N_2528);
nand U3465 (N_3465,N_2846,N_2542);
or U3466 (N_3466,N_2595,N_2802);
nand U3467 (N_3467,N_2987,N_2646);
nand U3468 (N_3468,N_2590,N_2897);
or U3469 (N_3469,N_2835,N_2716);
xor U3470 (N_3470,N_2819,N_2861);
or U3471 (N_3471,N_2532,N_2708);
nor U3472 (N_3472,N_2994,N_2888);
nand U3473 (N_3473,N_2727,N_2847);
nand U3474 (N_3474,N_2779,N_2683);
nor U3475 (N_3475,N_2568,N_2813);
and U3476 (N_3476,N_2645,N_2814);
nor U3477 (N_3477,N_2587,N_2926);
and U3478 (N_3478,N_2859,N_2836);
and U3479 (N_3479,N_2842,N_2896);
nor U3480 (N_3480,N_2808,N_2881);
or U3481 (N_3481,N_2535,N_2791);
nor U3482 (N_3482,N_2599,N_2658);
or U3483 (N_3483,N_2724,N_2967);
nor U3484 (N_3484,N_2730,N_2744);
xnor U3485 (N_3485,N_2812,N_2721);
xor U3486 (N_3486,N_2732,N_2533);
and U3487 (N_3487,N_2702,N_2545);
and U3488 (N_3488,N_2759,N_2831);
or U3489 (N_3489,N_2641,N_2691);
or U3490 (N_3490,N_2676,N_2836);
or U3491 (N_3491,N_2556,N_2580);
or U3492 (N_3492,N_2947,N_2891);
or U3493 (N_3493,N_2510,N_2660);
nand U3494 (N_3494,N_2976,N_2649);
or U3495 (N_3495,N_2744,N_2864);
or U3496 (N_3496,N_2791,N_2848);
xor U3497 (N_3497,N_2754,N_2859);
and U3498 (N_3498,N_2890,N_2854);
xor U3499 (N_3499,N_2947,N_2794);
or U3500 (N_3500,N_3162,N_3264);
nand U3501 (N_3501,N_3132,N_3265);
and U3502 (N_3502,N_3401,N_3225);
nor U3503 (N_3503,N_3087,N_3209);
or U3504 (N_3504,N_3484,N_3410);
and U3505 (N_3505,N_3421,N_3324);
and U3506 (N_3506,N_3081,N_3373);
or U3507 (N_3507,N_3221,N_3359);
and U3508 (N_3508,N_3153,N_3305);
and U3509 (N_3509,N_3455,N_3480);
nor U3510 (N_3510,N_3156,N_3267);
nand U3511 (N_3511,N_3037,N_3031);
nor U3512 (N_3512,N_3308,N_3251);
nand U3513 (N_3513,N_3317,N_3263);
or U3514 (N_3514,N_3366,N_3259);
nor U3515 (N_3515,N_3417,N_3041);
nand U3516 (N_3516,N_3312,N_3282);
xnor U3517 (N_3517,N_3418,N_3186);
and U3518 (N_3518,N_3059,N_3285);
nand U3519 (N_3519,N_3304,N_3451);
nand U3520 (N_3520,N_3495,N_3077);
and U3521 (N_3521,N_3217,N_3065);
and U3522 (N_3522,N_3486,N_3235);
and U3523 (N_3523,N_3050,N_3319);
nor U3524 (N_3524,N_3361,N_3136);
or U3525 (N_3525,N_3159,N_3039);
nand U3526 (N_3526,N_3262,N_3015);
and U3527 (N_3527,N_3320,N_3470);
nor U3528 (N_3528,N_3405,N_3155);
and U3529 (N_3529,N_3193,N_3295);
nor U3530 (N_3530,N_3169,N_3390);
nor U3531 (N_3531,N_3211,N_3073);
or U3532 (N_3532,N_3404,N_3271);
and U3533 (N_3533,N_3190,N_3161);
nor U3534 (N_3534,N_3179,N_3110);
and U3535 (N_3535,N_3004,N_3042);
or U3536 (N_3536,N_3465,N_3227);
xor U3537 (N_3537,N_3009,N_3206);
and U3538 (N_3538,N_3184,N_3007);
or U3539 (N_3539,N_3144,N_3414);
and U3540 (N_3540,N_3198,N_3102);
nor U3541 (N_3541,N_3469,N_3456);
or U3542 (N_3542,N_3107,N_3177);
xor U3543 (N_3543,N_3071,N_3115);
nor U3544 (N_3544,N_3082,N_3260);
or U3545 (N_3545,N_3049,N_3446);
or U3546 (N_3546,N_3488,N_3151);
xor U3547 (N_3547,N_3038,N_3109);
and U3548 (N_3548,N_3284,N_3386);
or U3549 (N_3549,N_3377,N_3126);
and U3550 (N_3550,N_3388,N_3306);
and U3551 (N_3551,N_3105,N_3220);
xnor U3552 (N_3552,N_3234,N_3463);
nand U3553 (N_3553,N_3230,N_3160);
and U3554 (N_3554,N_3164,N_3340);
xor U3555 (N_3555,N_3076,N_3316);
or U3556 (N_3556,N_3165,N_3182);
or U3557 (N_3557,N_3010,N_3497);
nor U3558 (N_3558,N_3123,N_3172);
xor U3559 (N_3559,N_3084,N_3429);
xor U3560 (N_3560,N_3171,N_3074);
xnor U3561 (N_3561,N_3166,N_3315);
and U3562 (N_3562,N_3419,N_3427);
nand U3563 (N_3563,N_3134,N_3464);
or U3564 (N_3564,N_3467,N_3492);
nand U3565 (N_3565,N_3149,N_3033);
nand U3566 (N_3566,N_3482,N_3348);
and U3567 (N_3567,N_3409,N_3300);
nand U3568 (N_3568,N_3310,N_3239);
and U3569 (N_3569,N_3002,N_3104);
xnor U3570 (N_3570,N_3222,N_3301);
nor U3571 (N_3571,N_3453,N_3238);
and U3572 (N_3572,N_3422,N_3428);
nand U3573 (N_3573,N_3406,N_3399);
or U3574 (N_3574,N_3273,N_3266);
nor U3575 (N_3575,N_3120,N_3474);
and U3576 (N_3576,N_3337,N_3342);
and U3577 (N_3577,N_3122,N_3085);
and U3578 (N_3578,N_3255,N_3344);
or U3579 (N_3579,N_3350,N_3243);
and U3580 (N_3580,N_3472,N_3437);
and U3581 (N_3581,N_3351,N_3100);
or U3582 (N_3582,N_3261,N_3139);
or U3583 (N_3583,N_3152,N_3311);
nand U3584 (N_3584,N_3420,N_3116);
and U3585 (N_3585,N_3064,N_3332);
nor U3586 (N_3586,N_3281,N_3449);
or U3587 (N_3587,N_3097,N_3157);
and U3588 (N_3588,N_3011,N_3147);
or U3589 (N_3589,N_3489,N_3223);
xnor U3590 (N_3590,N_3207,N_3013);
nand U3591 (N_3591,N_3499,N_3313);
and U3592 (N_3592,N_3103,N_3204);
and U3593 (N_3593,N_3400,N_3345);
xnor U3594 (N_3594,N_3016,N_3445);
xnor U3595 (N_3595,N_3188,N_3240);
and U3596 (N_3596,N_3170,N_3133);
nand U3597 (N_3597,N_3258,N_3127);
nor U3598 (N_3598,N_3358,N_3382);
and U3599 (N_3599,N_3490,N_3403);
xnor U3600 (N_3600,N_3444,N_3117);
nand U3601 (N_3601,N_3473,N_3331);
or U3602 (N_3602,N_3346,N_3001);
xor U3603 (N_3603,N_3062,N_3121);
or U3604 (N_3604,N_3129,N_3195);
or U3605 (N_3605,N_3466,N_3236);
or U3606 (N_3606,N_3462,N_3280);
xnor U3607 (N_3607,N_3086,N_3439);
xnor U3608 (N_3608,N_3199,N_3289);
nand U3609 (N_3609,N_3079,N_3035);
nand U3610 (N_3610,N_3231,N_3216);
xor U3611 (N_3611,N_3232,N_3075);
nand U3612 (N_3612,N_3343,N_3355);
or U3613 (N_3613,N_3214,N_3047);
or U3614 (N_3614,N_3443,N_3440);
nor U3615 (N_3615,N_3070,N_3416);
and U3616 (N_3616,N_3286,N_3391);
and U3617 (N_3617,N_3108,N_3349);
nand U3618 (N_3618,N_3402,N_3352);
xnor U3619 (N_3619,N_3131,N_3299);
nand U3620 (N_3620,N_3094,N_3442);
nor U3621 (N_3621,N_3244,N_3224);
xor U3622 (N_3622,N_3425,N_3360);
xnor U3623 (N_3623,N_3053,N_3118);
and U3624 (N_3624,N_3183,N_3392);
xnor U3625 (N_3625,N_3329,N_3202);
nor U3626 (N_3626,N_3479,N_3093);
and U3627 (N_3627,N_3297,N_3369);
nand U3628 (N_3628,N_3432,N_3130);
and U3629 (N_3629,N_3174,N_3438);
or U3630 (N_3630,N_3458,N_3175);
or U3631 (N_3631,N_3246,N_3447);
nor U3632 (N_3632,N_3226,N_3167);
nand U3633 (N_3633,N_3242,N_3278);
xor U3634 (N_3634,N_3066,N_3080);
or U3635 (N_3635,N_3413,N_3368);
or U3636 (N_3636,N_3005,N_3022);
nand U3637 (N_3637,N_3367,N_3485);
nor U3638 (N_3638,N_3253,N_3212);
xnor U3639 (N_3639,N_3483,N_3218);
nand U3640 (N_3640,N_3203,N_3378);
nor U3641 (N_3641,N_3487,N_3326);
nor U3642 (N_3642,N_3335,N_3434);
nand U3643 (N_3643,N_3114,N_3051);
and U3644 (N_3644,N_3000,N_3208);
and U3645 (N_3645,N_3370,N_3277);
or U3646 (N_3646,N_3189,N_3090);
nor U3647 (N_3647,N_3385,N_3135);
nand U3648 (N_3648,N_3112,N_3288);
nor U3649 (N_3649,N_3063,N_3494);
nand U3650 (N_3650,N_3389,N_3101);
nor U3651 (N_3651,N_3096,N_3394);
and U3652 (N_3652,N_3459,N_3396);
or U3653 (N_3653,N_3054,N_3380);
xnor U3654 (N_3654,N_3347,N_3374);
nand U3655 (N_3655,N_3338,N_3365);
nand U3656 (N_3656,N_3393,N_3142);
or U3657 (N_3657,N_3026,N_3468);
nand U3658 (N_3658,N_3137,N_3356);
nand U3659 (N_3659,N_3012,N_3061);
or U3660 (N_3660,N_3032,N_3387);
or U3661 (N_3661,N_3200,N_3291);
and U3662 (N_3662,N_3491,N_3302);
nor U3663 (N_3663,N_3197,N_3067);
xnor U3664 (N_3664,N_3248,N_3426);
xnor U3665 (N_3665,N_3014,N_3268);
or U3666 (N_3666,N_3191,N_3254);
nor U3667 (N_3667,N_3296,N_3353);
xnor U3668 (N_3668,N_3364,N_3415);
xor U3669 (N_3669,N_3287,N_3140);
and U3670 (N_3670,N_3150,N_3196);
nor U3671 (N_3671,N_3215,N_3325);
nand U3672 (N_3672,N_3017,N_3292);
and U3673 (N_3673,N_3028,N_3036);
or U3674 (N_3674,N_3412,N_3057);
nand U3675 (N_3675,N_3341,N_3431);
nand U3676 (N_3676,N_3092,N_3052);
or U3677 (N_3677,N_3457,N_3233);
xnor U3678 (N_3678,N_3424,N_3141);
and U3679 (N_3679,N_3083,N_3187);
nor U3680 (N_3680,N_3241,N_3176);
nand U3681 (N_3681,N_3219,N_3398);
or U3682 (N_3682,N_3269,N_3397);
xor U3683 (N_3683,N_3498,N_3068);
and U3684 (N_3684,N_3481,N_3072);
nand U3685 (N_3685,N_3069,N_3247);
xor U3686 (N_3686,N_3168,N_3008);
xnor U3687 (N_3687,N_3095,N_3383);
nand U3688 (N_3688,N_3205,N_3452);
xnor U3689 (N_3689,N_3314,N_3138);
xor U3690 (N_3690,N_3275,N_3148);
nor U3691 (N_3691,N_3475,N_3256);
and U3692 (N_3692,N_3146,N_3328);
nand U3693 (N_3693,N_3143,N_3357);
xor U3694 (N_3694,N_3089,N_3030);
and U3695 (N_3695,N_3124,N_3270);
xor U3696 (N_3696,N_3323,N_3379);
or U3697 (N_3697,N_3433,N_3372);
nor U3698 (N_3698,N_3376,N_3336);
xnor U3699 (N_3699,N_3245,N_3318);
xnor U3700 (N_3700,N_3043,N_3290);
xor U3701 (N_3701,N_3003,N_3294);
and U3702 (N_3702,N_3023,N_3249);
nor U3703 (N_3703,N_3321,N_3450);
nor U3704 (N_3704,N_3435,N_3471);
nand U3705 (N_3705,N_3430,N_3154);
nand U3706 (N_3706,N_3213,N_3363);
xor U3707 (N_3707,N_3252,N_3210);
or U3708 (N_3708,N_3185,N_3309);
and U3709 (N_3709,N_3322,N_3091);
nor U3710 (N_3710,N_3060,N_3045);
xor U3711 (N_3711,N_3362,N_3034);
xnor U3712 (N_3712,N_3478,N_3411);
and U3713 (N_3713,N_3111,N_3044);
nor U3714 (N_3714,N_3407,N_3078);
xor U3715 (N_3715,N_3441,N_3293);
or U3716 (N_3716,N_3099,N_3119);
or U3717 (N_3717,N_3476,N_3493);
nor U3718 (N_3718,N_3145,N_3283);
xnor U3719 (N_3719,N_3496,N_3025);
xor U3720 (N_3720,N_3029,N_3040);
nand U3721 (N_3721,N_3448,N_3019);
xor U3722 (N_3722,N_3113,N_3381);
and U3723 (N_3723,N_3272,N_3454);
and U3724 (N_3724,N_3327,N_3354);
and U3725 (N_3725,N_3178,N_3021);
xnor U3726 (N_3726,N_3228,N_3307);
and U3727 (N_3727,N_3056,N_3181);
xor U3728 (N_3728,N_3384,N_3194);
nor U3729 (N_3729,N_3173,N_3461);
or U3730 (N_3730,N_3020,N_3276);
nand U3731 (N_3731,N_3477,N_3303);
xnor U3732 (N_3732,N_3250,N_3279);
xnor U3733 (N_3733,N_3055,N_3375);
xor U3734 (N_3734,N_3024,N_3018);
or U3735 (N_3735,N_3006,N_3334);
nand U3736 (N_3736,N_3098,N_3058);
or U3737 (N_3737,N_3128,N_3274);
or U3738 (N_3738,N_3395,N_3163);
nor U3739 (N_3739,N_3423,N_3371);
or U3740 (N_3740,N_3046,N_3330);
xor U3741 (N_3741,N_3106,N_3257);
nand U3742 (N_3742,N_3460,N_3237);
or U3743 (N_3743,N_3158,N_3048);
and U3744 (N_3744,N_3408,N_3088);
xor U3745 (N_3745,N_3298,N_3339);
nor U3746 (N_3746,N_3229,N_3125);
xnor U3747 (N_3747,N_3180,N_3333);
nor U3748 (N_3748,N_3201,N_3436);
or U3749 (N_3749,N_3027,N_3192);
or U3750 (N_3750,N_3449,N_3240);
nor U3751 (N_3751,N_3136,N_3379);
or U3752 (N_3752,N_3448,N_3260);
or U3753 (N_3753,N_3293,N_3443);
xnor U3754 (N_3754,N_3247,N_3028);
or U3755 (N_3755,N_3414,N_3130);
and U3756 (N_3756,N_3169,N_3148);
nor U3757 (N_3757,N_3389,N_3031);
and U3758 (N_3758,N_3425,N_3493);
nor U3759 (N_3759,N_3462,N_3199);
or U3760 (N_3760,N_3105,N_3262);
nand U3761 (N_3761,N_3132,N_3177);
nand U3762 (N_3762,N_3350,N_3253);
xnor U3763 (N_3763,N_3328,N_3297);
and U3764 (N_3764,N_3037,N_3192);
nand U3765 (N_3765,N_3074,N_3105);
and U3766 (N_3766,N_3195,N_3271);
or U3767 (N_3767,N_3238,N_3329);
nand U3768 (N_3768,N_3109,N_3265);
nand U3769 (N_3769,N_3180,N_3378);
and U3770 (N_3770,N_3437,N_3073);
xnor U3771 (N_3771,N_3251,N_3177);
or U3772 (N_3772,N_3139,N_3362);
and U3773 (N_3773,N_3430,N_3417);
nor U3774 (N_3774,N_3103,N_3396);
nor U3775 (N_3775,N_3223,N_3378);
or U3776 (N_3776,N_3424,N_3078);
nand U3777 (N_3777,N_3302,N_3374);
nand U3778 (N_3778,N_3024,N_3417);
nand U3779 (N_3779,N_3217,N_3122);
and U3780 (N_3780,N_3210,N_3377);
nand U3781 (N_3781,N_3185,N_3211);
and U3782 (N_3782,N_3262,N_3205);
and U3783 (N_3783,N_3235,N_3428);
xnor U3784 (N_3784,N_3301,N_3228);
and U3785 (N_3785,N_3130,N_3298);
nand U3786 (N_3786,N_3230,N_3410);
or U3787 (N_3787,N_3321,N_3388);
xor U3788 (N_3788,N_3312,N_3410);
xor U3789 (N_3789,N_3434,N_3084);
or U3790 (N_3790,N_3021,N_3492);
and U3791 (N_3791,N_3153,N_3187);
nor U3792 (N_3792,N_3155,N_3350);
and U3793 (N_3793,N_3126,N_3057);
and U3794 (N_3794,N_3497,N_3328);
or U3795 (N_3795,N_3479,N_3268);
or U3796 (N_3796,N_3331,N_3263);
or U3797 (N_3797,N_3484,N_3354);
nand U3798 (N_3798,N_3044,N_3496);
nor U3799 (N_3799,N_3325,N_3059);
or U3800 (N_3800,N_3219,N_3092);
xnor U3801 (N_3801,N_3032,N_3490);
xnor U3802 (N_3802,N_3163,N_3313);
or U3803 (N_3803,N_3297,N_3065);
or U3804 (N_3804,N_3368,N_3211);
or U3805 (N_3805,N_3327,N_3263);
nor U3806 (N_3806,N_3425,N_3326);
or U3807 (N_3807,N_3050,N_3359);
xnor U3808 (N_3808,N_3009,N_3475);
and U3809 (N_3809,N_3375,N_3154);
nand U3810 (N_3810,N_3128,N_3173);
or U3811 (N_3811,N_3431,N_3138);
nor U3812 (N_3812,N_3239,N_3037);
nor U3813 (N_3813,N_3368,N_3221);
or U3814 (N_3814,N_3355,N_3103);
and U3815 (N_3815,N_3403,N_3460);
or U3816 (N_3816,N_3043,N_3087);
xor U3817 (N_3817,N_3070,N_3088);
nor U3818 (N_3818,N_3009,N_3490);
or U3819 (N_3819,N_3303,N_3220);
nand U3820 (N_3820,N_3279,N_3193);
nor U3821 (N_3821,N_3128,N_3007);
nor U3822 (N_3822,N_3196,N_3278);
nor U3823 (N_3823,N_3089,N_3309);
nand U3824 (N_3824,N_3213,N_3207);
or U3825 (N_3825,N_3426,N_3017);
or U3826 (N_3826,N_3417,N_3015);
xnor U3827 (N_3827,N_3279,N_3091);
or U3828 (N_3828,N_3323,N_3159);
and U3829 (N_3829,N_3362,N_3320);
or U3830 (N_3830,N_3319,N_3255);
nand U3831 (N_3831,N_3440,N_3159);
nand U3832 (N_3832,N_3473,N_3245);
or U3833 (N_3833,N_3141,N_3088);
nand U3834 (N_3834,N_3470,N_3168);
and U3835 (N_3835,N_3427,N_3256);
or U3836 (N_3836,N_3026,N_3018);
and U3837 (N_3837,N_3092,N_3225);
xor U3838 (N_3838,N_3128,N_3102);
xnor U3839 (N_3839,N_3230,N_3225);
nand U3840 (N_3840,N_3100,N_3369);
nand U3841 (N_3841,N_3326,N_3494);
xnor U3842 (N_3842,N_3343,N_3080);
nand U3843 (N_3843,N_3059,N_3001);
or U3844 (N_3844,N_3242,N_3383);
xnor U3845 (N_3845,N_3439,N_3373);
or U3846 (N_3846,N_3080,N_3180);
xnor U3847 (N_3847,N_3006,N_3275);
or U3848 (N_3848,N_3341,N_3429);
nand U3849 (N_3849,N_3375,N_3069);
nor U3850 (N_3850,N_3040,N_3264);
nand U3851 (N_3851,N_3313,N_3364);
and U3852 (N_3852,N_3259,N_3400);
nor U3853 (N_3853,N_3070,N_3019);
xnor U3854 (N_3854,N_3104,N_3102);
xnor U3855 (N_3855,N_3275,N_3147);
and U3856 (N_3856,N_3290,N_3136);
xor U3857 (N_3857,N_3016,N_3086);
nand U3858 (N_3858,N_3324,N_3320);
nand U3859 (N_3859,N_3461,N_3314);
xor U3860 (N_3860,N_3281,N_3210);
and U3861 (N_3861,N_3063,N_3466);
xnor U3862 (N_3862,N_3456,N_3425);
nor U3863 (N_3863,N_3123,N_3012);
xnor U3864 (N_3864,N_3262,N_3450);
and U3865 (N_3865,N_3421,N_3107);
xor U3866 (N_3866,N_3331,N_3286);
or U3867 (N_3867,N_3335,N_3160);
nand U3868 (N_3868,N_3118,N_3078);
nand U3869 (N_3869,N_3353,N_3415);
or U3870 (N_3870,N_3425,N_3486);
and U3871 (N_3871,N_3104,N_3393);
nor U3872 (N_3872,N_3450,N_3040);
nand U3873 (N_3873,N_3395,N_3239);
nand U3874 (N_3874,N_3185,N_3357);
and U3875 (N_3875,N_3139,N_3366);
nor U3876 (N_3876,N_3155,N_3487);
nor U3877 (N_3877,N_3080,N_3120);
and U3878 (N_3878,N_3058,N_3039);
nand U3879 (N_3879,N_3085,N_3010);
and U3880 (N_3880,N_3270,N_3242);
nand U3881 (N_3881,N_3410,N_3356);
and U3882 (N_3882,N_3421,N_3330);
or U3883 (N_3883,N_3096,N_3304);
nand U3884 (N_3884,N_3190,N_3122);
nand U3885 (N_3885,N_3161,N_3372);
and U3886 (N_3886,N_3332,N_3292);
and U3887 (N_3887,N_3121,N_3399);
xor U3888 (N_3888,N_3238,N_3498);
and U3889 (N_3889,N_3367,N_3424);
xor U3890 (N_3890,N_3205,N_3392);
and U3891 (N_3891,N_3014,N_3180);
and U3892 (N_3892,N_3252,N_3270);
xor U3893 (N_3893,N_3291,N_3228);
or U3894 (N_3894,N_3084,N_3331);
or U3895 (N_3895,N_3047,N_3365);
and U3896 (N_3896,N_3140,N_3227);
xnor U3897 (N_3897,N_3024,N_3149);
nand U3898 (N_3898,N_3086,N_3080);
nor U3899 (N_3899,N_3202,N_3189);
xnor U3900 (N_3900,N_3373,N_3482);
nor U3901 (N_3901,N_3390,N_3033);
xor U3902 (N_3902,N_3456,N_3026);
nor U3903 (N_3903,N_3290,N_3440);
or U3904 (N_3904,N_3373,N_3097);
xor U3905 (N_3905,N_3362,N_3401);
nor U3906 (N_3906,N_3138,N_3141);
nor U3907 (N_3907,N_3000,N_3264);
or U3908 (N_3908,N_3445,N_3243);
and U3909 (N_3909,N_3144,N_3443);
nand U3910 (N_3910,N_3413,N_3279);
xor U3911 (N_3911,N_3093,N_3158);
and U3912 (N_3912,N_3307,N_3432);
nand U3913 (N_3913,N_3372,N_3217);
and U3914 (N_3914,N_3244,N_3320);
or U3915 (N_3915,N_3117,N_3254);
xor U3916 (N_3916,N_3021,N_3465);
nor U3917 (N_3917,N_3380,N_3156);
nor U3918 (N_3918,N_3003,N_3078);
or U3919 (N_3919,N_3442,N_3305);
and U3920 (N_3920,N_3171,N_3498);
xnor U3921 (N_3921,N_3405,N_3315);
xor U3922 (N_3922,N_3384,N_3447);
nor U3923 (N_3923,N_3117,N_3136);
and U3924 (N_3924,N_3094,N_3227);
or U3925 (N_3925,N_3368,N_3021);
nand U3926 (N_3926,N_3447,N_3361);
xor U3927 (N_3927,N_3398,N_3005);
nand U3928 (N_3928,N_3232,N_3103);
and U3929 (N_3929,N_3451,N_3289);
or U3930 (N_3930,N_3005,N_3481);
nand U3931 (N_3931,N_3067,N_3096);
nor U3932 (N_3932,N_3200,N_3185);
xnor U3933 (N_3933,N_3498,N_3360);
nand U3934 (N_3934,N_3141,N_3015);
or U3935 (N_3935,N_3286,N_3344);
xor U3936 (N_3936,N_3242,N_3453);
or U3937 (N_3937,N_3482,N_3224);
nor U3938 (N_3938,N_3116,N_3347);
nand U3939 (N_3939,N_3228,N_3021);
or U3940 (N_3940,N_3272,N_3295);
xnor U3941 (N_3941,N_3369,N_3232);
nor U3942 (N_3942,N_3309,N_3446);
and U3943 (N_3943,N_3053,N_3046);
nor U3944 (N_3944,N_3463,N_3304);
and U3945 (N_3945,N_3307,N_3009);
nand U3946 (N_3946,N_3466,N_3100);
and U3947 (N_3947,N_3325,N_3212);
and U3948 (N_3948,N_3413,N_3264);
nor U3949 (N_3949,N_3081,N_3225);
nand U3950 (N_3950,N_3018,N_3196);
xnor U3951 (N_3951,N_3033,N_3401);
nor U3952 (N_3952,N_3367,N_3239);
or U3953 (N_3953,N_3018,N_3390);
nand U3954 (N_3954,N_3409,N_3057);
xor U3955 (N_3955,N_3472,N_3474);
xor U3956 (N_3956,N_3436,N_3302);
nand U3957 (N_3957,N_3425,N_3061);
nand U3958 (N_3958,N_3493,N_3025);
or U3959 (N_3959,N_3395,N_3406);
or U3960 (N_3960,N_3343,N_3498);
nand U3961 (N_3961,N_3038,N_3012);
xor U3962 (N_3962,N_3159,N_3040);
and U3963 (N_3963,N_3215,N_3129);
xnor U3964 (N_3964,N_3174,N_3045);
and U3965 (N_3965,N_3281,N_3345);
and U3966 (N_3966,N_3347,N_3004);
nand U3967 (N_3967,N_3280,N_3394);
or U3968 (N_3968,N_3498,N_3280);
nand U3969 (N_3969,N_3460,N_3247);
nor U3970 (N_3970,N_3388,N_3426);
and U3971 (N_3971,N_3480,N_3182);
nor U3972 (N_3972,N_3430,N_3174);
and U3973 (N_3973,N_3362,N_3269);
and U3974 (N_3974,N_3397,N_3424);
nor U3975 (N_3975,N_3021,N_3099);
nor U3976 (N_3976,N_3216,N_3235);
and U3977 (N_3977,N_3268,N_3269);
nor U3978 (N_3978,N_3008,N_3407);
and U3979 (N_3979,N_3219,N_3387);
and U3980 (N_3980,N_3063,N_3460);
xnor U3981 (N_3981,N_3413,N_3240);
nand U3982 (N_3982,N_3110,N_3300);
xor U3983 (N_3983,N_3196,N_3416);
xnor U3984 (N_3984,N_3253,N_3321);
nor U3985 (N_3985,N_3374,N_3096);
xor U3986 (N_3986,N_3101,N_3139);
xnor U3987 (N_3987,N_3009,N_3195);
and U3988 (N_3988,N_3032,N_3220);
and U3989 (N_3989,N_3133,N_3460);
and U3990 (N_3990,N_3489,N_3147);
xor U3991 (N_3991,N_3424,N_3355);
xnor U3992 (N_3992,N_3112,N_3399);
nand U3993 (N_3993,N_3136,N_3174);
and U3994 (N_3994,N_3362,N_3431);
xor U3995 (N_3995,N_3325,N_3483);
xor U3996 (N_3996,N_3123,N_3481);
or U3997 (N_3997,N_3118,N_3057);
nor U3998 (N_3998,N_3112,N_3369);
nand U3999 (N_3999,N_3005,N_3102);
or U4000 (N_4000,N_3691,N_3582);
and U4001 (N_4001,N_3803,N_3608);
or U4002 (N_4002,N_3556,N_3952);
nand U4003 (N_4003,N_3598,N_3671);
or U4004 (N_4004,N_3868,N_3580);
and U4005 (N_4005,N_3869,N_3754);
nor U4006 (N_4006,N_3966,N_3950);
xor U4007 (N_4007,N_3888,N_3688);
or U4008 (N_4008,N_3786,N_3679);
nor U4009 (N_4009,N_3631,N_3854);
nand U4010 (N_4010,N_3731,N_3719);
or U4011 (N_4011,N_3817,N_3938);
and U4012 (N_4012,N_3625,N_3532);
nor U4013 (N_4013,N_3785,N_3519);
nand U4014 (N_4014,N_3958,N_3725);
nand U4015 (N_4015,N_3630,N_3991);
nor U4016 (N_4016,N_3792,N_3993);
nand U4017 (N_4017,N_3537,N_3695);
and U4018 (N_4018,N_3975,N_3937);
and U4019 (N_4019,N_3827,N_3555);
and U4020 (N_4020,N_3896,N_3920);
nand U4021 (N_4021,N_3621,N_3899);
or U4022 (N_4022,N_3887,N_3825);
and U4023 (N_4023,N_3609,N_3759);
nor U4024 (N_4024,N_3956,N_3901);
or U4025 (N_4025,N_3738,N_3793);
and U4026 (N_4026,N_3806,N_3932);
nand U4027 (N_4027,N_3907,N_3654);
or U4028 (N_4028,N_3961,N_3665);
nand U4029 (N_4029,N_3779,N_3981);
nor U4030 (N_4030,N_3992,N_3940);
nor U4031 (N_4031,N_3984,N_3585);
or U4032 (N_4032,N_3930,N_3667);
and U4033 (N_4033,N_3965,N_3846);
nand U4034 (N_4034,N_3748,N_3894);
xnor U4035 (N_4035,N_3712,N_3505);
xnor U4036 (N_4036,N_3977,N_3925);
or U4037 (N_4037,N_3622,N_3749);
nand U4038 (N_4038,N_3739,N_3575);
and U4039 (N_4039,N_3639,N_3633);
or U4040 (N_4040,N_3919,N_3834);
xor U4041 (N_4041,N_3865,N_3886);
or U4042 (N_4042,N_3670,N_3676);
and U4043 (N_4043,N_3543,N_3685);
nor U4044 (N_4044,N_3566,N_3998);
nor U4045 (N_4045,N_3840,N_3637);
and U4046 (N_4046,N_3509,N_3742);
xnor U4047 (N_4047,N_3948,N_3905);
or U4048 (N_4048,N_3953,N_3851);
or U4049 (N_4049,N_3976,N_3847);
nor U4050 (N_4050,N_3576,N_3507);
xor U4051 (N_4051,N_3546,N_3583);
nor U4052 (N_4052,N_3650,N_3681);
nand U4053 (N_4053,N_3897,N_3772);
nand U4054 (N_4054,N_3577,N_3512);
or U4055 (N_4055,N_3893,N_3799);
or U4056 (N_4056,N_3983,N_3548);
nand U4057 (N_4057,N_3736,N_3636);
nand U4058 (N_4058,N_3955,N_3587);
xor U4059 (N_4059,N_3680,N_3592);
and U4060 (N_4060,N_3570,N_3737);
xnor U4061 (N_4061,N_3658,N_3879);
and U4062 (N_4062,N_3723,N_3524);
and U4063 (N_4063,N_3508,N_3849);
and U4064 (N_4064,N_3878,N_3777);
nor U4065 (N_4065,N_3594,N_3780);
xor U4066 (N_4066,N_3672,N_3623);
nand U4067 (N_4067,N_3941,N_3766);
nand U4068 (N_4068,N_3696,N_3970);
and U4069 (N_4069,N_3588,N_3812);
and U4070 (N_4070,N_3782,N_3673);
and U4071 (N_4071,N_3969,N_3842);
xnor U4072 (N_4072,N_3722,N_3918);
and U4073 (N_4073,N_3765,N_3525);
or U4074 (N_4074,N_3662,N_3890);
xnor U4075 (N_4075,N_3557,N_3960);
nor U4076 (N_4076,N_3820,N_3891);
xor U4077 (N_4077,N_3593,N_3682);
or U4078 (N_4078,N_3789,N_3578);
or U4079 (N_4079,N_3558,N_3657);
and U4080 (N_4080,N_3613,N_3568);
and U4081 (N_4081,N_3763,N_3724);
xor U4082 (N_4082,N_3787,N_3906);
xor U4083 (N_4083,N_3607,N_3503);
xnor U4084 (N_4084,N_3990,N_3808);
xor U4085 (N_4085,N_3721,N_3844);
or U4086 (N_4086,N_3822,N_3559);
nand U4087 (N_4087,N_3752,N_3921);
nand U4088 (N_4088,N_3963,N_3602);
or U4089 (N_4089,N_3776,N_3644);
nand U4090 (N_4090,N_3554,N_3994);
nor U4091 (N_4091,N_3506,N_3610);
or U4092 (N_4092,N_3973,N_3732);
nand U4093 (N_4093,N_3617,N_3616);
nor U4094 (N_4094,N_3746,N_3802);
nand U4095 (N_4095,N_3874,N_3678);
and U4096 (N_4096,N_3515,N_3563);
nor U4097 (N_4097,N_3744,N_3523);
or U4098 (N_4098,N_3596,N_3968);
nand U4099 (N_4099,N_3936,N_3510);
or U4100 (N_4100,N_3804,N_3694);
nand U4101 (N_4101,N_3884,N_3862);
nand U4102 (N_4102,N_3999,N_3767);
xnor U4103 (N_4103,N_3527,N_3861);
nor U4104 (N_4104,N_3801,N_3857);
or U4105 (N_4105,N_3618,N_3597);
nor U4106 (N_4106,N_3705,N_3669);
xor U4107 (N_4107,N_3720,N_3912);
and U4108 (N_4108,N_3653,N_3735);
and U4109 (N_4109,N_3951,N_3611);
nor U4110 (N_4110,N_3795,N_3550);
nand U4111 (N_4111,N_3648,N_3651);
and U4112 (N_4112,N_3915,N_3604);
or U4113 (N_4113,N_3987,N_3771);
nand U4114 (N_4114,N_3917,N_3895);
nor U4115 (N_4115,N_3860,N_3944);
and U4116 (N_4116,N_3675,N_3818);
or U4117 (N_4117,N_3674,N_3743);
nand U4118 (N_4118,N_3699,N_3769);
or U4119 (N_4119,N_3640,N_3781);
and U4120 (N_4120,N_3980,N_3518);
or U4121 (N_4121,N_3707,N_3858);
nor U4122 (N_4122,N_3845,N_3927);
nand U4123 (N_4123,N_3828,N_3957);
nor U4124 (N_4124,N_3996,N_3635);
and U4125 (N_4125,N_3606,N_3706);
nand U4126 (N_4126,N_3520,N_3883);
nand U4127 (N_4127,N_3934,N_3750);
nor U4128 (N_4128,N_3985,N_3626);
or U4129 (N_4129,N_3646,N_3536);
nor U4130 (N_4130,N_3945,N_3656);
xor U4131 (N_4131,N_3659,N_3870);
and U4132 (N_4132,N_3708,N_3796);
or U4133 (N_4133,N_3791,N_3541);
nor U4134 (N_4134,N_3882,N_3881);
nand U4135 (N_4135,N_3762,N_3815);
and U4136 (N_4136,N_3713,N_3764);
nor U4137 (N_4137,N_3848,N_3829);
nor U4138 (N_4138,N_3931,N_3605);
nor U4139 (N_4139,N_3768,N_3761);
and U4140 (N_4140,N_3689,N_3692);
or U4141 (N_4141,N_3502,N_3979);
xor U4142 (N_4142,N_3833,N_3574);
nor U4143 (N_4143,N_3624,N_3995);
nor U4144 (N_4144,N_3783,N_3903);
or U4145 (N_4145,N_3838,N_3726);
nor U4146 (N_4146,N_3521,N_3758);
nor U4147 (N_4147,N_3875,N_3552);
or U4148 (N_4148,N_3734,N_3584);
and U4149 (N_4149,N_3562,N_3939);
nor U4150 (N_4150,N_3733,N_3997);
or U4151 (N_4151,N_3700,N_3704);
xnor U4152 (N_4152,N_3628,N_3811);
and U4153 (N_4153,N_3741,N_3949);
nand U4154 (N_4154,N_3839,N_3821);
and U4155 (N_4155,N_3599,N_3926);
nand U4156 (N_4156,N_3855,N_3740);
nand U4157 (N_4157,N_3770,N_3911);
xor U4158 (N_4158,N_3962,N_3560);
or U4159 (N_4159,N_3549,N_3914);
or U4160 (N_4160,N_3889,N_3972);
xnor U4161 (N_4161,N_3774,N_3661);
nor U4162 (N_4162,N_3876,N_3620);
nand U4163 (N_4163,N_3564,N_3986);
nor U4164 (N_4164,N_3711,N_3843);
nand U4165 (N_4165,N_3864,N_3501);
nand U4166 (N_4166,N_3614,N_3745);
nor U4167 (N_4167,N_3850,N_3747);
or U4168 (N_4168,N_3666,N_3629);
and U4169 (N_4169,N_3978,N_3529);
nor U4170 (N_4170,N_3794,N_3638);
or U4171 (N_4171,N_3810,N_3729);
and U4172 (N_4172,N_3590,N_3800);
nand U4173 (N_4173,N_3909,N_3971);
nor U4174 (N_4174,N_3517,N_3573);
and U4175 (N_4175,N_3756,N_3908);
xor U4176 (N_4176,N_3634,N_3534);
and U4177 (N_4177,N_3863,N_3579);
nor U4178 (N_4178,N_3871,N_3511);
nor U4179 (N_4179,N_3535,N_3819);
and U4180 (N_4180,N_3668,N_3916);
nand U4181 (N_4181,N_3814,N_3540);
nand U4182 (N_4182,N_3683,N_3660);
xor U4183 (N_4183,N_3947,N_3619);
xor U4184 (N_4184,N_3778,N_3885);
nor U4185 (N_4185,N_3526,N_3928);
nand U4186 (N_4186,N_3601,N_3572);
nor U4187 (N_4187,N_3652,N_3728);
or U4188 (N_4188,N_3982,N_3836);
nand U4189 (N_4189,N_3788,N_3933);
and U4190 (N_4190,N_3816,N_3600);
or U4191 (N_4191,N_3504,N_3831);
and U4192 (N_4192,N_3716,N_3935);
or U4193 (N_4193,N_3872,N_3751);
and U4194 (N_4194,N_3841,N_3565);
xnor U4195 (N_4195,N_3797,N_3852);
or U4196 (N_4196,N_3904,N_3589);
xor U4197 (N_4197,N_3547,N_3826);
xor U4198 (N_4198,N_3542,N_3701);
or U4199 (N_4199,N_3798,N_3595);
nor U4200 (N_4200,N_3757,N_3545);
nor U4201 (N_4201,N_3513,N_3530);
or U4202 (N_4202,N_3528,N_3942);
nand U4203 (N_4203,N_3586,N_3727);
xor U4204 (N_4204,N_3643,N_3790);
and U4205 (N_4205,N_3709,N_3824);
or U4206 (N_4206,N_3697,N_3567);
xor U4207 (N_4207,N_3964,N_3551);
or U4208 (N_4208,N_3612,N_3892);
nor U4209 (N_4209,N_3603,N_3553);
and U4210 (N_4210,N_3641,N_3866);
nand U4211 (N_4211,N_3538,N_3853);
xnor U4212 (N_4212,N_3877,N_3898);
xnor U4213 (N_4213,N_3686,N_3663);
xnor U4214 (N_4214,N_3703,N_3561);
or U4215 (N_4215,N_3591,N_3755);
nand U4216 (N_4216,N_3922,N_3946);
and U4217 (N_4217,N_3698,N_3809);
xnor U4218 (N_4218,N_3569,N_3880);
xnor U4219 (N_4219,N_3835,N_3813);
and U4220 (N_4220,N_3760,N_3924);
or U4221 (N_4221,N_3823,N_3544);
xor U4222 (N_4222,N_3859,N_3967);
nor U4223 (N_4223,N_3514,N_3522);
nand U4224 (N_4224,N_3687,N_3581);
and U4225 (N_4225,N_3655,N_3539);
xor U4226 (N_4226,N_3649,N_3710);
nand U4227 (N_4227,N_3805,N_3753);
xor U4228 (N_4228,N_3690,N_3684);
nand U4229 (N_4229,N_3627,N_3988);
nand U4230 (N_4230,N_3773,N_3571);
nor U4231 (N_4231,N_3867,N_3902);
and U4232 (N_4232,N_3873,N_3784);
nand U4233 (N_4233,N_3677,N_3856);
xor U4234 (N_4234,N_3929,N_3832);
and U4235 (N_4235,N_3718,N_3500);
or U4236 (N_4236,N_3954,N_3837);
or U4237 (N_4237,N_3730,N_3632);
xnor U4238 (N_4238,N_3959,N_3900);
nor U4239 (N_4239,N_3775,N_3715);
and U4240 (N_4240,N_3615,N_3647);
and U4241 (N_4241,N_3642,N_3531);
xnor U4242 (N_4242,N_3974,N_3989);
or U4243 (N_4243,N_3533,N_3830);
and U4244 (N_4244,N_3910,N_3645);
and U4245 (N_4245,N_3943,N_3807);
xnor U4246 (N_4246,N_3702,N_3693);
nor U4247 (N_4247,N_3714,N_3923);
and U4248 (N_4248,N_3913,N_3717);
or U4249 (N_4249,N_3664,N_3516);
and U4250 (N_4250,N_3572,N_3585);
or U4251 (N_4251,N_3845,N_3954);
or U4252 (N_4252,N_3981,N_3989);
and U4253 (N_4253,N_3773,N_3712);
or U4254 (N_4254,N_3972,N_3525);
nand U4255 (N_4255,N_3950,N_3989);
or U4256 (N_4256,N_3845,N_3783);
and U4257 (N_4257,N_3663,N_3648);
and U4258 (N_4258,N_3783,N_3643);
nor U4259 (N_4259,N_3952,N_3748);
nand U4260 (N_4260,N_3796,N_3638);
and U4261 (N_4261,N_3651,N_3587);
xor U4262 (N_4262,N_3674,N_3666);
and U4263 (N_4263,N_3892,N_3964);
or U4264 (N_4264,N_3645,N_3665);
nor U4265 (N_4265,N_3796,N_3872);
xnor U4266 (N_4266,N_3809,N_3895);
xor U4267 (N_4267,N_3692,N_3810);
nand U4268 (N_4268,N_3686,N_3524);
or U4269 (N_4269,N_3826,N_3843);
nor U4270 (N_4270,N_3584,N_3788);
or U4271 (N_4271,N_3923,N_3730);
or U4272 (N_4272,N_3589,N_3677);
and U4273 (N_4273,N_3851,N_3793);
and U4274 (N_4274,N_3683,N_3757);
nor U4275 (N_4275,N_3583,N_3570);
and U4276 (N_4276,N_3635,N_3709);
xnor U4277 (N_4277,N_3570,N_3999);
nand U4278 (N_4278,N_3943,N_3751);
or U4279 (N_4279,N_3742,N_3682);
nand U4280 (N_4280,N_3788,N_3913);
nor U4281 (N_4281,N_3862,N_3850);
and U4282 (N_4282,N_3950,N_3568);
nor U4283 (N_4283,N_3915,N_3738);
nand U4284 (N_4284,N_3962,N_3670);
and U4285 (N_4285,N_3603,N_3988);
nor U4286 (N_4286,N_3524,N_3777);
and U4287 (N_4287,N_3999,N_3713);
xor U4288 (N_4288,N_3983,N_3945);
xnor U4289 (N_4289,N_3581,N_3772);
or U4290 (N_4290,N_3654,N_3909);
xnor U4291 (N_4291,N_3715,N_3913);
and U4292 (N_4292,N_3665,N_3764);
xor U4293 (N_4293,N_3772,N_3987);
nor U4294 (N_4294,N_3907,N_3770);
and U4295 (N_4295,N_3931,N_3960);
or U4296 (N_4296,N_3635,N_3827);
xnor U4297 (N_4297,N_3847,N_3791);
and U4298 (N_4298,N_3707,N_3559);
xnor U4299 (N_4299,N_3613,N_3631);
nor U4300 (N_4300,N_3993,N_3893);
and U4301 (N_4301,N_3994,N_3962);
and U4302 (N_4302,N_3725,N_3662);
or U4303 (N_4303,N_3967,N_3518);
nor U4304 (N_4304,N_3852,N_3617);
nand U4305 (N_4305,N_3525,N_3539);
or U4306 (N_4306,N_3802,N_3981);
nand U4307 (N_4307,N_3772,N_3965);
nor U4308 (N_4308,N_3986,N_3967);
or U4309 (N_4309,N_3853,N_3565);
nand U4310 (N_4310,N_3659,N_3586);
nor U4311 (N_4311,N_3876,N_3564);
or U4312 (N_4312,N_3940,N_3697);
nor U4313 (N_4313,N_3592,N_3617);
nand U4314 (N_4314,N_3946,N_3834);
xor U4315 (N_4315,N_3701,N_3891);
nand U4316 (N_4316,N_3542,N_3761);
and U4317 (N_4317,N_3685,N_3861);
and U4318 (N_4318,N_3958,N_3674);
and U4319 (N_4319,N_3558,N_3633);
nor U4320 (N_4320,N_3695,N_3637);
and U4321 (N_4321,N_3920,N_3742);
or U4322 (N_4322,N_3598,N_3712);
xor U4323 (N_4323,N_3762,N_3970);
or U4324 (N_4324,N_3615,N_3838);
nand U4325 (N_4325,N_3688,N_3527);
or U4326 (N_4326,N_3550,N_3704);
nor U4327 (N_4327,N_3892,N_3513);
or U4328 (N_4328,N_3586,N_3764);
or U4329 (N_4329,N_3919,N_3810);
or U4330 (N_4330,N_3575,N_3660);
xor U4331 (N_4331,N_3965,N_3538);
nor U4332 (N_4332,N_3890,N_3976);
nand U4333 (N_4333,N_3716,N_3560);
xnor U4334 (N_4334,N_3709,N_3837);
xor U4335 (N_4335,N_3881,N_3870);
xnor U4336 (N_4336,N_3755,N_3673);
xnor U4337 (N_4337,N_3939,N_3532);
nor U4338 (N_4338,N_3805,N_3802);
and U4339 (N_4339,N_3607,N_3765);
nor U4340 (N_4340,N_3631,N_3795);
and U4341 (N_4341,N_3671,N_3911);
or U4342 (N_4342,N_3856,N_3662);
nand U4343 (N_4343,N_3816,N_3758);
xor U4344 (N_4344,N_3847,N_3636);
xor U4345 (N_4345,N_3905,N_3529);
nand U4346 (N_4346,N_3638,N_3918);
nor U4347 (N_4347,N_3760,N_3513);
nand U4348 (N_4348,N_3764,N_3601);
nand U4349 (N_4349,N_3601,N_3829);
nand U4350 (N_4350,N_3775,N_3661);
or U4351 (N_4351,N_3517,N_3800);
nor U4352 (N_4352,N_3610,N_3846);
and U4353 (N_4353,N_3545,N_3509);
nor U4354 (N_4354,N_3558,N_3883);
or U4355 (N_4355,N_3648,N_3790);
and U4356 (N_4356,N_3858,N_3525);
or U4357 (N_4357,N_3506,N_3790);
xnor U4358 (N_4358,N_3863,N_3908);
or U4359 (N_4359,N_3968,N_3899);
or U4360 (N_4360,N_3939,N_3992);
nor U4361 (N_4361,N_3723,N_3739);
xor U4362 (N_4362,N_3575,N_3868);
nand U4363 (N_4363,N_3906,N_3984);
nor U4364 (N_4364,N_3683,N_3978);
nand U4365 (N_4365,N_3524,N_3914);
nand U4366 (N_4366,N_3834,N_3775);
xnor U4367 (N_4367,N_3989,N_3632);
nand U4368 (N_4368,N_3881,N_3641);
nand U4369 (N_4369,N_3837,N_3633);
nor U4370 (N_4370,N_3756,N_3916);
nor U4371 (N_4371,N_3862,N_3688);
nand U4372 (N_4372,N_3945,N_3588);
nor U4373 (N_4373,N_3592,N_3557);
or U4374 (N_4374,N_3898,N_3901);
nor U4375 (N_4375,N_3675,N_3848);
xor U4376 (N_4376,N_3867,N_3868);
and U4377 (N_4377,N_3824,N_3888);
nand U4378 (N_4378,N_3786,N_3790);
and U4379 (N_4379,N_3782,N_3803);
and U4380 (N_4380,N_3533,N_3678);
xor U4381 (N_4381,N_3641,N_3985);
or U4382 (N_4382,N_3771,N_3866);
xor U4383 (N_4383,N_3760,N_3686);
nand U4384 (N_4384,N_3997,N_3914);
xor U4385 (N_4385,N_3777,N_3728);
or U4386 (N_4386,N_3848,N_3564);
nand U4387 (N_4387,N_3922,N_3843);
nor U4388 (N_4388,N_3956,N_3715);
nand U4389 (N_4389,N_3586,N_3899);
and U4390 (N_4390,N_3962,N_3744);
nand U4391 (N_4391,N_3993,N_3850);
xnor U4392 (N_4392,N_3624,N_3947);
or U4393 (N_4393,N_3705,N_3624);
nand U4394 (N_4394,N_3792,N_3748);
nor U4395 (N_4395,N_3763,N_3953);
or U4396 (N_4396,N_3597,N_3952);
and U4397 (N_4397,N_3952,N_3879);
nand U4398 (N_4398,N_3655,N_3825);
xnor U4399 (N_4399,N_3514,N_3985);
nand U4400 (N_4400,N_3507,N_3897);
or U4401 (N_4401,N_3829,N_3666);
nand U4402 (N_4402,N_3816,N_3779);
nand U4403 (N_4403,N_3777,N_3991);
nor U4404 (N_4404,N_3657,N_3721);
nand U4405 (N_4405,N_3580,N_3975);
xnor U4406 (N_4406,N_3573,N_3732);
nand U4407 (N_4407,N_3739,N_3832);
nand U4408 (N_4408,N_3609,N_3541);
xor U4409 (N_4409,N_3523,N_3897);
xor U4410 (N_4410,N_3804,N_3638);
or U4411 (N_4411,N_3813,N_3580);
nand U4412 (N_4412,N_3614,N_3775);
nor U4413 (N_4413,N_3647,N_3560);
nand U4414 (N_4414,N_3570,N_3912);
and U4415 (N_4415,N_3707,N_3878);
and U4416 (N_4416,N_3659,N_3934);
nor U4417 (N_4417,N_3551,N_3815);
nand U4418 (N_4418,N_3592,N_3645);
and U4419 (N_4419,N_3883,N_3976);
or U4420 (N_4420,N_3817,N_3875);
nand U4421 (N_4421,N_3901,N_3561);
xor U4422 (N_4422,N_3999,N_3703);
nor U4423 (N_4423,N_3817,N_3837);
xnor U4424 (N_4424,N_3522,N_3580);
or U4425 (N_4425,N_3908,N_3889);
and U4426 (N_4426,N_3814,N_3624);
nand U4427 (N_4427,N_3995,N_3686);
or U4428 (N_4428,N_3536,N_3990);
nand U4429 (N_4429,N_3704,N_3625);
and U4430 (N_4430,N_3949,N_3599);
nand U4431 (N_4431,N_3824,N_3775);
or U4432 (N_4432,N_3509,N_3692);
nor U4433 (N_4433,N_3980,N_3947);
or U4434 (N_4434,N_3893,N_3815);
xor U4435 (N_4435,N_3676,N_3600);
and U4436 (N_4436,N_3812,N_3633);
xor U4437 (N_4437,N_3833,N_3608);
xor U4438 (N_4438,N_3853,N_3705);
and U4439 (N_4439,N_3634,N_3632);
xor U4440 (N_4440,N_3922,N_3517);
nand U4441 (N_4441,N_3994,N_3869);
nor U4442 (N_4442,N_3812,N_3831);
or U4443 (N_4443,N_3714,N_3943);
or U4444 (N_4444,N_3972,N_3683);
or U4445 (N_4445,N_3811,N_3887);
nand U4446 (N_4446,N_3717,N_3994);
and U4447 (N_4447,N_3689,N_3591);
and U4448 (N_4448,N_3880,N_3721);
nor U4449 (N_4449,N_3818,N_3951);
nand U4450 (N_4450,N_3687,N_3648);
and U4451 (N_4451,N_3924,N_3912);
and U4452 (N_4452,N_3548,N_3861);
or U4453 (N_4453,N_3961,N_3901);
nor U4454 (N_4454,N_3588,N_3690);
or U4455 (N_4455,N_3802,N_3983);
nor U4456 (N_4456,N_3563,N_3633);
or U4457 (N_4457,N_3526,N_3680);
xor U4458 (N_4458,N_3758,N_3988);
xor U4459 (N_4459,N_3566,N_3673);
and U4460 (N_4460,N_3786,N_3707);
xor U4461 (N_4461,N_3584,N_3505);
or U4462 (N_4462,N_3900,N_3655);
xnor U4463 (N_4463,N_3586,N_3724);
nor U4464 (N_4464,N_3568,N_3881);
and U4465 (N_4465,N_3987,N_3548);
nor U4466 (N_4466,N_3840,N_3721);
nor U4467 (N_4467,N_3966,N_3997);
xnor U4468 (N_4468,N_3578,N_3701);
xor U4469 (N_4469,N_3795,N_3927);
nor U4470 (N_4470,N_3927,N_3637);
and U4471 (N_4471,N_3886,N_3717);
xor U4472 (N_4472,N_3794,N_3624);
and U4473 (N_4473,N_3614,N_3582);
nor U4474 (N_4474,N_3761,N_3854);
and U4475 (N_4475,N_3656,N_3779);
xor U4476 (N_4476,N_3922,N_3739);
nand U4477 (N_4477,N_3634,N_3527);
nor U4478 (N_4478,N_3834,N_3635);
or U4479 (N_4479,N_3831,N_3745);
nor U4480 (N_4480,N_3706,N_3902);
and U4481 (N_4481,N_3627,N_3825);
nor U4482 (N_4482,N_3840,N_3752);
nor U4483 (N_4483,N_3832,N_3915);
or U4484 (N_4484,N_3720,N_3641);
nand U4485 (N_4485,N_3748,N_3879);
or U4486 (N_4486,N_3790,N_3538);
and U4487 (N_4487,N_3615,N_3919);
or U4488 (N_4488,N_3639,N_3519);
and U4489 (N_4489,N_3802,N_3756);
and U4490 (N_4490,N_3756,N_3544);
or U4491 (N_4491,N_3540,N_3738);
and U4492 (N_4492,N_3888,N_3933);
xnor U4493 (N_4493,N_3613,N_3676);
or U4494 (N_4494,N_3874,N_3563);
or U4495 (N_4495,N_3889,N_3840);
xnor U4496 (N_4496,N_3817,N_3714);
and U4497 (N_4497,N_3570,N_3586);
nor U4498 (N_4498,N_3539,N_3585);
or U4499 (N_4499,N_3691,N_3926);
and U4500 (N_4500,N_4307,N_4091);
or U4501 (N_4501,N_4042,N_4048);
and U4502 (N_4502,N_4184,N_4209);
and U4503 (N_4503,N_4479,N_4336);
or U4504 (N_4504,N_4190,N_4341);
or U4505 (N_4505,N_4276,N_4296);
nand U4506 (N_4506,N_4470,N_4034);
or U4507 (N_4507,N_4331,N_4410);
nor U4508 (N_4508,N_4208,N_4004);
nand U4509 (N_4509,N_4013,N_4137);
xor U4510 (N_4510,N_4468,N_4449);
nand U4511 (N_4511,N_4061,N_4332);
nand U4512 (N_4512,N_4471,N_4085);
nand U4513 (N_4513,N_4437,N_4128);
nand U4514 (N_4514,N_4459,N_4023);
and U4515 (N_4515,N_4441,N_4130);
nand U4516 (N_4516,N_4419,N_4363);
xnor U4517 (N_4517,N_4308,N_4068);
nor U4518 (N_4518,N_4025,N_4466);
xor U4519 (N_4519,N_4492,N_4411);
nand U4520 (N_4520,N_4159,N_4440);
or U4521 (N_4521,N_4149,N_4260);
xnor U4522 (N_4522,N_4206,N_4291);
nor U4523 (N_4523,N_4392,N_4300);
or U4524 (N_4524,N_4325,N_4305);
nor U4525 (N_4525,N_4142,N_4063);
or U4526 (N_4526,N_4314,N_4233);
xor U4527 (N_4527,N_4046,N_4187);
nor U4528 (N_4528,N_4253,N_4380);
nand U4529 (N_4529,N_4255,N_4108);
nor U4530 (N_4530,N_4098,N_4350);
nor U4531 (N_4531,N_4258,N_4216);
nand U4532 (N_4532,N_4489,N_4249);
xnor U4533 (N_4533,N_4207,N_4328);
nand U4534 (N_4534,N_4185,N_4121);
nand U4535 (N_4535,N_4175,N_4056);
or U4536 (N_4536,N_4480,N_4227);
nor U4537 (N_4537,N_4272,N_4084);
or U4538 (N_4538,N_4431,N_4181);
or U4539 (N_4539,N_4111,N_4211);
xnor U4540 (N_4540,N_4408,N_4490);
xnor U4541 (N_4541,N_4297,N_4204);
nor U4542 (N_4542,N_4228,N_4484);
nor U4543 (N_4543,N_4434,N_4106);
nor U4544 (N_4544,N_4226,N_4167);
nand U4545 (N_4545,N_4372,N_4021);
nand U4546 (N_4546,N_4497,N_4095);
xor U4547 (N_4547,N_4442,N_4409);
nand U4548 (N_4548,N_4451,N_4357);
nor U4549 (N_4549,N_4349,N_4165);
or U4550 (N_4550,N_4005,N_4265);
and U4551 (N_4551,N_4244,N_4127);
xnor U4552 (N_4552,N_4330,N_4213);
xor U4553 (N_4553,N_4032,N_4317);
xor U4554 (N_4554,N_4065,N_4112);
nor U4555 (N_4555,N_4231,N_4214);
xor U4556 (N_4556,N_4456,N_4358);
and U4557 (N_4557,N_4155,N_4124);
xnor U4558 (N_4558,N_4424,N_4163);
and U4559 (N_4559,N_4453,N_4039);
and U4560 (N_4560,N_4284,N_4270);
or U4561 (N_4561,N_4309,N_4279);
nor U4562 (N_4562,N_4205,N_4047);
xor U4563 (N_4563,N_4457,N_4476);
and U4564 (N_4564,N_4026,N_4014);
or U4565 (N_4565,N_4282,N_4413);
and U4566 (N_4566,N_4134,N_4290);
nand U4567 (N_4567,N_4403,N_4221);
nor U4568 (N_4568,N_4340,N_4261);
or U4569 (N_4569,N_4323,N_4469);
or U4570 (N_4570,N_4082,N_4200);
nor U4571 (N_4571,N_4103,N_4031);
and U4572 (N_4572,N_4289,N_4060);
xor U4573 (N_4573,N_4009,N_4241);
nand U4574 (N_4574,N_4493,N_4474);
nand U4575 (N_4575,N_4024,N_4237);
and U4576 (N_4576,N_4377,N_4368);
nand U4577 (N_4577,N_4080,N_4388);
and U4578 (N_4578,N_4355,N_4102);
nor U4579 (N_4579,N_4460,N_4417);
or U4580 (N_4580,N_4280,N_4045);
or U4581 (N_4581,N_4180,N_4389);
and U4582 (N_4582,N_4071,N_4016);
nor U4583 (N_4583,N_4361,N_4105);
nor U4584 (N_4584,N_4110,N_4438);
nor U4585 (N_4585,N_4275,N_4346);
nor U4586 (N_4586,N_4375,N_4138);
nand U4587 (N_4587,N_4343,N_4230);
nor U4588 (N_4588,N_4088,N_4294);
nand U4589 (N_4589,N_4057,N_4172);
nor U4590 (N_4590,N_4354,N_4051);
or U4591 (N_4591,N_4401,N_4433);
or U4592 (N_4592,N_4381,N_4311);
or U4593 (N_4593,N_4306,N_4269);
xor U4594 (N_4594,N_4464,N_4139);
nor U4595 (N_4595,N_4263,N_4423);
nand U4596 (N_4596,N_4104,N_4010);
nor U4597 (N_4597,N_4268,N_4076);
xor U4598 (N_4598,N_4271,N_4083);
xnor U4599 (N_4599,N_4292,N_4310);
and U4600 (N_4600,N_4369,N_4416);
nand U4601 (N_4601,N_4498,N_4015);
or U4602 (N_4602,N_4406,N_4096);
nor U4603 (N_4603,N_4176,N_4259);
nor U4604 (N_4604,N_4006,N_4179);
nand U4605 (N_4605,N_4298,N_4073);
xor U4606 (N_4606,N_4017,N_4146);
nor U4607 (N_4607,N_4089,N_4362);
xnor U4608 (N_4608,N_4435,N_4475);
nor U4609 (N_4609,N_4000,N_4444);
nand U4610 (N_4610,N_4277,N_4266);
and U4611 (N_4611,N_4193,N_4174);
xor U4612 (N_4612,N_4356,N_4397);
nor U4613 (N_4613,N_4191,N_4278);
or U4614 (N_4614,N_4001,N_4011);
nor U4615 (N_4615,N_4118,N_4147);
or U4616 (N_4616,N_4069,N_4201);
xor U4617 (N_4617,N_4114,N_4171);
xnor U4618 (N_4618,N_4251,N_4168);
xnor U4619 (N_4619,N_4315,N_4186);
nor U4620 (N_4620,N_4339,N_4232);
xnor U4621 (N_4621,N_4151,N_4148);
nand U4622 (N_4622,N_4443,N_4288);
nor U4623 (N_4623,N_4412,N_4030);
and U4624 (N_4624,N_4432,N_4132);
and U4625 (N_4625,N_4342,N_4100);
nor U4626 (N_4626,N_4383,N_4324);
and U4627 (N_4627,N_4422,N_4072);
or U4628 (N_4628,N_4123,N_4020);
xnor U4629 (N_4629,N_4087,N_4295);
xor U4630 (N_4630,N_4119,N_4491);
or U4631 (N_4631,N_4229,N_4360);
xnor U4632 (N_4632,N_4224,N_4386);
and U4633 (N_4633,N_4283,N_4164);
xnor U4634 (N_4634,N_4420,N_4402);
or U4635 (N_4635,N_4371,N_4390);
nand U4636 (N_4636,N_4486,N_4160);
nand U4637 (N_4637,N_4055,N_4002);
or U4638 (N_4638,N_4304,N_4379);
nand U4639 (N_4639,N_4188,N_4079);
nor U4640 (N_4640,N_4094,N_4238);
and U4641 (N_4641,N_4086,N_4302);
and U4642 (N_4642,N_4344,N_4418);
and U4643 (N_4643,N_4036,N_4029);
xor U4644 (N_4644,N_4140,N_4252);
or U4645 (N_4645,N_4326,N_4463);
nand U4646 (N_4646,N_4445,N_4143);
nor U4647 (N_4647,N_4334,N_4235);
or U4648 (N_4648,N_4236,N_4487);
nand U4649 (N_4649,N_4043,N_4131);
xnor U4650 (N_4650,N_4202,N_4178);
nand U4651 (N_4651,N_4387,N_4478);
or U4652 (N_4652,N_4246,N_4250);
and U4653 (N_4653,N_4092,N_4152);
nor U4654 (N_4654,N_4393,N_4059);
xor U4655 (N_4655,N_4367,N_4345);
xnor U4656 (N_4656,N_4382,N_4448);
and U4657 (N_4657,N_4194,N_4173);
nor U4658 (N_4658,N_4287,N_4447);
nor U4659 (N_4659,N_4376,N_4012);
xnor U4660 (N_4660,N_4414,N_4038);
nand U4661 (N_4661,N_4396,N_4153);
nand U4662 (N_4662,N_4049,N_4462);
and U4663 (N_4663,N_4273,N_4415);
nand U4664 (N_4664,N_4220,N_4243);
or U4665 (N_4665,N_4019,N_4197);
nor U4666 (N_4666,N_4133,N_4482);
and U4667 (N_4667,N_4477,N_4135);
xnor U4668 (N_4668,N_4141,N_4481);
and U4669 (N_4669,N_4223,N_4018);
xnor U4670 (N_4670,N_4054,N_4041);
and U4671 (N_4671,N_4008,N_4301);
xor U4672 (N_4672,N_4099,N_4192);
and U4673 (N_4673,N_4274,N_4081);
nor U4674 (N_4674,N_4198,N_4439);
nand U4675 (N_4675,N_4312,N_4007);
and U4676 (N_4676,N_4117,N_4101);
or U4677 (N_4677,N_4407,N_4078);
nor U4678 (N_4678,N_4113,N_4318);
xnor U4679 (N_4679,N_4066,N_4428);
nand U4680 (N_4680,N_4446,N_4264);
and U4681 (N_4681,N_4203,N_4267);
nand U4682 (N_4682,N_4116,N_4157);
or U4683 (N_4683,N_4210,N_4240);
or U4684 (N_4684,N_4070,N_4347);
or U4685 (N_4685,N_4254,N_4337);
nor U4686 (N_4686,N_4215,N_4450);
nor U4687 (N_4687,N_4373,N_4234);
nand U4688 (N_4688,N_4385,N_4027);
nand U4689 (N_4689,N_4483,N_4090);
or U4690 (N_4690,N_4351,N_4496);
nor U4691 (N_4691,N_4189,N_4495);
and U4692 (N_4692,N_4281,N_4370);
nor U4693 (N_4693,N_4129,N_4458);
or U4694 (N_4694,N_4256,N_4322);
and U4695 (N_4695,N_4405,N_4126);
or U4696 (N_4696,N_4212,N_4473);
nand U4697 (N_4697,N_4299,N_4109);
and U4698 (N_4698,N_4144,N_4257);
or U4699 (N_4699,N_4391,N_4286);
nand U4700 (N_4700,N_4313,N_4404);
or U4701 (N_4701,N_4075,N_4161);
or U4702 (N_4702,N_4052,N_4040);
xnor U4703 (N_4703,N_4427,N_4120);
xnor U4704 (N_4704,N_4394,N_4378);
nor U4705 (N_4705,N_4320,N_4150);
nor U4706 (N_4706,N_4293,N_4425);
or U4707 (N_4707,N_4365,N_4053);
nand U4708 (N_4708,N_4097,N_4158);
xnor U4709 (N_4709,N_4316,N_4199);
nand U4710 (N_4710,N_4122,N_4454);
or U4711 (N_4711,N_4429,N_4064);
or U4712 (N_4712,N_4400,N_4145);
or U4713 (N_4713,N_4050,N_4125);
or U4714 (N_4714,N_4177,N_4366);
and U4715 (N_4715,N_4154,N_4384);
and U4716 (N_4716,N_4395,N_4303);
and U4717 (N_4717,N_4219,N_4222);
and U4718 (N_4718,N_4033,N_4472);
nor U4719 (N_4719,N_4003,N_4499);
xor U4720 (N_4720,N_4058,N_4035);
and U4721 (N_4721,N_4022,N_4426);
or U4722 (N_4722,N_4115,N_4430);
xor U4723 (N_4723,N_4353,N_4170);
nand U4724 (N_4724,N_4248,N_4028);
or U4725 (N_4725,N_4352,N_4327);
or U4726 (N_4726,N_4245,N_4319);
nor U4727 (N_4727,N_4093,N_4399);
nor U4728 (N_4728,N_4166,N_4348);
nand U4729 (N_4729,N_4077,N_4461);
nor U4730 (N_4730,N_4374,N_4338);
or U4731 (N_4731,N_4455,N_4044);
or U4732 (N_4732,N_4037,N_4107);
xnor U4733 (N_4733,N_4182,N_4335);
and U4734 (N_4734,N_4218,N_4239);
nor U4735 (N_4735,N_4452,N_4162);
or U4736 (N_4736,N_4074,N_4329);
and U4737 (N_4737,N_4333,N_4247);
nand U4738 (N_4738,N_4067,N_4398);
and U4739 (N_4739,N_4136,N_4364);
xor U4740 (N_4740,N_4195,N_4285);
nor U4741 (N_4741,N_4062,N_4436);
nor U4742 (N_4742,N_4156,N_4421);
and U4743 (N_4743,N_4488,N_4262);
and U4744 (N_4744,N_4321,N_4467);
nor U4745 (N_4745,N_4359,N_4494);
nor U4746 (N_4746,N_4217,N_4485);
and U4747 (N_4747,N_4465,N_4183);
nor U4748 (N_4748,N_4225,N_4242);
nor U4749 (N_4749,N_4169,N_4196);
xnor U4750 (N_4750,N_4441,N_4131);
nand U4751 (N_4751,N_4110,N_4351);
nand U4752 (N_4752,N_4239,N_4039);
and U4753 (N_4753,N_4325,N_4120);
or U4754 (N_4754,N_4188,N_4322);
and U4755 (N_4755,N_4397,N_4313);
xnor U4756 (N_4756,N_4224,N_4473);
xnor U4757 (N_4757,N_4111,N_4221);
and U4758 (N_4758,N_4231,N_4198);
and U4759 (N_4759,N_4051,N_4140);
or U4760 (N_4760,N_4373,N_4238);
xor U4761 (N_4761,N_4410,N_4374);
nand U4762 (N_4762,N_4367,N_4497);
nor U4763 (N_4763,N_4486,N_4480);
nand U4764 (N_4764,N_4448,N_4014);
or U4765 (N_4765,N_4227,N_4094);
or U4766 (N_4766,N_4281,N_4322);
nand U4767 (N_4767,N_4042,N_4311);
nand U4768 (N_4768,N_4436,N_4014);
xnor U4769 (N_4769,N_4189,N_4185);
or U4770 (N_4770,N_4114,N_4101);
xnor U4771 (N_4771,N_4402,N_4366);
or U4772 (N_4772,N_4121,N_4284);
nand U4773 (N_4773,N_4414,N_4189);
nor U4774 (N_4774,N_4021,N_4441);
and U4775 (N_4775,N_4153,N_4156);
nand U4776 (N_4776,N_4100,N_4289);
and U4777 (N_4777,N_4315,N_4308);
xnor U4778 (N_4778,N_4038,N_4150);
xor U4779 (N_4779,N_4169,N_4401);
nor U4780 (N_4780,N_4402,N_4105);
xnor U4781 (N_4781,N_4176,N_4227);
and U4782 (N_4782,N_4140,N_4058);
nand U4783 (N_4783,N_4058,N_4301);
xor U4784 (N_4784,N_4474,N_4119);
xnor U4785 (N_4785,N_4432,N_4044);
nor U4786 (N_4786,N_4099,N_4437);
and U4787 (N_4787,N_4067,N_4114);
or U4788 (N_4788,N_4351,N_4024);
or U4789 (N_4789,N_4187,N_4372);
or U4790 (N_4790,N_4060,N_4098);
and U4791 (N_4791,N_4151,N_4060);
and U4792 (N_4792,N_4160,N_4149);
nor U4793 (N_4793,N_4304,N_4001);
and U4794 (N_4794,N_4065,N_4270);
or U4795 (N_4795,N_4086,N_4207);
nor U4796 (N_4796,N_4034,N_4142);
or U4797 (N_4797,N_4045,N_4219);
or U4798 (N_4798,N_4313,N_4387);
xnor U4799 (N_4799,N_4493,N_4023);
nand U4800 (N_4800,N_4167,N_4093);
xnor U4801 (N_4801,N_4368,N_4465);
nand U4802 (N_4802,N_4402,N_4475);
and U4803 (N_4803,N_4148,N_4361);
and U4804 (N_4804,N_4480,N_4137);
nor U4805 (N_4805,N_4360,N_4396);
xor U4806 (N_4806,N_4218,N_4458);
or U4807 (N_4807,N_4151,N_4395);
nor U4808 (N_4808,N_4121,N_4231);
or U4809 (N_4809,N_4460,N_4293);
nor U4810 (N_4810,N_4028,N_4295);
nand U4811 (N_4811,N_4043,N_4482);
nor U4812 (N_4812,N_4032,N_4143);
nand U4813 (N_4813,N_4003,N_4273);
nand U4814 (N_4814,N_4429,N_4111);
nor U4815 (N_4815,N_4027,N_4007);
or U4816 (N_4816,N_4172,N_4279);
and U4817 (N_4817,N_4062,N_4479);
xnor U4818 (N_4818,N_4392,N_4255);
and U4819 (N_4819,N_4165,N_4352);
and U4820 (N_4820,N_4019,N_4214);
nand U4821 (N_4821,N_4397,N_4296);
xor U4822 (N_4822,N_4456,N_4173);
xor U4823 (N_4823,N_4309,N_4012);
nor U4824 (N_4824,N_4210,N_4074);
and U4825 (N_4825,N_4337,N_4371);
and U4826 (N_4826,N_4155,N_4446);
or U4827 (N_4827,N_4097,N_4340);
nor U4828 (N_4828,N_4445,N_4105);
nand U4829 (N_4829,N_4099,N_4244);
nor U4830 (N_4830,N_4198,N_4262);
or U4831 (N_4831,N_4201,N_4453);
nand U4832 (N_4832,N_4336,N_4195);
or U4833 (N_4833,N_4252,N_4112);
nor U4834 (N_4834,N_4347,N_4374);
xor U4835 (N_4835,N_4278,N_4447);
and U4836 (N_4836,N_4175,N_4418);
nand U4837 (N_4837,N_4441,N_4399);
nor U4838 (N_4838,N_4129,N_4427);
nand U4839 (N_4839,N_4464,N_4336);
or U4840 (N_4840,N_4079,N_4243);
xnor U4841 (N_4841,N_4339,N_4494);
nand U4842 (N_4842,N_4480,N_4278);
and U4843 (N_4843,N_4288,N_4034);
nor U4844 (N_4844,N_4180,N_4186);
or U4845 (N_4845,N_4337,N_4451);
nand U4846 (N_4846,N_4139,N_4387);
nor U4847 (N_4847,N_4426,N_4344);
or U4848 (N_4848,N_4427,N_4345);
nor U4849 (N_4849,N_4281,N_4331);
and U4850 (N_4850,N_4493,N_4236);
or U4851 (N_4851,N_4125,N_4173);
nor U4852 (N_4852,N_4162,N_4473);
xor U4853 (N_4853,N_4060,N_4376);
nor U4854 (N_4854,N_4409,N_4300);
nand U4855 (N_4855,N_4470,N_4413);
and U4856 (N_4856,N_4334,N_4088);
and U4857 (N_4857,N_4297,N_4458);
nand U4858 (N_4858,N_4008,N_4365);
and U4859 (N_4859,N_4407,N_4310);
nor U4860 (N_4860,N_4194,N_4093);
xnor U4861 (N_4861,N_4379,N_4326);
xor U4862 (N_4862,N_4492,N_4065);
nor U4863 (N_4863,N_4116,N_4192);
nand U4864 (N_4864,N_4031,N_4209);
nand U4865 (N_4865,N_4420,N_4140);
or U4866 (N_4866,N_4050,N_4305);
xor U4867 (N_4867,N_4354,N_4277);
or U4868 (N_4868,N_4343,N_4124);
or U4869 (N_4869,N_4141,N_4166);
xnor U4870 (N_4870,N_4367,N_4205);
xor U4871 (N_4871,N_4271,N_4049);
nand U4872 (N_4872,N_4181,N_4264);
nand U4873 (N_4873,N_4098,N_4033);
and U4874 (N_4874,N_4425,N_4165);
nand U4875 (N_4875,N_4199,N_4463);
xor U4876 (N_4876,N_4279,N_4196);
and U4877 (N_4877,N_4403,N_4103);
nand U4878 (N_4878,N_4385,N_4404);
nand U4879 (N_4879,N_4427,N_4177);
or U4880 (N_4880,N_4439,N_4116);
nor U4881 (N_4881,N_4385,N_4172);
nand U4882 (N_4882,N_4147,N_4172);
nor U4883 (N_4883,N_4370,N_4240);
nor U4884 (N_4884,N_4059,N_4282);
xnor U4885 (N_4885,N_4382,N_4162);
xor U4886 (N_4886,N_4443,N_4333);
and U4887 (N_4887,N_4477,N_4456);
xnor U4888 (N_4888,N_4263,N_4112);
nand U4889 (N_4889,N_4497,N_4051);
nand U4890 (N_4890,N_4206,N_4366);
and U4891 (N_4891,N_4174,N_4018);
nor U4892 (N_4892,N_4341,N_4160);
xor U4893 (N_4893,N_4072,N_4252);
and U4894 (N_4894,N_4413,N_4280);
or U4895 (N_4895,N_4398,N_4428);
nand U4896 (N_4896,N_4473,N_4167);
nor U4897 (N_4897,N_4208,N_4118);
or U4898 (N_4898,N_4384,N_4115);
or U4899 (N_4899,N_4213,N_4000);
and U4900 (N_4900,N_4454,N_4123);
nand U4901 (N_4901,N_4136,N_4237);
nand U4902 (N_4902,N_4381,N_4461);
nand U4903 (N_4903,N_4444,N_4099);
nand U4904 (N_4904,N_4361,N_4415);
and U4905 (N_4905,N_4022,N_4068);
or U4906 (N_4906,N_4109,N_4410);
or U4907 (N_4907,N_4112,N_4336);
and U4908 (N_4908,N_4383,N_4086);
nor U4909 (N_4909,N_4273,N_4203);
xnor U4910 (N_4910,N_4045,N_4036);
or U4911 (N_4911,N_4343,N_4175);
and U4912 (N_4912,N_4246,N_4230);
or U4913 (N_4913,N_4027,N_4079);
xor U4914 (N_4914,N_4129,N_4044);
or U4915 (N_4915,N_4052,N_4393);
nor U4916 (N_4916,N_4058,N_4323);
xnor U4917 (N_4917,N_4080,N_4344);
nand U4918 (N_4918,N_4210,N_4078);
xnor U4919 (N_4919,N_4059,N_4279);
xnor U4920 (N_4920,N_4331,N_4158);
nand U4921 (N_4921,N_4128,N_4216);
nor U4922 (N_4922,N_4084,N_4306);
xor U4923 (N_4923,N_4320,N_4109);
nor U4924 (N_4924,N_4138,N_4221);
or U4925 (N_4925,N_4148,N_4214);
and U4926 (N_4926,N_4143,N_4487);
nand U4927 (N_4927,N_4072,N_4028);
and U4928 (N_4928,N_4441,N_4341);
or U4929 (N_4929,N_4211,N_4499);
or U4930 (N_4930,N_4370,N_4253);
and U4931 (N_4931,N_4234,N_4393);
nor U4932 (N_4932,N_4279,N_4092);
or U4933 (N_4933,N_4191,N_4442);
nor U4934 (N_4934,N_4056,N_4034);
nand U4935 (N_4935,N_4340,N_4452);
nor U4936 (N_4936,N_4086,N_4325);
nor U4937 (N_4937,N_4074,N_4158);
and U4938 (N_4938,N_4115,N_4371);
nand U4939 (N_4939,N_4208,N_4113);
and U4940 (N_4940,N_4445,N_4460);
and U4941 (N_4941,N_4052,N_4367);
and U4942 (N_4942,N_4387,N_4140);
nor U4943 (N_4943,N_4382,N_4230);
nand U4944 (N_4944,N_4076,N_4236);
nand U4945 (N_4945,N_4266,N_4313);
xor U4946 (N_4946,N_4116,N_4041);
nand U4947 (N_4947,N_4416,N_4421);
nor U4948 (N_4948,N_4005,N_4107);
nand U4949 (N_4949,N_4051,N_4473);
nor U4950 (N_4950,N_4298,N_4432);
nand U4951 (N_4951,N_4200,N_4475);
nor U4952 (N_4952,N_4054,N_4457);
or U4953 (N_4953,N_4034,N_4118);
or U4954 (N_4954,N_4371,N_4378);
or U4955 (N_4955,N_4113,N_4309);
nand U4956 (N_4956,N_4031,N_4328);
xor U4957 (N_4957,N_4069,N_4353);
nor U4958 (N_4958,N_4389,N_4158);
or U4959 (N_4959,N_4195,N_4351);
or U4960 (N_4960,N_4235,N_4091);
nand U4961 (N_4961,N_4060,N_4425);
and U4962 (N_4962,N_4184,N_4110);
nor U4963 (N_4963,N_4034,N_4243);
and U4964 (N_4964,N_4101,N_4221);
nand U4965 (N_4965,N_4492,N_4358);
nor U4966 (N_4966,N_4174,N_4255);
nand U4967 (N_4967,N_4446,N_4374);
xnor U4968 (N_4968,N_4099,N_4426);
and U4969 (N_4969,N_4286,N_4480);
nand U4970 (N_4970,N_4436,N_4198);
nor U4971 (N_4971,N_4210,N_4410);
nor U4972 (N_4972,N_4495,N_4206);
nand U4973 (N_4973,N_4238,N_4044);
or U4974 (N_4974,N_4430,N_4160);
nor U4975 (N_4975,N_4345,N_4452);
nor U4976 (N_4976,N_4379,N_4310);
and U4977 (N_4977,N_4487,N_4142);
nor U4978 (N_4978,N_4349,N_4380);
and U4979 (N_4979,N_4176,N_4389);
and U4980 (N_4980,N_4432,N_4159);
xnor U4981 (N_4981,N_4005,N_4301);
or U4982 (N_4982,N_4014,N_4090);
nand U4983 (N_4983,N_4411,N_4240);
and U4984 (N_4984,N_4298,N_4373);
nor U4985 (N_4985,N_4326,N_4495);
nor U4986 (N_4986,N_4084,N_4429);
xnor U4987 (N_4987,N_4105,N_4121);
or U4988 (N_4988,N_4387,N_4038);
xnor U4989 (N_4989,N_4431,N_4420);
xor U4990 (N_4990,N_4282,N_4065);
nand U4991 (N_4991,N_4264,N_4436);
nor U4992 (N_4992,N_4233,N_4461);
or U4993 (N_4993,N_4485,N_4057);
nand U4994 (N_4994,N_4336,N_4155);
nand U4995 (N_4995,N_4221,N_4321);
nor U4996 (N_4996,N_4096,N_4356);
and U4997 (N_4997,N_4433,N_4316);
and U4998 (N_4998,N_4327,N_4044);
or U4999 (N_4999,N_4437,N_4019);
nand U5000 (N_5000,N_4571,N_4562);
and U5001 (N_5001,N_4937,N_4727);
or U5002 (N_5002,N_4600,N_4776);
or U5003 (N_5003,N_4744,N_4775);
nand U5004 (N_5004,N_4558,N_4541);
nand U5005 (N_5005,N_4979,N_4871);
xnor U5006 (N_5006,N_4750,N_4816);
or U5007 (N_5007,N_4517,N_4985);
nor U5008 (N_5008,N_4971,N_4608);
and U5009 (N_5009,N_4934,N_4585);
xnor U5010 (N_5010,N_4714,N_4789);
nor U5011 (N_5011,N_4689,N_4784);
nor U5012 (N_5012,N_4567,N_4901);
xor U5013 (N_5013,N_4959,N_4722);
or U5014 (N_5014,N_4768,N_4576);
nor U5015 (N_5015,N_4657,N_4659);
xor U5016 (N_5016,N_4919,N_4592);
xor U5017 (N_5017,N_4552,N_4640);
or U5018 (N_5018,N_4580,N_4831);
and U5019 (N_5019,N_4693,N_4596);
and U5020 (N_5020,N_4728,N_4876);
or U5021 (N_5021,N_4634,N_4879);
nor U5022 (N_5022,N_4760,N_4621);
nand U5023 (N_5023,N_4664,N_4606);
nand U5024 (N_5024,N_4795,N_4595);
and U5025 (N_5025,N_4837,N_4527);
or U5026 (N_5026,N_4745,N_4683);
or U5027 (N_5027,N_4601,N_4681);
xor U5028 (N_5028,N_4720,N_4636);
xnor U5029 (N_5029,N_4582,N_4854);
or U5030 (N_5030,N_4617,N_4822);
nand U5031 (N_5031,N_4607,N_4533);
xnor U5032 (N_5032,N_4642,N_4836);
nor U5033 (N_5033,N_4992,N_4652);
or U5034 (N_5034,N_4654,N_4612);
nor U5035 (N_5035,N_4902,N_4883);
and U5036 (N_5036,N_4954,N_4802);
nand U5037 (N_5037,N_4856,N_4785);
nand U5038 (N_5038,N_4885,N_4998);
xor U5039 (N_5039,N_4578,N_4629);
nor U5040 (N_5040,N_4920,N_4922);
and U5041 (N_5041,N_4535,N_4525);
xnor U5042 (N_5042,N_4806,N_4833);
or U5043 (N_5043,N_4872,N_4912);
nand U5044 (N_5044,N_4790,N_4788);
or U5045 (N_5045,N_4889,N_4530);
nor U5046 (N_5046,N_4874,N_4953);
and U5047 (N_5047,N_4544,N_4951);
nand U5048 (N_5048,N_4752,N_4882);
or U5049 (N_5049,N_4986,N_4633);
xor U5050 (N_5050,N_4812,N_4781);
xor U5051 (N_5051,N_4767,N_4529);
nand U5052 (N_5052,N_4565,N_4554);
and U5053 (N_5053,N_4829,N_4620);
xnor U5054 (N_5054,N_4656,N_4555);
and U5055 (N_5055,N_4515,N_4805);
nand U5056 (N_5056,N_4888,N_4605);
and U5057 (N_5057,N_4755,N_4748);
nand U5058 (N_5058,N_4778,N_4809);
nand U5059 (N_5059,N_4947,N_4814);
nand U5060 (N_5060,N_4539,N_4893);
nand U5061 (N_5061,N_4686,N_4740);
or U5062 (N_5062,N_4678,N_4690);
and U5063 (N_5063,N_4512,N_4761);
xor U5064 (N_5064,N_4756,N_4534);
xor U5065 (N_5065,N_4944,N_4993);
or U5066 (N_5066,N_4625,N_4598);
nor U5067 (N_5067,N_4671,N_4647);
xnor U5068 (N_5068,N_4749,N_4930);
and U5069 (N_5069,N_4797,N_4845);
nor U5070 (N_5070,N_4637,N_4653);
or U5071 (N_5071,N_4618,N_4697);
and U5072 (N_5072,N_4923,N_4713);
nand U5073 (N_5073,N_4643,N_4691);
or U5074 (N_5074,N_4589,N_4670);
nor U5075 (N_5075,N_4873,N_4884);
and U5076 (N_5076,N_4970,N_4549);
xor U5077 (N_5077,N_4855,N_4830);
and U5078 (N_5078,N_4905,N_4961);
and U5079 (N_5079,N_4746,N_4940);
and U5080 (N_5080,N_4560,N_4649);
nand U5081 (N_5081,N_4646,N_4863);
xor U5082 (N_5082,N_4556,N_4997);
nor U5083 (N_5083,N_4536,N_4559);
and U5084 (N_5084,N_4502,N_4886);
or U5085 (N_5085,N_4540,N_4957);
and U5086 (N_5086,N_4584,N_4772);
xnor U5087 (N_5087,N_4835,N_4615);
nor U5088 (N_5088,N_4894,N_4878);
and U5089 (N_5089,N_4890,N_4843);
xor U5090 (N_5090,N_4561,N_4751);
xnor U5091 (N_5091,N_4810,N_4907);
and U5092 (N_5092,N_4553,N_4839);
and U5093 (N_5093,N_4604,N_4769);
nand U5094 (N_5094,N_4990,N_4955);
or U5095 (N_5095,N_4983,N_4794);
and U5096 (N_5096,N_4943,N_4861);
nor U5097 (N_5097,N_4548,N_4932);
xor U5098 (N_5098,N_4906,N_4583);
and U5099 (N_5099,N_4631,N_4658);
nor U5100 (N_5100,N_4757,N_4887);
nand U5101 (N_5101,N_4516,N_4729);
nand U5102 (N_5102,N_4648,N_4774);
nand U5103 (N_5103,N_4602,N_4818);
and U5104 (N_5104,N_4586,N_4591);
nand U5105 (N_5105,N_4570,N_4577);
and U5106 (N_5106,N_4715,N_4904);
or U5107 (N_5107,N_4825,N_4733);
nor U5108 (N_5108,N_4635,N_4739);
and U5109 (N_5109,N_4510,N_4526);
xor U5110 (N_5110,N_4661,N_4771);
nor U5111 (N_5111,N_4817,N_4588);
xnor U5112 (N_5112,N_4865,N_4566);
nor U5113 (N_5113,N_4786,N_4844);
or U5114 (N_5114,N_4551,N_4903);
and U5115 (N_5115,N_4813,N_4572);
and U5116 (N_5116,N_4603,N_4834);
nor U5117 (N_5117,N_4868,N_4613);
xor U5118 (N_5118,N_4791,N_4505);
nand U5119 (N_5119,N_4832,N_4827);
nor U5120 (N_5120,N_4796,N_4507);
nor U5121 (N_5121,N_4685,N_4960);
nand U5122 (N_5122,N_4969,N_4931);
nor U5123 (N_5123,N_4972,N_4911);
or U5124 (N_5124,N_4880,N_4842);
nand U5125 (N_5125,N_4680,N_4568);
and U5126 (N_5126,N_4864,N_4910);
xor U5127 (N_5127,N_4838,N_4973);
or U5128 (N_5128,N_4866,N_4917);
nor U5129 (N_5129,N_4674,N_4574);
xor U5130 (N_5130,N_4564,N_4964);
or U5131 (N_5131,N_4718,N_4857);
xnor U5132 (N_5132,N_4927,N_4523);
nand U5133 (N_5133,N_4765,N_4698);
nand U5134 (N_5134,N_4611,N_4736);
nor U5135 (N_5135,N_4754,N_4860);
xnor U5136 (N_5136,N_4895,N_4692);
xor U5137 (N_5137,N_4929,N_4668);
or U5138 (N_5138,N_4773,N_4694);
nand U5139 (N_5139,N_4734,N_4764);
and U5140 (N_5140,N_4594,N_4532);
nor U5141 (N_5141,N_4913,N_4935);
nor U5142 (N_5142,N_4547,N_4859);
and U5143 (N_5143,N_4747,N_4852);
nand U5144 (N_5144,N_4726,N_4853);
or U5145 (N_5145,N_4821,N_4725);
nand U5146 (N_5146,N_4963,N_4735);
xor U5147 (N_5147,N_4676,N_4504);
xnor U5148 (N_5148,N_4641,N_4696);
nand U5149 (N_5149,N_4627,N_4875);
xnor U5150 (N_5150,N_4703,N_4870);
or U5151 (N_5151,N_4522,N_4846);
xor U5152 (N_5152,N_4639,N_4848);
nand U5153 (N_5153,N_4841,N_4705);
nor U5154 (N_5154,N_4682,N_4501);
nand U5155 (N_5155,N_4780,N_4777);
nand U5156 (N_5156,N_4650,N_4952);
nand U5157 (N_5157,N_4675,N_4513);
or U5158 (N_5158,N_4862,N_4921);
nor U5159 (N_5159,N_4924,N_4741);
nand U5160 (N_5160,N_4926,N_4702);
or U5161 (N_5161,N_4801,N_4651);
and U5162 (N_5162,N_4779,N_4766);
or U5163 (N_5163,N_4925,N_4687);
xnor U5164 (N_5164,N_4847,N_4519);
nor U5165 (N_5165,N_4593,N_4975);
and U5166 (N_5166,N_4763,N_4731);
and U5167 (N_5167,N_4669,N_4695);
xor U5168 (N_5168,N_4939,N_4799);
nor U5169 (N_5169,N_4877,N_4826);
and U5170 (N_5170,N_4537,N_4867);
xor U5171 (N_5171,N_4949,N_4711);
or U5172 (N_5172,N_4717,N_4787);
nor U5173 (N_5173,N_4622,N_4614);
nand U5174 (N_5174,N_4978,N_4506);
or U5175 (N_5175,N_4938,N_4770);
or U5176 (N_5176,N_4914,N_4742);
xor U5177 (N_5177,N_4984,N_4798);
and U5178 (N_5178,N_4999,N_4897);
and U5179 (N_5179,N_4996,N_4753);
and U5180 (N_5180,N_4632,N_4758);
or U5181 (N_5181,N_4965,N_4974);
nor U5182 (N_5182,N_4803,N_4508);
xnor U5183 (N_5183,N_4933,N_4850);
and U5184 (N_5184,N_4709,N_4819);
nand U5185 (N_5185,N_4719,N_4968);
nand U5186 (N_5186,N_4503,N_4716);
and U5187 (N_5187,N_4967,N_4898);
nand U5188 (N_5188,N_4531,N_4673);
or U5189 (N_5189,N_4946,N_4958);
xor U5190 (N_5190,N_4916,N_4712);
and U5191 (N_5191,N_4956,N_4597);
and U5192 (N_5192,N_4936,N_4630);
and U5193 (N_5193,N_4950,N_4977);
nand U5194 (N_5194,N_4550,N_4987);
nand U5195 (N_5195,N_4645,N_4684);
nand U5196 (N_5196,N_4701,N_4737);
nand U5197 (N_5197,N_4679,N_4823);
nand U5198 (N_5198,N_4928,N_4660);
and U5199 (N_5199,N_4667,N_4518);
and U5200 (N_5200,N_4824,N_4840);
xnor U5201 (N_5201,N_4948,N_4581);
xnor U5202 (N_5202,N_4579,N_4994);
nor U5203 (N_5203,N_4509,N_4662);
nor U5204 (N_5204,N_4908,N_4546);
or U5205 (N_5205,N_4892,N_4655);
nand U5206 (N_5206,N_4966,N_4677);
nor U5207 (N_5207,N_4538,N_4665);
and U5208 (N_5208,N_4820,N_4616);
or U5209 (N_5209,N_4900,N_4909);
and U5210 (N_5210,N_4706,N_4800);
nor U5211 (N_5211,N_4976,N_4599);
and U5212 (N_5212,N_4783,N_4942);
nor U5213 (N_5213,N_4828,N_4891);
or U5214 (N_5214,N_4995,N_4524);
and U5215 (N_5215,N_4619,N_4980);
and U5216 (N_5216,N_4988,N_4896);
and U5217 (N_5217,N_4626,N_4962);
nor U5218 (N_5218,N_4609,N_4587);
nor U5219 (N_5219,N_4762,N_4918);
and U5220 (N_5220,N_4981,N_4707);
nor U5221 (N_5221,N_4869,N_4557);
and U5222 (N_5222,N_4699,N_4500);
xor U5223 (N_5223,N_4569,N_4521);
and U5224 (N_5224,N_4982,N_4663);
nor U5225 (N_5225,N_4573,N_4815);
nand U5226 (N_5226,N_4782,N_4849);
and U5227 (N_5227,N_4514,N_4666);
xor U5228 (N_5228,N_4623,N_4545);
and U5229 (N_5229,N_4808,N_4542);
or U5230 (N_5230,N_4759,N_4610);
nand U5231 (N_5231,N_4858,N_4941);
and U5232 (N_5232,N_4792,N_4672);
nand U5233 (N_5233,N_4710,N_4881);
nand U5234 (N_5234,N_4528,N_4624);
nor U5235 (N_5235,N_4628,N_4708);
xnor U5236 (N_5236,N_4520,N_4724);
nand U5237 (N_5237,N_4700,N_4738);
xor U5238 (N_5238,N_4899,N_4721);
nor U5239 (N_5239,N_4804,N_4575);
and U5240 (N_5240,N_4851,N_4543);
nor U5241 (N_5241,N_4793,N_4991);
nand U5242 (N_5242,N_4915,N_4945);
xnor U5243 (N_5243,N_4730,N_4638);
nor U5244 (N_5244,N_4590,N_4989);
nand U5245 (N_5245,N_4811,N_4563);
xor U5246 (N_5246,N_4807,N_4688);
or U5247 (N_5247,N_4511,N_4644);
nand U5248 (N_5248,N_4704,N_4743);
nand U5249 (N_5249,N_4732,N_4723);
nand U5250 (N_5250,N_4724,N_4745);
nand U5251 (N_5251,N_4624,N_4900);
or U5252 (N_5252,N_4869,N_4671);
xor U5253 (N_5253,N_4760,N_4776);
nor U5254 (N_5254,N_4977,N_4816);
xor U5255 (N_5255,N_4725,N_4777);
nor U5256 (N_5256,N_4767,N_4750);
nor U5257 (N_5257,N_4971,N_4898);
and U5258 (N_5258,N_4737,N_4757);
nand U5259 (N_5259,N_4739,N_4714);
nor U5260 (N_5260,N_4989,N_4745);
nor U5261 (N_5261,N_4550,N_4622);
xor U5262 (N_5262,N_4985,N_4769);
nor U5263 (N_5263,N_4602,N_4822);
or U5264 (N_5264,N_4987,N_4974);
nand U5265 (N_5265,N_4582,N_4709);
nor U5266 (N_5266,N_4564,N_4919);
or U5267 (N_5267,N_4803,N_4619);
nor U5268 (N_5268,N_4972,N_4715);
or U5269 (N_5269,N_4568,N_4942);
nor U5270 (N_5270,N_4528,N_4883);
nor U5271 (N_5271,N_4763,N_4828);
and U5272 (N_5272,N_4661,N_4580);
nor U5273 (N_5273,N_4876,N_4688);
and U5274 (N_5274,N_4941,N_4662);
or U5275 (N_5275,N_4539,N_4722);
and U5276 (N_5276,N_4965,N_4690);
and U5277 (N_5277,N_4689,N_4556);
xor U5278 (N_5278,N_4535,N_4589);
nand U5279 (N_5279,N_4681,N_4732);
and U5280 (N_5280,N_4594,N_4756);
or U5281 (N_5281,N_4938,N_4753);
nand U5282 (N_5282,N_4564,N_4568);
nand U5283 (N_5283,N_4775,N_4573);
xnor U5284 (N_5284,N_4609,N_4634);
or U5285 (N_5285,N_4586,N_4738);
or U5286 (N_5286,N_4726,N_4944);
nand U5287 (N_5287,N_4642,N_4737);
xnor U5288 (N_5288,N_4867,N_4815);
and U5289 (N_5289,N_4817,N_4988);
nor U5290 (N_5290,N_4829,N_4516);
nand U5291 (N_5291,N_4875,N_4899);
or U5292 (N_5292,N_4767,N_4642);
nand U5293 (N_5293,N_4796,N_4579);
nor U5294 (N_5294,N_4785,N_4561);
or U5295 (N_5295,N_4688,N_4639);
xor U5296 (N_5296,N_4896,N_4568);
or U5297 (N_5297,N_4691,N_4781);
or U5298 (N_5298,N_4688,N_4682);
xor U5299 (N_5299,N_4809,N_4916);
xor U5300 (N_5300,N_4934,N_4959);
xor U5301 (N_5301,N_4564,N_4864);
xnor U5302 (N_5302,N_4797,N_4765);
and U5303 (N_5303,N_4536,N_4779);
nand U5304 (N_5304,N_4577,N_4981);
and U5305 (N_5305,N_4944,N_4702);
nor U5306 (N_5306,N_4864,N_4603);
xnor U5307 (N_5307,N_4898,N_4932);
and U5308 (N_5308,N_4830,N_4633);
nand U5309 (N_5309,N_4699,N_4763);
xnor U5310 (N_5310,N_4943,N_4671);
nor U5311 (N_5311,N_4825,N_4506);
nand U5312 (N_5312,N_4615,N_4627);
nand U5313 (N_5313,N_4980,N_4941);
xor U5314 (N_5314,N_4526,N_4987);
or U5315 (N_5315,N_4936,N_4579);
xnor U5316 (N_5316,N_4927,N_4579);
xnor U5317 (N_5317,N_4916,N_4866);
and U5318 (N_5318,N_4544,N_4861);
xnor U5319 (N_5319,N_4905,N_4914);
nand U5320 (N_5320,N_4628,N_4505);
nand U5321 (N_5321,N_4723,N_4876);
and U5322 (N_5322,N_4577,N_4812);
and U5323 (N_5323,N_4919,N_4863);
nor U5324 (N_5324,N_4528,N_4681);
or U5325 (N_5325,N_4734,N_4678);
and U5326 (N_5326,N_4891,N_4545);
nand U5327 (N_5327,N_4623,N_4939);
nor U5328 (N_5328,N_4723,N_4800);
xnor U5329 (N_5329,N_4939,N_4728);
nand U5330 (N_5330,N_4527,N_4912);
xnor U5331 (N_5331,N_4597,N_4665);
nand U5332 (N_5332,N_4505,N_4957);
and U5333 (N_5333,N_4977,N_4548);
nand U5334 (N_5334,N_4864,N_4593);
xnor U5335 (N_5335,N_4660,N_4751);
nand U5336 (N_5336,N_4600,N_4806);
nor U5337 (N_5337,N_4606,N_4710);
and U5338 (N_5338,N_4827,N_4569);
and U5339 (N_5339,N_4734,N_4521);
xor U5340 (N_5340,N_4701,N_4612);
nand U5341 (N_5341,N_4565,N_4747);
xor U5342 (N_5342,N_4967,N_4915);
xnor U5343 (N_5343,N_4967,N_4974);
nor U5344 (N_5344,N_4916,N_4683);
xnor U5345 (N_5345,N_4576,N_4778);
or U5346 (N_5346,N_4656,N_4878);
nor U5347 (N_5347,N_4704,N_4515);
and U5348 (N_5348,N_4960,N_4598);
nand U5349 (N_5349,N_4651,N_4760);
nor U5350 (N_5350,N_4689,N_4667);
or U5351 (N_5351,N_4549,N_4564);
nor U5352 (N_5352,N_4842,N_4614);
nand U5353 (N_5353,N_4821,N_4940);
and U5354 (N_5354,N_4813,N_4785);
xor U5355 (N_5355,N_4724,N_4585);
nor U5356 (N_5356,N_4617,N_4778);
xnor U5357 (N_5357,N_4643,N_4509);
nor U5358 (N_5358,N_4956,N_4801);
xor U5359 (N_5359,N_4703,N_4616);
nand U5360 (N_5360,N_4762,N_4713);
nor U5361 (N_5361,N_4592,N_4910);
or U5362 (N_5362,N_4551,N_4641);
nor U5363 (N_5363,N_4796,N_4629);
and U5364 (N_5364,N_4507,N_4693);
nand U5365 (N_5365,N_4591,N_4750);
or U5366 (N_5366,N_4536,N_4512);
or U5367 (N_5367,N_4659,N_4982);
xor U5368 (N_5368,N_4733,N_4859);
and U5369 (N_5369,N_4635,N_4849);
xnor U5370 (N_5370,N_4967,N_4671);
nand U5371 (N_5371,N_4976,N_4731);
nand U5372 (N_5372,N_4657,N_4625);
or U5373 (N_5373,N_4607,N_4866);
nand U5374 (N_5374,N_4967,N_4971);
or U5375 (N_5375,N_4905,N_4956);
nor U5376 (N_5376,N_4582,N_4978);
xor U5377 (N_5377,N_4578,N_4888);
xnor U5378 (N_5378,N_4799,N_4547);
nor U5379 (N_5379,N_4637,N_4535);
and U5380 (N_5380,N_4621,N_4752);
nand U5381 (N_5381,N_4924,N_4675);
or U5382 (N_5382,N_4751,N_4771);
nand U5383 (N_5383,N_4934,N_4648);
nor U5384 (N_5384,N_4999,N_4843);
or U5385 (N_5385,N_4960,N_4728);
and U5386 (N_5386,N_4908,N_4928);
and U5387 (N_5387,N_4728,N_4969);
or U5388 (N_5388,N_4872,N_4784);
nand U5389 (N_5389,N_4904,N_4649);
xor U5390 (N_5390,N_4633,N_4968);
and U5391 (N_5391,N_4636,N_4888);
xnor U5392 (N_5392,N_4782,N_4823);
xnor U5393 (N_5393,N_4848,N_4866);
xor U5394 (N_5394,N_4885,N_4700);
xor U5395 (N_5395,N_4817,N_4783);
and U5396 (N_5396,N_4707,N_4848);
xor U5397 (N_5397,N_4752,N_4632);
nor U5398 (N_5398,N_4789,N_4681);
xor U5399 (N_5399,N_4570,N_4553);
nor U5400 (N_5400,N_4609,N_4599);
xor U5401 (N_5401,N_4531,N_4911);
nor U5402 (N_5402,N_4638,N_4720);
or U5403 (N_5403,N_4698,N_4762);
or U5404 (N_5404,N_4842,N_4800);
nand U5405 (N_5405,N_4753,N_4536);
nand U5406 (N_5406,N_4859,N_4611);
and U5407 (N_5407,N_4620,N_4537);
and U5408 (N_5408,N_4654,N_4505);
nor U5409 (N_5409,N_4819,N_4600);
nand U5410 (N_5410,N_4615,N_4910);
or U5411 (N_5411,N_4893,N_4908);
or U5412 (N_5412,N_4629,N_4621);
and U5413 (N_5413,N_4922,N_4519);
nor U5414 (N_5414,N_4556,N_4777);
and U5415 (N_5415,N_4950,N_4876);
nand U5416 (N_5416,N_4658,N_4644);
and U5417 (N_5417,N_4503,N_4755);
or U5418 (N_5418,N_4945,N_4907);
or U5419 (N_5419,N_4927,N_4829);
and U5420 (N_5420,N_4565,N_4644);
and U5421 (N_5421,N_4527,N_4885);
nand U5422 (N_5422,N_4514,N_4725);
xnor U5423 (N_5423,N_4922,N_4862);
and U5424 (N_5424,N_4523,N_4892);
nor U5425 (N_5425,N_4554,N_4874);
or U5426 (N_5426,N_4865,N_4789);
nor U5427 (N_5427,N_4766,N_4611);
and U5428 (N_5428,N_4568,N_4988);
nand U5429 (N_5429,N_4801,N_4782);
nand U5430 (N_5430,N_4691,N_4763);
xor U5431 (N_5431,N_4700,N_4538);
and U5432 (N_5432,N_4973,N_4830);
xor U5433 (N_5433,N_4701,N_4943);
or U5434 (N_5434,N_4934,N_4768);
xnor U5435 (N_5435,N_4986,N_4907);
nand U5436 (N_5436,N_4518,N_4992);
and U5437 (N_5437,N_4868,N_4859);
nand U5438 (N_5438,N_4541,N_4524);
nand U5439 (N_5439,N_4679,N_4730);
and U5440 (N_5440,N_4879,N_4899);
xor U5441 (N_5441,N_4539,N_4688);
or U5442 (N_5442,N_4748,N_4664);
or U5443 (N_5443,N_4833,N_4881);
xor U5444 (N_5444,N_4760,N_4983);
and U5445 (N_5445,N_4718,N_4871);
or U5446 (N_5446,N_4930,N_4685);
xnor U5447 (N_5447,N_4645,N_4960);
and U5448 (N_5448,N_4821,N_4997);
nand U5449 (N_5449,N_4590,N_4707);
nand U5450 (N_5450,N_4707,N_4800);
and U5451 (N_5451,N_4791,N_4935);
nor U5452 (N_5452,N_4994,N_4510);
nor U5453 (N_5453,N_4521,N_4744);
xor U5454 (N_5454,N_4685,N_4900);
and U5455 (N_5455,N_4956,N_4687);
nor U5456 (N_5456,N_4977,N_4933);
or U5457 (N_5457,N_4528,N_4546);
or U5458 (N_5458,N_4762,N_4881);
xor U5459 (N_5459,N_4673,N_4837);
nand U5460 (N_5460,N_4677,N_4583);
nor U5461 (N_5461,N_4751,N_4911);
xor U5462 (N_5462,N_4846,N_4934);
or U5463 (N_5463,N_4844,N_4600);
or U5464 (N_5464,N_4546,N_4841);
or U5465 (N_5465,N_4739,N_4683);
xor U5466 (N_5466,N_4955,N_4768);
nand U5467 (N_5467,N_4519,N_4678);
xnor U5468 (N_5468,N_4933,N_4822);
and U5469 (N_5469,N_4780,N_4839);
and U5470 (N_5470,N_4649,N_4728);
or U5471 (N_5471,N_4633,N_4741);
nor U5472 (N_5472,N_4765,N_4703);
nand U5473 (N_5473,N_4676,N_4983);
and U5474 (N_5474,N_4551,N_4775);
and U5475 (N_5475,N_4839,N_4650);
nand U5476 (N_5476,N_4544,N_4857);
nand U5477 (N_5477,N_4959,N_4730);
nand U5478 (N_5478,N_4880,N_4567);
nand U5479 (N_5479,N_4707,N_4545);
xnor U5480 (N_5480,N_4624,N_4656);
or U5481 (N_5481,N_4700,N_4634);
and U5482 (N_5482,N_4910,N_4626);
and U5483 (N_5483,N_4973,N_4844);
nand U5484 (N_5484,N_4742,N_4578);
nor U5485 (N_5485,N_4618,N_4830);
or U5486 (N_5486,N_4553,N_4507);
xnor U5487 (N_5487,N_4520,N_4510);
nor U5488 (N_5488,N_4619,N_4899);
or U5489 (N_5489,N_4541,N_4919);
nor U5490 (N_5490,N_4553,N_4921);
and U5491 (N_5491,N_4845,N_4633);
xnor U5492 (N_5492,N_4794,N_4560);
xor U5493 (N_5493,N_4895,N_4878);
and U5494 (N_5494,N_4669,N_4988);
and U5495 (N_5495,N_4668,N_4619);
and U5496 (N_5496,N_4957,N_4941);
xnor U5497 (N_5497,N_4868,N_4588);
xnor U5498 (N_5498,N_4912,N_4669);
nand U5499 (N_5499,N_4938,N_4897);
nor U5500 (N_5500,N_5383,N_5172);
nor U5501 (N_5501,N_5347,N_5211);
or U5502 (N_5502,N_5319,N_5270);
nand U5503 (N_5503,N_5258,N_5047);
nand U5504 (N_5504,N_5001,N_5108);
or U5505 (N_5505,N_5360,N_5042);
nand U5506 (N_5506,N_5326,N_5216);
xnor U5507 (N_5507,N_5345,N_5123);
nand U5508 (N_5508,N_5025,N_5200);
or U5509 (N_5509,N_5139,N_5105);
nor U5510 (N_5510,N_5014,N_5133);
and U5511 (N_5511,N_5438,N_5463);
xnor U5512 (N_5512,N_5128,N_5066);
or U5513 (N_5513,N_5155,N_5412);
xor U5514 (N_5514,N_5013,N_5080);
or U5515 (N_5515,N_5441,N_5387);
nand U5516 (N_5516,N_5353,N_5004);
nand U5517 (N_5517,N_5000,N_5465);
and U5518 (N_5518,N_5402,N_5174);
and U5519 (N_5519,N_5269,N_5473);
and U5520 (N_5520,N_5430,N_5286);
nand U5521 (N_5521,N_5194,N_5079);
nand U5522 (N_5522,N_5418,N_5295);
nor U5523 (N_5523,N_5135,N_5264);
xor U5524 (N_5524,N_5459,N_5164);
nand U5525 (N_5525,N_5146,N_5343);
nand U5526 (N_5526,N_5087,N_5218);
and U5527 (N_5527,N_5284,N_5043);
nand U5528 (N_5528,N_5197,N_5027);
xor U5529 (N_5529,N_5092,N_5364);
and U5530 (N_5530,N_5140,N_5190);
or U5531 (N_5531,N_5202,N_5196);
and U5532 (N_5532,N_5136,N_5103);
and U5533 (N_5533,N_5424,N_5228);
and U5534 (N_5534,N_5131,N_5121);
nand U5535 (N_5535,N_5254,N_5086);
or U5536 (N_5536,N_5476,N_5165);
nand U5537 (N_5537,N_5354,N_5210);
and U5538 (N_5538,N_5395,N_5049);
or U5539 (N_5539,N_5415,N_5166);
or U5540 (N_5540,N_5127,N_5491);
xnor U5541 (N_5541,N_5321,N_5130);
and U5542 (N_5542,N_5431,N_5367);
and U5543 (N_5543,N_5330,N_5485);
xnor U5544 (N_5544,N_5192,N_5024);
nor U5545 (N_5545,N_5104,N_5420);
xor U5546 (N_5546,N_5428,N_5094);
nand U5547 (N_5547,N_5339,N_5052);
xor U5548 (N_5548,N_5062,N_5177);
nor U5549 (N_5549,N_5058,N_5113);
xnor U5550 (N_5550,N_5309,N_5300);
nor U5551 (N_5551,N_5159,N_5229);
nor U5552 (N_5552,N_5257,N_5016);
nor U5553 (N_5553,N_5214,N_5436);
nor U5554 (N_5554,N_5322,N_5288);
nor U5555 (N_5555,N_5278,N_5296);
nor U5556 (N_5556,N_5102,N_5088);
nand U5557 (N_5557,N_5150,N_5203);
and U5558 (N_5558,N_5209,N_5022);
and U5559 (N_5559,N_5020,N_5070);
nor U5560 (N_5560,N_5496,N_5276);
nand U5561 (N_5561,N_5224,N_5391);
and U5562 (N_5562,N_5084,N_5499);
and U5563 (N_5563,N_5290,N_5186);
and U5564 (N_5564,N_5494,N_5472);
nor U5565 (N_5565,N_5077,N_5124);
and U5566 (N_5566,N_5028,N_5002);
nor U5567 (N_5567,N_5467,N_5265);
xor U5568 (N_5568,N_5031,N_5495);
nand U5569 (N_5569,N_5149,N_5493);
and U5570 (N_5570,N_5095,N_5452);
xor U5571 (N_5571,N_5312,N_5289);
nor U5572 (N_5572,N_5437,N_5114);
xnor U5573 (N_5573,N_5247,N_5026);
xnor U5574 (N_5574,N_5169,N_5248);
nor U5575 (N_5575,N_5018,N_5010);
nor U5576 (N_5576,N_5335,N_5032);
and U5577 (N_5577,N_5435,N_5446);
xnor U5578 (N_5578,N_5481,N_5413);
nor U5579 (N_5579,N_5372,N_5241);
or U5580 (N_5580,N_5157,N_5313);
and U5581 (N_5581,N_5484,N_5426);
nor U5582 (N_5582,N_5199,N_5451);
or U5583 (N_5583,N_5362,N_5225);
xor U5584 (N_5584,N_5255,N_5337);
and U5585 (N_5585,N_5294,N_5320);
nand U5586 (N_5586,N_5408,N_5332);
xnor U5587 (N_5587,N_5386,N_5423);
or U5588 (N_5588,N_5129,N_5480);
and U5589 (N_5589,N_5434,N_5110);
or U5590 (N_5590,N_5015,N_5223);
nor U5591 (N_5591,N_5277,N_5138);
nand U5592 (N_5592,N_5279,N_5275);
nor U5593 (N_5593,N_5120,N_5447);
and U5594 (N_5594,N_5245,N_5093);
nor U5595 (N_5595,N_5268,N_5097);
and U5596 (N_5596,N_5057,N_5083);
nand U5597 (N_5597,N_5204,N_5274);
nor U5598 (N_5598,N_5271,N_5310);
nand U5599 (N_5599,N_5250,N_5444);
and U5600 (N_5600,N_5338,N_5324);
xnor U5601 (N_5601,N_5464,N_5369);
xnor U5602 (N_5602,N_5398,N_5375);
or U5603 (N_5603,N_5163,N_5302);
or U5604 (N_5604,N_5023,N_5053);
nor U5605 (N_5605,N_5282,N_5403);
and U5606 (N_5606,N_5063,N_5041);
and U5607 (N_5607,N_5045,N_5407);
xor U5608 (N_5608,N_5030,N_5429);
nand U5609 (N_5609,N_5244,N_5189);
nand U5610 (N_5610,N_5346,N_5448);
nand U5611 (N_5611,N_5478,N_5389);
nor U5612 (N_5612,N_5055,N_5073);
nand U5613 (N_5613,N_5409,N_5401);
xor U5614 (N_5614,N_5201,N_5344);
nand U5615 (N_5615,N_5005,N_5239);
or U5616 (N_5616,N_5267,N_5126);
nand U5617 (N_5617,N_5176,N_5457);
xnor U5618 (N_5618,N_5205,N_5370);
nand U5619 (N_5619,N_5230,N_5217);
nand U5620 (N_5620,N_5327,N_5068);
or U5621 (N_5621,N_5242,N_5100);
and U5622 (N_5622,N_5143,N_5411);
nor U5623 (N_5623,N_5263,N_5078);
xor U5624 (N_5624,N_5328,N_5109);
nand U5625 (N_5625,N_5112,N_5158);
xor U5626 (N_5626,N_5445,N_5272);
and U5627 (N_5627,N_5237,N_5019);
and U5628 (N_5628,N_5154,N_5184);
nand U5629 (N_5629,N_5060,N_5222);
nand U5630 (N_5630,N_5396,N_5323);
and U5631 (N_5631,N_5082,N_5456);
nand U5632 (N_5632,N_5293,N_5074);
or U5633 (N_5633,N_5308,N_5450);
or U5634 (N_5634,N_5352,N_5151);
nand U5635 (N_5635,N_5051,N_5388);
and U5636 (N_5636,N_5171,N_5231);
nand U5637 (N_5637,N_5365,N_5221);
nand U5638 (N_5638,N_5035,N_5116);
and U5639 (N_5639,N_5492,N_5260);
nand U5640 (N_5640,N_5208,N_5153);
and U5641 (N_5641,N_5317,N_5351);
nor U5642 (N_5642,N_5475,N_5356);
nand U5643 (N_5643,N_5009,N_5181);
and U5644 (N_5644,N_5368,N_5329);
nand U5645 (N_5645,N_5243,N_5119);
or U5646 (N_5646,N_5477,N_5469);
or U5647 (N_5647,N_5262,N_5291);
or U5648 (N_5648,N_5331,N_5350);
nor U5649 (N_5649,N_5357,N_5067);
xnor U5650 (N_5650,N_5029,N_5099);
xnor U5651 (N_5651,N_5318,N_5349);
or U5652 (N_5652,N_5012,N_5482);
nand U5653 (N_5653,N_5191,N_5301);
and U5654 (N_5654,N_5311,N_5392);
xor U5655 (N_5655,N_5361,N_5161);
nand U5656 (N_5656,N_5316,N_5050);
nor U5657 (N_5657,N_5363,N_5393);
and U5658 (N_5658,N_5195,N_5238);
and U5659 (N_5659,N_5040,N_5474);
and U5660 (N_5660,N_5152,N_5442);
and U5661 (N_5661,N_5213,N_5334);
or U5662 (N_5662,N_5054,N_5366);
xor U5663 (N_5663,N_5240,N_5090);
xnor U5664 (N_5664,N_5283,N_5227);
xor U5665 (N_5665,N_5410,N_5377);
nor U5666 (N_5666,N_5468,N_5376);
nand U5667 (N_5667,N_5417,N_5175);
or U5668 (N_5668,N_5137,N_5458);
nor U5669 (N_5669,N_5185,N_5056);
and U5670 (N_5670,N_5454,N_5416);
xor U5671 (N_5671,N_5106,N_5433);
xor U5672 (N_5672,N_5285,N_5215);
or U5673 (N_5673,N_5179,N_5098);
and U5674 (N_5674,N_5385,N_5384);
xnor U5675 (N_5675,N_5359,N_5156);
nand U5676 (N_5676,N_5399,N_5455);
or U5677 (N_5677,N_5183,N_5443);
nor U5678 (N_5678,N_5497,N_5479);
nor U5679 (N_5679,N_5358,N_5091);
nand U5680 (N_5680,N_5460,N_5287);
or U5681 (N_5681,N_5008,N_5315);
nand U5682 (N_5682,N_5065,N_5187);
or U5683 (N_5683,N_5142,N_5414);
and U5684 (N_5684,N_5305,N_5406);
nand U5685 (N_5685,N_5132,N_5235);
nand U5686 (N_5686,N_5397,N_5044);
xnor U5687 (N_5687,N_5036,N_5096);
or U5688 (N_5688,N_5355,N_5168);
xnor U5689 (N_5689,N_5011,N_5348);
xor U5690 (N_5690,N_5076,N_5226);
nand U5691 (N_5691,N_5341,N_5382);
and U5692 (N_5692,N_5303,N_5483);
xor U5693 (N_5693,N_5118,N_5232);
nand U5694 (N_5694,N_5380,N_5003);
xor U5695 (N_5695,N_5234,N_5390);
and U5696 (N_5696,N_5085,N_5182);
or U5697 (N_5697,N_5251,N_5212);
nor U5698 (N_5698,N_5404,N_5148);
nand U5699 (N_5699,N_5374,N_5160);
nor U5700 (N_5700,N_5034,N_5314);
or U5701 (N_5701,N_5256,N_5466);
nor U5702 (N_5702,N_5236,N_5178);
nand U5703 (N_5703,N_5486,N_5421);
xnor U5704 (N_5704,N_5340,N_5147);
or U5705 (N_5705,N_5273,N_5453);
xnor U5706 (N_5706,N_5081,N_5115);
nand U5707 (N_5707,N_5427,N_5281);
nand U5708 (N_5708,N_5432,N_5069);
nor U5709 (N_5709,N_5373,N_5259);
and U5710 (N_5710,N_5048,N_5233);
nand U5711 (N_5711,N_5198,N_5145);
and U5712 (N_5712,N_5336,N_5007);
nor U5713 (N_5713,N_5122,N_5333);
nor U5714 (N_5714,N_5266,N_5280);
xnor U5715 (N_5715,N_5379,N_5101);
nor U5716 (N_5716,N_5246,N_5206);
xnor U5717 (N_5717,N_5461,N_5173);
xnor U5718 (N_5718,N_5072,N_5371);
or U5719 (N_5719,N_5180,N_5046);
nand U5720 (N_5720,N_5075,N_5449);
or U5721 (N_5721,N_5306,N_5117);
nor U5722 (N_5722,N_5419,N_5470);
nor U5723 (N_5723,N_5219,N_5342);
and U5724 (N_5724,N_5249,N_5089);
and U5725 (N_5725,N_5033,N_5193);
or U5726 (N_5726,N_5298,N_5021);
nor U5727 (N_5727,N_5498,N_5207);
xnor U5728 (N_5728,N_5440,N_5299);
nand U5729 (N_5729,N_5170,N_5039);
nor U5730 (N_5730,N_5292,N_5107);
nand U5731 (N_5731,N_5006,N_5425);
and U5732 (N_5732,N_5422,N_5071);
or U5733 (N_5733,N_5111,N_5261);
nand U5734 (N_5734,N_5167,N_5188);
or U5735 (N_5735,N_5141,N_5125);
and U5736 (N_5736,N_5325,N_5059);
nand U5737 (N_5737,N_5490,N_5405);
nor U5738 (N_5738,N_5017,N_5144);
xor U5739 (N_5739,N_5307,N_5297);
xnor U5740 (N_5740,N_5064,N_5394);
and U5741 (N_5741,N_5304,N_5400);
or U5742 (N_5742,N_5162,N_5253);
xor U5743 (N_5743,N_5252,N_5381);
nor U5744 (N_5744,N_5487,N_5471);
xnor U5745 (N_5745,N_5489,N_5488);
and U5746 (N_5746,N_5220,N_5378);
nor U5747 (N_5747,N_5061,N_5038);
or U5748 (N_5748,N_5037,N_5134);
and U5749 (N_5749,N_5439,N_5462);
and U5750 (N_5750,N_5168,N_5254);
nand U5751 (N_5751,N_5115,N_5323);
and U5752 (N_5752,N_5257,N_5238);
and U5753 (N_5753,N_5019,N_5470);
or U5754 (N_5754,N_5426,N_5082);
nand U5755 (N_5755,N_5261,N_5483);
and U5756 (N_5756,N_5075,N_5316);
nor U5757 (N_5757,N_5404,N_5253);
nand U5758 (N_5758,N_5433,N_5393);
and U5759 (N_5759,N_5139,N_5054);
xnor U5760 (N_5760,N_5486,N_5479);
or U5761 (N_5761,N_5206,N_5196);
nor U5762 (N_5762,N_5226,N_5004);
or U5763 (N_5763,N_5177,N_5024);
nor U5764 (N_5764,N_5028,N_5189);
and U5765 (N_5765,N_5408,N_5181);
or U5766 (N_5766,N_5013,N_5372);
and U5767 (N_5767,N_5050,N_5068);
or U5768 (N_5768,N_5193,N_5270);
xor U5769 (N_5769,N_5077,N_5455);
or U5770 (N_5770,N_5139,N_5377);
xor U5771 (N_5771,N_5457,N_5014);
or U5772 (N_5772,N_5414,N_5021);
or U5773 (N_5773,N_5154,N_5053);
nand U5774 (N_5774,N_5304,N_5050);
or U5775 (N_5775,N_5012,N_5454);
xor U5776 (N_5776,N_5150,N_5184);
xor U5777 (N_5777,N_5073,N_5165);
and U5778 (N_5778,N_5233,N_5251);
nand U5779 (N_5779,N_5198,N_5335);
nand U5780 (N_5780,N_5468,N_5476);
xnor U5781 (N_5781,N_5309,N_5495);
nand U5782 (N_5782,N_5324,N_5303);
and U5783 (N_5783,N_5376,N_5115);
xor U5784 (N_5784,N_5044,N_5078);
or U5785 (N_5785,N_5178,N_5367);
or U5786 (N_5786,N_5084,N_5145);
or U5787 (N_5787,N_5147,N_5166);
or U5788 (N_5788,N_5293,N_5003);
xor U5789 (N_5789,N_5104,N_5351);
and U5790 (N_5790,N_5010,N_5334);
or U5791 (N_5791,N_5476,N_5176);
or U5792 (N_5792,N_5263,N_5175);
and U5793 (N_5793,N_5052,N_5422);
nor U5794 (N_5794,N_5212,N_5122);
or U5795 (N_5795,N_5176,N_5213);
nand U5796 (N_5796,N_5285,N_5150);
nor U5797 (N_5797,N_5184,N_5442);
nor U5798 (N_5798,N_5236,N_5075);
xor U5799 (N_5799,N_5022,N_5289);
nand U5800 (N_5800,N_5117,N_5249);
nand U5801 (N_5801,N_5014,N_5409);
xor U5802 (N_5802,N_5267,N_5487);
and U5803 (N_5803,N_5223,N_5276);
and U5804 (N_5804,N_5291,N_5071);
nand U5805 (N_5805,N_5113,N_5004);
or U5806 (N_5806,N_5452,N_5384);
or U5807 (N_5807,N_5213,N_5347);
and U5808 (N_5808,N_5425,N_5455);
nand U5809 (N_5809,N_5102,N_5013);
nor U5810 (N_5810,N_5417,N_5119);
xnor U5811 (N_5811,N_5384,N_5130);
and U5812 (N_5812,N_5377,N_5233);
and U5813 (N_5813,N_5097,N_5008);
nand U5814 (N_5814,N_5328,N_5187);
nand U5815 (N_5815,N_5098,N_5431);
or U5816 (N_5816,N_5075,N_5201);
and U5817 (N_5817,N_5372,N_5416);
or U5818 (N_5818,N_5294,N_5157);
xor U5819 (N_5819,N_5415,N_5115);
nand U5820 (N_5820,N_5058,N_5117);
or U5821 (N_5821,N_5199,N_5394);
or U5822 (N_5822,N_5363,N_5065);
nor U5823 (N_5823,N_5423,N_5469);
nor U5824 (N_5824,N_5051,N_5078);
xor U5825 (N_5825,N_5365,N_5387);
and U5826 (N_5826,N_5372,N_5205);
or U5827 (N_5827,N_5108,N_5181);
or U5828 (N_5828,N_5100,N_5438);
and U5829 (N_5829,N_5489,N_5293);
nand U5830 (N_5830,N_5358,N_5065);
nor U5831 (N_5831,N_5006,N_5166);
xor U5832 (N_5832,N_5372,N_5068);
nand U5833 (N_5833,N_5446,N_5004);
nor U5834 (N_5834,N_5183,N_5305);
or U5835 (N_5835,N_5304,N_5142);
xnor U5836 (N_5836,N_5330,N_5128);
nand U5837 (N_5837,N_5069,N_5113);
and U5838 (N_5838,N_5012,N_5440);
and U5839 (N_5839,N_5418,N_5095);
and U5840 (N_5840,N_5414,N_5403);
or U5841 (N_5841,N_5418,N_5025);
xor U5842 (N_5842,N_5438,N_5246);
and U5843 (N_5843,N_5122,N_5136);
or U5844 (N_5844,N_5243,N_5448);
nor U5845 (N_5845,N_5176,N_5159);
nor U5846 (N_5846,N_5279,N_5494);
and U5847 (N_5847,N_5360,N_5464);
or U5848 (N_5848,N_5321,N_5397);
nor U5849 (N_5849,N_5497,N_5054);
or U5850 (N_5850,N_5194,N_5008);
nor U5851 (N_5851,N_5038,N_5437);
nand U5852 (N_5852,N_5458,N_5087);
or U5853 (N_5853,N_5487,N_5059);
nand U5854 (N_5854,N_5391,N_5078);
or U5855 (N_5855,N_5065,N_5371);
xor U5856 (N_5856,N_5258,N_5431);
nor U5857 (N_5857,N_5414,N_5101);
nor U5858 (N_5858,N_5382,N_5292);
xnor U5859 (N_5859,N_5454,N_5412);
and U5860 (N_5860,N_5112,N_5343);
xnor U5861 (N_5861,N_5335,N_5116);
or U5862 (N_5862,N_5164,N_5426);
xnor U5863 (N_5863,N_5418,N_5240);
or U5864 (N_5864,N_5279,N_5122);
and U5865 (N_5865,N_5008,N_5080);
or U5866 (N_5866,N_5247,N_5178);
xor U5867 (N_5867,N_5248,N_5181);
xnor U5868 (N_5868,N_5031,N_5013);
and U5869 (N_5869,N_5086,N_5413);
xor U5870 (N_5870,N_5323,N_5138);
xor U5871 (N_5871,N_5447,N_5149);
xnor U5872 (N_5872,N_5396,N_5219);
nor U5873 (N_5873,N_5222,N_5195);
xnor U5874 (N_5874,N_5225,N_5128);
or U5875 (N_5875,N_5182,N_5258);
nor U5876 (N_5876,N_5010,N_5341);
or U5877 (N_5877,N_5226,N_5184);
nand U5878 (N_5878,N_5155,N_5206);
and U5879 (N_5879,N_5283,N_5082);
nor U5880 (N_5880,N_5309,N_5323);
nand U5881 (N_5881,N_5253,N_5024);
and U5882 (N_5882,N_5104,N_5413);
and U5883 (N_5883,N_5178,N_5093);
nand U5884 (N_5884,N_5057,N_5388);
or U5885 (N_5885,N_5003,N_5140);
xnor U5886 (N_5886,N_5204,N_5093);
nor U5887 (N_5887,N_5068,N_5091);
and U5888 (N_5888,N_5100,N_5188);
or U5889 (N_5889,N_5039,N_5084);
nor U5890 (N_5890,N_5480,N_5178);
and U5891 (N_5891,N_5229,N_5336);
nor U5892 (N_5892,N_5101,N_5269);
nand U5893 (N_5893,N_5114,N_5409);
nand U5894 (N_5894,N_5353,N_5381);
xnor U5895 (N_5895,N_5450,N_5098);
nor U5896 (N_5896,N_5042,N_5488);
xnor U5897 (N_5897,N_5038,N_5326);
and U5898 (N_5898,N_5298,N_5011);
xnor U5899 (N_5899,N_5382,N_5158);
and U5900 (N_5900,N_5188,N_5445);
and U5901 (N_5901,N_5329,N_5209);
nor U5902 (N_5902,N_5069,N_5293);
or U5903 (N_5903,N_5238,N_5422);
and U5904 (N_5904,N_5033,N_5007);
nand U5905 (N_5905,N_5280,N_5371);
xnor U5906 (N_5906,N_5030,N_5168);
nor U5907 (N_5907,N_5295,N_5412);
or U5908 (N_5908,N_5485,N_5030);
or U5909 (N_5909,N_5180,N_5397);
nand U5910 (N_5910,N_5198,N_5105);
or U5911 (N_5911,N_5244,N_5042);
nand U5912 (N_5912,N_5138,N_5272);
nand U5913 (N_5913,N_5439,N_5384);
nand U5914 (N_5914,N_5246,N_5083);
and U5915 (N_5915,N_5387,N_5282);
or U5916 (N_5916,N_5100,N_5352);
nand U5917 (N_5917,N_5169,N_5275);
nand U5918 (N_5918,N_5041,N_5304);
xnor U5919 (N_5919,N_5297,N_5490);
nand U5920 (N_5920,N_5311,N_5242);
and U5921 (N_5921,N_5031,N_5429);
and U5922 (N_5922,N_5016,N_5336);
and U5923 (N_5923,N_5310,N_5449);
nand U5924 (N_5924,N_5244,N_5105);
nor U5925 (N_5925,N_5219,N_5290);
nand U5926 (N_5926,N_5188,N_5000);
nand U5927 (N_5927,N_5371,N_5118);
xnor U5928 (N_5928,N_5445,N_5093);
or U5929 (N_5929,N_5064,N_5401);
xnor U5930 (N_5930,N_5228,N_5034);
xnor U5931 (N_5931,N_5235,N_5267);
and U5932 (N_5932,N_5161,N_5135);
xor U5933 (N_5933,N_5076,N_5038);
nor U5934 (N_5934,N_5485,N_5328);
xor U5935 (N_5935,N_5428,N_5404);
nor U5936 (N_5936,N_5434,N_5302);
nand U5937 (N_5937,N_5165,N_5487);
nand U5938 (N_5938,N_5103,N_5457);
or U5939 (N_5939,N_5343,N_5262);
nor U5940 (N_5940,N_5126,N_5113);
and U5941 (N_5941,N_5175,N_5454);
nor U5942 (N_5942,N_5112,N_5240);
or U5943 (N_5943,N_5101,N_5049);
nor U5944 (N_5944,N_5348,N_5342);
nand U5945 (N_5945,N_5368,N_5080);
nor U5946 (N_5946,N_5230,N_5050);
xor U5947 (N_5947,N_5261,N_5205);
nor U5948 (N_5948,N_5271,N_5329);
or U5949 (N_5949,N_5480,N_5477);
nor U5950 (N_5950,N_5051,N_5025);
or U5951 (N_5951,N_5166,N_5237);
xnor U5952 (N_5952,N_5298,N_5147);
nor U5953 (N_5953,N_5100,N_5472);
nor U5954 (N_5954,N_5052,N_5396);
nand U5955 (N_5955,N_5293,N_5231);
xor U5956 (N_5956,N_5485,N_5494);
or U5957 (N_5957,N_5165,N_5259);
and U5958 (N_5958,N_5155,N_5064);
nor U5959 (N_5959,N_5421,N_5133);
nor U5960 (N_5960,N_5357,N_5249);
nand U5961 (N_5961,N_5237,N_5099);
nand U5962 (N_5962,N_5487,N_5294);
and U5963 (N_5963,N_5437,N_5331);
nor U5964 (N_5964,N_5490,N_5477);
xnor U5965 (N_5965,N_5262,N_5298);
xor U5966 (N_5966,N_5224,N_5383);
nor U5967 (N_5967,N_5009,N_5344);
xnor U5968 (N_5968,N_5365,N_5437);
nand U5969 (N_5969,N_5186,N_5103);
nor U5970 (N_5970,N_5179,N_5042);
or U5971 (N_5971,N_5325,N_5130);
nor U5972 (N_5972,N_5077,N_5319);
xnor U5973 (N_5973,N_5301,N_5003);
or U5974 (N_5974,N_5468,N_5400);
or U5975 (N_5975,N_5020,N_5218);
and U5976 (N_5976,N_5053,N_5320);
nor U5977 (N_5977,N_5015,N_5389);
and U5978 (N_5978,N_5243,N_5126);
and U5979 (N_5979,N_5163,N_5011);
nor U5980 (N_5980,N_5011,N_5178);
nand U5981 (N_5981,N_5429,N_5112);
or U5982 (N_5982,N_5448,N_5095);
and U5983 (N_5983,N_5132,N_5301);
nand U5984 (N_5984,N_5197,N_5028);
and U5985 (N_5985,N_5220,N_5178);
nor U5986 (N_5986,N_5489,N_5037);
nand U5987 (N_5987,N_5374,N_5198);
nand U5988 (N_5988,N_5301,N_5361);
nand U5989 (N_5989,N_5115,N_5225);
xnor U5990 (N_5990,N_5282,N_5073);
nand U5991 (N_5991,N_5313,N_5387);
nand U5992 (N_5992,N_5192,N_5158);
and U5993 (N_5993,N_5442,N_5315);
and U5994 (N_5994,N_5114,N_5405);
or U5995 (N_5995,N_5475,N_5327);
nor U5996 (N_5996,N_5245,N_5097);
xnor U5997 (N_5997,N_5236,N_5281);
and U5998 (N_5998,N_5488,N_5069);
nand U5999 (N_5999,N_5201,N_5043);
and U6000 (N_6000,N_5851,N_5788);
xnor U6001 (N_6001,N_5961,N_5684);
nor U6002 (N_6002,N_5725,N_5667);
nor U6003 (N_6003,N_5565,N_5824);
and U6004 (N_6004,N_5838,N_5839);
xnor U6005 (N_6005,N_5945,N_5853);
or U6006 (N_6006,N_5847,N_5624);
or U6007 (N_6007,N_5514,N_5934);
nor U6008 (N_6008,N_5694,N_5748);
nand U6009 (N_6009,N_5596,N_5644);
nor U6010 (N_6010,N_5737,N_5680);
nand U6011 (N_6011,N_5549,N_5799);
or U6012 (N_6012,N_5807,N_5515);
xor U6013 (N_6013,N_5783,N_5670);
xnor U6014 (N_6014,N_5500,N_5995);
or U6015 (N_6015,N_5903,N_5960);
nor U6016 (N_6016,N_5637,N_5912);
or U6017 (N_6017,N_5560,N_5883);
and U6018 (N_6018,N_5774,N_5917);
or U6019 (N_6019,N_5869,N_5908);
and U6020 (N_6020,N_5622,N_5700);
nor U6021 (N_6021,N_5587,N_5522);
and U6022 (N_6022,N_5724,N_5742);
nand U6023 (N_6023,N_5863,N_5829);
or U6024 (N_6024,N_5875,N_5593);
xnor U6025 (N_6025,N_5821,N_5982);
xor U6026 (N_6026,N_5603,N_5764);
or U6027 (N_6027,N_5765,N_5709);
nand U6028 (N_6028,N_5915,N_5517);
nand U6029 (N_6029,N_5999,N_5729);
or U6030 (N_6030,N_5502,N_5755);
xnor U6031 (N_6031,N_5609,N_5954);
and U6032 (N_6032,N_5744,N_5556);
nand U6033 (N_6033,N_5928,N_5859);
xnor U6034 (N_6034,N_5902,N_5842);
nor U6035 (N_6035,N_5761,N_5657);
or U6036 (N_6036,N_5930,N_5526);
nor U6037 (N_6037,N_5787,N_5938);
nand U6038 (N_6038,N_5980,N_5538);
or U6039 (N_6039,N_5595,N_5998);
nor U6040 (N_6040,N_5758,N_5846);
and U6041 (N_6041,N_5527,N_5638);
or U6042 (N_6042,N_5707,N_5586);
and U6043 (N_6043,N_5837,N_5688);
or U6044 (N_6044,N_5958,N_5594);
and U6045 (N_6045,N_5918,N_5813);
nor U6046 (N_6046,N_5802,N_5905);
nand U6047 (N_6047,N_5721,N_5735);
nor U6048 (N_6048,N_5582,N_5981);
and U6049 (N_6049,N_5641,N_5857);
and U6050 (N_6050,N_5743,N_5723);
or U6051 (N_6051,N_5592,N_5814);
and U6052 (N_6052,N_5898,N_5965);
nor U6053 (N_6053,N_5642,N_5844);
nor U6054 (N_6054,N_5551,N_5574);
xor U6055 (N_6055,N_5550,N_5886);
or U6056 (N_6056,N_5907,N_5553);
nand U6057 (N_6057,N_5727,N_5955);
nand U6058 (N_6058,N_5873,N_5800);
nand U6059 (N_6059,N_5913,N_5614);
xor U6060 (N_6060,N_5932,N_5579);
or U6061 (N_6061,N_5703,N_5664);
nand U6062 (N_6062,N_5936,N_5541);
nand U6063 (N_6063,N_5880,N_5504);
and U6064 (N_6064,N_5510,N_5796);
and U6065 (N_6065,N_5752,N_5557);
nand U6066 (N_6066,N_5793,N_5805);
or U6067 (N_6067,N_5507,N_5652);
nand U6068 (N_6068,N_5823,N_5605);
nand U6069 (N_6069,N_5786,N_5740);
or U6070 (N_6070,N_5810,N_5732);
or U6071 (N_6071,N_5705,N_5525);
xor U6072 (N_6072,N_5792,N_5992);
xnor U6073 (N_6073,N_5971,N_5834);
nand U6074 (N_6074,N_5542,N_5922);
nand U6075 (N_6075,N_5711,N_5983);
and U6076 (N_6076,N_5626,N_5921);
or U6077 (N_6077,N_5619,N_5690);
xnor U6078 (N_6078,N_5756,N_5884);
or U6079 (N_6079,N_5675,N_5899);
nor U6080 (N_6080,N_5896,N_5655);
nand U6081 (N_6081,N_5762,N_5658);
nand U6082 (N_6082,N_5734,N_5686);
or U6083 (N_6083,N_5720,N_5760);
and U6084 (N_6084,N_5841,N_5589);
nor U6085 (N_6085,N_5996,N_5620);
xor U6086 (N_6086,N_5662,N_5848);
and U6087 (N_6087,N_5911,N_5830);
nand U6088 (N_6088,N_5598,N_5833);
and U6089 (N_6089,N_5763,N_5768);
or U6090 (N_6090,N_5575,N_5512);
and U6091 (N_6091,N_5570,N_5816);
xnor U6092 (N_6092,N_5716,N_5590);
nand U6093 (N_6093,N_5822,N_5754);
or U6094 (N_6094,N_5613,N_5858);
and U6095 (N_6095,N_5910,N_5519);
xor U6096 (N_6096,N_5818,N_5781);
nor U6097 (N_6097,N_5803,N_5804);
or U6098 (N_6098,N_5782,N_5789);
xor U6099 (N_6099,N_5618,N_5511);
and U6100 (N_6100,N_5649,N_5948);
nor U6101 (N_6101,N_5564,N_5651);
nand U6102 (N_6102,N_5989,N_5860);
nor U6103 (N_6103,N_5719,N_5940);
or U6104 (N_6104,N_5682,N_5591);
nand U6105 (N_6105,N_5806,N_5604);
and U6106 (N_6106,N_5997,N_5600);
nand U6107 (N_6107,N_5628,N_5632);
nor U6108 (N_6108,N_5673,N_5862);
and U6109 (N_6109,N_5672,N_5656);
nor U6110 (N_6110,N_5654,N_5866);
nor U6111 (N_6111,N_5695,N_5828);
and U6112 (N_6112,N_5558,N_5665);
nor U6113 (N_6113,N_5933,N_5972);
and U6114 (N_6114,N_5925,N_5881);
xor U6115 (N_6115,N_5530,N_5710);
nand U6116 (N_6116,N_5636,N_5518);
nand U6117 (N_6117,N_5949,N_5906);
or U6118 (N_6118,N_5617,N_5701);
or U6119 (N_6119,N_5878,N_5947);
xor U6120 (N_6120,N_5819,N_5931);
or U6121 (N_6121,N_5820,N_5661);
or U6122 (N_6122,N_5766,N_5890);
or U6123 (N_6123,N_5685,N_5887);
or U6124 (N_6124,N_5699,N_5785);
xnor U6125 (N_6125,N_5795,N_5750);
or U6126 (N_6126,N_5533,N_5585);
nor U6127 (N_6127,N_5916,N_5660);
nand U6128 (N_6128,N_5865,N_5769);
nand U6129 (N_6129,N_5731,N_5777);
or U6130 (N_6130,N_5825,N_5676);
nor U6131 (N_6131,N_5775,N_5508);
or U6132 (N_6132,N_5943,N_5942);
and U6133 (N_6133,N_5726,N_5715);
and U6134 (N_6134,N_5689,N_5856);
xnor U6135 (N_6135,N_5864,N_5536);
nand U6136 (N_6136,N_5580,N_5950);
nand U6137 (N_6137,N_5513,N_5611);
and U6138 (N_6138,N_5736,N_5767);
xor U6139 (N_6139,N_5581,N_5872);
xor U6140 (N_6140,N_5966,N_5683);
nor U6141 (N_6141,N_5634,N_5547);
xnor U6142 (N_6142,N_5607,N_5555);
or U6143 (N_6143,N_5879,N_5751);
and U6144 (N_6144,N_5854,N_5631);
xnor U6145 (N_6145,N_5576,N_5693);
xnor U6146 (N_6146,N_5811,N_5956);
nor U6147 (N_6147,N_5653,N_5868);
or U6148 (N_6148,N_5691,N_5979);
or U6149 (N_6149,N_5733,N_5988);
or U6150 (N_6150,N_5718,N_5509);
nand U6151 (N_6151,N_5779,N_5772);
nor U6152 (N_6152,N_5633,N_5924);
and U6153 (N_6153,N_5974,N_5569);
xnor U6154 (N_6154,N_5648,N_5738);
nor U6155 (N_6155,N_5554,N_5871);
or U6156 (N_6156,N_5987,N_5937);
nor U6157 (N_6157,N_5893,N_5669);
nor U6158 (N_6158,N_5832,N_5753);
nand U6159 (N_6159,N_5749,N_5745);
xnor U6160 (N_6160,N_5602,N_5967);
xnor U6161 (N_6161,N_5840,N_5534);
and U6162 (N_6162,N_5537,N_5717);
xor U6163 (N_6163,N_5612,N_5708);
xor U6164 (N_6164,N_5601,N_5874);
nand U6165 (N_6165,N_5535,N_5901);
xor U6166 (N_6166,N_5876,N_5870);
or U6167 (N_6167,N_5927,N_5888);
and U6168 (N_6168,N_5826,N_5608);
xor U6169 (N_6169,N_5935,N_5704);
xnor U6170 (N_6170,N_5546,N_5698);
nand U6171 (N_6171,N_5559,N_5953);
or U6172 (N_6172,N_5714,N_5650);
nor U6173 (N_6173,N_5757,N_5571);
nand U6174 (N_6174,N_5895,N_5817);
xnor U6175 (N_6175,N_5706,N_5978);
nand U6176 (N_6176,N_5894,N_5797);
xor U6177 (N_6177,N_5794,N_5520);
xnor U6178 (N_6178,N_5835,N_5900);
or U6179 (N_6179,N_5759,N_5973);
nand U6180 (N_6180,N_5926,N_5990);
or U6181 (N_6181,N_5827,N_5929);
and U6182 (N_6182,N_5852,N_5531);
and U6183 (N_6183,N_5572,N_5728);
nand U6184 (N_6184,N_5712,N_5970);
or U6185 (N_6185,N_5503,N_5532);
and U6186 (N_6186,N_5643,N_5798);
or U6187 (N_6187,N_5677,N_5645);
and U6188 (N_6188,N_5616,N_5573);
xnor U6189 (N_6189,N_5791,N_5944);
or U6190 (N_6190,N_5597,N_5505);
xnor U6191 (N_6191,N_5599,N_5778);
or U6192 (N_6192,N_5666,N_5584);
or U6193 (N_6193,N_5625,N_5516);
and U6194 (N_6194,N_5784,N_5747);
nor U6195 (N_6195,N_5528,N_5615);
or U6196 (N_6196,N_5681,N_5563);
nand U6197 (N_6197,N_5882,N_5836);
and U6198 (N_6198,N_5663,N_5831);
nor U6199 (N_6199,N_5964,N_5968);
or U6200 (N_6200,N_5845,N_5952);
or U6201 (N_6201,N_5877,N_5773);
nand U6202 (N_6202,N_5909,N_5889);
xor U6203 (N_6203,N_5539,N_5780);
xnor U6204 (N_6204,N_5543,N_5976);
and U6205 (N_6205,N_5739,N_5850);
xnor U6206 (N_6206,N_5588,N_5812);
xor U6207 (N_6207,N_5963,N_5977);
nand U6208 (N_6208,N_5891,N_5969);
and U6209 (N_6209,N_5920,N_5696);
nor U6210 (N_6210,N_5627,N_5746);
and U6211 (N_6211,N_5545,N_5986);
xor U6212 (N_6212,N_5523,N_5951);
and U6213 (N_6213,N_5771,N_5959);
nor U6214 (N_6214,N_5640,N_5561);
nor U6215 (N_6215,N_5776,N_5692);
xor U6216 (N_6216,N_5741,N_5668);
nor U6217 (N_6217,N_5578,N_5897);
nor U6218 (N_6218,N_5730,N_5702);
or U6219 (N_6219,N_5548,N_5809);
nor U6220 (N_6220,N_5529,N_5985);
or U6221 (N_6221,N_5506,N_5659);
or U6222 (N_6222,N_5904,N_5639);
nor U6223 (N_6223,N_5713,N_5994);
xor U6224 (N_6224,N_5957,N_5674);
and U6225 (N_6225,N_5962,N_5861);
nor U6226 (N_6226,N_5501,N_5843);
or U6227 (N_6227,N_5566,N_5849);
and U6228 (N_6228,N_5524,N_5583);
and U6229 (N_6229,N_5540,N_5671);
and U6230 (N_6230,N_5647,N_5679);
nand U6231 (N_6231,N_5867,N_5623);
nor U6232 (N_6232,N_5770,N_5790);
xnor U6233 (N_6233,N_5919,N_5808);
and U6234 (N_6234,N_5687,N_5521);
and U6235 (N_6235,N_5939,N_5562);
and U6236 (N_6236,N_5568,N_5606);
nand U6237 (N_6237,N_5914,N_5815);
nor U6238 (N_6238,N_5567,N_5635);
nor U6239 (N_6239,N_5577,N_5984);
or U6240 (N_6240,N_5646,N_5544);
xor U6241 (N_6241,N_5975,N_5885);
nand U6242 (N_6242,N_5629,N_5678);
or U6243 (N_6243,N_5993,N_5610);
nand U6244 (N_6244,N_5923,N_5697);
nor U6245 (N_6245,N_5892,N_5941);
nor U6246 (N_6246,N_5722,N_5855);
xor U6247 (N_6247,N_5630,N_5801);
or U6248 (N_6248,N_5621,N_5946);
and U6249 (N_6249,N_5991,N_5552);
nor U6250 (N_6250,N_5790,N_5549);
nor U6251 (N_6251,N_5886,N_5925);
nor U6252 (N_6252,N_5787,N_5670);
or U6253 (N_6253,N_5699,N_5745);
or U6254 (N_6254,N_5552,N_5973);
or U6255 (N_6255,N_5558,N_5603);
nor U6256 (N_6256,N_5775,N_5597);
nand U6257 (N_6257,N_5820,N_5934);
nand U6258 (N_6258,N_5757,N_5507);
nand U6259 (N_6259,N_5906,N_5979);
xor U6260 (N_6260,N_5557,N_5654);
or U6261 (N_6261,N_5825,N_5500);
and U6262 (N_6262,N_5631,N_5509);
xor U6263 (N_6263,N_5674,N_5845);
nand U6264 (N_6264,N_5835,N_5593);
nor U6265 (N_6265,N_5845,N_5924);
xor U6266 (N_6266,N_5932,N_5925);
nand U6267 (N_6267,N_5606,N_5857);
nand U6268 (N_6268,N_5684,N_5753);
nand U6269 (N_6269,N_5675,N_5522);
nor U6270 (N_6270,N_5971,N_5753);
or U6271 (N_6271,N_5821,N_5850);
or U6272 (N_6272,N_5750,N_5892);
xnor U6273 (N_6273,N_5852,N_5952);
nand U6274 (N_6274,N_5577,N_5857);
nor U6275 (N_6275,N_5751,N_5987);
and U6276 (N_6276,N_5581,N_5610);
nand U6277 (N_6277,N_5760,N_5509);
and U6278 (N_6278,N_5761,N_5986);
and U6279 (N_6279,N_5957,N_5551);
nor U6280 (N_6280,N_5743,N_5703);
and U6281 (N_6281,N_5570,N_5589);
and U6282 (N_6282,N_5607,N_5897);
nor U6283 (N_6283,N_5961,N_5520);
xnor U6284 (N_6284,N_5554,N_5601);
nand U6285 (N_6285,N_5568,N_5908);
or U6286 (N_6286,N_5579,N_5667);
nand U6287 (N_6287,N_5635,N_5613);
nor U6288 (N_6288,N_5989,N_5923);
nand U6289 (N_6289,N_5893,N_5766);
nand U6290 (N_6290,N_5597,N_5610);
nor U6291 (N_6291,N_5980,N_5639);
nand U6292 (N_6292,N_5935,N_5793);
and U6293 (N_6293,N_5503,N_5980);
or U6294 (N_6294,N_5627,N_5753);
or U6295 (N_6295,N_5996,N_5694);
xnor U6296 (N_6296,N_5868,N_5517);
nand U6297 (N_6297,N_5871,N_5699);
nor U6298 (N_6298,N_5756,N_5532);
nor U6299 (N_6299,N_5700,N_5767);
and U6300 (N_6300,N_5522,N_5659);
or U6301 (N_6301,N_5949,N_5702);
or U6302 (N_6302,N_5821,N_5863);
or U6303 (N_6303,N_5859,N_5962);
nand U6304 (N_6304,N_5693,N_5762);
or U6305 (N_6305,N_5530,N_5543);
or U6306 (N_6306,N_5752,N_5665);
nor U6307 (N_6307,N_5666,N_5951);
or U6308 (N_6308,N_5880,N_5537);
xor U6309 (N_6309,N_5789,N_5506);
and U6310 (N_6310,N_5930,N_5906);
nand U6311 (N_6311,N_5814,N_5557);
and U6312 (N_6312,N_5905,N_5919);
nand U6313 (N_6313,N_5510,N_5921);
and U6314 (N_6314,N_5771,N_5803);
xnor U6315 (N_6315,N_5936,N_5754);
and U6316 (N_6316,N_5823,N_5565);
xnor U6317 (N_6317,N_5556,N_5874);
nand U6318 (N_6318,N_5688,N_5575);
and U6319 (N_6319,N_5863,N_5563);
xor U6320 (N_6320,N_5649,N_5554);
nor U6321 (N_6321,N_5677,N_5508);
nor U6322 (N_6322,N_5735,N_5673);
nand U6323 (N_6323,N_5857,N_5570);
and U6324 (N_6324,N_5733,N_5804);
xor U6325 (N_6325,N_5640,N_5548);
nand U6326 (N_6326,N_5650,N_5687);
xor U6327 (N_6327,N_5638,N_5779);
or U6328 (N_6328,N_5853,N_5906);
xnor U6329 (N_6329,N_5590,N_5776);
and U6330 (N_6330,N_5949,N_5684);
nand U6331 (N_6331,N_5809,N_5534);
nand U6332 (N_6332,N_5825,N_5811);
or U6333 (N_6333,N_5908,N_5712);
or U6334 (N_6334,N_5672,N_5646);
xor U6335 (N_6335,N_5952,N_5802);
and U6336 (N_6336,N_5613,N_5678);
nand U6337 (N_6337,N_5576,N_5774);
nand U6338 (N_6338,N_5981,N_5742);
and U6339 (N_6339,N_5724,N_5714);
nor U6340 (N_6340,N_5840,N_5929);
nand U6341 (N_6341,N_5794,N_5732);
nor U6342 (N_6342,N_5818,N_5833);
or U6343 (N_6343,N_5605,N_5592);
or U6344 (N_6344,N_5778,N_5654);
or U6345 (N_6345,N_5967,N_5541);
xnor U6346 (N_6346,N_5943,N_5658);
xnor U6347 (N_6347,N_5595,N_5702);
nor U6348 (N_6348,N_5714,N_5522);
nand U6349 (N_6349,N_5585,N_5921);
and U6350 (N_6350,N_5857,N_5802);
or U6351 (N_6351,N_5748,N_5799);
nor U6352 (N_6352,N_5571,N_5985);
and U6353 (N_6353,N_5570,N_5594);
xor U6354 (N_6354,N_5704,N_5875);
nor U6355 (N_6355,N_5620,N_5682);
and U6356 (N_6356,N_5535,N_5974);
or U6357 (N_6357,N_5965,N_5535);
nor U6358 (N_6358,N_5796,N_5945);
xor U6359 (N_6359,N_5689,N_5503);
xor U6360 (N_6360,N_5524,N_5531);
and U6361 (N_6361,N_5879,N_5999);
or U6362 (N_6362,N_5760,N_5950);
and U6363 (N_6363,N_5799,N_5820);
nor U6364 (N_6364,N_5666,N_5519);
and U6365 (N_6365,N_5908,N_5649);
xnor U6366 (N_6366,N_5622,N_5610);
xnor U6367 (N_6367,N_5896,N_5608);
or U6368 (N_6368,N_5702,N_5602);
xor U6369 (N_6369,N_5556,N_5814);
nor U6370 (N_6370,N_5850,N_5859);
and U6371 (N_6371,N_5892,N_5809);
nor U6372 (N_6372,N_5773,N_5546);
xor U6373 (N_6373,N_5927,N_5857);
nand U6374 (N_6374,N_5650,N_5583);
or U6375 (N_6375,N_5825,N_5935);
xnor U6376 (N_6376,N_5958,N_5502);
nand U6377 (N_6377,N_5708,N_5726);
nand U6378 (N_6378,N_5528,N_5506);
xnor U6379 (N_6379,N_5614,N_5872);
and U6380 (N_6380,N_5840,N_5633);
nor U6381 (N_6381,N_5738,N_5737);
nand U6382 (N_6382,N_5536,N_5692);
xnor U6383 (N_6383,N_5826,N_5752);
xor U6384 (N_6384,N_5806,N_5983);
nand U6385 (N_6385,N_5952,N_5922);
nand U6386 (N_6386,N_5825,N_5630);
nand U6387 (N_6387,N_5520,N_5877);
nand U6388 (N_6388,N_5660,N_5885);
xor U6389 (N_6389,N_5732,N_5697);
xnor U6390 (N_6390,N_5962,N_5714);
xor U6391 (N_6391,N_5550,N_5675);
nand U6392 (N_6392,N_5748,N_5813);
xnor U6393 (N_6393,N_5665,N_5667);
and U6394 (N_6394,N_5647,N_5633);
nor U6395 (N_6395,N_5904,N_5553);
xnor U6396 (N_6396,N_5530,N_5787);
nand U6397 (N_6397,N_5580,N_5628);
nand U6398 (N_6398,N_5576,N_5905);
xor U6399 (N_6399,N_5936,N_5904);
and U6400 (N_6400,N_5851,N_5818);
and U6401 (N_6401,N_5739,N_5938);
xnor U6402 (N_6402,N_5522,N_5669);
nor U6403 (N_6403,N_5884,N_5762);
nor U6404 (N_6404,N_5751,N_5511);
xor U6405 (N_6405,N_5892,N_5846);
xor U6406 (N_6406,N_5554,N_5982);
and U6407 (N_6407,N_5732,N_5793);
nand U6408 (N_6408,N_5860,N_5780);
nor U6409 (N_6409,N_5963,N_5633);
or U6410 (N_6410,N_5542,N_5872);
and U6411 (N_6411,N_5710,N_5747);
and U6412 (N_6412,N_5595,N_5915);
and U6413 (N_6413,N_5797,N_5853);
xnor U6414 (N_6414,N_5666,N_5912);
and U6415 (N_6415,N_5533,N_5726);
xnor U6416 (N_6416,N_5557,N_5827);
nor U6417 (N_6417,N_5772,N_5719);
xnor U6418 (N_6418,N_5698,N_5607);
and U6419 (N_6419,N_5857,N_5867);
xnor U6420 (N_6420,N_5965,N_5652);
or U6421 (N_6421,N_5785,N_5908);
and U6422 (N_6422,N_5881,N_5569);
and U6423 (N_6423,N_5723,N_5594);
and U6424 (N_6424,N_5597,N_5637);
xnor U6425 (N_6425,N_5655,N_5996);
and U6426 (N_6426,N_5896,N_5783);
and U6427 (N_6427,N_5903,N_5577);
or U6428 (N_6428,N_5739,N_5932);
and U6429 (N_6429,N_5755,N_5654);
or U6430 (N_6430,N_5782,N_5787);
or U6431 (N_6431,N_5824,N_5561);
nand U6432 (N_6432,N_5869,N_5627);
xor U6433 (N_6433,N_5991,N_5855);
or U6434 (N_6434,N_5928,N_5611);
nand U6435 (N_6435,N_5674,N_5867);
and U6436 (N_6436,N_5768,N_5548);
nand U6437 (N_6437,N_5719,N_5711);
and U6438 (N_6438,N_5790,N_5716);
or U6439 (N_6439,N_5956,N_5935);
and U6440 (N_6440,N_5738,N_5820);
xnor U6441 (N_6441,N_5762,N_5967);
or U6442 (N_6442,N_5876,N_5585);
or U6443 (N_6443,N_5525,N_5844);
xor U6444 (N_6444,N_5944,N_5934);
xor U6445 (N_6445,N_5822,N_5562);
nand U6446 (N_6446,N_5845,N_5560);
and U6447 (N_6447,N_5884,N_5934);
xnor U6448 (N_6448,N_5812,N_5524);
nor U6449 (N_6449,N_5595,N_5849);
or U6450 (N_6450,N_5508,N_5784);
nand U6451 (N_6451,N_5945,N_5670);
or U6452 (N_6452,N_5539,N_5868);
and U6453 (N_6453,N_5865,N_5733);
or U6454 (N_6454,N_5753,N_5820);
nand U6455 (N_6455,N_5516,N_5673);
xnor U6456 (N_6456,N_5613,N_5694);
nor U6457 (N_6457,N_5780,N_5850);
or U6458 (N_6458,N_5912,N_5893);
nand U6459 (N_6459,N_5774,N_5877);
xor U6460 (N_6460,N_5576,N_5811);
nand U6461 (N_6461,N_5808,N_5681);
and U6462 (N_6462,N_5778,N_5829);
nor U6463 (N_6463,N_5837,N_5979);
nor U6464 (N_6464,N_5801,N_5893);
nor U6465 (N_6465,N_5787,N_5659);
nand U6466 (N_6466,N_5677,N_5594);
xnor U6467 (N_6467,N_5702,N_5998);
nand U6468 (N_6468,N_5992,N_5553);
and U6469 (N_6469,N_5873,N_5946);
or U6470 (N_6470,N_5978,N_5842);
nand U6471 (N_6471,N_5761,N_5556);
or U6472 (N_6472,N_5519,N_5995);
nor U6473 (N_6473,N_5764,N_5886);
and U6474 (N_6474,N_5956,N_5839);
or U6475 (N_6475,N_5619,N_5822);
xnor U6476 (N_6476,N_5909,N_5739);
nor U6477 (N_6477,N_5811,N_5750);
nor U6478 (N_6478,N_5821,N_5667);
and U6479 (N_6479,N_5529,N_5947);
nor U6480 (N_6480,N_5934,N_5881);
nor U6481 (N_6481,N_5681,N_5713);
and U6482 (N_6482,N_5651,N_5853);
nand U6483 (N_6483,N_5565,N_5902);
xnor U6484 (N_6484,N_5571,N_5594);
nand U6485 (N_6485,N_5724,N_5739);
and U6486 (N_6486,N_5763,N_5636);
nand U6487 (N_6487,N_5565,N_5641);
and U6488 (N_6488,N_5852,N_5656);
nand U6489 (N_6489,N_5728,N_5653);
or U6490 (N_6490,N_5534,N_5689);
nand U6491 (N_6491,N_5500,N_5763);
or U6492 (N_6492,N_5524,N_5796);
xnor U6493 (N_6493,N_5520,N_5938);
and U6494 (N_6494,N_5988,N_5819);
nor U6495 (N_6495,N_5587,N_5572);
nor U6496 (N_6496,N_5882,N_5738);
and U6497 (N_6497,N_5972,N_5918);
xnor U6498 (N_6498,N_5527,N_5740);
nor U6499 (N_6499,N_5935,N_5981);
or U6500 (N_6500,N_6045,N_6380);
nand U6501 (N_6501,N_6484,N_6324);
and U6502 (N_6502,N_6462,N_6261);
xnor U6503 (N_6503,N_6478,N_6094);
nand U6504 (N_6504,N_6059,N_6170);
nand U6505 (N_6505,N_6432,N_6134);
and U6506 (N_6506,N_6471,N_6158);
xor U6507 (N_6507,N_6041,N_6202);
nand U6508 (N_6508,N_6099,N_6294);
and U6509 (N_6509,N_6358,N_6066);
and U6510 (N_6510,N_6239,N_6068);
or U6511 (N_6511,N_6269,N_6145);
or U6512 (N_6512,N_6057,N_6424);
nor U6513 (N_6513,N_6402,N_6119);
nand U6514 (N_6514,N_6397,N_6191);
xnor U6515 (N_6515,N_6043,N_6051);
or U6516 (N_6516,N_6328,N_6496);
nand U6517 (N_6517,N_6002,N_6296);
nor U6518 (N_6518,N_6105,N_6179);
or U6519 (N_6519,N_6480,N_6448);
xor U6520 (N_6520,N_6076,N_6477);
xor U6521 (N_6521,N_6089,N_6123);
xor U6522 (N_6522,N_6102,N_6166);
and U6523 (N_6523,N_6423,N_6137);
nor U6524 (N_6524,N_6273,N_6193);
nand U6525 (N_6525,N_6443,N_6385);
or U6526 (N_6526,N_6309,N_6131);
nand U6527 (N_6527,N_6052,N_6081);
nor U6528 (N_6528,N_6064,N_6310);
and U6529 (N_6529,N_6135,N_6155);
and U6530 (N_6530,N_6121,N_6330);
nor U6531 (N_6531,N_6214,N_6195);
and U6532 (N_6532,N_6409,N_6001);
nand U6533 (N_6533,N_6047,N_6283);
nor U6534 (N_6534,N_6483,N_6469);
nand U6535 (N_6535,N_6108,N_6168);
nor U6536 (N_6536,N_6097,N_6071);
nand U6537 (N_6537,N_6410,N_6067);
nor U6538 (N_6538,N_6388,N_6357);
nor U6539 (N_6539,N_6046,N_6184);
xor U6540 (N_6540,N_6420,N_6014);
xnor U6541 (N_6541,N_6061,N_6023);
nand U6542 (N_6542,N_6055,N_6378);
nor U6543 (N_6543,N_6449,N_6444);
or U6544 (N_6544,N_6271,N_6189);
xor U6545 (N_6545,N_6229,N_6264);
nand U6546 (N_6546,N_6418,N_6147);
xor U6547 (N_6547,N_6298,N_6178);
nand U6548 (N_6548,N_6116,N_6465);
xnor U6549 (N_6549,N_6242,N_6441);
nand U6550 (N_6550,N_6476,N_6115);
or U6551 (N_6551,N_6408,N_6005);
or U6552 (N_6552,N_6257,N_6212);
xnor U6553 (N_6553,N_6042,N_6025);
or U6554 (N_6554,N_6437,N_6350);
nor U6555 (N_6555,N_6054,N_6162);
xnor U6556 (N_6556,N_6232,N_6245);
xor U6557 (N_6557,N_6314,N_6139);
nand U6558 (N_6558,N_6204,N_6405);
or U6559 (N_6559,N_6467,N_6101);
xor U6560 (N_6560,N_6266,N_6348);
xnor U6561 (N_6561,N_6086,N_6370);
nand U6562 (N_6562,N_6197,N_6451);
and U6563 (N_6563,N_6060,N_6156);
nand U6564 (N_6564,N_6065,N_6485);
or U6565 (N_6565,N_6126,N_6369);
nand U6566 (N_6566,N_6459,N_6015);
or U6567 (N_6567,N_6498,N_6285);
xor U6568 (N_6568,N_6417,N_6299);
nand U6569 (N_6569,N_6491,N_6473);
and U6570 (N_6570,N_6048,N_6182);
nor U6571 (N_6571,N_6365,N_6474);
xnor U6572 (N_6572,N_6203,N_6492);
and U6573 (N_6573,N_6083,N_6332);
and U6574 (N_6574,N_6461,N_6305);
or U6575 (N_6575,N_6185,N_6497);
or U6576 (N_6576,N_6406,N_6237);
xor U6577 (N_6577,N_6211,N_6371);
nand U6578 (N_6578,N_6219,N_6367);
or U6579 (N_6579,N_6340,N_6333);
nand U6580 (N_6580,N_6109,N_6248);
nand U6581 (N_6581,N_6347,N_6428);
and U6582 (N_6582,N_6173,N_6130);
and U6583 (N_6583,N_6208,N_6251);
nor U6584 (N_6584,N_6436,N_6470);
and U6585 (N_6585,N_6413,N_6016);
and U6586 (N_6586,N_6021,N_6072);
or U6587 (N_6587,N_6148,N_6411);
nand U6588 (N_6588,N_6398,N_6177);
or U6589 (N_6589,N_6372,N_6058);
and U6590 (N_6590,N_6151,N_6475);
or U6591 (N_6591,N_6138,N_6128);
and U6592 (N_6592,N_6037,N_6289);
or U6593 (N_6593,N_6243,N_6217);
or U6594 (N_6594,N_6260,N_6090);
xor U6595 (N_6595,N_6141,N_6396);
or U6596 (N_6596,N_6114,N_6488);
nand U6597 (N_6597,N_6049,N_6263);
or U6598 (N_6598,N_6323,N_6092);
nand U6599 (N_6599,N_6075,N_6327);
or U6600 (N_6600,N_6206,N_6414);
and U6601 (N_6601,N_6176,N_6150);
nor U6602 (N_6602,N_6387,N_6454);
or U6603 (N_6603,N_6028,N_6201);
nand U6604 (N_6604,N_6456,N_6040);
nor U6605 (N_6605,N_6079,N_6034);
nor U6606 (N_6606,N_6308,N_6249);
nand U6607 (N_6607,N_6044,N_6440);
nor U6608 (N_6608,N_6355,N_6181);
and U6609 (N_6609,N_6425,N_6319);
xnor U6610 (N_6610,N_6012,N_6117);
or U6611 (N_6611,N_6167,N_6032);
nand U6612 (N_6612,N_6062,N_6499);
nand U6613 (N_6613,N_6122,N_6165);
and U6614 (N_6614,N_6172,N_6088);
and U6615 (N_6615,N_6352,N_6258);
nor U6616 (N_6616,N_6133,N_6278);
xnor U6617 (N_6617,N_6169,N_6335);
nor U6618 (N_6618,N_6407,N_6368);
or U6619 (N_6619,N_6228,N_6460);
and U6620 (N_6620,N_6140,N_6284);
xnor U6621 (N_6621,N_6112,N_6056);
nor U6622 (N_6622,N_6174,N_6144);
nor U6623 (N_6623,N_6399,N_6149);
nand U6624 (N_6624,N_6146,N_6254);
or U6625 (N_6625,N_6297,N_6143);
or U6626 (N_6626,N_6275,N_6213);
nor U6627 (N_6627,N_6106,N_6279);
or U6628 (N_6628,N_6224,N_6194);
nand U6629 (N_6629,N_6003,N_6430);
and U6630 (N_6630,N_6455,N_6438);
and U6631 (N_6631,N_6494,N_6427);
xor U6632 (N_6632,N_6389,N_6349);
nor U6633 (N_6633,N_6199,N_6036);
xnor U6634 (N_6634,N_6033,N_6029);
nor U6635 (N_6635,N_6104,N_6220);
or U6636 (N_6636,N_6362,N_6103);
nand U6637 (N_6637,N_6325,N_6196);
xnor U6638 (N_6638,N_6070,N_6267);
or U6639 (N_6639,N_6274,N_6452);
xnor U6640 (N_6640,N_6439,N_6136);
xnor U6641 (N_6641,N_6160,N_6223);
nor U6642 (N_6642,N_6354,N_6486);
nor U6643 (N_6643,N_6447,N_6482);
nor U6644 (N_6644,N_6205,N_6394);
xor U6645 (N_6645,N_6277,N_6069);
nand U6646 (N_6646,N_6290,N_6487);
xnor U6647 (N_6647,N_6154,N_6111);
nand U6648 (N_6648,N_6415,N_6050);
nor U6649 (N_6649,N_6010,N_6233);
and U6650 (N_6650,N_6422,N_6026);
and U6651 (N_6651,N_6256,N_6142);
nand U6652 (N_6652,N_6481,N_6164);
nand U6653 (N_6653,N_6188,N_6035);
nand U6654 (N_6654,N_6391,N_6311);
nand U6655 (N_6655,N_6019,N_6458);
and U6656 (N_6656,N_6157,N_6082);
xnor U6657 (N_6657,N_6286,N_6226);
xor U6658 (N_6658,N_6240,N_6353);
and U6659 (N_6659,N_6343,N_6303);
nor U6660 (N_6660,N_6030,N_6009);
and U6661 (N_6661,N_6288,N_6363);
and U6662 (N_6662,N_6401,N_6073);
nand U6663 (N_6663,N_6376,N_6007);
nand U6664 (N_6664,N_6313,N_6078);
nand U6665 (N_6665,N_6329,N_6281);
nor U6666 (N_6666,N_6107,N_6316);
nand U6667 (N_6667,N_6207,N_6318);
nor U6668 (N_6668,N_6342,N_6011);
nand U6669 (N_6669,N_6024,N_6027);
nand U6670 (N_6670,N_6495,N_6171);
xor U6671 (N_6671,N_6433,N_6493);
xor U6672 (N_6672,N_6464,N_6215);
nand U6673 (N_6673,N_6466,N_6063);
or U6674 (N_6674,N_6221,N_6093);
nand U6675 (N_6675,N_6183,N_6341);
nor U6676 (N_6676,N_6100,N_6361);
nand U6677 (N_6677,N_6091,N_6084);
or U6678 (N_6678,N_6346,N_6390);
nor U6679 (N_6679,N_6360,N_6489);
and U6680 (N_6680,N_6113,N_6375);
nand U6681 (N_6681,N_6295,N_6020);
nor U6682 (N_6682,N_6293,N_6315);
and U6683 (N_6683,N_6312,N_6472);
nor U6684 (N_6684,N_6320,N_6180);
xnor U6685 (N_6685,N_6379,N_6351);
xor U6686 (N_6686,N_6393,N_6234);
and U6687 (N_6687,N_6227,N_6490);
xnor U6688 (N_6688,N_6110,N_6334);
xnor U6689 (N_6689,N_6302,N_6085);
or U6690 (N_6690,N_6331,N_6255);
xnor U6691 (N_6691,N_6236,N_6307);
and U6692 (N_6692,N_6377,N_6374);
xnor U6693 (N_6693,N_6384,N_6426);
and U6694 (N_6694,N_6445,N_6345);
or U6695 (N_6695,N_6022,N_6095);
and U6696 (N_6696,N_6087,N_6175);
xor U6697 (N_6697,N_6317,N_6186);
nand U6698 (N_6698,N_6080,N_6000);
nor U6699 (N_6699,N_6431,N_6247);
or U6700 (N_6700,N_6321,N_6225);
or U6701 (N_6701,N_6198,N_6268);
or U6702 (N_6702,N_6457,N_6270);
nand U6703 (N_6703,N_6479,N_6244);
nand U6704 (N_6704,N_6287,N_6230);
or U6705 (N_6705,N_6209,N_6442);
xor U6706 (N_6706,N_6053,N_6463);
nor U6707 (N_6707,N_6192,N_6280);
or U6708 (N_6708,N_6404,N_6468);
nand U6709 (N_6709,N_6190,N_6039);
xor U6710 (N_6710,N_6218,N_6004);
nor U6711 (N_6711,N_6118,N_6222);
or U6712 (N_6712,N_6241,N_6006);
and U6713 (N_6713,N_6074,N_6253);
xor U6714 (N_6714,N_6125,N_6453);
and U6715 (N_6715,N_6098,N_6373);
nand U6716 (N_6716,N_6031,N_6339);
or U6717 (N_6717,N_6416,N_6250);
xor U6718 (N_6718,N_6161,N_6359);
or U6719 (N_6719,N_6152,N_6336);
nand U6720 (N_6720,N_6306,N_6216);
xnor U6721 (N_6721,N_6364,N_6392);
nor U6722 (N_6722,N_6210,N_6292);
or U6723 (N_6723,N_6127,N_6124);
or U6724 (N_6724,N_6163,N_6338);
and U6725 (N_6725,N_6159,N_6187);
xnor U6726 (N_6726,N_6259,N_6403);
nor U6727 (N_6727,N_6265,N_6252);
nor U6728 (N_6728,N_6326,N_6008);
and U6729 (N_6729,N_6435,N_6262);
xor U6730 (N_6730,N_6304,N_6096);
nor U6731 (N_6731,N_6238,N_6120);
and U6732 (N_6732,N_6018,N_6301);
nor U6733 (N_6733,N_6412,N_6381);
and U6734 (N_6734,N_6386,N_6235);
nand U6735 (N_6735,N_6450,N_6395);
nor U6736 (N_6736,N_6272,N_6291);
and U6737 (N_6737,N_6429,N_6132);
and U6738 (N_6738,N_6282,N_6300);
or U6739 (N_6739,N_6077,N_6383);
or U6740 (N_6740,N_6382,N_6231);
nor U6741 (N_6741,N_6200,N_6038);
nand U6742 (N_6742,N_6419,N_6337);
nand U6743 (N_6743,N_6446,N_6013);
and U6744 (N_6744,N_6246,N_6322);
xor U6745 (N_6745,N_6153,N_6017);
or U6746 (N_6746,N_6344,N_6276);
xor U6747 (N_6747,N_6356,N_6129);
nand U6748 (N_6748,N_6421,N_6434);
nand U6749 (N_6749,N_6400,N_6366);
nand U6750 (N_6750,N_6351,N_6059);
nand U6751 (N_6751,N_6068,N_6222);
nor U6752 (N_6752,N_6227,N_6013);
xor U6753 (N_6753,N_6354,N_6347);
or U6754 (N_6754,N_6421,N_6181);
or U6755 (N_6755,N_6253,N_6073);
or U6756 (N_6756,N_6291,N_6268);
or U6757 (N_6757,N_6319,N_6190);
nand U6758 (N_6758,N_6182,N_6276);
and U6759 (N_6759,N_6432,N_6079);
nand U6760 (N_6760,N_6428,N_6183);
or U6761 (N_6761,N_6314,N_6230);
or U6762 (N_6762,N_6477,N_6446);
and U6763 (N_6763,N_6365,N_6304);
and U6764 (N_6764,N_6176,N_6251);
or U6765 (N_6765,N_6036,N_6146);
nor U6766 (N_6766,N_6093,N_6452);
or U6767 (N_6767,N_6070,N_6266);
nor U6768 (N_6768,N_6350,N_6017);
xor U6769 (N_6769,N_6201,N_6475);
or U6770 (N_6770,N_6057,N_6390);
nor U6771 (N_6771,N_6240,N_6438);
nand U6772 (N_6772,N_6374,N_6483);
xnor U6773 (N_6773,N_6257,N_6145);
and U6774 (N_6774,N_6015,N_6099);
xor U6775 (N_6775,N_6070,N_6382);
and U6776 (N_6776,N_6366,N_6266);
xor U6777 (N_6777,N_6066,N_6195);
nand U6778 (N_6778,N_6422,N_6014);
or U6779 (N_6779,N_6083,N_6067);
or U6780 (N_6780,N_6342,N_6055);
nand U6781 (N_6781,N_6087,N_6276);
nand U6782 (N_6782,N_6234,N_6420);
and U6783 (N_6783,N_6254,N_6326);
and U6784 (N_6784,N_6423,N_6031);
and U6785 (N_6785,N_6495,N_6055);
nand U6786 (N_6786,N_6367,N_6476);
nor U6787 (N_6787,N_6247,N_6079);
or U6788 (N_6788,N_6182,N_6108);
and U6789 (N_6789,N_6331,N_6073);
nand U6790 (N_6790,N_6208,N_6419);
or U6791 (N_6791,N_6166,N_6432);
nand U6792 (N_6792,N_6183,N_6309);
nor U6793 (N_6793,N_6252,N_6311);
or U6794 (N_6794,N_6275,N_6093);
nor U6795 (N_6795,N_6122,N_6356);
nand U6796 (N_6796,N_6060,N_6474);
or U6797 (N_6797,N_6005,N_6433);
and U6798 (N_6798,N_6296,N_6361);
or U6799 (N_6799,N_6408,N_6292);
or U6800 (N_6800,N_6139,N_6442);
nor U6801 (N_6801,N_6156,N_6385);
xnor U6802 (N_6802,N_6199,N_6072);
and U6803 (N_6803,N_6311,N_6067);
nand U6804 (N_6804,N_6088,N_6011);
or U6805 (N_6805,N_6011,N_6496);
and U6806 (N_6806,N_6202,N_6063);
and U6807 (N_6807,N_6494,N_6482);
or U6808 (N_6808,N_6395,N_6435);
nor U6809 (N_6809,N_6004,N_6158);
xnor U6810 (N_6810,N_6128,N_6283);
nand U6811 (N_6811,N_6237,N_6383);
nand U6812 (N_6812,N_6204,N_6200);
nor U6813 (N_6813,N_6115,N_6064);
and U6814 (N_6814,N_6025,N_6406);
and U6815 (N_6815,N_6443,N_6196);
and U6816 (N_6816,N_6023,N_6126);
nor U6817 (N_6817,N_6251,N_6459);
nor U6818 (N_6818,N_6034,N_6471);
nor U6819 (N_6819,N_6223,N_6254);
and U6820 (N_6820,N_6286,N_6468);
nand U6821 (N_6821,N_6016,N_6253);
or U6822 (N_6822,N_6131,N_6328);
xor U6823 (N_6823,N_6387,N_6239);
nand U6824 (N_6824,N_6085,N_6114);
nor U6825 (N_6825,N_6246,N_6015);
xnor U6826 (N_6826,N_6295,N_6268);
and U6827 (N_6827,N_6037,N_6310);
nor U6828 (N_6828,N_6087,N_6157);
and U6829 (N_6829,N_6156,N_6155);
xor U6830 (N_6830,N_6337,N_6331);
nor U6831 (N_6831,N_6263,N_6185);
or U6832 (N_6832,N_6401,N_6256);
xor U6833 (N_6833,N_6135,N_6291);
and U6834 (N_6834,N_6398,N_6157);
nand U6835 (N_6835,N_6365,N_6157);
nand U6836 (N_6836,N_6479,N_6093);
xor U6837 (N_6837,N_6385,N_6322);
nand U6838 (N_6838,N_6432,N_6126);
xor U6839 (N_6839,N_6391,N_6085);
xnor U6840 (N_6840,N_6498,N_6183);
nand U6841 (N_6841,N_6185,N_6239);
xnor U6842 (N_6842,N_6034,N_6276);
nand U6843 (N_6843,N_6240,N_6383);
or U6844 (N_6844,N_6206,N_6351);
nor U6845 (N_6845,N_6047,N_6248);
xnor U6846 (N_6846,N_6093,N_6475);
or U6847 (N_6847,N_6493,N_6482);
nor U6848 (N_6848,N_6277,N_6116);
and U6849 (N_6849,N_6491,N_6480);
nand U6850 (N_6850,N_6415,N_6180);
and U6851 (N_6851,N_6345,N_6048);
or U6852 (N_6852,N_6034,N_6312);
xnor U6853 (N_6853,N_6226,N_6204);
nor U6854 (N_6854,N_6060,N_6281);
and U6855 (N_6855,N_6016,N_6382);
nor U6856 (N_6856,N_6291,N_6391);
and U6857 (N_6857,N_6138,N_6140);
nand U6858 (N_6858,N_6116,N_6260);
nor U6859 (N_6859,N_6410,N_6114);
xnor U6860 (N_6860,N_6453,N_6296);
nor U6861 (N_6861,N_6151,N_6158);
nand U6862 (N_6862,N_6054,N_6276);
and U6863 (N_6863,N_6114,N_6038);
and U6864 (N_6864,N_6089,N_6117);
or U6865 (N_6865,N_6042,N_6376);
and U6866 (N_6866,N_6234,N_6236);
nand U6867 (N_6867,N_6380,N_6492);
and U6868 (N_6868,N_6054,N_6466);
nor U6869 (N_6869,N_6263,N_6363);
nor U6870 (N_6870,N_6404,N_6259);
or U6871 (N_6871,N_6428,N_6128);
or U6872 (N_6872,N_6001,N_6286);
xor U6873 (N_6873,N_6091,N_6100);
xor U6874 (N_6874,N_6157,N_6020);
nor U6875 (N_6875,N_6261,N_6447);
or U6876 (N_6876,N_6180,N_6023);
xnor U6877 (N_6877,N_6171,N_6262);
nand U6878 (N_6878,N_6287,N_6090);
or U6879 (N_6879,N_6364,N_6321);
and U6880 (N_6880,N_6084,N_6105);
nand U6881 (N_6881,N_6343,N_6085);
xor U6882 (N_6882,N_6371,N_6477);
and U6883 (N_6883,N_6278,N_6240);
nand U6884 (N_6884,N_6259,N_6489);
xnor U6885 (N_6885,N_6303,N_6154);
or U6886 (N_6886,N_6065,N_6384);
nand U6887 (N_6887,N_6483,N_6207);
nand U6888 (N_6888,N_6154,N_6159);
and U6889 (N_6889,N_6227,N_6446);
and U6890 (N_6890,N_6101,N_6453);
and U6891 (N_6891,N_6118,N_6315);
nand U6892 (N_6892,N_6348,N_6246);
nand U6893 (N_6893,N_6259,N_6048);
or U6894 (N_6894,N_6316,N_6322);
nand U6895 (N_6895,N_6449,N_6346);
and U6896 (N_6896,N_6135,N_6067);
nand U6897 (N_6897,N_6459,N_6384);
xor U6898 (N_6898,N_6178,N_6044);
xnor U6899 (N_6899,N_6223,N_6494);
nand U6900 (N_6900,N_6441,N_6076);
or U6901 (N_6901,N_6358,N_6113);
and U6902 (N_6902,N_6099,N_6349);
xnor U6903 (N_6903,N_6273,N_6102);
xor U6904 (N_6904,N_6187,N_6367);
nand U6905 (N_6905,N_6127,N_6307);
xor U6906 (N_6906,N_6001,N_6484);
or U6907 (N_6907,N_6348,N_6498);
xnor U6908 (N_6908,N_6018,N_6225);
nand U6909 (N_6909,N_6251,N_6047);
and U6910 (N_6910,N_6116,N_6436);
nand U6911 (N_6911,N_6056,N_6365);
nand U6912 (N_6912,N_6190,N_6246);
nor U6913 (N_6913,N_6279,N_6186);
nor U6914 (N_6914,N_6292,N_6180);
and U6915 (N_6915,N_6319,N_6432);
xor U6916 (N_6916,N_6493,N_6276);
and U6917 (N_6917,N_6291,N_6352);
nor U6918 (N_6918,N_6152,N_6192);
or U6919 (N_6919,N_6376,N_6498);
or U6920 (N_6920,N_6033,N_6212);
xnor U6921 (N_6921,N_6044,N_6004);
or U6922 (N_6922,N_6228,N_6306);
nand U6923 (N_6923,N_6201,N_6467);
nand U6924 (N_6924,N_6123,N_6005);
nor U6925 (N_6925,N_6050,N_6374);
and U6926 (N_6926,N_6365,N_6246);
nand U6927 (N_6927,N_6388,N_6167);
or U6928 (N_6928,N_6353,N_6024);
nand U6929 (N_6929,N_6182,N_6424);
or U6930 (N_6930,N_6325,N_6285);
or U6931 (N_6931,N_6413,N_6160);
xnor U6932 (N_6932,N_6086,N_6026);
and U6933 (N_6933,N_6108,N_6397);
nor U6934 (N_6934,N_6186,N_6100);
nor U6935 (N_6935,N_6069,N_6494);
xnor U6936 (N_6936,N_6266,N_6115);
and U6937 (N_6937,N_6384,N_6225);
and U6938 (N_6938,N_6228,N_6081);
nand U6939 (N_6939,N_6492,N_6394);
xnor U6940 (N_6940,N_6341,N_6041);
nor U6941 (N_6941,N_6213,N_6416);
xnor U6942 (N_6942,N_6210,N_6053);
nor U6943 (N_6943,N_6034,N_6065);
xor U6944 (N_6944,N_6086,N_6478);
or U6945 (N_6945,N_6262,N_6127);
xor U6946 (N_6946,N_6391,N_6463);
nand U6947 (N_6947,N_6493,N_6090);
nand U6948 (N_6948,N_6014,N_6137);
xnor U6949 (N_6949,N_6107,N_6054);
nand U6950 (N_6950,N_6481,N_6088);
nand U6951 (N_6951,N_6250,N_6484);
nor U6952 (N_6952,N_6050,N_6213);
and U6953 (N_6953,N_6481,N_6438);
nand U6954 (N_6954,N_6316,N_6487);
xnor U6955 (N_6955,N_6492,N_6162);
or U6956 (N_6956,N_6148,N_6452);
and U6957 (N_6957,N_6143,N_6283);
xnor U6958 (N_6958,N_6226,N_6020);
and U6959 (N_6959,N_6166,N_6408);
and U6960 (N_6960,N_6102,N_6130);
or U6961 (N_6961,N_6372,N_6201);
nand U6962 (N_6962,N_6141,N_6355);
nor U6963 (N_6963,N_6007,N_6326);
nor U6964 (N_6964,N_6221,N_6227);
xor U6965 (N_6965,N_6038,N_6327);
and U6966 (N_6966,N_6017,N_6060);
xnor U6967 (N_6967,N_6391,N_6371);
xor U6968 (N_6968,N_6376,N_6184);
xor U6969 (N_6969,N_6080,N_6176);
nor U6970 (N_6970,N_6155,N_6043);
or U6971 (N_6971,N_6218,N_6344);
and U6972 (N_6972,N_6156,N_6208);
nor U6973 (N_6973,N_6198,N_6105);
nand U6974 (N_6974,N_6226,N_6200);
nor U6975 (N_6975,N_6214,N_6419);
nor U6976 (N_6976,N_6431,N_6471);
or U6977 (N_6977,N_6380,N_6371);
nand U6978 (N_6978,N_6431,N_6481);
xor U6979 (N_6979,N_6446,N_6358);
xor U6980 (N_6980,N_6032,N_6242);
xor U6981 (N_6981,N_6135,N_6484);
nor U6982 (N_6982,N_6291,N_6486);
or U6983 (N_6983,N_6120,N_6171);
nor U6984 (N_6984,N_6033,N_6498);
nand U6985 (N_6985,N_6263,N_6101);
nor U6986 (N_6986,N_6150,N_6323);
nor U6987 (N_6987,N_6134,N_6139);
or U6988 (N_6988,N_6243,N_6104);
and U6989 (N_6989,N_6232,N_6181);
nand U6990 (N_6990,N_6152,N_6469);
nor U6991 (N_6991,N_6179,N_6163);
xor U6992 (N_6992,N_6265,N_6314);
xnor U6993 (N_6993,N_6167,N_6312);
or U6994 (N_6994,N_6136,N_6198);
xor U6995 (N_6995,N_6276,N_6302);
and U6996 (N_6996,N_6059,N_6131);
xor U6997 (N_6997,N_6479,N_6450);
nor U6998 (N_6998,N_6129,N_6205);
nor U6999 (N_6999,N_6122,N_6437);
xnor U7000 (N_7000,N_6687,N_6922);
xnor U7001 (N_7001,N_6958,N_6898);
xor U7002 (N_7002,N_6528,N_6733);
xnor U7003 (N_7003,N_6559,N_6682);
or U7004 (N_7004,N_6547,N_6765);
nor U7005 (N_7005,N_6673,N_6757);
nor U7006 (N_7006,N_6943,N_6589);
nor U7007 (N_7007,N_6884,N_6758);
nand U7008 (N_7008,N_6883,N_6523);
nor U7009 (N_7009,N_6726,N_6764);
nor U7010 (N_7010,N_6507,N_6852);
or U7011 (N_7011,N_6580,N_6778);
xnor U7012 (N_7012,N_6761,N_6524);
or U7013 (N_7013,N_6644,N_6667);
xnor U7014 (N_7014,N_6745,N_6739);
xnor U7015 (N_7015,N_6796,N_6754);
and U7016 (N_7016,N_6822,N_6649);
nand U7017 (N_7017,N_6808,N_6723);
and U7018 (N_7018,N_6521,N_6517);
or U7019 (N_7019,N_6707,N_6620);
or U7020 (N_7020,N_6813,N_6776);
and U7021 (N_7021,N_6818,N_6593);
or U7022 (N_7022,N_6692,N_6640);
nand U7023 (N_7023,N_6970,N_6738);
nor U7024 (N_7024,N_6914,N_6994);
and U7025 (N_7025,N_6828,N_6982);
xnor U7026 (N_7026,N_6749,N_6552);
or U7027 (N_7027,N_6718,N_6572);
and U7028 (N_7028,N_6956,N_6777);
or U7029 (N_7029,N_6939,N_6964);
or U7030 (N_7030,N_6954,N_6836);
or U7031 (N_7031,N_6872,N_6621);
or U7032 (N_7032,N_6693,N_6591);
and U7033 (N_7033,N_6999,N_6503);
or U7034 (N_7034,N_6961,N_6587);
nor U7035 (N_7035,N_6633,N_6569);
or U7036 (N_7036,N_6893,N_6830);
nor U7037 (N_7037,N_6769,N_6965);
and U7038 (N_7038,N_6990,N_6535);
nand U7039 (N_7039,N_6751,N_6696);
nor U7040 (N_7040,N_6741,N_6955);
or U7041 (N_7041,N_6534,N_6960);
and U7042 (N_7042,N_6558,N_6564);
or U7043 (N_7043,N_6937,N_6923);
nor U7044 (N_7044,N_6537,N_6968);
nand U7045 (N_7045,N_6632,N_6921);
or U7046 (N_7046,N_6689,N_6936);
or U7047 (N_7047,N_6695,N_6832);
nor U7048 (N_7048,N_6785,N_6529);
and U7049 (N_7049,N_6721,N_6834);
or U7050 (N_7050,N_6942,N_6973);
nor U7051 (N_7051,N_6816,N_6715);
and U7052 (N_7052,N_6952,N_6634);
and U7053 (N_7053,N_6806,N_6779);
and U7054 (N_7054,N_6815,N_6799);
xnor U7055 (N_7055,N_6599,N_6677);
and U7056 (N_7056,N_6853,N_6859);
or U7057 (N_7057,N_6878,N_6623);
nand U7058 (N_7058,N_6594,N_6807);
nand U7059 (N_7059,N_6541,N_6561);
nor U7060 (N_7060,N_6533,N_6501);
and U7061 (N_7061,N_6981,N_6639);
xor U7062 (N_7062,N_6905,N_6658);
nor U7063 (N_7063,N_6752,N_6582);
xnor U7064 (N_7064,N_6906,N_6988);
xnor U7065 (N_7065,N_6946,N_6877);
and U7066 (N_7066,N_6676,N_6895);
or U7067 (N_7067,N_6728,N_6825);
and U7068 (N_7068,N_6505,N_6803);
and U7069 (N_7069,N_6911,N_6920);
nor U7070 (N_7070,N_6710,N_6903);
or U7071 (N_7071,N_6890,N_6879);
xor U7072 (N_7072,N_6628,N_6606);
and U7073 (N_7073,N_6627,N_6930);
or U7074 (N_7074,N_6550,N_6910);
and U7075 (N_7075,N_6519,N_6694);
or U7076 (N_7076,N_6588,N_6876);
xor U7077 (N_7077,N_6917,N_6536);
nor U7078 (N_7078,N_6838,N_6743);
xor U7079 (N_7079,N_6983,N_6735);
nand U7080 (N_7080,N_6951,N_6858);
or U7081 (N_7081,N_6656,N_6849);
nor U7082 (N_7082,N_6788,N_6899);
and U7083 (N_7083,N_6887,N_6985);
nor U7084 (N_7084,N_6657,N_6748);
nand U7085 (N_7085,N_6763,N_6925);
xnor U7086 (N_7086,N_6556,N_6753);
nor U7087 (N_7087,N_6842,N_6902);
nor U7088 (N_7088,N_6913,N_6708);
and U7089 (N_7089,N_6618,N_6542);
or U7090 (N_7090,N_6648,N_6548);
or U7091 (N_7091,N_6671,N_6881);
xnor U7092 (N_7092,N_6768,N_6868);
and U7093 (N_7093,N_6518,N_6549);
xnor U7094 (N_7094,N_6650,N_6613);
xnor U7095 (N_7095,N_6714,N_6719);
and U7096 (N_7096,N_6947,N_6509);
nand U7097 (N_7097,N_6844,N_6989);
and U7098 (N_7098,N_6575,N_6651);
nor U7099 (N_7099,N_6576,N_6997);
and U7100 (N_7100,N_6678,N_6551);
nand U7101 (N_7101,N_6790,N_6516);
nand U7102 (N_7102,N_6510,N_6670);
or U7103 (N_7103,N_6848,N_6630);
or U7104 (N_7104,N_6760,N_6854);
nand U7105 (N_7105,N_6686,N_6767);
nand U7106 (N_7106,N_6713,N_6531);
or U7107 (N_7107,N_6861,N_6938);
and U7108 (N_7108,N_6798,N_6756);
nor U7109 (N_7109,N_6809,N_6864);
and U7110 (N_7110,N_6904,N_6579);
xor U7111 (N_7111,N_6929,N_6941);
xnor U7112 (N_7112,N_6730,N_6664);
xnor U7113 (N_7113,N_6571,N_6619);
nand U7114 (N_7114,N_6993,N_6794);
nor U7115 (N_7115,N_6833,N_6775);
nand U7116 (N_7116,N_6638,N_6646);
and U7117 (N_7117,N_6966,N_6601);
xnor U7118 (N_7118,N_6722,N_6625);
nor U7119 (N_7119,N_6544,N_6998);
or U7120 (N_7120,N_6892,N_6986);
nand U7121 (N_7121,N_6637,N_6894);
and U7122 (N_7122,N_6885,N_6538);
xor U7123 (N_7123,N_6962,N_6725);
or U7124 (N_7124,N_6847,N_6802);
xor U7125 (N_7125,N_6814,N_6782);
or U7126 (N_7126,N_6927,N_6605);
nor U7127 (N_7127,N_6786,N_6978);
xnor U7128 (N_7128,N_6597,N_6540);
or U7129 (N_7129,N_6980,N_6774);
xnor U7130 (N_7130,N_6916,N_6724);
nand U7131 (N_7131,N_6963,N_6700);
nor U7132 (N_7132,N_6685,N_6856);
nor U7133 (N_7133,N_6669,N_6697);
xor U7134 (N_7134,N_6731,N_6539);
nor U7135 (N_7135,N_6635,N_6585);
or U7136 (N_7136,N_6846,N_6959);
or U7137 (N_7137,N_6869,N_6975);
or U7138 (N_7138,N_6543,N_6727);
or U7139 (N_7139,N_6683,N_6530);
nor U7140 (N_7140,N_6555,N_6770);
and U7141 (N_7141,N_6690,N_6957);
and U7142 (N_7142,N_6795,N_6643);
or U7143 (N_7143,N_6566,N_6821);
nand U7144 (N_7144,N_6565,N_6502);
nand U7145 (N_7145,N_6850,N_6866);
xnor U7146 (N_7146,N_6609,N_6520);
xnor U7147 (N_7147,N_6652,N_6631);
nor U7148 (N_7148,N_6860,N_6712);
nand U7149 (N_7149,N_6773,N_6679);
nand U7150 (N_7150,N_6840,N_6616);
xor U7151 (N_7151,N_6950,N_6826);
xor U7152 (N_7152,N_6734,N_6800);
or U7153 (N_7153,N_6532,N_6611);
xnor U7154 (N_7154,N_6668,N_6573);
nor U7155 (N_7155,N_6949,N_6839);
and U7156 (N_7156,N_6655,N_6602);
or U7157 (N_7157,N_6789,N_6805);
xnor U7158 (N_7158,N_6772,N_6940);
and U7159 (N_7159,N_6513,N_6971);
xor U7160 (N_7160,N_6875,N_6680);
and U7161 (N_7161,N_6598,N_6600);
nand U7162 (N_7162,N_6603,N_6545);
or U7163 (N_7163,N_6992,N_6912);
nand U7164 (N_7164,N_6684,N_6653);
nand U7165 (N_7165,N_6604,N_6873);
nor U7166 (N_7166,N_6546,N_6703);
and U7167 (N_7167,N_6608,N_6515);
nor U7168 (N_7168,N_6865,N_6900);
or U7169 (N_7169,N_6934,N_6863);
and U7170 (N_7170,N_6500,N_6918);
nand U7171 (N_7171,N_6557,N_6793);
and U7172 (N_7172,N_6976,N_6924);
and U7173 (N_7173,N_6701,N_6972);
and U7174 (N_7174,N_6706,N_6750);
nor U7175 (N_7175,N_6874,N_6504);
xor U7176 (N_7176,N_6811,N_6666);
xor U7177 (N_7177,N_6967,N_6596);
nor U7178 (N_7178,N_6953,N_6583);
xor U7179 (N_7179,N_6996,N_6584);
nand U7180 (N_7180,N_6662,N_6762);
xnor U7181 (N_7181,N_6674,N_6527);
xor U7182 (N_7182,N_6919,N_6736);
xor U7183 (N_7183,N_6979,N_6506);
xnor U7184 (N_7184,N_6792,N_6897);
nor U7185 (N_7185,N_6823,N_6948);
xnor U7186 (N_7186,N_6974,N_6699);
nand U7187 (N_7187,N_6665,N_6737);
nand U7188 (N_7188,N_6562,N_6636);
xor U7189 (N_7189,N_6553,N_6780);
and U7190 (N_7190,N_6812,N_6817);
nor U7191 (N_7191,N_6931,N_6801);
nor U7192 (N_7192,N_6675,N_6622);
xnor U7193 (N_7193,N_6717,N_6791);
nand U7194 (N_7194,N_6862,N_6574);
and U7195 (N_7195,N_6581,N_6827);
xnor U7196 (N_7196,N_6577,N_6935);
nand U7197 (N_7197,N_6784,N_6889);
xnor U7198 (N_7198,N_6716,N_6732);
nor U7199 (N_7199,N_6511,N_6568);
nand U7200 (N_7200,N_6804,N_6567);
and U7201 (N_7201,N_6888,N_6831);
nand U7202 (N_7202,N_6659,N_6871);
xor U7203 (N_7203,N_6755,N_6698);
xor U7204 (N_7204,N_6570,N_6661);
or U7205 (N_7205,N_6945,N_6720);
and U7206 (N_7206,N_6578,N_6820);
xnor U7207 (N_7207,N_6514,N_6907);
nand U7208 (N_7208,N_6554,N_6704);
xor U7209 (N_7209,N_6508,N_6691);
xor U7210 (N_7210,N_6891,N_6740);
and U7211 (N_7211,N_6746,N_6641);
or U7212 (N_7212,N_6642,N_6909);
xnor U7213 (N_7213,N_6747,N_6742);
or U7214 (N_7214,N_6969,N_6995);
or U7215 (N_7215,N_6928,N_6522);
nor U7216 (N_7216,N_6926,N_6586);
nor U7217 (N_7217,N_6851,N_6629);
and U7218 (N_7218,N_6835,N_6824);
nor U7219 (N_7219,N_6612,N_6595);
nor U7220 (N_7220,N_6592,N_6787);
nand U7221 (N_7221,N_6645,N_6660);
or U7222 (N_7222,N_6915,N_6819);
nor U7223 (N_7223,N_6702,N_6560);
or U7224 (N_7224,N_6843,N_6781);
nand U7225 (N_7225,N_6624,N_6797);
or U7226 (N_7226,N_6563,N_6896);
nand U7227 (N_7227,N_6810,N_6759);
xnor U7228 (N_7228,N_6855,N_6837);
xnor U7229 (N_7229,N_6709,N_6615);
nor U7230 (N_7230,N_6729,N_6705);
nor U7231 (N_7231,N_6783,N_6525);
and U7232 (N_7232,N_6590,N_6744);
nand U7233 (N_7233,N_6617,N_6841);
xnor U7234 (N_7234,N_6607,N_6688);
nor U7235 (N_7235,N_6610,N_6857);
nor U7236 (N_7236,N_6614,N_6829);
and U7237 (N_7237,N_6880,N_6987);
or U7238 (N_7238,N_6672,N_6626);
nand U7239 (N_7239,N_6932,N_6882);
or U7240 (N_7240,N_6886,N_6654);
and U7241 (N_7241,N_6681,N_6991);
and U7242 (N_7242,N_6867,N_6977);
nor U7243 (N_7243,N_6771,N_6663);
nand U7244 (N_7244,N_6908,N_6984);
nor U7245 (N_7245,N_6944,N_6933);
nand U7246 (N_7246,N_6647,N_6711);
xnor U7247 (N_7247,N_6526,N_6870);
or U7248 (N_7248,N_6766,N_6845);
nor U7249 (N_7249,N_6512,N_6901);
and U7250 (N_7250,N_6623,N_6626);
and U7251 (N_7251,N_6935,N_6716);
nand U7252 (N_7252,N_6899,N_6698);
xor U7253 (N_7253,N_6863,N_6986);
nor U7254 (N_7254,N_6798,N_6831);
and U7255 (N_7255,N_6634,N_6696);
xor U7256 (N_7256,N_6824,N_6753);
or U7257 (N_7257,N_6521,N_6596);
and U7258 (N_7258,N_6751,N_6951);
or U7259 (N_7259,N_6649,N_6996);
nor U7260 (N_7260,N_6790,N_6895);
nor U7261 (N_7261,N_6747,N_6823);
or U7262 (N_7262,N_6698,N_6706);
nand U7263 (N_7263,N_6739,N_6591);
and U7264 (N_7264,N_6767,N_6985);
or U7265 (N_7265,N_6607,N_6997);
or U7266 (N_7266,N_6675,N_6583);
nand U7267 (N_7267,N_6526,N_6820);
nor U7268 (N_7268,N_6679,N_6961);
xor U7269 (N_7269,N_6927,N_6731);
and U7270 (N_7270,N_6984,N_6588);
nor U7271 (N_7271,N_6894,N_6728);
nand U7272 (N_7272,N_6718,N_6923);
nand U7273 (N_7273,N_6572,N_6746);
and U7274 (N_7274,N_6853,N_6625);
nand U7275 (N_7275,N_6931,N_6703);
xnor U7276 (N_7276,N_6747,N_6793);
nand U7277 (N_7277,N_6996,N_6967);
xnor U7278 (N_7278,N_6969,N_6601);
nand U7279 (N_7279,N_6830,N_6819);
nor U7280 (N_7280,N_6716,N_6811);
and U7281 (N_7281,N_6702,N_6718);
nand U7282 (N_7282,N_6769,N_6730);
nand U7283 (N_7283,N_6847,N_6681);
or U7284 (N_7284,N_6557,N_6823);
xor U7285 (N_7285,N_6513,N_6502);
nor U7286 (N_7286,N_6808,N_6947);
nand U7287 (N_7287,N_6677,N_6666);
or U7288 (N_7288,N_6693,N_6694);
or U7289 (N_7289,N_6874,N_6765);
nor U7290 (N_7290,N_6599,N_6800);
and U7291 (N_7291,N_6793,N_6977);
nand U7292 (N_7292,N_6579,N_6531);
nand U7293 (N_7293,N_6785,N_6853);
or U7294 (N_7294,N_6657,N_6519);
or U7295 (N_7295,N_6619,N_6544);
or U7296 (N_7296,N_6860,N_6533);
and U7297 (N_7297,N_6630,N_6556);
or U7298 (N_7298,N_6772,N_6828);
nand U7299 (N_7299,N_6750,N_6878);
nor U7300 (N_7300,N_6821,N_6841);
xor U7301 (N_7301,N_6681,N_6820);
and U7302 (N_7302,N_6807,N_6649);
xnor U7303 (N_7303,N_6540,N_6671);
or U7304 (N_7304,N_6775,N_6807);
or U7305 (N_7305,N_6912,N_6701);
nor U7306 (N_7306,N_6578,N_6880);
nor U7307 (N_7307,N_6875,N_6621);
and U7308 (N_7308,N_6972,N_6567);
and U7309 (N_7309,N_6918,N_6846);
xor U7310 (N_7310,N_6917,N_6957);
nor U7311 (N_7311,N_6907,N_6593);
xnor U7312 (N_7312,N_6790,N_6553);
nand U7313 (N_7313,N_6976,N_6934);
xor U7314 (N_7314,N_6506,N_6556);
and U7315 (N_7315,N_6855,N_6819);
nand U7316 (N_7316,N_6954,N_6833);
nor U7317 (N_7317,N_6506,N_6693);
xor U7318 (N_7318,N_6506,N_6691);
and U7319 (N_7319,N_6659,N_6796);
nor U7320 (N_7320,N_6997,N_6541);
nand U7321 (N_7321,N_6867,N_6834);
or U7322 (N_7322,N_6643,N_6984);
nor U7323 (N_7323,N_6629,N_6974);
and U7324 (N_7324,N_6576,N_6569);
or U7325 (N_7325,N_6676,N_6752);
or U7326 (N_7326,N_6599,N_6522);
and U7327 (N_7327,N_6738,N_6888);
nand U7328 (N_7328,N_6865,N_6964);
nor U7329 (N_7329,N_6765,N_6761);
xor U7330 (N_7330,N_6879,N_6850);
nand U7331 (N_7331,N_6562,N_6643);
or U7332 (N_7332,N_6696,N_6707);
nand U7333 (N_7333,N_6693,N_6839);
nor U7334 (N_7334,N_6867,N_6502);
or U7335 (N_7335,N_6991,N_6709);
nor U7336 (N_7336,N_6631,N_6788);
nand U7337 (N_7337,N_6730,N_6993);
nand U7338 (N_7338,N_6994,N_6962);
nor U7339 (N_7339,N_6775,N_6926);
nand U7340 (N_7340,N_6725,N_6521);
xor U7341 (N_7341,N_6850,N_6568);
nor U7342 (N_7342,N_6506,N_6938);
and U7343 (N_7343,N_6520,N_6894);
xnor U7344 (N_7344,N_6998,N_6523);
and U7345 (N_7345,N_6926,N_6529);
and U7346 (N_7346,N_6802,N_6771);
xnor U7347 (N_7347,N_6664,N_6774);
nor U7348 (N_7348,N_6821,N_6742);
nand U7349 (N_7349,N_6880,N_6512);
and U7350 (N_7350,N_6883,N_6754);
xor U7351 (N_7351,N_6986,N_6741);
nor U7352 (N_7352,N_6795,N_6719);
nand U7353 (N_7353,N_6993,N_6532);
xnor U7354 (N_7354,N_6693,N_6620);
or U7355 (N_7355,N_6941,N_6851);
xnor U7356 (N_7356,N_6586,N_6619);
nand U7357 (N_7357,N_6698,N_6536);
nor U7358 (N_7358,N_6959,N_6833);
nand U7359 (N_7359,N_6835,N_6707);
nor U7360 (N_7360,N_6746,N_6846);
nand U7361 (N_7361,N_6585,N_6957);
nor U7362 (N_7362,N_6737,N_6803);
nand U7363 (N_7363,N_6895,N_6767);
nand U7364 (N_7364,N_6608,N_6924);
nor U7365 (N_7365,N_6673,N_6683);
xnor U7366 (N_7366,N_6549,N_6753);
and U7367 (N_7367,N_6529,N_6911);
nor U7368 (N_7368,N_6674,N_6954);
nand U7369 (N_7369,N_6582,N_6543);
xnor U7370 (N_7370,N_6670,N_6760);
and U7371 (N_7371,N_6947,N_6904);
nor U7372 (N_7372,N_6686,N_6734);
and U7373 (N_7373,N_6686,N_6530);
nand U7374 (N_7374,N_6509,N_6933);
xor U7375 (N_7375,N_6986,N_6645);
and U7376 (N_7376,N_6774,N_6992);
nand U7377 (N_7377,N_6917,N_6937);
nor U7378 (N_7378,N_6987,N_6740);
and U7379 (N_7379,N_6548,N_6970);
xor U7380 (N_7380,N_6691,N_6874);
and U7381 (N_7381,N_6530,N_6732);
nor U7382 (N_7382,N_6665,N_6655);
nand U7383 (N_7383,N_6531,N_6971);
nor U7384 (N_7384,N_6509,N_6953);
or U7385 (N_7385,N_6590,N_6756);
xor U7386 (N_7386,N_6872,N_6531);
nand U7387 (N_7387,N_6815,N_6741);
xnor U7388 (N_7388,N_6831,N_6803);
nor U7389 (N_7389,N_6635,N_6696);
nand U7390 (N_7390,N_6807,N_6692);
or U7391 (N_7391,N_6924,N_6739);
or U7392 (N_7392,N_6802,N_6628);
nor U7393 (N_7393,N_6942,N_6931);
nand U7394 (N_7394,N_6879,N_6874);
nand U7395 (N_7395,N_6809,N_6673);
and U7396 (N_7396,N_6626,N_6612);
nor U7397 (N_7397,N_6542,N_6820);
nand U7398 (N_7398,N_6913,N_6957);
nor U7399 (N_7399,N_6838,N_6727);
nor U7400 (N_7400,N_6711,N_6580);
nor U7401 (N_7401,N_6848,N_6911);
or U7402 (N_7402,N_6545,N_6975);
or U7403 (N_7403,N_6978,N_6971);
nand U7404 (N_7404,N_6866,N_6787);
or U7405 (N_7405,N_6772,N_6707);
xor U7406 (N_7406,N_6505,N_6869);
nor U7407 (N_7407,N_6614,N_6740);
nor U7408 (N_7408,N_6610,N_6938);
nand U7409 (N_7409,N_6658,N_6647);
xnor U7410 (N_7410,N_6979,N_6950);
nand U7411 (N_7411,N_6643,N_6671);
and U7412 (N_7412,N_6696,N_6725);
xor U7413 (N_7413,N_6948,N_6822);
xor U7414 (N_7414,N_6843,N_6818);
and U7415 (N_7415,N_6624,N_6783);
or U7416 (N_7416,N_6528,N_6820);
and U7417 (N_7417,N_6740,N_6536);
nor U7418 (N_7418,N_6627,N_6644);
nand U7419 (N_7419,N_6664,N_6644);
and U7420 (N_7420,N_6730,N_6719);
nand U7421 (N_7421,N_6992,N_6539);
nor U7422 (N_7422,N_6948,N_6583);
and U7423 (N_7423,N_6883,N_6503);
xor U7424 (N_7424,N_6812,N_6990);
and U7425 (N_7425,N_6632,N_6604);
xnor U7426 (N_7426,N_6737,N_6950);
nor U7427 (N_7427,N_6731,N_6999);
nand U7428 (N_7428,N_6831,N_6675);
nand U7429 (N_7429,N_6993,N_6641);
nor U7430 (N_7430,N_6793,N_6552);
xor U7431 (N_7431,N_6908,N_6501);
nor U7432 (N_7432,N_6671,N_6523);
xor U7433 (N_7433,N_6551,N_6535);
nor U7434 (N_7434,N_6619,N_6718);
or U7435 (N_7435,N_6830,N_6800);
nor U7436 (N_7436,N_6810,N_6859);
xnor U7437 (N_7437,N_6811,N_6796);
and U7438 (N_7438,N_6743,N_6624);
and U7439 (N_7439,N_6716,N_6844);
and U7440 (N_7440,N_6524,N_6784);
or U7441 (N_7441,N_6832,N_6760);
or U7442 (N_7442,N_6538,N_6661);
or U7443 (N_7443,N_6907,N_6729);
nor U7444 (N_7444,N_6631,N_6980);
xnor U7445 (N_7445,N_6660,N_6575);
nand U7446 (N_7446,N_6586,N_6863);
and U7447 (N_7447,N_6797,N_6510);
xor U7448 (N_7448,N_6681,N_6636);
and U7449 (N_7449,N_6534,N_6723);
and U7450 (N_7450,N_6517,N_6609);
or U7451 (N_7451,N_6819,N_6536);
nand U7452 (N_7452,N_6871,N_6758);
xnor U7453 (N_7453,N_6570,N_6644);
nor U7454 (N_7454,N_6804,N_6849);
or U7455 (N_7455,N_6720,N_6851);
xor U7456 (N_7456,N_6555,N_6549);
nand U7457 (N_7457,N_6630,N_6853);
or U7458 (N_7458,N_6590,N_6587);
and U7459 (N_7459,N_6769,N_6867);
nor U7460 (N_7460,N_6697,N_6525);
xnor U7461 (N_7461,N_6662,N_6607);
and U7462 (N_7462,N_6732,N_6714);
nor U7463 (N_7463,N_6699,N_6646);
xor U7464 (N_7464,N_6885,N_6686);
xnor U7465 (N_7465,N_6585,N_6678);
xnor U7466 (N_7466,N_6887,N_6923);
or U7467 (N_7467,N_6806,N_6591);
nor U7468 (N_7468,N_6625,N_6973);
xor U7469 (N_7469,N_6553,N_6670);
nor U7470 (N_7470,N_6740,N_6617);
nor U7471 (N_7471,N_6640,N_6891);
nand U7472 (N_7472,N_6903,N_6500);
xnor U7473 (N_7473,N_6693,N_6827);
or U7474 (N_7474,N_6584,N_6766);
nor U7475 (N_7475,N_6789,N_6950);
nand U7476 (N_7476,N_6754,N_6555);
and U7477 (N_7477,N_6604,N_6816);
nor U7478 (N_7478,N_6501,N_6665);
nor U7479 (N_7479,N_6849,N_6607);
and U7480 (N_7480,N_6590,N_6581);
or U7481 (N_7481,N_6688,N_6734);
nand U7482 (N_7482,N_6848,N_6855);
xnor U7483 (N_7483,N_6743,N_6540);
or U7484 (N_7484,N_6550,N_6549);
nor U7485 (N_7485,N_6552,N_6520);
nor U7486 (N_7486,N_6739,N_6746);
or U7487 (N_7487,N_6917,N_6828);
nor U7488 (N_7488,N_6715,N_6896);
nand U7489 (N_7489,N_6819,N_6965);
and U7490 (N_7490,N_6978,N_6581);
and U7491 (N_7491,N_6970,N_6891);
nand U7492 (N_7492,N_6999,N_6929);
or U7493 (N_7493,N_6811,N_6812);
or U7494 (N_7494,N_6973,N_6999);
nand U7495 (N_7495,N_6804,N_6816);
nand U7496 (N_7496,N_6581,N_6896);
or U7497 (N_7497,N_6801,N_6860);
nor U7498 (N_7498,N_6829,N_6776);
and U7499 (N_7499,N_6695,N_6651);
and U7500 (N_7500,N_7444,N_7428);
or U7501 (N_7501,N_7049,N_7301);
and U7502 (N_7502,N_7284,N_7405);
xor U7503 (N_7503,N_7144,N_7384);
xnor U7504 (N_7504,N_7246,N_7108);
and U7505 (N_7505,N_7421,N_7309);
nand U7506 (N_7506,N_7299,N_7475);
and U7507 (N_7507,N_7400,N_7230);
xnor U7508 (N_7508,N_7035,N_7157);
xnor U7509 (N_7509,N_7149,N_7419);
xor U7510 (N_7510,N_7156,N_7344);
and U7511 (N_7511,N_7223,N_7490);
and U7512 (N_7512,N_7467,N_7452);
nand U7513 (N_7513,N_7377,N_7043);
nand U7514 (N_7514,N_7069,N_7141);
and U7515 (N_7515,N_7196,N_7132);
nand U7516 (N_7516,N_7127,N_7101);
nand U7517 (N_7517,N_7292,N_7100);
and U7518 (N_7518,N_7115,N_7031);
xnor U7519 (N_7519,N_7109,N_7232);
nand U7520 (N_7520,N_7039,N_7496);
and U7521 (N_7521,N_7426,N_7410);
nand U7522 (N_7522,N_7205,N_7263);
nand U7523 (N_7523,N_7018,N_7298);
or U7524 (N_7524,N_7057,N_7480);
nor U7525 (N_7525,N_7110,N_7199);
xor U7526 (N_7526,N_7225,N_7046);
nand U7527 (N_7527,N_7354,N_7423);
xnor U7528 (N_7528,N_7155,N_7059);
and U7529 (N_7529,N_7258,N_7139);
xnor U7530 (N_7530,N_7450,N_7341);
or U7531 (N_7531,N_7310,N_7076);
or U7532 (N_7532,N_7151,N_7180);
and U7533 (N_7533,N_7104,N_7021);
xor U7534 (N_7534,N_7081,N_7231);
nand U7535 (N_7535,N_7206,N_7133);
or U7536 (N_7536,N_7193,N_7413);
nand U7537 (N_7537,N_7086,N_7497);
or U7538 (N_7538,N_7473,N_7150);
nor U7539 (N_7539,N_7068,N_7058);
xor U7540 (N_7540,N_7433,N_7129);
or U7541 (N_7541,N_7342,N_7369);
or U7542 (N_7542,N_7427,N_7219);
nand U7543 (N_7543,N_7213,N_7125);
nor U7544 (N_7544,N_7164,N_7243);
nor U7545 (N_7545,N_7434,N_7272);
or U7546 (N_7546,N_7145,N_7366);
nand U7547 (N_7547,N_7078,N_7107);
xnor U7548 (N_7548,N_7353,N_7367);
nand U7549 (N_7549,N_7083,N_7430);
nor U7550 (N_7550,N_7439,N_7262);
and U7551 (N_7551,N_7061,N_7457);
xnor U7552 (N_7552,N_7192,N_7460);
nand U7553 (N_7553,N_7422,N_7052);
nor U7554 (N_7554,N_7064,N_7355);
and U7555 (N_7555,N_7040,N_7245);
or U7556 (N_7556,N_7368,N_7331);
xor U7557 (N_7557,N_7195,N_7348);
xor U7558 (N_7558,N_7340,N_7338);
nor U7559 (N_7559,N_7106,N_7337);
nand U7560 (N_7560,N_7389,N_7171);
nand U7561 (N_7561,N_7260,N_7293);
and U7562 (N_7562,N_7412,N_7112);
or U7563 (N_7563,N_7168,N_7166);
nand U7564 (N_7564,N_7070,N_7013);
nand U7565 (N_7565,N_7461,N_7240);
nand U7566 (N_7566,N_7385,N_7463);
nor U7567 (N_7567,N_7488,N_7295);
xnor U7568 (N_7568,N_7278,N_7316);
nor U7569 (N_7569,N_7188,N_7218);
and U7570 (N_7570,N_7220,N_7318);
or U7571 (N_7571,N_7097,N_7248);
and U7572 (N_7572,N_7431,N_7204);
nor U7573 (N_7573,N_7143,N_7200);
nand U7574 (N_7574,N_7015,N_7000);
and U7575 (N_7575,N_7014,N_7054);
or U7576 (N_7576,N_7401,N_7053);
nand U7577 (N_7577,N_7487,N_7235);
nand U7578 (N_7578,N_7126,N_7175);
nand U7579 (N_7579,N_7297,N_7183);
nand U7580 (N_7580,N_7075,N_7343);
nor U7581 (N_7581,N_7119,N_7425);
or U7582 (N_7582,N_7087,N_7312);
xnor U7583 (N_7583,N_7362,N_7073);
or U7584 (N_7584,N_7447,N_7379);
nor U7585 (N_7585,N_7095,N_7334);
or U7586 (N_7586,N_7409,N_7210);
and U7587 (N_7587,N_7438,N_7357);
nand U7588 (N_7588,N_7275,N_7216);
xnor U7589 (N_7589,N_7261,N_7314);
nand U7590 (N_7590,N_7130,N_7313);
and U7591 (N_7591,N_7209,N_7392);
or U7592 (N_7592,N_7019,N_7167);
xor U7593 (N_7593,N_7174,N_7026);
nor U7594 (N_7594,N_7397,N_7282);
xnor U7595 (N_7595,N_7215,N_7315);
nor U7596 (N_7596,N_7288,N_7492);
nand U7597 (N_7597,N_7178,N_7446);
and U7598 (N_7598,N_7038,N_7091);
xnor U7599 (N_7599,N_7010,N_7006);
nor U7600 (N_7600,N_7255,N_7416);
and U7601 (N_7601,N_7328,N_7254);
and U7602 (N_7602,N_7468,N_7203);
nand U7603 (N_7603,N_7402,N_7084);
or U7604 (N_7604,N_7465,N_7296);
nand U7605 (N_7605,N_7271,N_7207);
or U7606 (N_7606,N_7267,N_7499);
nor U7607 (N_7607,N_7462,N_7451);
nand U7608 (N_7608,N_7257,N_7453);
nor U7609 (N_7609,N_7339,N_7391);
xnor U7610 (N_7610,N_7214,N_7408);
nor U7611 (N_7611,N_7085,N_7077);
nor U7612 (N_7612,N_7459,N_7387);
or U7613 (N_7613,N_7056,N_7351);
nor U7614 (N_7614,N_7388,N_7202);
nand U7615 (N_7615,N_7103,N_7036);
or U7616 (N_7616,N_7148,N_7226);
nor U7617 (N_7617,N_7186,N_7009);
and U7618 (N_7618,N_7088,N_7436);
or U7619 (N_7619,N_7491,N_7432);
or U7620 (N_7620,N_7320,N_7037);
and U7621 (N_7621,N_7184,N_7324);
or U7622 (N_7622,N_7363,N_7134);
nand U7623 (N_7623,N_7269,N_7033);
nor U7624 (N_7624,N_7277,N_7050);
nand U7625 (N_7625,N_7264,N_7376);
nor U7626 (N_7626,N_7165,N_7411);
nand U7627 (N_7627,N_7445,N_7352);
xnor U7628 (N_7628,N_7071,N_7227);
or U7629 (N_7629,N_7283,N_7306);
nand U7630 (N_7630,N_7025,N_7335);
nand U7631 (N_7631,N_7259,N_7152);
and U7632 (N_7632,N_7212,N_7102);
and U7633 (N_7633,N_7382,N_7455);
xor U7634 (N_7634,N_7360,N_7198);
or U7635 (N_7635,N_7398,N_7474);
xor U7636 (N_7636,N_7381,N_7208);
nand U7637 (N_7637,N_7442,N_7279);
and U7638 (N_7638,N_7182,N_7290);
or U7639 (N_7639,N_7329,N_7370);
nand U7640 (N_7640,N_7495,N_7250);
or U7641 (N_7641,N_7333,N_7001);
xnor U7642 (N_7642,N_7177,N_7111);
and U7643 (N_7643,N_7336,N_7222);
nor U7644 (N_7644,N_7233,N_7435);
and U7645 (N_7645,N_7317,N_7270);
nand U7646 (N_7646,N_7194,N_7099);
xor U7647 (N_7647,N_7374,N_7493);
or U7648 (N_7648,N_7161,N_7027);
nor U7649 (N_7649,N_7378,N_7330);
and U7650 (N_7650,N_7236,N_7345);
or U7651 (N_7651,N_7448,N_7280);
xor U7652 (N_7652,N_7242,N_7023);
nor U7653 (N_7653,N_7063,N_7420);
nor U7654 (N_7654,N_7191,N_7386);
xnor U7655 (N_7655,N_7485,N_7291);
xor U7656 (N_7656,N_7470,N_7396);
or U7657 (N_7657,N_7454,N_7276);
xor U7658 (N_7658,N_7373,N_7029);
and U7659 (N_7659,N_7065,N_7098);
and U7660 (N_7660,N_7221,N_7414);
xnor U7661 (N_7661,N_7197,N_7147);
nand U7662 (N_7662,N_7090,N_7137);
or U7663 (N_7663,N_7266,N_7007);
nand U7664 (N_7664,N_7325,N_7241);
and U7665 (N_7665,N_7079,N_7484);
and U7666 (N_7666,N_7466,N_7486);
or U7667 (N_7667,N_7172,N_7281);
xnor U7668 (N_7668,N_7494,N_7116);
nor U7669 (N_7669,N_7289,N_7011);
nor U7670 (N_7670,N_7124,N_7356);
nor U7671 (N_7671,N_7321,N_7142);
or U7672 (N_7672,N_7286,N_7066);
and U7673 (N_7673,N_7440,N_7140);
nor U7674 (N_7674,N_7022,N_7089);
xor U7675 (N_7675,N_7238,N_7123);
and U7676 (N_7676,N_7211,N_7358);
and U7677 (N_7677,N_7136,N_7375);
nand U7678 (N_7678,N_7481,N_7449);
and U7679 (N_7679,N_7105,N_7159);
and U7680 (N_7680,N_7287,N_7224);
nor U7681 (N_7681,N_7042,N_7472);
nor U7682 (N_7682,N_7326,N_7252);
nor U7683 (N_7683,N_7476,N_7332);
nor U7684 (N_7684,N_7458,N_7265);
xnor U7685 (N_7685,N_7469,N_7304);
nand U7686 (N_7686,N_7135,N_7160);
nand U7687 (N_7687,N_7190,N_7128);
and U7688 (N_7688,N_7062,N_7201);
xor U7689 (N_7689,N_7350,N_7311);
nor U7690 (N_7690,N_7359,N_7179);
and U7691 (N_7691,N_7154,N_7234);
or U7692 (N_7692,N_7189,N_7187);
xnor U7693 (N_7693,N_7228,N_7093);
and U7694 (N_7694,N_7045,N_7285);
nor U7695 (N_7695,N_7482,N_7244);
or U7696 (N_7696,N_7307,N_7364);
and U7697 (N_7697,N_7256,N_7479);
and U7698 (N_7698,N_7096,N_7403);
xor U7699 (N_7699,N_7268,N_7173);
nor U7700 (N_7700,N_7163,N_7114);
xnor U7701 (N_7701,N_7380,N_7016);
xnor U7702 (N_7702,N_7051,N_7138);
or U7703 (N_7703,N_7158,N_7118);
or U7704 (N_7704,N_7020,N_7371);
nor U7705 (N_7705,N_7055,N_7395);
or U7706 (N_7706,N_7008,N_7404);
or U7707 (N_7707,N_7170,N_7300);
or U7708 (N_7708,N_7483,N_7464);
or U7709 (N_7709,N_7032,N_7074);
or U7710 (N_7710,N_7072,N_7004);
nor U7711 (N_7711,N_7498,N_7017);
or U7712 (N_7712,N_7478,N_7417);
xor U7713 (N_7713,N_7229,N_7305);
nor U7714 (N_7714,N_7247,N_7024);
nor U7715 (N_7715,N_7181,N_7456);
nand U7716 (N_7716,N_7030,N_7003);
nor U7717 (N_7717,N_7217,N_7060);
and U7718 (N_7718,N_7153,N_7146);
or U7719 (N_7719,N_7044,N_7308);
nor U7720 (N_7720,N_7239,N_7121);
or U7721 (N_7721,N_7176,N_7424);
nand U7722 (N_7722,N_7346,N_7349);
nor U7723 (N_7723,N_7390,N_7067);
and U7724 (N_7724,N_7302,N_7273);
and U7725 (N_7725,N_7319,N_7322);
xnor U7726 (N_7726,N_7274,N_7048);
nor U7727 (N_7727,N_7406,N_7251);
or U7728 (N_7728,N_7394,N_7012);
nor U7729 (N_7729,N_7294,N_7477);
nor U7730 (N_7730,N_7303,N_7162);
nand U7731 (N_7731,N_7082,N_7122);
and U7732 (N_7732,N_7047,N_7415);
xor U7733 (N_7733,N_7489,N_7092);
xnor U7734 (N_7734,N_7393,N_7383);
nand U7735 (N_7735,N_7117,N_7365);
nand U7736 (N_7736,N_7002,N_7113);
xor U7737 (N_7737,N_7169,N_7028);
nor U7738 (N_7738,N_7185,N_7094);
nor U7739 (N_7739,N_7253,N_7372);
nor U7740 (N_7740,N_7437,N_7399);
and U7741 (N_7741,N_7327,N_7131);
or U7742 (N_7742,N_7471,N_7429);
xnor U7743 (N_7743,N_7237,N_7443);
and U7744 (N_7744,N_7361,N_7441);
and U7745 (N_7745,N_7347,N_7323);
or U7746 (N_7746,N_7041,N_7080);
xnor U7747 (N_7747,N_7034,N_7407);
or U7748 (N_7748,N_7418,N_7005);
xor U7749 (N_7749,N_7249,N_7120);
xor U7750 (N_7750,N_7469,N_7269);
and U7751 (N_7751,N_7132,N_7479);
nor U7752 (N_7752,N_7268,N_7225);
nand U7753 (N_7753,N_7223,N_7203);
nand U7754 (N_7754,N_7287,N_7206);
or U7755 (N_7755,N_7327,N_7497);
and U7756 (N_7756,N_7139,N_7366);
nand U7757 (N_7757,N_7149,N_7002);
and U7758 (N_7758,N_7418,N_7135);
nor U7759 (N_7759,N_7318,N_7491);
xnor U7760 (N_7760,N_7272,N_7287);
nor U7761 (N_7761,N_7236,N_7334);
nor U7762 (N_7762,N_7432,N_7357);
nor U7763 (N_7763,N_7086,N_7046);
nand U7764 (N_7764,N_7319,N_7385);
or U7765 (N_7765,N_7348,N_7499);
and U7766 (N_7766,N_7080,N_7394);
nand U7767 (N_7767,N_7212,N_7261);
nor U7768 (N_7768,N_7387,N_7170);
nand U7769 (N_7769,N_7262,N_7027);
nor U7770 (N_7770,N_7383,N_7021);
or U7771 (N_7771,N_7381,N_7283);
or U7772 (N_7772,N_7211,N_7074);
or U7773 (N_7773,N_7071,N_7404);
nand U7774 (N_7774,N_7374,N_7123);
nand U7775 (N_7775,N_7473,N_7204);
xor U7776 (N_7776,N_7384,N_7261);
or U7777 (N_7777,N_7299,N_7125);
xnor U7778 (N_7778,N_7022,N_7135);
nor U7779 (N_7779,N_7294,N_7460);
nor U7780 (N_7780,N_7342,N_7214);
xnor U7781 (N_7781,N_7183,N_7365);
nor U7782 (N_7782,N_7272,N_7309);
or U7783 (N_7783,N_7027,N_7383);
nand U7784 (N_7784,N_7414,N_7481);
nor U7785 (N_7785,N_7366,N_7138);
or U7786 (N_7786,N_7182,N_7004);
and U7787 (N_7787,N_7313,N_7133);
and U7788 (N_7788,N_7267,N_7089);
and U7789 (N_7789,N_7258,N_7192);
nor U7790 (N_7790,N_7344,N_7064);
nor U7791 (N_7791,N_7022,N_7457);
and U7792 (N_7792,N_7272,N_7337);
xnor U7793 (N_7793,N_7081,N_7147);
xor U7794 (N_7794,N_7414,N_7067);
xnor U7795 (N_7795,N_7304,N_7296);
and U7796 (N_7796,N_7254,N_7435);
nand U7797 (N_7797,N_7156,N_7395);
nor U7798 (N_7798,N_7205,N_7492);
and U7799 (N_7799,N_7361,N_7202);
nor U7800 (N_7800,N_7472,N_7467);
or U7801 (N_7801,N_7114,N_7451);
or U7802 (N_7802,N_7280,N_7439);
nand U7803 (N_7803,N_7236,N_7466);
or U7804 (N_7804,N_7103,N_7238);
nor U7805 (N_7805,N_7093,N_7049);
or U7806 (N_7806,N_7379,N_7070);
or U7807 (N_7807,N_7213,N_7409);
or U7808 (N_7808,N_7268,N_7033);
nor U7809 (N_7809,N_7182,N_7256);
and U7810 (N_7810,N_7395,N_7217);
xor U7811 (N_7811,N_7205,N_7490);
nor U7812 (N_7812,N_7377,N_7052);
nor U7813 (N_7813,N_7456,N_7156);
and U7814 (N_7814,N_7275,N_7371);
or U7815 (N_7815,N_7140,N_7165);
xor U7816 (N_7816,N_7068,N_7179);
nand U7817 (N_7817,N_7118,N_7153);
nor U7818 (N_7818,N_7131,N_7389);
or U7819 (N_7819,N_7099,N_7342);
nor U7820 (N_7820,N_7397,N_7405);
and U7821 (N_7821,N_7169,N_7290);
or U7822 (N_7822,N_7101,N_7228);
or U7823 (N_7823,N_7252,N_7077);
or U7824 (N_7824,N_7150,N_7489);
or U7825 (N_7825,N_7255,N_7287);
nand U7826 (N_7826,N_7477,N_7293);
or U7827 (N_7827,N_7460,N_7496);
or U7828 (N_7828,N_7306,N_7143);
or U7829 (N_7829,N_7405,N_7334);
xor U7830 (N_7830,N_7493,N_7485);
xor U7831 (N_7831,N_7450,N_7221);
nand U7832 (N_7832,N_7267,N_7273);
nor U7833 (N_7833,N_7129,N_7080);
nor U7834 (N_7834,N_7423,N_7412);
and U7835 (N_7835,N_7061,N_7379);
and U7836 (N_7836,N_7166,N_7135);
or U7837 (N_7837,N_7066,N_7071);
nor U7838 (N_7838,N_7143,N_7420);
nor U7839 (N_7839,N_7422,N_7199);
xor U7840 (N_7840,N_7263,N_7380);
and U7841 (N_7841,N_7434,N_7487);
nor U7842 (N_7842,N_7426,N_7414);
nor U7843 (N_7843,N_7375,N_7389);
nand U7844 (N_7844,N_7045,N_7420);
or U7845 (N_7845,N_7234,N_7332);
nand U7846 (N_7846,N_7009,N_7421);
nand U7847 (N_7847,N_7358,N_7381);
and U7848 (N_7848,N_7220,N_7062);
and U7849 (N_7849,N_7433,N_7028);
and U7850 (N_7850,N_7325,N_7209);
xor U7851 (N_7851,N_7485,N_7442);
and U7852 (N_7852,N_7199,N_7177);
and U7853 (N_7853,N_7207,N_7394);
nand U7854 (N_7854,N_7333,N_7426);
nand U7855 (N_7855,N_7168,N_7253);
or U7856 (N_7856,N_7243,N_7306);
nor U7857 (N_7857,N_7320,N_7069);
nor U7858 (N_7858,N_7393,N_7451);
xor U7859 (N_7859,N_7115,N_7414);
or U7860 (N_7860,N_7364,N_7346);
or U7861 (N_7861,N_7185,N_7031);
xnor U7862 (N_7862,N_7235,N_7362);
nor U7863 (N_7863,N_7051,N_7201);
or U7864 (N_7864,N_7432,N_7445);
nor U7865 (N_7865,N_7203,N_7377);
or U7866 (N_7866,N_7421,N_7178);
or U7867 (N_7867,N_7022,N_7209);
nor U7868 (N_7868,N_7309,N_7056);
nand U7869 (N_7869,N_7055,N_7282);
and U7870 (N_7870,N_7196,N_7284);
nor U7871 (N_7871,N_7074,N_7287);
and U7872 (N_7872,N_7140,N_7414);
nor U7873 (N_7873,N_7452,N_7428);
xnor U7874 (N_7874,N_7489,N_7459);
and U7875 (N_7875,N_7257,N_7393);
or U7876 (N_7876,N_7441,N_7135);
or U7877 (N_7877,N_7209,N_7412);
or U7878 (N_7878,N_7228,N_7140);
and U7879 (N_7879,N_7295,N_7271);
nand U7880 (N_7880,N_7401,N_7499);
nand U7881 (N_7881,N_7226,N_7199);
xnor U7882 (N_7882,N_7445,N_7085);
nor U7883 (N_7883,N_7287,N_7399);
and U7884 (N_7884,N_7274,N_7405);
and U7885 (N_7885,N_7158,N_7122);
nor U7886 (N_7886,N_7488,N_7103);
xor U7887 (N_7887,N_7175,N_7213);
nand U7888 (N_7888,N_7050,N_7191);
or U7889 (N_7889,N_7470,N_7452);
nand U7890 (N_7890,N_7001,N_7228);
nand U7891 (N_7891,N_7434,N_7322);
or U7892 (N_7892,N_7256,N_7359);
nand U7893 (N_7893,N_7074,N_7343);
or U7894 (N_7894,N_7201,N_7181);
and U7895 (N_7895,N_7138,N_7242);
nand U7896 (N_7896,N_7104,N_7053);
xnor U7897 (N_7897,N_7224,N_7249);
nand U7898 (N_7898,N_7132,N_7452);
xor U7899 (N_7899,N_7071,N_7438);
and U7900 (N_7900,N_7494,N_7486);
or U7901 (N_7901,N_7124,N_7422);
or U7902 (N_7902,N_7340,N_7081);
and U7903 (N_7903,N_7312,N_7144);
nand U7904 (N_7904,N_7438,N_7241);
nand U7905 (N_7905,N_7346,N_7345);
nor U7906 (N_7906,N_7368,N_7429);
nor U7907 (N_7907,N_7228,N_7434);
nand U7908 (N_7908,N_7253,N_7292);
nor U7909 (N_7909,N_7209,N_7319);
nand U7910 (N_7910,N_7227,N_7457);
xnor U7911 (N_7911,N_7231,N_7037);
xnor U7912 (N_7912,N_7049,N_7001);
or U7913 (N_7913,N_7179,N_7045);
and U7914 (N_7914,N_7221,N_7193);
and U7915 (N_7915,N_7393,N_7317);
xnor U7916 (N_7916,N_7295,N_7454);
nand U7917 (N_7917,N_7388,N_7299);
nand U7918 (N_7918,N_7352,N_7238);
nor U7919 (N_7919,N_7347,N_7438);
nor U7920 (N_7920,N_7296,N_7232);
nor U7921 (N_7921,N_7091,N_7366);
nand U7922 (N_7922,N_7084,N_7045);
or U7923 (N_7923,N_7406,N_7465);
and U7924 (N_7924,N_7065,N_7400);
or U7925 (N_7925,N_7286,N_7012);
xor U7926 (N_7926,N_7455,N_7306);
and U7927 (N_7927,N_7015,N_7290);
xnor U7928 (N_7928,N_7145,N_7192);
xor U7929 (N_7929,N_7022,N_7447);
xnor U7930 (N_7930,N_7144,N_7350);
nand U7931 (N_7931,N_7295,N_7480);
nor U7932 (N_7932,N_7154,N_7140);
nor U7933 (N_7933,N_7440,N_7004);
xor U7934 (N_7934,N_7312,N_7106);
xnor U7935 (N_7935,N_7471,N_7089);
xnor U7936 (N_7936,N_7113,N_7412);
nor U7937 (N_7937,N_7356,N_7226);
nand U7938 (N_7938,N_7436,N_7361);
nand U7939 (N_7939,N_7204,N_7282);
or U7940 (N_7940,N_7364,N_7320);
nor U7941 (N_7941,N_7073,N_7243);
and U7942 (N_7942,N_7115,N_7374);
and U7943 (N_7943,N_7124,N_7207);
nand U7944 (N_7944,N_7204,N_7192);
nor U7945 (N_7945,N_7188,N_7172);
or U7946 (N_7946,N_7402,N_7072);
xnor U7947 (N_7947,N_7093,N_7392);
xor U7948 (N_7948,N_7452,N_7406);
nand U7949 (N_7949,N_7360,N_7060);
nand U7950 (N_7950,N_7367,N_7403);
xor U7951 (N_7951,N_7424,N_7480);
xnor U7952 (N_7952,N_7229,N_7178);
nand U7953 (N_7953,N_7070,N_7214);
xor U7954 (N_7954,N_7167,N_7040);
or U7955 (N_7955,N_7313,N_7085);
xnor U7956 (N_7956,N_7445,N_7372);
or U7957 (N_7957,N_7109,N_7406);
xnor U7958 (N_7958,N_7155,N_7397);
nor U7959 (N_7959,N_7170,N_7261);
nor U7960 (N_7960,N_7406,N_7048);
or U7961 (N_7961,N_7065,N_7419);
xnor U7962 (N_7962,N_7390,N_7007);
nor U7963 (N_7963,N_7304,N_7383);
and U7964 (N_7964,N_7395,N_7308);
xor U7965 (N_7965,N_7116,N_7394);
nand U7966 (N_7966,N_7053,N_7472);
and U7967 (N_7967,N_7031,N_7184);
nor U7968 (N_7968,N_7348,N_7283);
and U7969 (N_7969,N_7239,N_7227);
and U7970 (N_7970,N_7491,N_7151);
xor U7971 (N_7971,N_7012,N_7071);
and U7972 (N_7972,N_7412,N_7417);
xor U7973 (N_7973,N_7400,N_7394);
xor U7974 (N_7974,N_7007,N_7177);
or U7975 (N_7975,N_7394,N_7366);
nor U7976 (N_7976,N_7498,N_7440);
nand U7977 (N_7977,N_7019,N_7077);
or U7978 (N_7978,N_7484,N_7057);
xor U7979 (N_7979,N_7287,N_7453);
xnor U7980 (N_7980,N_7143,N_7128);
nor U7981 (N_7981,N_7187,N_7226);
or U7982 (N_7982,N_7292,N_7424);
xor U7983 (N_7983,N_7160,N_7418);
or U7984 (N_7984,N_7425,N_7486);
nor U7985 (N_7985,N_7448,N_7274);
and U7986 (N_7986,N_7435,N_7407);
or U7987 (N_7987,N_7369,N_7185);
or U7988 (N_7988,N_7258,N_7462);
xor U7989 (N_7989,N_7280,N_7456);
or U7990 (N_7990,N_7392,N_7083);
nor U7991 (N_7991,N_7150,N_7452);
nand U7992 (N_7992,N_7312,N_7141);
nor U7993 (N_7993,N_7326,N_7136);
or U7994 (N_7994,N_7022,N_7056);
nor U7995 (N_7995,N_7242,N_7448);
or U7996 (N_7996,N_7386,N_7480);
nor U7997 (N_7997,N_7463,N_7254);
or U7998 (N_7998,N_7235,N_7216);
nand U7999 (N_7999,N_7138,N_7354);
nand U8000 (N_8000,N_7651,N_7613);
nand U8001 (N_8001,N_7784,N_7942);
or U8002 (N_8002,N_7883,N_7557);
xnor U8003 (N_8003,N_7639,N_7568);
xnor U8004 (N_8004,N_7527,N_7904);
xor U8005 (N_8005,N_7760,N_7727);
nand U8006 (N_8006,N_7655,N_7931);
or U8007 (N_8007,N_7956,N_7567);
nor U8008 (N_8008,N_7729,N_7675);
or U8009 (N_8009,N_7552,N_7555);
and U8010 (N_8010,N_7737,N_7914);
xor U8011 (N_8011,N_7906,N_7860);
and U8012 (N_8012,N_7669,N_7505);
nor U8013 (N_8013,N_7665,N_7879);
and U8014 (N_8014,N_7550,N_7963);
or U8015 (N_8015,N_7977,N_7654);
or U8016 (N_8016,N_7582,N_7620);
or U8017 (N_8017,N_7941,N_7743);
or U8018 (N_8018,N_7578,N_7803);
and U8019 (N_8019,N_7797,N_7966);
nand U8020 (N_8020,N_7717,N_7616);
nand U8021 (N_8021,N_7626,N_7512);
xnor U8022 (N_8022,N_7907,N_7520);
nor U8023 (N_8023,N_7529,N_7916);
nand U8024 (N_8024,N_7896,N_7607);
or U8025 (N_8025,N_7998,N_7969);
xor U8026 (N_8026,N_7682,N_7551);
nor U8027 (N_8027,N_7658,N_7545);
nor U8028 (N_8028,N_7726,N_7518);
or U8029 (N_8029,N_7838,N_7762);
and U8030 (N_8030,N_7674,N_7656);
nand U8031 (N_8031,N_7662,N_7779);
or U8032 (N_8032,N_7902,N_7842);
nand U8033 (N_8033,N_7792,N_7570);
nor U8034 (N_8034,N_7770,N_7772);
xor U8035 (N_8035,N_7757,N_7575);
nor U8036 (N_8036,N_7563,N_7648);
or U8037 (N_8037,N_7560,N_7895);
nand U8038 (N_8038,N_7764,N_7927);
or U8039 (N_8039,N_7601,N_7795);
and U8040 (N_8040,N_7507,N_7704);
and U8041 (N_8041,N_7517,N_7775);
nor U8042 (N_8042,N_7844,N_7572);
and U8043 (N_8043,N_7522,N_7731);
and U8044 (N_8044,N_7548,N_7554);
and U8045 (N_8045,N_7589,N_7994);
or U8046 (N_8046,N_7872,N_7962);
xnor U8047 (N_8047,N_7787,N_7930);
nand U8048 (N_8048,N_7897,N_7983);
nor U8049 (N_8049,N_7511,N_7873);
xor U8050 (N_8050,N_7749,N_7861);
and U8051 (N_8051,N_7821,N_7853);
nand U8052 (N_8052,N_7753,N_7810);
or U8053 (N_8053,N_7680,N_7986);
and U8054 (N_8054,N_7577,N_7818);
nand U8055 (N_8055,N_7869,N_7558);
and U8056 (N_8056,N_7628,N_7791);
or U8057 (N_8057,N_7928,N_7523);
and U8058 (N_8058,N_7964,N_7666);
nand U8059 (N_8059,N_7719,N_7694);
nand U8060 (N_8060,N_7980,N_7826);
or U8061 (N_8061,N_7542,N_7696);
nor U8062 (N_8062,N_7864,N_7837);
nor U8063 (N_8063,N_7796,N_7801);
and U8064 (N_8064,N_7503,N_7936);
xnor U8065 (N_8065,N_7663,N_7659);
or U8066 (N_8066,N_7687,N_7829);
nor U8067 (N_8067,N_7874,N_7752);
nand U8068 (N_8068,N_7950,N_7627);
xnor U8069 (N_8069,N_7886,N_7723);
xor U8070 (N_8070,N_7676,N_7769);
and U8071 (N_8071,N_7871,N_7611);
nand U8072 (N_8072,N_7934,N_7865);
nor U8073 (N_8073,N_7711,N_7703);
nand U8074 (N_8074,N_7644,N_7541);
xor U8075 (N_8075,N_7825,N_7649);
xnor U8076 (N_8076,N_7882,N_7850);
nor U8077 (N_8077,N_7985,N_7773);
nor U8078 (N_8078,N_7599,N_7820);
xor U8079 (N_8079,N_7546,N_7705);
nand U8080 (N_8080,N_7580,N_7815);
and U8081 (N_8081,N_7991,N_7746);
nand U8082 (N_8082,N_7724,N_7521);
or U8083 (N_8083,N_7816,N_7640);
and U8084 (N_8084,N_7718,N_7693);
xnor U8085 (N_8085,N_7852,N_7932);
nand U8086 (N_8086,N_7984,N_7707);
and U8087 (N_8087,N_7615,N_7510);
nor U8088 (N_8088,N_7596,N_7828);
nor U8089 (N_8089,N_7780,N_7993);
or U8090 (N_8090,N_7535,N_7786);
nand U8091 (N_8091,N_7949,N_7889);
nand U8092 (N_8092,N_7681,N_7562);
nor U8093 (N_8093,N_7925,N_7894);
and U8094 (N_8094,N_7678,N_7595);
or U8095 (N_8095,N_7885,N_7530);
or U8096 (N_8096,N_7793,N_7835);
nand U8097 (N_8097,N_7622,N_7996);
xnor U8098 (N_8098,N_7621,N_7851);
and U8099 (N_8099,N_7822,N_7642);
nand U8100 (N_8100,N_7933,N_7939);
nor U8101 (N_8101,N_7641,N_7594);
nand U8102 (N_8102,N_7929,N_7576);
nor U8103 (N_8103,N_7800,N_7847);
xnor U8104 (N_8104,N_7736,N_7987);
nor U8105 (N_8105,N_7968,N_7631);
nand U8106 (N_8106,N_7892,N_7876);
xnor U8107 (N_8107,N_7982,N_7880);
and U8108 (N_8108,N_7667,N_7586);
and U8109 (N_8109,N_7893,N_7908);
nor U8110 (N_8110,N_7978,N_7782);
xor U8111 (N_8111,N_7989,N_7758);
nor U8112 (N_8112,N_7602,N_7878);
and U8113 (N_8113,N_7765,N_7961);
and U8114 (N_8114,N_7598,N_7652);
nand U8115 (N_8115,N_7597,N_7559);
nand U8116 (N_8116,N_7972,N_7856);
or U8117 (N_8117,N_7553,N_7526);
nor U8118 (N_8118,N_7730,N_7776);
and U8119 (N_8119,N_7695,N_7509);
or U8120 (N_8120,N_7664,N_7556);
xor U8121 (N_8121,N_7608,N_7735);
or U8122 (N_8122,N_7646,N_7733);
nor U8123 (N_8123,N_7960,N_7940);
xor U8124 (N_8124,N_7988,N_7643);
or U8125 (N_8125,N_7912,N_7513);
and U8126 (N_8126,N_7971,N_7630);
or U8127 (N_8127,N_7683,N_7915);
nor U8128 (N_8128,N_7836,N_7635);
or U8129 (N_8129,N_7574,N_7637);
xor U8130 (N_8130,N_7973,N_7827);
nor U8131 (N_8131,N_7650,N_7888);
nor U8132 (N_8132,N_7585,N_7617);
xnor U8133 (N_8133,N_7702,N_7911);
nand U8134 (N_8134,N_7809,N_7759);
xor U8135 (N_8135,N_7661,N_7807);
nand U8136 (N_8136,N_7877,N_7684);
or U8137 (N_8137,N_7740,N_7709);
nand U8138 (N_8138,N_7591,N_7539);
and U8139 (N_8139,N_7858,N_7806);
xor U8140 (N_8140,N_7525,N_7975);
nand U8141 (N_8141,N_7812,N_7697);
nor U8142 (N_8142,N_7913,N_7632);
xnor U8143 (N_8143,N_7751,N_7672);
or U8144 (N_8144,N_7862,N_7890);
and U8145 (N_8145,N_7745,N_7609);
and U8146 (N_8146,N_7919,N_7938);
and U8147 (N_8147,N_7706,N_7708);
xor U8148 (N_8148,N_7584,N_7742);
xnor U8149 (N_8149,N_7725,N_7824);
or U8150 (N_8150,N_7834,N_7698);
or U8151 (N_8151,N_7625,N_7804);
nor U8152 (N_8152,N_7571,N_7504);
or U8153 (N_8153,N_7830,N_7618);
nand U8154 (N_8154,N_7700,N_7965);
nand U8155 (N_8155,N_7848,N_7954);
or U8156 (N_8156,N_7688,N_7549);
or U8157 (N_8157,N_7689,N_7910);
nor U8158 (N_8158,N_7997,N_7813);
nor U8159 (N_8159,N_7900,N_7502);
nand U8160 (N_8160,N_7957,N_7612);
or U8161 (N_8161,N_7995,N_7840);
xnor U8162 (N_8162,N_7794,N_7519);
nand U8163 (N_8163,N_7788,N_7923);
nor U8164 (N_8164,N_7633,N_7747);
or U8165 (N_8165,N_7715,N_7538);
or U8166 (N_8166,N_7917,N_7720);
or U8167 (N_8167,N_7638,N_7831);
nor U8168 (N_8168,N_7778,N_7921);
nor U8169 (N_8169,N_7691,N_7817);
and U8170 (N_8170,N_7866,N_7606);
xor U8171 (N_8171,N_7660,N_7524);
or U8172 (N_8172,N_7561,N_7605);
or U8173 (N_8173,N_7564,N_7692);
xor U8174 (N_8174,N_7755,N_7543);
and U8175 (N_8175,N_7744,N_7774);
xnor U8176 (N_8176,N_7952,N_7528);
nor U8177 (N_8177,N_7540,N_7699);
and U8178 (N_8178,N_7722,N_7600);
nor U8179 (N_8179,N_7920,N_7783);
nor U8180 (N_8180,N_7768,N_7671);
and U8181 (N_8181,N_7868,N_7935);
nor U8182 (N_8182,N_7867,N_7992);
nand U8183 (N_8183,N_7855,N_7845);
xor U8184 (N_8184,N_7944,N_7958);
nand U8185 (N_8185,N_7645,N_7590);
or U8186 (N_8186,N_7839,N_7716);
nor U8187 (N_8187,N_7981,N_7514);
nor U8188 (N_8188,N_7531,N_7785);
nor U8189 (N_8189,N_7501,N_7629);
or U8190 (N_8190,N_7500,N_7647);
nand U8191 (N_8191,N_7905,N_7686);
xor U8192 (N_8192,N_7738,N_7710);
xor U8193 (N_8193,N_7634,N_7901);
nand U8194 (N_8194,N_7970,N_7581);
or U8195 (N_8195,N_7891,N_7506);
nor U8196 (N_8196,N_7841,N_7566);
nand U8197 (N_8197,N_7802,N_7734);
and U8198 (N_8198,N_7859,N_7653);
nor U8199 (N_8199,N_7604,N_7955);
xor U8200 (N_8200,N_7823,N_7573);
nand U8201 (N_8201,N_7677,N_7516);
nor U8202 (N_8202,N_7761,N_7690);
nand U8203 (N_8203,N_7610,N_7670);
and U8204 (N_8204,N_7593,N_7887);
or U8205 (N_8205,N_7943,N_7741);
xor U8206 (N_8206,N_7767,N_7739);
nor U8207 (N_8207,N_7854,N_7614);
and U8208 (N_8208,N_7771,N_7508);
and U8209 (N_8209,N_7766,N_7668);
and U8210 (N_8210,N_7849,N_7903);
nand U8211 (N_8211,N_7990,N_7870);
or U8212 (N_8212,N_7899,N_7713);
xor U8213 (N_8213,N_7979,N_7756);
or U8214 (N_8214,N_7721,N_7789);
and U8215 (N_8215,N_7732,N_7857);
and U8216 (N_8216,N_7951,N_7799);
and U8217 (N_8217,N_7763,N_7603);
or U8218 (N_8218,N_7953,N_7832);
and U8219 (N_8219,N_7843,N_7909);
or U8220 (N_8220,N_7536,N_7587);
xor U8221 (N_8221,N_7999,N_7881);
nor U8222 (N_8222,N_7636,N_7515);
xnor U8223 (N_8223,N_7565,N_7833);
xnor U8224 (N_8224,N_7846,N_7777);
xnor U8225 (N_8225,N_7926,N_7798);
or U8226 (N_8226,N_7948,N_7728);
or U8227 (N_8227,N_7808,N_7967);
or U8228 (N_8228,N_7619,N_7534);
nand U8229 (N_8229,N_7947,N_7748);
nor U8230 (N_8230,N_7583,N_7544);
xor U8231 (N_8231,N_7805,N_7946);
nand U8232 (N_8232,N_7679,N_7863);
and U8233 (N_8233,N_7673,N_7898);
nor U8234 (N_8234,N_7547,N_7814);
or U8235 (N_8235,N_7569,N_7945);
and U8236 (N_8236,N_7918,N_7701);
nand U8237 (N_8237,N_7623,N_7781);
xor U8238 (N_8238,N_7922,N_7790);
and U8239 (N_8239,N_7959,N_7924);
xor U8240 (N_8240,N_7974,N_7532);
xor U8241 (N_8241,N_7884,N_7811);
xnor U8242 (N_8242,N_7875,N_7624);
xor U8243 (N_8243,N_7588,N_7976);
or U8244 (N_8244,N_7750,N_7685);
xnor U8245 (N_8245,N_7937,N_7592);
and U8246 (N_8246,N_7657,N_7537);
xnor U8247 (N_8247,N_7754,N_7714);
and U8248 (N_8248,N_7579,N_7819);
xor U8249 (N_8249,N_7712,N_7533);
and U8250 (N_8250,N_7762,N_7706);
and U8251 (N_8251,N_7520,N_7623);
xor U8252 (N_8252,N_7608,N_7695);
nand U8253 (N_8253,N_7532,N_7589);
nand U8254 (N_8254,N_7956,N_7740);
xor U8255 (N_8255,N_7908,N_7744);
or U8256 (N_8256,N_7848,N_7653);
xor U8257 (N_8257,N_7743,N_7512);
xor U8258 (N_8258,N_7806,N_7747);
and U8259 (N_8259,N_7581,N_7952);
or U8260 (N_8260,N_7505,N_7824);
and U8261 (N_8261,N_7583,N_7841);
nand U8262 (N_8262,N_7701,N_7858);
and U8263 (N_8263,N_7907,N_7562);
nand U8264 (N_8264,N_7861,N_7626);
and U8265 (N_8265,N_7744,N_7799);
nor U8266 (N_8266,N_7528,N_7978);
xor U8267 (N_8267,N_7888,N_7736);
or U8268 (N_8268,N_7696,N_7528);
xnor U8269 (N_8269,N_7789,N_7851);
xor U8270 (N_8270,N_7515,N_7904);
and U8271 (N_8271,N_7706,N_7732);
nor U8272 (N_8272,N_7756,N_7970);
or U8273 (N_8273,N_7772,N_7671);
or U8274 (N_8274,N_7763,N_7675);
nand U8275 (N_8275,N_7878,N_7780);
nor U8276 (N_8276,N_7744,N_7755);
nand U8277 (N_8277,N_7835,N_7805);
xor U8278 (N_8278,N_7969,N_7607);
and U8279 (N_8279,N_7690,N_7684);
nor U8280 (N_8280,N_7569,N_7904);
and U8281 (N_8281,N_7601,N_7976);
and U8282 (N_8282,N_7971,N_7517);
or U8283 (N_8283,N_7796,N_7967);
and U8284 (N_8284,N_7532,N_7854);
nor U8285 (N_8285,N_7994,N_7881);
nand U8286 (N_8286,N_7693,N_7853);
or U8287 (N_8287,N_7594,N_7876);
xnor U8288 (N_8288,N_7547,N_7516);
and U8289 (N_8289,N_7882,N_7943);
nand U8290 (N_8290,N_7909,N_7642);
and U8291 (N_8291,N_7908,N_7732);
nor U8292 (N_8292,N_7806,N_7667);
nand U8293 (N_8293,N_7873,N_7621);
or U8294 (N_8294,N_7693,N_7927);
nand U8295 (N_8295,N_7945,N_7547);
or U8296 (N_8296,N_7688,N_7566);
nor U8297 (N_8297,N_7909,N_7854);
nand U8298 (N_8298,N_7701,N_7781);
and U8299 (N_8299,N_7779,N_7769);
xor U8300 (N_8300,N_7630,N_7688);
and U8301 (N_8301,N_7523,N_7767);
or U8302 (N_8302,N_7747,N_7544);
and U8303 (N_8303,N_7745,N_7614);
or U8304 (N_8304,N_7889,N_7668);
nand U8305 (N_8305,N_7782,N_7728);
nor U8306 (N_8306,N_7613,N_7758);
or U8307 (N_8307,N_7744,N_7825);
or U8308 (N_8308,N_7995,N_7521);
or U8309 (N_8309,N_7980,N_7638);
nand U8310 (N_8310,N_7792,N_7931);
and U8311 (N_8311,N_7720,N_7819);
nand U8312 (N_8312,N_7604,N_7553);
or U8313 (N_8313,N_7996,N_7709);
xor U8314 (N_8314,N_7921,N_7811);
xnor U8315 (N_8315,N_7697,N_7605);
nor U8316 (N_8316,N_7593,N_7868);
and U8317 (N_8317,N_7709,N_7932);
nand U8318 (N_8318,N_7763,N_7988);
nand U8319 (N_8319,N_7507,N_7703);
or U8320 (N_8320,N_7545,N_7982);
nand U8321 (N_8321,N_7886,N_7827);
xor U8322 (N_8322,N_7813,N_7729);
and U8323 (N_8323,N_7926,N_7660);
or U8324 (N_8324,N_7545,N_7555);
xnor U8325 (N_8325,N_7788,N_7670);
or U8326 (N_8326,N_7756,N_7644);
nand U8327 (N_8327,N_7849,N_7526);
nand U8328 (N_8328,N_7509,N_7521);
and U8329 (N_8329,N_7538,N_7754);
nand U8330 (N_8330,N_7585,N_7896);
nand U8331 (N_8331,N_7900,N_7860);
nor U8332 (N_8332,N_7554,N_7757);
nor U8333 (N_8333,N_7980,N_7881);
nand U8334 (N_8334,N_7620,N_7648);
and U8335 (N_8335,N_7896,N_7858);
nand U8336 (N_8336,N_7667,N_7711);
and U8337 (N_8337,N_7997,N_7764);
xnor U8338 (N_8338,N_7655,N_7816);
nor U8339 (N_8339,N_7711,N_7967);
xnor U8340 (N_8340,N_7750,N_7733);
nand U8341 (N_8341,N_7805,N_7583);
xnor U8342 (N_8342,N_7720,N_7727);
xor U8343 (N_8343,N_7788,N_7969);
xor U8344 (N_8344,N_7969,N_7648);
xnor U8345 (N_8345,N_7881,N_7933);
nand U8346 (N_8346,N_7722,N_7684);
and U8347 (N_8347,N_7781,N_7528);
or U8348 (N_8348,N_7761,N_7911);
nand U8349 (N_8349,N_7542,N_7954);
nand U8350 (N_8350,N_7783,N_7884);
or U8351 (N_8351,N_7800,N_7822);
nor U8352 (N_8352,N_7954,N_7839);
or U8353 (N_8353,N_7670,N_7636);
and U8354 (N_8354,N_7738,N_7833);
xnor U8355 (N_8355,N_7615,N_7974);
xor U8356 (N_8356,N_7660,N_7535);
xor U8357 (N_8357,N_7624,N_7872);
and U8358 (N_8358,N_7731,N_7758);
xnor U8359 (N_8359,N_7715,N_7840);
nand U8360 (N_8360,N_7542,N_7646);
or U8361 (N_8361,N_7906,N_7688);
or U8362 (N_8362,N_7774,N_7511);
and U8363 (N_8363,N_7681,N_7769);
nor U8364 (N_8364,N_7877,N_7537);
nand U8365 (N_8365,N_7973,N_7509);
nor U8366 (N_8366,N_7962,N_7710);
nand U8367 (N_8367,N_7516,N_7766);
nor U8368 (N_8368,N_7624,N_7850);
nand U8369 (N_8369,N_7602,N_7547);
xor U8370 (N_8370,N_7950,N_7747);
and U8371 (N_8371,N_7725,N_7894);
xnor U8372 (N_8372,N_7566,N_7514);
nor U8373 (N_8373,N_7519,N_7546);
nor U8374 (N_8374,N_7958,N_7995);
xor U8375 (N_8375,N_7991,N_7695);
and U8376 (N_8376,N_7662,N_7898);
nand U8377 (N_8377,N_7891,N_7863);
xor U8378 (N_8378,N_7710,N_7579);
and U8379 (N_8379,N_7636,N_7951);
and U8380 (N_8380,N_7657,N_7935);
nand U8381 (N_8381,N_7610,N_7770);
or U8382 (N_8382,N_7665,N_7878);
nor U8383 (N_8383,N_7747,N_7613);
and U8384 (N_8384,N_7784,N_7768);
nor U8385 (N_8385,N_7543,N_7677);
nor U8386 (N_8386,N_7884,N_7905);
nor U8387 (N_8387,N_7631,N_7578);
xnor U8388 (N_8388,N_7584,N_7831);
nand U8389 (N_8389,N_7883,N_7766);
nand U8390 (N_8390,N_7502,N_7934);
nand U8391 (N_8391,N_7663,N_7651);
nor U8392 (N_8392,N_7788,N_7762);
and U8393 (N_8393,N_7807,N_7674);
nor U8394 (N_8394,N_7869,N_7947);
nand U8395 (N_8395,N_7566,N_7952);
nor U8396 (N_8396,N_7584,N_7614);
nor U8397 (N_8397,N_7627,N_7870);
xnor U8398 (N_8398,N_7968,N_7928);
and U8399 (N_8399,N_7873,N_7941);
nand U8400 (N_8400,N_7872,N_7983);
and U8401 (N_8401,N_7778,N_7797);
nor U8402 (N_8402,N_7652,N_7922);
and U8403 (N_8403,N_7735,N_7558);
and U8404 (N_8404,N_7518,N_7606);
nor U8405 (N_8405,N_7858,N_7978);
xor U8406 (N_8406,N_7705,N_7515);
and U8407 (N_8407,N_7952,N_7665);
xnor U8408 (N_8408,N_7605,N_7644);
nand U8409 (N_8409,N_7960,N_7577);
and U8410 (N_8410,N_7677,N_7814);
or U8411 (N_8411,N_7964,N_7908);
nor U8412 (N_8412,N_7873,N_7959);
nor U8413 (N_8413,N_7866,N_7992);
or U8414 (N_8414,N_7847,N_7953);
or U8415 (N_8415,N_7833,N_7917);
and U8416 (N_8416,N_7730,N_7672);
and U8417 (N_8417,N_7839,N_7668);
and U8418 (N_8418,N_7515,N_7890);
nor U8419 (N_8419,N_7961,N_7678);
xnor U8420 (N_8420,N_7840,N_7846);
nor U8421 (N_8421,N_7743,N_7932);
nor U8422 (N_8422,N_7520,N_7541);
and U8423 (N_8423,N_7881,N_7887);
and U8424 (N_8424,N_7772,N_7859);
nand U8425 (N_8425,N_7649,N_7536);
xor U8426 (N_8426,N_7873,N_7568);
or U8427 (N_8427,N_7670,N_7828);
nor U8428 (N_8428,N_7629,N_7791);
and U8429 (N_8429,N_7553,N_7909);
and U8430 (N_8430,N_7997,N_7683);
xnor U8431 (N_8431,N_7641,N_7686);
nand U8432 (N_8432,N_7558,N_7954);
nand U8433 (N_8433,N_7736,N_7914);
and U8434 (N_8434,N_7597,N_7502);
nand U8435 (N_8435,N_7726,N_7732);
xor U8436 (N_8436,N_7502,N_7702);
xor U8437 (N_8437,N_7722,N_7608);
xor U8438 (N_8438,N_7517,N_7526);
and U8439 (N_8439,N_7963,N_7609);
nor U8440 (N_8440,N_7925,N_7623);
xor U8441 (N_8441,N_7629,N_7731);
or U8442 (N_8442,N_7755,N_7722);
xnor U8443 (N_8443,N_7708,N_7859);
nor U8444 (N_8444,N_7702,N_7635);
and U8445 (N_8445,N_7831,N_7578);
xnor U8446 (N_8446,N_7842,N_7697);
or U8447 (N_8447,N_7740,N_7565);
and U8448 (N_8448,N_7661,N_7626);
nand U8449 (N_8449,N_7710,N_7924);
nor U8450 (N_8450,N_7995,N_7868);
or U8451 (N_8451,N_7929,N_7554);
and U8452 (N_8452,N_7963,N_7886);
xnor U8453 (N_8453,N_7897,N_7560);
nand U8454 (N_8454,N_7530,N_7749);
xnor U8455 (N_8455,N_7748,N_7837);
or U8456 (N_8456,N_7777,N_7939);
nand U8457 (N_8457,N_7697,N_7633);
and U8458 (N_8458,N_7949,N_7538);
xnor U8459 (N_8459,N_7959,N_7530);
and U8460 (N_8460,N_7825,N_7765);
and U8461 (N_8461,N_7904,N_7635);
and U8462 (N_8462,N_7793,N_7763);
and U8463 (N_8463,N_7884,N_7991);
or U8464 (N_8464,N_7916,N_7805);
nor U8465 (N_8465,N_7777,N_7914);
or U8466 (N_8466,N_7845,N_7534);
and U8467 (N_8467,N_7992,N_7539);
xor U8468 (N_8468,N_7732,N_7645);
nor U8469 (N_8469,N_7807,N_7994);
nand U8470 (N_8470,N_7783,N_7643);
and U8471 (N_8471,N_7824,N_7780);
nor U8472 (N_8472,N_7929,N_7744);
xnor U8473 (N_8473,N_7867,N_7894);
nor U8474 (N_8474,N_7970,N_7818);
and U8475 (N_8475,N_7611,N_7589);
xnor U8476 (N_8476,N_7897,N_7861);
nor U8477 (N_8477,N_7557,N_7643);
and U8478 (N_8478,N_7998,N_7729);
and U8479 (N_8479,N_7685,N_7857);
or U8480 (N_8480,N_7827,N_7540);
or U8481 (N_8481,N_7585,N_7565);
xnor U8482 (N_8482,N_7794,N_7504);
or U8483 (N_8483,N_7803,N_7859);
xnor U8484 (N_8484,N_7826,N_7725);
nand U8485 (N_8485,N_7764,N_7703);
and U8486 (N_8486,N_7543,N_7549);
or U8487 (N_8487,N_7609,N_7593);
and U8488 (N_8488,N_7920,N_7816);
and U8489 (N_8489,N_7614,N_7821);
xnor U8490 (N_8490,N_7621,N_7575);
and U8491 (N_8491,N_7869,N_7962);
nor U8492 (N_8492,N_7706,N_7981);
nand U8493 (N_8493,N_7561,N_7673);
and U8494 (N_8494,N_7901,N_7531);
or U8495 (N_8495,N_7797,N_7595);
xor U8496 (N_8496,N_7825,N_7965);
nand U8497 (N_8497,N_7865,N_7811);
or U8498 (N_8498,N_7703,N_7583);
xnor U8499 (N_8499,N_7610,N_7970);
nand U8500 (N_8500,N_8091,N_8395);
xnor U8501 (N_8501,N_8238,N_8101);
and U8502 (N_8502,N_8059,N_8448);
xor U8503 (N_8503,N_8440,N_8452);
or U8504 (N_8504,N_8411,N_8247);
nor U8505 (N_8505,N_8172,N_8011);
xnor U8506 (N_8506,N_8202,N_8266);
and U8507 (N_8507,N_8294,N_8430);
nor U8508 (N_8508,N_8005,N_8392);
nand U8509 (N_8509,N_8475,N_8278);
nand U8510 (N_8510,N_8189,N_8180);
and U8511 (N_8511,N_8296,N_8456);
or U8512 (N_8512,N_8056,N_8303);
nand U8513 (N_8513,N_8227,N_8451);
or U8514 (N_8514,N_8040,N_8201);
nor U8515 (N_8515,N_8494,N_8467);
or U8516 (N_8516,N_8268,N_8207);
nor U8517 (N_8517,N_8106,N_8142);
and U8518 (N_8518,N_8433,N_8048);
and U8519 (N_8519,N_8254,N_8442);
and U8520 (N_8520,N_8031,N_8118);
and U8521 (N_8521,N_8480,N_8140);
nor U8522 (N_8522,N_8054,N_8316);
xor U8523 (N_8523,N_8282,N_8065);
nor U8524 (N_8524,N_8079,N_8021);
nor U8525 (N_8525,N_8166,N_8214);
nand U8526 (N_8526,N_8099,N_8152);
or U8527 (N_8527,N_8043,N_8212);
and U8528 (N_8528,N_8388,N_8309);
and U8529 (N_8529,N_8276,N_8478);
nor U8530 (N_8530,N_8449,N_8137);
and U8531 (N_8531,N_8485,N_8330);
and U8532 (N_8532,N_8499,N_8439);
nor U8533 (N_8533,N_8029,N_8389);
or U8534 (N_8534,N_8125,N_8258);
xnor U8535 (N_8535,N_8299,N_8413);
and U8536 (N_8536,N_8138,N_8374);
or U8537 (N_8537,N_8130,N_8195);
xnor U8538 (N_8538,N_8127,N_8100);
nor U8539 (N_8539,N_8486,N_8492);
and U8540 (N_8540,N_8487,N_8306);
xor U8541 (N_8541,N_8033,N_8012);
or U8542 (N_8542,N_8421,N_8200);
nor U8543 (N_8543,N_8081,N_8329);
nor U8544 (N_8544,N_8162,N_8479);
nand U8545 (N_8545,N_8169,N_8277);
xnor U8546 (N_8546,N_8148,N_8382);
and U8547 (N_8547,N_8213,N_8211);
xnor U8548 (N_8548,N_8004,N_8481);
nand U8549 (N_8549,N_8006,N_8473);
or U8550 (N_8550,N_8197,N_8075);
or U8551 (N_8551,N_8024,N_8412);
or U8552 (N_8552,N_8185,N_8359);
and U8553 (N_8553,N_8019,N_8154);
nor U8554 (N_8554,N_8049,N_8241);
nand U8555 (N_8555,N_8318,N_8377);
nor U8556 (N_8556,N_8465,N_8369);
nand U8557 (N_8557,N_8074,N_8469);
nand U8558 (N_8558,N_8186,N_8236);
nand U8559 (N_8559,N_8003,N_8471);
and U8560 (N_8560,N_8490,N_8151);
or U8561 (N_8561,N_8260,N_8067);
nor U8562 (N_8562,N_8443,N_8016);
xor U8563 (N_8563,N_8115,N_8007);
nor U8564 (N_8564,N_8176,N_8349);
xor U8565 (N_8565,N_8183,N_8437);
xnor U8566 (N_8566,N_8105,N_8089);
xnor U8567 (N_8567,N_8410,N_8322);
xor U8568 (N_8568,N_8163,N_8310);
xnor U8569 (N_8569,N_8270,N_8466);
nor U8570 (N_8570,N_8356,N_8333);
nor U8571 (N_8571,N_8293,N_8221);
and U8572 (N_8572,N_8290,N_8464);
and U8573 (N_8573,N_8351,N_8233);
xor U8574 (N_8574,N_8405,N_8242);
and U8575 (N_8575,N_8263,N_8335);
nor U8576 (N_8576,N_8041,N_8387);
nor U8577 (N_8577,N_8325,N_8145);
nand U8578 (N_8578,N_8379,N_8331);
xor U8579 (N_8579,N_8368,N_8171);
or U8580 (N_8580,N_8143,N_8231);
nand U8581 (N_8581,N_8086,N_8435);
nor U8582 (N_8582,N_8354,N_8234);
nor U8583 (N_8583,N_8337,N_8248);
nand U8584 (N_8584,N_8170,N_8450);
nand U8585 (N_8585,N_8446,N_8253);
and U8586 (N_8586,N_8257,N_8239);
nand U8587 (N_8587,N_8396,N_8085);
and U8588 (N_8588,N_8216,N_8114);
and U8589 (N_8589,N_8121,N_8493);
nand U8590 (N_8590,N_8256,N_8157);
or U8591 (N_8591,N_8230,N_8414);
nor U8592 (N_8592,N_8308,N_8052);
nand U8593 (N_8593,N_8066,N_8340);
xnor U8594 (N_8594,N_8071,N_8319);
xor U8595 (N_8595,N_8491,N_8057);
nor U8596 (N_8596,N_8397,N_8039);
or U8597 (N_8597,N_8399,N_8243);
xor U8598 (N_8598,N_8376,N_8002);
nand U8599 (N_8599,N_8470,N_8431);
nor U8600 (N_8600,N_8317,N_8275);
and U8601 (N_8601,N_8196,N_8014);
or U8602 (N_8602,N_8198,N_8417);
nand U8603 (N_8603,N_8080,N_8217);
xnor U8604 (N_8604,N_8098,N_8459);
xor U8605 (N_8605,N_8441,N_8182);
xnor U8606 (N_8606,N_8334,N_8199);
or U8607 (N_8607,N_8476,N_8267);
nor U8608 (N_8608,N_8280,N_8461);
or U8609 (N_8609,N_8482,N_8312);
and U8610 (N_8610,N_8281,N_8174);
nor U8611 (N_8611,N_8009,N_8111);
nand U8612 (N_8612,N_8249,N_8053);
and U8613 (N_8613,N_8336,N_8190);
nor U8614 (N_8614,N_8415,N_8062);
and U8615 (N_8615,N_8072,N_8133);
or U8616 (N_8616,N_8323,N_8032);
or U8617 (N_8617,N_8285,N_8068);
nand U8618 (N_8618,N_8432,N_8372);
xor U8619 (N_8619,N_8426,N_8167);
xor U8620 (N_8620,N_8168,N_8010);
nand U8621 (N_8621,N_8416,N_8371);
xor U8622 (N_8622,N_8300,N_8025);
nor U8623 (N_8623,N_8283,N_8135);
and U8624 (N_8624,N_8398,N_8287);
nand U8625 (N_8625,N_8188,N_8423);
nand U8626 (N_8626,N_8246,N_8204);
or U8627 (N_8627,N_8366,N_8077);
and U8628 (N_8628,N_8453,N_8206);
xnor U8629 (N_8629,N_8209,N_8373);
and U8630 (N_8630,N_8307,N_8360);
nor U8631 (N_8631,N_8403,N_8288);
xnor U8632 (N_8632,N_8215,N_8332);
xor U8633 (N_8633,N_8208,N_8424);
xor U8634 (N_8634,N_8223,N_8327);
nand U8635 (N_8635,N_8386,N_8017);
xnor U8636 (N_8636,N_8347,N_8191);
xnor U8637 (N_8637,N_8484,N_8164);
or U8638 (N_8638,N_8401,N_8272);
nand U8639 (N_8639,N_8244,N_8344);
nand U8640 (N_8640,N_8455,N_8020);
nor U8641 (N_8641,N_8084,N_8314);
or U8642 (N_8642,N_8255,N_8123);
or U8643 (N_8643,N_8144,N_8358);
or U8644 (N_8644,N_8124,N_8245);
xnor U8645 (N_8645,N_8063,N_8434);
nor U8646 (N_8646,N_8346,N_8261);
or U8647 (N_8647,N_8076,N_8109);
nor U8648 (N_8648,N_8390,N_8116);
xor U8649 (N_8649,N_8418,N_8292);
and U8650 (N_8650,N_8165,N_8311);
nand U8651 (N_8651,N_8146,N_8113);
and U8652 (N_8652,N_8226,N_8220);
nor U8653 (N_8653,N_8402,N_8419);
or U8654 (N_8654,N_8134,N_8218);
or U8655 (N_8655,N_8122,N_8385);
xor U8656 (N_8656,N_8219,N_8128);
or U8657 (N_8657,N_8436,N_8400);
xnor U8658 (N_8658,N_8097,N_8210);
nor U8659 (N_8659,N_8407,N_8046);
xor U8660 (N_8660,N_8147,N_8082);
or U8661 (N_8661,N_8297,N_8015);
and U8662 (N_8662,N_8050,N_8051);
xor U8663 (N_8663,N_8107,N_8184);
xnor U8664 (N_8664,N_8380,N_8315);
nand U8665 (N_8665,N_8187,N_8000);
nand U8666 (N_8666,N_8240,N_8295);
nor U8667 (N_8667,N_8409,N_8090);
or U8668 (N_8668,N_8286,N_8394);
nor U8669 (N_8669,N_8047,N_8279);
and U8670 (N_8670,N_8444,N_8458);
or U8671 (N_8671,N_8013,N_8108);
nor U8672 (N_8672,N_8381,N_8445);
xor U8673 (N_8673,N_8222,N_8305);
and U8674 (N_8674,N_8044,N_8361);
xnor U8675 (N_8675,N_8362,N_8205);
and U8676 (N_8676,N_8406,N_8422);
nor U8677 (N_8677,N_8357,N_8259);
nand U8678 (N_8678,N_8438,N_8364);
xor U8679 (N_8679,N_8110,N_8095);
and U8680 (N_8680,N_8161,N_8028);
nand U8681 (N_8681,N_8173,N_8141);
or U8682 (N_8682,N_8060,N_8262);
xor U8683 (N_8683,N_8037,N_8391);
nand U8684 (N_8684,N_8393,N_8289);
and U8685 (N_8685,N_8178,N_8120);
or U8686 (N_8686,N_8030,N_8045);
or U8687 (N_8687,N_8181,N_8155);
or U8688 (N_8688,N_8192,N_8355);
xnor U8689 (N_8689,N_8078,N_8136);
or U8690 (N_8690,N_8427,N_8265);
xnor U8691 (N_8691,N_8193,N_8363);
xnor U8692 (N_8692,N_8179,N_8027);
or U8693 (N_8693,N_8008,N_8149);
nand U8694 (N_8694,N_8343,N_8061);
nor U8695 (N_8695,N_8001,N_8150);
or U8696 (N_8696,N_8301,N_8158);
and U8697 (N_8697,N_8269,N_8420);
or U8698 (N_8698,N_8474,N_8273);
nor U8699 (N_8699,N_8497,N_8404);
nand U8700 (N_8700,N_8264,N_8104);
nor U8701 (N_8701,N_8058,N_8064);
nand U8702 (N_8702,N_8468,N_8018);
or U8703 (N_8703,N_8225,N_8083);
or U8704 (N_8704,N_8129,N_8119);
or U8705 (N_8705,N_8271,N_8425);
xor U8706 (N_8706,N_8320,N_8378);
nor U8707 (N_8707,N_8353,N_8087);
and U8708 (N_8708,N_8177,N_8291);
nand U8709 (N_8709,N_8088,N_8023);
xnor U8710 (N_8710,N_8462,N_8022);
nand U8711 (N_8711,N_8313,N_8338);
xor U8712 (N_8712,N_8350,N_8384);
nand U8713 (N_8713,N_8203,N_8348);
or U8714 (N_8714,N_8339,N_8408);
xnor U8715 (N_8715,N_8228,N_8472);
nand U8716 (N_8716,N_8498,N_8495);
nor U8717 (N_8717,N_8457,N_8092);
or U8718 (N_8718,N_8232,N_8042);
or U8719 (N_8719,N_8463,N_8126);
nand U8720 (N_8720,N_8038,N_8447);
nand U8721 (N_8721,N_8345,N_8159);
nor U8722 (N_8722,N_8194,N_8073);
nor U8723 (N_8723,N_8321,N_8304);
xor U8724 (N_8724,N_8352,N_8160);
or U8725 (N_8725,N_8117,N_8365);
or U8726 (N_8726,N_8034,N_8454);
nor U8727 (N_8727,N_8036,N_8460);
nor U8728 (N_8728,N_8055,N_8341);
nor U8729 (N_8729,N_8175,N_8139);
and U8730 (N_8730,N_8274,N_8237);
xor U8731 (N_8731,N_8250,N_8035);
nor U8732 (N_8732,N_8112,N_8094);
or U8733 (N_8733,N_8131,N_8069);
nor U8734 (N_8734,N_8252,N_8375);
and U8735 (N_8735,N_8235,N_8153);
or U8736 (N_8736,N_8428,N_8483);
or U8737 (N_8737,N_8102,N_8383);
xnor U8738 (N_8738,N_8298,N_8489);
xnor U8739 (N_8739,N_8477,N_8488);
nor U8740 (N_8740,N_8132,N_8429);
or U8741 (N_8741,N_8224,N_8367);
xnor U8742 (N_8742,N_8370,N_8342);
or U8743 (N_8743,N_8324,N_8093);
xnor U8744 (N_8744,N_8302,N_8026);
and U8745 (N_8745,N_8496,N_8328);
xnor U8746 (N_8746,N_8284,N_8103);
and U8747 (N_8747,N_8251,N_8156);
nand U8748 (N_8748,N_8229,N_8096);
nor U8749 (N_8749,N_8326,N_8070);
or U8750 (N_8750,N_8124,N_8440);
and U8751 (N_8751,N_8489,N_8038);
or U8752 (N_8752,N_8006,N_8432);
nand U8753 (N_8753,N_8324,N_8401);
nand U8754 (N_8754,N_8184,N_8261);
nand U8755 (N_8755,N_8101,N_8379);
xor U8756 (N_8756,N_8182,N_8281);
nor U8757 (N_8757,N_8353,N_8039);
nand U8758 (N_8758,N_8388,N_8116);
xor U8759 (N_8759,N_8031,N_8412);
nor U8760 (N_8760,N_8431,N_8201);
or U8761 (N_8761,N_8402,N_8092);
nor U8762 (N_8762,N_8241,N_8376);
and U8763 (N_8763,N_8148,N_8025);
xor U8764 (N_8764,N_8120,N_8457);
nand U8765 (N_8765,N_8061,N_8328);
and U8766 (N_8766,N_8177,N_8145);
nand U8767 (N_8767,N_8108,N_8360);
nand U8768 (N_8768,N_8347,N_8438);
nor U8769 (N_8769,N_8398,N_8083);
xor U8770 (N_8770,N_8283,N_8318);
nand U8771 (N_8771,N_8061,N_8337);
nor U8772 (N_8772,N_8482,N_8212);
or U8773 (N_8773,N_8092,N_8148);
and U8774 (N_8774,N_8401,N_8276);
nor U8775 (N_8775,N_8194,N_8334);
nor U8776 (N_8776,N_8241,N_8047);
nand U8777 (N_8777,N_8493,N_8216);
or U8778 (N_8778,N_8093,N_8051);
nor U8779 (N_8779,N_8307,N_8309);
nand U8780 (N_8780,N_8039,N_8071);
or U8781 (N_8781,N_8102,N_8054);
nor U8782 (N_8782,N_8100,N_8309);
and U8783 (N_8783,N_8345,N_8237);
and U8784 (N_8784,N_8200,N_8328);
or U8785 (N_8785,N_8480,N_8337);
nor U8786 (N_8786,N_8298,N_8103);
xnor U8787 (N_8787,N_8487,N_8377);
and U8788 (N_8788,N_8315,N_8204);
nand U8789 (N_8789,N_8285,N_8168);
and U8790 (N_8790,N_8355,N_8118);
nand U8791 (N_8791,N_8191,N_8092);
and U8792 (N_8792,N_8220,N_8102);
and U8793 (N_8793,N_8326,N_8448);
nor U8794 (N_8794,N_8372,N_8309);
nand U8795 (N_8795,N_8403,N_8338);
and U8796 (N_8796,N_8387,N_8252);
nand U8797 (N_8797,N_8053,N_8449);
nor U8798 (N_8798,N_8178,N_8492);
nor U8799 (N_8799,N_8051,N_8129);
nand U8800 (N_8800,N_8409,N_8184);
or U8801 (N_8801,N_8248,N_8153);
or U8802 (N_8802,N_8028,N_8353);
nand U8803 (N_8803,N_8154,N_8010);
nor U8804 (N_8804,N_8182,N_8015);
xnor U8805 (N_8805,N_8270,N_8062);
nand U8806 (N_8806,N_8271,N_8236);
xnor U8807 (N_8807,N_8139,N_8153);
or U8808 (N_8808,N_8225,N_8331);
xnor U8809 (N_8809,N_8242,N_8155);
or U8810 (N_8810,N_8189,N_8213);
or U8811 (N_8811,N_8472,N_8443);
nor U8812 (N_8812,N_8013,N_8309);
xor U8813 (N_8813,N_8341,N_8219);
nand U8814 (N_8814,N_8415,N_8370);
and U8815 (N_8815,N_8123,N_8222);
nor U8816 (N_8816,N_8157,N_8424);
or U8817 (N_8817,N_8475,N_8194);
nand U8818 (N_8818,N_8035,N_8106);
or U8819 (N_8819,N_8373,N_8052);
xor U8820 (N_8820,N_8260,N_8232);
xor U8821 (N_8821,N_8412,N_8035);
or U8822 (N_8822,N_8480,N_8235);
xnor U8823 (N_8823,N_8401,N_8381);
and U8824 (N_8824,N_8177,N_8125);
xnor U8825 (N_8825,N_8006,N_8068);
and U8826 (N_8826,N_8082,N_8329);
or U8827 (N_8827,N_8219,N_8070);
and U8828 (N_8828,N_8317,N_8319);
or U8829 (N_8829,N_8020,N_8066);
nand U8830 (N_8830,N_8451,N_8357);
nand U8831 (N_8831,N_8212,N_8381);
xor U8832 (N_8832,N_8423,N_8399);
nand U8833 (N_8833,N_8062,N_8042);
nand U8834 (N_8834,N_8277,N_8241);
nor U8835 (N_8835,N_8321,N_8153);
nand U8836 (N_8836,N_8465,N_8275);
and U8837 (N_8837,N_8216,N_8116);
xor U8838 (N_8838,N_8342,N_8059);
nor U8839 (N_8839,N_8333,N_8472);
xnor U8840 (N_8840,N_8148,N_8464);
and U8841 (N_8841,N_8239,N_8358);
xnor U8842 (N_8842,N_8085,N_8260);
nand U8843 (N_8843,N_8461,N_8324);
nor U8844 (N_8844,N_8281,N_8175);
nor U8845 (N_8845,N_8187,N_8313);
or U8846 (N_8846,N_8152,N_8106);
or U8847 (N_8847,N_8156,N_8013);
xnor U8848 (N_8848,N_8168,N_8264);
nand U8849 (N_8849,N_8040,N_8433);
xnor U8850 (N_8850,N_8147,N_8300);
nand U8851 (N_8851,N_8321,N_8446);
xnor U8852 (N_8852,N_8301,N_8219);
and U8853 (N_8853,N_8200,N_8196);
nand U8854 (N_8854,N_8213,N_8114);
nor U8855 (N_8855,N_8289,N_8411);
nor U8856 (N_8856,N_8232,N_8098);
and U8857 (N_8857,N_8011,N_8370);
nand U8858 (N_8858,N_8258,N_8015);
and U8859 (N_8859,N_8488,N_8460);
nor U8860 (N_8860,N_8217,N_8390);
and U8861 (N_8861,N_8487,N_8027);
nand U8862 (N_8862,N_8462,N_8148);
or U8863 (N_8863,N_8223,N_8393);
and U8864 (N_8864,N_8052,N_8471);
nor U8865 (N_8865,N_8066,N_8279);
or U8866 (N_8866,N_8364,N_8304);
nand U8867 (N_8867,N_8373,N_8151);
or U8868 (N_8868,N_8357,N_8225);
or U8869 (N_8869,N_8382,N_8259);
or U8870 (N_8870,N_8481,N_8064);
nor U8871 (N_8871,N_8057,N_8243);
and U8872 (N_8872,N_8286,N_8413);
and U8873 (N_8873,N_8009,N_8211);
nand U8874 (N_8874,N_8078,N_8345);
xnor U8875 (N_8875,N_8431,N_8303);
and U8876 (N_8876,N_8319,N_8253);
or U8877 (N_8877,N_8270,N_8471);
nor U8878 (N_8878,N_8313,N_8148);
and U8879 (N_8879,N_8038,N_8388);
nand U8880 (N_8880,N_8352,N_8440);
nor U8881 (N_8881,N_8483,N_8081);
xnor U8882 (N_8882,N_8087,N_8130);
nor U8883 (N_8883,N_8054,N_8268);
nand U8884 (N_8884,N_8000,N_8401);
xnor U8885 (N_8885,N_8278,N_8125);
xor U8886 (N_8886,N_8476,N_8132);
and U8887 (N_8887,N_8448,N_8106);
and U8888 (N_8888,N_8310,N_8471);
xor U8889 (N_8889,N_8100,N_8171);
nand U8890 (N_8890,N_8013,N_8385);
or U8891 (N_8891,N_8150,N_8238);
nand U8892 (N_8892,N_8357,N_8342);
nor U8893 (N_8893,N_8097,N_8390);
nor U8894 (N_8894,N_8089,N_8409);
xor U8895 (N_8895,N_8258,N_8470);
and U8896 (N_8896,N_8252,N_8411);
nor U8897 (N_8897,N_8330,N_8082);
nand U8898 (N_8898,N_8089,N_8318);
xor U8899 (N_8899,N_8151,N_8116);
xnor U8900 (N_8900,N_8363,N_8284);
xor U8901 (N_8901,N_8102,N_8461);
and U8902 (N_8902,N_8204,N_8285);
nand U8903 (N_8903,N_8409,N_8358);
nand U8904 (N_8904,N_8463,N_8484);
nor U8905 (N_8905,N_8246,N_8082);
nand U8906 (N_8906,N_8136,N_8469);
xor U8907 (N_8907,N_8258,N_8262);
nor U8908 (N_8908,N_8031,N_8320);
nand U8909 (N_8909,N_8229,N_8458);
and U8910 (N_8910,N_8331,N_8238);
xnor U8911 (N_8911,N_8308,N_8109);
nand U8912 (N_8912,N_8245,N_8280);
xnor U8913 (N_8913,N_8424,N_8204);
xnor U8914 (N_8914,N_8145,N_8078);
or U8915 (N_8915,N_8357,N_8263);
nor U8916 (N_8916,N_8058,N_8209);
nand U8917 (N_8917,N_8445,N_8069);
nand U8918 (N_8918,N_8026,N_8241);
nor U8919 (N_8919,N_8333,N_8427);
xor U8920 (N_8920,N_8197,N_8278);
nor U8921 (N_8921,N_8020,N_8169);
or U8922 (N_8922,N_8427,N_8306);
or U8923 (N_8923,N_8048,N_8316);
and U8924 (N_8924,N_8109,N_8050);
nand U8925 (N_8925,N_8454,N_8100);
nand U8926 (N_8926,N_8241,N_8083);
xnor U8927 (N_8927,N_8084,N_8309);
nor U8928 (N_8928,N_8171,N_8446);
nor U8929 (N_8929,N_8089,N_8305);
or U8930 (N_8930,N_8023,N_8438);
and U8931 (N_8931,N_8456,N_8250);
and U8932 (N_8932,N_8346,N_8160);
nand U8933 (N_8933,N_8060,N_8197);
and U8934 (N_8934,N_8469,N_8356);
xnor U8935 (N_8935,N_8127,N_8012);
nor U8936 (N_8936,N_8172,N_8447);
or U8937 (N_8937,N_8407,N_8356);
and U8938 (N_8938,N_8297,N_8277);
nor U8939 (N_8939,N_8068,N_8219);
or U8940 (N_8940,N_8401,N_8169);
xnor U8941 (N_8941,N_8020,N_8466);
and U8942 (N_8942,N_8146,N_8310);
nand U8943 (N_8943,N_8320,N_8005);
nand U8944 (N_8944,N_8013,N_8426);
nor U8945 (N_8945,N_8158,N_8087);
or U8946 (N_8946,N_8177,N_8294);
nand U8947 (N_8947,N_8093,N_8400);
xor U8948 (N_8948,N_8484,N_8340);
nand U8949 (N_8949,N_8002,N_8172);
xnor U8950 (N_8950,N_8433,N_8423);
xnor U8951 (N_8951,N_8374,N_8484);
or U8952 (N_8952,N_8309,N_8178);
xor U8953 (N_8953,N_8181,N_8206);
or U8954 (N_8954,N_8453,N_8153);
or U8955 (N_8955,N_8448,N_8081);
or U8956 (N_8956,N_8412,N_8279);
nor U8957 (N_8957,N_8468,N_8174);
xnor U8958 (N_8958,N_8181,N_8320);
xnor U8959 (N_8959,N_8188,N_8080);
or U8960 (N_8960,N_8353,N_8095);
nor U8961 (N_8961,N_8331,N_8307);
nand U8962 (N_8962,N_8230,N_8115);
nor U8963 (N_8963,N_8429,N_8311);
or U8964 (N_8964,N_8195,N_8477);
nor U8965 (N_8965,N_8086,N_8174);
nor U8966 (N_8966,N_8076,N_8258);
or U8967 (N_8967,N_8311,N_8152);
nand U8968 (N_8968,N_8280,N_8035);
and U8969 (N_8969,N_8270,N_8459);
and U8970 (N_8970,N_8150,N_8023);
or U8971 (N_8971,N_8060,N_8164);
nand U8972 (N_8972,N_8328,N_8347);
or U8973 (N_8973,N_8473,N_8392);
xor U8974 (N_8974,N_8108,N_8405);
or U8975 (N_8975,N_8034,N_8328);
xor U8976 (N_8976,N_8359,N_8191);
xor U8977 (N_8977,N_8161,N_8266);
xnor U8978 (N_8978,N_8193,N_8124);
nand U8979 (N_8979,N_8400,N_8402);
and U8980 (N_8980,N_8370,N_8129);
and U8981 (N_8981,N_8401,N_8418);
or U8982 (N_8982,N_8143,N_8473);
or U8983 (N_8983,N_8127,N_8270);
xor U8984 (N_8984,N_8089,N_8493);
and U8985 (N_8985,N_8221,N_8149);
xnor U8986 (N_8986,N_8105,N_8111);
and U8987 (N_8987,N_8127,N_8219);
nand U8988 (N_8988,N_8410,N_8150);
xnor U8989 (N_8989,N_8457,N_8130);
or U8990 (N_8990,N_8193,N_8369);
nor U8991 (N_8991,N_8050,N_8118);
xor U8992 (N_8992,N_8461,N_8203);
xor U8993 (N_8993,N_8317,N_8230);
xnor U8994 (N_8994,N_8324,N_8231);
nor U8995 (N_8995,N_8365,N_8051);
and U8996 (N_8996,N_8010,N_8279);
nor U8997 (N_8997,N_8390,N_8459);
or U8998 (N_8998,N_8309,N_8072);
nor U8999 (N_8999,N_8177,N_8355);
nor U9000 (N_9000,N_8898,N_8659);
or U9001 (N_9001,N_8909,N_8977);
nand U9002 (N_9002,N_8609,N_8925);
xor U9003 (N_9003,N_8825,N_8502);
and U9004 (N_9004,N_8641,N_8830);
or U9005 (N_9005,N_8796,N_8892);
and U9006 (N_9006,N_8788,N_8700);
or U9007 (N_9007,N_8776,N_8970);
nand U9008 (N_9008,N_8561,N_8553);
or U9009 (N_9009,N_8602,N_8521);
or U9010 (N_9010,N_8777,N_8538);
and U9011 (N_9011,N_8670,N_8893);
nor U9012 (N_9012,N_8965,N_8587);
or U9013 (N_9013,N_8944,N_8960);
nand U9014 (N_9014,N_8604,N_8613);
and U9015 (N_9015,N_8639,N_8720);
and U9016 (N_9016,N_8527,N_8867);
xor U9017 (N_9017,N_8590,N_8769);
or U9018 (N_9018,N_8738,N_8576);
or U9019 (N_9019,N_8837,N_8882);
nand U9020 (N_9020,N_8993,N_8775);
xor U9021 (N_9021,N_8808,N_8983);
or U9022 (N_9022,N_8801,N_8517);
and U9023 (N_9023,N_8969,N_8821);
nor U9024 (N_9024,N_8530,N_8608);
or U9025 (N_9025,N_8935,N_8795);
nor U9026 (N_9026,N_8577,N_8570);
xnor U9027 (N_9027,N_8809,N_8884);
nand U9028 (N_9028,N_8961,N_8774);
nand U9029 (N_9029,N_8971,N_8828);
or U9030 (N_9030,N_8900,N_8792);
and U9031 (N_9031,N_8584,N_8683);
xor U9032 (N_9032,N_8981,N_8621);
nor U9033 (N_9033,N_8747,N_8630);
xnor U9034 (N_9034,N_8885,N_8948);
nor U9035 (N_9035,N_8928,N_8655);
and U9036 (N_9036,N_8735,N_8695);
nor U9037 (N_9037,N_8758,N_8542);
nor U9038 (N_9038,N_8878,N_8618);
nand U9039 (N_9039,N_8813,N_8514);
xor U9040 (N_9040,N_8790,N_8725);
nor U9041 (N_9041,N_8930,N_8671);
nor U9042 (N_9042,N_8847,N_8840);
and U9043 (N_9043,N_8525,N_8889);
nor U9044 (N_9044,N_8508,N_8660);
xnor U9045 (N_9045,N_8708,N_8888);
nor U9046 (N_9046,N_8994,N_8690);
xnor U9047 (N_9047,N_8642,N_8619);
and U9048 (N_9048,N_8819,N_8558);
nor U9049 (N_9049,N_8824,N_8681);
nand U9050 (N_9050,N_8543,N_8927);
or U9051 (N_9051,N_8728,N_8833);
xnor U9052 (N_9052,N_8737,N_8754);
nor U9053 (N_9053,N_8890,N_8665);
xnor U9054 (N_9054,N_8835,N_8805);
xnor U9055 (N_9055,N_8924,N_8583);
nor U9056 (N_9056,N_8581,N_8586);
or U9057 (N_9057,N_8854,N_8875);
or U9058 (N_9058,N_8629,N_8532);
or U9059 (N_9059,N_8549,N_8512);
nand U9060 (N_9060,N_8863,N_8667);
and U9061 (N_9061,N_8915,N_8964);
and U9062 (N_9062,N_8816,N_8533);
and U9063 (N_9063,N_8919,N_8832);
nor U9064 (N_9064,N_8741,N_8922);
nor U9065 (N_9065,N_8931,N_8736);
nand U9066 (N_9066,N_8614,N_8666);
or U9067 (N_9067,N_8858,N_8963);
or U9068 (N_9068,N_8731,N_8519);
nor U9069 (N_9069,N_8691,N_8680);
and U9070 (N_9070,N_8992,N_8950);
and U9071 (N_9071,N_8559,N_8810);
nand U9072 (N_9072,N_8723,N_8877);
and U9073 (N_9073,N_8803,N_8669);
xor U9074 (N_9074,N_8946,N_8988);
or U9075 (N_9075,N_8941,N_8640);
xnor U9076 (N_9076,N_8607,N_8886);
nor U9077 (N_9077,N_8540,N_8504);
nand U9078 (N_9078,N_8507,N_8582);
and U9079 (N_9079,N_8516,N_8763);
and U9080 (N_9080,N_8696,N_8566);
nand U9081 (N_9081,N_8851,N_8568);
nand U9082 (N_9082,N_8596,N_8715);
or U9083 (N_9083,N_8580,N_8780);
xnor U9084 (N_9084,N_8980,N_8622);
xnor U9085 (N_9085,N_8697,N_8673);
nor U9086 (N_9086,N_8500,N_8779);
xor U9087 (N_9087,N_8879,N_8637);
or U9088 (N_9088,N_8743,N_8501);
xor U9089 (N_9089,N_8784,N_8675);
or U9090 (N_9090,N_8766,N_8672);
and U9091 (N_9091,N_8520,N_8511);
or U9092 (N_9092,N_8987,N_8555);
or U9093 (N_9093,N_8979,N_8638);
xnor U9094 (N_9094,N_8649,N_8903);
and U9095 (N_9095,N_8518,N_8906);
and U9096 (N_9096,N_8554,N_8986);
nand U9097 (N_9097,N_8579,N_8949);
and U9098 (N_9098,N_8818,N_8881);
and U9099 (N_9099,N_8959,N_8611);
or U9100 (N_9100,N_8645,N_8615);
nor U9101 (N_9101,N_8545,N_8872);
or U9102 (N_9102,N_8745,N_8907);
nand U9103 (N_9103,N_8902,N_8564);
nor U9104 (N_9104,N_8871,N_8546);
xor U9105 (N_9105,N_8727,N_8541);
nor U9106 (N_9106,N_8764,N_8967);
or U9107 (N_9107,N_8975,N_8913);
or U9108 (N_9108,N_8524,N_8855);
or U9109 (N_9109,N_8591,N_8605);
and U9110 (N_9110,N_8709,N_8815);
nor U9111 (N_9111,N_8874,N_8701);
nor U9112 (N_9112,N_8678,N_8684);
nor U9113 (N_9113,N_8523,N_8560);
nand U9114 (N_9114,N_8556,N_8938);
nand U9115 (N_9115,N_8998,N_8823);
nand U9116 (N_9116,N_8714,N_8995);
or U9117 (N_9117,N_8749,N_8997);
nor U9118 (N_9118,N_8510,N_8911);
and U9119 (N_9119,N_8850,N_8651);
nor U9120 (N_9120,N_8838,N_8771);
and U9121 (N_9121,N_8572,N_8712);
nor U9122 (N_9122,N_8534,N_8646);
nor U9123 (N_9123,N_8624,N_8866);
and U9124 (N_9124,N_8748,N_8899);
nor U9125 (N_9125,N_8952,N_8929);
xnor U9126 (N_9126,N_8940,N_8968);
nand U9127 (N_9127,N_8706,N_8954);
nor U9128 (N_9128,N_8601,N_8772);
nand U9129 (N_9129,N_8908,N_8565);
nor U9130 (N_9130,N_8513,N_8578);
xor U9131 (N_9131,N_8632,N_8793);
or U9132 (N_9132,N_8933,N_8845);
or U9133 (N_9133,N_8785,N_8797);
xor U9134 (N_9134,N_8734,N_8921);
or U9135 (N_9135,N_8569,N_8563);
xor U9136 (N_9136,N_8873,N_8635);
xor U9137 (N_9137,N_8936,N_8852);
nand U9138 (N_9138,N_8916,N_8778);
nand U9139 (N_9139,N_8689,N_8699);
nor U9140 (N_9140,N_8599,N_8860);
nor U9141 (N_9141,N_8751,N_8827);
nor U9142 (N_9142,N_8917,N_8759);
nand U9143 (N_9143,N_8550,N_8990);
nand U9144 (N_9144,N_8687,N_8647);
nor U9145 (N_9145,N_8802,N_8552);
and U9146 (N_9146,N_8923,N_8868);
or U9147 (N_9147,N_8829,N_8600);
or U9148 (N_9148,N_8826,N_8726);
nand U9149 (N_9149,N_8679,N_8702);
and U9150 (N_9150,N_8627,N_8870);
nor U9151 (N_9151,N_8656,N_8861);
nand U9152 (N_9152,N_8710,N_8806);
xor U9153 (N_9153,N_8891,N_8713);
xor U9154 (N_9154,N_8616,N_8551);
xor U9155 (N_9155,N_8887,N_8703);
or U9156 (N_9156,N_8798,N_8592);
or U9157 (N_9157,N_8762,N_8973);
or U9158 (N_9158,N_8999,N_8634);
xor U9159 (N_9159,N_8989,N_8739);
nand U9160 (N_9160,N_8844,N_8658);
nor U9161 (N_9161,N_8531,N_8991);
nor U9162 (N_9162,N_8529,N_8515);
or U9163 (N_9163,N_8814,N_8953);
xor U9164 (N_9164,N_8588,N_8742);
nor U9165 (N_9165,N_8732,N_8905);
nand U9166 (N_9166,N_8982,N_8768);
xor U9167 (N_9167,N_8528,N_8765);
or U9168 (N_9168,N_8603,N_8760);
nor U9169 (N_9169,N_8733,N_8939);
and U9170 (N_9170,N_8914,N_8834);
nor U9171 (N_9171,N_8722,N_8926);
or U9172 (N_9172,N_8910,N_8620);
xor U9173 (N_9173,N_8562,N_8755);
and U9174 (N_9174,N_8985,N_8897);
nand U9175 (N_9175,N_8643,N_8962);
nor U9176 (N_9176,N_8957,N_8794);
nand U9177 (N_9177,N_8682,N_8846);
nor U9178 (N_9178,N_8756,N_8869);
or U9179 (N_9179,N_8817,N_8623);
and U9180 (N_9180,N_8839,N_8894);
nor U9181 (N_9181,N_8978,N_8781);
and U9182 (N_9182,N_8544,N_8506);
nand U9183 (N_9183,N_8711,N_8676);
and U9184 (N_9184,N_8585,N_8597);
and U9185 (N_9185,N_8606,N_8744);
xnor U9186 (N_9186,N_8761,N_8920);
nand U9187 (N_9187,N_8698,N_8862);
nand U9188 (N_9188,N_8942,N_8804);
and U9189 (N_9189,N_8901,N_8589);
xnor U9190 (N_9190,N_8557,N_8896);
nor U9191 (N_9191,N_8654,N_8664);
or U9192 (N_9192,N_8571,N_8753);
nand U9193 (N_9193,N_8791,N_8996);
xor U9194 (N_9194,N_8943,N_8612);
or U9195 (N_9195,N_8865,N_8856);
and U9196 (N_9196,N_8843,N_8598);
nor U9197 (N_9197,N_8574,N_8807);
nand U9198 (N_9198,N_8536,N_8841);
nand U9199 (N_9199,N_8800,N_8822);
or U9200 (N_9200,N_8767,N_8853);
xnor U9201 (N_9201,N_8773,N_8648);
or U9202 (N_9202,N_8705,N_8718);
or U9203 (N_9203,N_8610,N_8918);
nor U9204 (N_9204,N_8674,N_8663);
nor U9205 (N_9205,N_8704,N_8811);
nor U9206 (N_9206,N_8812,N_8535);
xnor U9207 (N_9207,N_8787,N_8857);
nor U9208 (N_9208,N_8864,N_8668);
nor U9209 (N_9209,N_8876,N_8686);
nor U9210 (N_9210,N_8974,N_8724);
and U9211 (N_9211,N_8836,N_8522);
nand U9212 (N_9212,N_8677,N_8692);
or U9213 (N_9213,N_8625,N_8904);
xor U9214 (N_9214,N_8955,N_8958);
nand U9215 (N_9215,N_8650,N_8782);
or U9216 (N_9216,N_8859,N_8548);
nor U9217 (N_9217,N_8783,N_8626);
nor U9218 (N_9218,N_8831,N_8757);
nor U9219 (N_9219,N_8595,N_8842);
nor U9220 (N_9220,N_8746,N_8883);
nor U9221 (N_9221,N_8657,N_8567);
or U9222 (N_9222,N_8770,N_8593);
nor U9223 (N_9223,N_8934,N_8912);
or U9224 (N_9224,N_8721,N_8537);
nand U9225 (N_9225,N_8547,N_8661);
or U9226 (N_9226,N_8932,N_8505);
xnor U9227 (N_9227,N_8895,N_8789);
nand U9228 (N_9228,N_8631,N_8509);
or U9229 (N_9229,N_8539,N_8628);
or U9230 (N_9230,N_8972,N_8820);
nand U9231 (N_9231,N_8740,N_8693);
nor U9232 (N_9232,N_8503,N_8937);
nor U9233 (N_9233,N_8594,N_8880);
or U9234 (N_9234,N_8685,N_8752);
or U9235 (N_9235,N_8786,N_8717);
nand U9236 (N_9236,N_8662,N_8750);
nand U9237 (N_9237,N_8688,N_8644);
nand U9238 (N_9238,N_8947,N_8799);
or U9239 (N_9239,N_8633,N_8653);
nand U9240 (N_9240,N_8984,N_8945);
and U9241 (N_9241,N_8849,N_8652);
and U9242 (N_9242,N_8617,N_8976);
nor U9243 (N_9243,N_8719,N_8729);
nand U9244 (N_9244,N_8526,N_8707);
nand U9245 (N_9245,N_8956,N_8730);
nor U9246 (N_9246,N_8848,N_8716);
nor U9247 (N_9247,N_8636,N_8694);
nand U9248 (N_9248,N_8573,N_8966);
and U9249 (N_9249,N_8575,N_8951);
and U9250 (N_9250,N_8999,N_8522);
nand U9251 (N_9251,N_8812,N_8932);
nor U9252 (N_9252,N_8689,N_8971);
nor U9253 (N_9253,N_8838,N_8787);
and U9254 (N_9254,N_8829,N_8670);
and U9255 (N_9255,N_8669,N_8696);
nand U9256 (N_9256,N_8766,N_8683);
and U9257 (N_9257,N_8945,N_8664);
nand U9258 (N_9258,N_8534,N_8934);
or U9259 (N_9259,N_8763,N_8569);
nand U9260 (N_9260,N_8654,N_8513);
and U9261 (N_9261,N_8682,N_8917);
or U9262 (N_9262,N_8853,N_8932);
or U9263 (N_9263,N_8891,N_8941);
nor U9264 (N_9264,N_8738,N_8997);
nor U9265 (N_9265,N_8598,N_8681);
nand U9266 (N_9266,N_8539,N_8588);
or U9267 (N_9267,N_8622,N_8803);
xnor U9268 (N_9268,N_8807,N_8776);
nand U9269 (N_9269,N_8600,N_8779);
nand U9270 (N_9270,N_8940,N_8695);
or U9271 (N_9271,N_8522,N_8650);
or U9272 (N_9272,N_8784,N_8917);
nor U9273 (N_9273,N_8977,N_8817);
or U9274 (N_9274,N_8693,N_8746);
nand U9275 (N_9275,N_8838,N_8918);
and U9276 (N_9276,N_8662,N_8600);
and U9277 (N_9277,N_8733,N_8823);
xnor U9278 (N_9278,N_8533,N_8970);
or U9279 (N_9279,N_8856,N_8807);
xnor U9280 (N_9280,N_8746,N_8729);
nand U9281 (N_9281,N_8881,N_8778);
nor U9282 (N_9282,N_8575,N_8690);
or U9283 (N_9283,N_8910,N_8827);
nor U9284 (N_9284,N_8915,N_8901);
or U9285 (N_9285,N_8954,N_8999);
or U9286 (N_9286,N_8603,N_8655);
xor U9287 (N_9287,N_8599,N_8805);
and U9288 (N_9288,N_8826,N_8905);
and U9289 (N_9289,N_8875,N_8869);
xor U9290 (N_9290,N_8733,N_8554);
xor U9291 (N_9291,N_8594,N_8569);
or U9292 (N_9292,N_8582,N_8664);
and U9293 (N_9293,N_8886,N_8532);
nor U9294 (N_9294,N_8519,N_8997);
xnor U9295 (N_9295,N_8629,N_8513);
and U9296 (N_9296,N_8560,N_8984);
nor U9297 (N_9297,N_8605,N_8559);
nor U9298 (N_9298,N_8869,N_8710);
nand U9299 (N_9299,N_8910,N_8817);
nor U9300 (N_9300,N_8790,N_8987);
xnor U9301 (N_9301,N_8796,N_8529);
or U9302 (N_9302,N_8508,N_8690);
xor U9303 (N_9303,N_8866,N_8916);
xor U9304 (N_9304,N_8716,N_8986);
or U9305 (N_9305,N_8984,N_8806);
and U9306 (N_9306,N_8853,N_8575);
xnor U9307 (N_9307,N_8659,N_8917);
nand U9308 (N_9308,N_8888,N_8979);
or U9309 (N_9309,N_8642,N_8862);
and U9310 (N_9310,N_8806,N_8574);
and U9311 (N_9311,N_8688,N_8918);
and U9312 (N_9312,N_8538,N_8817);
nand U9313 (N_9313,N_8985,N_8689);
or U9314 (N_9314,N_8620,N_8929);
nand U9315 (N_9315,N_8831,N_8776);
nor U9316 (N_9316,N_8879,N_8869);
xnor U9317 (N_9317,N_8998,N_8500);
nand U9318 (N_9318,N_8927,N_8721);
and U9319 (N_9319,N_8616,N_8595);
or U9320 (N_9320,N_8992,N_8769);
nand U9321 (N_9321,N_8727,N_8835);
xor U9322 (N_9322,N_8580,N_8862);
and U9323 (N_9323,N_8902,N_8535);
nor U9324 (N_9324,N_8973,N_8621);
or U9325 (N_9325,N_8642,N_8595);
nand U9326 (N_9326,N_8901,N_8900);
or U9327 (N_9327,N_8719,N_8899);
or U9328 (N_9328,N_8627,N_8594);
and U9329 (N_9329,N_8985,N_8800);
or U9330 (N_9330,N_8642,N_8881);
xnor U9331 (N_9331,N_8913,N_8878);
or U9332 (N_9332,N_8826,N_8722);
nor U9333 (N_9333,N_8590,N_8991);
nor U9334 (N_9334,N_8632,N_8664);
or U9335 (N_9335,N_8857,N_8681);
or U9336 (N_9336,N_8690,N_8788);
or U9337 (N_9337,N_8828,N_8741);
xor U9338 (N_9338,N_8520,N_8999);
or U9339 (N_9339,N_8534,N_8617);
xnor U9340 (N_9340,N_8793,N_8781);
and U9341 (N_9341,N_8953,N_8715);
or U9342 (N_9342,N_8885,N_8891);
nor U9343 (N_9343,N_8762,N_8525);
and U9344 (N_9344,N_8716,N_8971);
nor U9345 (N_9345,N_8914,N_8502);
and U9346 (N_9346,N_8776,N_8600);
nand U9347 (N_9347,N_8559,N_8729);
nand U9348 (N_9348,N_8942,N_8941);
nand U9349 (N_9349,N_8935,N_8759);
and U9350 (N_9350,N_8818,N_8590);
xnor U9351 (N_9351,N_8973,N_8880);
nor U9352 (N_9352,N_8630,N_8790);
nand U9353 (N_9353,N_8604,N_8699);
nand U9354 (N_9354,N_8854,N_8930);
and U9355 (N_9355,N_8757,N_8563);
and U9356 (N_9356,N_8807,N_8603);
nand U9357 (N_9357,N_8692,N_8552);
or U9358 (N_9358,N_8601,N_8734);
xnor U9359 (N_9359,N_8844,N_8582);
or U9360 (N_9360,N_8841,N_8916);
and U9361 (N_9361,N_8877,N_8569);
and U9362 (N_9362,N_8591,N_8576);
nor U9363 (N_9363,N_8921,N_8571);
xnor U9364 (N_9364,N_8920,N_8977);
nor U9365 (N_9365,N_8977,N_8635);
or U9366 (N_9366,N_8878,N_8539);
nand U9367 (N_9367,N_8683,N_8908);
or U9368 (N_9368,N_8630,N_8516);
nor U9369 (N_9369,N_8806,N_8543);
nand U9370 (N_9370,N_8582,N_8637);
and U9371 (N_9371,N_8871,N_8592);
nand U9372 (N_9372,N_8554,N_8843);
nand U9373 (N_9373,N_8880,N_8834);
or U9374 (N_9374,N_8582,N_8860);
xor U9375 (N_9375,N_8718,N_8678);
nand U9376 (N_9376,N_8608,N_8534);
nor U9377 (N_9377,N_8730,N_8650);
or U9378 (N_9378,N_8530,N_8955);
nand U9379 (N_9379,N_8828,N_8670);
nor U9380 (N_9380,N_8567,N_8845);
nand U9381 (N_9381,N_8747,N_8514);
nor U9382 (N_9382,N_8773,N_8926);
xnor U9383 (N_9383,N_8950,N_8655);
nand U9384 (N_9384,N_8641,N_8918);
or U9385 (N_9385,N_8520,N_8525);
nand U9386 (N_9386,N_8941,N_8766);
and U9387 (N_9387,N_8662,N_8983);
nor U9388 (N_9388,N_8852,N_8543);
nand U9389 (N_9389,N_8761,N_8811);
and U9390 (N_9390,N_8650,N_8871);
xor U9391 (N_9391,N_8757,N_8662);
or U9392 (N_9392,N_8899,N_8990);
xnor U9393 (N_9393,N_8754,N_8794);
or U9394 (N_9394,N_8812,N_8938);
and U9395 (N_9395,N_8537,N_8588);
nand U9396 (N_9396,N_8884,N_8502);
nor U9397 (N_9397,N_8907,N_8636);
and U9398 (N_9398,N_8699,N_8668);
nor U9399 (N_9399,N_8755,N_8549);
xnor U9400 (N_9400,N_8607,N_8817);
xnor U9401 (N_9401,N_8860,N_8688);
or U9402 (N_9402,N_8594,N_8866);
nor U9403 (N_9403,N_8599,N_8882);
xnor U9404 (N_9404,N_8558,N_8549);
xnor U9405 (N_9405,N_8871,N_8945);
xnor U9406 (N_9406,N_8873,N_8523);
nor U9407 (N_9407,N_8827,N_8573);
nand U9408 (N_9408,N_8866,N_8595);
nor U9409 (N_9409,N_8875,N_8526);
or U9410 (N_9410,N_8728,N_8718);
nand U9411 (N_9411,N_8587,N_8981);
or U9412 (N_9412,N_8712,N_8996);
and U9413 (N_9413,N_8712,N_8500);
nor U9414 (N_9414,N_8592,N_8975);
and U9415 (N_9415,N_8805,N_8593);
xor U9416 (N_9416,N_8688,N_8818);
and U9417 (N_9417,N_8991,N_8779);
nand U9418 (N_9418,N_8651,N_8670);
nand U9419 (N_9419,N_8835,N_8713);
or U9420 (N_9420,N_8821,N_8828);
nand U9421 (N_9421,N_8839,N_8564);
xor U9422 (N_9422,N_8909,N_8781);
nand U9423 (N_9423,N_8812,N_8750);
or U9424 (N_9424,N_8680,N_8641);
xnor U9425 (N_9425,N_8548,N_8944);
xor U9426 (N_9426,N_8967,N_8611);
xnor U9427 (N_9427,N_8761,N_8712);
nor U9428 (N_9428,N_8590,N_8754);
nand U9429 (N_9429,N_8758,N_8614);
and U9430 (N_9430,N_8978,N_8533);
or U9431 (N_9431,N_8712,N_8558);
nor U9432 (N_9432,N_8672,N_8514);
and U9433 (N_9433,N_8780,N_8617);
nand U9434 (N_9434,N_8512,N_8973);
and U9435 (N_9435,N_8613,N_8881);
xor U9436 (N_9436,N_8848,N_8895);
nor U9437 (N_9437,N_8588,N_8862);
or U9438 (N_9438,N_8876,N_8920);
nand U9439 (N_9439,N_8792,N_8977);
nand U9440 (N_9440,N_8878,N_8923);
nand U9441 (N_9441,N_8905,N_8892);
and U9442 (N_9442,N_8919,N_8859);
xnor U9443 (N_9443,N_8772,N_8940);
nand U9444 (N_9444,N_8622,N_8935);
and U9445 (N_9445,N_8972,N_8973);
and U9446 (N_9446,N_8973,N_8746);
nor U9447 (N_9447,N_8923,N_8873);
xor U9448 (N_9448,N_8999,N_8738);
or U9449 (N_9449,N_8568,N_8750);
xnor U9450 (N_9450,N_8741,N_8914);
nand U9451 (N_9451,N_8563,N_8647);
and U9452 (N_9452,N_8538,N_8910);
and U9453 (N_9453,N_8511,N_8692);
or U9454 (N_9454,N_8951,N_8628);
nand U9455 (N_9455,N_8516,N_8654);
nand U9456 (N_9456,N_8870,N_8699);
xor U9457 (N_9457,N_8572,N_8587);
nor U9458 (N_9458,N_8573,N_8854);
and U9459 (N_9459,N_8517,N_8799);
nor U9460 (N_9460,N_8977,N_8713);
nor U9461 (N_9461,N_8577,N_8582);
nor U9462 (N_9462,N_8500,N_8705);
and U9463 (N_9463,N_8903,N_8644);
xnor U9464 (N_9464,N_8593,N_8707);
or U9465 (N_9465,N_8586,N_8510);
nand U9466 (N_9466,N_8880,N_8615);
xor U9467 (N_9467,N_8884,N_8603);
nor U9468 (N_9468,N_8740,N_8899);
or U9469 (N_9469,N_8984,N_8627);
or U9470 (N_9470,N_8678,N_8942);
nand U9471 (N_9471,N_8707,N_8636);
and U9472 (N_9472,N_8716,N_8981);
nor U9473 (N_9473,N_8597,N_8844);
xnor U9474 (N_9474,N_8660,N_8565);
nor U9475 (N_9475,N_8965,N_8980);
xnor U9476 (N_9476,N_8748,N_8882);
xor U9477 (N_9477,N_8515,N_8983);
and U9478 (N_9478,N_8858,N_8691);
and U9479 (N_9479,N_8624,N_8794);
or U9480 (N_9480,N_8570,N_8546);
or U9481 (N_9481,N_8609,N_8802);
or U9482 (N_9482,N_8689,N_8706);
or U9483 (N_9483,N_8937,N_8596);
or U9484 (N_9484,N_8803,N_8734);
or U9485 (N_9485,N_8881,N_8666);
nor U9486 (N_9486,N_8541,N_8536);
nor U9487 (N_9487,N_8913,N_8600);
xor U9488 (N_9488,N_8882,N_8937);
xor U9489 (N_9489,N_8707,N_8559);
and U9490 (N_9490,N_8853,N_8630);
xnor U9491 (N_9491,N_8849,N_8643);
and U9492 (N_9492,N_8705,N_8999);
nor U9493 (N_9493,N_8811,N_8599);
and U9494 (N_9494,N_8775,N_8545);
or U9495 (N_9495,N_8938,N_8834);
nand U9496 (N_9496,N_8512,N_8960);
nor U9497 (N_9497,N_8665,N_8724);
and U9498 (N_9498,N_8874,N_8781);
nand U9499 (N_9499,N_8667,N_8507);
xor U9500 (N_9500,N_9477,N_9388);
xnor U9501 (N_9501,N_9338,N_9305);
or U9502 (N_9502,N_9250,N_9099);
or U9503 (N_9503,N_9365,N_9128);
and U9504 (N_9504,N_9419,N_9283);
nand U9505 (N_9505,N_9176,N_9225);
nand U9506 (N_9506,N_9348,N_9003);
nor U9507 (N_9507,N_9385,N_9401);
or U9508 (N_9508,N_9321,N_9229);
or U9509 (N_9509,N_9200,N_9312);
nor U9510 (N_9510,N_9123,N_9342);
nand U9511 (N_9511,N_9032,N_9344);
nor U9512 (N_9512,N_9166,N_9150);
nand U9513 (N_9513,N_9400,N_9202);
xor U9514 (N_9514,N_9011,N_9278);
nor U9515 (N_9515,N_9377,N_9062);
nand U9516 (N_9516,N_9289,N_9423);
nor U9517 (N_9517,N_9366,N_9258);
xor U9518 (N_9518,N_9059,N_9075);
nor U9519 (N_9519,N_9384,N_9493);
nand U9520 (N_9520,N_9345,N_9104);
nor U9521 (N_9521,N_9374,N_9389);
or U9522 (N_9522,N_9380,N_9251);
and U9523 (N_9523,N_9252,N_9387);
nand U9524 (N_9524,N_9192,N_9030);
xnor U9525 (N_9525,N_9358,N_9432);
or U9526 (N_9526,N_9240,N_9210);
or U9527 (N_9527,N_9051,N_9332);
nand U9528 (N_9528,N_9163,N_9143);
nor U9529 (N_9529,N_9067,N_9077);
xnor U9530 (N_9530,N_9456,N_9110);
and U9531 (N_9531,N_9390,N_9415);
or U9532 (N_9532,N_9406,N_9352);
or U9533 (N_9533,N_9125,N_9159);
nor U9534 (N_9534,N_9084,N_9096);
xnor U9535 (N_9535,N_9023,N_9160);
xnor U9536 (N_9536,N_9187,N_9324);
nand U9537 (N_9537,N_9444,N_9040);
or U9538 (N_9538,N_9437,N_9412);
nand U9539 (N_9539,N_9363,N_9318);
and U9540 (N_9540,N_9362,N_9281);
xnor U9541 (N_9541,N_9114,N_9413);
or U9542 (N_9542,N_9111,N_9264);
and U9543 (N_9543,N_9426,N_9103);
and U9544 (N_9544,N_9214,N_9292);
xor U9545 (N_9545,N_9145,N_9325);
or U9546 (N_9546,N_9147,N_9036);
or U9547 (N_9547,N_9495,N_9431);
or U9548 (N_9548,N_9138,N_9155);
nand U9549 (N_9549,N_9314,N_9022);
nand U9550 (N_9550,N_9248,N_9140);
and U9551 (N_9551,N_9317,N_9007);
and U9552 (N_9552,N_9304,N_9121);
xor U9553 (N_9553,N_9204,N_9439);
and U9554 (N_9554,N_9127,N_9405);
and U9555 (N_9555,N_9162,N_9326);
xor U9556 (N_9556,N_9486,N_9279);
or U9557 (N_9557,N_9336,N_9260);
nand U9558 (N_9558,N_9115,N_9467);
xor U9559 (N_9559,N_9201,N_9037);
or U9560 (N_9560,N_9015,N_9347);
and U9561 (N_9561,N_9466,N_9130);
nor U9562 (N_9562,N_9141,N_9284);
or U9563 (N_9563,N_9424,N_9392);
xor U9564 (N_9564,N_9106,N_9095);
nand U9565 (N_9565,N_9409,N_9257);
nand U9566 (N_9566,N_9013,N_9208);
or U9567 (N_9567,N_9183,N_9033);
and U9568 (N_9568,N_9158,N_9256);
nand U9569 (N_9569,N_9116,N_9083);
nand U9570 (N_9570,N_9132,N_9061);
xnor U9571 (N_9571,N_9349,N_9451);
nand U9572 (N_9572,N_9148,N_9499);
nand U9573 (N_9573,N_9286,N_9319);
or U9574 (N_9574,N_9496,N_9422);
and U9575 (N_9575,N_9274,N_9381);
or U9576 (N_9576,N_9494,N_9194);
nand U9577 (N_9577,N_9177,N_9359);
and U9578 (N_9578,N_9025,N_9246);
and U9579 (N_9579,N_9006,N_9203);
nor U9580 (N_9580,N_9307,N_9418);
or U9581 (N_9581,N_9399,N_9055);
xor U9582 (N_9582,N_9393,N_9049);
xnor U9583 (N_9583,N_9243,N_9330);
xor U9584 (N_9584,N_9222,N_9092);
nand U9585 (N_9585,N_9100,N_9382);
nor U9586 (N_9586,N_9164,N_9275);
nor U9587 (N_9587,N_9199,N_9396);
xor U9588 (N_9588,N_9124,N_9320);
nand U9589 (N_9589,N_9196,N_9403);
xnor U9590 (N_9590,N_9476,N_9178);
or U9591 (N_9591,N_9433,N_9218);
and U9592 (N_9592,N_9453,N_9249);
nor U9593 (N_9593,N_9310,N_9149);
nor U9594 (N_9594,N_9153,N_9017);
nand U9595 (N_9595,N_9063,N_9410);
nor U9596 (N_9596,N_9407,N_9489);
xnor U9597 (N_9597,N_9072,N_9161);
nor U9598 (N_9598,N_9438,N_9480);
and U9599 (N_9599,N_9420,N_9473);
nand U9600 (N_9600,N_9404,N_9282);
or U9601 (N_9601,N_9000,N_9491);
or U9602 (N_9602,N_9171,N_9212);
nor U9603 (N_9603,N_9378,N_9078);
and U9604 (N_9604,N_9105,N_9157);
or U9605 (N_9605,N_9335,N_9024);
xnor U9606 (N_9606,N_9101,N_9117);
or U9607 (N_9607,N_9300,N_9154);
xor U9608 (N_9608,N_9226,N_9206);
or U9609 (N_9609,N_9056,N_9402);
nand U9610 (N_9610,N_9221,N_9189);
xor U9611 (N_9611,N_9004,N_9265);
xnor U9612 (N_9612,N_9268,N_9361);
and U9613 (N_9613,N_9175,N_9233);
xnor U9614 (N_9614,N_9207,N_9168);
or U9615 (N_9615,N_9058,N_9440);
nand U9616 (N_9616,N_9383,N_9186);
and U9617 (N_9617,N_9459,N_9443);
xnor U9618 (N_9618,N_9395,N_9098);
xnor U9619 (N_9619,N_9454,N_9146);
nor U9620 (N_9620,N_9241,N_9446);
nand U9621 (N_9621,N_9089,N_9370);
xor U9622 (N_9622,N_9090,N_9118);
nor U9623 (N_9623,N_9375,N_9427);
xor U9624 (N_9624,N_9185,N_9215);
nand U9625 (N_9625,N_9244,N_9340);
xor U9626 (N_9626,N_9434,N_9134);
nor U9627 (N_9627,N_9193,N_9041);
nor U9628 (N_9628,N_9452,N_9216);
nand U9629 (N_9629,N_9197,N_9137);
nand U9630 (N_9630,N_9180,N_9122);
xor U9631 (N_9631,N_9231,N_9093);
xnor U9632 (N_9632,N_9356,N_9429);
xnor U9633 (N_9633,N_9047,N_9136);
or U9634 (N_9634,N_9054,N_9277);
and U9635 (N_9635,N_9042,N_9205);
or U9636 (N_9636,N_9060,N_9211);
nor U9637 (N_9637,N_9082,N_9035);
nor U9638 (N_9638,N_9045,N_9167);
nor U9639 (N_9639,N_9485,N_9328);
xor U9640 (N_9640,N_9273,N_9014);
and U9641 (N_9641,N_9367,N_9027);
xor U9642 (N_9642,N_9043,N_9308);
xor U9643 (N_9643,N_9253,N_9369);
or U9644 (N_9644,N_9497,N_9169);
nand U9645 (N_9645,N_9484,N_9165);
xor U9646 (N_9646,N_9131,N_9009);
or U9647 (N_9647,N_9492,N_9181);
and U9648 (N_9648,N_9087,N_9213);
or U9649 (N_9649,N_9425,N_9010);
and U9650 (N_9650,N_9309,N_9120);
xnor U9651 (N_9651,N_9228,N_9088);
or U9652 (N_9652,N_9302,N_9259);
nor U9653 (N_9653,N_9331,N_9235);
nor U9654 (N_9654,N_9044,N_9152);
nor U9655 (N_9655,N_9303,N_9108);
nand U9656 (N_9656,N_9269,N_9109);
xor U9657 (N_9657,N_9239,N_9364);
xnor U9658 (N_9658,N_9018,N_9301);
xnor U9659 (N_9659,N_9139,N_9291);
and U9660 (N_9660,N_9488,N_9074);
or U9661 (N_9661,N_9133,N_9463);
or U9662 (N_9662,N_9091,N_9073);
nand U9663 (N_9663,N_9034,N_9411);
nor U9664 (N_9664,N_9234,N_9262);
nand U9665 (N_9665,N_9053,N_9195);
nor U9666 (N_9666,N_9315,N_9064);
xnor U9667 (N_9667,N_9080,N_9442);
nor U9668 (N_9668,N_9144,N_9297);
nor U9669 (N_9669,N_9271,N_9019);
or U9670 (N_9670,N_9479,N_9126);
nand U9671 (N_9671,N_9232,N_9005);
xnor U9672 (N_9672,N_9272,N_9142);
or U9673 (N_9673,N_9245,N_9094);
and U9674 (N_9674,N_9065,N_9428);
or U9675 (N_9675,N_9327,N_9290);
nand U9676 (N_9676,N_9316,N_9386);
nand U9677 (N_9677,N_9227,N_9468);
and U9678 (N_9678,N_9028,N_9371);
nand U9679 (N_9679,N_9230,N_9474);
nor U9680 (N_9680,N_9191,N_9172);
or U9681 (N_9681,N_9391,N_9002);
nand U9682 (N_9682,N_9285,N_9470);
and U9683 (N_9683,N_9322,N_9217);
nor U9684 (N_9684,N_9416,N_9112);
or U9685 (N_9685,N_9306,N_9334);
nor U9686 (N_9686,N_9038,N_9031);
xnor U9687 (N_9687,N_9295,N_9066);
nand U9688 (N_9688,N_9490,N_9135);
and U9689 (N_9689,N_9398,N_9255);
nor U9690 (N_9690,N_9076,N_9263);
or U9691 (N_9691,N_9293,N_9313);
or U9692 (N_9692,N_9483,N_9458);
nand U9693 (N_9693,N_9498,N_9224);
xor U9694 (N_9694,N_9280,N_9461);
nand U9695 (N_9695,N_9057,N_9294);
nand U9696 (N_9696,N_9357,N_9350);
or U9697 (N_9697,N_9001,N_9299);
nand U9698 (N_9698,N_9460,N_9276);
and U9699 (N_9699,N_9351,N_9156);
and U9700 (N_9700,N_9346,N_9012);
or U9701 (N_9701,N_9086,N_9353);
nor U9702 (N_9702,N_9417,N_9329);
or U9703 (N_9703,N_9457,N_9081);
and U9704 (N_9704,N_9449,N_9287);
nor U9705 (N_9705,N_9198,N_9052);
nor U9706 (N_9706,N_9482,N_9464);
xor U9707 (N_9707,N_9029,N_9469);
and U9708 (N_9708,N_9070,N_9323);
nand U9709 (N_9709,N_9267,N_9119);
nand U9710 (N_9710,N_9487,N_9339);
and U9711 (N_9711,N_9209,N_9179);
nor U9712 (N_9712,N_9296,N_9237);
and U9713 (N_9713,N_9450,N_9462);
or U9714 (N_9714,N_9341,N_9071);
nand U9715 (N_9715,N_9472,N_9008);
or U9716 (N_9716,N_9173,N_9333);
and U9717 (N_9717,N_9298,N_9343);
nor U9718 (N_9718,N_9220,N_9242);
xnor U9719 (N_9719,N_9397,N_9107);
or U9720 (N_9720,N_9085,N_9079);
xnor U9721 (N_9721,N_9266,N_9430);
nand U9722 (N_9722,N_9021,N_9188);
nand U9723 (N_9723,N_9447,N_9129);
and U9724 (N_9724,N_9184,N_9376);
xnor U9725 (N_9725,N_9478,N_9436);
or U9726 (N_9726,N_9475,N_9182);
xnor U9727 (N_9727,N_9219,N_9039);
nand U9728 (N_9728,N_9372,N_9238);
nand U9729 (N_9729,N_9113,N_9379);
and U9730 (N_9730,N_9097,N_9190);
and U9731 (N_9731,N_9360,N_9445);
or U9732 (N_9732,N_9471,N_9020);
nand U9733 (N_9733,N_9311,N_9394);
or U9734 (N_9734,N_9448,N_9354);
or U9735 (N_9735,N_9337,N_9069);
and U9736 (N_9736,N_9016,N_9441);
nor U9737 (N_9737,N_9046,N_9151);
xnor U9738 (N_9738,N_9102,N_9026);
nand U9739 (N_9739,N_9368,N_9455);
xnor U9740 (N_9740,N_9355,N_9254);
or U9741 (N_9741,N_9223,N_9174);
nor U9742 (N_9742,N_9408,N_9170);
xor U9743 (N_9743,N_9236,N_9465);
nor U9744 (N_9744,N_9261,N_9048);
nor U9745 (N_9745,N_9288,N_9481);
or U9746 (N_9746,N_9435,N_9050);
xor U9747 (N_9747,N_9414,N_9068);
nand U9748 (N_9748,N_9373,N_9270);
nor U9749 (N_9749,N_9421,N_9247);
nand U9750 (N_9750,N_9302,N_9339);
xnor U9751 (N_9751,N_9262,N_9466);
xnor U9752 (N_9752,N_9085,N_9212);
nor U9753 (N_9753,N_9069,N_9175);
or U9754 (N_9754,N_9303,N_9365);
xor U9755 (N_9755,N_9322,N_9478);
nor U9756 (N_9756,N_9203,N_9137);
xnor U9757 (N_9757,N_9490,N_9101);
nand U9758 (N_9758,N_9385,N_9311);
nand U9759 (N_9759,N_9127,N_9465);
and U9760 (N_9760,N_9318,N_9219);
or U9761 (N_9761,N_9301,N_9326);
and U9762 (N_9762,N_9013,N_9457);
and U9763 (N_9763,N_9401,N_9499);
nand U9764 (N_9764,N_9123,N_9053);
xnor U9765 (N_9765,N_9102,N_9036);
and U9766 (N_9766,N_9172,N_9155);
xor U9767 (N_9767,N_9337,N_9432);
nand U9768 (N_9768,N_9092,N_9164);
nand U9769 (N_9769,N_9129,N_9336);
and U9770 (N_9770,N_9431,N_9194);
xnor U9771 (N_9771,N_9040,N_9260);
nor U9772 (N_9772,N_9149,N_9493);
nand U9773 (N_9773,N_9093,N_9333);
xnor U9774 (N_9774,N_9155,N_9179);
or U9775 (N_9775,N_9223,N_9287);
or U9776 (N_9776,N_9285,N_9258);
nor U9777 (N_9777,N_9269,N_9126);
and U9778 (N_9778,N_9123,N_9310);
and U9779 (N_9779,N_9105,N_9487);
nor U9780 (N_9780,N_9142,N_9196);
xnor U9781 (N_9781,N_9395,N_9237);
nand U9782 (N_9782,N_9041,N_9155);
and U9783 (N_9783,N_9164,N_9465);
nand U9784 (N_9784,N_9103,N_9350);
and U9785 (N_9785,N_9049,N_9080);
xor U9786 (N_9786,N_9280,N_9265);
nor U9787 (N_9787,N_9285,N_9455);
nand U9788 (N_9788,N_9300,N_9431);
xnor U9789 (N_9789,N_9180,N_9219);
and U9790 (N_9790,N_9462,N_9142);
or U9791 (N_9791,N_9088,N_9129);
and U9792 (N_9792,N_9331,N_9304);
xor U9793 (N_9793,N_9303,N_9128);
xnor U9794 (N_9794,N_9145,N_9075);
nand U9795 (N_9795,N_9493,N_9119);
or U9796 (N_9796,N_9065,N_9347);
or U9797 (N_9797,N_9472,N_9387);
nand U9798 (N_9798,N_9121,N_9136);
xor U9799 (N_9799,N_9377,N_9461);
and U9800 (N_9800,N_9478,N_9376);
or U9801 (N_9801,N_9026,N_9198);
or U9802 (N_9802,N_9295,N_9385);
xor U9803 (N_9803,N_9423,N_9425);
nand U9804 (N_9804,N_9384,N_9203);
nor U9805 (N_9805,N_9423,N_9356);
or U9806 (N_9806,N_9073,N_9041);
nor U9807 (N_9807,N_9492,N_9260);
xor U9808 (N_9808,N_9058,N_9246);
nor U9809 (N_9809,N_9078,N_9488);
and U9810 (N_9810,N_9449,N_9496);
nor U9811 (N_9811,N_9261,N_9398);
xor U9812 (N_9812,N_9478,N_9307);
or U9813 (N_9813,N_9284,N_9364);
nand U9814 (N_9814,N_9348,N_9181);
and U9815 (N_9815,N_9388,N_9274);
xor U9816 (N_9816,N_9009,N_9112);
xnor U9817 (N_9817,N_9234,N_9448);
or U9818 (N_9818,N_9494,N_9259);
or U9819 (N_9819,N_9055,N_9197);
nor U9820 (N_9820,N_9345,N_9241);
or U9821 (N_9821,N_9340,N_9099);
nand U9822 (N_9822,N_9350,N_9090);
or U9823 (N_9823,N_9404,N_9430);
nand U9824 (N_9824,N_9470,N_9219);
and U9825 (N_9825,N_9071,N_9301);
or U9826 (N_9826,N_9263,N_9383);
nand U9827 (N_9827,N_9476,N_9318);
xor U9828 (N_9828,N_9102,N_9316);
and U9829 (N_9829,N_9136,N_9466);
nand U9830 (N_9830,N_9122,N_9193);
nand U9831 (N_9831,N_9307,N_9084);
nand U9832 (N_9832,N_9191,N_9019);
and U9833 (N_9833,N_9468,N_9248);
nand U9834 (N_9834,N_9400,N_9394);
xor U9835 (N_9835,N_9494,N_9190);
or U9836 (N_9836,N_9385,N_9461);
nand U9837 (N_9837,N_9033,N_9252);
or U9838 (N_9838,N_9010,N_9101);
nand U9839 (N_9839,N_9262,N_9235);
or U9840 (N_9840,N_9138,N_9483);
nand U9841 (N_9841,N_9039,N_9464);
xnor U9842 (N_9842,N_9320,N_9034);
nand U9843 (N_9843,N_9144,N_9188);
and U9844 (N_9844,N_9207,N_9197);
and U9845 (N_9845,N_9433,N_9148);
xor U9846 (N_9846,N_9254,N_9139);
nand U9847 (N_9847,N_9483,N_9440);
nand U9848 (N_9848,N_9316,N_9416);
xor U9849 (N_9849,N_9214,N_9088);
and U9850 (N_9850,N_9417,N_9126);
and U9851 (N_9851,N_9461,N_9116);
or U9852 (N_9852,N_9307,N_9107);
or U9853 (N_9853,N_9257,N_9038);
nand U9854 (N_9854,N_9253,N_9024);
xnor U9855 (N_9855,N_9117,N_9172);
nand U9856 (N_9856,N_9078,N_9271);
nor U9857 (N_9857,N_9411,N_9063);
and U9858 (N_9858,N_9482,N_9132);
xnor U9859 (N_9859,N_9253,N_9363);
xnor U9860 (N_9860,N_9478,N_9480);
xnor U9861 (N_9861,N_9073,N_9430);
and U9862 (N_9862,N_9188,N_9321);
xnor U9863 (N_9863,N_9001,N_9112);
xor U9864 (N_9864,N_9438,N_9050);
nand U9865 (N_9865,N_9163,N_9091);
nand U9866 (N_9866,N_9052,N_9083);
nor U9867 (N_9867,N_9325,N_9081);
or U9868 (N_9868,N_9246,N_9111);
nand U9869 (N_9869,N_9088,N_9055);
and U9870 (N_9870,N_9265,N_9368);
and U9871 (N_9871,N_9108,N_9004);
nand U9872 (N_9872,N_9148,N_9337);
nor U9873 (N_9873,N_9313,N_9067);
or U9874 (N_9874,N_9221,N_9259);
or U9875 (N_9875,N_9122,N_9009);
or U9876 (N_9876,N_9436,N_9447);
nor U9877 (N_9877,N_9246,N_9273);
xor U9878 (N_9878,N_9017,N_9444);
nor U9879 (N_9879,N_9493,N_9379);
nor U9880 (N_9880,N_9361,N_9127);
or U9881 (N_9881,N_9117,N_9022);
xor U9882 (N_9882,N_9133,N_9233);
or U9883 (N_9883,N_9484,N_9408);
nand U9884 (N_9884,N_9476,N_9089);
and U9885 (N_9885,N_9127,N_9259);
nand U9886 (N_9886,N_9296,N_9031);
and U9887 (N_9887,N_9265,N_9376);
or U9888 (N_9888,N_9462,N_9488);
xor U9889 (N_9889,N_9081,N_9342);
and U9890 (N_9890,N_9144,N_9171);
nor U9891 (N_9891,N_9340,N_9438);
and U9892 (N_9892,N_9164,N_9037);
xnor U9893 (N_9893,N_9359,N_9363);
nand U9894 (N_9894,N_9468,N_9357);
nor U9895 (N_9895,N_9068,N_9436);
and U9896 (N_9896,N_9145,N_9061);
nor U9897 (N_9897,N_9040,N_9167);
nor U9898 (N_9898,N_9269,N_9423);
or U9899 (N_9899,N_9075,N_9019);
and U9900 (N_9900,N_9144,N_9332);
nor U9901 (N_9901,N_9374,N_9426);
xor U9902 (N_9902,N_9042,N_9314);
or U9903 (N_9903,N_9186,N_9042);
nand U9904 (N_9904,N_9136,N_9325);
or U9905 (N_9905,N_9127,N_9464);
and U9906 (N_9906,N_9340,N_9168);
nor U9907 (N_9907,N_9172,N_9075);
xor U9908 (N_9908,N_9488,N_9371);
nand U9909 (N_9909,N_9336,N_9170);
or U9910 (N_9910,N_9164,N_9314);
and U9911 (N_9911,N_9161,N_9099);
or U9912 (N_9912,N_9168,N_9484);
and U9913 (N_9913,N_9376,N_9042);
or U9914 (N_9914,N_9366,N_9192);
xor U9915 (N_9915,N_9279,N_9336);
and U9916 (N_9916,N_9002,N_9208);
nand U9917 (N_9917,N_9347,N_9031);
nand U9918 (N_9918,N_9295,N_9459);
nor U9919 (N_9919,N_9002,N_9468);
or U9920 (N_9920,N_9150,N_9138);
or U9921 (N_9921,N_9462,N_9329);
nor U9922 (N_9922,N_9402,N_9232);
nand U9923 (N_9923,N_9456,N_9287);
nor U9924 (N_9924,N_9351,N_9342);
nand U9925 (N_9925,N_9187,N_9280);
nand U9926 (N_9926,N_9075,N_9052);
and U9927 (N_9927,N_9299,N_9246);
nor U9928 (N_9928,N_9147,N_9482);
nor U9929 (N_9929,N_9286,N_9264);
nand U9930 (N_9930,N_9201,N_9428);
nand U9931 (N_9931,N_9332,N_9283);
and U9932 (N_9932,N_9056,N_9095);
and U9933 (N_9933,N_9401,N_9303);
or U9934 (N_9934,N_9163,N_9422);
or U9935 (N_9935,N_9211,N_9294);
or U9936 (N_9936,N_9069,N_9290);
nand U9937 (N_9937,N_9344,N_9389);
xnor U9938 (N_9938,N_9032,N_9172);
nor U9939 (N_9939,N_9087,N_9235);
and U9940 (N_9940,N_9432,N_9029);
nand U9941 (N_9941,N_9019,N_9228);
nand U9942 (N_9942,N_9022,N_9398);
nor U9943 (N_9943,N_9209,N_9460);
or U9944 (N_9944,N_9415,N_9062);
nor U9945 (N_9945,N_9423,N_9498);
xnor U9946 (N_9946,N_9055,N_9151);
nand U9947 (N_9947,N_9025,N_9189);
or U9948 (N_9948,N_9164,N_9040);
nand U9949 (N_9949,N_9082,N_9090);
xnor U9950 (N_9950,N_9118,N_9177);
or U9951 (N_9951,N_9396,N_9221);
xor U9952 (N_9952,N_9371,N_9081);
xnor U9953 (N_9953,N_9212,N_9434);
nor U9954 (N_9954,N_9096,N_9278);
and U9955 (N_9955,N_9107,N_9304);
nand U9956 (N_9956,N_9136,N_9102);
xnor U9957 (N_9957,N_9199,N_9448);
or U9958 (N_9958,N_9063,N_9208);
xnor U9959 (N_9959,N_9121,N_9487);
and U9960 (N_9960,N_9322,N_9030);
and U9961 (N_9961,N_9200,N_9434);
nor U9962 (N_9962,N_9278,N_9050);
xnor U9963 (N_9963,N_9117,N_9331);
xnor U9964 (N_9964,N_9474,N_9001);
nor U9965 (N_9965,N_9112,N_9127);
nand U9966 (N_9966,N_9213,N_9151);
nor U9967 (N_9967,N_9399,N_9325);
and U9968 (N_9968,N_9034,N_9161);
nor U9969 (N_9969,N_9220,N_9194);
nand U9970 (N_9970,N_9382,N_9459);
nor U9971 (N_9971,N_9184,N_9303);
or U9972 (N_9972,N_9031,N_9167);
and U9973 (N_9973,N_9490,N_9189);
and U9974 (N_9974,N_9227,N_9148);
nor U9975 (N_9975,N_9068,N_9381);
nor U9976 (N_9976,N_9408,N_9177);
nor U9977 (N_9977,N_9320,N_9127);
nor U9978 (N_9978,N_9142,N_9333);
or U9979 (N_9979,N_9429,N_9478);
xor U9980 (N_9980,N_9465,N_9388);
nand U9981 (N_9981,N_9407,N_9458);
nor U9982 (N_9982,N_9188,N_9200);
xnor U9983 (N_9983,N_9172,N_9329);
and U9984 (N_9984,N_9145,N_9367);
nor U9985 (N_9985,N_9449,N_9373);
nor U9986 (N_9986,N_9028,N_9387);
xor U9987 (N_9987,N_9277,N_9242);
and U9988 (N_9988,N_9274,N_9438);
or U9989 (N_9989,N_9090,N_9105);
nor U9990 (N_9990,N_9185,N_9168);
nand U9991 (N_9991,N_9180,N_9001);
and U9992 (N_9992,N_9033,N_9421);
nand U9993 (N_9993,N_9163,N_9027);
nor U9994 (N_9994,N_9042,N_9230);
and U9995 (N_9995,N_9375,N_9404);
xor U9996 (N_9996,N_9448,N_9425);
xnor U9997 (N_9997,N_9176,N_9081);
or U9998 (N_9998,N_9474,N_9044);
nand U9999 (N_9999,N_9084,N_9377);
nor U10000 (N_10000,N_9985,N_9755);
nor U10001 (N_10001,N_9927,N_9775);
nand U10002 (N_10002,N_9915,N_9617);
nand U10003 (N_10003,N_9949,N_9627);
nor U10004 (N_10004,N_9631,N_9685);
xnor U10005 (N_10005,N_9901,N_9771);
xor U10006 (N_10006,N_9897,N_9858);
or U10007 (N_10007,N_9524,N_9651);
nor U10008 (N_10008,N_9522,N_9893);
nand U10009 (N_10009,N_9774,N_9788);
nand U10010 (N_10010,N_9963,N_9698);
nor U10011 (N_10011,N_9847,N_9970);
or U10012 (N_10012,N_9831,N_9916);
nor U10013 (N_10013,N_9909,N_9845);
xnor U10014 (N_10014,N_9607,N_9700);
and U10015 (N_10015,N_9853,N_9795);
and U10016 (N_10016,N_9641,N_9514);
nand U10017 (N_10017,N_9940,N_9951);
nand U10018 (N_10018,N_9792,N_9834);
xor U10019 (N_10019,N_9878,N_9835);
and U10020 (N_10020,N_9842,N_9529);
nand U10021 (N_10021,N_9681,N_9677);
nor U10022 (N_10022,N_9886,N_9604);
nand U10023 (N_10023,N_9948,N_9567);
xnor U10024 (N_10024,N_9768,N_9544);
and U10025 (N_10025,N_9862,N_9877);
or U10026 (N_10026,N_9563,N_9809);
nor U10027 (N_10027,N_9666,N_9959);
and U10028 (N_10028,N_9679,N_9982);
nand U10029 (N_10029,N_9599,N_9947);
nand U10030 (N_10030,N_9630,N_9532);
xnor U10031 (N_10031,N_9918,N_9872);
nor U10032 (N_10032,N_9787,N_9958);
nor U10033 (N_10033,N_9729,N_9518);
and U10034 (N_10034,N_9819,N_9707);
nand U10035 (N_10035,N_9600,N_9944);
nand U10036 (N_10036,N_9505,N_9924);
nand U10037 (N_10037,N_9705,N_9817);
nor U10038 (N_10038,N_9621,N_9742);
or U10039 (N_10039,N_9512,N_9682);
xnor U10040 (N_10040,N_9789,N_9608);
xnor U10041 (N_10041,N_9971,N_9715);
xor U10042 (N_10042,N_9805,N_9592);
and U10043 (N_10043,N_9815,N_9606);
xnor U10044 (N_10044,N_9989,N_9704);
nor U10045 (N_10045,N_9731,N_9688);
nand U10046 (N_10046,N_9937,N_9585);
nor U10047 (N_10047,N_9697,N_9867);
nand U10048 (N_10048,N_9968,N_9780);
nand U10049 (N_10049,N_9992,N_9902);
or U10050 (N_10050,N_9905,N_9808);
nor U10051 (N_10051,N_9501,N_9995);
or U10052 (N_10052,N_9786,N_9620);
or U10053 (N_10053,N_9781,N_9675);
and U10054 (N_10054,N_9738,N_9527);
xor U10055 (N_10055,N_9693,N_9706);
nor U10056 (N_10056,N_9748,N_9973);
nor U10057 (N_10057,N_9619,N_9578);
nand U10058 (N_10058,N_9943,N_9827);
nand U10059 (N_10059,N_9998,N_9660);
and U10060 (N_10060,N_9838,N_9588);
and U10061 (N_10061,N_9717,N_9868);
and U10062 (N_10062,N_9581,N_9587);
or U10063 (N_10063,N_9926,N_9637);
xnor U10064 (N_10064,N_9743,N_9644);
or U10065 (N_10065,N_9727,N_9560);
xnor U10066 (N_10066,N_9552,N_9804);
xor U10067 (N_10067,N_9938,N_9624);
and U10068 (N_10068,N_9903,N_9642);
nand U10069 (N_10069,N_9720,N_9674);
or U10070 (N_10070,N_9779,N_9852);
or U10071 (N_10071,N_9836,N_9987);
xor U10072 (N_10072,N_9952,N_9639);
xnor U10073 (N_10073,N_9713,N_9961);
xnor U10074 (N_10074,N_9823,N_9864);
xor U10075 (N_10075,N_9721,N_9718);
nand U10076 (N_10076,N_9690,N_9602);
or U10077 (N_10077,N_9668,N_9785);
nor U10078 (N_10078,N_9555,N_9672);
nor U10079 (N_10079,N_9507,N_9545);
or U10080 (N_10080,N_9671,N_9670);
nand U10081 (N_10081,N_9665,N_9647);
nand U10082 (N_10082,N_9692,N_9757);
or U10083 (N_10083,N_9974,N_9913);
nor U10084 (N_10084,N_9869,N_9571);
nand U10085 (N_10085,N_9582,N_9941);
nor U10086 (N_10086,N_9556,N_9843);
nor U10087 (N_10087,N_9699,N_9882);
nor U10088 (N_10088,N_9701,N_9596);
and U10089 (N_10089,N_9550,N_9984);
and U10090 (N_10090,N_9538,N_9508);
xor U10091 (N_10091,N_9841,N_9656);
and U10092 (N_10092,N_9859,N_9589);
xor U10093 (N_10093,N_9575,N_9509);
or U10094 (N_10094,N_9730,N_9954);
xor U10095 (N_10095,N_9816,N_9760);
and U10096 (N_10096,N_9623,N_9603);
nor U10097 (N_10097,N_9521,N_9871);
nand U10098 (N_10098,N_9914,N_9939);
nand U10099 (N_10099,N_9653,N_9540);
nor U10100 (N_10100,N_9646,N_9504);
nor U10101 (N_10101,N_9648,N_9999);
nor U10102 (N_10102,N_9908,N_9626);
nand U10103 (N_10103,N_9917,N_9863);
and U10104 (N_10104,N_9751,N_9813);
xnor U10105 (N_10105,N_9541,N_9519);
xnor U10106 (N_10106,N_9680,N_9702);
nand U10107 (N_10107,N_9513,N_9900);
nor U10108 (N_10108,N_9942,N_9810);
xor U10109 (N_10109,N_9752,N_9851);
nand U10110 (N_10110,N_9764,N_9754);
xnor U10111 (N_10111,N_9737,N_9605);
and U10112 (N_10112,N_9733,N_9956);
nor U10113 (N_10113,N_9534,N_9573);
xor U10114 (N_10114,N_9708,N_9734);
and U10115 (N_10115,N_9977,N_9802);
xnor U10116 (N_10116,N_9911,N_9611);
and U10117 (N_10117,N_9561,N_9723);
or U10118 (N_10118,N_9655,N_9500);
xor U10119 (N_10119,N_9662,N_9857);
nand U10120 (N_10120,N_9981,N_9874);
xor U10121 (N_10121,N_9988,N_9687);
or U10122 (N_10122,N_9866,N_9628);
nand U10123 (N_10123,N_9722,N_9579);
or U10124 (N_10124,N_9828,N_9849);
or U10125 (N_10125,N_9770,N_9996);
and U10126 (N_10126,N_9844,N_9983);
or U10127 (N_10127,N_9664,N_9576);
xnor U10128 (N_10128,N_9846,N_9972);
and U10129 (N_10129,N_9568,N_9549);
nor U10130 (N_10130,N_9881,N_9837);
nor U10131 (N_10131,N_9962,N_9965);
nand U10132 (N_10132,N_9833,N_9726);
nor U10133 (N_10133,N_9643,N_9750);
nand U10134 (N_10134,N_9526,N_9691);
nor U10135 (N_10135,N_9953,N_9811);
and U10136 (N_10136,N_9920,N_9800);
xnor U10137 (N_10137,N_9840,N_9669);
nor U10138 (N_10138,N_9537,N_9612);
nand U10139 (N_10139,N_9758,N_9906);
or U10140 (N_10140,N_9898,N_9883);
or U10141 (N_10141,N_9543,N_9856);
xnor U10142 (N_10142,N_9976,N_9967);
or U10143 (N_10143,N_9632,N_9885);
nor U10144 (N_10144,N_9986,N_9551);
nor U10145 (N_10145,N_9876,N_9930);
nor U10146 (N_10146,N_9638,N_9601);
nor U10147 (N_10147,N_9732,N_9564);
nor U10148 (N_10148,N_9523,N_9772);
xor U10149 (N_10149,N_9583,N_9546);
and U10150 (N_10150,N_9610,N_9899);
or U10151 (N_10151,N_9525,N_9855);
and U10152 (N_10152,N_9889,N_9574);
nand U10153 (N_10153,N_9714,N_9661);
or U10154 (N_10154,N_9929,N_9761);
xor U10155 (N_10155,N_9812,N_9746);
xor U10156 (N_10156,N_9654,N_9773);
or U10157 (N_10157,N_9609,N_9783);
xor U10158 (N_10158,N_9892,N_9839);
and U10159 (N_10159,N_9895,N_9650);
nor U10160 (N_10160,N_9594,N_9558);
xnor U10161 (N_10161,N_9794,N_9659);
or U10162 (N_10162,N_9736,N_9689);
nand U10163 (N_10163,N_9910,N_9991);
or U10164 (N_10164,N_9536,N_9584);
nand U10165 (N_10165,N_9934,N_9622);
xor U10166 (N_10166,N_9873,N_9921);
nand U10167 (N_10167,N_9801,N_9645);
or U10168 (N_10168,N_9784,N_9957);
nor U10169 (N_10169,N_9511,N_9888);
xor U10170 (N_10170,N_9912,N_9932);
or U10171 (N_10171,N_9814,N_9649);
nor U10172 (N_10172,N_9880,N_9562);
xnor U10173 (N_10173,N_9826,N_9928);
and U10174 (N_10174,N_9535,N_9667);
or U10175 (N_10175,N_9925,N_9894);
nor U10176 (N_10176,N_9745,N_9753);
nor U10177 (N_10177,N_9955,N_9678);
nand U10178 (N_10178,N_9572,N_9547);
nand U10179 (N_10179,N_9975,N_9739);
xor U10180 (N_10180,N_9791,N_9799);
or U10181 (N_10181,N_9598,N_9591);
nor U10182 (N_10182,N_9663,N_9502);
nand U10183 (N_10183,N_9553,N_9740);
xnor U10184 (N_10184,N_9728,N_9636);
nand U10185 (N_10185,N_9747,N_9586);
xnor U10186 (N_10186,N_9597,N_9767);
or U10187 (N_10187,N_9884,N_9593);
xnor U10188 (N_10188,N_9520,N_9694);
or U10189 (N_10189,N_9506,N_9798);
nand U10190 (N_10190,N_9763,N_9990);
xor U10191 (N_10191,N_9533,N_9635);
xnor U10192 (N_10192,N_9861,N_9559);
and U10193 (N_10193,N_9933,N_9807);
or U10194 (N_10194,N_9539,N_9615);
or U10195 (N_10195,N_9935,N_9633);
and U10196 (N_10196,N_9709,N_9565);
xnor U10197 (N_10197,N_9832,N_9516);
or U10198 (N_10198,N_9825,N_9616);
nand U10199 (N_10199,N_9657,N_9820);
or U10200 (N_10200,N_9821,N_9640);
or U10201 (N_10201,N_9629,N_9580);
xnor U10202 (N_10202,N_9950,N_9945);
or U10203 (N_10203,N_9614,N_9830);
xnor U10204 (N_10204,N_9725,N_9960);
or U10205 (N_10205,N_9756,N_9759);
xnor U10206 (N_10206,N_9946,N_9696);
and U10207 (N_10207,N_9854,N_9969);
and U10208 (N_10208,N_9936,N_9793);
nand U10209 (N_10209,N_9964,N_9978);
nand U10210 (N_10210,N_9618,N_9676);
nand U10211 (N_10211,N_9762,N_9890);
and U10212 (N_10212,N_9530,N_9870);
and U10213 (N_10213,N_9776,N_9879);
or U10214 (N_10214,N_9510,N_9684);
nor U10215 (N_10215,N_9577,N_9503);
nand U10216 (N_10216,N_9904,N_9848);
xnor U10217 (N_10217,N_9818,N_9922);
nand U10218 (N_10218,N_9769,N_9796);
or U10219 (N_10219,N_9994,N_9860);
nand U10220 (N_10220,N_9531,N_9744);
xor U10221 (N_10221,N_9517,N_9797);
nor U10222 (N_10222,N_9735,N_9778);
xor U10223 (N_10223,N_9790,N_9806);
and U10224 (N_10224,N_9570,N_9703);
or U10225 (N_10225,N_9528,N_9822);
nand U10226 (N_10226,N_9658,N_9875);
or U10227 (N_10227,N_9931,N_9686);
nand U10228 (N_10228,N_9966,N_9741);
nand U10229 (N_10229,N_9907,N_9766);
nor U10230 (N_10230,N_9993,N_9652);
nand U10231 (N_10231,N_9765,N_9782);
and U10232 (N_10232,N_9896,N_9569);
nor U10233 (N_10233,N_9548,N_9613);
or U10234 (N_10234,N_9712,N_9542);
and U10235 (N_10235,N_9590,N_9829);
or U10236 (N_10236,N_9980,N_9557);
xor U10237 (N_10237,N_9683,N_9850);
and U10238 (N_10238,N_9710,N_9566);
or U10239 (N_10239,N_9887,N_9595);
and U10240 (N_10240,N_9997,N_9625);
nand U10241 (N_10241,N_9515,N_9979);
nand U10242 (N_10242,N_9923,N_9719);
and U10243 (N_10243,N_9749,N_9554);
xnor U10244 (N_10244,N_9634,N_9891);
xnor U10245 (N_10245,N_9695,N_9865);
nor U10246 (N_10246,N_9716,N_9673);
nand U10247 (N_10247,N_9724,N_9777);
and U10248 (N_10248,N_9824,N_9919);
or U10249 (N_10249,N_9803,N_9711);
nand U10250 (N_10250,N_9609,N_9678);
or U10251 (N_10251,N_9692,N_9931);
xnor U10252 (N_10252,N_9704,N_9556);
or U10253 (N_10253,N_9540,N_9752);
xnor U10254 (N_10254,N_9558,N_9792);
xnor U10255 (N_10255,N_9941,N_9750);
nand U10256 (N_10256,N_9903,N_9725);
xor U10257 (N_10257,N_9629,N_9670);
xnor U10258 (N_10258,N_9595,N_9894);
nor U10259 (N_10259,N_9938,N_9976);
and U10260 (N_10260,N_9671,N_9892);
nand U10261 (N_10261,N_9947,N_9741);
nor U10262 (N_10262,N_9756,N_9637);
nand U10263 (N_10263,N_9897,N_9809);
nor U10264 (N_10264,N_9546,N_9609);
nand U10265 (N_10265,N_9969,N_9580);
xnor U10266 (N_10266,N_9622,N_9583);
or U10267 (N_10267,N_9651,N_9919);
and U10268 (N_10268,N_9523,N_9980);
or U10269 (N_10269,N_9969,N_9809);
and U10270 (N_10270,N_9520,N_9644);
or U10271 (N_10271,N_9886,N_9832);
nor U10272 (N_10272,N_9555,N_9512);
xor U10273 (N_10273,N_9588,N_9735);
and U10274 (N_10274,N_9660,N_9618);
or U10275 (N_10275,N_9874,N_9557);
nand U10276 (N_10276,N_9658,N_9964);
xnor U10277 (N_10277,N_9705,N_9629);
or U10278 (N_10278,N_9582,N_9874);
nor U10279 (N_10279,N_9920,N_9587);
nor U10280 (N_10280,N_9834,N_9896);
and U10281 (N_10281,N_9853,N_9537);
or U10282 (N_10282,N_9750,N_9817);
nand U10283 (N_10283,N_9828,N_9580);
nand U10284 (N_10284,N_9531,N_9765);
or U10285 (N_10285,N_9516,N_9787);
nor U10286 (N_10286,N_9526,N_9523);
nor U10287 (N_10287,N_9527,N_9590);
and U10288 (N_10288,N_9564,N_9740);
or U10289 (N_10289,N_9891,N_9754);
and U10290 (N_10290,N_9841,N_9653);
nor U10291 (N_10291,N_9915,N_9673);
and U10292 (N_10292,N_9936,N_9807);
xor U10293 (N_10293,N_9609,N_9605);
nor U10294 (N_10294,N_9743,N_9960);
or U10295 (N_10295,N_9939,N_9514);
nand U10296 (N_10296,N_9785,N_9821);
and U10297 (N_10297,N_9631,N_9848);
nand U10298 (N_10298,N_9851,N_9592);
xor U10299 (N_10299,N_9855,N_9619);
or U10300 (N_10300,N_9896,N_9890);
xnor U10301 (N_10301,N_9592,N_9524);
and U10302 (N_10302,N_9554,N_9861);
or U10303 (N_10303,N_9792,N_9718);
and U10304 (N_10304,N_9939,N_9980);
nor U10305 (N_10305,N_9985,N_9735);
nand U10306 (N_10306,N_9966,N_9982);
xnor U10307 (N_10307,N_9529,N_9909);
and U10308 (N_10308,N_9611,N_9969);
xor U10309 (N_10309,N_9820,N_9689);
or U10310 (N_10310,N_9994,N_9713);
nand U10311 (N_10311,N_9618,N_9828);
nand U10312 (N_10312,N_9795,N_9978);
nor U10313 (N_10313,N_9838,N_9560);
and U10314 (N_10314,N_9745,N_9875);
xnor U10315 (N_10315,N_9934,N_9554);
or U10316 (N_10316,N_9916,N_9702);
nand U10317 (N_10317,N_9652,N_9789);
and U10318 (N_10318,N_9580,N_9842);
xnor U10319 (N_10319,N_9692,N_9844);
xor U10320 (N_10320,N_9838,N_9815);
xor U10321 (N_10321,N_9845,N_9501);
xnor U10322 (N_10322,N_9501,N_9947);
nand U10323 (N_10323,N_9764,N_9526);
xnor U10324 (N_10324,N_9725,N_9729);
nor U10325 (N_10325,N_9815,N_9787);
and U10326 (N_10326,N_9811,N_9894);
and U10327 (N_10327,N_9637,N_9621);
xnor U10328 (N_10328,N_9968,N_9538);
and U10329 (N_10329,N_9749,N_9744);
nand U10330 (N_10330,N_9910,N_9770);
and U10331 (N_10331,N_9662,N_9546);
nor U10332 (N_10332,N_9971,N_9722);
nand U10333 (N_10333,N_9664,N_9786);
nor U10334 (N_10334,N_9883,N_9597);
or U10335 (N_10335,N_9561,N_9864);
xor U10336 (N_10336,N_9644,N_9715);
or U10337 (N_10337,N_9746,N_9713);
or U10338 (N_10338,N_9692,N_9952);
nand U10339 (N_10339,N_9670,N_9935);
and U10340 (N_10340,N_9521,N_9893);
xor U10341 (N_10341,N_9816,N_9792);
nand U10342 (N_10342,N_9763,N_9516);
nor U10343 (N_10343,N_9510,N_9749);
nor U10344 (N_10344,N_9964,N_9914);
nor U10345 (N_10345,N_9809,N_9566);
or U10346 (N_10346,N_9876,N_9789);
or U10347 (N_10347,N_9974,N_9761);
nor U10348 (N_10348,N_9505,N_9798);
nand U10349 (N_10349,N_9855,N_9891);
or U10350 (N_10350,N_9778,N_9695);
and U10351 (N_10351,N_9540,N_9753);
nor U10352 (N_10352,N_9956,N_9981);
nand U10353 (N_10353,N_9539,N_9880);
or U10354 (N_10354,N_9674,N_9781);
or U10355 (N_10355,N_9889,N_9939);
or U10356 (N_10356,N_9891,N_9888);
or U10357 (N_10357,N_9545,N_9535);
nand U10358 (N_10358,N_9710,N_9968);
or U10359 (N_10359,N_9632,N_9624);
or U10360 (N_10360,N_9743,N_9886);
xnor U10361 (N_10361,N_9732,N_9859);
xor U10362 (N_10362,N_9535,N_9528);
or U10363 (N_10363,N_9823,N_9910);
nand U10364 (N_10364,N_9846,N_9876);
xnor U10365 (N_10365,N_9760,N_9947);
nor U10366 (N_10366,N_9551,N_9949);
or U10367 (N_10367,N_9541,N_9934);
nor U10368 (N_10368,N_9879,N_9538);
xor U10369 (N_10369,N_9728,N_9530);
nand U10370 (N_10370,N_9896,N_9615);
and U10371 (N_10371,N_9529,N_9512);
and U10372 (N_10372,N_9891,N_9951);
and U10373 (N_10373,N_9664,N_9785);
nand U10374 (N_10374,N_9662,N_9514);
xor U10375 (N_10375,N_9732,N_9974);
nand U10376 (N_10376,N_9956,N_9716);
and U10377 (N_10377,N_9757,N_9714);
nor U10378 (N_10378,N_9746,N_9591);
nor U10379 (N_10379,N_9728,N_9755);
or U10380 (N_10380,N_9507,N_9622);
nand U10381 (N_10381,N_9760,N_9998);
or U10382 (N_10382,N_9658,N_9695);
or U10383 (N_10383,N_9972,N_9608);
nor U10384 (N_10384,N_9818,N_9976);
and U10385 (N_10385,N_9957,N_9682);
nor U10386 (N_10386,N_9964,N_9984);
or U10387 (N_10387,N_9681,N_9693);
or U10388 (N_10388,N_9746,N_9936);
nand U10389 (N_10389,N_9799,N_9794);
xor U10390 (N_10390,N_9951,N_9826);
or U10391 (N_10391,N_9655,N_9833);
nor U10392 (N_10392,N_9839,N_9521);
or U10393 (N_10393,N_9577,N_9895);
and U10394 (N_10394,N_9924,N_9785);
nand U10395 (N_10395,N_9555,N_9621);
nor U10396 (N_10396,N_9675,N_9847);
xnor U10397 (N_10397,N_9962,N_9745);
and U10398 (N_10398,N_9711,N_9549);
nand U10399 (N_10399,N_9700,N_9781);
nand U10400 (N_10400,N_9635,N_9768);
and U10401 (N_10401,N_9634,N_9585);
or U10402 (N_10402,N_9800,N_9877);
xor U10403 (N_10403,N_9551,N_9743);
xor U10404 (N_10404,N_9813,N_9551);
or U10405 (N_10405,N_9584,N_9766);
nand U10406 (N_10406,N_9652,N_9691);
and U10407 (N_10407,N_9550,N_9830);
nand U10408 (N_10408,N_9559,N_9968);
or U10409 (N_10409,N_9926,N_9652);
nand U10410 (N_10410,N_9602,N_9713);
nor U10411 (N_10411,N_9502,N_9920);
nand U10412 (N_10412,N_9617,N_9710);
nand U10413 (N_10413,N_9880,N_9695);
or U10414 (N_10414,N_9763,N_9525);
nand U10415 (N_10415,N_9784,N_9572);
nor U10416 (N_10416,N_9881,N_9703);
or U10417 (N_10417,N_9542,N_9696);
or U10418 (N_10418,N_9759,N_9927);
nor U10419 (N_10419,N_9534,N_9730);
xor U10420 (N_10420,N_9740,N_9691);
nor U10421 (N_10421,N_9626,N_9761);
or U10422 (N_10422,N_9993,N_9939);
nor U10423 (N_10423,N_9970,N_9504);
nand U10424 (N_10424,N_9622,N_9516);
or U10425 (N_10425,N_9568,N_9786);
and U10426 (N_10426,N_9782,N_9763);
nand U10427 (N_10427,N_9933,N_9844);
xnor U10428 (N_10428,N_9814,N_9523);
and U10429 (N_10429,N_9835,N_9561);
xnor U10430 (N_10430,N_9866,N_9665);
nand U10431 (N_10431,N_9712,N_9901);
and U10432 (N_10432,N_9668,N_9661);
and U10433 (N_10433,N_9621,N_9901);
xor U10434 (N_10434,N_9693,N_9914);
xor U10435 (N_10435,N_9718,N_9787);
nand U10436 (N_10436,N_9628,N_9578);
xnor U10437 (N_10437,N_9729,N_9766);
nand U10438 (N_10438,N_9915,N_9713);
nor U10439 (N_10439,N_9953,N_9565);
nand U10440 (N_10440,N_9530,N_9848);
xor U10441 (N_10441,N_9631,N_9966);
nand U10442 (N_10442,N_9887,N_9529);
or U10443 (N_10443,N_9819,N_9649);
or U10444 (N_10444,N_9950,N_9788);
xnor U10445 (N_10445,N_9918,N_9984);
nor U10446 (N_10446,N_9637,N_9690);
nand U10447 (N_10447,N_9557,N_9548);
nor U10448 (N_10448,N_9622,N_9867);
nand U10449 (N_10449,N_9903,N_9675);
nor U10450 (N_10450,N_9574,N_9508);
xnor U10451 (N_10451,N_9950,N_9563);
xnor U10452 (N_10452,N_9717,N_9576);
or U10453 (N_10453,N_9841,N_9508);
or U10454 (N_10454,N_9602,N_9889);
nand U10455 (N_10455,N_9949,N_9959);
xnor U10456 (N_10456,N_9525,N_9638);
and U10457 (N_10457,N_9837,N_9993);
nand U10458 (N_10458,N_9683,N_9785);
nand U10459 (N_10459,N_9840,N_9971);
nor U10460 (N_10460,N_9799,N_9682);
and U10461 (N_10461,N_9525,N_9543);
nor U10462 (N_10462,N_9625,N_9540);
or U10463 (N_10463,N_9533,N_9556);
nor U10464 (N_10464,N_9815,N_9564);
xnor U10465 (N_10465,N_9817,N_9584);
xor U10466 (N_10466,N_9967,N_9568);
nand U10467 (N_10467,N_9742,N_9617);
and U10468 (N_10468,N_9808,N_9546);
nor U10469 (N_10469,N_9955,N_9941);
and U10470 (N_10470,N_9611,N_9915);
and U10471 (N_10471,N_9635,N_9514);
and U10472 (N_10472,N_9532,N_9837);
xor U10473 (N_10473,N_9899,N_9923);
and U10474 (N_10474,N_9601,N_9538);
or U10475 (N_10475,N_9737,N_9634);
nor U10476 (N_10476,N_9972,N_9780);
nand U10477 (N_10477,N_9871,N_9921);
nand U10478 (N_10478,N_9507,N_9601);
or U10479 (N_10479,N_9896,N_9504);
nand U10480 (N_10480,N_9668,N_9609);
and U10481 (N_10481,N_9831,N_9976);
nor U10482 (N_10482,N_9802,N_9776);
nor U10483 (N_10483,N_9562,N_9672);
or U10484 (N_10484,N_9907,N_9540);
nor U10485 (N_10485,N_9843,N_9716);
or U10486 (N_10486,N_9541,N_9659);
nand U10487 (N_10487,N_9604,N_9769);
xor U10488 (N_10488,N_9542,N_9731);
xor U10489 (N_10489,N_9822,N_9717);
xnor U10490 (N_10490,N_9693,N_9763);
nor U10491 (N_10491,N_9710,N_9559);
and U10492 (N_10492,N_9841,N_9679);
nor U10493 (N_10493,N_9986,N_9925);
and U10494 (N_10494,N_9691,N_9570);
xor U10495 (N_10495,N_9699,N_9602);
or U10496 (N_10496,N_9874,N_9923);
xor U10497 (N_10497,N_9758,N_9676);
xor U10498 (N_10498,N_9773,N_9739);
nor U10499 (N_10499,N_9865,N_9962);
and U10500 (N_10500,N_10473,N_10177);
xor U10501 (N_10501,N_10434,N_10384);
nor U10502 (N_10502,N_10187,N_10356);
nand U10503 (N_10503,N_10368,N_10181);
nor U10504 (N_10504,N_10430,N_10084);
xor U10505 (N_10505,N_10426,N_10361);
nand U10506 (N_10506,N_10262,N_10245);
nand U10507 (N_10507,N_10333,N_10247);
or U10508 (N_10508,N_10485,N_10488);
nand U10509 (N_10509,N_10120,N_10387);
nor U10510 (N_10510,N_10355,N_10342);
xnor U10511 (N_10511,N_10271,N_10125);
and U10512 (N_10512,N_10311,N_10055);
xor U10513 (N_10513,N_10082,N_10281);
nor U10514 (N_10514,N_10135,N_10462);
or U10515 (N_10515,N_10119,N_10312);
and U10516 (N_10516,N_10284,N_10027);
nor U10517 (N_10517,N_10369,N_10464);
xnor U10518 (N_10518,N_10366,N_10447);
nor U10519 (N_10519,N_10225,N_10231);
and U10520 (N_10520,N_10171,N_10074);
and U10521 (N_10521,N_10413,N_10338);
and U10522 (N_10522,N_10063,N_10222);
nand U10523 (N_10523,N_10188,N_10388);
or U10524 (N_10524,N_10443,N_10374);
nor U10525 (N_10525,N_10010,N_10183);
nand U10526 (N_10526,N_10046,N_10307);
nor U10527 (N_10527,N_10427,N_10129);
nor U10528 (N_10528,N_10197,N_10062);
nand U10529 (N_10529,N_10180,N_10286);
nor U10530 (N_10530,N_10493,N_10498);
xnor U10531 (N_10531,N_10345,N_10399);
and U10532 (N_10532,N_10215,N_10480);
nor U10533 (N_10533,N_10034,N_10411);
xnor U10534 (N_10534,N_10377,N_10250);
and U10535 (N_10535,N_10386,N_10364);
or U10536 (N_10536,N_10373,N_10154);
nand U10537 (N_10537,N_10325,N_10344);
or U10538 (N_10538,N_10418,N_10398);
and U10539 (N_10539,N_10244,N_10168);
nor U10540 (N_10540,N_10172,N_10491);
or U10541 (N_10541,N_10270,N_10045);
nor U10542 (N_10542,N_10459,N_10436);
or U10543 (N_10543,N_10030,N_10152);
nor U10544 (N_10544,N_10007,N_10486);
xor U10545 (N_10545,N_10004,N_10446);
xnor U10546 (N_10546,N_10224,N_10107);
and U10547 (N_10547,N_10397,N_10132);
xor U10548 (N_10548,N_10448,N_10047);
xor U10549 (N_10549,N_10001,N_10256);
xor U10550 (N_10550,N_10263,N_10196);
xor U10551 (N_10551,N_10077,N_10020);
and U10552 (N_10552,N_10445,N_10349);
nand U10553 (N_10553,N_10415,N_10057);
nand U10554 (N_10554,N_10341,N_10309);
nor U10555 (N_10555,N_10011,N_10456);
nand U10556 (N_10556,N_10460,N_10463);
nor U10557 (N_10557,N_10461,N_10035);
or U10558 (N_10558,N_10064,N_10496);
nor U10559 (N_10559,N_10324,N_10381);
and U10560 (N_10560,N_10289,N_10218);
xor U10561 (N_10561,N_10482,N_10201);
nor U10562 (N_10562,N_10070,N_10216);
and U10563 (N_10563,N_10230,N_10126);
and U10564 (N_10564,N_10259,N_10008);
nand U10565 (N_10565,N_10412,N_10394);
or U10566 (N_10566,N_10149,N_10167);
or U10567 (N_10567,N_10232,N_10272);
nand U10568 (N_10568,N_10039,N_10053);
xor U10569 (N_10569,N_10058,N_10076);
or U10570 (N_10570,N_10127,N_10449);
nand U10571 (N_10571,N_10142,N_10300);
nand U10572 (N_10572,N_10110,N_10367);
nor U10573 (N_10573,N_10242,N_10475);
xnor U10574 (N_10574,N_10383,N_10274);
and U10575 (N_10575,N_10437,N_10200);
or U10576 (N_10576,N_10068,N_10229);
and U10577 (N_10577,N_10065,N_10465);
or U10578 (N_10578,N_10433,N_10357);
or U10579 (N_10579,N_10254,N_10321);
nor U10580 (N_10580,N_10371,N_10202);
nor U10581 (N_10581,N_10260,N_10292);
nand U10582 (N_10582,N_10117,N_10056);
or U10583 (N_10583,N_10170,N_10251);
or U10584 (N_10584,N_10164,N_10050);
xnor U10585 (N_10585,N_10269,N_10320);
nor U10586 (N_10586,N_10192,N_10100);
nor U10587 (N_10587,N_10490,N_10179);
and U10588 (N_10588,N_10089,N_10018);
and U10589 (N_10589,N_10479,N_10315);
xnor U10590 (N_10590,N_10078,N_10416);
nor U10591 (N_10591,N_10112,N_10489);
xor U10592 (N_10592,N_10305,N_10404);
nand U10593 (N_10593,N_10113,N_10067);
and U10594 (N_10594,N_10162,N_10212);
and U10595 (N_10595,N_10499,N_10441);
or U10596 (N_10596,N_10432,N_10478);
nor U10597 (N_10597,N_10024,N_10458);
xor U10598 (N_10598,N_10438,N_10417);
and U10599 (N_10599,N_10026,N_10086);
nand U10600 (N_10600,N_10348,N_10096);
xor U10601 (N_10601,N_10336,N_10114);
xor U10602 (N_10602,N_10198,N_10176);
or U10603 (N_10603,N_10214,N_10165);
nand U10604 (N_10604,N_10327,N_10104);
and U10605 (N_10605,N_10435,N_10028);
xnor U10606 (N_10606,N_10049,N_10331);
or U10607 (N_10607,N_10227,N_10283);
or U10608 (N_10608,N_10440,N_10032);
and U10609 (N_10609,N_10472,N_10267);
xnor U10610 (N_10610,N_10022,N_10444);
nor U10611 (N_10611,N_10081,N_10408);
xor U10612 (N_10612,N_10012,N_10234);
or U10613 (N_10613,N_10299,N_10091);
xnor U10614 (N_10614,N_10048,N_10407);
nor U10615 (N_10615,N_10005,N_10195);
nor U10616 (N_10616,N_10391,N_10352);
xor U10617 (N_10617,N_10173,N_10006);
nand U10618 (N_10618,N_10494,N_10487);
nand U10619 (N_10619,N_10332,N_10334);
nor U10620 (N_10620,N_10233,N_10221);
or U10621 (N_10621,N_10452,N_10092);
and U10622 (N_10622,N_10343,N_10296);
nand U10623 (N_10623,N_10451,N_10470);
and U10624 (N_10624,N_10380,N_10476);
nand U10625 (N_10625,N_10205,N_10157);
or U10626 (N_10626,N_10450,N_10239);
or U10627 (N_10627,N_10097,N_10279);
nor U10628 (N_10628,N_10322,N_10217);
and U10629 (N_10629,N_10278,N_10016);
nand U10630 (N_10630,N_10249,N_10087);
or U10631 (N_10631,N_10280,N_10042);
nand U10632 (N_10632,N_10191,N_10392);
nor U10633 (N_10633,N_10178,N_10040);
nor U10634 (N_10634,N_10453,N_10317);
nor U10635 (N_10635,N_10144,N_10358);
xor U10636 (N_10636,N_10423,N_10146);
or U10637 (N_10637,N_10354,N_10481);
or U10638 (N_10638,N_10137,N_10403);
or U10639 (N_10639,N_10109,N_10264);
nor U10640 (N_10640,N_10273,N_10454);
and U10641 (N_10641,N_10069,N_10308);
and U10642 (N_10642,N_10038,N_10013);
nor U10643 (N_10643,N_10306,N_10071);
xor U10644 (N_10644,N_10303,N_10455);
or U10645 (N_10645,N_10375,N_10497);
xor U10646 (N_10646,N_10253,N_10287);
nand U10647 (N_10647,N_10258,N_10031);
nand U10648 (N_10648,N_10036,N_10340);
nor U10649 (N_10649,N_10115,N_10052);
and U10650 (N_10650,N_10017,N_10277);
nand U10651 (N_10651,N_10099,N_10108);
nand U10652 (N_10652,N_10237,N_10166);
nand U10653 (N_10653,N_10106,N_10248);
nand U10654 (N_10654,N_10243,N_10484);
or U10655 (N_10655,N_10213,N_10169);
or U10656 (N_10656,N_10133,N_10098);
xnor U10657 (N_10657,N_10372,N_10138);
and U10658 (N_10658,N_10134,N_10326);
xnor U10659 (N_10659,N_10059,N_10429);
nand U10660 (N_10660,N_10301,N_10136);
or U10661 (N_10661,N_10468,N_10226);
and U10662 (N_10662,N_10147,N_10457);
nor U10663 (N_10663,N_10353,N_10095);
xor U10664 (N_10664,N_10153,N_10409);
or U10665 (N_10665,N_10379,N_10313);
xor U10666 (N_10666,N_10402,N_10376);
nand U10667 (N_10667,N_10405,N_10002);
and U10668 (N_10668,N_10335,N_10174);
xnor U10669 (N_10669,N_10240,N_10101);
and U10670 (N_10670,N_10420,N_10393);
nor U10671 (N_10671,N_10339,N_10290);
xor U10672 (N_10672,N_10206,N_10060);
nor U10673 (N_10673,N_10009,N_10298);
and U10674 (N_10674,N_10211,N_10186);
or U10675 (N_10675,N_10466,N_10037);
xnor U10676 (N_10676,N_10346,N_10370);
xor U10677 (N_10677,N_10093,N_10073);
nand U10678 (N_10678,N_10094,N_10439);
and U10679 (N_10679,N_10184,N_10130);
and U10680 (N_10680,N_10304,N_10246);
or U10681 (N_10681,N_10021,N_10351);
nor U10682 (N_10682,N_10257,N_10148);
nor U10683 (N_10683,N_10079,N_10156);
nand U10684 (N_10684,N_10185,N_10276);
xnor U10685 (N_10685,N_10421,N_10425);
or U10686 (N_10686,N_10123,N_10223);
nor U10687 (N_10687,N_10295,N_10401);
xnor U10688 (N_10688,N_10385,N_10314);
nor U10689 (N_10689,N_10467,N_10102);
and U10690 (N_10690,N_10143,N_10066);
and U10691 (N_10691,N_10328,N_10209);
nand U10692 (N_10692,N_10474,N_10075);
or U10693 (N_10693,N_10442,N_10406);
nor U10694 (N_10694,N_10139,N_10422);
and U10695 (N_10695,N_10318,N_10072);
or U10696 (N_10696,N_10360,N_10241);
and U10697 (N_10697,N_10302,N_10193);
nor U10698 (N_10698,N_10492,N_10033);
nor U10699 (N_10699,N_10061,N_10431);
xor U10700 (N_10700,N_10310,N_10359);
xnor U10701 (N_10701,N_10275,N_10396);
or U10702 (N_10702,N_10378,N_10235);
nor U10703 (N_10703,N_10203,N_10350);
nand U10704 (N_10704,N_10291,N_10228);
nand U10705 (N_10705,N_10323,N_10252);
nor U10706 (N_10706,N_10015,N_10190);
and U10707 (N_10707,N_10118,N_10051);
and U10708 (N_10708,N_10023,N_10189);
and U10709 (N_10709,N_10266,N_10151);
or U10710 (N_10710,N_10330,N_10207);
or U10711 (N_10711,N_10219,N_10199);
xnor U10712 (N_10712,N_10158,N_10141);
nor U10713 (N_10713,N_10477,N_10238);
nor U10714 (N_10714,N_10208,N_10365);
nor U10715 (N_10715,N_10090,N_10428);
nand U10716 (N_10716,N_10145,N_10210);
and U10717 (N_10717,N_10088,N_10105);
nand U10718 (N_10718,N_10161,N_10103);
nor U10719 (N_10719,N_10029,N_10410);
nor U10720 (N_10720,N_10194,N_10400);
or U10721 (N_10721,N_10204,N_10159);
or U10722 (N_10722,N_10182,N_10268);
or U10723 (N_10723,N_10085,N_10236);
nand U10724 (N_10724,N_10390,N_10414);
nand U10725 (N_10725,N_10319,N_10128);
xor U10726 (N_10726,N_10255,N_10175);
xor U10727 (N_10727,N_10261,N_10122);
nand U10728 (N_10728,N_10362,N_10155);
or U10729 (N_10729,N_10419,N_10337);
and U10730 (N_10730,N_10121,N_10288);
nor U10731 (N_10731,N_10471,N_10347);
nand U10732 (N_10732,N_10140,N_10054);
xnor U10733 (N_10733,N_10160,N_10163);
or U10734 (N_10734,N_10083,N_10363);
and U10735 (N_10735,N_10000,N_10395);
nor U10736 (N_10736,N_10080,N_10124);
xor U10737 (N_10737,N_10316,N_10297);
nand U10738 (N_10738,N_10282,N_10019);
xor U10739 (N_10739,N_10424,N_10469);
nand U10740 (N_10740,N_10265,N_10044);
nor U10741 (N_10741,N_10285,N_10329);
xor U10742 (N_10742,N_10131,N_10150);
nor U10743 (N_10743,N_10220,N_10389);
nand U10744 (N_10744,N_10014,N_10294);
and U10745 (N_10745,N_10116,N_10483);
xor U10746 (N_10746,N_10495,N_10382);
nor U10747 (N_10747,N_10043,N_10025);
xor U10748 (N_10748,N_10293,N_10003);
or U10749 (N_10749,N_10041,N_10111);
xor U10750 (N_10750,N_10179,N_10356);
xor U10751 (N_10751,N_10385,N_10128);
and U10752 (N_10752,N_10281,N_10127);
nand U10753 (N_10753,N_10496,N_10138);
nor U10754 (N_10754,N_10130,N_10087);
xor U10755 (N_10755,N_10341,N_10194);
nor U10756 (N_10756,N_10456,N_10450);
or U10757 (N_10757,N_10131,N_10424);
xnor U10758 (N_10758,N_10216,N_10439);
nor U10759 (N_10759,N_10352,N_10473);
or U10760 (N_10760,N_10143,N_10404);
or U10761 (N_10761,N_10336,N_10111);
xnor U10762 (N_10762,N_10400,N_10333);
nor U10763 (N_10763,N_10058,N_10063);
or U10764 (N_10764,N_10365,N_10142);
xor U10765 (N_10765,N_10442,N_10351);
or U10766 (N_10766,N_10208,N_10437);
nor U10767 (N_10767,N_10488,N_10281);
nand U10768 (N_10768,N_10327,N_10111);
xor U10769 (N_10769,N_10433,N_10228);
xor U10770 (N_10770,N_10029,N_10284);
nor U10771 (N_10771,N_10140,N_10431);
and U10772 (N_10772,N_10325,N_10195);
or U10773 (N_10773,N_10309,N_10201);
nor U10774 (N_10774,N_10360,N_10228);
xnor U10775 (N_10775,N_10254,N_10116);
and U10776 (N_10776,N_10493,N_10118);
nand U10777 (N_10777,N_10174,N_10272);
and U10778 (N_10778,N_10266,N_10354);
or U10779 (N_10779,N_10442,N_10357);
and U10780 (N_10780,N_10400,N_10494);
nand U10781 (N_10781,N_10198,N_10343);
and U10782 (N_10782,N_10266,N_10249);
xor U10783 (N_10783,N_10068,N_10190);
and U10784 (N_10784,N_10485,N_10204);
and U10785 (N_10785,N_10494,N_10020);
nor U10786 (N_10786,N_10270,N_10474);
xor U10787 (N_10787,N_10137,N_10079);
nor U10788 (N_10788,N_10093,N_10198);
nand U10789 (N_10789,N_10234,N_10197);
or U10790 (N_10790,N_10253,N_10179);
or U10791 (N_10791,N_10144,N_10101);
or U10792 (N_10792,N_10051,N_10049);
nor U10793 (N_10793,N_10022,N_10449);
nand U10794 (N_10794,N_10142,N_10162);
or U10795 (N_10795,N_10327,N_10054);
or U10796 (N_10796,N_10355,N_10370);
nor U10797 (N_10797,N_10078,N_10123);
and U10798 (N_10798,N_10457,N_10051);
xor U10799 (N_10799,N_10302,N_10036);
or U10800 (N_10800,N_10110,N_10222);
nor U10801 (N_10801,N_10405,N_10099);
xnor U10802 (N_10802,N_10468,N_10217);
nor U10803 (N_10803,N_10464,N_10419);
nand U10804 (N_10804,N_10205,N_10359);
nor U10805 (N_10805,N_10276,N_10494);
and U10806 (N_10806,N_10281,N_10047);
nand U10807 (N_10807,N_10020,N_10352);
or U10808 (N_10808,N_10366,N_10206);
xnor U10809 (N_10809,N_10003,N_10093);
and U10810 (N_10810,N_10046,N_10235);
xor U10811 (N_10811,N_10285,N_10311);
nand U10812 (N_10812,N_10300,N_10467);
xor U10813 (N_10813,N_10483,N_10025);
nand U10814 (N_10814,N_10173,N_10050);
xnor U10815 (N_10815,N_10403,N_10079);
xnor U10816 (N_10816,N_10436,N_10352);
nor U10817 (N_10817,N_10260,N_10105);
nand U10818 (N_10818,N_10468,N_10208);
nand U10819 (N_10819,N_10306,N_10356);
nor U10820 (N_10820,N_10245,N_10043);
xor U10821 (N_10821,N_10466,N_10139);
nor U10822 (N_10822,N_10463,N_10428);
xnor U10823 (N_10823,N_10012,N_10388);
or U10824 (N_10824,N_10141,N_10444);
and U10825 (N_10825,N_10273,N_10469);
nand U10826 (N_10826,N_10412,N_10472);
nor U10827 (N_10827,N_10210,N_10050);
xnor U10828 (N_10828,N_10396,N_10112);
nor U10829 (N_10829,N_10105,N_10371);
xor U10830 (N_10830,N_10059,N_10007);
and U10831 (N_10831,N_10186,N_10239);
and U10832 (N_10832,N_10428,N_10078);
and U10833 (N_10833,N_10150,N_10470);
or U10834 (N_10834,N_10493,N_10260);
nand U10835 (N_10835,N_10189,N_10220);
nand U10836 (N_10836,N_10170,N_10073);
or U10837 (N_10837,N_10233,N_10178);
or U10838 (N_10838,N_10432,N_10240);
or U10839 (N_10839,N_10476,N_10408);
or U10840 (N_10840,N_10146,N_10491);
nand U10841 (N_10841,N_10258,N_10248);
nand U10842 (N_10842,N_10288,N_10400);
xnor U10843 (N_10843,N_10152,N_10346);
and U10844 (N_10844,N_10378,N_10156);
xor U10845 (N_10845,N_10423,N_10435);
xor U10846 (N_10846,N_10050,N_10139);
nor U10847 (N_10847,N_10125,N_10056);
xnor U10848 (N_10848,N_10114,N_10433);
and U10849 (N_10849,N_10039,N_10249);
nand U10850 (N_10850,N_10174,N_10200);
nand U10851 (N_10851,N_10492,N_10127);
nor U10852 (N_10852,N_10263,N_10269);
nand U10853 (N_10853,N_10302,N_10489);
nor U10854 (N_10854,N_10393,N_10289);
and U10855 (N_10855,N_10195,N_10332);
xor U10856 (N_10856,N_10006,N_10366);
nand U10857 (N_10857,N_10305,N_10004);
nor U10858 (N_10858,N_10280,N_10490);
nand U10859 (N_10859,N_10064,N_10049);
nand U10860 (N_10860,N_10341,N_10124);
and U10861 (N_10861,N_10264,N_10287);
nor U10862 (N_10862,N_10317,N_10017);
nor U10863 (N_10863,N_10246,N_10012);
nand U10864 (N_10864,N_10336,N_10383);
xor U10865 (N_10865,N_10034,N_10345);
and U10866 (N_10866,N_10242,N_10099);
and U10867 (N_10867,N_10465,N_10024);
and U10868 (N_10868,N_10022,N_10220);
nand U10869 (N_10869,N_10063,N_10173);
nand U10870 (N_10870,N_10318,N_10281);
nor U10871 (N_10871,N_10069,N_10081);
xor U10872 (N_10872,N_10101,N_10018);
xnor U10873 (N_10873,N_10287,N_10226);
nand U10874 (N_10874,N_10181,N_10344);
or U10875 (N_10875,N_10098,N_10012);
nand U10876 (N_10876,N_10309,N_10286);
xor U10877 (N_10877,N_10067,N_10200);
nor U10878 (N_10878,N_10177,N_10221);
or U10879 (N_10879,N_10487,N_10139);
nand U10880 (N_10880,N_10227,N_10395);
xnor U10881 (N_10881,N_10254,N_10157);
and U10882 (N_10882,N_10077,N_10462);
xor U10883 (N_10883,N_10123,N_10385);
or U10884 (N_10884,N_10366,N_10425);
and U10885 (N_10885,N_10124,N_10404);
and U10886 (N_10886,N_10377,N_10350);
and U10887 (N_10887,N_10373,N_10224);
nor U10888 (N_10888,N_10377,N_10223);
or U10889 (N_10889,N_10282,N_10432);
nand U10890 (N_10890,N_10041,N_10076);
xor U10891 (N_10891,N_10076,N_10110);
xor U10892 (N_10892,N_10195,N_10232);
xnor U10893 (N_10893,N_10241,N_10078);
nor U10894 (N_10894,N_10236,N_10090);
xor U10895 (N_10895,N_10165,N_10159);
and U10896 (N_10896,N_10466,N_10123);
and U10897 (N_10897,N_10145,N_10064);
or U10898 (N_10898,N_10241,N_10133);
nand U10899 (N_10899,N_10016,N_10133);
and U10900 (N_10900,N_10396,N_10073);
nor U10901 (N_10901,N_10043,N_10049);
nor U10902 (N_10902,N_10376,N_10423);
nand U10903 (N_10903,N_10311,N_10438);
nand U10904 (N_10904,N_10397,N_10381);
nand U10905 (N_10905,N_10369,N_10152);
nand U10906 (N_10906,N_10179,N_10126);
nand U10907 (N_10907,N_10222,N_10191);
xnor U10908 (N_10908,N_10468,N_10012);
nand U10909 (N_10909,N_10124,N_10069);
nand U10910 (N_10910,N_10071,N_10095);
xor U10911 (N_10911,N_10214,N_10114);
nand U10912 (N_10912,N_10170,N_10129);
or U10913 (N_10913,N_10012,N_10221);
nor U10914 (N_10914,N_10461,N_10388);
or U10915 (N_10915,N_10052,N_10401);
xnor U10916 (N_10916,N_10373,N_10455);
xor U10917 (N_10917,N_10313,N_10404);
or U10918 (N_10918,N_10392,N_10262);
and U10919 (N_10919,N_10153,N_10447);
xor U10920 (N_10920,N_10491,N_10206);
nor U10921 (N_10921,N_10471,N_10140);
nor U10922 (N_10922,N_10141,N_10407);
xnor U10923 (N_10923,N_10252,N_10236);
xnor U10924 (N_10924,N_10336,N_10433);
and U10925 (N_10925,N_10281,N_10188);
or U10926 (N_10926,N_10498,N_10121);
xnor U10927 (N_10927,N_10351,N_10342);
or U10928 (N_10928,N_10321,N_10031);
nor U10929 (N_10929,N_10086,N_10282);
nor U10930 (N_10930,N_10429,N_10441);
and U10931 (N_10931,N_10498,N_10276);
or U10932 (N_10932,N_10014,N_10133);
xor U10933 (N_10933,N_10409,N_10444);
nor U10934 (N_10934,N_10349,N_10166);
nor U10935 (N_10935,N_10370,N_10077);
xnor U10936 (N_10936,N_10079,N_10436);
or U10937 (N_10937,N_10332,N_10243);
or U10938 (N_10938,N_10304,N_10333);
xor U10939 (N_10939,N_10388,N_10488);
nor U10940 (N_10940,N_10113,N_10299);
xor U10941 (N_10941,N_10129,N_10059);
nand U10942 (N_10942,N_10217,N_10244);
and U10943 (N_10943,N_10257,N_10195);
or U10944 (N_10944,N_10185,N_10354);
nand U10945 (N_10945,N_10423,N_10246);
nand U10946 (N_10946,N_10241,N_10308);
nor U10947 (N_10947,N_10425,N_10298);
or U10948 (N_10948,N_10239,N_10179);
and U10949 (N_10949,N_10195,N_10406);
xnor U10950 (N_10950,N_10281,N_10122);
xnor U10951 (N_10951,N_10166,N_10331);
nand U10952 (N_10952,N_10134,N_10253);
nand U10953 (N_10953,N_10095,N_10026);
xor U10954 (N_10954,N_10009,N_10284);
xnor U10955 (N_10955,N_10064,N_10289);
nor U10956 (N_10956,N_10291,N_10352);
xor U10957 (N_10957,N_10009,N_10010);
and U10958 (N_10958,N_10465,N_10055);
and U10959 (N_10959,N_10118,N_10137);
or U10960 (N_10960,N_10143,N_10365);
or U10961 (N_10961,N_10067,N_10016);
nor U10962 (N_10962,N_10433,N_10203);
and U10963 (N_10963,N_10268,N_10025);
or U10964 (N_10964,N_10152,N_10011);
nor U10965 (N_10965,N_10366,N_10304);
and U10966 (N_10966,N_10189,N_10241);
xnor U10967 (N_10967,N_10058,N_10435);
xnor U10968 (N_10968,N_10139,N_10219);
and U10969 (N_10969,N_10158,N_10327);
nor U10970 (N_10970,N_10215,N_10234);
or U10971 (N_10971,N_10449,N_10121);
or U10972 (N_10972,N_10231,N_10026);
nand U10973 (N_10973,N_10218,N_10153);
and U10974 (N_10974,N_10378,N_10313);
or U10975 (N_10975,N_10121,N_10224);
or U10976 (N_10976,N_10157,N_10387);
and U10977 (N_10977,N_10161,N_10191);
nor U10978 (N_10978,N_10048,N_10150);
nand U10979 (N_10979,N_10352,N_10023);
nor U10980 (N_10980,N_10448,N_10405);
or U10981 (N_10981,N_10405,N_10489);
or U10982 (N_10982,N_10075,N_10359);
nand U10983 (N_10983,N_10238,N_10342);
nand U10984 (N_10984,N_10469,N_10345);
nor U10985 (N_10985,N_10218,N_10236);
nor U10986 (N_10986,N_10164,N_10258);
or U10987 (N_10987,N_10444,N_10178);
nand U10988 (N_10988,N_10214,N_10212);
or U10989 (N_10989,N_10121,N_10351);
nor U10990 (N_10990,N_10251,N_10167);
or U10991 (N_10991,N_10021,N_10078);
or U10992 (N_10992,N_10287,N_10247);
and U10993 (N_10993,N_10015,N_10455);
or U10994 (N_10994,N_10032,N_10454);
xor U10995 (N_10995,N_10064,N_10259);
xnor U10996 (N_10996,N_10127,N_10056);
and U10997 (N_10997,N_10103,N_10178);
nor U10998 (N_10998,N_10301,N_10050);
or U10999 (N_10999,N_10313,N_10141);
nand U11000 (N_11000,N_10666,N_10855);
xor U11001 (N_11001,N_10750,N_10562);
or U11002 (N_11002,N_10647,N_10643);
nor U11003 (N_11003,N_10617,N_10600);
xor U11004 (N_11004,N_10628,N_10866);
or U11005 (N_11005,N_10763,N_10556);
or U11006 (N_11006,N_10873,N_10657);
nand U11007 (N_11007,N_10594,N_10904);
and U11008 (N_11008,N_10805,N_10799);
xor U11009 (N_11009,N_10792,N_10755);
or U11010 (N_11010,N_10886,N_10630);
or U11011 (N_11011,N_10777,N_10868);
nand U11012 (N_11012,N_10642,N_10512);
xnor U11013 (N_11013,N_10874,N_10583);
nand U11014 (N_11014,N_10925,N_10638);
or U11015 (N_11015,N_10681,N_10716);
nand U11016 (N_11016,N_10570,N_10902);
or U11017 (N_11017,N_10964,N_10685);
xor U11018 (N_11018,N_10559,N_10542);
or U11019 (N_11019,N_10606,N_10553);
or U11020 (N_11020,N_10650,N_10587);
and U11021 (N_11021,N_10834,N_10845);
nand U11022 (N_11022,N_10895,N_10725);
nand U11023 (N_11023,N_10742,N_10804);
nor U11024 (N_11024,N_10621,N_10765);
nand U11025 (N_11025,N_10673,N_10974);
and U11026 (N_11026,N_10539,N_10979);
or U11027 (N_11027,N_10893,N_10880);
or U11028 (N_11028,N_10667,N_10596);
xnor U11029 (N_11029,N_10508,N_10905);
nor U11030 (N_11030,N_10669,N_10857);
nand U11031 (N_11031,N_10535,N_10926);
xnor U11032 (N_11032,N_10527,N_10514);
and U11033 (N_11033,N_10578,N_10821);
and U11034 (N_11034,N_10809,N_10887);
xnor U11035 (N_11035,N_10551,N_10814);
or U11036 (N_11036,N_10714,N_10770);
and U11037 (N_11037,N_10826,N_10573);
nand U11038 (N_11038,N_10953,N_10919);
nor U11039 (N_11039,N_10790,N_10747);
nor U11040 (N_11040,N_10783,N_10862);
nor U11041 (N_11041,N_10989,N_10848);
or U11042 (N_11042,N_10636,N_10737);
nand U11043 (N_11043,N_10815,N_10724);
xnor U11044 (N_11044,N_10852,N_10661);
nor U11045 (N_11045,N_10710,N_10867);
or U11046 (N_11046,N_10812,N_10516);
nor U11047 (N_11047,N_10720,N_10611);
and U11048 (N_11048,N_10718,N_10824);
xor U11049 (N_11049,N_10693,N_10787);
nor U11050 (N_11050,N_10973,N_10665);
nor U11051 (N_11051,N_10995,N_10978);
and U11052 (N_11052,N_10908,N_10761);
nand U11053 (N_11053,N_10865,N_10762);
or U11054 (N_11054,N_10913,N_10746);
nor U11055 (N_11055,N_10706,N_10697);
or U11056 (N_11056,N_10590,N_10757);
xor U11057 (N_11057,N_10567,N_10938);
xor U11058 (N_11058,N_10684,N_10603);
nor U11059 (N_11059,N_10536,N_10923);
nor U11060 (N_11060,N_10807,N_10911);
and U11061 (N_11061,N_10533,N_10549);
xnor U11062 (N_11062,N_10952,N_10963);
and U11063 (N_11063,N_10550,N_10956);
nand U11064 (N_11064,N_10994,N_10589);
xor U11065 (N_11065,N_10591,N_10727);
xnor U11066 (N_11066,N_10751,N_10878);
nand U11067 (N_11067,N_10932,N_10959);
nor U11068 (N_11068,N_10827,N_10829);
and U11069 (N_11069,N_10945,N_10561);
or U11070 (N_11070,N_10768,N_10990);
nand U11071 (N_11071,N_10592,N_10711);
and U11072 (N_11072,N_10564,N_10613);
nor U11073 (N_11073,N_10789,N_10988);
or U11074 (N_11074,N_10916,N_10851);
nand U11075 (N_11075,N_10840,N_10883);
or U11076 (N_11076,N_10912,N_10877);
or U11077 (N_11077,N_10506,N_10608);
or U11078 (N_11078,N_10601,N_10985);
and U11079 (N_11079,N_10502,N_10655);
nor U11080 (N_11080,N_10580,N_10889);
nor U11081 (N_11081,N_10781,N_10609);
nor U11082 (N_11082,N_10728,N_10772);
and U11083 (N_11083,N_10907,N_10691);
nor U11084 (N_11084,N_10644,N_10951);
nor U11085 (N_11085,N_10802,N_10610);
nand U11086 (N_11086,N_10800,N_10860);
and U11087 (N_11087,N_10664,N_10870);
xnor U11088 (N_11088,N_10723,N_10803);
nand U11089 (N_11089,N_10631,N_10841);
nand U11090 (N_11090,N_10869,N_10922);
xor U11091 (N_11091,N_10838,N_10897);
nand U11092 (N_11092,N_10884,N_10704);
or U11093 (N_11093,N_10853,N_10517);
or U11094 (N_11094,N_10776,N_10702);
or U11095 (N_11095,N_10983,N_10901);
and U11096 (N_11096,N_10523,N_10795);
or U11097 (N_11097,N_10962,N_10961);
nand U11098 (N_11098,N_10986,N_10722);
or U11099 (N_11099,N_10620,N_10876);
xnor U11100 (N_11100,N_10607,N_10552);
nand U11101 (N_11101,N_10575,N_10936);
xnor U11102 (N_11102,N_10987,N_10577);
and U11103 (N_11103,N_10659,N_10612);
and U11104 (N_11104,N_10641,N_10977);
or U11105 (N_11105,N_10520,N_10504);
xnor U11106 (N_11106,N_10858,N_10957);
nor U11107 (N_11107,N_10859,N_10784);
or U11108 (N_11108,N_10689,N_10721);
or U11109 (N_11109,N_10984,N_10934);
nand U11110 (N_11110,N_10531,N_10888);
nor U11111 (N_11111,N_10672,N_10519);
and U11112 (N_11112,N_10705,N_10965);
xor U11113 (N_11113,N_10909,N_10939);
or U11114 (N_11114,N_10663,N_10712);
or U11115 (N_11115,N_10856,N_10754);
and U11116 (N_11116,N_10822,N_10576);
nand U11117 (N_11117,N_10811,N_10696);
nand U11118 (N_11118,N_10782,N_10971);
nor U11119 (N_11119,N_10688,N_10891);
nor U11120 (N_11120,N_10844,N_10633);
nand U11121 (N_11121,N_10692,N_10579);
nand U11122 (N_11122,N_10568,N_10538);
xnor U11123 (N_11123,N_10726,N_10529);
or U11124 (N_11124,N_10813,N_10654);
or U11125 (N_11125,N_10832,N_10791);
and U11126 (N_11126,N_10753,N_10769);
xnor U11127 (N_11127,N_10645,N_10894);
nand U11128 (N_11128,N_10678,N_10930);
xor U11129 (N_11129,N_10543,N_10937);
nor U11130 (N_11130,N_10920,N_10810);
xnor U11131 (N_11131,N_10980,N_10554);
or U11132 (N_11132,N_10545,N_10586);
nor U11133 (N_11133,N_10565,N_10839);
nor U11134 (N_11134,N_10569,N_10574);
or U11135 (N_11135,N_10794,N_10875);
or U11136 (N_11136,N_10816,N_10540);
nor U11137 (N_11137,N_10732,N_10864);
nand U11138 (N_11138,N_10557,N_10749);
and U11139 (N_11139,N_10509,N_10882);
or U11140 (N_11140,N_10534,N_10639);
xor U11141 (N_11141,N_10744,N_10560);
nand U11142 (N_11142,N_10892,N_10879);
or U11143 (N_11143,N_10597,N_10975);
nand U11144 (N_11144,N_10501,N_10532);
or U11145 (N_11145,N_10566,N_10899);
and U11146 (N_11146,N_10863,N_10652);
nor U11147 (N_11147,N_10677,N_10555);
or U11148 (N_11148,N_10843,N_10760);
nand U11149 (N_11149,N_10670,N_10739);
nor U11150 (N_11150,N_10849,N_10831);
xor U11151 (N_11151,N_10825,N_10730);
nor U11152 (N_11152,N_10954,N_10703);
nor U11153 (N_11153,N_10940,N_10699);
nand U11154 (N_11154,N_10637,N_10518);
nand U11155 (N_11155,N_10996,N_10695);
and U11156 (N_11156,N_10806,N_10854);
or U11157 (N_11157,N_10896,N_10694);
or U11158 (N_11158,N_10819,N_10779);
or U11159 (N_11159,N_10708,N_10949);
or U11160 (N_11160,N_10798,N_10521);
nand U11161 (N_11161,N_10547,N_10595);
nor U11162 (N_11162,N_10752,N_10513);
nand U11163 (N_11163,N_10717,N_10872);
or U11164 (N_11164,N_10615,N_10946);
or U11165 (N_11165,N_10653,N_10731);
and U11166 (N_11166,N_10500,N_10778);
nand U11167 (N_11167,N_10915,N_10709);
or U11168 (N_11168,N_10830,N_10528);
nand U11169 (N_11169,N_10503,N_10871);
nor U11170 (N_11170,N_10788,N_10786);
and U11171 (N_11171,N_10808,N_10736);
or U11172 (N_11172,N_10982,N_10823);
xor U11173 (N_11173,N_10847,N_10616);
and U11174 (N_11174,N_10976,N_10649);
nand U11175 (N_11175,N_10968,N_10698);
nor U11176 (N_11176,N_10548,N_10525);
nor U11177 (N_11177,N_10793,N_10690);
and U11178 (N_11178,N_10676,N_10625);
xnor U11179 (N_11179,N_10679,N_10623);
nor U11180 (N_11180,N_10917,N_10598);
or U11181 (N_11181,N_10960,N_10947);
xor U11182 (N_11182,N_10950,N_10571);
nand U11183 (N_11183,N_10740,N_10683);
and U11184 (N_11184,N_10572,N_10671);
xor U11185 (N_11185,N_10967,N_10687);
nand U11186 (N_11186,N_10646,N_10526);
xnor U11187 (N_11187,N_10584,N_10675);
and U11188 (N_11188,N_10581,N_10593);
xor U11189 (N_11189,N_10921,N_10756);
and U11190 (N_11190,N_10944,N_10748);
and U11191 (N_11191,N_10614,N_10660);
or U11192 (N_11192,N_10828,N_10972);
and U11193 (N_11193,N_10632,N_10624);
nand U11194 (N_11194,N_10797,N_10619);
xor U11195 (N_11195,N_10966,N_10943);
xnor U11196 (N_11196,N_10942,N_10668);
and U11197 (N_11197,N_10758,N_10510);
nand U11198 (N_11198,N_10817,N_10935);
xnor U11199 (N_11199,N_10729,N_10998);
and U11200 (N_11200,N_10928,N_10993);
nor U11201 (N_11201,N_10970,N_10801);
nor U11202 (N_11202,N_10741,N_10767);
and U11203 (N_11203,N_10686,N_10846);
or U11204 (N_11204,N_10515,N_10733);
nand U11205 (N_11205,N_10780,N_10544);
nand U11206 (N_11206,N_10651,N_10850);
or U11207 (N_11207,N_10766,N_10898);
nand U11208 (N_11208,N_10713,N_10861);
xor U11209 (N_11209,N_10719,N_10818);
xnor U11210 (N_11210,N_10629,N_10820);
nand U11211 (N_11211,N_10524,N_10836);
and U11212 (N_11212,N_10507,N_10738);
xnor U11213 (N_11213,N_10715,N_10537);
nor U11214 (N_11214,N_10842,N_10764);
nand U11215 (N_11215,N_10785,N_10910);
xor U11216 (N_11216,N_10835,N_10734);
nor U11217 (N_11217,N_10918,N_10622);
xor U11218 (N_11218,N_10948,N_10837);
nand U11219 (N_11219,N_10599,N_10627);
nor U11220 (N_11220,N_10604,N_10796);
nand U11221 (N_11221,N_10981,N_10969);
nor U11222 (N_11222,N_10759,N_10635);
or U11223 (N_11223,N_10626,N_10997);
xnor U11224 (N_11224,N_10530,N_10774);
nor U11225 (N_11225,N_10773,N_10658);
or U11226 (N_11226,N_10680,N_10900);
nand U11227 (N_11227,N_10582,N_10618);
and U11228 (N_11228,N_10588,N_10707);
nor U11229 (N_11229,N_10924,N_10634);
xnor U11230 (N_11230,N_10941,N_10585);
nand U11231 (N_11231,N_10640,N_10992);
or U11232 (N_11232,N_10511,N_10914);
nand U11233 (N_11233,N_10546,N_10743);
and U11234 (N_11234,N_10833,N_10735);
or U11235 (N_11235,N_10602,N_10881);
xor U11236 (N_11236,N_10674,N_10927);
nand U11237 (N_11237,N_10906,N_10991);
and U11238 (N_11238,N_10522,N_10958);
xor U11239 (N_11239,N_10563,N_10929);
xor U11240 (N_11240,N_10931,N_10999);
nor U11241 (N_11241,N_10955,N_10885);
nand U11242 (N_11242,N_10701,N_10558);
and U11243 (N_11243,N_10662,N_10682);
nand U11244 (N_11244,N_10605,N_10505);
and U11245 (N_11245,N_10745,N_10775);
or U11246 (N_11246,N_10890,N_10771);
xor U11247 (N_11247,N_10933,N_10903);
nand U11248 (N_11248,N_10700,N_10656);
xnor U11249 (N_11249,N_10541,N_10648);
and U11250 (N_11250,N_10956,N_10873);
or U11251 (N_11251,N_10857,N_10614);
or U11252 (N_11252,N_10644,N_10679);
nand U11253 (N_11253,N_10827,N_10976);
and U11254 (N_11254,N_10529,N_10783);
or U11255 (N_11255,N_10843,N_10533);
and U11256 (N_11256,N_10758,N_10674);
and U11257 (N_11257,N_10618,N_10713);
or U11258 (N_11258,N_10695,N_10751);
nand U11259 (N_11259,N_10979,N_10616);
nand U11260 (N_11260,N_10720,N_10881);
xor U11261 (N_11261,N_10914,N_10722);
xnor U11262 (N_11262,N_10839,N_10649);
nand U11263 (N_11263,N_10807,N_10568);
nor U11264 (N_11264,N_10806,N_10821);
nor U11265 (N_11265,N_10690,N_10758);
and U11266 (N_11266,N_10556,N_10540);
xor U11267 (N_11267,N_10503,N_10855);
nor U11268 (N_11268,N_10612,N_10550);
xor U11269 (N_11269,N_10572,N_10813);
and U11270 (N_11270,N_10809,N_10504);
nand U11271 (N_11271,N_10940,N_10520);
or U11272 (N_11272,N_10723,N_10560);
xnor U11273 (N_11273,N_10871,N_10658);
or U11274 (N_11274,N_10923,N_10721);
nand U11275 (N_11275,N_10945,N_10685);
xor U11276 (N_11276,N_10740,N_10511);
nor U11277 (N_11277,N_10926,N_10741);
nand U11278 (N_11278,N_10999,N_10939);
xor U11279 (N_11279,N_10943,N_10827);
or U11280 (N_11280,N_10733,N_10857);
nand U11281 (N_11281,N_10528,N_10764);
and U11282 (N_11282,N_10857,N_10688);
or U11283 (N_11283,N_10605,N_10563);
or U11284 (N_11284,N_10690,N_10778);
nand U11285 (N_11285,N_10641,N_10590);
nand U11286 (N_11286,N_10845,N_10929);
nand U11287 (N_11287,N_10547,N_10571);
xor U11288 (N_11288,N_10891,N_10985);
or U11289 (N_11289,N_10953,N_10923);
and U11290 (N_11290,N_10925,N_10975);
xor U11291 (N_11291,N_10933,N_10668);
nand U11292 (N_11292,N_10699,N_10886);
nand U11293 (N_11293,N_10705,N_10945);
or U11294 (N_11294,N_10818,N_10865);
or U11295 (N_11295,N_10513,N_10821);
xor U11296 (N_11296,N_10755,N_10867);
or U11297 (N_11297,N_10529,N_10894);
or U11298 (N_11298,N_10649,N_10621);
nand U11299 (N_11299,N_10812,N_10980);
nor U11300 (N_11300,N_10735,N_10803);
nor U11301 (N_11301,N_10752,N_10683);
nor U11302 (N_11302,N_10631,N_10937);
xor U11303 (N_11303,N_10672,N_10942);
or U11304 (N_11304,N_10704,N_10854);
nand U11305 (N_11305,N_10635,N_10613);
xnor U11306 (N_11306,N_10770,N_10986);
or U11307 (N_11307,N_10578,N_10513);
xor U11308 (N_11308,N_10730,N_10857);
nand U11309 (N_11309,N_10816,N_10584);
nand U11310 (N_11310,N_10814,N_10505);
nor U11311 (N_11311,N_10755,N_10947);
nand U11312 (N_11312,N_10692,N_10824);
nand U11313 (N_11313,N_10666,N_10583);
xor U11314 (N_11314,N_10544,N_10918);
or U11315 (N_11315,N_10578,N_10522);
nor U11316 (N_11316,N_10932,N_10560);
nand U11317 (N_11317,N_10949,N_10726);
and U11318 (N_11318,N_10568,N_10628);
nor U11319 (N_11319,N_10997,N_10589);
nand U11320 (N_11320,N_10913,N_10769);
or U11321 (N_11321,N_10945,N_10847);
nand U11322 (N_11322,N_10529,N_10930);
nor U11323 (N_11323,N_10627,N_10527);
xnor U11324 (N_11324,N_10525,N_10845);
and U11325 (N_11325,N_10592,N_10849);
nor U11326 (N_11326,N_10805,N_10594);
nor U11327 (N_11327,N_10770,N_10797);
or U11328 (N_11328,N_10624,N_10541);
xnor U11329 (N_11329,N_10664,N_10726);
nand U11330 (N_11330,N_10963,N_10555);
nand U11331 (N_11331,N_10651,N_10581);
xor U11332 (N_11332,N_10850,N_10749);
or U11333 (N_11333,N_10992,N_10553);
nand U11334 (N_11334,N_10720,N_10764);
and U11335 (N_11335,N_10548,N_10731);
or U11336 (N_11336,N_10918,N_10984);
or U11337 (N_11337,N_10681,N_10826);
xnor U11338 (N_11338,N_10635,N_10958);
or U11339 (N_11339,N_10582,N_10924);
xnor U11340 (N_11340,N_10596,N_10745);
nand U11341 (N_11341,N_10994,N_10873);
or U11342 (N_11342,N_10590,N_10679);
or U11343 (N_11343,N_10672,N_10660);
nor U11344 (N_11344,N_10586,N_10579);
and U11345 (N_11345,N_10949,N_10857);
xnor U11346 (N_11346,N_10969,N_10702);
and U11347 (N_11347,N_10909,N_10812);
or U11348 (N_11348,N_10539,N_10544);
xnor U11349 (N_11349,N_10754,N_10537);
xnor U11350 (N_11350,N_10977,N_10936);
xnor U11351 (N_11351,N_10577,N_10930);
nor U11352 (N_11352,N_10944,N_10568);
nand U11353 (N_11353,N_10958,N_10739);
nand U11354 (N_11354,N_10593,N_10971);
nand U11355 (N_11355,N_10901,N_10663);
nor U11356 (N_11356,N_10595,N_10575);
xor U11357 (N_11357,N_10862,N_10945);
nand U11358 (N_11358,N_10716,N_10828);
or U11359 (N_11359,N_10514,N_10558);
nand U11360 (N_11360,N_10592,N_10643);
and U11361 (N_11361,N_10916,N_10573);
or U11362 (N_11362,N_10612,N_10843);
and U11363 (N_11363,N_10764,N_10824);
and U11364 (N_11364,N_10752,N_10967);
nor U11365 (N_11365,N_10809,N_10890);
and U11366 (N_11366,N_10695,N_10807);
and U11367 (N_11367,N_10937,N_10679);
nor U11368 (N_11368,N_10643,N_10554);
or U11369 (N_11369,N_10703,N_10579);
or U11370 (N_11370,N_10769,N_10520);
and U11371 (N_11371,N_10546,N_10535);
nor U11372 (N_11372,N_10969,N_10668);
and U11373 (N_11373,N_10525,N_10729);
nand U11374 (N_11374,N_10859,N_10830);
or U11375 (N_11375,N_10787,N_10745);
xor U11376 (N_11376,N_10978,N_10738);
nor U11377 (N_11377,N_10593,N_10816);
or U11378 (N_11378,N_10861,N_10668);
nor U11379 (N_11379,N_10578,N_10637);
or U11380 (N_11380,N_10622,N_10553);
or U11381 (N_11381,N_10678,N_10896);
nor U11382 (N_11382,N_10530,N_10593);
or U11383 (N_11383,N_10921,N_10575);
xor U11384 (N_11384,N_10575,N_10604);
or U11385 (N_11385,N_10661,N_10560);
and U11386 (N_11386,N_10731,N_10765);
or U11387 (N_11387,N_10562,N_10599);
nand U11388 (N_11388,N_10971,N_10663);
or U11389 (N_11389,N_10903,N_10738);
and U11390 (N_11390,N_10864,N_10608);
or U11391 (N_11391,N_10939,N_10947);
nand U11392 (N_11392,N_10826,N_10736);
and U11393 (N_11393,N_10721,N_10943);
nand U11394 (N_11394,N_10965,N_10686);
or U11395 (N_11395,N_10673,N_10922);
nor U11396 (N_11396,N_10678,N_10873);
or U11397 (N_11397,N_10986,N_10783);
nand U11398 (N_11398,N_10597,N_10591);
or U11399 (N_11399,N_10864,N_10535);
xnor U11400 (N_11400,N_10832,N_10683);
or U11401 (N_11401,N_10765,N_10981);
or U11402 (N_11402,N_10928,N_10593);
xor U11403 (N_11403,N_10927,N_10764);
nand U11404 (N_11404,N_10592,N_10520);
nand U11405 (N_11405,N_10775,N_10909);
nor U11406 (N_11406,N_10760,N_10846);
and U11407 (N_11407,N_10920,N_10645);
nor U11408 (N_11408,N_10610,N_10809);
nor U11409 (N_11409,N_10699,N_10984);
and U11410 (N_11410,N_10500,N_10825);
and U11411 (N_11411,N_10903,N_10536);
nand U11412 (N_11412,N_10688,N_10975);
nand U11413 (N_11413,N_10795,N_10819);
or U11414 (N_11414,N_10812,N_10741);
nor U11415 (N_11415,N_10731,N_10785);
or U11416 (N_11416,N_10582,N_10551);
nor U11417 (N_11417,N_10708,N_10587);
or U11418 (N_11418,N_10970,N_10507);
nor U11419 (N_11419,N_10868,N_10508);
and U11420 (N_11420,N_10739,N_10982);
and U11421 (N_11421,N_10892,N_10518);
nand U11422 (N_11422,N_10540,N_10861);
and U11423 (N_11423,N_10573,N_10510);
nor U11424 (N_11424,N_10929,N_10783);
xor U11425 (N_11425,N_10777,N_10715);
nand U11426 (N_11426,N_10997,N_10999);
and U11427 (N_11427,N_10533,N_10644);
nand U11428 (N_11428,N_10839,N_10528);
nor U11429 (N_11429,N_10781,N_10545);
or U11430 (N_11430,N_10548,N_10554);
or U11431 (N_11431,N_10869,N_10719);
and U11432 (N_11432,N_10546,N_10604);
nand U11433 (N_11433,N_10776,N_10913);
nand U11434 (N_11434,N_10770,N_10864);
nand U11435 (N_11435,N_10556,N_10517);
nor U11436 (N_11436,N_10933,N_10959);
or U11437 (N_11437,N_10562,N_10534);
or U11438 (N_11438,N_10875,N_10500);
or U11439 (N_11439,N_10851,N_10996);
or U11440 (N_11440,N_10552,N_10573);
xor U11441 (N_11441,N_10899,N_10967);
or U11442 (N_11442,N_10654,N_10566);
and U11443 (N_11443,N_10535,N_10788);
and U11444 (N_11444,N_10727,N_10714);
nor U11445 (N_11445,N_10660,N_10849);
and U11446 (N_11446,N_10579,N_10764);
nand U11447 (N_11447,N_10860,N_10625);
or U11448 (N_11448,N_10847,N_10611);
xor U11449 (N_11449,N_10709,N_10590);
xnor U11450 (N_11450,N_10703,N_10894);
and U11451 (N_11451,N_10978,N_10538);
nand U11452 (N_11452,N_10517,N_10915);
and U11453 (N_11453,N_10503,N_10606);
or U11454 (N_11454,N_10548,N_10843);
or U11455 (N_11455,N_10606,N_10943);
nor U11456 (N_11456,N_10605,N_10815);
or U11457 (N_11457,N_10633,N_10511);
nor U11458 (N_11458,N_10753,N_10967);
nor U11459 (N_11459,N_10503,N_10678);
xor U11460 (N_11460,N_10913,N_10582);
xor U11461 (N_11461,N_10714,N_10588);
and U11462 (N_11462,N_10832,N_10961);
or U11463 (N_11463,N_10665,N_10893);
xnor U11464 (N_11464,N_10738,N_10958);
nor U11465 (N_11465,N_10578,N_10928);
nor U11466 (N_11466,N_10996,N_10977);
and U11467 (N_11467,N_10968,N_10623);
xnor U11468 (N_11468,N_10895,N_10938);
nor U11469 (N_11469,N_10603,N_10670);
nor U11470 (N_11470,N_10672,N_10525);
xor U11471 (N_11471,N_10660,N_10896);
nand U11472 (N_11472,N_10970,N_10832);
nand U11473 (N_11473,N_10660,N_10798);
and U11474 (N_11474,N_10839,N_10948);
or U11475 (N_11475,N_10988,N_10599);
or U11476 (N_11476,N_10614,N_10942);
nand U11477 (N_11477,N_10755,N_10986);
or U11478 (N_11478,N_10789,N_10517);
nor U11479 (N_11479,N_10894,N_10813);
nand U11480 (N_11480,N_10502,N_10695);
and U11481 (N_11481,N_10782,N_10997);
and U11482 (N_11482,N_10979,N_10706);
nor U11483 (N_11483,N_10595,N_10689);
and U11484 (N_11484,N_10947,N_10846);
and U11485 (N_11485,N_10860,N_10862);
and U11486 (N_11486,N_10869,N_10516);
and U11487 (N_11487,N_10570,N_10764);
or U11488 (N_11488,N_10609,N_10617);
nor U11489 (N_11489,N_10553,N_10578);
or U11490 (N_11490,N_10615,N_10514);
and U11491 (N_11491,N_10840,N_10748);
nor U11492 (N_11492,N_10987,N_10529);
and U11493 (N_11493,N_10685,N_10543);
and U11494 (N_11494,N_10788,N_10991);
and U11495 (N_11495,N_10998,N_10894);
or U11496 (N_11496,N_10763,N_10854);
and U11497 (N_11497,N_10885,N_10860);
nand U11498 (N_11498,N_10648,N_10706);
nor U11499 (N_11499,N_10740,N_10753);
nand U11500 (N_11500,N_11038,N_11406);
or U11501 (N_11501,N_11092,N_11272);
xor U11502 (N_11502,N_11158,N_11482);
nor U11503 (N_11503,N_11095,N_11198);
xor U11504 (N_11504,N_11480,N_11395);
or U11505 (N_11505,N_11326,N_11112);
nand U11506 (N_11506,N_11056,N_11386);
nand U11507 (N_11507,N_11379,N_11331);
and U11508 (N_11508,N_11321,N_11120);
nand U11509 (N_11509,N_11139,N_11297);
nand U11510 (N_11510,N_11143,N_11413);
xor U11511 (N_11511,N_11082,N_11409);
nand U11512 (N_11512,N_11383,N_11226);
and U11513 (N_11513,N_11387,N_11313);
and U11514 (N_11514,N_11020,N_11316);
nor U11515 (N_11515,N_11343,N_11123);
xnor U11516 (N_11516,N_11437,N_11129);
xnor U11517 (N_11517,N_11087,N_11006);
and U11518 (N_11518,N_11325,N_11348);
or U11519 (N_11519,N_11291,N_11097);
and U11520 (N_11520,N_11197,N_11116);
nor U11521 (N_11521,N_11019,N_11144);
xnor U11522 (N_11522,N_11213,N_11370);
nor U11523 (N_11523,N_11298,N_11474);
nor U11524 (N_11524,N_11396,N_11182);
and U11525 (N_11525,N_11430,N_11152);
xnor U11526 (N_11526,N_11187,N_11093);
nor U11527 (N_11527,N_11372,N_11074);
nand U11528 (N_11528,N_11353,N_11273);
and U11529 (N_11529,N_11276,N_11477);
nor U11530 (N_11530,N_11155,N_11090);
xnor U11531 (N_11531,N_11261,N_11128);
and U11532 (N_11532,N_11333,N_11339);
and U11533 (N_11533,N_11211,N_11171);
xor U11534 (N_11534,N_11418,N_11318);
xor U11535 (N_11535,N_11014,N_11328);
or U11536 (N_11536,N_11342,N_11345);
and U11537 (N_11537,N_11256,N_11141);
and U11538 (N_11538,N_11119,N_11300);
nor U11539 (N_11539,N_11266,N_11435);
or U11540 (N_11540,N_11186,N_11479);
nand U11541 (N_11541,N_11084,N_11384);
xnor U11542 (N_11542,N_11428,N_11420);
or U11543 (N_11543,N_11166,N_11100);
nand U11544 (N_11544,N_11490,N_11105);
nor U11545 (N_11545,N_11189,N_11471);
nor U11546 (N_11546,N_11337,N_11073);
xor U11547 (N_11547,N_11147,N_11125);
or U11548 (N_11548,N_11174,N_11391);
nand U11549 (N_11549,N_11350,N_11466);
nand U11550 (N_11550,N_11184,N_11003);
nand U11551 (N_11551,N_11239,N_11064);
xnor U11552 (N_11552,N_11111,N_11270);
nand U11553 (N_11553,N_11309,N_11140);
xor U11554 (N_11554,N_11269,N_11225);
xnor U11555 (N_11555,N_11277,N_11381);
nor U11556 (N_11556,N_11465,N_11089);
and U11557 (N_11557,N_11389,N_11069);
xnor U11558 (N_11558,N_11148,N_11445);
nor U11559 (N_11559,N_11335,N_11218);
nand U11560 (N_11560,N_11029,N_11427);
nor U11561 (N_11561,N_11290,N_11238);
nand U11562 (N_11562,N_11244,N_11248);
or U11563 (N_11563,N_11062,N_11072);
or U11564 (N_11564,N_11055,N_11150);
nor U11565 (N_11565,N_11071,N_11440);
and U11566 (N_11566,N_11026,N_11423);
and U11567 (N_11567,N_11118,N_11444);
nor U11568 (N_11568,N_11392,N_11401);
and U11569 (N_11569,N_11001,N_11004);
or U11570 (N_11570,N_11371,N_11067);
xor U11571 (N_11571,N_11173,N_11403);
nand U11572 (N_11572,N_11065,N_11322);
nor U11573 (N_11573,N_11405,N_11468);
and U11574 (N_11574,N_11484,N_11136);
and U11575 (N_11575,N_11412,N_11083);
and U11576 (N_11576,N_11134,N_11149);
nor U11577 (N_11577,N_11058,N_11271);
or U11578 (N_11578,N_11044,N_11416);
nand U11579 (N_11579,N_11126,N_11232);
or U11580 (N_11580,N_11181,N_11281);
and U11581 (N_11581,N_11469,N_11033);
nand U11582 (N_11582,N_11156,N_11208);
nor U11583 (N_11583,N_11414,N_11368);
xor U11584 (N_11584,N_11145,N_11461);
nand U11585 (N_11585,N_11485,N_11402);
xnor U11586 (N_11586,N_11340,N_11180);
and U11587 (N_11587,N_11421,N_11076);
nor U11588 (N_11588,N_11346,N_11049);
nor U11589 (N_11589,N_11305,N_11080);
and U11590 (N_11590,N_11324,N_11400);
and U11591 (N_11591,N_11191,N_11061);
and U11592 (N_11592,N_11036,N_11436);
xor U11593 (N_11593,N_11456,N_11453);
or U11594 (N_11594,N_11351,N_11251);
or U11595 (N_11595,N_11454,N_11274);
or U11596 (N_11596,N_11024,N_11317);
and U11597 (N_11597,N_11494,N_11268);
nand U11598 (N_11598,N_11382,N_11216);
nor U11599 (N_11599,N_11363,N_11415);
and U11600 (N_11600,N_11254,N_11397);
xor U11601 (N_11601,N_11323,N_11338);
or U11602 (N_11602,N_11091,N_11078);
and U11603 (N_11603,N_11175,N_11362);
nor U11604 (N_11604,N_11205,N_11288);
nand U11605 (N_11605,N_11230,N_11408);
nand U11606 (N_11606,N_11422,N_11374);
nor U11607 (N_11607,N_11443,N_11311);
nor U11608 (N_11608,N_11267,N_11446);
xnor U11609 (N_11609,N_11114,N_11472);
nor U11610 (N_11610,N_11098,N_11235);
or U11611 (N_11611,N_11434,N_11394);
and U11612 (N_11612,N_11354,N_11204);
xnor U11613 (N_11613,N_11194,N_11496);
or U11614 (N_11614,N_11369,N_11018);
and U11615 (N_11615,N_11282,N_11236);
nor U11616 (N_11616,N_11048,N_11177);
or U11617 (N_11617,N_11227,N_11497);
nor U11618 (N_11618,N_11219,N_11441);
nand U11619 (N_11619,N_11481,N_11028);
or U11620 (N_11620,N_11279,N_11320);
xor U11621 (N_11621,N_11260,N_11410);
nand U11622 (N_11622,N_11011,N_11070);
or U11623 (N_11623,N_11154,N_11110);
and U11624 (N_11624,N_11167,N_11259);
nor U11625 (N_11625,N_11299,N_11138);
and U11626 (N_11626,N_11385,N_11467);
or U11627 (N_11627,N_11046,N_11388);
nand U11628 (N_11628,N_11063,N_11492);
nor U11629 (N_11629,N_11068,N_11130);
and U11630 (N_11630,N_11366,N_11314);
nor U11631 (N_11631,N_11188,N_11442);
or U11632 (N_11632,N_11057,N_11278);
or U11633 (N_11633,N_11329,N_11476);
nor U11634 (N_11634,N_11168,N_11233);
or U11635 (N_11635,N_11117,N_11032);
or U11636 (N_11636,N_11310,N_11215);
and U11637 (N_11637,N_11304,N_11475);
xnor U11638 (N_11638,N_11301,N_11464);
nor U11639 (N_11639,N_11255,N_11122);
nor U11640 (N_11640,N_11263,N_11035);
xnor U11641 (N_11641,N_11356,N_11429);
or U11642 (N_11642,N_11463,N_11203);
and U11643 (N_11643,N_11361,N_11364);
or U11644 (N_11644,N_11241,N_11017);
nand U11645 (N_11645,N_11285,N_11220);
nand U11646 (N_11646,N_11040,N_11165);
nor U11647 (N_11647,N_11106,N_11142);
nor U11648 (N_11648,N_11393,N_11102);
nand U11649 (N_11649,N_11275,N_11498);
xnor U11650 (N_11650,N_11365,N_11210);
or U11651 (N_11651,N_11489,N_11153);
and U11652 (N_11652,N_11450,N_11081);
nor U11653 (N_11653,N_11021,N_11295);
nand U11654 (N_11654,N_11043,N_11200);
nand U11655 (N_11655,N_11280,N_11355);
nor U11656 (N_11656,N_11376,N_11257);
nor U11657 (N_11657,N_11127,N_11367);
xnor U11658 (N_11658,N_11432,N_11283);
and U11659 (N_11659,N_11002,N_11045);
and U11660 (N_11660,N_11289,N_11201);
or U11661 (N_11661,N_11495,N_11245);
and U11662 (N_11662,N_11390,N_11088);
nand U11663 (N_11663,N_11209,N_11193);
xnor U11664 (N_11664,N_11047,N_11109);
nand U11665 (N_11665,N_11341,N_11352);
and U11666 (N_11666,N_11212,N_11359);
xor U11667 (N_11667,N_11195,N_11192);
and U11668 (N_11668,N_11103,N_11160);
nor U11669 (N_11669,N_11448,N_11439);
or U11670 (N_11670,N_11380,N_11132);
nor U11671 (N_11671,N_11493,N_11096);
nor U11672 (N_11672,N_11399,N_11294);
nand U11673 (N_11673,N_11027,N_11411);
nand U11674 (N_11674,N_11258,N_11094);
and U11675 (N_11675,N_11470,N_11344);
xor U11676 (N_11676,N_11050,N_11039);
nor U11677 (N_11677,N_11242,N_11133);
and U11678 (N_11678,N_11086,N_11286);
xor U11679 (N_11679,N_11037,N_11499);
nor U11680 (N_11680,N_11234,N_11000);
nor U11681 (N_11681,N_11438,N_11185);
nand U11682 (N_11682,N_11099,N_11293);
nand U11683 (N_11683,N_11334,N_11085);
and U11684 (N_11684,N_11307,N_11373);
nor U11685 (N_11685,N_11431,N_11190);
nand U11686 (N_11686,N_11163,N_11012);
nand U11687 (N_11687,N_11240,N_11462);
or U11688 (N_11688,N_11228,N_11169);
xor U11689 (N_11689,N_11417,N_11164);
nand U11690 (N_11690,N_11053,N_11460);
or U11691 (N_11691,N_11115,N_11178);
and U11692 (N_11692,N_11358,N_11034);
nand U11693 (N_11693,N_11315,N_11287);
nor U11694 (N_11694,N_11237,N_11478);
or U11695 (N_11695,N_11170,N_11407);
xnor U11696 (N_11696,N_11250,N_11023);
and U11697 (N_11697,N_11146,N_11041);
nor U11698 (N_11698,N_11052,N_11229);
nand U11699 (N_11699,N_11451,N_11360);
nor U11700 (N_11700,N_11302,N_11183);
nand U11701 (N_11701,N_11005,N_11031);
nor U11702 (N_11702,N_11247,N_11378);
nor U11703 (N_11703,N_11457,N_11179);
and U11704 (N_11704,N_11455,N_11433);
and U11705 (N_11705,N_11025,N_11332);
and U11706 (N_11706,N_11319,N_11308);
nor U11707 (N_11707,N_11124,N_11243);
nand U11708 (N_11708,N_11013,N_11113);
xnor U11709 (N_11709,N_11296,N_11207);
nor U11710 (N_11710,N_11452,N_11199);
or U11711 (N_11711,N_11284,N_11010);
and U11712 (N_11712,N_11231,N_11176);
or U11713 (N_11713,N_11487,N_11224);
and U11714 (N_11714,N_11419,N_11357);
xnor U11715 (N_11715,N_11459,N_11425);
or U11716 (N_11716,N_11246,N_11030);
xnor U11717 (N_11717,N_11491,N_11424);
or U11718 (N_11718,N_11022,N_11473);
nor U11719 (N_11719,N_11108,N_11079);
xnor U11720 (N_11720,N_11066,N_11131);
and U11721 (N_11721,N_11016,N_11264);
and U11722 (N_11722,N_11253,N_11214);
and U11723 (N_11723,N_11202,N_11206);
nand U11724 (N_11724,N_11306,N_11249);
or U11725 (N_11725,N_11059,N_11488);
nand U11726 (N_11726,N_11172,N_11375);
xnor U11727 (N_11727,N_11262,N_11486);
xnor U11728 (N_11728,N_11060,N_11077);
or U11729 (N_11729,N_11159,N_11349);
nand U11730 (N_11730,N_11121,N_11336);
nand U11731 (N_11731,N_11009,N_11221);
or U11732 (N_11732,N_11449,N_11252);
nand U11733 (N_11733,N_11398,N_11051);
xor U11734 (N_11734,N_11042,N_11162);
nand U11735 (N_11735,N_11426,N_11054);
or U11736 (N_11736,N_11161,N_11377);
xnor U11737 (N_11737,N_11104,N_11157);
and U11738 (N_11738,N_11327,N_11196);
and U11739 (N_11739,N_11137,N_11404);
xnor U11740 (N_11740,N_11447,N_11151);
and U11741 (N_11741,N_11303,N_11222);
and U11742 (N_11742,N_11101,N_11075);
or U11743 (N_11743,N_11008,N_11135);
nor U11744 (N_11744,N_11312,N_11483);
xor U11745 (N_11745,N_11458,N_11347);
or U11746 (N_11746,N_11007,N_11330);
or U11747 (N_11747,N_11015,N_11265);
nand U11748 (N_11748,N_11292,N_11223);
xor U11749 (N_11749,N_11107,N_11217);
xnor U11750 (N_11750,N_11233,N_11100);
nor U11751 (N_11751,N_11450,N_11106);
nand U11752 (N_11752,N_11433,N_11182);
and U11753 (N_11753,N_11084,N_11090);
xor U11754 (N_11754,N_11255,N_11048);
xnor U11755 (N_11755,N_11053,N_11173);
xor U11756 (N_11756,N_11077,N_11404);
or U11757 (N_11757,N_11484,N_11045);
nor U11758 (N_11758,N_11295,N_11011);
nand U11759 (N_11759,N_11127,N_11199);
or U11760 (N_11760,N_11071,N_11423);
nor U11761 (N_11761,N_11114,N_11054);
nand U11762 (N_11762,N_11433,N_11144);
xnor U11763 (N_11763,N_11309,N_11081);
or U11764 (N_11764,N_11440,N_11121);
xor U11765 (N_11765,N_11205,N_11385);
xor U11766 (N_11766,N_11339,N_11117);
nand U11767 (N_11767,N_11136,N_11245);
xor U11768 (N_11768,N_11215,N_11458);
and U11769 (N_11769,N_11215,N_11213);
and U11770 (N_11770,N_11383,N_11172);
nor U11771 (N_11771,N_11417,N_11486);
xnor U11772 (N_11772,N_11288,N_11308);
nor U11773 (N_11773,N_11094,N_11185);
xor U11774 (N_11774,N_11037,N_11197);
and U11775 (N_11775,N_11098,N_11420);
xnor U11776 (N_11776,N_11309,N_11094);
or U11777 (N_11777,N_11478,N_11147);
nor U11778 (N_11778,N_11170,N_11252);
nor U11779 (N_11779,N_11235,N_11259);
and U11780 (N_11780,N_11019,N_11438);
nor U11781 (N_11781,N_11196,N_11356);
xnor U11782 (N_11782,N_11488,N_11273);
nor U11783 (N_11783,N_11486,N_11164);
nand U11784 (N_11784,N_11329,N_11425);
or U11785 (N_11785,N_11008,N_11065);
nor U11786 (N_11786,N_11233,N_11488);
and U11787 (N_11787,N_11173,N_11494);
nor U11788 (N_11788,N_11376,N_11451);
and U11789 (N_11789,N_11319,N_11082);
or U11790 (N_11790,N_11113,N_11155);
xor U11791 (N_11791,N_11321,N_11044);
and U11792 (N_11792,N_11010,N_11292);
nand U11793 (N_11793,N_11079,N_11433);
and U11794 (N_11794,N_11247,N_11189);
or U11795 (N_11795,N_11084,N_11468);
or U11796 (N_11796,N_11362,N_11298);
nand U11797 (N_11797,N_11163,N_11492);
and U11798 (N_11798,N_11026,N_11055);
or U11799 (N_11799,N_11489,N_11058);
nor U11800 (N_11800,N_11078,N_11291);
xor U11801 (N_11801,N_11485,N_11224);
nand U11802 (N_11802,N_11422,N_11437);
xor U11803 (N_11803,N_11450,N_11212);
or U11804 (N_11804,N_11413,N_11376);
and U11805 (N_11805,N_11222,N_11472);
nand U11806 (N_11806,N_11038,N_11413);
nor U11807 (N_11807,N_11286,N_11400);
and U11808 (N_11808,N_11319,N_11006);
xnor U11809 (N_11809,N_11459,N_11427);
or U11810 (N_11810,N_11474,N_11224);
nor U11811 (N_11811,N_11310,N_11320);
nor U11812 (N_11812,N_11497,N_11115);
nand U11813 (N_11813,N_11403,N_11294);
nor U11814 (N_11814,N_11017,N_11325);
xor U11815 (N_11815,N_11495,N_11139);
nor U11816 (N_11816,N_11335,N_11153);
nor U11817 (N_11817,N_11405,N_11103);
or U11818 (N_11818,N_11159,N_11370);
xor U11819 (N_11819,N_11370,N_11227);
xor U11820 (N_11820,N_11171,N_11172);
and U11821 (N_11821,N_11005,N_11184);
and U11822 (N_11822,N_11292,N_11457);
nand U11823 (N_11823,N_11158,N_11495);
xor U11824 (N_11824,N_11251,N_11412);
or U11825 (N_11825,N_11201,N_11428);
nand U11826 (N_11826,N_11334,N_11317);
and U11827 (N_11827,N_11484,N_11320);
xnor U11828 (N_11828,N_11103,N_11452);
or U11829 (N_11829,N_11151,N_11485);
nand U11830 (N_11830,N_11426,N_11021);
or U11831 (N_11831,N_11368,N_11314);
and U11832 (N_11832,N_11394,N_11134);
and U11833 (N_11833,N_11124,N_11366);
nor U11834 (N_11834,N_11115,N_11449);
nand U11835 (N_11835,N_11014,N_11111);
nor U11836 (N_11836,N_11139,N_11364);
and U11837 (N_11837,N_11033,N_11282);
and U11838 (N_11838,N_11157,N_11328);
xnor U11839 (N_11839,N_11145,N_11440);
nand U11840 (N_11840,N_11079,N_11307);
xor U11841 (N_11841,N_11049,N_11110);
xnor U11842 (N_11842,N_11424,N_11311);
and U11843 (N_11843,N_11333,N_11387);
and U11844 (N_11844,N_11320,N_11201);
xnor U11845 (N_11845,N_11198,N_11322);
nand U11846 (N_11846,N_11152,N_11181);
nor U11847 (N_11847,N_11257,N_11253);
nor U11848 (N_11848,N_11497,N_11201);
nand U11849 (N_11849,N_11460,N_11183);
xor U11850 (N_11850,N_11462,N_11027);
or U11851 (N_11851,N_11297,N_11347);
or U11852 (N_11852,N_11011,N_11067);
nand U11853 (N_11853,N_11100,N_11306);
nor U11854 (N_11854,N_11032,N_11370);
or U11855 (N_11855,N_11085,N_11116);
or U11856 (N_11856,N_11363,N_11109);
or U11857 (N_11857,N_11374,N_11493);
or U11858 (N_11858,N_11298,N_11366);
nor U11859 (N_11859,N_11025,N_11386);
nor U11860 (N_11860,N_11260,N_11052);
or U11861 (N_11861,N_11159,N_11322);
nand U11862 (N_11862,N_11137,N_11210);
or U11863 (N_11863,N_11091,N_11423);
xnor U11864 (N_11864,N_11384,N_11472);
nor U11865 (N_11865,N_11259,N_11222);
and U11866 (N_11866,N_11010,N_11380);
or U11867 (N_11867,N_11198,N_11046);
nand U11868 (N_11868,N_11074,N_11315);
nor U11869 (N_11869,N_11425,N_11029);
and U11870 (N_11870,N_11359,N_11312);
xnor U11871 (N_11871,N_11026,N_11226);
nand U11872 (N_11872,N_11098,N_11251);
nand U11873 (N_11873,N_11008,N_11038);
nand U11874 (N_11874,N_11040,N_11433);
or U11875 (N_11875,N_11495,N_11359);
or U11876 (N_11876,N_11297,N_11264);
or U11877 (N_11877,N_11166,N_11208);
or U11878 (N_11878,N_11151,N_11347);
or U11879 (N_11879,N_11368,N_11394);
nor U11880 (N_11880,N_11013,N_11080);
or U11881 (N_11881,N_11449,N_11269);
and U11882 (N_11882,N_11021,N_11292);
nor U11883 (N_11883,N_11039,N_11291);
or U11884 (N_11884,N_11116,N_11151);
xor U11885 (N_11885,N_11150,N_11264);
and U11886 (N_11886,N_11106,N_11273);
nand U11887 (N_11887,N_11387,N_11219);
or U11888 (N_11888,N_11173,N_11453);
and U11889 (N_11889,N_11275,N_11163);
or U11890 (N_11890,N_11237,N_11048);
xor U11891 (N_11891,N_11127,N_11185);
or U11892 (N_11892,N_11447,N_11287);
and U11893 (N_11893,N_11477,N_11254);
or U11894 (N_11894,N_11004,N_11436);
nor U11895 (N_11895,N_11239,N_11322);
or U11896 (N_11896,N_11006,N_11083);
nor U11897 (N_11897,N_11423,N_11364);
nand U11898 (N_11898,N_11053,N_11305);
nand U11899 (N_11899,N_11132,N_11021);
or U11900 (N_11900,N_11360,N_11483);
nand U11901 (N_11901,N_11440,N_11322);
xnor U11902 (N_11902,N_11140,N_11039);
nand U11903 (N_11903,N_11188,N_11372);
nor U11904 (N_11904,N_11134,N_11056);
nor U11905 (N_11905,N_11212,N_11478);
nor U11906 (N_11906,N_11099,N_11051);
and U11907 (N_11907,N_11415,N_11036);
xor U11908 (N_11908,N_11211,N_11183);
nor U11909 (N_11909,N_11244,N_11480);
xnor U11910 (N_11910,N_11166,N_11289);
nand U11911 (N_11911,N_11458,N_11208);
nand U11912 (N_11912,N_11182,N_11106);
or U11913 (N_11913,N_11482,N_11091);
nand U11914 (N_11914,N_11171,N_11271);
nand U11915 (N_11915,N_11271,N_11343);
nor U11916 (N_11916,N_11423,N_11388);
and U11917 (N_11917,N_11133,N_11307);
nor U11918 (N_11918,N_11101,N_11462);
nand U11919 (N_11919,N_11434,N_11202);
or U11920 (N_11920,N_11198,N_11246);
and U11921 (N_11921,N_11229,N_11344);
xnor U11922 (N_11922,N_11492,N_11356);
and U11923 (N_11923,N_11048,N_11415);
or U11924 (N_11924,N_11013,N_11419);
nor U11925 (N_11925,N_11241,N_11159);
and U11926 (N_11926,N_11429,N_11056);
or U11927 (N_11927,N_11493,N_11242);
nor U11928 (N_11928,N_11343,N_11188);
nor U11929 (N_11929,N_11124,N_11465);
and U11930 (N_11930,N_11437,N_11459);
or U11931 (N_11931,N_11493,N_11241);
xor U11932 (N_11932,N_11443,N_11476);
xnor U11933 (N_11933,N_11318,N_11072);
xor U11934 (N_11934,N_11287,N_11418);
nand U11935 (N_11935,N_11305,N_11379);
xnor U11936 (N_11936,N_11188,N_11495);
or U11937 (N_11937,N_11380,N_11303);
and U11938 (N_11938,N_11255,N_11185);
or U11939 (N_11939,N_11170,N_11493);
nand U11940 (N_11940,N_11128,N_11000);
nand U11941 (N_11941,N_11019,N_11109);
nor U11942 (N_11942,N_11017,N_11306);
xnor U11943 (N_11943,N_11466,N_11010);
nand U11944 (N_11944,N_11077,N_11121);
nor U11945 (N_11945,N_11149,N_11346);
or U11946 (N_11946,N_11334,N_11082);
nand U11947 (N_11947,N_11035,N_11299);
nor U11948 (N_11948,N_11059,N_11305);
or U11949 (N_11949,N_11068,N_11251);
xor U11950 (N_11950,N_11268,N_11489);
nor U11951 (N_11951,N_11401,N_11209);
nor U11952 (N_11952,N_11082,N_11107);
nand U11953 (N_11953,N_11211,N_11408);
xor U11954 (N_11954,N_11022,N_11235);
xor U11955 (N_11955,N_11019,N_11198);
and U11956 (N_11956,N_11005,N_11488);
or U11957 (N_11957,N_11013,N_11001);
nand U11958 (N_11958,N_11293,N_11149);
nor U11959 (N_11959,N_11444,N_11087);
and U11960 (N_11960,N_11057,N_11471);
xor U11961 (N_11961,N_11136,N_11157);
or U11962 (N_11962,N_11081,N_11090);
or U11963 (N_11963,N_11134,N_11100);
nand U11964 (N_11964,N_11102,N_11385);
or U11965 (N_11965,N_11026,N_11231);
nand U11966 (N_11966,N_11092,N_11108);
nor U11967 (N_11967,N_11334,N_11029);
and U11968 (N_11968,N_11316,N_11123);
or U11969 (N_11969,N_11325,N_11237);
nor U11970 (N_11970,N_11112,N_11225);
nor U11971 (N_11971,N_11245,N_11400);
nand U11972 (N_11972,N_11335,N_11044);
nand U11973 (N_11973,N_11296,N_11344);
nand U11974 (N_11974,N_11467,N_11012);
xor U11975 (N_11975,N_11424,N_11269);
and U11976 (N_11976,N_11303,N_11325);
or U11977 (N_11977,N_11279,N_11425);
nor U11978 (N_11978,N_11080,N_11437);
or U11979 (N_11979,N_11081,N_11100);
and U11980 (N_11980,N_11422,N_11012);
xor U11981 (N_11981,N_11459,N_11472);
and U11982 (N_11982,N_11119,N_11430);
or U11983 (N_11983,N_11149,N_11336);
nand U11984 (N_11984,N_11240,N_11445);
xor U11985 (N_11985,N_11251,N_11333);
nor U11986 (N_11986,N_11026,N_11352);
nand U11987 (N_11987,N_11134,N_11120);
or U11988 (N_11988,N_11199,N_11496);
nor U11989 (N_11989,N_11432,N_11444);
nand U11990 (N_11990,N_11018,N_11245);
nand U11991 (N_11991,N_11019,N_11482);
nor U11992 (N_11992,N_11194,N_11398);
nor U11993 (N_11993,N_11219,N_11434);
and U11994 (N_11994,N_11209,N_11276);
and U11995 (N_11995,N_11364,N_11269);
nand U11996 (N_11996,N_11087,N_11288);
nand U11997 (N_11997,N_11159,N_11472);
nand U11998 (N_11998,N_11356,N_11272);
or U11999 (N_11999,N_11155,N_11148);
nor U12000 (N_12000,N_11947,N_11966);
nand U12001 (N_12001,N_11528,N_11746);
xnor U12002 (N_12002,N_11571,N_11777);
xnor U12003 (N_12003,N_11896,N_11902);
xnor U12004 (N_12004,N_11523,N_11863);
xnor U12005 (N_12005,N_11520,N_11737);
xor U12006 (N_12006,N_11699,N_11789);
nand U12007 (N_12007,N_11706,N_11654);
nand U12008 (N_12008,N_11736,N_11908);
nand U12009 (N_12009,N_11683,N_11953);
or U12010 (N_12010,N_11888,N_11549);
nand U12011 (N_12011,N_11828,N_11677);
xnor U12012 (N_12012,N_11807,N_11997);
nor U12013 (N_12013,N_11821,N_11951);
nor U12014 (N_12014,N_11591,N_11916);
nor U12015 (N_12015,N_11536,N_11624);
nor U12016 (N_12016,N_11765,N_11854);
and U12017 (N_12017,N_11867,N_11885);
or U12018 (N_12018,N_11598,N_11511);
nor U12019 (N_12019,N_11954,N_11566);
xnor U12020 (N_12020,N_11880,N_11838);
or U12021 (N_12021,N_11559,N_11871);
and U12022 (N_12022,N_11592,N_11690);
nor U12023 (N_12023,N_11529,N_11812);
xor U12024 (N_12024,N_11974,N_11534);
xnor U12025 (N_12025,N_11819,N_11643);
nor U12026 (N_12026,N_11776,N_11538);
xnor U12027 (N_12027,N_11585,N_11873);
and U12028 (N_12028,N_11904,N_11719);
nand U12029 (N_12029,N_11785,N_11744);
or U12030 (N_12030,N_11957,N_11704);
nand U12031 (N_12031,N_11940,N_11717);
and U12032 (N_12032,N_11769,N_11797);
nor U12033 (N_12033,N_11970,N_11936);
and U12034 (N_12034,N_11517,N_11803);
nor U12035 (N_12035,N_11927,N_11600);
nor U12036 (N_12036,N_11682,N_11733);
nand U12037 (N_12037,N_11955,N_11647);
nand U12038 (N_12038,N_11894,N_11675);
nand U12039 (N_12039,N_11531,N_11987);
xnor U12040 (N_12040,N_11749,N_11623);
nand U12041 (N_12041,N_11800,N_11928);
xor U12042 (N_12042,N_11781,N_11962);
xor U12043 (N_12043,N_11790,N_11553);
xnor U12044 (N_12044,N_11825,N_11626);
nor U12045 (N_12045,N_11978,N_11676);
nor U12046 (N_12046,N_11935,N_11762);
xor U12047 (N_12047,N_11735,N_11831);
nor U12048 (N_12048,N_11969,N_11979);
nand U12049 (N_12049,N_11988,N_11607);
nor U12050 (N_12050,N_11716,N_11614);
nor U12051 (N_12051,N_11581,N_11778);
or U12052 (N_12052,N_11973,N_11664);
xnor U12053 (N_12053,N_11836,N_11758);
and U12054 (N_12054,N_11686,N_11731);
or U12055 (N_12055,N_11681,N_11535);
nand U12056 (N_12056,N_11640,N_11891);
nor U12057 (N_12057,N_11862,N_11567);
or U12058 (N_12058,N_11843,N_11972);
xor U12059 (N_12059,N_11665,N_11542);
or U12060 (N_12060,N_11701,N_11564);
or U12061 (N_12061,N_11563,N_11558);
or U12062 (N_12062,N_11939,N_11981);
xor U12063 (N_12063,N_11703,N_11864);
and U12064 (N_12064,N_11856,N_11850);
or U12065 (N_12065,N_11922,N_11810);
nor U12066 (N_12066,N_11832,N_11773);
xor U12067 (N_12067,N_11650,N_11985);
xnor U12068 (N_12068,N_11527,N_11726);
xnor U12069 (N_12069,N_11829,N_11872);
nor U12070 (N_12070,N_11753,N_11992);
xnor U12071 (N_12071,N_11898,N_11780);
or U12072 (N_12072,N_11619,N_11900);
and U12073 (N_12073,N_11949,N_11674);
or U12074 (N_12074,N_11795,N_11993);
and U12075 (N_12075,N_11760,N_11794);
nand U12076 (N_12076,N_11580,N_11646);
nand U12077 (N_12077,N_11596,N_11708);
xnor U12078 (N_12078,N_11818,N_11930);
and U12079 (N_12079,N_11870,N_11521);
xnor U12080 (N_12080,N_11608,N_11764);
nand U12081 (N_12081,N_11815,N_11657);
nor U12082 (N_12082,N_11501,N_11689);
xnor U12083 (N_12083,N_11560,N_11956);
nor U12084 (N_12084,N_11986,N_11967);
xor U12085 (N_12085,N_11541,N_11605);
nor U12086 (N_12086,N_11965,N_11813);
and U12087 (N_12087,N_11915,N_11857);
nor U12088 (N_12088,N_11865,N_11835);
and U12089 (N_12089,N_11628,N_11620);
xor U12090 (N_12090,N_11933,N_11866);
xnor U12091 (N_12091,N_11621,N_11526);
or U12092 (N_12092,N_11722,N_11505);
nand U12093 (N_12093,N_11879,N_11588);
nor U12094 (N_12094,N_11663,N_11757);
nand U12095 (N_12095,N_11651,N_11806);
or U12096 (N_12096,N_11705,N_11684);
nor U12097 (N_12097,N_11941,N_11811);
nand U12098 (N_12098,N_11590,N_11846);
and U12099 (N_12099,N_11878,N_11672);
or U12100 (N_12100,N_11509,N_11723);
xnor U12101 (N_12101,N_11653,N_11556);
or U12102 (N_12102,N_11976,N_11959);
nor U12103 (N_12103,N_11788,N_11575);
and U12104 (N_12104,N_11639,N_11612);
nand U12105 (N_12105,N_11855,N_11796);
nand U12106 (N_12106,N_11604,N_11923);
xor U12107 (N_12107,N_11804,N_11515);
xnor U12108 (N_12108,N_11938,N_11817);
or U12109 (N_12109,N_11884,N_11968);
xor U12110 (N_12110,N_11874,N_11645);
xnor U12111 (N_12111,N_11595,N_11768);
xnor U12112 (N_12112,N_11715,N_11673);
xor U12113 (N_12113,N_11518,N_11950);
nand U12114 (N_12114,N_11724,N_11748);
and U12115 (N_12115,N_11680,N_11917);
xnor U12116 (N_12116,N_11911,N_11635);
nor U12117 (N_12117,N_11887,N_11519);
nor U12118 (N_12118,N_11539,N_11603);
nor U12119 (N_12119,N_11814,N_11995);
or U12120 (N_12120,N_11696,N_11734);
nor U12121 (N_12121,N_11514,N_11990);
nor U12122 (N_12122,N_11783,N_11739);
nand U12123 (N_12123,N_11943,N_11532);
or U12124 (N_12124,N_11732,N_11573);
nand U12125 (N_12125,N_11617,N_11895);
and U12126 (N_12126,N_11569,N_11550);
and U12127 (N_12127,N_11709,N_11533);
xor U12128 (N_12128,N_11711,N_11606);
or U12129 (N_12129,N_11944,N_11537);
or U12130 (N_12130,N_11671,N_11741);
xnor U12131 (N_12131,N_11661,N_11989);
and U12132 (N_12132,N_11668,N_11510);
and U12133 (N_12133,N_11525,N_11721);
or U12134 (N_12134,N_11752,N_11679);
nor U12135 (N_12135,N_11840,N_11738);
xor U12136 (N_12136,N_11658,N_11574);
xor U12137 (N_12137,N_11925,N_11586);
nand U12138 (N_12138,N_11602,N_11907);
nor U12139 (N_12139,N_11755,N_11839);
nor U12140 (N_12140,N_11984,N_11975);
xnor U12141 (N_12141,N_11861,N_11912);
or U12142 (N_12142,N_11561,N_11655);
and U12143 (N_12143,N_11971,N_11568);
nand U12144 (N_12144,N_11552,N_11641);
nand U12145 (N_12145,N_11636,N_11868);
or U12146 (N_12146,N_11877,N_11890);
nor U12147 (N_12147,N_11714,N_11998);
nand U12148 (N_12148,N_11577,N_11851);
and U12149 (N_12149,N_11876,N_11827);
or U12150 (N_12150,N_11889,N_11599);
and U12151 (N_12151,N_11587,N_11906);
nand U12152 (N_12152,N_11784,N_11824);
nor U12153 (N_12153,N_11530,N_11615);
nor U12154 (N_12154,N_11662,N_11913);
xnor U12155 (N_12155,N_11743,N_11751);
and U12156 (N_12156,N_11772,N_11793);
or U12157 (N_12157,N_11801,N_11627);
and U12158 (N_12158,N_11934,N_11852);
nand U12159 (N_12159,N_11660,N_11594);
nand U12160 (N_12160,N_11634,N_11670);
xnor U12161 (N_12161,N_11618,N_11792);
and U12162 (N_12162,N_11656,N_11763);
nand U12163 (N_12163,N_11593,N_11918);
and U12164 (N_12164,N_11816,N_11754);
nor U12165 (N_12165,N_11562,N_11875);
or U12166 (N_12166,N_11892,N_11834);
nand U12167 (N_12167,N_11958,N_11774);
xnor U12168 (N_12168,N_11910,N_11767);
xor U12169 (N_12169,N_11691,N_11782);
and U12170 (N_12170,N_11808,N_11710);
nand U12171 (N_12171,N_11946,N_11678);
nor U12172 (N_12172,N_11557,N_11725);
nand U12173 (N_12173,N_11937,N_11921);
xnor U12174 (N_12174,N_11728,N_11747);
nand U12175 (N_12175,N_11848,N_11799);
nand U12176 (N_12176,N_11688,N_11630);
nor U12177 (N_12177,N_11637,N_11631);
or U12178 (N_12178,N_11932,N_11977);
xnor U12179 (N_12179,N_11584,N_11610);
or U12180 (N_12180,N_11698,N_11504);
xnor U12181 (N_12181,N_11695,N_11718);
or U12182 (N_12182,N_11632,N_11522);
xnor U12183 (N_12183,N_11576,N_11512);
nor U12184 (N_12184,N_11730,N_11565);
nor U12185 (N_12185,N_11707,N_11648);
and U12186 (N_12186,N_11853,N_11609);
and U12187 (N_12187,N_11572,N_11882);
nand U12188 (N_12188,N_11583,N_11826);
xor U12189 (N_12189,N_11500,N_11545);
nand U12190 (N_12190,N_11555,N_11540);
nand U12191 (N_12191,N_11761,N_11644);
and U12192 (N_12192,N_11845,N_11597);
nand U12193 (N_12193,N_11809,N_11770);
or U12194 (N_12194,N_11613,N_11750);
nand U12195 (N_12195,N_11860,N_11775);
xor U12196 (N_12196,N_11914,N_11638);
or U12197 (N_12197,N_11897,N_11837);
and U12198 (N_12198,N_11616,N_11508);
nand U12199 (N_12199,N_11948,N_11822);
nor U12200 (N_12200,N_11920,N_11859);
or U12201 (N_12201,N_11983,N_11841);
nand U12202 (N_12202,N_11830,N_11692);
and U12203 (N_12203,N_11554,N_11759);
nor U12204 (N_12204,N_11929,N_11712);
or U12205 (N_12205,N_11622,N_11931);
or U12206 (N_12206,N_11903,N_11694);
or U12207 (N_12207,N_11516,N_11766);
and U12208 (N_12208,N_11771,N_11963);
or U12209 (N_12209,N_11548,N_11729);
and U12210 (N_12210,N_11524,N_11601);
xor U12211 (N_12211,N_11996,N_11544);
and U12212 (N_12212,N_11507,N_11960);
nand U12213 (N_12213,N_11652,N_11700);
or U12214 (N_12214,N_11961,N_11551);
and U12215 (N_12215,N_11820,N_11582);
and U12216 (N_12216,N_11513,N_11849);
nor U12217 (N_12217,N_11740,N_11720);
or U12218 (N_12218,N_11858,N_11926);
and U12219 (N_12219,N_11802,N_11886);
nand U12220 (N_12220,N_11629,N_11924);
nand U12221 (N_12221,N_11503,N_11611);
or U12222 (N_12222,N_11899,N_11543);
and U12223 (N_12223,N_11506,N_11697);
nor U12224 (N_12224,N_11942,N_11666);
and U12225 (N_12225,N_11844,N_11756);
nor U12226 (N_12226,N_11847,N_11786);
nor U12227 (N_12227,N_11669,N_11625);
xor U12228 (N_12228,N_11869,N_11883);
or U12229 (N_12229,N_11579,N_11881);
xor U12230 (N_12230,N_11994,N_11578);
xnor U12231 (N_12231,N_11589,N_11687);
nand U12232 (N_12232,N_11964,N_11702);
xnor U12233 (N_12233,N_11991,N_11745);
nor U12234 (N_12234,N_11570,N_11547);
or U12235 (N_12235,N_11919,N_11779);
and U12236 (N_12236,N_11893,N_11909);
nand U12237 (N_12237,N_11667,N_11659);
or U12238 (N_12238,N_11791,N_11952);
nand U12239 (N_12239,N_11945,N_11842);
or U12240 (N_12240,N_11693,N_11823);
xor U12241 (N_12241,N_11685,N_11742);
nor U12242 (N_12242,N_11633,N_11502);
or U12243 (N_12243,N_11642,N_11999);
xnor U12244 (N_12244,N_11805,N_11833);
and U12245 (N_12245,N_11787,N_11905);
nor U12246 (N_12246,N_11727,N_11980);
nand U12247 (N_12247,N_11798,N_11649);
and U12248 (N_12248,N_11546,N_11713);
or U12249 (N_12249,N_11982,N_11901);
or U12250 (N_12250,N_11736,N_11615);
nand U12251 (N_12251,N_11841,N_11510);
xor U12252 (N_12252,N_11552,N_11606);
xnor U12253 (N_12253,N_11977,N_11548);
xnor U12254 (N_12254,N_11594,N_11663);
nor U12255 (N_12255,N_11966,N_11926);
and U12256 (N_12256,N_11719,N_11985);
nor U12257 (N_12257,N_11683,N_11962);
or U12258 (N_12258,N_11806,N_11925);
nor U12259 (N_12259,N_11798,N_11888);
or U12260 (N_12260,N_11949,N_11694);
nor U12261 (N_12261,N_11762,N_11719);
nor U12262 (N_12262,N_11965,N_11814);
xnor U12263 (N_12263,N_11622,N_11651);
and U12264 (N_12264,N_11767,N_11952);
xnor U12265 (N_12265,N_11621,N_11628);
nor U12266 (N_12266,N_11716,N_11692);
nor U12267 (N_12267,N_11877,N_11593);
nor U12268 (N_12268,N_11999,N_11943);
and U12269 (N_12269,N_11905,N_11817);
nor U12270 (N_12270,N_11572,N_11842);
xor U12271 (N_12271,N_11833,N_11773);
xor U12272 (N_12272,N_11697,N_11877);
and U12273 (N_12273,N_11559,N_11758);
nand U12274 (N_12274,N_11729,N_11657);
or U12275 (N_12275,N_11825,N_11932);
nor U12276 (N_12276,N_11948,N_11726);
or U12277 (N_12277,N_11753,N_11630);
nor U12278 (N_12278,N_11534,N_11745);
or U12279 (N_12279,N_11582,N_11909);
nor U12280 (N_12280,N_11737,N_11637);
xor U12281 (N_12281,N_11505,N_11947);
xnor U12282 (N_12282,N_11901,N_11539);
xnor U12283 (N_12283,N_11639,N_11713);
nor U12284 (N_12284,N_11562,N_11865);
xnor U12285 (N_12285,N_11985,N_11764);
or U12286 (N_12286,N_11954,N_11752);
and U12287 (N_12287,N_11602,N_11816);
or U12288 (N_12288,N_11927,N_11893);
or U12289 (N_12289,N_11983,N_11892);
nand U12290 (N_12290,N_11616,N_11805);
nor U12291 (N_12291,N_11581,N_11754);
nor U12292 (N_12292,N_11947,N_11986);
nor U12293 (N_12293,N_11839,N_11583);
nand U12294 (N_12294,N_11620,N_11640);
nor U12295 (N_12295,N_11906,N_11851);
and U12296 (N_12296,N_11772,N_11754);
nand U12297 (N_12297,N_11892,N_11643);
and U12298 (N_12298,N_11969,N_11706);
nand U12299 (N_12299,N_11675,N_11772);
nand U12300 (N_12300,N_11999,N_11909);
nor U12301 (N_12301,N_11837,N_11765);
xor U12302 (N_12302,N_11911,N_11915);
xor U12303 (N_12303,N_11540,N_11673);
and U12304 (N_12304,N_11739,N_11503);
or U12305 (N_12305,N_11879,N_11835);
or U12306 (N_12306,N_11757,N_11956);
nor U12307 (N_12307,N_11773,N_11783);
nand U12308 (N_12308,N_11706,N_11885);
or U12309 (N_12309,N_11527,N_11701);
nor U12310 (N_12310,N_11727,N_11531);
nor U12311 (N_12311,N_11979,N_11783);
xnor U12312 (N_12312,N_11663,N_11679);
nand U12313 (N_12313,N_11765,N_11902);
nor U12314 (N_12314,N_11964,N_11845);
nand U12315 (N_12315,N_11728,N_11681);
and U12316 (N_12316,N_11742,N_11778);
xnor U12317 (N_12317,N_11767,N_11914);
nand U12318 (N_12318,N_11539,N_11773);
nor U12319 (N_12319,N_11684,N_11916);
and U12320 (N_12320,N_11624,N_11543);
nand U12321 (N_12321,N_11642,N_11824);
nand U12322 (N_12322,N_11687,N_11665);
or U12323 (N_12323,N_11847,N_11596);
nand U12324 (N_12324,N_11690,N_11688);
nor U12325 (N_12325,N_11933,N_11767);
and U12326 (N_12326,N_11616,N_11828);
and U12327 (N_12327,N_11871,N_11683);
nand U12328 (N_12328,N_11691,N_11611);
nand U12329 (N_12329,N_11726,N_11923);
nor U12330 (N_12330,N_11603,N_11614);
nand U12331 (N_12331,N_11644,N_11821);
and U12332 (N_12332,N_11604,N_11779);
xor U12333 (N_12333,N_11855,N_11617);
nand U12334 (N_12334,N_11795,N_11794);
or U12335 (N_12335,N_11667,N_11710);
nor U12336 (N_12336,N_11725,N_11863);
or U12337 (N_12337,N_11989,N_11809);
nor U12338 (N_12338,N_11502,N_11773);
xnor U12339 (N_12339,N_11642,N_11945);
xor U12340 (N_12340,N_11643,N_11569);
nor U12341 (N_12341,N_11657,N_11637);
or U12342 (N_12342,N_11902,N_11972);
and U12343 (N_12343,N_11715,N_11900);
or U12344 (N_12344,N_11801,N_11763);
xor U12345 (N_12345,N_11698,N_11878);
and U12346 (N_12346,N_11590,N_11912);
xor U12347 (N_12347,N_11507,N_11845);
or U12348 (N_12348,N_11548,N_11986);
nand U12349 (N_12349,N_11794,N_11770);
or U12350 (N_12350,N_11762,N_11859);
nand U12351 (N_12351,N_11672,N_11766);
and U12352 (N_12352,N_11963,N_11757);
nor U12353 (N_12353,N_11874,N_11949);
and U12354 (N_12354,N_11906,N_11810);
nor U12355 (N_12355,N_11504,N_11549);
and U12356 (N_12356,N_11601,N_11605);
nand U12357 (N_12357,N_11643,N_11943);
nor U12358 (N_12358,N_11895,N_11691);
nand U12359 (N_12359,N_11836,N_11792);
or U12360 (N_12360,N_11852,N_11935);
nand U12361 (N_12361,N_11986,N_11867);
and U12362 (N_12362,N_11776,N_11619);
or U12363 (N_12363,N_11584,N_11691);
xor U12364 (N_12364,N_11578,N_11551);
nor U12365 (N_12365,N_11938,N_11841);
or U12366 (N_12366,N_11749,N_11768);
xor U12367 (N_12367,N_11743,N_11998);
xor U12368 (N_12368,N_11587,N_11938);
nand U12369 (N_12369,N_11521,N_11687);
or U12370 (N_12370,N_11824,N_11968);
or U12371 (N_12371,N_11527,N_11504);
nor U12372 (N_12372,N_11610,N_11887);
xnor U12373 (N_12373,N_11828,N_11755);
nand U12374 (N_12374,N_11673,N_11567);
nand U12375 (N_12375,N_11823,N_11642);
nand U12376 (N_12376,N_11662,N_11888);
nand U12377 (N_12377,N_11664,N_11592);
or U12378 (N_12378,N_11834,N_11558);
and U12379 (N_12379,N_11778,N_11976);
or U12380 (N_12380,N_11993,N_11977);
xor U12381 (N_12381,N_11978,N_11748);
or U12382 (N_12382,N_11603,N_11949);
or U12383 (N_12383,N_11963,N_11615);
nor U12384 (N_12384,N_11823,N_11981);
nand U12385 (N_12385,N_11777,N_11501);
nor U12386 (N_12386,N_11678,N_11902);
xor U12387 (N_12387,N_11646,N_11879);
and U12388 (N_12388,N_11909,N_11529);
and U12389 (N_12389,N_11976,N_11902);
nand U12390 (N_12390,N_11706,N_11763);
nand U12391 (N_12391,N_11538,N_11856);
nor U12392 (N_12392,N_11676,N_11977);
nor U12393 (N_12393,N_11879,N_11682);
and U12394 (N_12394,N_11712,N_11665);
nor U12395 (N_12395,N_11710,N_11821);
nor U12396 (N_12396,N_11641,N_11804);
or U12397 (N_12397,N_11666,N_11937);
or U12398 (N_12398,N_11633,N_11781);
nand U12399 (N_12399,N_11872,N_11933);
nor U12400 (N_12400,N_11726,N_11673);
nand U12401 (N_12401,N_11860,N_11511);
nand U12402 (N_12402,N_11737,N_11857);
and U12403 (N_12403,N_11759,N_11960);
and U12404 (N_12404,N_11680,N_11819);
xor U12405 (N_12405,N_11978,N_11842);
nor U12406 (N_12406,N_11787,N_11689);
nand U12407 (N_12407,N_11641,N_11568);
nand U12408 (N_12408,N_11702,N_11546);
xor U12409 (N_12409,N_11723,N_11569);
and U12410 (N_12410,N_11785,N_11933);
xor U12411 (N_12411,N_11982,N_11587);
xor U12412 (N_12412,N_11784,N_11878);
and U12413 (N_12413,N_11968,N_11541);
xnor U12414 (N_12414,N_11922,N_11820);
and U12415 (N_12415,N_11723,N_11969);
nand U12416 (N_12416,N_11638,N_11682);
and U12417 (N_12417,N_11876,N_11691);
nand U12418 (N_12418,N_11565,N_11641);
nand U12419 (N_12419,N_11673,N_11806);
xor U12420 (N_12420,N_11983,N_11862);
and U12421 (N_12421,N_11743,N_11888);
xor U12422 (N_12422,N_11504,N_11821);
or U12423 (N_12423,N_11628,N_11638);
xor U12424 (N_12424,N_11974,N_11855);
xor U12425 (N_12425,N_11944,N_11747);
or U12426 (N_12426,N_11614,N_11535);
nand U12427 (N_12427,N_11832,N_11690);
or U12428 (N_12428,N_11841,N_11951);
xor U12429 (N_12429,N_11642,N_11965);
xnor U12430 (N_12430,N_11956,N_11860);
nand U12431 (N_12431,N_11976,N_11754);
or U12432 (N_12432,N_11695,N_11531);
nand U12433 (N_12433,N_11786,N_11889);
and U12434 (N_12434,N_11580,N_11918);
xnor U12435 (N_12435,N_11560,N_11515);
or U12436 (N_12436,N_11850,N_11640);
nand U12437 (N_12437,N_11702,N_11730);
nand U12438 (N_12438,N_11855,N_11559);
nand U12439 (N_12439,N_11590,N_11571);
xor U12440 (N_12440,N_11698,N_11753);
and U12441 (N_12441,N_11629,N_11591);
or U12442 (N_12442,N_11677,N_11741);
xor U12443 (N_12443,N_11514,N_11537);
nor U12444 (N_12444,N_11631,N_11972);
or U12445 (N_12445,N_11724,N_11737);
nand U12446 (N_12446,N_11715,N_11935);
nand U12447 (N_12447,N_11774,N_11718);
and U12448 (N_12448,N_11802,N_11676);
and U12449 (N_12449,N_11883,N_11731);
and U12450 (N_12450,N_11547,N_11744);
nand U12451 (N_12451,N_11611,N_11782);
and U12452 (N_12452,N_11969,N_11857);
and U12453 (N_12453,N_11628,N_11635);
xnor U12454 (N_12454,N_11860,N_11558);
nor U12455 (N_12455,N_11551,N_11705);
nand U12456 (N_12456,N_11803,N_11928);
nor U12457 (N_12457,N_11605,N_11986);
nand U12458 (N_12458,N_11653,N_11510);
or U12459 (N_12459,N_11925,N_11685);
or U12460 (N_12460,N_11549,N_11934);
or U12461 (N_12461,N_11991,N_11689);
and U12462 (N_12462,N_11774,N_11637);
or U12463 (N_12463,N_11695,N_11843);
and U12464 (N_12464,N_11750,N_11600);
and U12465 (N_12465,N_11943,N_11575);
xnor U12466 (N_12466,N_11532,N_11995);
xnor U12467 (N_12467,N_11842,N_11561);
or U12468 (N_12468,N_11987,N_11954);
and U12469 (N_12469,N_11958,N_11745);
or U12470 (N_12470,N_11720,N_11996);
and U12471 (N_12471,N_11736,N_11776);
nand U12472 (N_12472,N_11660,N_11653);
nor U12473 (N_12473,N_11892,N_11733);
xnor U12474 (N_12474,N_11577,N_11951);
xor U12475 (N_12475,N_11668,N_11545);
nor U12476 (N_12476,N_11538,N_11610);
nor U12477 (N_12477,N_11648,N_11779);
or U12478 (N_12478,N_11728,N_11691);
and U12479 (N_12479,N_11829,N_11837);
nand U12480 (N_12480,N_11610,N_11896);
nand U12481 (N_12481,N_11755,N_11826);
and U12482 (N_12482,N_11616,N_11870);
xor U12483 (N_12483,N_11707,N_11729);
or U12484 (N_12484,N_11804,N_11796);
nor U12485 (N_12485,N_11897,N_11560);
and U12486 (N_12486,N_11957,N_11919);
and U12487 (N_12487,N_11778,N_11708);
xor U12488 (N_12488,N_11787,N_11593);
and U12489 (N_12489,N_11866,N_11857);
nor U12490 (N_12490,N_11550,N_11874);
xnor U12491 (N_12491,N_11549,N_11647);
nor U12492 (N_12492,N_11795,N_11740);
and U12493 (N_12493,N_11600,N_11896);
and U12494 (N_12494,N_11807,N_11906);
and U12495 (N_12495,N_11926,N_11701);
xnor U12496 (N_12496,N_11878,N_11688);
xor U12497 (N_12497,N_11688,N_11903);
or U12498 (N_12498,N_11581,N_11731);
nor U12499 (N_12499,N_11873,N_11887);
xnor U12500 (N_12500,N_12038,N_12481);
and U12501 (N_12501,N_12201,N_12160);
xor U12502 (N_12502,N_12475,N_12424);
xnor U12503 (N_12503,N_12295,N_12178);
or U12504 (N_12504,N_12110,N_12095);
and U12505 (N_12505,N_12252,N_12001);
and U12506 (N_12506,N_12230,N_12368);
nand U12507 (N_12507,N_12224,N_12087);
nor U12508 (N_12508,N_12044,N_12471);
or U12509 (N_12509,N_12444,N_12304);
xnor U12510 (N_12510,N_12359,N_12292);
xnor U12511 (N_12511,N_12243,N_12399);
nand U12512 (N_12512,N_12176,N_12460);
xnor U12513 (N_12513,N_12362,N_12188);
or U12514 (N_12514,N_12119,N_12045);
nand U12515 (N_12515,N_12375,N_12098);
nor U12516 (N_12516,N_12482,N_12476);
nand U12517 (N_12517,N_12318,N_12020);
xnor U12518 (N_12518,N_12313,N_12128);
nor U12519 (N_12519,N_12129,N_12299);
or U12520 (N_12520,N_12251,N_12382);
xor U12521 (N_12521,N_12259,N_12089);
or U12522 (N_12522,N_12076,N_12074);
nor U12523 (N_12523,N_12221,N_12497);
and U12524 (N_12524,N_12316,N_12369);
and U12525 (N_12525,N_12190,N_12101);
or U12526 (N_12526,N_12120,N_12172);
nor U12527 (N_12527,N_12083,N_12344);
or U12528 (N_12528,N_12385,N_12326);
nor U12529 (N_12529,N_12144,N_12389);
and U12530 (N_12530,N_12446,N_12216);
nand U12531 (N_12531,N_12409,N_12454);
or U12532 (N_12532,N_12191,N_12043);
or U12533 (N_12533,N_12315,N_12492);
or U12534 (N_12534,N_12012,N_12264);
or U12535 (N_12535,N_12240,N_12167);
or U12536 (N_12536,N_12286,N_12478);
nor U12537 (N_12537,N_12418,N_12195);
nand U12538 (N_12538,N_12103,N_12263);
nand U12539 (N_12539,N_12238,N_12206);
nor U12540 (N_12540,N_12467,N_12213);
and U12541 (N_12541,N_12016,N_12474);
and U12542 (N_12542,N_12331,N_12143);
nand U12543 (N_12543,N_12353,N_12033);
nor U12544 (N_12544,N_12047,N_12489);
and U12545 (N_12545,N_12072,N_12107);
or U12546 (N_12546,N_12105,N_12496);
nand U12547 (N_12547,N_12254,N_12293);
or U12548 (N_12548,N_12354,N_12180);
nor U12549 (N_12549,N_12197,N_12376);
and U12550 (N_12550,N_12408,N_12219);
nand U12551 (N_12551,N_12342,N_12077);
nor U12552 (N_12552,N_12260,N_12106);
nand U12553 (N_12553,N_12407,N_12168);
or U12554 (N_12554,N_12488,N_12395);
nand U12555 (N_12555,N_12136,N_12393);
and U12556 (N_12556,N_12388,N_12433);
nor U12557 (N_12557,N_12079,N_12123);
and U12558 (N_12558,N_12345,N_12170);
or U12559 (N_12559,N_12294,N_12413);
xnor U12560 (N_12560,N_12459,N_12035);
nor U12561 (N_12561,N_12245,N_12132);
nor U12562 (N_12562,N_12314,N_12056);
or U12563 (N_12563,N_12184,N_12466);
xnor U12564 (N_12564,N_12159,N_12411);
or U12565 (N_12565,N_12281,N_12343);
nand U12566 (N_12566,N_12085,N_12405);
nand U12567 (N_12567,N_12181,N_12270);
and U12568 (N_12568,N_12465,N_12429);
xor U12569 (N_12569,N_12464,N_12013);
xor U12570 (N_12570,N_12462,N_12147);
and U12571 (N_12571,N_12239,N_12027);
nand U12572 (N_12572,N_12302,N_12495);
or U12573 (N_12573,N_12112,N_12099);
xnor U12574 (N_12574,N_12084,N_12320);
nor U12575 (N_12575,N_12122,N_12361);
nor U12576 (N_12576,N_12059,N_12332);
and U12577 (N_12577,N_12493,N_12165);
and U12578 (N_12578,N_12447,N_12214);
and U12579 (N_12579,N_12064,N_12241);
nor U12580 (N_12580,N_12004,N_12211);
or U12581 (N_12581,N_12189,N_12058);
nand U12582 (N_12582,N_12406,N_12091);
and U12583 (N_12583,N_12068,N_12133);
xor U12584 (N_12584,N_12421,N_12031);
or U12585 (N_12585,N_12328,N_12096);
nor U12586 (N_12586,N_12307,N_12335);
and U12587 (N_12587,N_12440,N_12327);
or U12588 (N_12588,N_12480,N_12461);
and U12589 (N_12589,N_12289,N_12284);
xor U12590 (N_12590,N_12040,N_12185);
nor U12591 (N_12591,N_12111,N_12470);
nand U12592 (N_12592,N_12006,N_12257);
or U12593 (N_12593,N_12060,N_12014);
nand U12594 (N_12594,N_12055,N_12146);
nor U12595 (N_12595,N_12053,N_12126);
xnor U12596 (N_12596,N_12028,N_12486);
xor U12597 (N_12597,N_12265,N_12441);
xor U12598 (N_12598,N_12311,N_12138);
or U12599 (N_12599,N_12276,N_12403);
nand U12600 (N_12600,N_12499,N_12324);
or U12601 (N_12601,N_12435,N_12121);
and U12602 (N_12602,N_12357,N_12450);
or U12603 (N_12603,N_12155,N_12036);
and U12604 (N_12604,N_12253,N_12422);
nor U12605 (N_12605,N_12139,N_12341);
xor U12606 (N_12606,N_12391,N_12347);
or U12607 (N_12607,N_12222,N_12416);
or U12608 (N_12608,N_12337,N_12177);
xor U12609 (N_12609,N_12175,N_12434);
or U12610 (N_12610,N_12050,N_12023);
nand U12611 (N_12611,N_12140,N_12485);
or U12612 (N_12612,N_12005,N_12154);
nand U12613 (N_12613,N_12192,N_12234);
nand U12614 (N_12614,N_12237,N_12487);
nor U12615 (N_12615,N_12212,N_12017);
nand U12616 (N_12616,N_12379,N_12374);
and U12617 (N_12617,N_12007,N_12256);
nor U12618 (N_12618,N_12065,N_12080);
or U12619 (N_12619,N_12445,N_12271);
xnor U12620 (N_12620,N_12130,N_12291);
nor U12621 (N_12621,N_12372,N_12235);
nor U12622 (N_12622,N_12338,N_12458);
and U12623 (N_12623,N_12207,N_12280);
or U12624 (N_12624,N_12303,N_12498);
nor U12625 (N_12625,N_12090,N_12336);
nor U12626 (N_12626,N_12448,N_12108);
xnor U12627 (N_12627,N_12378,N_12402);
and U12628 (N_12628,N_12453,N_12456);
nor U12629 (N_12629,N_12198,N_12249);
nand U12630 (N_12630,N_12401,N_12246);
or U12631 (N_12631,N_12046,N_12350);
nand U12632 (N_12632,N_12484,N_12037);
and U12633 (N_12633,N_12003,N_12325);
nor U12634 (N_12634,N_12297,N_12386);
and U12635 (N_12635,N_12356,N_12226);
nor U12636 (N_12636,N_12000,N_12494);
xnor U12637 (N_12637,N_12363,N_12404);
and U12638 (N_12638,N_12309,N_12310);
xnor U12639 (N_12639,N_12209,N_12081);
or U12640 (N_12640,N_12164,N_12438);
nand U12641 (N_12641,N_12194,N_12118);
nand U12642 (N_12642,N_12171,N_12131);
xnor U12643 (N_12643,N_12269,N_12430);
nor U12644 (N_12644,N_12034,N_12449);
nand U12645 (N_12645,N_12329,N_12306);
or U12646 (N_12646,N_12452,N_12169);
and U12647 (N_12647,N_12082,N_12158);
and U12648 (N_12648,N_12048,N_12094);
nand U12649 (N_12649,N_12210,N_12152);
nor U12650 (N_12650,N_12199,N_12030);
and U12651 (N_12651,N_12063,N_12248);
nor U12652 (N_12652,N_12261,N_12223);
xor U12653 (N_12653,N_12109,N_12322);
nand U12654 (N_12654,N_12078,N_12145);
nor U12655 (N_12655,N_12228,N_12426);
and U12656 (N_12656,N_12351,N_12066);
nand U12657 (N_12657,N_12412,N_12032);
nor U12658 (N_12658,N_12193,N_12247);
and U12659 (N_12659,N_12420,N_12490);
and U12660 (N_12660,N_12323,N_12373);
or U12661 (N_12661,N_12062,N_12196);
xor U12662 (N_12662,N_12279,N_12266);
xor U12663 (N_12663,N_12010,N_12148);
xnor U12664 (N_12664,N_12015,N_12182);
xnor U12665 (N_12665,N_12054,N_12333);
and U12666 (N_12666,N_12300,N_12179);
nor U12667 (N_12667,N_12220,N_12437);
nand U12668 (N_12668,N_12009,N_12377);
nor U12669 (N_12669,N_12349,N_12319);
or U12670 (N_12670,N_12227,N_12419);
nor U12671 (N_12671,N_12455,N_12439);
nor U12672 (N_12672,N_12400,N_12383);
or U12673 (N_12673,N_12071,N_12039);
or U12674 (N_12674,N_12366,N_12340);
and U12675 (N_12675,N_12290,N_12092);
or U12676 (N_12676,N_12436,N_12355);
nor U12677 (N_12677,N_12301,N_12273);
nor U12678 (N_12678,N_12457,N_12267);
xnor U12679 (N_12679,N_12156,N_12149);
or U12680 (N_12680,N_12364,N_12468);
and U12681 (N_12681,N_12442,N_12125);
or U12682 (N_12682,N_12428,N_12473);
xor U12683 (N_12683,N_12255,N_12057);
nand U12684 (N_12684,N_12451,N_12029);
nor U12685 (N_12685,N_12163,N_12415);
or U12686 (N_12686,N_12367,N_12427);
nor U12687 (N_12687,N_12483,N_12208);
nand U12688 (N_12688,N_12443,N_12186);
nand U12689 (N_12689,N_12305,N_12115);
nand U12690 (N_12690,N_12049,N_12371);
nand U12691 (N_12691,N_12387,N_12153);
nand U12692 (N_12692,N_12365,N_12398);
xor U12693 (N_12693,N_12463,N_12086);
and U12694 (N_12694,N_12229,N_12308);
nor U12695 (N_12695,N_12124,N_12134);
nor U12696 (N_12696,N_12102,N_12285);
nand U12697 (N_12697,N_12200,N_12204);
nand U12698 (N_12698,N_12019,N_12348);
nor U12699 (N_12699,N_12067,N_12061);
or U12700 (N_12700,N_12022,N_12137);
nor U12701 (N_12701,N_12117,N_12024);
xnor U12702 (N_12702,N_12380,N_12151);
or U12703 (N_12703,N_12317,N_12161);
xor U12704 (N_12704,N_12069,N_12075);
and U12705 (N_12705,N_12205,N_12472);
and U12706 (N_12706,N_12173,N_12394);
and U12707 (N_12707,N_12042,N_12469);
or U12708 (N_12708,N_12116,N_12287);
or U12709 (N_12709,N_12321,N_12298);
nor U12710 (N_12710,N_12250,N_12150);
nand U12711 (N_12711,N_12268,N_12051);
nor U12712 (N_12712,N_12127,N_12296);
nor U12713 (N_12713,N_12113,N_12236);
or U12714 (N_12714,N_12423,N_12275);
nor U12715 (N_12715,N_12262,N_12183);
xor U12716 (N_12716,N_12417,N_12203);
or U12717 (N_12717,N_12202,N_12390);
or U12718 (N_12718,N_12358,N_12011);
and U12719 (N_12719,N_12231,N_12104);
or U12720 (N_12720,N_12258,N_12288);
and U12721 (N_12721,N_12346,N_12008);
xor U12722 (N_12722,N_12100,N_12166);
or U12723 (N_12723,N_12425,N_12088);
or U12724 (N_12724,N_12187,N_12274);
and U12725 (N_12725,N_12397,N_12135);
or U12726 (N_12726,N_12141,N_12174);
nor U12727 (N_12727,N_12360,N_12339);
and U12728 (N_12728,N_12097,N_12479);
or U12729 (N_12729,N_12041,N_12414);
or U12730 (N_12730,N_12070,N_12277);
nor U12731 (N_12731,N_12114,N_12002);
and U12732 (N_12732,N_12283,N_12396);
and U12733 (N_12733,N_12312,N_12157);
nor U12734 (N_12734,N_12093,N_12370);
xnor U12735 (N_12735,N_12018,N_12381);
and U12736 (N_12736,N_12244,N_12431);
or U12737 (N_12737,N_12218,N_12021);
nand U12738 (N_12738,N_12215,N_12217);
nand U12739 (N_12739,N_12232,N_12162);
or U12740 (N_12740,N_12233,N_12025);
or U12741 (N_12741,N_12352,N_12477);
nor U12742 (N_12742,N_12432,N_12278);
nand U12743 (N_12743,N_12225,N_12334);
nand U12744 (N_12744,N_12142,N_12384);
nand U12745 (N_12745,N_12242,N_12272);
xnor U12746 (N_12746,N_12026,N_12052);
or U12747 (N_12747,N_12330,N_12410);
nor U12748 (N_12748,N_12392,N_12282);
nor U12749 (N_12749,N_12073,N_12491);
or U12750 (N_12750,N_12379,N_12477);
and U12751 (N_12751,N_12480,N_12499);
and U12752 (N_12752,N_12123,N_12059);
or U12753 (N_12753,N_12309,N_12411);
nor U12754 (N_12754,N_12315,N_12164);
and U12755 (N_12755,N_12073,N_12153);
and U12756 (N_12756,N_12154,N_12309);
and U12757 (N_12757,N_12233,N_12217);
or U12758 (N_12758,N_12069,N_12338);
or U12759 (N_12759,N_12240,N_12129);
and U12760 (N_12760,N_12412,N_12133);
and U12761 (N_12761,N_12017,N_12470);
nor U12762 (N_12762,N_12088,N_12456);
and U12763 (N_12763,N_12330,N_12023);
nor U12764 (N_12764,N_12011,N_12095);
nor U12765 (N_12765,N_12473,N_12419);
or U12766 (N_12766,N_12320,N_12025);
xnor U12767 (N_12767,N_12380,N_12214);
and U12768 (N_12768,N_12194,N_12306);
nor U12769 (N_12769,N_12173,N_12459);
nor U12770 (N_12770,N_12202,N_12083);
and U12771 (N_12771,N_12133,N_12333);
and U12772 (N_12772,N_12284,N_12269);
nor U12773 (N_12773,N_12246,N_12458);
or U12774 (N_12774,N_12260,N_12499);
or U12775 (N_12775,N_12408,N_12224);
nand U12776 (N_12776,N_12358,N_12246);
nor U12777 (N_12777,N_12311,N_12033);
xor U12778 (N_12778,N_12238,N_12010);
nand U12779 (N_12779,N_12323,N_12208);
nand U12780 (N_12780,N_12337,N_12288);
nand U12781 (N_12781,N_12365,N_12178);
xor U12782 (N_12782,N_12426,N_12313);
nand U12783 (N_12783,N_12156,N_12125);
xnor U12784 (N_12784,N_12304,N_12094);
nand U12785 (N_12785,N_12478,N_12357);
nor U12786 (N_12786,N_12362,N_12404);
or U12787 (N_12787,N_12089,N_12116);
or U12788 (N_12788,N_12475,N_12450);
or U12789 (N_12789,N_12453,N_12483);
nand U12790 (N_12790,N_12106,N_12071);
or U12791 (N_12791,N_12386,N_12382);
nor U12792 (N_12792,N_12119,N_12195);
xnor U12793 (N_12793,N_12030,N_12073);
and U12794 (N_12794,N_12461,N_12412);
xor U12795 (N_12795,N_12015,N_12017);
and U12796 (N_12796,N_12136,N_12383);
or U12797 (N_12797,N_12086,N_12362);
nor U12798 (N_12798,N_12361,N_12226);
nor U12799 (N_12799,N_12441,N_12083);
nand U12800 (N_12800,N_12123,N_12319);
or U12801 (N_12801,N_12335,N_12442);
nand U12802 (N_12802,N_12205,N_12338);
nor U12803 (N_12803,N_12272,N_12414);
and U12804 (N_12804,N_12334,N_12006);
or U12805 (N_12805,N_12405,N_12466);
or U12806 (N_12806,N_12139,N_12033);
or U12807 (N_12807,N_12088,N_12295);
and U12808 (N_12808,N_12493,N_12355);
nand U12809 (N_12809,N_12167,N_12403);
nor U12810 (N_12810,N_12109,N_12269);
nand U12811 (N_12811,N_12368,N_12327);
nor U12812 (N_12812,N_12290,N_12177);
and U12813 (N_12813,N_12261,N_12441);
and U12814 (N_12814,N_12128,N_12355);
and U12815 (N_12815,N_12131,N_12225);
nand U12816 (N_12816,N_12487,N_12496);
nor U12817 (N_12817,N_12123,N_12142);
and U12818 (N_12818,N_12037,N_12269);
xor U12819 (N_12819,N_12152,N_12424);
xor U12820 (N_12820,N_12352,N_12343);
or U12821 (N_12821,N_12356,N_12322);
nor U12822 (N_12822,N_12253,N_12099);
or U12823 (N_12823,N_12362,N_12117);
nand U12824 (N_12824,N_12382,N_12414);
nand U12825 (N_12825,N_12042,N_12346);
nand U12826 (N_12826,N_12251,N_12361);
nand U12827 (N_12827,N_12377,N_12498);
and U12828 (N_12828,N_12198,N_12033);
nor U12829 (N_12829,N_12383,N_12373);
xor U12830 (N_12830,N_12181,N_12492);
nand U12831 (N_12831,N_12477,N_12265);
nand U12832 (N_12832,N_12018,N_12356);
and U12833 (N_12833,N_12339,N_12359);
and U12834 (N_12834,N_12398,N_12364);
or U12835 (N_12835,N_12476,N_12015);
xor U12836 (N_12836,N_12113,N_12440);
nor U12837 (N_12837,N_12044,N_12172);
and U12838 (N_12838,N_12024,N_12381);
xor U12839 (N_12839,N_12369,N_12294);
and U12840 (N_12840,N_12416,N_12286);
or U12841 (N_12841,N_12492,N_12116);
nand U12842 (N_12842,N_12175,N_12269);
xnor U12843 (N_12843,N_12128,N_12007);
or U12844 (N_12844,N_12128,N_12040);
nor U12845 (N_12845,N_12233,N_12110);
and U12846 (N_12846,N_12145,N_12392);
nand U12847 (N_12847,N_12373,N_12194);
nand U12848 (N_12848,N_12286,N_12100);
xor U12849 (N_12849,N_12335,N_12200);
xnor U12850 (N_12850,N_12497,N_12462);
or U12851 (N_12851,N_12253,N_12194);
nor U12852 (N_12852,N_12363,N_12181);
nand U12853 (N_12853,N_12074,N_12417);
xor U12854 (N_12854,N_12400,N_12485);
nand U12855 (N_12855,N_12347,N_12447);
xnor U12856 (N_12856,N_12003,N_12121);
or U12857 (N_12857,N_12334,N_12210);
nand U12858 (N_12858,N_12073,N_12139);
or U12859 (N_12859,N_12040,N_12021);
xor U12860 (N_12860,N_12073,N_12181);
xor U12861 (N_12861,N_12195,N_12311);
nand U12862 (N_12862,N_12004,N_12460);
or U12863 (N_12863,N_12272,N_12326);
or U12864 (N_12864,N_12009,N_12410);
nand U12865 (N_12865,N_12343,N_12430);
nand U12866 (N_12866,N_12104,N_12004);
xnor U12867 (N_12867,N_12207,N_12131);
or U12868 (N_12868,N_12322,N_12234);
or U12869 (N_12869,N_12282,N_12360);
or U12870 (N_12870,N_12168,N_12156);
nor U12871 (N_12871,N_12488,N_12026);
nand U12872 (N_12872,N_12353,N_12423);
and U12873 (N_12873,N_12244,N_12360);
nand U12874 (N_12874,N_12074,N_12123);
nand U12875 (N_12875,N_12355,N_12380);
and U12876 (N_12876,N_12440,N_12142);
nand U12877 (N_12877,N_12003,N_12336);
and U12878 (N_12878,N_12467,N_12229);
nand U12879 (N_12879,N_12283,N_12243);
nor U12880 (N_12880,N_12065,N_12354);
and U12881 (N_12881,N_12429,N_12057);
nor U12882 (N_12882,N_12196,N_12302);
nand U12883 (N_12883,N_12295,N_12102);
xnor U12884 (N_12884,N_12213,N_12228);
nor U12885 (N_12885,N_12109,N_12038);
nand U12886 (N_12886,N_12130,N_12366);
or U12887 (N_12887,N_12017,N_12433);
xor U12888 (N_12888,N_12326,N_12198);
nor U12889 (N_12889,N_12479,N_12319);
nor U12890 (N_12890,N_12396,N_12134);
nor U12891 (N_12891,N_12413,N_12326);
xor U12892 (N_12892,N_12292,N_12007);
or U12893 (N_12893,N_12133,N_12137);
nand U12894 (N_12894,N_12392,N_12180);
or U12895 (N_12895,N_12037,N_12302);
nor U12896 (N_12896,N_12061,N_12114);
nor U12897 (N_12897,N_12173,N_12029);
xor U12898 (N_12898,N_12257,N_12298);
nor U12899 (N_12899,N_12080,N_12022);
nor U12900 (N_12900,N_12306,N_12496);
and U12901 (N_12901,N_12147,N_12366);
xor U12902 (N_12902,N_12165,N_12144);
nand U12903 (N_12903,N_12133,N_12418);
and U12904 (N_12904,N_12026,N_12214);
nand U12905 (N_12905,N_12043,N_12088);
nand U12906 (N_12906,N_12112,N_12138);
or U12907 (N_12907,N_12263,N_12122);
nand U12908 (N_12908,N_12359,N_12326);
or U12909 (N_12909,N_12295,N_12127);
and U12910 (N_12910,N_12450,N_12254);
or U12911 (N_12911,N_12469,N_12316);
and U12912 (N_12912,N_12459,N_12394);
nor U12913 (N_12913,N_12437,N_12194);
xor U12914 (N_12914,N_12022,N_12498);
and U12915 (N_12915,N_12397,N_12443);
and U12916 (N_12916,N_12390,N_12357);
nand U12917 (N_12917,N_12096,N_12386);
nand U12918 (N_12918,N_12068,N_12418);
nand U12919 (N_12919,N_12327,N_12333);
or U12920 (N_12920,N_12441,N_12067);
nand U12921 (N_12921,N_12078,N_12155);
and U12922 (N_12922,N_12256,N_12020);
or U12923 (N_12923,N_12066,N_12077);
or U12924 (N_12924,N_12122,N_12034);
nor U12925 (N_12925,N_12002,N_12368);
or U12926 (N_12926,N_12424,N_12012);
or U12927 (N_12927,N_12118,N_12238);
and U12928 (N_12928,N_12488,N_12200);
nand U12929 (N_12929,N_12183,N_12419);
nor U12930 (N_12930,N_12307,N_12280);
or U12931 (N_12931,N_12369,N_12494);
xor U12932 (N_12932,N_12141,N_12203);
nor U12933 (N_12933,N_12413,N_12021);
and U12934 (N_12934,N_12385,N_12367);
nand U12935 (N_12935,N_12059,N_12420);
and U12936 (N_12936,N_12392,N_12172);
nor U12937 (N_12937,N_12098,N_12384);
nor U12938 (N_12938,N_12057,N_12161);
xnor U12939 (N_12939,N_12140,N_12268);
xor U12940 (N_12940,N_12088,N_12040);
and U12941 (N_12941,N_12458,N_12042);
nand U12942 (N_12942,N_12486,N_12496);
nor U12943 (N_12943,N_12077,N_12279);
and U12944 (N_12944,N_12310,N_12472);
and U12945 (N_12945,N_12025,N_12309);
and U12946 (N_12946,N_12076,N_12077);
nand U12947 (N_12947,N_12273,N_12453);
or U12948 (N_12948,N_12314,N_12171);
nor U12949 (N_12949,N_12121,N_12056);
nand U12950 (N_12950,N_12013,N_12188);
or U12951 (N_12951,N_12172,N_12272);
nor U12952 (N_12952,N_12389,N_12369);
nor U12953 (N_12953,N_12023,N_12047);
nor U12954 (N_12954,N_12113,N_12230);
xor U12955 (N_12955,N_12307,N_12180);
xor U12956 (N_12956,N_12260,N_12312);
nand U12957 (N_12957,N_12221,N_12043);
nand U12958 (N_12958,N_12061,N_12245);
nand U12959 (N_12959,N_12132,N_12355);
and U12960 (N_12960,N_12207,N_12398);
xnor U12961 (N_12961,N_12274,N_12067);
nor U12962 (N_12962,N_12229,N_12498);
or U12963 (N_12963,N_12459,N_12093);
nand U12964 (N_12964,N_12346,N_12307);
nor U12965 (N_12965,N_12414,N_12265);
or U12966 (N_12966,N_12095,N_12165);
or U12967 (N_12967,N_12134,N_12034);
nor U12968 (N_12968,N_12183,N_12460);
xnor U12969 (N_12969,N_12097,N_12328);
nor U12970 (N_12970,N_12464,N_12278);
nor U12971 (N_12971,N_12109,N_12382);
or U12972 (N_12972,N_12276,N_12039);
or U12973 (N_12973,N_12071,N_12385);
nand U12974 (N_12974,N_12318,N_12321);
nor U12975 (N_12975,N_12280,N_12268);
or U12976 (N_12976,N_12338,N_12030);
nor U12977 (N_12977,N_12354,N_12409);
or U12978 (N_12978,N_12321,N_12126);
or U12979 (N_12979,N_12056,N_12254);
and U12980 (N_12980,N_12265,N_12245);
xor U12981 (N_12981,N_12391,N_12011);
and U12982 (N_12982,N_12412,N_12376);
and U12983 (N_12983,N_12375,N_12019);
nor U12984 (N_12984,N_12359,N_12018);
nor U12985 (N_12985,N_12198,N_12242);
xor U12986 (N_12986,N_12203,N_12028);
xnor U12987 (N_12987,N_12233,N_12484);
and U12988 (N_12988,N_12313,N_12184);
or U12989 (N_12989,N_12404,N_12047);
nor U12990 (N_12990,N_12420,N_12409);
nor U12991 (N_12991,N_12191,N_12150);
or U12992 (N_12992,N_12327,N_12244);
or U12993 (N_12993,N_12351,N_12272);
and U12994 (N_12994,N_12044,N_12188);
nand U12995 (N_12995,N_12115,N_12333);
and U12996 (N_12996,N_12445,N_12329);
xnor U12997 (N_12997,N_12292,N_12433);
nand U12998 (N_12998,N_12081,N_12093);
nor U12999 (N_12999,N_12118,N_12251);
nand U13000 (N_13000,N_12712,N_12845);
or U13001 (N_13001,N_12838,N_12740);
nand U13002 (N_13002,N_12746,N_12965);
and U13003 (N_13003,N_12928,N_12634);
xnor U13004 (N_13004,N_12792,N_12807);
nand U13005 (N_13005,N_12821,N_12692);
and U13006 (N_13006,N_12733,N_12527);
nor U13007 (N_13007,N_12888,N_12585);
xor U13008 (N_13008,N_12829,N_12875);
or U13009 (N_13009,N_12649,N_12864);
or U13010 (N_13010,N_12988,N_12884);
and U13011 (N_13011,N_12617,N_12764);
nand U13012 (N_13012,N_12759,N_12936);
nand U13013 (N_13013,N_12950,N_12781);
nand U13014 (N_13014,N_12700,N_12620);
nand U13015 (N_13015,N_12701,N_12938);
nor U13016 (N_13016,N_12597,N_12921);
and U13017 (N_13017,N_12693,N_12686);
nor U13018 (N_13018,N_12559,N_12826);
nand U13019 (N_13019,N_12580,N_12849);
or U13020 (N_13020,N_12713,N_12677);
nor U13021 (N_13021,N_12635,N_12531);
or U13022 (N_13022,N_12916,N_12793);
nor U13023 (N_13023,N_12776,N_12905);
nor U13024 (N_13024,N_12751,N_12828);
nor U13025 (N_13025,N_12874,N_12524);
xnor U13026 (N_13026,N_12579,N_12754);
xor U13027 (N_13027,N_12638,N_12632);
or U13028 (N_13028,N_12548,N_12689);
or U13029 (N_13029,N_12798,N_12955);
or U13030 (N_13030,N_12629,N_12702);
nand U13031 (N_13031,N_12900,N_12815);
and U13032 (N_13032,N_12510,N_12668);
and U13033 (N_13033,N_12744,N_12783);
nand U13034 (N_13034,N_12523,N_12813);
or U13035 (N_13035,N_12671,N_12878);
nor U13036 (N_13036,N_12571,N_12515);
and U13037 (N_13037,N_12736,N_12806);
xnor U13038 (N_13038,N_12802,N_12964);
or U13039 (N_13039,N_12596,N_12985);
and U13040 (N_13040,N_12763,N_12765);
or U13041 (N_13041,N_12663,N_12768);
or U13042 (N_13042,N_12573,N_12881);
nor U13043 (N_13043,N_12778,N_12914);
and U13044 (N_13044,N_12834,N_12711);
nand U13045 (N_13045,N_12581,N_12823);
and U13046 (N_13046,N_12831,N_12636);
xor U13047 (N_13047,N_12511,N_12972);
nor U13048 (N_13048,N_12658,N_12787);
nor U13049 (N_13049,N_12930,N_12760);
nor U13050 (N_13050,N_12984,N_12614);
nand U13051 (N_13051,N_12625,N_12912);
nor U13052 (N_13052,N_12980,N_12879);
or U13053 (N_13053,N_12859,N_12537);
nand U13054 (N_13054,N_12642,N_12611);
and U13055 (N_13055,N_12534,N_12922);
xnor U13056 (N_13056,N_12791,N_12684);
xor U13057 (N_13057,N_12532,N_12851);
or U13058 (N_13058,N_12767,N_12973);
and U13059 (N_13059,N_12974,N_12971);
and U13060 (N_13060,N_12761,N_12946);
or U13061 (N_13061,N_12664,N_12825);
and U13062 (N_13062,N_12999,N_12691);
nor U13063 (N_13063,N_12709,N_12948);
or U13064 (N_13064,N_12725,N_12758);
and U13065 (N_13065,N_12683,N_12687);
nand U13066 (N_13066,N_12832,N_12707);
or U13067 (N_13067,N_12512,N_12956);
nor U13068 (N_13068,N_12503,N_12925);
or U13069 (N_13069,N_12616,N_12899);
nor U13070 (N_13070,N_12720,N_12766);
nand U13071 (N_13071,N_12848,N_12833);
nand U13072 (N_13072,N_12739,N_12587);
and U13073 (N_13073,N_12817,N_12883);
xnor U13074 (N_13074,N_12660,N_12530);
and U13075 (N_13075,N_12522,N_12835);
or U13076 (N_13076,N_12882,N_12591);
and U13077 (N_13077,N_12565,N_12749);
nand U13078 (N_13078,N_12622,N_12504);
nor U13079 (N_13079,N_12673,N_12771);
and U13080 (N_13080,N_12836,N_12646);
or U13081 (N_13081,N_12743,N_12890);
xnor U13082 (N_13082,N_12852,N_12871);
xnor U13083 (N_13083,N_12672,N_12880);
xnor U13084 (N_13084,N_12977,N_12841);
xnor U13085 (N_13085,N_12641,N_12872);
and U13086 (N_13086,N_12857,N_12556);
or U13087 (N_13087,N_12870,N_12607);
xor U13088 (N_13088,N_12590,N_12752);
nand U13089 (N_13089,N_12699,N_12891);
or U13090 (N_13090,N_12583,N_12514);
xnor U13091 (N_13091,N_12619,N_12794);
xnor U13092 (N_13092,N_12982,N_12850);
nand U13093 (N_13093,N_12885,N_12628);
and U13094 (N_13094,N_12932,N_12595);
or U13095 (N_13095,N_12991,N_12724);
nand U13096 (N_13096,N_12703,N_12732);
xnor U13097 (N_13097,N_12970,N_12969);
and U13098 (N_13098,N_12987,N_12947);
nor U13099 (N_13099,N_12500,N_12708);
and U13100 (N_13100,N_12533,N_12582);
and U13101 (N_13101,N_12839,N_12558);
nor U13102 (N_13102,N_12561,N_12650);
nand U13103 (N_13103,N_12519,N_12951);
and U13104 (N_13104,N_12697,N_12727);
or U13105 (N_13105,N_12570,N_12669);
or U13106 (N_13106,N_12804,N_12613);
xnor U13107 (N_13107,N_12989,N_12958);
xnor U13108 (N_13108,N_12680,N_12704);
nand U13109 (N_13109,N_12808,N_12506);
or U13110 (N_13110,N_12923,N_12997);
and U13111 (N_13111,N_12550,N_12645);
or U13112 (N_13112,N_12960,N_12602);
xnor U13113 (N_13113,N_12934,N_12608);
nand U13114 (N_13114,N_12953,N_12795);
xnor U13115 (N_13115,N_12893,N_12529);
or U13116 (N_13116,N_12865,N_12862);
or U13117 (N_13117,N_12690,N_12695);
and U13118 (N_13118,N_12762,N_12861);
xnor U13119 (N_13119,N_12846,N_12931);
xnor U13120 (N_13120,N_12566,N_12601);
nor U13121 (N_13121,N_12623,N_12705);
nand U13122 (N_13122,N_12741,N_12779);
nor U13123 (N_13123,N_12904,N_12654);
or U13124 (N_13124,N_12979,N_12735);
nor U13125 (N_13125,N_12726,N_12651);
and U13126 (N_13126,N_12995,N_12722);
nor U13127 (N_13127,N_12803,N_12992);
nor U13128 (N_13128,N_12978,N_12674);
xor U13129 (N_13129,N_12535,N_12889);
xor U13130 (N_13130,N_12860,N_12858);
nor U13131 (N_13131,N_12678,N_12539);
nand U13132 (N_13132,N_12661,N_12929);
nand U13133 (N_13133,N_12941,N_12715);
nor U13134 (N_13134,N_12513,N_12944);
or U13135 (N_13135,N_12568,N_12844);
nand U13136 (N_13136,N_12667,N_12589);
or U13137 (N_13137,N_12756,N_12775);
or U13138 (N_13138,N_12818,N_12785);
or U13139 (N_13139,N_12847,N_12631);
nor U13140 (N_13140,N_12981,N_12721);
or U13141 (N_13141,N_12837,N_12706);
nor U13142 (N_13142,N_12910,N_12896);
xor U13143 (N_13143,N_12755,N_12949);
xor U13144 (N_13144,N_12868,N_12569);
and U13145 (N_13145,N_12509,N_12894);
and U13146 (N_13146,N_12966,N_12586);
or U13147 (N_13147,N_12546,N_12560);
xnor U13148 (N_13148,N_12547,N_12576);
and U13149 (N_13149,N_12536,N_12747);
nand U13150 (N_13150,N_12520,N_12901);
xor U13151 (N_13151,N_12854,N_12907);
nand U13152 (N_13152,N_12717,N_12564);
or U13153 (N_13153,N_12643,N_12924);
nand U13154 (N_13154,N_12935,N_12603);
xor U13155 (N_13155,N_12915,N_12920);
nor U13156 (N_13156,N_12688,N_12954);
xor U13157 (N_13157,N_12545,N_12830);
nand U13158 (N_13158,N_12679,N_12877);
nand U13159 (N_13159,N_12962,N_12790);
and U13160 (N_13160,N_12729,N_12942);
nor U13161 (N_13161,N_12819,N_12918);
and U13162 (N_13162,N_12867,N_12659);
and U13163 (N_13163,N_12876,N_12940);
or U13164 (N_13164,N_12553,N_12737);
xor U13165 (N_13165,N_12563,N_12774);
xor U13166 (N_13166,N_12959,N_12723);
nor U13167 (N_13167,N_12549,N_12592);
or U13168 (N_13168,N_12994,N_12639);
nor U13169 (N_13169,N_12567,N_12612);
xnor U13170 (N_13170,N_12917,N_12577);
nand U13171 (N_13171,N_12502,N_12856);
xor U13172 (N_13172,N_12627,N_12606);
and U13173 (N_13173,N_12873,N_12605);
and U13174 (N_13174,N_12618,N_12753);
and U13175 (N_13175,N_12796,N_12963);
nand U13176 (N_13176,N_12685,N_12913);
nor U13177 (N_13177,N_12968,N_12811);
xnor U13178 (N_13178,N_12898,N_12554);
or U13179 (N_13179,N_12887,N_12853);
and U13180 (N_13180,N_12983,N_12657);
nand U13181 (N_13181,N_12769,N_12810);
nand U13182 (N_13182,N_12572,N_12788);
xnor U13183 (N_13183,N_12653,N_12521);
nor U13184 (N_13184,N_12528,N_12770);
xor U13185 (N_13185,N_12748,N_12757);
and U13186 (N_13186,N_12593,N_12630);
nor U13187 (N_13187,N_12742,N_12895);
nand U13188 (N_13188,N_12939,N_12902);
xnor U13189 (N_13189,N_12906,N_12816);
xnor U13190 (N_13190,N_12805,N_12599);
nor U13191 (N_13191,N_12897,N_12662);
xnor U13192 (N_13192,N_12655,N_12682);
and U13193 (N_13193,N_12694,N_12782);
xor U13194 (N_13194,N_12797,N_12990);
or U13195 (N_13195,N_12640,N_12908);
nand U13196 (N_13196,N_12578,N_12967);
nand U13197 (N_13197,N_12926,N_12675);
xnor U13198 (N_13198,N_12996,N_12866);
nor U13199 (N_13199,N_12738,N_12945);
nor U13200 (N_13200,N_12540,N_12594);
and U13201 (N_13201,N_12716,N_12615);
nand U13202 (N_13202,N_12919,N_12508);
or U13203 (N_13203,N_12598,N_12665);
nor U13204 (N_13204,N_12562,N_12551);
nand U13205 (N_13205,N_12892,N_12525);
or U13206 (N_13206,N_12538,N_12526);
or U13207 (N_13207,N_12555,N_12886);
xnor U13208 (N_13208,N_12843,N_12750);
xnor U13209 (N_13209,N_12574,N_12719);
xor U13210 (N_13210,N_12855,N_12772);
nand U13211 (N_13211,N_12718,N_12840);
or U13212 (N_13212,N_12728,N_12780);
xor U13213 (N_13213,N_12952,N_12610);
nor U13214 (N_13214,N_12927,N_12600);
nor U13215 (N_13215,N_12501,N_12666);
nor U13216 (N_13216,N_12975,N_12903);
or U13217 (N_13217,N_12820,N_12909);
or U13218 (N_13218,N_12812,N_12517);
xnor U13219 (N_13219,N_12863,N_12809);
xor U13220 (N_13220,N_12507,N_12696);
or U13221 (N_13221,N_12842,N_12745);
nor U13222 (N_13222,N_12731,N_12609);
nor U13223 (N_13223,N_12799,N_12933);
nand U13224 (N_13224,N_12543,N_12575);
nand U13225 (N_13225,N_12698,N_12827);
xor U13226 (N_13226,N_12961,N_12800);
nand U13227 (N_13227,N_12786,N_12604);
and U13228 (N_13228,N_12644,N_12943);
nor U13229 (N_13229,N_12993,N_12814);
and U13230 (N_13230,N_12710,N_12777);
nor U13231 (N_13231,N_12621,N_12998);
xnor U13232 (N_13232,N_12541,N_12588);
nor U13233 (N_13233,N_12647,N_12584);
or U13234 (N_13234,N_12789,N_12957);
nor U13235 (N_13235,N_12516,N_12670);
nand U13236 (N_13236,N_12937,N_12652);
nor U13237 (N_13237,N_12542,N_12656);
nand U13238 (N_13238,N_12801,N_12626);
nor U13239 (N_13239,N_12633,N_12681);
and U13240 (N_13240,N_12557,N_12773);
or U13241 (N_13241,N_12784,N_12822);
and U13242 (N_13242,N_12676,N_12518);
nor U13243 (N_13243,N_12730,N_12714);
or U13244 (N_13244,N_12911,N_12734);
xnor U13245 (N_13245,N_12824,N_12976);
nor U13246 (N_13246,N_12552,N_12624);
nand U13247 (N_13247,N_12544,N_12505);
xor U13248 (N_13248,N_12648,N_12986);
and U13249 (N_13249,N_12869,N_12637);
xnor U13250 (N_13250,N_12836,N_12532);
nor U13251 (N_13251,N_12609,N_12878);
xnor U13252 (N_13252,N_12900,N_12950);
or U13253 (N_13253,N_12548,N_12522);
or U13254 (N_13254,N_12555,N_12615);
and U13255 (N_13255,N_12869,N_12612);
and U13256 (N_13256,N_12828,N_12524);
and U13257 (N_13257,N_12654,N_12781);
and U13258 (N_13258,N_12957,N_12603);
or U13259 (N_13259,N_12562,N_12586);
or U13260 (N_13260,N_12742,N_12991);
or U13261 (N_13261,N_12876,N_12617);
and U13262 (N_13262,N_12664,N_12986);
and U13263 (N_13263,N_12626,N_12973);
or U13264 (N_13264,N_12744,N_12647);
or U13265 (N_13265,N_12738,N_12737);
nand U13266 (N_13266,N_12570,N_12566);
and U13267 (N_13267,N_12646,N_12639);
nor U13268 (N_13268,N_12990,N_12779);
nand U13269 (N_13269,N_12576,N_12694);
xor U13270 (N_13270,N_12786,N_12689);
or U13271 (N_13271,N_12648,N_12695);
nand U13272 (N_13272,N_12671,N_12570);
and U13273 (N_13273,N_12950,N_12862);
xor U13274 (N_13274,N_12799,N_12677);
nor U13275 (N_13275,N_12591,N_12782);
nand U13276 (N_13276,N_12934,N_12694);
and U13277 (N_13277,N_12611,N_12721);
nor U13278 (N_13278,N_12572,N_12747);
xnor U13279 (N_13279,N_12974,N_12782);
xor U13280 (N_13280,N_12935,N_12580);
and U13281 (N_13281,N_12522,N_12814);
nor U13282 (N_13282,N_12925,N_12960);
and U13283 (N_13283,N_12808,N_12952);
nand U13284 (N_13284,N_12617,N_12699);
nand U13285 (N_13285,N_12909,N_12671);
xnor U13286 (N_13286,N_12660,N_12815);
and U13287 (N_13287,N_12756,N_12664);
nand U13288 (N_13288,N_12858,N_12854);
or U13289 (N_13289,N_12992,N_12590);
nand U13290 (N_13290,N_12651,N_12539);
or U13291 (N_13291,N_12801,N_12567);
and U13292 (N_13292,N_12565,N_12945);
nor U13293 (N_13293,N_12899,N_12959);
nand U13294 (N_13294,N_12549,N_12587);
and U13295 (N_13295,N_12830,N_12784);
nand U13296 (N_13296,N_12921,N_12804);
and U13297 (N_13297,N_12850,N_12633);
xnor U13298 (N_13298,N_12890,N_12967);
nand U13299 (N_13299,N_12652,N_12701);
and U13300 (N_13300,N_12771,N_12539);
nand U13301 (N_13301,N_12885,N_12814);
xnor U13302 (N_13302,N_12913,N_12863);
nand U13303 (N_13303,N_12757,N_12684);
nand U13304 (N_13304,N_12870,N_12894);
nand U13305 (N_13305,N_12866,N_12717);
or U13306 (N_13306,N_12693,N_12566);
or U13307 (N_13307,N_12816,N_12799);
nor U13308 (N_13308,N_12967,N_12826);
or U13309 (N_13309,N_12693,N_12527);
xnor U13310 (N_13310,N_12614,N_12715);
and U13311 (N_13311,N_12518,N_12531);
xnor U13312 (N_13312,N_12606,N_12741);
nand U13313 (N_13313,N_12660,N_12707);
nor U13314 (N_13314,N_12662,N_12660);
or U13315 (N_13315,N_12642,N_12889);
and U13316 (N_13316,N_12766,N_12618);
nor U13317 (N_13317,N_12683,N_12952);
xor U13318 (N_13318,N_12548,N_12554);
xnor U13319 (N_13319,N_12847,N_12979);
or U13320 (N_13320,N_12627,N_12636);
and U13321 (N_13321,N_12828,N_12968);
or U13322 (N_13322,N_12698,N_12552);
nand U13323 (N_13323,N_12841,N_12908);
or U13324 (N_13324,N_12989,N_12643);
and U13325 (N_13325,N_12770,N_12971);
nor U13326 (N_13326,N_12929,N_12951);
and U13327 (N_13327,N_12998,N_12992);
and U13328 (N_13328,N_12965,N_12995);
and U13329 (N_13329,N_12910,N_12936);
or U13330 (N_13330,N_12508,N_12505);
or U13331 (N_13331,N_12827,N_12962);
and U13332 (N_13332,N_12746,N_12562);
nand U13333 (N_13333,N_12659,N_12897);
or U13334 (N_13334,N_12818,N_12919);
xor U13335 (N_13335,N_12711,N_12841);
xnor U13336 (N_13336,N_12715,N_12875);
nor U13337 (N_13337,N_12889,N_12849);
nand U13338 (N_13338,N_12630,N_12589);
xor U13339 (N_13339,N_12726,N_12660);
xnor U13340 (N_13340,N_12779,N_12584);
nand U13341 (N_13341,N_12627,N_12571);
nand U13342 (N_13342,N_12796,N_12555);
and U13343 (N_13343,N_12506,N_12505);
or U13344 (N_13344,N_12758,N_12671);
nor U13345 (N_13345,N_12955,N_12921);
nor U13346 (N_13346,N_12615,N_12810);
xnor U13347 (N_13347,N_12783,N_12937);
nand U13348 (N_13348,N_12925,N_12624);
nor U13349 (N_13349,N_12960,N_12697);
and U13350 (N_13350,N_12793,N_12838);
nor U13351 (N_13351,N_12696,N_12625);
and U13352 (N_13352,N_12797,N_12964);
or U13353 (N_13353,N_12585,N_12913);
nand U13354 (N_13354,N_12921,N_12721);
nor U13355 (N_13355,N_12655,N_12741);
xor U13356 (N_13356,N_12711,N_12673);
nor U13357 (N_13357,N_12743,N_12530);
nor U13358 (N_13358,N_12907,N_12867);
nand U13359 (N_13359,N_12931,N_12758);
xnor U13360 (N_13360,N_12677,N_12501);
or U13361 (N_13361,N_12891,N_12965);
nor U13362 (N_13362,N_12851,N_12984);
or U13363 (N_13363,N_12792,N_12843);
xor U13364 (N_13364,N_12970,N_12706);
nand U13365 (N_13365,N_12533,N_12657);
nor U13366 (N_13366,N_12545,N_12804);
nand U13367 (N_13367,N_12964,N_12786);
nand U13368 (N_13368,N_12515,N_12974);
nand U13369 (N_13369,N_12829,N_12621);
or U13370 (N_13370,N_12775,N_12860);
xnor U13371 (N_13371,N_12757,N_12593);
and U13372 (N_13372,N_12581,N_12590);
or U13373 (N_13373,N_12513,N_12527);
nor U13374 (N_13374,N_12880,N_12651);
nand U13375 (N_13375,N_12841,N_12833);
nor U13376 (N_13376,N_12973,N_12826);
xor U13377 (N_13377,N_12518,N_12798);
nor U13378 (N_13378,N_12820,N_12896);
and U13379 (N_13379,N_12939,N_12959);
or U13380 (N_13380,N_12710,N_12731);
or U13381 (N_13381,N_12934,N_12782);
or U13382 (N_13382,N_12967,N_12982);
nor U13383 (N_13383,N_12701,N_12808);
xor U13384 (N_13384,N_12886,N_12645);
or U13385 (N_13385,N_12735,N_12789);
or U13386 (N_13386,N_12665,N_12670);
xor U13387 (N_13387,N_12844,N_12879);
nor U13388 (N_13388,N_12901,N_12919);
or U13389 (N_13389,N_12722,N_12508);
nand U13390 (N_13390,N_12514,N_12577);
nand U13391 (N_13391,N_12600,N_12663);
or U13392 (N_13392,N_12623,N_12812);
xnor U13393 (N_13393,N_12829,N_12631);
or U13394 (N_13394,N_12672,N_12596);
xor U13395 (N_13395,N_12957,N_12573);
or U13396 (N_13396,N_12652,N_12634);
and U13397 (N_13397,N_12597,N_12605);
and U13398 (N_13398,N_12542,N_12863);
xor U13399 (N_13399,N_12622,N_12885);
nand U13400 (N_13400,N_12859,N_12576);
or U13401 (N_13401,N_12556,N_12594);
nand U13402 (N_13402,N_12792,N_12743);
or U13403 (N_13403,N_12617,N_12615);
xor U13404 (N_13404,N_12815,N_12735);
and U13405 (N_13405,N_12745,N_12541);
or U13406 (N_13406,N_12701,N_12871);
nand U13407 (N_13407,N_12650,N_12838);
xor U13408 (N_13408,N_12780,N_12501);
nand U13409 (N_13409,N_12529,N_12936);
nand U13410 (N_13410,N_12975,N_12844);
nand U13411 (N_13411,N_12705,N_12562);
nand U13412 (N_13412,N_12541,N_12908);
and U13413 (N_13413,N_12857,N_12587);
xor U13414 (N_13414,N_12531,N_12915);
and U13415 (N_13415,N_12754,N_12573);
nor U13416 (N_13416,N_12765,N_12565);
nor U13417 (N_13417,N_12522,N_12945);
xnor U13418 (N_13418,N_12604,N_12506);
xor U13419 (N_13419,N_12828,N_12675);
nor U13420 (N_13420,N_12635,N_12827);
xor U13421 (N_13421,N_12979,N_12696);
or U13422 (N_13422,N_12562,N_12736);
xor U13423 (N_13423,N_12629,N_12911);
xor U13424 (N_13424,N_12867,N_12608);
xor U13425 (N_13425,N_12666,N_12726);
and U13426 (N_13426,N_12650,N_12940);
nand U13427 (N_13427,N_12957,N_12566);
nor U13428 (N_13428,N_12996,N_12917);
nor U13429 (N_13429,N_12630,N_12742);
and U13430 (N_13430,N_12571,N_12808);
nand U13431 (N_13431,N_12542,N_12759);
xor U13432 (N_13432,N_12861,N_12986);
nand U13433 (N_13433,N_12666,N_12515);
nand U13434 (N_13434,N_12572,N_12771);
xor U13435 (N_13435,N_12923,N_12628);
xor U13436 (N_13436,N_12839,N_12761);
xor U13437 (N_13437,N_12933,N_12677);
xor U13438 (N_13438,N_12521,N_12510);
and U13439 (N_13439,N_12875,N_12601);
nor U13440 (N_13440,N_12754,N_12768);
nor U13441 (N_13441,N_12592,N_12614);
or U13442 (N_13442,N_12823,N_12679);
nand U13443 (N_13443,N_12655,N_12561);
xor U13444 (N_13444,N_12969,N_12727);
or U13445 (N_13445,N_12681,N_12924);
nand U13446 (N_13446,N_12831,N_12646);
xnor U13447 (N_13447,N_12683,N_12847);
and U13448 (N_13448,N_12774,N_12646);
xnor U13449 (N_13449,N_12797,N_12657);
and U13450 (N_13450,N_12502,N_12826);
and U13451 (N_13451,N_12572,N_12879);
nand U13452 (N_13452,N_12952,N_12964);
nand U13453 (N_13453,N_12591,N_12905);
xnor U13454 (N_13454,N_12857,N_12733);
nor U13455 (N_13455,N_12725,N_12730);
nor U13456 (N_13456,N_12584,N_12578);
xnor U13457 (N_13457,N_12540,N_12995);
and U13458 (N_13458,N_12522,N_12785);
nor U13459 (N_13459,N_12763,N_12564);
and U13460 (N_13460,N_12975,N_12912);
xnor U13461 (N_13461,N_12896,N_12518);
nand U13462 (N_13462,N_12679,N_12573);
xnor U13463 (N_13463,N_12777,N_12697);
nand U13464 (N_13464,N_12770,N_12621);
and U13465 (N_13465,N_12888,N_12881);
nor U13466 (N_13466,N_12712,N_12763);
or U13467 (N_13467,N_12728,N_12613);
xor U13468 (N_13468,N_12854,N_12544);
nor U13469 (N_13469,N_12737,N_12976);
nor U13470 (N_13470,N_12537,N_12959);
and U13471 (N_13471,N_12624,N_12537);
and U13472 (N_13472,N_12885,N_12587);
xnor U13473 (N_13473,N_12843,N_12747);
nand U13474 (N_13474,N_12915,N_12652);
or U13475 (N_13475,N_12841,N_12891);
nand U13476 (N_13476,N_12565,N_12580);
xor U13477 (N_13477,N_12864,N_12563);
and U13478 (N_13478,N_12912,N_12521);
nor U13479 (N_13479,N_12502,N_12844);
nor U13480 (N_13480,N_12831,N_12523);
and U13481 (N_13481,N_12950,N_12563);
and U13482 (N_13482,N_12900,N_12678);
nor U13483 (N_13483,N_12790,N_12564);
nand U13484 (N_13484,N_12553,N_12889);
or U13485 (N_13485,N_12889,N_12940);
and U13486 (N_13486,N_12777,N_12663);
nand U13487 (N_13487,N_12607,N_12939);
nand U13488 (N_13488,N_12928,N_12515);
nand U13489 (N_13489,N_12648,N_12951);
and U13490 (N_13490,N_12934,N_12847);
or U13491 (N_13491,N_12521,N_12899);
and U13492 (N_13492,N_12933,N_12731);
or U13493 (N_13493,N_12623,N_12999);
nand U13494 (N_13494,N_12658,N_12841);
and U13495 (N_13495,N_12762,N_12541);
xor U13496 (N_13496,N_12724,N_12539);
xor U13497 (N_13497,N_12515,N_12872);
and U13498 (N_13498,N_12626,N_12685);
nor U13499 (N_13499,N_12641,N_12777);
xor U13500 (N_13500,N_13481,N_13200);
and U13501 (N_13501,N_13070,N_13193);
xor U13502 (N_13502,N_13378,N_13090);
xor U13503 (N_13503,N_13368,N_13071);
and U13504 (N_13504,N_13337,N_13287);
nand U13505 (N_13505,N_13115,N_13398);
or U13506 (N_13506,N_13322,N_13492);
nor U13507 (N_13507,N_13136,N_13401);
or U13508 (N_13508,N_13180,N_13421);
nand U13509 (N_13509,N_13412,N_13268);
nand U13510 (N_13510,N_13402,N_13498);
nor U13511 (N_13511,N_13374,N_13280);
xor U13512 (N_13512,N_13106,N_13484);
nand U13513 (N_13513,N_13038,N_13244);
nor U13514 (N_13514,N_13255,N_13356);
nor U13515 (N_13515,N_13009,N_13300);
xnor U13516 (N_13516,N_13447,N_13393);
and U13517 (N_13517,N_13286,N_13445);
xnor U13518 (N_13518,N_13351,N_13105);
and U13519 (N_13519,N_13364,N_13143);
nand U13520 (N_13520,N_13146,N_13175);
or U13521 (N_13521,N_13452,N_13489);
and U13522 (N_13522,N_13097,N_13359);
or U13523 (N_13523,N_13462,N_13113);
and U13524 (N_13524,N_13050,N_13111);
nor U13525 (N_13525,N_13279,N_13026);
nand U13526 (N_13526,N_13198,N_13248);
or U13527 (N_13527,N_13389,N_13024);
or U13528 (N_13528,N_13446,N_13100);
xor U13529 (N_13529,N_13063,N_13144);
nor U13530 (N_13530,N_13301,N_13228);
nand U13531 (N_13531,N_13034,N_13207);
and U13532 (N_13532,N_13323,N_13273);
nor U13533 (N_13533,N_13027,N_13473);
and U13534 (N_13534,N_13283,N_13068);
nor U13535 (N_13535,N_13182,N_13429);
xnor U13536 (N_13536,N_13139,N_13159);
nor U13537 (N_13537,N_13056,N_13456);
xnor U13538 (N_13538,N_13078,N_13002);
nor U13539 (N_13539,N_13480,N_13367);
nor U13540 (N_13540,N_13474,N_13414);
xor U13541 (N_13541,N_13477,N_13203);
nor U13542 (N_13542,N_13016,N_13174);
nand U13543 (N_13543,N_13006,N_13208);
and U13544 (N_13544,N_13055,N_13032);
nand U13545 (N_13545,N_13297,N_13176);
or U13546 (N_13546,N_13017,N_13008);
nor U13547 (N_13547,N_13204,N_13443);
and U13548 (N_13548,N_13127,N_13355);
or U13549 (N_13549,N_13237,N_13256);
nand U13550 (N_13550,N_13296,N_13419);
nor U13551 (N_13551,N_13339,N_13298);
or U13552 (N_13552,N_13222,N_13425);
or U13553 (N_13553,N_13365,N_13250);
nand U13554 (N_13554,N_13338,N_13463);
nand U13555 (N_13555,N_13307,N_13453);
xor U13556 (N_13556,N_13080,N_13395);
or U13557 (N_13557,N_13199,N_13345);
or U13558 (N_13558,N_13158,N_13011);
nor U13559 (N_13559,N_13376,N_13360);
nand U13560 (N_13560,N_13232,N_13444);
and U13561 (N_13561,N_13242,N_13420);
nand U13562 (N_13562,N_13224,N_13133);
and U13563 (N_13563,N_13013,N_13385);
nand U13564 (N_13564,N_13109,N_13427);
nand U13565 (N_13565,N_13277,N_13004);
xor U13566 (N_13566,N_13449,N_13392);
nor U13567 (N_13567,N_13119,N_13142);
or U13568 (N_13568,N_13195,N_13214);
nand U13569 (N_13569,N_13494,N_13418);
nand U13570 (N_13570,N_13332,N_13226);
nand U13571 (N_13571,N_13346,N_13290);
xor U13572 (N_13572,N_13470,N_13375);
and U13573 (N_13573,N_13076,N_13309);
xor U13574 (N_13574,N_13285,N_13328);
or U13575 (N_13575,N_13305,N_13439);
and U13576 (N_13576,N_13157,N_13028);
and U13577 (N_13577,N_13344,N_13329);
or U13578 (N_13578,N_13137,N_13448);
nor U13579 (N_13579,N_13249,N_13259);
nand U13580 (N_13580,N_13052,N_13276);
and U13581 (N_13581,N_13441,N_13134);
xor U13582 (N_13582,N_13320,N_13123);
nand U13583 (N_13583,N_13014,N_13460);
xnor U13584 (N_13584,N_13152,N_13394);
xor U13585 (N_13585,N_13049,N_13030);
and U13586 (N_13586,N_13035,N_13251);
nor U13587 (N_13587,N_13170,N_13019);
nand U13588 (N_13588,N_13253,N_13150);
or U13589 (N_13589,N_13431,N_13424);
nand U13590 (N_13590,N_13223,N_13302);
nor U13591 (N_13591,N_13354,N_13162);
nor U13592 (N_13592,N_13262,N_13117);
nand U13593 (N_13593,N_13202,N_13010);
nand U13594 (N_13594,N_13304,N_13428);
nand U13595 (N_13595,N_13217,N_13317);
and U13596 (N_13596,N_13031,N_13267);
and U13597 (N_13597,N_13003,N_13281);
nand U13598 (N_13598,N_13330,N_13095);
nor U13599 (N_13599,N_13333,N_13475);
and U13600 (N_13600,N_13308,N_13291);
nor U13601 (N_13601,N_13386,N_13189);
nor U13602 (N_13602,N_13021,N_13036);
nand U13603 (N_13603,N_13227,N_13404);
nor U13604 (N_13604,N_13020,N_13400);
nand U13605 (N_13605,N_13172,N_13015);
xnor U13606 (N_13606,N_13265,N_13138);
nor U13607 (N_13607,N_13455,N_13377);
nor U13608 (N_13608,N_13153,N_13382);
xor U13609 (N_13609,N_13087,N_13496);
and U13610 (N_13610,N_13007,N_13335);
nand U13611 (N_13611,N_13183,N_13261);
and U13612 (N_13612,N_13260,N_13131);
or U13613 (N_13613,N_13350,N_13084);
xnor U13614 (N_13614,N_13233,N_13383);
or U13615 (N_13615,N_13210,N_13085);
nor U13616 (N_13616,N_13274,N_13275);
or U13617 (N_13617,N_13466,N_13083);
nor U13618 (N_13618,N_13091,N_13380);
or U13619 (N_13619,N_13229,N_13045);
nor U13620 (N_13620,N_13094,N_13327);
or U13621 (N_13621,N_13067,N_13497);
xnor U13622 (N_13622,N_13061,N_13343);
or U13623 (N_13623,N_13216,N_13155);
and U13624 (N_13624,N_13306,N_13079);
xnor U13625 (N_13625,N_13096,N_13409);
and U13626 (N_13626,N_13066,N_13154);
and U13627 (N_13627,N_13188,N_13417);
and U13628 (N_13628,N_13437,N_13235);
nand U13629 (N_13629,N_13403,N_13303);
and U13630 (N_13630,N_13060,N_13459);
and U13631 (N_13631,N_13411,N_13310);
nor U13632 (N_13632,N_13442,N_13212);
nand U13633 (N_13633,N_13039,N_13075);
nand U13634 (N_13634,N_13230,N_13331);
or U13635 (N_13635,N_13033,N_13349);
and U13636 (N_13636,N_13081,N_13201);
and U13637 (N_13637,N_13270,N_13363);
and U13638 (N_13638,N_13132,N_13299);
nand U13639 (N_13639,N_13352,N_13245);
xnor U13640 (N_13640,N_13179,N_13082);
nand U13641 (N_13641,N_13126,N_13289);
nor U13642 (N_13642,N_13361,N_13246);
nor U13643 (N_13643,N_13177,N_13370);
nand U13644 (N_13644,N_13171,N_13074);
nand U13645 (N_13645,N_13209,N_13482);
and U13646 (N_13646,N_13358,N_13041);
nor U13647 (N_13647,N_13163,N_13121);
and U13648 (N_13648,N_13342,N_13469);
nor U13649 (N_13649,N_13018,N_13476);
or U13650 (N_13650,N_13271,N_13314);
or U13651 (N_13651,N_13173,N_13215);
nand U13652 (N_13652,N_13321,N_13252);
nor U13653 (N_13653,N_13434,N_13488);
or U13654 (N_13654,N_13211,N_13430);
nand U13655 (N_13655,N_13348,N_13241);
and U13656 (N_13656,N_13347,N_13461);
or U13657 (N_13657,N_13040,N_13247);
or U13658 (N_13658,N_13435,N_13042);
xnor U13659 (N_13659,N_13220,N_13058);
xor U13660 (N_13660,N_13148,N_13098);
nor U13661 (N_13661,N_13110,N_13205);
and U13662 (N_13662,N_13168,N_13037);
and U13663 (N_13663,N_13292,N_13169);
xnor U13664 (N_13664,N_13107,N_13483);
nor U13665 (N_13665,N_13422,N_13238);
nor U13666 (N_13666,N_13099,N_13396);
nand U13667 (N_13667,N_13116,N_13114);
nor U13668 (N_13668,N_13318,N_13192);
nand U13669 (N_13669,N_13405,N_13093);
nand U13670 (N_13670,N_13315,N_13340);
or U13671 (N_13671,N_13499,N_13043);
nand U13672 (N_13672,N_13112,N_13046);
or U13673 (N_13673,N_13440,N_13379);
and U13674 (N_13674,N_13353,N_13324);
nand U13675 (N_13675,N_13001,N_13388);
or U13676 (N_13676,N_13390,N_13128);
nor U13677 (N_13677,N_13468,N_13051);
nor U13678 (N_13678,N_13069,N_13239);
and U13679 (N_13679,N_13293,N_13490);
nand U13680 (N_13680,N_13086,N_13130);
and U13681 (N_13681,N_13053,N_13196);
xnor U13682 (N_13682,N_13219,N_13384);
nor U13683 (N_13683,N_13311,N_13372);
or U13684 (N_13684,N_13149,N_13064);
nand U13685 (N_13685,N_13120,N_13181);
nand U13686 (N_13686,N_13478,N_13186);
nand U13687 (N_13687,N_13124,N_13151);
xor U13688 (N_13688,N_13156,N_13145);
nand U13689 (N_13689,N_13125,N_13325);
nand U13690 (N_13690,N_13406,N_13059);
and U13691 (N_13691,N_13465,N_13433);
xor U13692 (N_13692,N_13391,N_13413);
nor U13693 (N_13693,N_13454,N_13054);
nor U13694 (N_13694,N_13282,N_13161);
nor U13695 (N_13695,N_13326,N_13450);
xnor U13696 (N_13696,N_13101,N_13047);
and U13697 (N_13697,N_13479,N_13073);
or U13698 (N_13698,N_13258,N_13072);
and U13699 (N_13699,N_13213,N_13432);
nand U13700 (N_13700,N_13399,N_13458);
xnor U13701 (N_13701,N_13254,N_13263);
and U13702 (N_13702,N_13029,N_13102);
or U13703 (N_13703,N_13397,N_13464);
or U13704 (N_13704,N_13135,N_13407);
nor U13705 (N_13705,N_13104,N_13048);
and U13706 (N_13706,N_13234,N_13164);
xor U13707 (N_13707,N_13184,N_13022);
and U13708 (N_13708,N_13065,N_13140);
nor U13709 (N_13709,N_13472,N_13178);
nand U13710 (N_13710,N_13190,N_13197);
xnor U13711 (N_13711,N_13334,N_13451);
nand U13712 (N_13712,N_13272,N_13221);
nand U13713 (N_13713,N_13077,N_13295);
or U13714 (N_13714,N_13165,N_13257);
nor U13715 (N_13715,N_13141,N_13057);
xor U13716 (N_13716,N_13362,N_13166);
and U13717 (N_13717,N_13319,N_13092);
nand U13718 (N_13718,N_13000,N_13357);
or U13719 (N_13719,N_13025,N_13005);
nand U13720 (N_13720,N_13218,N_13341);
nand U13721 (N_13721,N_13167,N_13023);
nand U13722 (N_13722,N_13185,N_13243);
and U13723 (N_13723,N_13410,N_13416);
or U13724 (N_13724,N_13269,N_13313);
nand U13725 (N_13725,N_13264,N_13485);
xor U13726 (N_13726,N_13147,N_13194);
and U13727 (N_13727,N_13373,N_13231);
xnor U13728 (N_13728,N_13236,N_13108);
nor U13729 (N_13729,N_13088,N_13225);
nand U13730 (N_13730,N_13206,N_13012);
and U13731 (N_13731,N_13312,N_13288);
nor U13732 (N_13732,N_13129,N_13491);
xor U13733 (N_13733,N_13160,N_13387);
nor U13734 (N_13734,N_13336,N_13191);
nand U13735 (N_13735,N_13457,N_13103);
and U13736 (N_13736,N_13118,N_13415);
nand U13737 (N_13737,N_13426,N_13486);
and U13738 (N_13738,N_13294,N_13371);
nand U13739 (N_13739,N_13366,N_13487);
and U13740 (N_13740,N_13495,N_13187);
nor U13741 (N_13741,N_13278,N_13423);
and U13742 (N_13742,N_13493,N_13240);
and U13743 (N_13743,N_13316,N_13408);
nand U13744 (N_13744,N_13062,N_13089);
xnor U13745 (N_13745,N_13284,N_13471);
nor U13746 (N_13746,N_13436,N_13369);
and U13747 (N_13747,N_13044,N_13266);
xnor U13748 (N_13748,N_13467,N_13122);
xor U13749 (N_13749,N_13381,N_13438);
or U13750 (N_13750,N_13082,N_13456);
nor U13751 (N_13751,N_13163,N_13271);
and U13752 (N_13752,N_13353,N_13117);
and U13753 (N_13753,N_13131,N_13283);
nand U13754 (N_13754,N_13220,N_13383);
or U13755 (N_13755,N_13339,N_13422);
nand U13756 (N_13756,N_13192,N_13166);
and U13757 (N_13757,N_13489,N_13029);
xnor U13758 (N_13758,N_13017,N_13485);
or U13759 (N_13759,N_13159,N_13315);
and U13760 (N_13760,N_13243,N_13395);
nor U13761 (N_13761,N_13357,N_13166);
xor U13762 (N_13762,N_13484,N_13384);
and U13763 (N_13763,N_13388,N_13015);
xnor U13764 (N_13764,N_13320,N_13351);
nor U13765 (N_13765,N_13367,N_13385);
or U13766 (N_13766,N_13259,N_13031);
or U13767 (N_13767,N_13159,N_13153);
nor U13768 (N_13768,N_13407,N_13497);
nor U13769 (N_13769,N_13232,N_13305);
nor U13770 (N_13770,N_13159,N_13223);
or U13771 (N_13771,N_13109,N_13173);
xor U13772 (N_13772,N_13041,N_13256);
or U13773 (N_13773,N_13439,N_13003);
or U13774 (N_13774,N_13341,N_13480);
or U13775 (N_13775,N_13195,N_13145);
and U13776 (N_13776,N_13108,N_13435);
nor U13777 (N_13777,N_13377,N_13145);
or U13778 (N_13778,N_13431,N_13380);
xnor U13779 (N_13779,N_13387,N_13075);
and U13780 (N_13780,N_13241,N_13474);
and U13781 (N_13781,N_13486,N_13249);
xor U13782 (N_13782,N_13339,N_13160);
xnor U13783 (N_13783,N_13050,N_13070);
nand U13784 (N_13784,N_13190,N_13366);
nor U13785 (N_13785,N_13492,N_13382);
nand U13786 (N_13786,N_13239,N_13369);
nor U13787 (N_13787,N_13405,N_13190);
nor U13788 (N_13788,N_13451,N_13037);
xor U13789 (N_13789,N_13454,N_13399);
nand U13790 (N_13790,N_13395,N_13486);
xnor U13791 (N_13791,N_13450,N_13413);
nand U13792 (N_13792,N_13476,N_13209);
and U13793 (N_13793,N_13152,N_13468);
or U13794 (N_13794,N_13199,N_13164);
nor U13795 (N_13795,N_13329,N_13443);
nor U13796 (N_13796,N_13410,N_13423);
nor U13797 (N_13797,N_13118,N_13068);
nand U13798 (N_13798,N_13164,N_13287);
and U13799 (N_13799,N_13150,N_13428);
nor U13800 (N_13800,N_13125,N_13086);
or U13801 (N_13801,N_13156,N_13465);
and U13802 (N_13802,N_13053,N_13184);
nand U13803 (N_13803,N_13090,N_13420);
and U13804 (N_13804,N_13357,N_13132);
nand U13805 (N_13805,N_13158,N_13019);
nor U13806 (N_13806,N_13092,N_13093);
nand U13807 (N_13807,N_13487,N_13182);
or U13808 (N_13808,N_13459,N_13303);
or U13809 (N_13809,N_13353,N_13379);
nor U13810 (N_13810,N_13013,N_13024);
nor U13811 (N_13811,N_13012,N_13108);
nand U13812 (N_13812,N_13491,N_13251);
or U13813 (N_13813,N_13298,N_13382);
xnor U13814 (N_13814,N_13467,N_13322);
nor U13815 (N_13815,N_13384,N_13310);
nand U13816 (N_13816,N_13068,N_13059);
and U13817 (N_13817,N_13281,N_13023);
nor U13818 (N_13818,N_13079,N_13177);
and U13819 (N_13819,N_13378,N_13420);
nand U13820 (N_13820,N_13187,N_13037);
nor U13821 (N_13821,N_13257,N_13438);
and U13822 (N_13822,N_13311,N_13082);
and U13823 (N_13823,N_13262,N_13192);
nor U13824 (N_13824,N_13217,N_13153);
or U13825 (N_13825,N_13312,N_13221);
nor U13826 (N_13826,N_13090,N_13331);
or U13827 (N_13827,N_13283,N_13291);
nand U13828 (N_13828,N_13326,N_13007);
xor U13829 (N_13829,N_13360,N_13328);
and U13830 (N_13830,N_13307,N_13082);
nor U13831 (N_13831,N_13159,N_13463);
xor U13832 (N_13832,N_13140,N_13039);
or U13833 (N_13833,N_13195,N_13494);
xnor U13834 (N_13834,N_13193,N_13239);
nor U13835 (N_13835,N_13126,N_13097);
nand U13836 (N_13836,N_13304,N_13379);
and U13837 (N_13837,N_13359,N_13302);
or U13838 (N_13838,N_13215,N_13021);
and U13839 (N_13839,N_13473,N_13335);
and U13840 (N_13840,N_13224,N_13036);
nor U13841 (N_13841,N_13128,N_13189);
or U13842 (N_13842,N_13448,N_13386);
nor U13843 (N_13843,N_13210,N_13179);
and U13844 (N_13844,N_13137,N_13070);
and U13845 (N_13845,N_13188,N_13201);
or U13846 (N_13846,N_13308,N_13070);
nor U13847 (N_13847,N_13283,N_13391);
nor U13848 (N_13848,N_13103,N_13488);
xor U13849 (N_13849,N_13034,N_13143);
nor U13850 (N_13850,N_13163,N_13060);
nand U13851 (N_13851,N_13492,N_13362);
or U13852 (N_13852,N_13127,N_13314);
and U13853 (N_13853,N_13127,N_13236);
or U13854 (N_13854,N_13017,N_13111);
nor U13855 (N_13855,N_13143,N_13396);
nand U13856 (N_13856,N_13084,N_13358);
and U13857 (N_13857,N_13310,N_13047);
xnor U13858 (N_13858,N_13241,N_13151);
nor U13859 (N_13859,N_13263,N_13124);
nor U13860 (N_13860,N_13030,N_13181);
or U13861 (N_13861,N_13087,N_13362);
nor U13862 (N_13862,N_13265,N_13225);
or U13863 (N_13863,N_13234,N_13057);
nor U13864 (N_13864,N_13044,N_13244);
or U13865 (N_13865,N_13043,N_13220);
xnor U13866 (N_13866,N_13310,N_13266);
xor U13867 (N_13867,N_13287,N_13383);
xnor U13868 (N_13868,N_13011,N_13002);
and U13869 (N_13869,N_13149,N_13382);
xor U13870 (N_13870,N_13172,N_13188);
or U13871 (N_13871,N_13404,N_13032);
xnor U13872 (N_13872,N_13149,N_13155);
nand U13873 (N_13873,N_13115,N_13058);
nor U13874 (N_13874,N_13220,N_13448);
or U13875 (N_13875,N_13286,N_13171);
xnor U13876 (N_13876,N_13478,N_13485);
and U13877 (N_13877,N_13407,N_13179);
nand U13878 (N_13878,N_13047,N_13284);
nor U13879 (N_13879,N_13389,N_13474);
and U13880 (N_13880,N_13452,N_13329);
and U13881 (N_13881,N_13373,N_13498);
or U13882 (N_13882,N_13149,N_13399);
or U13883 (N_13883,N_13088,N_13318);
xnor U13884 (N_13884,N_13413,N_13410);
nor U13885 (N_13885,N_13227,N_13194);
xnor U13886 (N_13886,N_13205,N_13338);
and U13887 (N_13887,N_13439,N_13127);
and U13888 (N_13888,N_13344,N_13318);
nor U13889 (N_13889,N_13316,N_13447);
or U13890 (N_13890,N_13141,N_13089);
or U13891 (N_13891,N_13345,N_13325);
xor U13892 (N_13892,N_13320,N_13315);
and U13893 (N_13893,N_13432,N_13043);
nand U13894 (N_13894,N_13089,N_13202);
nand U13895 (N_13895,N_13272,N_13360);
and U13896 (N_13896,N_13244,N_13291);
or U13897 (N_13897,N_13131,N_13488);
and U13898 (N_13898,N_13258,N_13293);
and U13899 (N_13899,N_13286,N_13455);
or U13900 (N_13900,N_13164,N_13177);
or U13901 (N_13901,N_13125,N_13220);
and U13902 (N_13902,N_13101,N_13174);
nor U13903 (N_13903,N_13419,N_13363);
nand U13904 (N_13904,N_13410,N_13300);
nand U13905 (N_13905,N_13083,N_13051);
and U13906 (N_13906,N_13368,N_13051);
nor U13907 (N_13907,N_13245,N_13417);
and U13908 (N_13908,N_13049,N_13356);
nand U13909 (N_13909,N_13486,N_13065);
nor U13910 (N_13910,N_13322,N_13351);
nand U13911 (N_13911,N_13428,N_13190);
nand U13912 (N_13912,N_13370,N_13289);
or U13913 (N_13913,N_13013,N_13006);
nand U13914 (N_13914,N_13191,N_13205);
nor U13915 (N_13915,N_13177,N_13484);
or U13916 (N_13916,N_13032,N_13382);
nor U13917 (N_13917,N_13296,N_13035);
or U13918 (N_13918,N_13283,N_13145);
nor U13919 (N_13919,N_13333,N_13008);
xnor U13920 (N_13920,N_13421,N_13108);
nand U13921 (N_13921,N_13250,N_13194);
and U13922 (N_13922,N_13286,N_13384);
xnor U13923 (N_13923,N_13014,N_13100);
nand U13924 (N_13924,N_13344,N_13404);
xor U13925 (N_13925,N_13404,N_13195);
nand U13926 (N_13926,N_13414,N_13275);
nor U13927 (N_13927,N_13310,N_13034);
nor U13928 (N_13928,N_13445,N_13309);
and U13929 (N_13929,N_13309,N_13173);
nand U13930 (N_13930,N_13377,N_13129);
nand U13931 (N_13931,N_13249,N_13061);
and U13932 (N_13932,N_13065,N_13432);
and U13933 (N_13933,N_13105,N_13216);
nor U13934 (N_13934,N_13046,N_13128);
nand U13935 (N_13935,N_13198,N_13371);
or U13936 (N_13936,N_13150,N_13476);
nor U13937 (N_13937,N_13244,N_13448);
nand U13938 (N_13938,N_13290,N_13043);
xnor U13939 (N_13939,N_13232,N_13140);
nor U13940 (N_13940,N_13095,N_13479);
xor U13941 (N_13941,N_13120,N_13081);
xnor U13942 (N_13942,N_13498,N_13486);
xor U13943 (N_13943,N_13021,N_13066);
nand U13944 (N_13944,N_13167,N_13468);
nand U13945 (N_13945,N_13141,N_13436);
and U13946 (N_13946,N_13423,N_13050);
xor U13947 (N_13947,N_13031,N_13408);
and U13948 (N_13948,N_13155,N_13426);
or U13949 (N_13949,N_13038,N_13385);
nor U13950 (N_13950,N_13325,N_13220);
xor U13951 (N_13951,N_13202,N_13366);
or U13952 (N_13952,N_13455,N_13444);
and U13953 (N_13953,N_13452,N_13273);
nor U13954 (N_13954,N_13499,N_13082);
or U13955 (N_13955,N_13437,N_13356);
or U13956 (N_13956,N_13399,N_13086);
and U13957 (N_13957,N_13397,N_13120);
xor U13958 (N_13958,N_13210,N_13299);
xnor U13959 (N_13959,N_13470,N_13447);
and U13960 (N_13960,N_13124,N_13246);
nand U13961 (N_13961,N_13489,N_13465);
nand U13962 (N_13962,N_13485,N_13172);
nand U13963 (N_13963,N_13223,N_13136);
nand U13964 (N_13964,N_13273,N_13375);
xnor U13965 (N_13965,N_13277,N_13319);
or U13966 (N_13966,N_13167,N_13026);
nand U13967 (N_13967,N_13130,N_13327);
and U13968 (N_13968,N_13074,N_13038);
or U13969 (N_13969,N_13428,N_13193);
xnor U13970 (N_13970,N_13475,N_13228);
nand U13971 (N_13971,N_13094,N_13271);
or U13972 (N_13972,N_13357,N_13466);
xnor U13973 (N_13973,N_13329,N_13431);
nand U13974 (N_13974,N_13289,N_13227);
xnor U13975 (N_13975,N_13184,N_13411);
xnor U13976 (N_13976,N_13470,N_13238);
and U13977 (N_13977,N_13014,N_13163);
nand U13978 (N_13978,N_13419,N_13122);
and U13979 (N_13979,N_13119,N_13228);
and U13980 (N_13980,N_13452,N_13415);
nor U13981 (N_13981,N_13349,N_13168);
nor U13982 (N_13982,N_13481,N_13165);
nor U13983 (N_13983,N_13178,N_13002);
and U13984 (N_13984,N_13472,N_13087);
xnor U13985 (N_13985,N_13284,N_13338);
or U13986 (N_13986,N_13455,N_13387);
nor U13987 (N_13987,N_13302,N_13183);
or U13988 (N_13988,N_13037,N_13035);
xor U13989 (N_13989,N_13142,N_13228);
nand U13990 (N_13990,N_13259,N_13002);
xor U13991 (N_13991,N_13044,N_13320);
nand U13992 (N_13992,N_13345,N_13391);
nand U13993 (N_13993,N_13312,N_13032);
nor U13994 (N_13994,N_13454,N_13019);
nor U13995 (N_13995,N_13096,N_13327);
nand U13996 (N_13996,N_13463,N_13234);
nand U13997 (N_13997,N_13342,N_13004);
xnor U13998 (N_13998,N_13460,N_13119);
or U13999 (N_13999,N_13221,N_13464);
nor U14000 (N_14000,N_13703,N_13937);
nor U14001 (N_14001,N_13522,N_13887);
xnor U14002 (N_14002,N_13654,N_13899);
nor U14003 (N_14003,N_13769,N_13718);
and U14004 (N_14004,N_13627,N_13646);
nand U14005 (N_14005,N_13733,N_13904);
nor U14006 (N_14006,N_13530,N_13572);
or U14007 (N_14007,N_13551,N_13534);
or U14008 (N_14008,N_13704,N_13775);
or U14009 (N_14009,N_13818,N_13524);
nor U14010 (N_14010,N_13556,N_13568);
xor U14011 (N_14011,N_13675,N_13795);
nor U14012 (N_14012,N_13571,N_13777);
and U14013 (N_14013,N_13555,N_13976);
nand U14014 (N_14014,N_13631,N_13584);
and U14015 (N_14015,N_13518,N_13563);
or U14016 (N_14016,N_13826,N_13812);
and U14017 (N_14017,N_13544,N_13916);
nor U14018 (N_14018,N_13501,N_13954);
xnor U14019 (N_14019,N_13664,N_13784);
nor U14020 (N_14020,N_13810,N_13838);
and U14021 (N_14021,N_13925,N_13655);
nand U14022 (N_14022,N_13939,N_13787);
xnor U14023 (N_14023,N_13855,N_13756);
or U14024 (N_14024,N_13870,N_13837);
or U14025 (N_14025,N_13734,N_13510);
and U14026 (N_14026,N_13514,N_13749);
or U14027 (N_14027,N_13730,N_13578);
or U14028 (N_14028,N_13716,N_13809);
nor U14029 (N_14029,N_13594,N_13575);
xnor U14030 (N_14030,N_13850,N_13685);
nand U14031 (N_14031,N_13679,N_13545);
nand U14032 (N_14032,N_13695,N_13823);
xor U14033 (N_14033,N_13738,N_13634);
nand U14034 (N_14034,N_13677,N_13764);
and U14035 (N_14035,N_13592,N_13553);
or U14036 (N_14036,N_13640,N_13794);
or U14037 (N_14037,N_13877,N_13593);
nor U14038 (N_14038,N_13596,N_13540);
or U14039 (N_14039,N_13882,N_13909);
or U14040 (N_14040,N_13504,N_13755);
xor U14041 (N_14041,N_13625,N_13919);
and U14042 (N_14042,N_13933,N_13595);
and U14043 (N_14043,N_13583,N_13952);
or U14044 (N_14044,N_13624,N_13814);
and U14045 (N_14045,N_13918,N_13588);
nand U14046 (N_14046,N_13985,N_13961);
nand U14047 (N_14047,N_13732,N_13642);
xnor U14048 (N_14048,N_13758,N_13967);
xor U14049 (N_14049,N_13917,N_13561);
nor U14050 (N_14050,N_13955,N_13512);
or U14051 (N_14051,N_13715,N_13932);
nor U14052 (N_14052,N_13552,N_13519);
and U14053 (N_14053,N_13743,N_13891);
nand U14054 (N_14054,N_13778,N_13859);
nand U14055 (N_14055,N_13765,N_13987);
and U14056 (N_14056,N_13830,N_13963);
nor U14057 (N_14057,N_13774,N_13750);
and U14058 (N_14058,N_13740,N_13520);
nand U14059 (N_14059,N_13569,N_13876);
or U14060 (N_14060,N_13525,N_13745);
nand U14061 (N_14061,N_13880,N_13966);
nand U14062 (N_14062,N_13731,N_13742);
xor U14063 (N_14063,N_13537,N_13688);
or U14064 (N_14064,N_13705,N_13557);
xor U14065 (N_14065,N_13603,N_13943);
and U14066 (N_14066,N_13566,N_13879);
xor U14067 (N_14067,N_13529,N_13936);
or U14068 (N_14068,N_13687,N_13548);
nand U14069 (N_14069,N_13788,N_13969);
and U14070 (N_14070,N_13820,N_13934);
and U14071 (N_14071,N_13911,N_13808);
nand U14072 (N_14072,N_13698,N_13617);
and U14073 (N_14073,N_13727,N_13893);
nand U14074 (N_14074,N_13565,N_13509);
xor U14075 (N_14075,N_13856,N_13950);
nor U14076 (N_14076,N_13533,N_13801);
nor U14077 (N_14077,N_13999,N_13517);
and U14078 (N_14078,N_13921,N_13662);
nor U14079 (N_14079,N_13652,N_13725);
and U14080 (N_14080,N_13938,N_13948);
or U14081 (N_14081,N_13586,N_13729);
or U14082 (N_14082,N_13959,N_13549);
nor U14083 (N_14083,N_13598,N_13811);
and U14084 (N_14084,N_13960,N_13711);
and U14085 (N_14085,N_13979,N_13992);
or U14086 (N_14086,N_13860,N_13941);
and U14087 (N_14087,N_13721,N_13700);
and U14088 (N_14088,N_13828,N_13946);
nor U14089 (N_14089,N_13706,N_13739);
or U14090 (N_14090,N_13886,N_13709);
nand U14091 (N_14091,N_13589,N_13789);
xnor U14092 (N_14092,N_13993,N_13573);
or U14093 (N_14093,N_13892,N_13928);
xnor U14094 (N_14094,N_13958,N_13667);
nor U14095 (N_14095,N_13854,N_13682);
or U14096 (N_14096,N_13824,N_13831);
xor U14097 (N_14097,N_13951,N_13931);
xnor U14098 (N_14098,N_13577,N_13550);
nand U14099 (N_14099,N_13761,N_13659);
and U14100 (N_14100,N_13800,N_13815);
and U14101 (N_14101,N_13696,N_13945);
and U14102 (N_14102,N_13644,N_13723);
xnor U14103 (N_14103,N_13641,N_13957);
or U14104 (N_14104,N_13620,N_13773);
or U14105 (N_14105,N_13947,N_13615);
nor U14106 (N_14106,N_13591,N_13796);
xor U14107 (N_14107,N_13690,N_13759);
nor U14108 (N_14108,N_13744,N_13719);
nor U14109 (N_14109,N_13944,N_13962);
xnor U14110 (N_14110,N_13531,N_13871);
and U14111 (N_14111,N_13513,N_13600);
or U14112 (N_14112,N_13579,N_13748);
xor U14113 (N_14113,N_13559,N_13608);
nand U14114 (N_14114,N_13873,N_13968);
nand U14115 (N_14115,N_13606,N_13973);
nand U14116 (N_14116,N_13665,N_13768);
xnor U14117 (N_14117,N_13953,N_13663);
xor U14118 (N_14118,N_13940,N_13770);
or U14119 (N_14119,N_13956,N_13849);
and U14120 (N_14120,N_13636,N_13680);
xnor U14121 (N_14121,N_13635,N_13914);
nor U14122 (N_14122,N_13825,N_13997);
nor U14123 (N_14123,N_13762,N_13527);
or U14124 (N_14124,N_13532,N_13930);
nor U14125 (N_14125,N_13922,N_13853);
nor U14126 (N_14126,N_13839,N_13689);
or U14127 (N_14127,N_13741,N_13781);
nand U14128 (N_14128,N_13683,N_13657);
nand U14129 (N_14129,N_13907,N_13707);
and U14130 (N_14130,N_13701,N_13576);
or U14131 (N_14131,N_13862,N_13912);
nand U14132 (N_14132,N_13982,N_13543);
xnor U14133 (N_14133,N_13878,N_13666);
and U14134 (N_14134,N_13580,N_13981);
xnor U14135 (N_14135,N_13728,N_13602);
nor U14136 (N_14136,N_13697,N_13502);
nor U14137 (N_14137,N_13846,N_13998);
nand U14138 (N_14138,N_13511,N_13710);
xnor U14139 (N_14139,N_13851,N_13747);
and U14140 (N_14140,N_13714,N_13868);
xnor U14141 (N_14141,N_13638,N_13763);
nand U14142 (N_14142,N_13889,N_13791);
nor U14143 (N_14143,N_13622,N_13567);
xor U14144 (N_14144,N_13515,N_13673);
xnor U14145 (N_14145,N_13713,N_13793);
nand U14146 (N_14146,N_13807,N_13751);
or U14147 (N_14147,N_13819,N_13983);
xnor U14148 (N_14148,N_13900,N_13872);
nand U14149 (N_14149,N_13570,N_13726);
nor U14150 (N_14150,N_13735,N_13866);
nand U14151 (N_14151,N_13874,N_13536);
nand U14152 (N_14152,N_13970,N_13616);
xor U14153 (N_14153,N_13935,N_13564);
and U14154 (N_14154,N_13585,N_13975);
xor U14155 (N_14155,N_13516,N_13599);
nor U14156 (N_14156,N_13613,N_13581);
or U14157 (N_14157,N_13798,N_13782);
and U14158 (N_14158,N_13822,N_13843);
nor U14159 (N_14159,N_13712,N_13597);
nand U14160 (N_14160,N_13648,N_13857);
and U14161 (N_14161,N_13834,N_13990);
xnor U14162 (N_14162,N_13674,N_13858);
nor U14163 (N_14163,N_13977,N_13875);
xor U14164 (N_14164,N_13754,N_13864);
or U14165 (N_14165,N_13890,N_13653);
nor U14166 (N_14166,N_13628,N_13574);
nand U14167 (N_14167,N_13865,N_13996);
nand U14168 (N_14168,N_13994,N_13766);
and U14169 (N_14169,N_13546,N_13881);
nor U14170 (N_14170,N_13903,N_13560);
nor U14171 (N_14171,N_13724,N_13980);
nor U14172 (N_14172,N_13671,N_13651);
and U14173 (N_14173,N_13813,N_13924);
xor U14174 (N_14174,N_13772,N_13708);
nor U14175 (N_14175,N_13852,N_13799);
and U14176 (N_14176,N_13783,N_13737);
nor U14177 (N_14177,N_13978,N_13619);
or U14178 (N_14178,N_13604,N_13792);
nor U14179 (N_14179,N_13972,N_13630);
nand U14180 (N_14180,N_13895,N_13623);
or U14181 (N_14181,N_13647,N_13609);
nor U14182 (N_14182,N_13645,N_13612);
xor U14183 (N_14183,N_13684,N_13717);
xor U14184 (N_14184,N_13929,N_13670);
nand U14185 (N_14185,N_13842,N_13986);
nor U14186 (N_14186,N_13785,N_13582);
nand U14187 (N_14187,N_13720,N_13605);
nand U14188 (N_14188,N_13897,N_13554);
nand U14189 (N_14189,N_13505,N_13913);
or U14190 (N_14190,N_13614,N_13632);
nand U14191 (N_14191,N_13804,N_13649);
nor U14192 (N_14192,N_13643,N_13507);
xnor U14193 (N_14193,N_13780,N_13844);
nand U14194 (N_14194,N_13558,N_13503);
or U14195 (N_14195,N_13836,N_13500);
and U14196 (N_14196,N_13542,N_13869);
or U14197 (N_14197,N_13539,N_13521);
or U14198 (N_14198,N_13535,N_13757);
xor U14199 (N_14199,N_13526,N_13767);
or U14200 (N_14200,N_13984,N_13610);
xor U14201 (N_14201,N_13845,N_13686);
xor U14202 (N_14202,N_13746,N_13989);
and U14203 (N_14203,N_13906,N_13523);
nand U14204 (N_14204,N_13702,N_13833);
xnor U14205 (N_14205,N_13776,N_13910);
xnor U14206 (N_14206,N_13885,N_13668);
nand U14207 (N_14207,N_13621,N_13779);
xor U14208 (N_14208,N_13661,N_13816);
or U14209 (N_14209,N_13760,N_13965);
or U14210 (N_14210,N_13678,N_13607);
nand U14211 (N_14211,N_13506,N_13691);
nand U14212 (N_14212,N_13991,N_13867);
or U14213 (N_14213,N_13841,N_13541);
or U14214 (N_14214,N_13848,N_13672);
or U14215 (N_14215,N_13547,N_13988);
nor U14216 (N_14216,N_13650,N_13894);
nand U14217 (N_14217,N_13884,N_13806);
xor U14218 (N_14218,N_13883,N_13692);
and U14219 (N_14219,N_13508,N_13771);
or U14220 (N_14220,N_13656,N_13821);
xnor U14221 (N_14221,N_13902,N_13601);
nand U14222 (N_14222,N_13669,N_13786);
and U14223 (N_14223,N_13611,N_13920);
or U14224 (N_14224,N_13888,N_13949);
nand U14225 (N_14225,N_13736,N_13974);
nand U14226 (N_14226,N_13528,N_13639);
or U14227 (N_14227,N_13681,N_13618);
nor U14228 (N_14228,N_13829,N_13908);
and U14229 (N_14229,N_13840,N_13832);
nand U14230 (N_14230,N_13896,N_13964);
or U14231 (N_14231,N_13995,N_13926);
and U14232 (N_14232,N_13626,N_13722);
or U14233 (N_14233,N_13587,N_13658);
and U14234 (N_14234,N_13752,N_13693);
nand U14235 (N_14235,N_13633,N_13915);
or U14236 (N_14236,N_13861,N_13847);
nand U14237 (N_14237,N_13790,N_13905);
xor U14238 (N_14238,N_13817,N_13637);
xor U14239 (N_14239,N_13753,N_13797);
or U14240 (N_14240,N_13927,N_13863);
nand U14241 (N_14241,N_13590,N_13562);
xnor U14242 (N_14242,N_13676,N_13694);
xor U14243 (N_14243,N_13901,N_13803);
or U14244 (N_14244,N_13835,N_13629);
xor U14245 (N_14245,N_13802,N_13699);
nand U14246 (N_14246,N_13923,N_13827);
or U14247 (N_14247,N_13660,N_13538);
nor U14248 (N_14248,N_13942,N_13898);
xnor U14249 (N_14249,N_13805,N_13971);
nand U14250 (N_14250,N_13651,N_13644);
xnor U14251 (N_14251,N_13906,N_13698);
and U14252 (N_14252,N_13759,N_13556);
nor U14253 (N_14253,N_13694,N_13639);
xor U14254 (N_14254,N_13590,N_13710);
nand U14255 (N_14255,N_13993,N_13598);
nand U14256 (N_14256,N_13781,N_13594);
nor U14257 (N_14257,N_13911,N_13711);
nand U14258 (N_14258,N_13950,N_13971);
nor U14259 (N_14259,N_13586,N_13505);
nor U14260 (N_14260,N_13985,N_13514);
nor U14261 (N_14261,N_13832,N_13618);
or U14262 (N_14262,N_13747,N_13824);
or U14263 (N_14263,N_13595,N_13841);
xnor U14264 (N_14264,N_13763,N_13898);
nor U14265 (N_14265,N_13958,N_13620);
nand U14266 (N_14266,N_13695,N_13914);
or U14267 (N_14267,N_13547,N_13971);
nand U14268 (N_14268,N_13546,N_13552);
and U14269 (N_14269,N_13880,N_13519);
and U14270 (N_14270,N_13631,N_13550);
or U14271 (N_14271,N_13936,N_13577);
nand U14272 (N_14272,N_13865,N_13878);
and U14273 (N_14273,N_13908,N_13867);
nor U14274 (N_14274,N_13548,N_13506);
and U14275 (N_14275,N_13815,N_13746);
nand U14276 (N_14276,N_13957,N_13675);
or U14277 (N_14277,N_13696,N_13518);
nand U14278 (N_14278,N_13620,N_13748);
nor U14279 (N_14279,N_13950,N_13651);
nor U14280 (N_14280,N_13788,N_13855);
nor U14281 (N_14281,N_13564,N_13988);
nor U14282 (N_14282,N_13888,N_13729);
nand U14283 (N_14283,N_13686,N_13615);
xor U14284 (N_14284,N_13538,N_13531);
and U14285 (N_14285,N_13619,N_13547);
or U14286 (N_14286,N_13720,N_13861);
and U14287 (N_14287,N_13919,N_13803);
xnor U14288 (N_14288,N_13860,N_13867);
xor U14289 (N_14289,N_13813,N_13946);
nor U14290 (N_14290,N_13920,N_13927);
and U14291 (N_14291,N_13996,N_13560);
xnor U14292 (N_14292,N_13675,N_13710);
or U14293 (N_14293,N_13868,N_13560);
xor U14294 (N_14294,N_13715,N_13639);
xor U14295 (N_14295,N_13891,N_13574);
nor U14296 (N_14296,N_13543,N_13839);
or U14297 (N_14297,N_13685,N_13932);
nor U14298 (N_14298,N_13729,N_13749);
and U14299 (N_14299,N_13691,N_13629);
or U14300 (N_14300,N_13894,N_13836);
and U14301 (N_14301,N_13678,N_13748);
and U14302 (N_14302,N_13530,N_13763);
xnor U14303 (N_14303,N_13854,N_13717);
xnor U14304 (N_14304,N_13623,N_13659);
and U14305 (N_14305,N_13503,N_13705);
nand U14306 (N_14306,N_13960,N_13941);
nor U14307 (N_14307,N_13870,N_13674);
or U14308 (N_14308,N_13696,N_13821);
nand U14309 (N_14309,N_13879,N_13719);
nor U14310 (N_14310,N_13649,N_13982);
nand U14311 (N_14311,N_13825,N_13785);
xnor U14312 (N_14312,N_13908,N_13609);
and U14313 (N_14313,N_13573,N_13591);
xor U14314 (N_14314,N_13841,N_13648);
nand U14315 (N_14315,N_13907,N_13960);
nor U14316 (N_14316,N_13624,N_13905);
nand U14317 (N_14317,N_13932,N_13751);
nand U14318 (N_14318,N_13917,N_13777);
xor U14319 (N_14319,N_13782,N_13979);
or U14320 (N_14320,N_13851,N_13822);
nor U14321 (N_14321,N_13786,N_13711);
nand U14322 (N_14322,N_13578,N_13904);
nand U14323 (N_14323,N_13543,N_13591);
or U14324 (N_14324,N_13776,N_13863);
or U14325 (N_14325,N_13647,N_13614);
nor U14326 (N_14326,N_13832,N_13664);
nand U14327 (N_14327,N_13726,N_13649);
nand U14328 (N_14328,N_13886,N_13778);
and U14329 (N_14329,N_13958,N_13533);
xor U14330 (N_14330,N_13513,N_13807);
xor U14331 (N_14331,N_13586,N_13744);
or U14332 (N_14332,N_13919,N_13959);
or U14333 (N_14333,N_13512,N_13757);
or U14334 (N_14334,N_13538,N_13740);
xnor U14335 (N_14335,N_13905,N_13911);
and U14336 (N_14336,N_13542,N_13589);
or U14337 (N_14337,N_13693,N_13771);
xor U14338 (N_14338,N_13754,N_13729);
nand U14339 (N_14339,N_13636,N_13960);
nor U14340 (N_14340,N_13753,N_13947);
nor U14341 (N_14341,N_13502,N_13635);
or U14342 (N_14342,N_13666,N_13701);
nor U14343 (N_14343,N_13867,N_13677);
nor U14344 (N_14344,N_13662,N_13983);
nor U14345 (N_14345,N_13747,N_13759);
or U14346 (N_14346,N_13751,N_13654);
nand U14347 (N_14347,N_13806,N_13886);
xor U14348 (N_14348,N_13723,N_13607);
nor U14349 (N_14349,N_13871,N_13523);
nand U14350 (N_14350,N_13610,N_13944);
or U14351 (N_14351,N_13841,N_13855);
and U14352 (N_14352,N_13902,N_13611);
nand U14353 (N_14353,N_13958,N_13811);
and U14354 (N_14354,N_13560,N_13759);
and U14355 (N_14355,N_13952,N_13768);
nand U14356 (N_14356,N_13512,N_13951);
and U14357 (N_14357,N_13574,N_13543);
nor U14358 (N_14358,N_13758,N_13756);
nor U14359 (N_14359,N_13861,N_13505);
nand U14360 (N_14360,N_13739,N_13632);
nand U14361 (N_14361,N_13544,N_13659);
nand U14362 (N_14362,N_13552,N_13657);
nand U14363 (N_14363,N_13545,N_13749);
nand U14364 (N_14364,N_13751,N_13606);
nor U14365 (N_14365,N_13738,N_13675);
nand U14366 (N_14366,N_13908,N_13929);
nand U14367 (N_14367,N_13590,N_13683);
and U14368 (N_14368,N_13745,N_13768);
or U14369 (N_14369,N_13743,N_13881);
nand U14370 (N_14370,N_13652,N_13948);
xor U14371 (N_14371,N_13880,N_13515);
and U14372 (N_14372,N_13881,N_13717);
and U14373 (N_14373,N_13957,N_13838);
xnor U14374 (N_14374,N_13876,N_13568);
or U14375 (N_14375,N_13621,N_13768);
and U14376 (N_14376,N_13972,N_13652);
or U14377 (N_14377,N_13514,N_13501);
nand U14378 (N_14378,N_13621,N_13514);
and U14379 (N_14379,N_13580,N_13821);
nor U14380 (N_14380,N_13570,N_13996);
and U14381 (N_14381,N_13581,N_13745);
or U14382 (N_14382,N_13874,N_13519);
xnor U14383 (N_14383,N_13909,N_13985);
and U14384 (N_14384,N_13842,N_13863);
or U14385 (N_14385,N_13695,N_13866);
xnor U14386 (N_14386,N_13629,N_13807);
or U14387 (N_14387,N_13859,N_13759);
nand U14388 (N_14388,N_13893,N_13885);
nand U14389 (N_14389,N_13687,N_13787);
or U14390 (N_14390,N_13592,N_13991);
xor U14391 (N_14391,N_13531,N_13738);
or U14392 (N_14392,N_13721,N_13788);
xor U14393 (N_14393,N_13529,N_13915);
or U14394 (N_14394,N_13782,N_13727);
or U14395 (N_14395,N_13619,N_13818);
or U14396 (N_14396,N_13581,N_13898);
and U14397 (N_14397,N_13992,N_13676);
and U14398 (N_14398,N_13500,N_13668);
nor U14399 (N_14399,N_13625,N_13791);
or U14400 (N_14400,N_13710,N_13505);
nand U14401 (N_14401,N_13605,N_13648);
xnor U14402 (N_14402,N_13663,N_13704);
xnor U14403 (N_14403,N_13674,N_13536);
xnor U14404 (N_14404,N_13652,N_13643);
or U14405 (N_14405,N_13947,N_13529);
xor U14406 (N_14406,N_13921,N_13566);
and U14407 (N_14407,N_13786,N_13526);
or U14408 (N_14408,N_13977,N_13937);
nand U14409 (N_14409,N_13651,N_13888);
or U14410 (N_14410,N_13949,N_13566);
nand U14411 (N_14411,N_13521,N_13624);
nor U14412 (N_14412,N_13950,N_13613);
nor U14413 (N_14413,N_13538,N_13706);
xnor U14414 (N_14414,N_13539,N_13546);
and U14415 (N_14415,N_13501,N_13947);
xnor U14416 (N_14416,N_13688,N_13545);
or U14417 (N_14417,N_13852,N_13919);
or U14418 (N_14418,N_13829,N_13722);
and U14419 (N_14419,N_13966,N_13848);
nand U14420 (N_14420,N_13863,N_13690);
nor U14421 (N_14421,N_13615,N_13501);
and U14422 (N_14422,N_13596,N_13949);
nor U14423 (N_14423,N_13777,N_13842);
xnor U14424 (N_14424,N_13796,N_13668);
nor U14425 (N_14425,N_13876,N_13550);
nor U14426 (N_14426,N_13978,N_13774);
and U14427 (N_14427,N_13566,N_13920);
or U14428 (N_14428,N_13828,N_13723);
nand U14429 (N_14429,N_13865,N_13704);
or U14430 (N_14430,N_13950,N_13796);
nor U14431 (N_14431,N_13697,N_13957);
nand U14432 (N_14432,N_13859,N_13632);
or U14433 (N_14433,N_13589,N_13638);
or U14434 (N_14434,N_13770,N_13780);
or U14435 (N_14435,N_13615,N_13605);
nor U14436 (N_14436,N_13718,N_13532);
xor U14437 (N_14437,N_13615,N_13838);
or U14438 (N_14438,N_13842,N_13970);
and U14439 (N_14439,N_13758,N_13552);
nor U14440 (N_14440,N_13832,N_13922);
nand U14441 (N_14441,N_13955,N_13672);
nor U14442 (N_14442,N_13714,N_13528);
and U14443 (N_14443,N_13790,N_13660);
or U14444 (N_14444,N_13861,N_13903);
nor U14445 (N_14445,N_13989,N_13991);
nand U14446 (N_14446,N_13995,N_13789);
and U14447 (N_14447,N_13856,N_13864);
and U14448 (N_14448,N_13570,N_13956);
nand U14449 (N_14449,N_13885,N_13501);
or U14450 (N_14450,N_13542,N_13520);
or U14451 (N_14451,N_13983,N_13546);
xnor U14452 (N_14452,N_13812,N_13671);
xor U14453 (N_14453,N_13942,N_13545);
and U14454 (N_14454,N_13756,N_13654);
nand U14455 (N_14455,N_13833,N_13540);
or U14456 (N_14456,N_13677,N_13930);
or U14457 (N_14457,N_13770,N_13797);
or U14458 (N_14458,N_13527,N_13669);
nor U14459 (N_14459,N_13950,N_13829);
and U14460 (N_14460,N_13884,N_13632);
nand U14461 (N_14461,N_13733,N_13778);
or U14462 (N_14462,N_13738,N_13878);
xor U14463 (N_14463,N_13505,N_13655);
and U14464 (N_14464,N_13915,N_13631);
xor U14465 (N_14465,N_13820,N_13597);
or U14466 (N_14466,N_13824,N_13615);
nor U14467 (N_14467,N_13823,N_13912);
nand U14468 (N_14468,N_13939,N_13732);
nand U14469 (N_14469,N_13673,N_13781);
or U14470 (N_14470,N_13715,N_13588);
xnor U14471 (N_14471,N_13707,N_13658);
nand U14472 (N_14472,N_13882,N_13830);
or U14473 (N_14473,N_13574,N_13690);
xnor U14474 (N_14474,N_13662,N_13674);
xor U14475 (N_14475,N_13748,N_13773);
or U14476 (N_14476,N_13906,N_13628);
and U14477 (N_14477,N_13705,N_13747);
xnor U14478 (N_14478,N_13677,N_13520);
nor U14479 (N_14479,N_13574,N_13713);
nor U14480 (N_14480,N_13957,N_13514);
and U14481 (N_14481,N_13791,N_13728);
xor U14482 (N_14482,N_13570,N_13896);
nand U14483 (N_14483,N_13736,N_13786);
and U14484 (N_14484,N_13798,N_13932);
or U14485 (N_14485,N_13703,N_13848);
xor U14486 (N_14486,N_13619,N_13612);
nand U14487 (N_14487,N_13717,N_13572);
xor U14488 (N_14488,N_13862,N_13510);
or U14489 (N_14489,N_13694,N_13926);
nand U14490 (N_14490,N_13883,N_13737);
xor U14491 (N_14491,N_13665,N_13714);
nand U14492 (N_14492,N_13607,N_13575);
xor U14493 (N_14493,N_13637,N_13795);
nand U14494 (N_14494,N_13619,N_13993);
nor U14495 (N_14495,N_13891,N_13972);
nor U14496 (N_14496,N_13662,N_13727);
nand U14497 (N_14497,N_13969,N_13710);
nor U14498 (N_14498,N_13964,N_13750);
xnor U14499 (N_14499,N_13861,N_13979);
and U14500 (N_14500,N_14449,N_14422);
xor U14501 (N_14501,N_14218,N_14053);
nor U14502 (N_14502,N_14272,N_14370);
nor U14503 (N_14503,N_14323,N_14016);
or U14504 (N_14504,N_14222,N_14459);
xor U14505 (N_14505,N_14132,N_14011);
xnor U14506 (N_14506,N_14072,N_14262);
and U14507 (N_14507,N_14090,N_14234);
or U14508 (N_14508,N_14484,N_14056);
and U14509 (N_14509,N_14337,N_14278);
xnor U14510 (N_14510,N_14380,N_14019);
xor U14511 (N_14511,N_14462,N_14361);
xor U14512 (N_14512,N_14313,N_14372);
or U14513 (N_14513,N_14465,N_14017);
and U14514 (N_14514,N_14386,N_14379);
and U14515 (N_14515,N_14267,N_14478);
nand U14516 (N_14516,N_14051,N_14038);
nand U14517 (N_14517,N_14271,N_14345);
nand U14518 (N_14518,N_14029,N_14020);
and U14519 (N_14519,N_14421,N_14163);
nor U14520 (N_14520,N_14282,N_14155);
xnor U14521 (N_14521,N_14466,N_14169);
nor U14522 (N_14522,N_14081,N_14371);
and U14523 (N_14523,N_14205,N_14416);
and U14524 (N_14524,N_14480,N_14398);
and U14525 (N_14525,N_14110,N_14173);
and U14526 (N_14526,N_14447,N_14197);
nor U14527 (N_14527,N_14297,N_14327);
xnor U14528 (N_14528,N_14036,N_14015);
nand U14529 (N_14529,N_14409,N_14333);
and U14530 (N_14530,N_14369,N_14171);
nor U14531 (N_14531,N_14049,N_14025);
nor U14532 (N_14532,N_14292,N_14253);
nor U14533 (N_14533,N_14077,N_14136);
or U14534 (N_14534,N_14027,N_14092);
and U14535 (N_14535,N_14360,N_14074);
nand U14536 (N_14536,N_14300,N_14184);
nand U14537 (N_14537,N_14102,N_14358);
and U14538 (N_14538,N_14128,N_14474);
nand U14539 (N_14539,N_14123,N_14178);
nor U14540 (N_14540,N_14022,N_14150);
nand U14541 (N_14541,N_14080,N_14427);
xor U14542 (N_14542,N_14160,N_14387);
nand U14543 (N_14543,N_14131,N_14158);
and U14544 (N_14544,N_14341,N_14041);
nor U14545 (N_14545,N_14431,N_14194);
nand U14546 (N_14546,N_14340,N_14463);
or U14547 (N_14547,N_14349,N_14104);
or U14548 (N_14548,N_14335,N_14406);
nor U14549 (N_14549,N_14330,N_14224);
xor U14550 (N_14550,N_14185,N_14499);
nand U14551 (N_14551,N_14402,N_14070);
and U14552 (N_14552,N_14154,N_14486);
xnor U14553 (N_14553,N_14105,N_14279);
nand U14554 (N_14554,N_14035,N_14225);
and U14555 (N_14555,N_14207,N_14429);
nand U14556 (N_14556,N_14124,N_14309);
nor U14557 (N_14557,N_14311,N_14107);
and U14558 (N_14558,N_14250,N_14256);
nand U14559 (N_14559,N_14393,N_14003);
nand U14560 (N_14560,N_14277,N_14006);
nand U14561 (N_14561,N_14425,N_14164);
and U14562 (N_14562,N_14456,N_14452);
xnor U14563 (N_14563,N_14091,N_14211);
xnor U14564 (N_14564,N_14244,N_14389);
nand U14565 (N_14565,N_14426,N_14063);
or U14566 (N_14566,N_14214,N_14274);
nor U14567 (N_14567,N_14438,N_14242);
or U14568 (N_14568,N_14007,N_14415);
or U14569 (N_14569,N_14411,N_14385);
xor U14570 (N_14570,N_14428,N_14419);
or U14571 (N_14571,N_14472,N_14442);
xnor U14572 (N_14572,N_14494,N_14298);
nand U14573 (N_14573,N_14433,N_14059);
xnor U14574 (N_14574,N_14165,N_14137);
nand U14575 (N_14575,N_14336,N_14144);
nand U14576 (N_14576,N_14089,N_14210);
or U14577 (N_14577,N_14328,N_14334);
and U14578 (N_14578,N_14404,N_14170);
nor U14579 (N_14579,N_14203,N_14255);
nor U14580 (N_14580,N_14012,N_14407);
xor U14581 (N_14581,N_14257,N_14108);
or U14582 (N_14582,N_14347,N_14373);
nand U14583 (N_14583,N_14343,N_14014);
and U14584 (N_14584,N_14191,N_14451);
or U14585 (N_14585,N_14441,N_14146);
and U14586 (N_14586,N_14286,N_14213);
or U14587 (N_14587,N_14096,N_14176);
and U14588 (N_14588,N_14399,N_14045);
nor U14589 (N_14589,N_14151,N_14209);
or U14590 (N_14590,N_14078,N_14236);
xor U14591 (N_14591,N_14352,N_14457);
or U14592 (N_14592,N_14348,N_14353);
xnor U14593 (N_14593,N_14111,N_14153);
and U14594 (N_14594,N_14322,N_14062);
nor U14595 (N_14595,N_14338,N_14388);
xor U14596 (N_14596,N_14125,N_14177);
nand U14597 (N_14597,N_14187,N_14005);
nand U14598 (N_14598,N_14087,N_14375);
or U14599 (N_14599,N_14227,N_14159);
and U14600 (N_14600,N_14392,N_14147);
nor U14601 (N_14601,N_14367,N_14157);
nor U14602 (N_14602,N_14002,N_14339);
nor U14603 (N_14603,N_14182,N_14455);
nand U14604 (N_14604,N_14066,N_14445);
or U14605 (N_14605,N_14042,N_14162);
nor U14606 (N_14606,N_14302,N_14052);
or U14607 (N_14607,N_14239,N_14308);
and U14608 (N_14608,N_14305,N_14103);
or U14609 (N_14609,N_14028,N_14295);
nor U14610 (N_14610,N_14212,N_14440);
and U14611 (N_14611,N_14233,N_14098);
or U14612 (N_14612,N_14050,N_14384);
or U14613 (N_14613,N_14381,N_14307);
or U14614 (N_14614,N_14446,N_14228);
nor U14615 (N_14615,N_14405,N_14289);
nor U14616 (N_14616,N_14179,N_14458);
and U14617 (N_14617,N_14208,N_14247);
or U14618 (N_14618,N_14488,N_14057);
xnor U14619 (N_14619,N_14198,N_14116);
and U14620 (N_14620,N_14093,N_14126);
or U14621 (N_14621,N_14226,N_14134);
nor U14622 (N_14622,N_14296,N_14167);
or U14623 (N_14623,N_14493,N_14142);
and U14624 (N_14624,N_14048,N_14496);
xor U14625 (N_14625,N_14202,N_14044);
xnor U14626 (N_14626,N_14139,N_14008);
nand U14627 (N_14627,N_14265,N_14097);
nor U14628 (N_14628,N_14023,N_14141);
xnor U14629 (N_14629,N_14119,N_14100);
nor U14630 (N_14630,N_14481,N_14413);
nand U14631 (N_14631,N_14329,N_14346);
nor U14632 (N_14632,N_14362,N_14306);
nand U14633 (N_14633,N_14420,N_14200);
nor U14634 (N_14634,N_14483,N_14127);
nor U14635 (N_14635,N_14403,N_14275);
nand U14636 (N_14636,N_14396,N_14082);
or U14637 (N_14637,N_14498,N_14201);
nand U14638 (N_14638,N_14223,N_14476);
and U14639 (N_14639,N_14076,N_14193);
and U14640 (N_14640,N_14189,N_14118);
or U14641 (N_14641,N_14174,N_14383);
or U14642 (N_14642,N_14231,N_14437);
nand U14643 (N_14643,N_14248,N_14412);
nor U14644 (N_14644,N_14374,N_14460);
nand U14645 (N_14645,N_14047,N_14314);
nor U14646 (N_14646,N_14001,N_14064);
and U14647 (N_14647,N_14079,N_14325);
and U14648 (N_14648,N_14068,N_14106);
nand U14649 (N_14649,N_14432,N_14354);
nand U14650 (N_14650,N_14094,N_14206);
and U14651 (N_14651,N_14299,N_14394);
nor U14652 (N_14652,N_14312,N_14135);
or U14653 (N_14653,N_14417,N_14229);
xnor U14654 (N_14654,N_14195,N_14221);
and U14655 (N_14655,N_14324,N_14166);
nand U14656 (N_14656,N_14190,N_14254);
nand U14657 (N_14657,N_14261,N_14477);
and U14658 (N_14658,N_14161,N_14145);
and U14659 (N_14659,N_14034,N_14114);
or U14660 (N_14660,N_14469,N_14410);
xnor U14661 (N_14661,N_14320,N_14475);
and U14662 (N_14662,N_14482,N_14013);
or U14663 (N_14663,N_14054,N_14084);
or U14664 (N_14664,N_14240,N_14117);
xor U14665 (N_14665,N_14120,N_14283);
and U14666 (N_14666,N_14263,N_14192);
nor U14667 (N_14667,N_14284,N_14243);
or U14668 (N_14668,N_14268,N_14021);
xnor U14669 (N_14669,N_14138,N_14285);
nor U14670 (N_14670,N_14495,N_14026);
nor U14671 (N_14671,N_14464,N_14009);
and U14672 (N_14672,N_14378,N_14318);
nor U14673 (N_14673,N_14471,N_14342);
and U14674 (N_14674,N_14260,N_14276);
and U14675 (N_14675,N_14397,N_14390);
nand U14676 (N_14676,N_14235,N_14485);
or U14677 (N_14677,N_14215,N_14301);
nand U14678 (N_14678,N_14377,N_14293);
or U14679 (N_14679,N_14149,N_14450);
and U14680 (N_14680,N_14376,N_14326);
nand U14681 (N_14681,N_14288,N_14216);
nand U14682 (N_14682,N_14055,N_14408);
nand U14683 (N_14683,N_14434,N_14453);
or U14684 (N_14684,N_14303,N_14291);
and U14685 (N_14685,N_14246,N_14357);
and U14686 (N_14686,N_14492,N_14232);
nor U14687 (N_14687,N_14310,N_14133);
nor U14688 (N_14688,N_14363,N_14344);
nand U14689 (N_14689,N_14030,N_14061);
and U14690 (N_14690,N_14065,N_14251);
and U14691 (N_14691,N_14043,N_14109);
or U14692 (N_14692,N_14400,N_14148);
or U14693 (N_14693,N_14351,N_14004);
nand U14694 (N_14694,N_14101,N_14196);
and U14695 (N_14695,N_14270,N_14152);
and U14696 (N_14696,N_14085,N_14414);
or U14697 (N_14697,N_14401,N_14491);
or U14698 (N_14698,N_14060,N_14071);
xnor U14699 (N_14699,N_14058,N_14294);
or U14700 (N_14700,N_14454,N_14317);
and U14701 (N_14701,N_14368,N_14461);
nand U14702 (N_14702,N_14130,N_14467);
xor U14703 (N_14703,N_14418,N_14473);
nand U14704 (N_14704,N_14448,N_14183);
xnor U14705 (N_14705,N_14332,N_14037);
and U14706 (N_14706,N_14199,N_14252);
xor U14707 (N_14707,N_14237,N_14319);
nor U14708 (N_14708,N_14470,N_14140);
nor U14709 (N_14709,N_14356,N_14266);
and U14710 (N_14710,N_14032,N_14024);
nand U14711 (N_14711,N_14444,N_14031);
nor U14712 (N_14712,N_14439,N_14487);
nand U14713 (N_14713,N_14069,N_14040);
xnor U14714 (N_14714,N_14281,N_14249);
nand U14715 (N_14715,N_14204,N_14259);
and U14716 (N_14716,N_14315,N_14269);
nand U14717 (N_14717,N_14188,N_14287);
nor U14718 (N_14718,N_14304,N_14489);
nor U14719 (N_14719,N_14436,N_14264);
nand U14720 (N_14720,N_14331,N_14122);
or U14721 (N_14721,N_14230,N_14219);
nor U14722 (N_14722,N_14115,N_14490);
xor U14723 (N_14723,N_14443,N_14424);
or U14724 (N_14724,N_14273,N_14086);
nand U14725 (N_14725,N_14186,N_14181);
or U14726 (N_14726,N_14258,N_14172);
nand U14727 (N_14727,N_14000,N_14391);
and U14728 (N_14728,N_14121,N_14099);
nand U14729 (N_14729,N_14217,N_14479);
xnor U14730 (N_14730,N_14497,N_14083);
nand U14731 (N_14731,N_14018,N_14290);
or U14732 (N_14732,N_14046,N_14280);
nand U14733 (N_14733,N_14143,N_14220);
xor U14734 (N_14734,N_14180,N_14112);
xnor U14735 (N_14735,N_14039,N_14382);
nand U14736 (N_14736,N_14156,N_14168);
nor U14737 (N_14737,N_14241,N_14113);
or U14738 (N_14738,N_14350,N_14073);
nor U14739 (N_14739,N_14033,N_14088);
nor U14740 (N_14740,N_14366,N_14321);
nand U14741 (N_14741,N_14067,N_14075);
nand U14742 (N_14742,N_14364,N_14468);
nor U14743 (N_14743,N_14423,N_14175);
and U14744 (N_14744,N_14359,N_14238);
xnor U14745 (N_14745,N_14245,N_14435);
and U14746 (N_14746,N_14395,N_14430);
nand U14747 (N_14747,N_14129,N_14355);
nor U14748 (N_14748,N_14095,N_14010);
or U14749 (N_14749,N_14365,N_14316);
or U14750 (N_14750,N_14197,N_14104);
xnor U14751 (N_14751,N_14407,N_14325);
nor U14752 (N_14752,N_14217,N_14193);
and U14753 (N_14753,N_14298,N_14168);
nor U14754 (N_14754,N_14410,N_14039);
nand U14755 (N_14755,N_14395,N_14297);
nand U14756 (N_14756,N_14190,N_14414);
and U14757 (N_14757,N_14393,N_14184);
or U14758 (N_14758,N_14106,N_14432);
xnor U14759 (N_14759,N_14324,N_14126);
and U14760 (N_14760,N_14089,N_14380);
nand U14761 (N_14761,N_14378,N_14014);
or U14762 (N_14762,N_14274,N_14444);
or U14763 (N_14763,N_14144,N_14323);
and U14764 (N_14764,N_14390,N_14349);
xnor U14765 (N_14765,N_14242,N_14255);
or U14766 (N_14766,N_14222,N_14341);
nand U14767 (N_14767,N_14019,N_14287);
and U14768 (N_14768,N_14144,N_14051);
xor U14769 (N_14769,N_14363,N_14045);
and U14770 (N_14770,N_14014,N_14236);
xor U14771 (N_14771,N_14421,N_14494);
nor U14772 (N_14772,N_14420,N_14036);
and U14773 (N_14773,N_14405,N_14029);
xor U14774 (N_14774,N_14096,N_14144);
or U14775 (N_14775,N_14028,N_14031);
and U14776 (N_14776,N_14126,N_14104);
nor U14777 (N_14777,N_14375,N_14148);
xnor U14778 (N_14778,N_14022,N_14444);
and U14779 (N_14779,N_14204,N_14146);
nor U14780 (N_14780,N_14317,N_14044);
nand U14781 (N_14781,N_14394,N_14318);
xor U14782 (N_14782,N_14209,N_14412);
nor U14783 (N_14783,N_14444,N_14277);
nand U14784 (N_14784,N_14243,N_14113);
nand U14785 (N_14785,N_14250,N_14026);
nand U14786 (N_14786,N_14476,N_14019);
nand U14787 (N_14787,N_14441,N_14464);
and U14788 (N_14788,N_14177,N_14106);
nor U14789 (N_14789,N_14106,N_14497);
or U14790 (N_14790,N_14375,N_14068);
or U14791 (N_14791,N_14476,N_14493);
nand U14792 (N_14792,N_14220,N_14185);
and U14793 (N_14793,N_14200,N_14210);
nor U14794 (N_14794,N_14187,N_14351);
or U14795 (N_14795,N_14419,N_14483);
nor U14796 (N_14796,N_14485,N_14166);
or U14797 (N_14797,N_14026,N_14412);
and U14798 (N_14798,N_14191,N_14403);
nor U14799 (N_14799,N_14466,N_14342);
nand U14800 (N_14800,N_14114,N_14200);
nor U14801 (N_14801,N_14365,N_14040);
and U14802 (N_14802,N_14478,N_14159);
or U14803 (N_14803,N_14124,N_14206);
or U14804 (N_14804,N_14456,N_14438);
nand U14805 (N_14805,N_14179,N_14180);
xnor U14806 (N_14806,N_14274,N_14466);
and U14807 (N_14807,N_14476,N_14459);
xor U14808 (N_14808,N_14135,N_14314);
nand U14809 (N_14809,N_14075,N_14463);
and U14810 (N_14810,N_14246,N_14093);
or U14811 (N_14811,N_14090,N_14380);
nor U14812 (N_14812,N_14001,N_14404);
xnor U14813 (N_14813,N_14479,N_14457);
nand U14814 (N_14814,N_14271,N_14428);
nor U14815 (N_14815,N_14423,N_14387);
or U14816 (N_14816,N_14378,N_14248);
and U14817 (N_14817,N_14496,N_14061);
and U14818 (N_14818,N_14245,N_14013);
xnor U14819 (N_14819,N_14491,N_14178);
nand U14820 (N_14820,N_14031,N_14085);
nor U14821 (N_14821,N_14469,N_14449);
nor U14822 (N_14822,N_14167,N_14494);
nor U14823 (N_14823,N_14268,N_14214);
or U14824 (N_14824,N_14483,N_14365);
nor U14825 (N_14825,N_14174,N_14422);
and U14826 (N_14826,N_14382,N_14378);
xor U14827 (N_14827,N_14152,N_14109);
nand U14828 (N_14828,N_14032,N_14482);
xnor U14829 (N_14829,N_14353,N_14054);
nand U14830 (N_14830,N_14194,N_14391);
xor U14831 (N_14831,N_14109,N_14061);
and U14832 (N_14832,N_14282,N_14222);
nand U14833 (N_14833,N_14465,N_14210);
nand U14834 (N_14834,N_14359,N_14083);
xor U14835 (N_14835,N_14384,N_14096);
or U14836 (N_14836,N_14461,N_14082);
or U14837 (N_14837,N_14082,N_14466);
nand U14838 (N_14838,N_14030,N_14083);
nor U14839 (N_14839,N_14106,N_14210);
nor U14840 (N_14840,N_14432,N_14350);
and U14841 (N_14841,N_14169,N_14495);
and U14842 (N_14842,N_14183,N_14331);
and U14843 (N_14843,N_14087,N_14222);
and U14844 (N_14844,N_14347,N_14250);
or U14845 (N_14845,N_14211,N_14409);
nand U14846 (N_14846,N_14425,N_14271);
or U14847 (N_14847,N_14407,N_14143);
nand U14848 (N_14848,N_14062,N_14104);
and U14849 (N_14849,N_14095,N_14470);
nor U14850 (N_14850,N_14239,N_14046);
and U14851 (N_14851,N_14493,N_14498);
nor U14852 (N_14852,N_14460,N_14407);
and U14853 (N_14853,N_14400,N_14377);
or U14854 (N_14854,N_14238,N_14376);
and U14855 (N_14855,N_14185,N_14483);
or U14856 (N_14856,N_14039,N_14254);
and U14857 (N_14857,N_14206,N_14275);
or U14858 (N_14858,N_14457,N_14203);
xor U14859 (N_14859,N_14461,N_14165);
xor U14860 (N_14860,N_14233,N_14131);
nand U14861 (N_14861,N_14357,N_14468);
or U14862 (N_14862,N_14285,N_14053);
and U14863 (N_14863,N_14311,N_14040);
or U14864 (N_14864,N_14371,N_14415);
xor U14865 (N_14865,N_14426,N_14393);
xor U14866 (N_14866,N_14442,N_14379);
and U14867 (N_14867,N_14495,N_14393);
nor U14868 (N_14868,N_14181,N_14348);
nor U14869 (N_14869,N_14403,N_14442);
and U14870 (N_14870,N_14297,N_14210);
and U14871 (N_14871,N_14477,N_14134);
and U14872 (N_14872,N_14034,N_14391);
and U14873 (N_14873,N_14283,N_14076);
nand U14874 (N_14874,N_14290,N_14197);
or U14875 (N_14875,N_14349,N_14050);
nand U14876 (N_14876,N_14130,N_14410);
or U14877 (N_14877,N_14252,N_14450);
and U14878 (N_14878,N_14065,N_14302);
or U14879 (N_14879,N_14162,N_14257);
xor U14880 (N_14880,N_14098,N_14274);
xnor U14881 (N_14881,N_14433,N_14005);
nand U14882 (N_14882,N_14350,N_14365);
or U14883 (N_14883,N_14104,N_14107);
nor U14884 (N_14884,N_14008,N_14217);
nor U14885 (N_14885,N_14371,N_14243);
and U14886 (N_14886,N_14019,N_14135);
nor U14887 (N_14887,N_14260,N_14358);
and U14888 (N_14888,N_14172,N_14370);
nand U14889 (N_14889,N_14198,N_14315);
nor U14890 (N_14890,N_14361,N_14489);
xor U14891 (N_14891,N_14274,N_14199);
nand U14892 (N_14892,N_14072,N_14415);
or U14893 (N_14893,N_14236,N_14345);
and U14894 (N_14894,N_14059,N_14476);
nand U14895 (N_14895,N_14247,N_14417);
xnor U14896 (N_14896,N_14147,N_14361);
and U14897 (N_14897,N_14281,N_14158);
nand U14898 (N_14898,N_14273,N_14471);
xor U14899 (N_14899,N_14163,N_14447);
nor U14900 (N_14900,N_14210,N_14293);
nor U14901 (N_14901,N_14272,N_14075);
and U14902 (N_14902,N_14361,N_14381);
and U14903 (N_14903,N_14444,N_14491);
nand U14904 (N_14904,N_14237,N_14158);
and U14905 (N_14905,N_14298,N_14485);
or U14906 (N_14906,N_14464,N_14081);
nand U14907 (N_14907,N_14087,N_14249);
nor U14908 (N_14908,N_14074,N_14368);
nor U14909 (N_14909,N_14211,N_14210);
nor U14910 (N_14910,N_14177,N_14116);
nand U14911 (N_14911,N_14296,N_14465);
nor U14912 (N_14912,N_14091,N_14272);
nor U14913 (N_14913,N_14054,N_14278);
xor U14914 (N_14914,N_14421,N_14159);
nor U14915 (N_14915,N_14211,N_14215);
nor U14916 (N_14916,N_14276,N_14064);
nor U14917 (N_14917,N_14478,N_14074);
nand U14918 (N_14918,N_14203,N_14079);
nor U14919 (N_14919,N_14129,N_14087);
or U14920 (N_14920,N_14028,N_14098);
nor U14921 (N_14921,N_14210,N_14366);
or U14922 (N_14922,N_14463,N_14074);
xnor U14923 (N_14923,N_14440,N_14256);
and U14924 (N_14924,N_14496,N_14494);
nor U14925 (N_14925,N_14018,N_14394);
nor U14926 (N_14926,N_14475,N_14080);
nand U14927 (N_14927,N_14262,N_14226);
xnor U14928 (N_14928,N_14362,N_14028);
xor U14929 (N_14929,N_14376,N_14438);
and U14930 (N_14930,N_14349,N_14132);
nor U14931 (N_14931,N_14385,N_14077);
and U14932 (N_14932,N_14099,N_14039);
or U14933 (N_14933,N_14299,N_14338);
nand U14934 (N_14934,N_14321,N_14211);
nor U14935 (N_14935,N_14279,N_14041);
xor U14936 (N_14936,N_14176,N_14498);
xor U14937 (N_14937,N_14165,N_14490);
xnor U14938 (N_14938,N_14338,N_14402);
nand U14939 (N_14939,N_14020,N_14024);
or U14940 (N_14940,N_14100,N_14183);
or U14941 (N_14941,N_14190,N_14453);
xor U14942 (N_14942,N_14473,N_14037);
xor U14943 (N_14943,N_14316,N_14145);
and U14944 (N_14944,N_14491,N_14032);
and U14945 (N_14945,N_14228,N_14102);
nand U14946 (N_14946,N_14187,N_14119);
and U14947 (N_14947,N_14368,N_14448);
nor U14948 (N_14948,N_14021,N_14255);
nor U14949 (N_14949,N_14331,N_14141);
xnor U14950 (N_14950,N_14167,N_14364);
nor U14951 (N_14951,N_14369,N_14282);
or U14952 (N_14952,N_14270,N_14029);
nand U14953 (N_14953,N_14230,N_14066);
nor U14954 (N_14954,N_14010,N_14277);
nand U14955 (N_14955,N_14325,N_14269);
xnor U14956 (N_14956,N_14361,N_14188);
and U14957 (N_14957,N_14148,N_14327);
nor U14958 (N_14958,N_14031,N_14027);
nor U14959 (N_14959,N_14346,N_14130);
nand U14960 (N_14960,N_14414,N_14231);
and U14961 (N_14961,N_14157,N_14232);
nor U14962 (N_14962,N_14310,N_14197);
or U14963 (N_14963,N_14047,N_14202);
nand U14964 (N_14964,N_14159,N_14049);
xnor U14965 (N_14965,N_14477,N_14346);
nor U14966 (N_14966,N_14126,N_14391);
xor U14967 (N_14967,N_14434,N_14473);
or U14968 (N_14968,N_14143,N_14285);
and U14969 (N_14969,N_14411,N_14168);
and U14970 (N_14970,N_14068,N_14308);
xor U14971 (N_14971,N_14226,N_14310);
and U14972 (N_14972,N_14369,N_14017);
nor U14973 (N_14973,N_14000,N_14205);
and U14974 (N_14974,N_14089,N_14367);
xnor U14975 (N_14975,N_14330,N_14137);
nand U14976 (N_14976,N_14030,N_14420);
and U14977 (N_14977,N_14401,N_14488);
nor U14978 (N_14978,N_14348,N_14082);
and U14979 (N_14979,N_14105,N_14224);
and U14980 (N_14980,N_14018,N_14434);
and U14981 (N_14981,N_14016,N_14070);
nand U14982 (N_14982,N_14051,N_14192);
and U14983 (N_14983,N_14146,N_14346);
nand U14984 (N_14984,N_14112,N_14138);
and U14985 (N_14985,N_14364,N_14290);
xnor U14986 (N_14986,N_14210,N_14480);
nor U14987 (N_14987,N_14452,N_14059);
and U14988 (N_14988,N_14387,N_14351);
and U14989 (N_14989,N_14155,N_14103);
and U14990 (N_14990,N_14142,N_14342);
nand U14991 (N_14991,N_14424,N_14295);
xnor U14992 (N_14992,N_14478,N_14472);
nor U14993 (N_14993,N_14422,N_14415);
nand U14994 (N_14994,N_14480,N_14253);
or U14995 (N_14995,N_14494,N_14417);
and U14996 (N_14996,N_14485,N_14014);
and U14997 (N_14997,N_14257,N_14237);
nor U14998 (N_14998,N_14041,N_14241);
nor U14999 (N_14999,N_14450,N_14456);
xnor U15000 (N_15000,N_14942,N_14982);
nor U15001 (N_15001,N_14936,N_14823);
nor U15002 (N_15002,N_14712,N_14891);
nand U15003 (N_15003,N_14993,N_14553);
nor U15004 (N_15004,N_14659,N_14690);
and U15005 (N_15005,N_14632,N_14846);
nor U15006 (N_15006,N_14839,N_14827);
xnor U15007 (N_15007,N_14603,N_14835);
xor U15008 (N_15008,N_14888,N_14913);
or U15009 (N_15009,N_14918,N_14604);
and U15010 (N_15010,N_14554,N_14564);
or U15011 (N_15011,N_14962,N_14524);
xnor U15012 (N_15012,N_14831,N_14565);
nand U15013 (N_15013,N_14915,N_14987);
or U15014 (N_15014,N_14645,N_14613);
or U15015 (N_15015,N_14621,N_14601);
or U15016 (N_15016,N_14841,N_14507);
nor U15017 (N_15017,N_14964,N_14711);
nand U15018 (N_15018,N_14568,N_14671);
xnor U15019 (N_15019,N_14676,N_14515);
xor U15020 (N_15020,N_14658,N_14505);
and U15021 (N_15021,N_14673,N_14630);
and U15022 (N_15022,N_14984,N_14956);
nor U15023 (N_15023,N_14559,N_14876);
or U15024 (N_15024,N_14957,N_14769);
or U15025 (N_15025,N_14895,N_14502);
or U15026 (N_15026,N_14781,N_14725);
and U15027 (N_15027,N_14715,N_14561);
nor U15028 (N_15028,N_14872,N_14926);
nand U15029 (N_15029,N_14900,N_14910);
xnor U15030 (N_15030,N_14871,N_14723);
nor U15031 (N_15031,N_14751,N_14950);
or U15032 (N_15032,N_14503,N_14695);
nand U15033 (N_15033,N_14892,N_14633);
and U15034 (N_15034,N_14612,N_14593);
xor U15035 (N_15035,N_14579,N_14834);
nand U15036 (N_15036,N_14665,N_14698);
xor U15037 (N_15037,N_14865,N_14727);
nor U15038 (N_15038,N_14909,N_14605);
nand U15039 (N_15039,N_14762,N_14506);
nor U15040 (N_15040,N_14704,N_14517);
nand U15041 (N_15041,N_14634,N_14577);
nor U15042 (N_15042,N_14618,N_14560);
xor U15043 (N_15043,N_14741,N_14851);
and U15044 (N_15044,N_14920,N_14819);
nand U15045 (N_15045,N_14528,N_14792);
or U15046 (N_15046,N_14784,N_14951);
and U15047 (N_15047,N_14525,N_14804);
nand U15048 (N_15048,N_14991,N_14664);
xnor U15049 (N_15049,N_14687,N_14575);
nand U15050 (N_15050,N_14948,N_14759);
and U15051 (N_15051,N_14666,N_14663);
or U15052 (N_15052,N_14754,N_14767);
nand U15053 (N_15053,N_14939,N_14952);
nand U15054 (N_15054,N_14521,N_14642);
or U15055 (N_15055,N_14898,N_14821);
or U15056 (N_15056,N_14945,N_14735);
nor U15057 (N_15057,N_14897,N_14683);
nor U15058 (N_15058,N_14961,N_14674);
nor U15059 (N_15059,N_14944,N_14739);
and U15060 (N_15060,N_14861,N_14679);
nor U15061 (N_15061,N_14975,N_14999);
or U15062 (N_15062,N_14534,N_14787);
or U15063 (N_15063,N_14662,N_14989);
nand U15064 (N_15064,N_14855,N_14550);
nor U15065 (N_15065,N_14903,N_14894);
xnor U15066 (N_15066,N_14817,N_14627);
nor U15067 (N_15067,N_14914,N_14636);
or U15068 (N_15068,N_14800,N_14607);
or U15069 (N_15069,N_14513,N_14919);
or U15070 (N_15070,N_14598,N_14746);
xnor U15071 (N_15071,N_14996,N_14809);
nand U15072 (N_15072,N_14551,N_14978);
nand U15073 (N_15073,N_14748,N_14912);
nand U15074 (N_15074,N_14668,N_14925);
and U15075 (N_15075,N_14907,N_14937);
nand U15076 (N_15076,N_14816,N_14829);
xnor U15077 (N_15077,N_14790,N_14705);
nor U15078 (N_15078,N_14845,N_14563);
or U15079 (N_15079,N_14558,N_14686);
xor U15080 (N_15080,N_14721,N_14752);
and U15081 (N_15081,N_14765,N_14611);
nand U15082 (N_15082,N_14775,N_14976);
nor U15083 (N_15083,N_14610,N_14637);
nand U15084 (N_15084,N_14796,N_14998);
nor U15085 (N_15085,N_14880,N_14701);
xor U15086 (N_15086,N_14896,N_14955);
or U15087 (N_15087,N_14737,N_14713);
nand U15088 (N_15088,N_14539,N_14847);
or U15089 (N_15089,N_14931,N_14660);
and U15090 (N_15090,N_14772,N_14814);
and U15091 (N_15091,N_14875,N_14706);
and U15092 (N_15092,N_14818,N_14902);
or U15093 (N_15093,N_14828,N_14731);
or U15094 (N_15094,N_14904,N_14968);
or U15095 (N_15095,N_14549,N_14771);
or U15096 (N_15096,N_14794,N_14667);
and U15097 (N_15097,N_14670,N_14868);
and U15098 (N_15098,N_14863,N_14608);
xnor U15099 (N_15099,N_14609,N_14960);
nand U15100 (N_15100,N_14661,N_14578);
and U15101 (N_15101,N_14867,N_14647);
nand U15102 (N_15102,N_14520,N_14877);
nor U15103 (N_15103,N_14805,N_14720);
and U15104 (N_15104,N_14570,N_14548);
xnor U15105 (N_15105,N_14724,N_14890);
nor U15106 (N_15106,N_14714,N_14718);
nor U15107 (N_15107,N_14783,N_14722);
nor U15108 (N_15108,N_14908,N_14531);
nor U15109 (N_15109,N_14820,N_14807);
nor U15110 (N_15110,N_14932,N_14826);
nor U15111 (N_15111,N_14921,N_14592);
xor U15112 (N_15112,N_14789,N_14512);
nand U15113 (N_15113,N_14617,N_14822);
xnor U15114 (N_15114,N_14806,N_14878);
nor U15115 (N_15115,N_14730,N_14833);
nand U15116 (N_15116,N_14614,N_14791);
xnor U15117 (N_15117,N_14940,N_14750);
nor U15118 (N_15118,N_14646,N_14916);
nand U15119 (N_15119,N_14547,N_14911);
xor U15120 (N_15120,N_14744,N_14747);
and U15121 (N_15121,N_14699,N_14963);
xnor U15122 (N_15122,N_14859,N_14793);
and U15123 (N_15123,N_14626,N_14858);
xnor U15124 (N_15124,N_14774,N_14717);
xnor U15125 (N_15125,N_14591,N_14696);
xor U15126 (N_15126,N_14749,N_14555);
nor U15127 (N_15127,N_14700,N_14588);
nor U15128 (N_15128,N_14743,N_14523);
and U15129 (N_15129,N_14997,N_14967);
nor U15130 (N_15130,N_14905,N_14813);
nand U15131 (N_15131,N_14873,N_14654);
xor U15132 (N_15132,N_14803,N_14732);
xnor U15133 (N_15133,N_14947,N_14596);
or U15134 (N_15134,N_14682,N_14799);
nand U15135 (N_15135,N_14538,N_14753);
and U15136 (N_15136,N_14980,N_14795);
or U15137 (N_15137,N_14546,N_14651);
xor U15138 (N_15138,N_14934,N_14677);
nor U15139 (N_15139,N_14842,N_14639);
or U15140 (N_15140,N_14641,N_14622);
xor U15141 (N_15141,N_14756,N_14776);
xnor U15142 (N_15142,N_14536,N_14624);
nand U15143 (N_15143,N_14930,N_14586);
nand U15144 (N_15144,N_14979,N_14572);
nand U15145 (N_15145,N_14556,N_14879);
nor U15146 (N_15146,N_14869,N_14562);
nand U15147 (N_15147,N_14620,N_14901);
nand U15148 (N_15148,N_14681,N_14599);
nor U15149 (N_15149,N_14526,N_14552);
and U15150 (N_15150,N_14519,N_14619);
or U15151 (N_15151,N_14689,N_14537);
or U15152 (N_15152,N_14511,N_14943);
and U15153 (N_15153,N_14848,N_14927);
or U15154 (N_15154,N_14606,N_14832);
xor U15155 (N_15155,N_14889,N_14972);
xor U15156 (N_15156,N_14837,N_14881);
or U15157 (N_15157,N_14985,N_14992);
and U15158 (N_15158,N_14786,N_14929);
xor U15159 (N_15159,N_14535,N_14779);
nor U15160 (N_15160,N_14516,N_14815);
or U15161 (N_15161,N_14583,N_14567);
xor U15162 (N_15162,N_14856,N_14542);
or U15163 (N_15163,N_14691,N_14981);
nor U15164 (N_15164,N_14514,N_14740);
or U15165 (N_15165,N_14885,N_14933);
xnor U15166 (N_15166,N_14569,N_14571);
nor U15167 (N_15167,N_14798,N_14703);
and U15168 (N_15168,N_14785,N_14849);
xnor U15169 (N_15169,N_14709,N_14649);
or U15170 (N_15170,N_14693,N_14953);
xor U15171 (N_15171,N_14778,N_14625);
or U15172 (N_15172,N_14958,N_14576);
nand U15173 (N_15173,N_14760,N_14893);
nor U15174 (N_15174,N_14600,N_14640);
and U15175 (N_15175,N_14580,N_14938);
and U15176 (N_15176,N_14616,N_14504);
nor U15177 (N_15177,N_14527,N_14986);
nor U15178 (N_15178,N_14518,N_14811);
and U15179 (N_15179,N_14917,N_14540);
or U15180 (N_15180,N_14684,N_14899);
nor U15181 (N_15181,N_14678,N_14923);
or U15182 (N_15182,N_14812,N_14860);
and U15183 (N_15183,N_14850,N_14782);
nor U15184 (N_15184,N_14761,N_14707);
and U15185 (N_15185,N_14946,N_14702);
xnor U15186 (N_15186,N_14742,N_14764);
or U15187 (N_15187,N_14949,N_14655);
nand U15188 (N_15188,N_14648,N_14589);
nand U15189 (N_15189,N_14853,N_14597);
or U15190 (N_15190,N_14862,N_14728);
or U15191 (N_15191,N_14770,N_14797);
or U15192 (N_15192,N_14988,N_14510);
nand U15193 (N_15193,N_14595,N_14854);
and U15194 (N_15194,N_14594,N_14602);
nand U15195 (N_15195,N_14808,N_14716);
nand U15196 (N_15196,N_14810,N_14763);
nor U15197 (N_15197,N_14644,N_14965);
xnor U15198 (N_15198,N_14969,N_14843);
nand U15199 (N_15199,N_14631,N_14864);
or U15200 (N_15200,N_14587,N_14685);
or U15201 (N_15201,N_14543,N_14973);
xnor U15202 (N_15202,N_14830,N_14755);
or U15203 (N_15203,N_14638,N_14657);
and U15204 (N_15204,N_14887,N_14736);
or U15205 (N_15205,N_14941,N_14557);
nand U15206 (N_15206,N_14585,N_14874);
nand U15207 (N_15207,N_14780,N_14582);
nor U15208 (N_15208,N_14710,N_14733);
or U15209 (N_15209,N_14694,N_14669);
or U15210 (N_15210,N_14533,N_14758);
nand U15211 (N_15211,N_14726,N_14688);
xnor U15212 (N_15212,N_14844,N_14882);
nor U15213 (N_15213,N_14971,N_14970);
nor U15214 (N_15214,N_14824,N_14773);
and U15215 (N_15215,N_14734,N_14501);
or U15216 (N_15216,N_14836,N_14522);
nand U15217 (N_15217,N_14672,N_14857);
nor U15218 (N_15218,N_14544,N_14990);
nor U15219 (N_15219,N_14697,N_14777);
nor U15220 (N_15220,N_14825,N_14532);
xor U15221 (N_15221,N_14906,N_14866);
nand U15222 (N_15222,N_14883,N_14768);
or U15223 (N_15223,N_14788,N_14623);
xor U15224 (N_15224,N_14653,N_14574);
nand U15225 (N_15225,N_14922,N_14545);
xnor U15226 (N_15226,N_14635,N_14954);
nand U15227 (N_15227,N_14615,N_14708);
nand U15228 (N_15228,N_14870,N_14508);
nor U15229 (N_15229,N_14692,N_14959);
nand U15230 (N_15230,N_14643,N_14566);
nor U15231 (N_15231,N_14573,N_14529);
nand U15232 (N_15232,N_14738,N_14994);
and U15233 (N_15233,N_14966,N_14983);
nor U15234 (N_15234,N_14928,N_14650);
or U15235 (N_15235,N_14924,N_14766);
and U15236 (N_15236,N_14852,N_14838);
nand U15237 (N_15237,N_14840,N_14719);
or U15238 (N_15238,N_14581,N_14680);
nor U15239 (N_15239,N_14509,N_14884);
or U15240 (N_15240,N_14974,N_14530);
and U15241 (N_15241,N_14675,N_14628);
nor U15242 (N_15242,N_14541,N_14629);
xor U15243 (N_15243,N_14801,N_14995);
and U15244 (N_15244,N_14500,N_14729);
nand U15245 (N_15245,N_14802,N_14652);
nor U15246 (N_15246,N_14656,N_14590);
or U15247 (N_15247,N_14745,N_14977);
and U15248 (N_15248,N_14886,N_14757);
or U15249 (N_15249,N_14584,N_14935);
xnor U15250 (N_15250,N_14808,N_14981);
or U15251 (N_15251,N_14703,N_14866);
nor U15252 (N_15252,N_14978,N_14573);
nand U15253 (N_15253,N_14587,N_14816);
and U15254 (N_15254,N_14886,N_14632);
xor U15255 (N_15255,N_14760,N_14572);
nand U15256 (N_15256,N_14809,N_14693);
and U15257 (N_15257,N_14748,N_14714);
nor U15258 (N_15258,N_14673,N_14796);
nand U15259 (N_15259,N_14598,N_14838);
and U15260 (N_15260,N_14678,N_14662);
and U15261 (N_15261,N_14915,N_14684);
and U15262 (N_15262,N_14861,N_14953);
xnor U15263 (N_15263,N_14732,N_14999);
nor U15264 (N_15264,N_14854,N_14632);
nand U15265 (N_15265,N_14704,N_14614);
and U15266 (N_15266,N_14656,N_14511);
nand U15267 (N_15267,N_14827,N_14724);
and U15268 (N_15268,N_14623,N_14985);
nand U15269 (N_15269,N_14904,N_14950);
xnor U15270 (N_15270,N_14717,N_14746);
nor U15271 (N_15271,N_14988,N_14657);
or U15272 (N_15272,N_14679,N_14609);
xnor U15273 (N_15273,N_14549,N_14631);
nor U15274 (N_15274,N_14909,N_14785);
or U15275 (N_15275,N_14925,N_14534);
nor U15276 (N_15276,N_14526,N_14944);
nand U15277 (N_15277,N_14754,N_14969);
or U15278 (N_15278,N_14874,N_14875);
nand U15279 (N_15279,N_14775,N_14585);
or U15280 (N_15280,N_14890,N_14945);
nor U15281 (N_15281,N_14528,N_14743);
nand U15282 (N_15282,N_14649,N_14990);
and U15283 (N_15283,N_14755,N_14899);
nand U15284 (N_15284,N_14799,N_14699);
xor U15285 (N_15285,N_14675,N_14770);
nand U15286 (N_15286,N_14778,N_14772);
and U15287 (N_15287,N_14933,N_14684);
or U15288 (N_15288,N_14901,N_14859);
nor U15289 (N_15289,N_14568,N_14586);
xnor U15290 (N_15290,N_14899,N_14982);
nor U15291 (N_15291,N_14578,N_14973);
nand U15292 (N_15292,N_14568,N_14953);
and U15293 (N_15293,N_14951,N_14979);
or U15294 (N_15294,N_14601,N_14757);
and U15295 (N_15295,N_14595,N_14763);
or U15296 (N_15296,N_14584,N_14571);
xor U15297 (N_15297,N_14525,N_14740);
nand U15298 (N_15298,N_14596,N_14546);
or U15299 (N_15299,N_14710,N_14611);
or U15300 (N_15300,N_14761,N_14929);
nand U15301 (N_15301,N_14543,N_14536);
or U15302 (N_15302,N_14623,N_14699);
and U15303 (N_15303,N_14979,N_14815);
nand U15304 (N_15304,N_14752,N_14590);
and U15305 (N_15305,N_14726,N_14738);
nor U15306 (N_15306,N_14870,N_14861);
nand U15307 (N_15307,N_14532,N_14707);
nor U15308 (N_15308,N_14968,N_14909);
and U15309 (N_15309,N_14964,N_14651);
or U15310 (N_15310,N_14527,N_14512);
or U15311 (N_15311,N_14938,N_14511);
nor U15312 (N_15312,N_14835,N_14516);
nor U15313 (N_15313,N_14995,N_14523);
or U15314 (N_15314,N_14640,N_14576);
and U15315 (N_15315,N_14513,N_14591);
nor U15316 (N_15316,N_14859,N_14891);
or U15317 (N_15317,N_14550,N_14864);
xnor U15318 (N_15318,N_14702,N_14658);
nand U15319 (N_15319,N_14992,N_14982);
nor U15320 (N_15320,N_14863,N_14753);
and U15321 (N_15321,N_14779,N_14533);
or U15322 (N_15322,N_14637,N_14706);
nor U15323 (N_15323,N_14714,N_14865);
and U15324 (N_15324,N_14652,N_14702);
and U15325 (N_15325,N_14549,N_14925);
nand U15326 (N_15326,N_14812,N_14548);
and U15327 (N_15327,N_14615,N_14528);
nand U15328 (N_15328,N_14760,N_14535);
nand U15329 (N_15329,N_14534,N_14996);
nor U15330 (N_15330,N_14777,N_14765);
or U15331 (N_15331,N_14848,N_14894);
and U15332 (N_15332,N_14574,N_14740);
nor U15333 (N_15333,N_14689,N_14679);
xnor U15334 (N_15334,N_14822,N_14636);
nor U15335 (N_15335,N_14639,N_14684);
xor U15336 (N_15336,N_14918,N_14984);
xnor U15337 (N_15337,N_14840,N_14980);
xor U15338 (N_15338,N_14582,N_14811);
xor U15339 (N_15339,N_14854,N_14975);
nand U15340 (N_15340,N_14739,N_14721);
xor U15341 (N_15341,N_14562,N_14508);
and U15342 (N_15342,N_14909,N_14832);
nor U15343 (N_15343,N_14995,N_14613);
xor U15344 (N_15344,N_14930,N_14731);
nand U15345 (N_15345,N_14893,N_14618);
or U15346 (N_15346,N_14922,N_14920);
nor U15347 (N_15347,N_14702,N_14814);
or U15348 (N_15348,N_14626,N_14896);
nand U15349 (N_15349,N_14923,N_14696);
nand U15350 (N_15350,N_14621,N_14840);
nor U15351 (N_15351,N_14835,N_14520);
or U15352 (N_15352,N_14695,N_14586);
or U15353 (N_15353,N_14620,N_14618);
nor U15354 (N_15354,N_14856,N_14623);
nand U15355 (N_15355,N_14519,N_14917);
or U15356 (N_15356,N_14745,N_14784);
nor U15357 (N_15357,N_14921,N_14718);
nand U15358 (N_15358,N_14621,N_14986);
or U15359 (N_15359,N_14622,N_14756);
or U15360 (N_15360,N_14656,N_14824);
and U15361 (N_15361,N_14802,N_14544);
or U15362 (N_15362,N_14973,N_14535);
nor U15363 (N_15363,N_14888,N_14739);
nand U15364 (N_15364,N_14844,N_14842);
nand U15365 (N_15365,N_14908,N_14791);
and U15366 (N_15366,N_14943,N_14676);
xnor U15367 (N_15367,N_14513,N_14945);
or U15368 (N_15368,N_14615,N_14955);
xnor U15369 (N_15369,N_14907,N_14686);
nor U15370 (N_15370,N_14600,N_14728);
nor U15371 (N_15371,N_14944,N_14885);
xnor U15372 (N_15372,N_14784,N_14597);
nor U15373 (N_15373,N_14847,N_14980);
nor U15374 (N_15374,N_14844,N_14561);
nor U15375 (N_15375,N_14918,N_14798);
or U15376 (N_15376,N_14844,N_14992);
and U15377 (N_15377,N_14571,N_14941);
or U15378 (N_15378,N_14512,N_14654);
nor U15379 (N_15379,N_14701,N_14634);
or U15380 (N_15380,N_14864,N_14647);
xor U15381 (N_15381,N_14677,N_14923);
and U15382 (N_15382,N_14512,N_14826);
or U15383 (N_15383,N_14907,N_14627);
and U15384 (N_15384,N_14937,N_14668);
or U15385 (N_15385,N_14853,N_14955);
xor U15386 (N_15386,N_14940,N_14558);
and U15387 (N_15387,N_14667,N_14860);
nor U15388 (N_15388,N_14705,N_14800);
and U15389 (N_15389,N_14612,N_14722);
nor U15390 (N_15390,N_14518,N_14848);
xor U15391 (N_15391,N_14934,N_14662);
nand U15392 (N_15392,N_14858,N_14607);
nand U15393 (N_15393,N_14896,N_14640);
nor U15394 (N_15394,N_14573,N_14641);
or U15395 (N_15395,N_14523,N_14563);
and U15396 (N_15396,N_14799,N_14782);
nor U15397 (N_15397,N_14664,N_14673);
nand U15398 (N_15398,N_14716,N_14816);
or U15399 (N_15399,N_14879,N_14559);
nor U15400 (N_15400,N_14844,N_14607);
xor U15401 (N_15401,N_14527,N_14989);
or U15402 (N_15402,N_14977,N_14936);
xnor U15403 (N_15403,N_14965,N_14819);
or U15404 (N_15404,N_14900,N_14827);
nand U15405 (N_15405,N_14651,N_14785);
xnor U15406 (N_15406,N_14900,N_14742);
nand U15407 (N_15407,N_14672,N_14754);
nand U15408 (N_15408,N_14515,N_14879);
xor U15409 (N_15409,N_14610,N_14674);
nor U15410 (N_15410,N_14749,N_14914);
or U15411 (N_15411,N_14512,N_14683);
nand U15412 (N_15412,N_14911,N_14746);
and U15413 (N_15413,N_14811,N_14640);
and U15414 (N_15414,N_14584,N_14662);
nor U15415 (N_15415,N_14995,N_14533);
or U15416 (N_15416,N_14683,N_14694);
or U15417 (N_15417,N_14797,N_14858);
and U15418 (N_15418,N_14688,N_14945);
xor U15419 (N_15419,N_14975,N_14950);
or U15420 (N_15420,N_14561,N_14900);
nand U15421 (N_15421,N_14809,N_14531);
or U15422 (N_15422,N_14916,N_14932);
or U15423 (N_15423,N_14623,N_14937);
or U15424 (N_15424,N_14559,N_14564);
nand U15425 (N_15425,N_14689,N_14631);
nand U15426 (N_15426,N_14642,N_14547);
and U15427 (N_15427,N_14827,N_14606);
nor U15428 (N_15428,N_14848,N_14542);
xor U15429 (N_15429,N_14566,N_14844);
nand U15430 (N_15430,N_14671,N_14543);
or U15431 (N_15431,N_14885,N_14920);
nor U15432 (N_15432,N_14988,N_14887);
xnor U15433 (N_15433,N_14737,N_14592);
xor U15434 (N_15434,N_14661,N_14946);
xor U15435 (N_15435,N_14955,N_14905);
nand U15436 (N_15436,N_14811,N_14787);
xnor U15437 (N_15437,N_14652,N_14977);
or U15438 (N_15438,N_14760,N_14739);
xor U15439 (N_15439,N_14605,N_14896);
nand U15440 (N_15440,N_14569,N_14874);
and U15441 (N_15441,N_14713,N_14991);
nand U15442 (N_15442,N_14978,N_14684);
and U15443 (N_15443,N_14560,N_14775);
xnor U15444 (N_15444,N_14822,N_14930);
nor U15445 (N_15445,N_14923,N_14739);
xnor U15446 (N_15446,N_14715,N_14853);
xnor U15447 (N_15447,N_14891,N_14885);
nand U15448 (N_15448,N_14921,N_14851);
xor U15449 (N_15449,N_14784,N_14720);
or U15450 (N_15450,N_14672,N_14832);
and U15451 (N_15451,N_14786,N_14818);
nand U15452 (N_15452,N_14737,N_14760);
nor U15453 (N_15453,N_14869,N_14956);
and U15454 (N_15454,N_14726,N_14598);
nor U15455 (N_15455,N_14745,N_14623);
nand U15456 (N_15456,N_14733,N_14514);
xor U15457 (N_15457,N_14839,N_14826);
or U15458 (N_15458,N_14953,N_14902);
xor U15459 (N_15459,N_14648,N_14546);
and U15460 (N_15460,N_14528,N_14852);
xnor U15461 (N_15461,N_14542,N_14573);
nor U15462 (N_15462,N_14688,N_14970);
and U15463 (N_15463,N_14842,N_14987);
nand U15464 (N_15464,N_14815,N_14772);
or U15465 (N_15465,N_14734,N_14698);
nor U15466 (N_15466,N_14669,N_14717);
nand U15467 (N_15467,N_14584,N_14936);
xor U15468 (N_15468,N_14705,N_14516);
or U15469 (N_15469,N_14837,N_14657);
and U15470 (N_15470,N_14879,N_14725);
or U15471 (N_15471,N_14799,N_14648);
xnor U15472 (N_15472,N_14986,N_14550);
nor U15473 (N_15473,N_14930,N_14518);
xnor U15474 (N_15474,N_14728,N_14546);
nand U15475 (N_15475,N_14943,N_14959);
nor U15476 (N_15476,N_14930,N_14932);
nand U15477 (N_15477,N_14767,N_14565);
and U15478 (N_15478,N_14727,N_14729);
or U15479 (N_15479,N_14677,N_14760);
nand U15480 (N_15480,N_14923,N_14825);
nor U15481 (N_15481,N_14682,N_14629);
nor U15482 (N_15482,N_14693,N_14815);
nand U15483 (N_15483,N_14917,N_14812);
or U15484 (N_15484,N_14692,N_14930);
and U15485 (N_15485,N_14936,N_14821);
nand U15486 (N_15486,N_14555,N_14550);
nand U15487 (N_15487,N_14502,N_14500);
or U15488 (N_15488,N_14937,N_14574);
or U15489 (N_15489,N_14787,N_14945);
nand U15490 (N_15490,N_14755,N_14798);
or U15491 (N_15491,N_14639,N_14933);
nor U15492 (N_15492,N_14876,N_14671);
nor U15493 (N_15493,N_14962,N_14654);
nand U15494 (N_15494,N_14958,N_14858);
and U15495 (N_15495,N_14663,N_14988);
and U15496 (N_15496,N_14722,N_14672);
xor U15497 (N_15497,N_14993,N_14968);
or U15498 (N_15498,N_14777,N_14622);
or U15499 (N_15499,N_14593,N_14619);
xnor U15500 (N_15500,N_15140,N_15429);
nand U15501 (N_15501,N_15130,N_15408);
or U15502 (N_15502,N_15092,N_15494);
nand U15503 (N_15503,N_15045,N_15451);
nor U15504 (N_15504,N_15264,N_15276);
and U15505 (N_15505,N_15129,N_15213);
and U15506 (N_15506,N_15031,N_15118);
or U15507 (N_15507,N_15392,N_15255);
and U15508 (N_15508,N_15176,N_15001);
or U15509 (N_15509,N_15158,N_15268);
nor U15510 (N_15510,N_15230,N_15220);
and U15511 (N_15511,N_15362,N_15063);
nor U15512 (N_15512,N_15409,N_15047);
or U15513 (N_15513,N_15361,N_15443);
or U15514 (N_15514,N_15175,N_15330);
xnor U15515 (N_15515,N_15208,N_15271);
xnor U15516 (N_15516,N_15126,N_15036);
xnor U15517 (N_15517,N_15133,N_15394);
nand U15518 (N_15518,N_15046,N_15337);
or U15519 (N_15519,N_15114,N_15439);
nand U15520 (N_15520,N_15436,N_15009);
xnor U15521 (N_15521,N_15037,N_15192);
nor U15522 (N_15522,N_15059,N_15442);
nor U15523 (N_15523,N_15180,N_15177);
or U15524 (N_15524,N_15101,N_15084);
nand U15525 (N_15525,N_15363,N_15194);
xor U15526 (N_15526,N_15300,N_15316);
or U15527 (N_15527,N_15259,N_15309);
or U15528 (N_15528,N_15313,N_15042);
nand U15529 (N_15529,N_15106,N_15139);
nand U15530 (N_15530,N_15326,N_15079);
and U15531 (N_15531,N_15496,N_15007);
nor U15532 (N_15532,N_15413,N_15170);
or U15533 (N_15533,N_15102,N_15141);
nand U15534 (N_15534,N_15017,N_15228);
nor U15535 (N_15535,N_15488,N_15367);
nand U15536 (N_15536,N_15098,N_15399);
nand U15537 (N_15537,N_15277,N_15446);
or U15538 (N_15538,N_15467,N_15146);
xor U15539 (N_15539,N_15317,N_15174);
and U15540 (N_15540,N_15324,N_15088);
nand U15541 (N_15541,N_15152,N_15297);
and U15542 (N_15542,N_15186,N_15293);
or U15543 (N_15543,N_15061,N_15252);
xor U15544 (N_15544,N_15280,N_15191);
and U15545 (N_15545,N_15035,N_15380);
xnor U15546 (N_15546,N_15469,N_15193);
nor U15547 (N_15547,N_15331,N_15103);
or U15548 (N_15548,N_15159,N_15357);
and U15549 (N_15549,N_15072,N_15403);
and U15550 (N_15550,N_15188,N_15232);
nand U15551 (N_15551,N_15085,N_15342);
and U15552 (N_15552,N_15241,N_15110);
nand U15553 (N_15553,N_15325,N_15049);
and U15554 (N_15554,N_15381,N_15263);
nand U15555 (N_15555,N_15097,N_15348);
nand U15556 (N_15556,N_15181,N_15395);
and U15557 (N_15557,N_15299,N_15265);
xnor U15558 (N_15558,N_15183,N_15428);
xnor U15559 (N_15559,N_15267,N_15308);
xor U15560 (N_15560,N_15044,N_15425);
xor U15561 (N_15561,N_15025,N_15447);
and U15562 (N_15562,N_15053,N_15303);
nor U15563 (N_15563,N_15206,N_15444);
nand U15564 (N_15564,N_15421,N_15195);
xnor U15565 (N_15565,N_15334,N_15080);
nor U15566 (N_15566,N_15209,N_15014);
xnor U15567 (N_15567,N_15369,N_15090);
nand U15568 (N_15568,N_15167,N_15078);
nand U15569 (N_15569,N_15026,N_15246);
nand U15570 (N_15570,N_15462,N_15423);
nand U15571 (N_15571,N_15360,N_15430);
nor U15572 (N_15572,N_15284,N_15003);
xnor U15573 (N_15573,N_15131,N_15273);
xor U15574 (N_15574,N_15449,N_15144);
xor U15575 (N_15575,N_15163,N_15125);
xnor U15576 (N_15576,N_15082,N_15002);
nand U15577 (N_15577,N_15005,N_15269);
and U15578 (N_15578,N_15455,N_15022);
nand U15579 (N_15579,N_15134,N_15214);
or U15580 (N_15580,N_15116,N_15450);
nor U15581 (N_15581,N_15288,N_15073);
or U15582 (N_15582,N_15379,N_15096);
xnor U15583 (N_15583,N_15456,N_15388);
or U15584 (N_15584,N_15201,N_15472);
or U15585 (N_15585,N_15405,N_15328);
and U15586 (N_15586,N_15477,N_15240);
or U15587 (N_15587,N_15081,N_15157);
nand U15588 (N_15588,N_15233,N_15242);
or U15589 (N_15589,N_15249,N_15190);
nor U15590 (N_15590,N_15067,N_15060);
and U15591 (N_15591,N_15011,N_15172);
nand U15592 (N_15592,N_15312,N_15321);
or U15593 (N_15593,N_15283,N_15262);
or U15594 (N_15594,N_15437,N_15480);
or U15595 (N_15595,N_15121,N_15296);
or U15596 (N_15596,N_15153,N_15327);
and U15597 (N_15597,N_15256,N_15484);
nand U15598 (N_15598,N_15371,N_15030);
xor U15599 (N_15599,N_15458,N_15016);
xor U15600 (N_15600,N_15499,N_15120);
nor U15601 (N_15601,N_15020,N_15278);
or U15602 (N_15602,N_15266,N_15132);
nand U15603 (N_15603,N_15113,N_15389);
or U15604 (N_15604,N_15124,N_15064);
nand U15605 (N_15605,N_15295,N_15332);
nand U15606 (N_15606,N_15204,N_15459);
nor U15607 (N_15607,N_15358,N_15223);
nand U15608 (N_15608,N_15401,N_15086);
xor U15609 (N_15609,N_15353,N_15162);
xor U15610 (N_15610,N_15178,N_15419);
or U15611 (N_15611,N_15471,N_15225);
xnor U15612 (N_15612,N_15111,N_15048);
nand U15613 (N_15613,N_15479,N_15311);
or U15614 (N_15614,N_15032,N_15136);
nand U15615 (N_15615,N_15491,N_15010);
nor U15616 (N_15616,N_15200,N_15226);
or U15617 (N_15617,N_15122,N_15235);
or U15618 (N_15618,N_15473,N_15245);
xnor U15619 (N_15619,N_15107,N_15013);
xor U15620 (N_15620,N_15282,N_15169);
nand U15621 (N_15621,N_15094,N_15237);
nand U15622 (N_15622,N_15258,N_15340);
or U15623 (N_15623,N_15427,N_15221);
and U15624 (N_15624,N_15222,N_15274);
xnor U15625 (N_15625,N_15386,N_15154);
nor U15626 (N_15626,N_15057,N_15410);
and U15627 (N_15627,N_15123,N_15234);
and U15628 (N_15628,N_15215,N_15091);
nand U15629 (N_15629,N_15149,N_15108);
nor U15630 (N_15630,N_15292,N_15100);
and U15631 (N_15631,N_15257,N_15341);
xnor U15632 (N_15632,N_15093,N_15095);
nand U15633 (N_15633,N_15375,N_15441);
and U15634 (N_15634,N_15117,N_15187);
xor U15635 (N_15635,N_15171,N_15355);
or U15636 (N_15636,N_15272,N_15468);
or U15637 (N_15637,N_15483,N_15112);
and U15638 (N_15638,N_15104,N_15412);
and U15639 (N_15639,N_15454,N_15376);
nand U15640 (N_15640,N_15414,N_15485);
nand U15641 (N_15641,N_15416,N_15127);
nand U15642 (N_15642,N_15071,N_15138);
nor U15643 (N_15643,N_15004,N_15055);
nor U15644 (N_15644,N_15145,N_15012);
nor U15645 (N_15645,N_15453,N_15099);
or U15646 (N_15646,N_15075,N_15404);
and U15647 (N_15647,N_15493,N_15445);
and U15648 (N_15648,N_15433,N_15420);
nor U15649 (N_15649,N_15343,N_15089);
nand U15650 (N_15650,N_15398,N_15281);
or U15651 (N_15651,N_15474,N_15142);
xor U15652 (N_15652,N_15290,N_15260);
xnor U15653 (N_15653,N_15418,N_15038);
nor U15654 (N_15654,N_15393,N_15054);
or U15655 (N_15655,N_15440,N_15155);
and U15656 (N_15656,N_15000,N_15087);
nor U15657 (N_15657,N_15147,N_15066);
or U15658 (N_15658,N_15323,N_15351);
or U15659 (N_15659,N_15068,N_15105);
nor U15660 (N_15660,N_15076,N_15248);
xnor U15661 (N_15661,N_15490,N_15211);
or U15662 (N_15662,N_15302,N_15254);
xor U15663 (N_15663,N_15197,N_15426);
nand U15664 (N_15664,N_15270,N_15040);
and U15665 (N_15665,N_15058,N_15498);
or U15666 (N_15666,N_15006,N_15244);
xnor U15667 (N_15667,N_15345,N_15109);
xor U15668 (N_15668,N_15021,N_15203);
nand U15669 (N_15669,N_15356,N_15383);
and U15670 (N_15670,N_15062,N_15497);
xor U15671 (N_15671,N_15359,N_15352);
or U15672 (N_15672,N_15148,N_15229);
nor U15673 (N_15673,N_15050,N_15407);
nand U15674 (N_15674,N_15434,N_15184);
nand U15675 (N_15675,N_15238,N_15043);
xor U15676 (N_15676,N_15207,N_15261);
or U15677 (N_15677,N_15382,N_15305);
xor U15678 (N_15678,N_15052,N_15335);
or U15679 (N_15679,N_15336,N_15024);
and U15680 (N_15680,N_15310,N_15318);
and U15681 (N_15681,N_15438,N_15065);
nor U15682 (N_15682,N_15150,N_15370);
xnor U15683 (N_15683,N_15354,N_15033);
nor U15684 (N_15684,N_15406,N_15198);
nand U15685 (N_15685,N_15189,N_15349);
nor U15686 (N_15686,N_15294,N_15478);
nor U15687 (N_15687,N_15492,N_15227);
xnor U15688 (N_15688,N_15486,N_15431);
xor U15689 (N_15689,N_15306,N_15275);
nand U15690 (N_15690,N_15448,N_15074);
and U15691 (N_15691,N_15285,N_15231);
or U15692 (N_15692,N_15156,N_15298);
nor U15693 (N_15693,N_15339,N_15253);
nand U15694 (N_15694,N_15160,N_15374);
or U15695 (N_15695,N_15029,N_15481);
xnor U15696 (N_15696,N_15164,N_15051);
nand U15697 (N_15697,N_15373,N_15411);
and U15698 (N_15698,N_15417,N_15077);
and U15699 (N_15699,N_15018,N_15432);
or U15700 (N_15700,N_15173,N_15396);
nor U15701 (N_15701,N_15219,N_15333);
and U15702 (N_15702,N_15243,N_15143);
xnor U15703 (N_15703,N_15039,N_15015);
nor U15704 (N_15704,N_15346,N_15387);
nand U15705 (N_15705,N_15344,N_15475);
nor U15706 (N_15706,N_15239,N_15415);
xnor U15707 (N_15707,N_15487,N_15464);
nand U15708 (N_15708,N_15165,N_15202);
xor U15709 (N_15709,N_15301,N_15041);
nor U15710 (N_15710,N_15287,N_15320);
and U15711 (N_15711,N_15185,N_15385);
and U15712 (N_15712,N_15470,N_15023);
nand U15713 (N_15713,N_15210,N_15366);
nor U15714 (N_15714,N_15070,N_15314);
or U15715 (N_15715,N_15402,N_15028);
and U15716 (N_15716,N_15247,N_15476);
nor U15717 (N_15717,N_15400,N_15390);
xnor U15718 (N_15718,N_15212,N_15435);
nand U15719 (N_15719,N_15137,N_15384);
nand U15720 (N_15720,N_15424,N_15466);
or U15721 (N_15721,N_15489,N_15027);
and U15722 (N_15722,N_15119,N_15205);
and U15723 (N_15723,N_15378,N_15461);
nor U15724 (N_15724,N_15135,N_15304);
nand U15725 (N_15725,N_15166,N_15368);
nand U15726 (N_15726,N_15377,N_15457);
nand U15727 (N_15727,N_15217,N_15196);
or U15728 (N_15728,N_15460,N_15465);
xor U15729 (N_15729,N_15291,N_15199);
and U15730 (N_15730,N_15083,N_15008);
and U15731 (N_15731,N_15329,N_15236);
nand U15732 (N_15732,N_15338,N_15034);
and U15733 (N_15733,N_15251,N_15279);
xor U15734 (N_15734,N_15365,N_15069);
nand U15735 (N_15735,N_15218,N_15322);
nand U15736 (N_15736,N_15495,N_15350);
xor U15737 (N_15737,N_15307,N_15397);
nand U15738 (N_15738,N_15224,N_15019);
nand U15739 (N_15739,N_15482,N_15182);
and U15740 (N_15740,N_15216,N_15347);
nor U15741 (N_15741,N_15128,N_15286);
nor U15742 (N_15742,N_15364,N_15315);
and U15743 (N_15743,N_15422,N_15391);
and U15744 (N_15744,N_15289,N_15179);
nor U15745 (N_15745,N_15168,N_15161);
nand U15746 (N_15746,N_15250,N_15056);
nand U15747 (N_15747,N_15319,N_15372);
nor U15748 (N_15748,N_15452,N_15463);
nand U15749 (N_15749,N_15151,N_15115);
nor U15750 (N_15750,N_15013,N_15280);
and U15751 (N_15751,N_15294,N_15316);
and U15752 (N_15752,N_15330,N_15113);
xor U15753 (N_15753,N_15091,N_15239);
nor U15754 (N_15754,N_15259,N_15131);
and U15755 (N_15755,N_15292,N_15480);
or U15756 (N_15756,N_15085,N_15248);
nand U15757 (N_15757,N_15130,N_15355);
and U15758 (N_15758,N_15099,N_15068);
nor U15759 (N_15759,N_15407,N_15031);
nand U15760 (N_15760,N_15150,N_15279);
xor U15761 (N_15761,N_15110,N_15391);
or U15762 (N_15762,N_15211,N_15209);
xor U15763 (N_15763,N_15292,N_15489);
xnor U15764 (N_15764,N_15353,N_15086);
and U15765 (N_15765,N_15134,N_15288);
and U15766 (N_15766,N_15267,N_15006);
nor U15767 (N_15767,N_15298,N_15087);
or U15768 (N_15768,N_15330,N_15262);
and U15769 (N_15769,N_15484,N_15173);
or U15770 (N_15770,N_15145,N_15302);
or U15771 (N_15771,N_15416,N_15066);
and U15772 (N_15772,N_15362,N_15448);
xor U15773 (N_15773,N_15233,N_15453);
nand U15774 (N_15774,N_15057,N_15245);
and U15775 (N_15775,N_15201,N_15059);
and U15776 (N_15776,N_15133,N_15125);
and U15777 (N_15777,N_15153,N_15096);
xor U15778 (N_15778,N_15330,N_15450);
xnor U15779 (N_15779,N_15432,N_15465);
nor U15780 (N_15780,N_15149,N_15408);
nand U15781 (N_15781,N_15318,N_15207);
nor U15782 (N_15782,N_15020,N_15442);
and U15783 (N_15783,N_15297,N_15298);
nand U15784 (N_15784,N_15219,N_15493);
or U15785 (N_15785,N_15469,N_15273);
or U15786 (N_15786,N_15046,N_15315);
xor U15787 (N_15787,N_15209,N_15164);
nand U15788 (N_15788,N_15374,N_15277);
nor U15789 (N_15789,N_15342,N_15311);
and U15790 (N_15790,N_15303,N_15157);
and U15791 (N_15791,N_15015,N_15166);
nor U15792 (N_15792,N_15485,N_15344);
nand U15793 (N_15793,N_15037,N_15061);
nand U15794 (N_15794,N_15351,N_15475);
and U15795 (N_15795,N_15084,N_15322);
nand U15796 (N_15796,N_15153,N_15465);
nand U15797 (N_15797,N_15193,N_15119);
xor U15798 (N_15798,N_15135,N_15374);
or U15799 (N_15799,N_15338,N_15317);
xor U15800 (N_15800,N_15310,N_15484);
nor U15801 (N_15801,N_15249,N_15223);
or U15802 (N_15802,N_15490,N_15449);
or U15803 (N_15803,N_15455,N_15282);
nand U15804 (N_15804,N_15176,N_15257);
nand U15805 (N_15805,N_15392,N_15166);
or U15806 (N_15806,N_15060,N_15038);
nor U15807 (N_15807,N_15006,N_15331);
or U15808 (N_15808,N_15406,N_15207);
nand U15809 (N_15809,N_15158,N_15328);
and U15810 (N_15810,N_15218,N_15158);
nand U15811 (N_15811,N_15126,N_15073);
or U15812 (N_15812,N_15472,N_15371);
xor U15813 (N_15813,N_15469,N_15048);
or U15814 (N_15814,N_15003,N_15335);
xnor U15815 (N_15815,N_15403,N_15229);
nand U15816 (N_15816,N_15497,N_15060);
xor U15817 (N_15817,N_15119,N_15200);
nor U15818 (N_15818,N_15448,N_15281);
xnor U15819 (N_15819,N_15219,N_15475);
nand U15820 (N_15820,N_15006,N_15288);
or U15821 (N_15821,N_15436,N_15448);
xor U15822 (N_15822,N_15428,N_15468);
or U15823 (N_15823,N_15246,N_15089);
and U15824 (N_15824,N_15398,N_15325);
or U15825 (N_15825,N_15499,N_15448);
or U15826 (N_15826,N_15105,N_15416);
xor U15827 (N_15827,N_15012,N_15480);
nor U15828 (N_15828,N_15260,N_15315);
or U15829 (N_15829,N_15276,N_15446);
xnor U15830 (N_15830,N_15387,N_15472);
xnor U15831 (N_15831,N_15383,N_15246);
xor U15832 (N_15832,N_15386,N_15277);
xnor U15833 (N_15833,N_15304,N_15137);
nor U15834 (N_15834,N_15231,N_15088);
or U15835 (N_15835,N_15352,N_15214);
or U15836 (N_15836,N_15114,N_15237);
nand U15837 (N_15837,N_15487,N_15322);
nor U15838 (N_15838,N_15487,N_15145);
xnor U15839 (N_15839,N_15231,N_15041);
nor U15840 (N_15840,N_15465,N_15354);
and U15841 (N_15841,N_15339,N_15199);
and U15842 (N_15842,N_15205,N_15176);
xor U15843 (N_15843,N_15157,N_15071);
nor U15844 (N_15844,N_15229,N_15357);
nand U15845 (N_15845,N_15131,N_15373);
and U15846 (N_15846,N_15376,N_15213);
xnor U15847 (N_15847,N_15338,N_15427);
and U15848 (N_15848,N_15301,N_15441);
xnor U15849 (N_15849,N_15329,N_15300);
nor U15850 (N_15850,N_15368,N_15429);
xor U15851 (N_15851,N_15282,N_15384);
nand U15852 (N_15852,N_15019,N_15398);
xnor U15853 (N_15853,N_15436,N_15485);
and U15854 (N_15854,N_15420,N_15276);
or U15855 (N_15855,N_15069,N_15072);
xor U15856 (N_15856,N_15413,N_15047);
nor U15857 (N_15857,N_15256,N_15187);
and U15858 (N_15858,N_15135,N_15009);
nor U15859 (N_15859,N_15161,N_15475);
nor U15860 (N_15860,N_15236,N_15330);
and U15861 (N_15861,N_15245,N_15162);
and U15862 (N_15862,N_15240,N_15242);
or U15863 (N_15863,N_15312,N_15040);
nor U15864 (N_15864,N_15257,N_15282);
nand U15865 (N_15865,N_15325,N_15223);
and U15866 (N_15866,N_15094,N_15235);
and U15867 (N_15867,N_15265,N_15007);
nand U15868 (N_15868,N_15024,N_15236);
xnor U15869 (N_15869,N_15213,N_15049);
or U15870 (N_15870,N_15197,N_15438);
and U15871 (N_15871,N_15311,N_15489);
nand U15872 (N_15872,N_15463,N_15454);
nor U15873 (N_15873,N_15025,N_15203);
nand U15874 (N_15874,N_15231,N_15205);
nand U15875 (N_15875,N_15430,N_15445);
nor U15876 (N_15876,N_15370,N_15012);
and U15877 (N_15877,N_15301,N_15395);
and U15878 (N_15878,N_15335,N_15169);
xor U15879 (N_15879,N_15429,N_15122);
xnor U15880 (N_15880,N_15181,N_15326);
nand U15881 (N_15881,N_15157,N_15316);
nand U15882 (N_15882,N_15207,N_15321);
nor U15883 (N_15883,N_15108,N_15244);
nor U15884 (N_15884,N_15147,N_15415);
nand U15885 (N_15885,N_15347,N_15430);
and U15886 (N_15886,N_15166,N_15038);
or U15887 (N_15887,N_15108,N_15397);
or U15888 (N_15888,N_15051,N_15087);
xor U15889 (N_15889,N_15466,N_15280);
nor U15890 (N_15890,N_15280,N_15451);
nand U15891 (N_15891,N_15248,N_15188);
nand U15892 (N_15892,N_15116,N_15270);
and U15893 (N_15893,N_15090,N_15191);
and U15894 (N_15894,N_15282,N_15035);
and U15895 (N_15895,N_15346,N_15253);
or U15896 (N_15896,N_15379,N_15487);
and U15897 (N_15897,N_15265,N_15367);
nand U15898 (N_15898,N_15126,N_15028);
nor U15899 (N_15899,N_15309,N_15456);
or U15900 (N_15900,N_15231,N_15115);
nor U15901 (N_15901,N_15367,N_15406);
xnor U15902 (N_15902,N_15161,N_15342);
xnor U15903 (N_15903,N_15101,N_15311);
nor U15904 (N_15904,N_15319,N_15365);
nor U15905 (N_15905,N_15310,N_15113);
and U15906 (N_15906,N_15227,N_15082);
nor U15907 (N_15907,N_15002,N_15303);
xnor U15908 (N_15908,N_15291,N_15043);
and U15909 (N_15909,N_15446,N_15432);
nand U15910 (N_15910,N_15394,N_15080);
nand U15911 (N_15911,N_15206,N_15005);
or U15912 (N_15912,N_15360,N_15017);
xor U15913 (N_15913,N_15146,N_15223);
nor U15914 (N_15914,N_15402,N_15267);
and U15915 (N_15915,N_15144,N_15293);
and U15916 (N_15916,N_15449,N_15038);
or U15917 (N_15917,N_15450,N_15047);
nor U15918 (N_15918,N_15056,N_15089);
and U15919 (N_15919,N_15450,N_15052);
nor U15920 (N_15920,N_15377,N_15134);
or U15921 (N_15921,N_15043,N_15316);
and U15922 (N_15922,N_15409,N_15387);
and U15923 (N_15923,N_15354,N_15211);
nand U15924 (N_15924,N_15316,N_15035);
and U15925 (N_15925,N_15471,N_15414);
or U15926 (N_15926,N_15487,N_15386);
nor U15927 (N_15927,N_15104,N_15169);
and U15928 (N_15928,N_15461,N_15153);
xnor U15929 (N_15929,N_15394,N_15313);
nand U15930 (N_15930,N_15240,N_15209);
nand U15931 (N_15931,N_15141,N_15486);
or U15932 (N_15932,N_15481,N_15347);
nor U15933 (N_15933,N_15161,N_15482);
nor U15934 (N_15934,N_15475,N_15293);
nand U15935 (N_15935,N_15454,N_15025);
nand U15936 (N_15936,N_15104,N_15069);
or U15937 (N_15937,N_15329,N_15497);
or U15938 (N_15938,N_15363,N_15425);
and U15939 (N_15939,N_15406,N_15126);
and U15940 (N_15940,N_15086,N_15263);
nand U15941 (N_15941,N_15288,N_15408);
nand U15942 (N_15942,N_15185,N_15440);
and U15943 (N_15943,N_15190,N_15210);
xor U15944 (N_15944,N_15149,N_15418);
or U15945 (N_15945,N_15064,N_15313);
nor U15946 (N_15946,N_15033,N_15191);
and U15947 (N_15947,N_15497,N_15195);
nand U15948 (N_15948,N_15125,N_15433);
and U15949 (N_15949,N_15166,N_15006);
nand U15950 (N_15950,N_15172,N_15115);
or U15951 (N_15951,N_15366,N_15166);
nand U15952 (N_15952,N_15078,N_15049);
and U15953 (N_15953,N_15204,N_15345);
or U15954 (N_15954,N_15178,N_15395);
and U15955 (N_15955,N_15136,N_15094);
or U15956 (N_15956,N_15263,N_15290);
nand U15957 (N_15957,N_15091,N_15342);
or U15958 (N_15958,N_15295,N_15161);
and U15959 (N_15959,N_15029,N_15373);
nor U15960 (N_15960,N_15374,N_15454);
nand U15961 (N_15961,N_15292,N_15062);
nand U15962 (N_15962,N_15328,N_15112);
xnor U15963 (N_15963,N_15474,N_15095);
nand U15964 (N_15964,N_15013,N_15083);
or U15965 (N_15965,N_15052,N_15230);
and U15966 (N_15966,N_15130,N_15441);
nor U15967 (N_15967,N_15340,N_15462);
nor U15968 (N_15968,N_15448,N_15279);
nand U15969 (N_15969,N_15301,N_15373);
and U15970 (N_15970,N_15293,N_15075);
nor U15971 (N_15971,N_15438,N_15335);
and U15972 (N_15972,N_15490,N_15383);
or U15973 (N_15973,N_15341,N_15189);
nand U15974 (N_15974,N_15135,N_15063);
nor U15975 (N_15975,N_15002,N_15325);
nand U15976 (N_15976,N_15079,N_15486);
nand U15977 (N_15977,N_15089,N_15353);
xor U15978 (N_15978,N_15054,N_15375);
nand U15979 (N_15979,N_15478,N_15368);
or U15980 (N_15980,N_15231,N_15120);
and U15981 (N_15981,N_15435,N_15391);
nand U15982 (N_15982,N_15387,N_15005);
nor U15983 (N_15983,N_15293,N_15333);
and U15984 (N_15984,N_15155,N_15270);
nand U15985 (N_15985,N_15026,N_15281);
nand U15986 (N_15986,N_15077,N_15123);
nand U15987 (N_15987,N_15111,N_15450);
nand U15988 (N_15988,N_15478,N_15418);
nand U15989 (N_15989,N_15417,N_15019);
nand U15990 (N_15990,N_15407,N_15079);
or U15991 (N_15991,N_15285,N_15027);
or U15992 (N_15992,N_15033,N_15050);
xnor U15993 (N_15993,N_15209,N_15232);
xnor U15994 (N_15994,N_15349,N_15278);
nor U15995 (N_15995,N_15217,N_15261);
and U15996 (N_15996,N_15182,N_15262);
nor U15997 (N_15997,N_15229,N_15290);
or U15998 (N_15998,N_15332,N_15425);
nor U15999 (N_15999,N_15152,N_15169);
xor U16000 (N_16000,N_15686,N_15768);
or U16001 (N_16001,N_15822,N_15631);
xnor U16002 (N_16002,N_15524,N_15875);
and U16003 (N_16003,N_15873,N_15698);
nor U16004 (N_16004,N_15780,N_15771);
and U16005 (N_16005,N_15630,N_15810);
xnor U16006 (N_16006,N_15702,N_15739);
or U16007 (N_16007,N_15654,N_15525);
xor U16008 (N_16008,N_15815,N_15639);
nor U16009 (N_16009,N_15658,N_15920);
xnor U16010 (N_16010,N_15939,N_15899);
nand U16011 (N_16011,N_15648,N_15688);
xor U16012 (N_16012,N_15730,N_15779);
xnor U16013 (N_16013,N_15552,N_15904);
nand U16014 (N_16014,N_15576,N_15689);
and U16015 (N_16015,N_15617,N_15667);
nand U16016 (N_16016,N_15990,N_15878);
and U16017 (N_16017,N_15529,N_15677);
nand U16018 (N_16018,N_15944,N_15930);
or U16019 (N_16019,N_15790,N_15752);
and U16020 (N_16020,N_15851,N_15574);
nor U16021 (N_16021,N_15567,N_15636);
xnor U16022 (N_16022,N_15547,N_15751);
or U16023 (N_16023,N_15870,N_15620);
or U16024 (N_16024,N_15653,N_15600);
nand U16025 (N_16025,N_15535,N_15956);
and U16026 (N_16026,N_15823,N_15788);
nand U16027 (N_16027,N_15932,N_15936);
nand U16028 (N_16028,N_15963,N_15989);
and U16029 (N_16029,N_15858,N_15545);
nand U16030 (N_16030,N_15760,N_15531);
nand U16031 (N_16031,N_15972,N_15901);
and U16032 (N_16032,N_15804,N_15881);
nand U16033 (N_16033,N_15616,N_15781);
or U16034 (N_16034,N_15664,N_15729);
nand U16035 (N_16035,N_15763,N_15610);
nor U16036 (N_16036,N_15697,N_15625);
nand U16037 (N_16037,N_15766,N_15871);
xor U16038 (N_16038,N_15755,N_15805);
and U16039 (N_16039,N_15782,N_15794);
or U16040 (N_16040,N_15951,N_15738);
and U16041 (N_16041,N_15706,N_15940);
xnor U16042 (N_16042,N_15573,N_15575);
xor U16043 (N_16043,N_15609,N_15937);
xor U16044 (N_16044,N_15721,N_15618);
nor U16045 (N_16045,N_15716,N_15743);
nand U16046 (N_16046,N_15627,N_15913);
or U16047 (N_16047,N_15519,N_15628);
xnor U16048 (N_16048,N_15701,N_15869);
or U16049 (N_16049,N_15731,N_15923);
xnor U16050 (N_16050,N_15744,N_15874);
or U16051 (N_16051,N_15590,N_15570);
xor U16052 (N_16052,N_15910,N_15727);
or U16053 (N_16053,N_15579,N_15872);
and U16054 (N_16054,N_15624,N_15934);
nor U16055 (N_16055,N_15943,N_15704);
xor U16056 (N_16056,N_15812,N_15546);
xor U16057 (N_16057,N_15839,N_15974);
and U16058 (N_16058,N_15537,N_15880);
or U16059 (N_16059,N_15971,N_15959);
xor U16060 (N_16060,N_15868,N_15829);
or U16061 (N_16061,N_15840,N_15973);
nor U16062 (N_16062,N_15824,N_15663);
nor U16063 (N_16063,N_15778,N_15997);
or U16064 (N_16064,N_15955,N_15544);
nor U16065 (N_16065,N_15717,N_15587);
and U16066 (N_16066,N_15911,N_15512);
nor U16067 (N_16067,N_15562,N_15542);
nor U16068 (N_16068,N_15853,N_15582);
or U16069 (N_16069,N_15977,N_15996);
nor U16070 (N_16070,N_15987,N_15789);
nand U16071 (N_16071,N_15854,N_15993);
xnor U16072 (N_16072,N_15611,N_15929);
or U16073 (N_16073,N_15994,N_15675);
nor U16074 (N_16074,N_15846,N_15799);
or U16075 (N_16075,N_15718,N_15680);
nand U16076 (N_16076,N_15979,N_15541);
or U16077 (N_16077,N_15841,N_15500);
and U16078 (N_16078,N_15563,N_15795);
nor U16079 (N_16079,N_15733,N_15510);
nand U16080 (N_16080,N_15598,N_15820);
or U16081 (N_16081,N_15926,N_15933);
nor U16082 (N_16082,N_15606,N_15695);
xor U16083 (N_16083,N_15999,N_15879);
nor U16084 (N_16084,N_15509,N_15608);
nor U16085 (N_16085,N_15859,N_15737);
or U16086 (N_16086,N_15862,N_15792);
or U16087 (N_16087,N_15539,N_15536);
or U16088 (N_16088,N_15641,N_15594);
nor U16089 (N_16089,N_15965,N_15674);
nand U16090 (N_16090,N_15523,N_15775);
or U16091 (N_16091,N_15821,N_15916);
nor U16092 (N_16092,N_15530,N_15762);
nor U16093 (N_16093,N_15534,N_15984);
nand U16094 (N_16094,N_15709,N_15960);
nand U16095 (N_16095,N_15982,N_15811);
nor U16096 (N_16096,N_15921,N_15572);
xnor U16097 (N_16097,N_15682,N_15985);
or U16098 (N_16098,N_15684,N_15734);
xnor U16099 (N_16099,N_15890,N_15966);
and U16100 (N_16100,N_15601,N_15801);
or U16101 (N_16101,N_15844,N_15903);
nand U16102 (N_16102,N_15833,N_15646);
nor U16103 (N_16103,N_15728,N_15758);
and U16104 (N_16104,N_15809,N_15816);
nand U16105 (N_16105,N_15679,N_15902);
xor U16106 (N_16106,N_15817,N_15668);
xnor U16107 (N_16107,N_15662,N_15976);
xnor U16108 (N_16108,N_15749,N_15818);
and U16109 (N_16109,N_15550,N_15660);
nand U16110 (N_16110,N_15741,N_15591);
nand U16111 (N_16111,N_15671,N_15757);
or U16112 (N_16112,N_15863,N_15520);
xnor U16113 (N_16113,N_15849,N_15998);
xor U16114 (N_16114,N_15597,N_15711);
and U16115 (N_16115,N_15707,N_15516);
or U16116 (N_16116,N_15569,N_15557);
xor U16117 (N_16117,N_15565,N_15586);
nand U16118 (N_16118,N_15918,N_15967);
or U16119 (N_16119,N_15772,N_15856);
or U16120 (N_16120,N_15885,N_15961);
and U16121 (N_16121,N_15835,N_15938);
and U16122 (N_16122,N_15619,N_15764);
or U16123 (N_16123,N_15538,N_15970);
xnor U16124 (N_16124,N_15896,N_15651);
xor U16125 (N_16125,N_15917,N_15696);
or U16126 (N_16126,N_15501,N_15725);
nand U16127 (N_16127,N_15533,N_15953);
nand U16128 (N_16128,N_15802,N_15640);
xor U16129 (N_16129,N_15831,N_15746);
nor U16130 (N_16130,N_15797,N_15635);
or U16131 (N_16131,N_15935,N_15908);
and U16132 (N_16132,N_15898,N_15687);
or U16133 (N_16133,N_15647,N_15946);
nor U16134 (N_16134,N_15566,N_15589);
nor U16135 (N_16135,N_15514,N_15740);
nor U16136 (N_16136,N_15643,N_15784);
nand U16137 (N_16137,N_15592,N_15753);
nor U16138 (N_16138,N_15596,N_15765);
and U16139 (N_16139,N_15588,N_15622);
and U16140 (N_16140,N_15659,N_15678);
nand U16141 (N_16141,N_15681,N_15876);
nor U16142 (N_16142,N_15549,N_15767);
xor U16143 (N_16143,N_15796,N_15694);
nand U16144 (N_16144,N_15852,N_15634);
xnor U16145 (N_16145,N_15700,N_15931);
or U16146 (N_16146,N_15585,N_15528);
nor U16147 (N_16147,N_15912,N_15507);
nand U16148 (N_16148,N_15632,N_15968);
xor U16149 (N_16149,N_15893,N_15756);
xnor U16150 (N_16150,N_15543,N_15564);
nand U16151 (N_16151,N_15715,N_15644);
xnor U16152 (N_16152,N_15515,N_15556);
nor U16153 (N_16153,N_15877,N_15607);
nor U16154 (N_16154,N_15978,N_15883);
or U16155 (N_16155,N_15814,N_15614);
or U16156 (N_16156,N_15922,N_15950);
xnor U16157 (N_16157,N_15992,N_15958);
and U16158 (N_16158,N_15577,N_15947);
or U16159 (N_16159,N_15626,N_15773);
nand U16160 (N_16160,N_15623,N_15754);
xor U16161 (N_16161,N_15941,N_15791);
nand U16162 (N_16162,N_15669,N_15793);
nand U16163 (N_16163,N_15558,N_15842);
or U16164 (N_16164,N_15672,N_15732);
xor U16165 (N_16165,N_15666,N_15602);
nor U16166 (N_16166,N_15712,N_15986);
and U16167 (N_16167,N_15551,N_15889);
and U16168 (N_16168,N_15806,N_15962);
and U16169 (N_16169,N_15866,N_15710);
nor U16170 (N_16170,N_15724,N_15895);
and U16171 (N_16171,N_15719,N_15803);
nand U16172 (N_16172,N_15919,N_15578);
xnor U16173 (N_16173,N_15526,N_15770);
or U16174 (N_16174,N_15703,N_15750);
nand U16175 (N_16175,N_15580,N_15857);
nor U16176 (N_16176,N_15900,N_15942);
or U16177 (N_16177,N_15786,N_15830);
or U16178 (N_16178,N_15532,N_15548);
or U16179 (N_16179,N_15502,N_15655);
xnor U16180 (N_16180,N_15522,N_15584);
or U16181 (N_16181,N_15503,N_15828);
nand U16182 (N_16182,N_15723,N_15665);
or U16183 (N_16183,N_15891,N_15774);
or U16184 (N_16184,N_15713,N_15670);
nor U16185 (N_16185,N_15924,N_15560);
nand U16186 (N_16186,N_15983,N_15692);
nand U16187 (N_16187,N_15508,N_15906);
nand U16188 (N_16188,N_15894,N_15554);
xor U16189 (N_16189,N_15599,N_15845);
or U16190 (N_16190,N_15887,N_15948);
nand U16191 (N_16191,N_15785,N_15981);
or U16192 (N_16192,N_15555,N_15553);
nor U16193 (N_16193,N_15540,N_15897);
and U16194 (N_16194,N_15783,N_15603);
or U16195 (N_16195,N_15988,N_15798);
and U16196 (N_16196,N_15800,N_15807);
and U16197 (N_16197,N_15676,N_15720);
nand U16198 (N_16198,N_15847,N_15886);
nor U16199 (N_16199,N_15595,N_15604);
or U16200 (N_16200,N_15691,N_15685);
and U16201 (N_16201,N_15907,N_15690);
nand U16202 (N_16202,N_15504,N_15884);
and U16203 (N_16203,N_15834,N_15980);
and U16204 (N_16204,N_15683,N_15642);
xnor U16205 (N_16205,N_15511,N_15559);
and U16206 (N_16206,N_15892,N_15527);
nand U16207 (N_16207,N_15615,N_15661);
xor U16208 (N_16208,N_15759,N_15928);
and U16209 (N_16209,N_15964,N_15518);
or U16210 (N_16210,N_15673,N_15745);
nor U16211 (N_16211,N_15952,N_15699);
and U16212 (N_16212,N_15949,N_15517);
xnor U16213 (N_16213,N_15726,N_15593);
nor U16214 (N_16214,N_15777,N_15705);
xor U16215 (N_16215,N_15819,N_15629);
nand U16216 (N_16216,N_15633,N_15568);
and U16217 (N_16217,N_15736,N_15832);
or U16218 (N_16218,N_15882,N_15905);
or U16219 (N_16219,N_15850,N_15969);
or U16220 (N_16220,N_15506,N_15776);
nor U16221 (N_16221,N_15722,N_15864);
nor U16222 (N_16222,N_15649,N_15714);
and U16223 (N_16223,N_15748,N_15915);
or U16224 (N_16224,N_15645,N_15927);
nand U16225 (N_16225,N_15652,N_15975);
nor U16226 (N_16226,N_15914,N_15865);
nor U16227 (N_16227,N_15827,N_15954);
nor U16228 (N_16228,N_15787,N_15761);
or U16229 (N_16229,N_15656,N_15708);
and U16230 (N_16230,N_15909,N_15769);
xnor U16231 (N_16231,N_15995,N_15808);
nand U16232 (N_16232,N_15735,N_15561);
and U16233 (N_16233,N_15657,N_15855);
xnor U16234 (N_16234,N_15513,N_15861);
nand U16235 (N_16235,N_15843,N_15867);
or U16236 (N_16236,N_15505,N_15621);
or U16237 (N_16237,N_15888,N_15742);
nand U16238 (N_16238,N_15612,N_15991);
xor U16239 (N_16239,N_15837,N_15957);
xnor U16240 (N_16240,N_15836,N_15945);
and U16241 (N_16241,N_15826,N_15650);
and U16242 (N_16242,N_15693,N_15848);
xor U16243 (N_16243,N_15825,N_15638);
nand U16244 (N_16244,N_15813,N_15605);
nor U16245 (N_16245,N_15571,N_15637);
nand U16246 (N_16246,N_15613,N_15860);
or U16247 (N_16247,N_15925,N_15747);
or U16248 (N_16248,N_15583,N_15838);
xnor U16249 (N_16249,N_15521,N_15581);
nor U16250 (N_16250,N_15921,N_15765);
nor U16251 (N_16251,N_15813,N_15993);
xor U16252 (N_16252,N_15671,N_15587);
nand U16253 (N_16253,N_15696,N_15597);
and U16254 (N_16254,N_15706,N_15928);
nor U16255 (N_16255,N_15581,N_15799);
nor U16256 (N_16256,N_15993,N_15947);
and U16257 (N_16257,N_15742,N_15525);
nand U16258 (N_16258,N_15898,N_15666);
and U16259 (N_16259,N_15695,N_15517);
nor U16260 (N_16260,N_15875,N_15528);
or U16261 (N_16261,N_15697,N_15658);
xor U16262 (N_16262,N_15508,N_15543);
and U16263 (N_16263,N_15739,N_15970);
or U16264 (N_16264,N_15926,N_15973);
nand U16265 (N_16265,N_15646,N_15936);
and U16266 (N_16266,N_15513,N_15729);
nor U16267 (N_16267,N_15893,N_15768);
nor U16268 (N_16268,N_15622,N_15694);
xnor U16269 (N_16269,N_15719,N_15908);
nor U16270 (N_16270,N_15546,N_15995);
xor U16271 (N_16271,N_15530,N_15732);
nand U16272 (N_16272,N_15696,N_15773);
or U16273 (N_16273,N_15511,N_15553);
or U16274 (N_16274,N_15952,N_15555);
xor U16275 (N_16275,N_15642,N_15901);
xor U16276 (N_16276,N_15890,N_15661);
nor U16277 (N_16277,N_15874,N_15551);
nor U16278 (N_16278,N_15619,N_15751);
and U16279 (N_16279,N_15509,N_15852);
nor U16280 (N_16280,N_15915,N_15668);
and U16281 (N_16281,N_15810,N_15579);
and U16282 (N_16282,N_15960,N_15656);
xor U16283 (N_16283,N_15629,N_15684);
and U16284 (N_16284,N_15881,N_15793);
or U16285 (N_16285,N_15951,N_15952);
xnor U16286 (N_16286,N_15918,N_15663);
nand U16287 (N_16287,N_15511,N_15883);
nand U16288 (N_16288,N_15707,N_15684);
nor U16289 (N_16289,N_15700,N_15868);
or U16290 (N_16290,N_15835,N_15771);
xor U16291 (N_16291,N_15698,N_15761);
xor U16292 (N_16292,N_15644,N_15983);
nand U16293 (N_16293,N_15758,N_15656);
xor U16294 (N_16294,N_15502,N_15522);
nor U16295 (N_16295,N_15630,N_15610);
nor U16296 (N_16296,N_15553,N_15876);
or U16297 (N_16297,N_15985,N_15765);
or U16298 (N_16298,N_15964,N_15756);
xnor U16299 (N_16299,N_15681,N_15960);
or U16300 (N_16300,N_15963,N_15829);
nor U16301 (N_16301,N_15920,N_15903);
nand U16302 (N_16302,N_15933,N_15895);
and U16303 (N_16303,N_15995,N_15832);
and U16304 (N_16304,N_15651,N_15759);
and U16305 (N_16305,N_15622,N_15536);
xor U16306 (N_16306,N_15678,N_15602);
or U16307 (N_16307,N_15697,N_15642);
and U16308 (N_16308,N_15602,N_15932);
or U16309 (N_16309,N_15965,N_15818);
or U16310 (N_16310,N_15708,N_15798);
nand U16311 (N_16311,N_15663,N_15572);
nand U16312 (N_16312,N_15690,N_15985);
nand U16313 (N_16313,N_15555,N_15542);
nand U16314 (N_16314,N_15726,N_15658);
nand U16315 (N_16315,N_15652,N_15809);
nor U16316 (N_16316,N_15783,N_15770);
and U16317 (N_16317,N_15633,N_15938);
and U16318 (N_16318,N_15675,N_15950);
xor U16319 (N_16319,N_15713,N_15681);
or U16320 (N_16320,N_15916,N_15751);
xnor U16321 (N_16321,N_15991,N_15804);
nor U16322 (N_16322,N_15821,N_15987);
xor U16323 (N_16323,N_15625,N_15894);
nor U16324 (N_16324,N_15948,N_15910);
xnor U16325 (N_16325,N_15743,N_15696);
xor U16326 (N_16326,N_15652,N_15830);
nor U16327 (N_16327,N_15679,N_15743);
or U16328 (N_16328,N_15864,N_15981);
nand U16329 (N_16329,N_15747,N_15965);
nor U16330 (N_16330,N_15810,N_15655);
and U16331 (N_16331,N_15723,N_15506);
xor U16332 (N_16332,N_15669,N_15765);
nand U16333 (N_16333,N_15788,N_15690);
nor U16334 (N_16334,N_15848,N_15780);
nor U16335 (N_16335,N_15955,N_15958);
or U16336 (N_16336,N_15585,N_15747);
or U16337 (N_16337,N_15835,N_15918);
xnor U16338 (N_16338,N_15993,N_15949);
and U16339 (N_16339,N_15667,N_15516);
nand U16340 (N_16340,N_15694,N_15764);
or U16341 (N_16341,N_15681,N_15801);
xnor U16342 (N_16342,N_15816,N_15751);
xor U16343 (N_16343,N_15973,N_15986);
nand U16344 (N_16344,N_15880,N_15840);
nand U16345 (N_16345,N_15748,N_15561);
or U16346 (N_16346,N_15829,N_15885);
nand U16347 (N_16347,N_15931,N_15757);
xor U16348 (N_16348,N_15959,N_15828);
or U16349 (N_16349,N_15900,N_15794);
or U16350 (N_16350,N_15504,N_15750);
xnor U16351 (N_16351,N_15510,N_15567);
nand U16352 (N_16352,N_15723,N_15712);
nand U16353 (N_16353,N_15560,N_15554);
nor U16354 (N_16354,N_15828,N_15985);
nand U16355 (N_16355,N_15638,N_15798);
and U16356 (N_16356,N_15876,N_15513);
and U16357 (N_16357,N_15870,N_15854);
nor U16358 (N_16358,N_15559,N_15764);
xnor U16359 (N_16359,N_15613,N_15624);
nand U16360 (N_16360,N_15525,N_15703);
nand U16361 (N_16361,N_15710,N_15781);
and U16362 (N_16362,N_15728,N_15648);
xnor U16363 (N_16363,N_15574,N_15923);
nand U16364 (N_16364,N_15643,N_15591);
and U16365 (N_16365,N_15938,N_15943);
and U16366 (N_16366,N_15529,N_15754);
xor U16367 (N_16367,N_15807,N_15933);
or U16368 (N_16368,N_15871,N_15893);
xnor U16369 (N_16369,N_15811,N_15637);
or U16370 (N_16370,N_15976,N_15936);
or U16371 (N_16371,N_15678,N_15570);
nor U16372 (N_16372,N_15818,N_15832);
or U16373 (N_16373,N_15980,N_15749);
or U16374 (N_16374,N_15886,N_15549);
nand U16375 (N_16375,N_15807,N_15633);
or U16376 (N_16376,N_15680,N_15618);
xnor U16377 (N_16377,N_15895,N_15700);
and U16378 (N_16378,N_15789,N_15630);
xnor U16379 (N_16379,N_15745,N_15833);
and U16380 (N_16380,N_15529,N_15730);
nand U16381 (N_16381,N_15553,N_15809);
nor U16382 (N_16382,N_15608,N_15901);
xor U16383 (N_16383,N_15760,N_15567);
nand U16384 (N_16384,N_15795,N_15951);
xnor U16385 (N_16385,N_15684,N_15903);
nand U16386 (N_16386,N_15907,N_15830);
or U16387 (N_16387,N_15778,N_15676);
nor U16388 (N_16388,N_15904,N_15876);
nor U16389 (N_16389,N_15505,N_15773);
xnor U16390 (N_16390,N_15577,N_15851);
nand U16391 (N_16391,N_15901,N_15895);
nor U16392 (N_16392,N_15501,N_15538);
nand U16393 (N_16393,N_15885,N_15667);
or U16394 (N_16394,N_15812,N_15754);
xor U16395 (N_16395,N_15537,N_15785);
and U16396 (N_16396,N_15740,N_15780);
or U16397 (N_16397,N_15969,N_15778);
nand U16398 (N_16398,N_15868,N_15977);
xor U16399 (N_16399,N_15918,N_15953);
or U16400 (N_16400,N_15706,N_15852);
or U16401 (N_16401,N_15712,N_15724);
nand U16402 (N_16402,N_15763,N_15768);
xnor U16403 (N_16403,N_15857,N_15642);
or U16404 (N_16404,N_15915,N_15565);
nor U16405 (N_16405,N_15583,N_15875);
nor U16406 (N_16406,N_15522,N_15702);
nor U16407 (N_16407,N_15633,N_15827);
nand U16408 (N_16408,N_15911,N_15537);
nand U16409 (N_16409,N_15992,N_15976);
nand U16410 (N_16410,N_15588,N_15747);
nand U16411 (N_16411,N_15762,N_15774);
xor U16412 (N_16412,N_15654,N_15608);
xnor U16413 (N_16413,N_15878,N_15526);
nor U16414 (N_16414,N_15635,N_15814);
xor U16415 (N_16415,N_15586,N_15546);
nor U16416 (N_16416,N_15528,N_15854);
nand U16417 (N_16417,N_15855,N_15690);
and U16418 (N_16418,N_15891,N_15818);
and U16419 (N_16419,N_15648,N_15558);
or U16420 (N_16420,N_15619,N_15591);
xnor U16421 (N_16421,N_15539,N_15923);
nor U16422 (N_16422,N_15960,N_15894);
nor U16423 (N_16423,N_15887,N_15954);
nor U16424 (N_16424,N_15569,N_15782);
nor U16425 (N_16425,N_15740,N_15980);
or U16426 (N_16426,N_15837,N_15721);
nor U16427 (N_16427,N_15608,N_15725);
and U16428 (N_16428,N_15817,N_15842);
nand U16429 (N_16429,N_15646,N_15985);
or U16430 (N_16430,N_15659,N_15663);
and U16431 (N_16431,N_15576,N_15750);
xor U16432 (N_16432,N_15507,N_15941);
nand U16433 (N_16433,N_15743,N_15795);
or U16434 (N_16434,N_15691,N_15821);
or U16435 (N_16435,N_15985,N_15752);
or U16436 (N_16436,N_15928,N_15838);
nor U16437 (N_16437,N_15652,N_15822);
nor U16438 (N_16438,N_15598,N_15662);
nor U16439 (N_16439,N_15862,N_15807);
or U16440 (N_16440,N_15918,N_15777);
nor U16441 (N_16441,N_15636,N_15953);
nand U16442 (N_16442,N_15675,N_15755);
nand U16443 (N_16443,N_15912,N_15589);
xnor U16444 (N_16444,N_15819,N_15620);
xor U16445 (N_16445,N_15527,N_15768);
nand U16446 (N_16446,N_15938,N_15521);
nand U16447 (N_16447,N_15756,N_15801);
and U16448 (N_16448,N_15737,N_15590);
nand U16449 (N_16449,N_15971,N_15675);
and U16450 (N_16450,N_15738,N_15984);
nor U16451 (N_16451,N_15575,N_15902);
nand U16452 (N_16452,N_15565,N_15576);
xnor U16453 (N_16453,N_15619,N_15980);
or U16454 (N_16454,N_15656,N_15543);
nor U16455 (N_16455,N_15815,N_15596);
and U16456 (N_16456,N_15836,N_15841);
and U16457 (N_16457,N_15538,N_15903);
xor U16458 (N_16458,N_15809,N_15868);
nor U16459 (N_16459,N_15865,N_15527);
and U16460 (N_16460,N_15639,N_15631);
nor U16461 (N_16461,N_15955,N_15590);
or U16462 (N_16462,N_15950,N_15944);
nor U16463 (N_16463,N_15927,N_15585);
nor U16464 (N_16464,N_15754,N_15677);
nor U16465 (N_16465,N_15938,N_15813);
nor U16466 (N_16466,N_15887,N_15763);
or U16467 (N_16467,N_15642,N_15742);
or U16468 (N_16468,N_15995,N_15565);
xnor U16469 (N_16469,N_15741,N_15926);
nand U16470 (N_16470,N_15870,N_15662);
and U16471 (N_16471,N_15521,N_15691);
nand U16472 (N_16472,N_15599,N_15961);
nor U16473 (N_16473,N_15758,N_15849);
nor U16474 (N_16474,N_15852,N_15666);
nor U16475 (N_16475,N_15819,N_15539);
nor U16476 (N_16476,N_15672,N_15760);
nor U16477 (N_16477,N_15889,N_15627);
nand U16478 (N_16478,N_15943,N_15920);
or U16479 (N_16479,N_15778,N_15693);
xor U16480 (N_16480,N_15788,N_15560);
or U16481 (N_16481,N_15659,N_15510);
xor U16482 (N_16482,N_15655,N_15660);
or U16483 (N_16483,N_15704,N_15511);
or U16484 (N_16484,N_15723,N_15735);
or U16485 (N_16485,N_15590,N_15663);
or U16486 (N_16486,N_15557,N_15920);
xnor U16487 (N_16487,N_15637,N_15517);
or U16488 (N_16488,N_15773,N_15877);
nand U16489 (N_16489,N_15533,N_15885);
and U16490 (N_16490,N_15688,N_15697);
xor U16491 (N_16491,N_15683,N_15890);
and U16492 (N_16492,N_15587,N_15743);
nor U16493 (N_16493,N_15620,N_15884);
or U16494 (N_16494,N_15585,N_15804);
xnor U16495 (N_16495,N_15960,N_15926);
and U16496 (N_16496,N_15642,N_15576);
or U16497 (N_16497,N_15969,N_15537);
or U16498 (N_16498,N_15619,N_15748);
nand U16499 (N_16499,N_15743,N_15885);
and U16500 (N_16500,N_16015,N_16431);
or U16501 (N_16501,N_16047,N_16325);
nor U16502 (N_16502,N_16154,N_16253);
or U16503 (N_16503,N_16311,N_16211);
nor U16504 (N_16504,N_16316,N_16274);
and U16505 (N_16505,N_16169,N_16062);
nand U16506 (N_16506,N_16018,N_16330);
xor U16507 (N_16507,N_16455,N_16328);
xor U16508 (N_16508,N_16232,N_16382);
nor U16509 (N_16509,N_16057,N_16304);
nor U16510 (N_16510,N_16161,N_16288);
or U16511 (N_16511,N_16172,N_16081);
nor U16512 (N_16512,N_16291,N_16261);
and U16513 (N_16513,N_16195,N_16343);
or U16514 (N_16514,N_16397,N_16315);
nand U16515 (N_16515,N_16077,N_16359);
and U16516 (N_16516,N_16386,N_16190);
nor U16517 (N_16517,N_16108,N_16162);
nor U16518 (N_16518,N_16177,N_16473);
and U16519 (N_16519,N_16220,N_16210);
nand U16520 (N_16520,N_16034,N_16410);
nand U16521 (N_16521,N_16224,N_16284);
or U16522 (N_16522,N_16490,N_16050);
or U16523 (N_16523,N_16024,N_16332);
xor U16524 (N_16524,N_16353,N_16061);
nor U16525 (N_16525,N_16206,N_16404);
xnor U16526 (N_16526,N_16339,N_16028);
xnor U16527 (N_16527,N_16046,N_16358);
and U16528 (N_16528,N_16064,N_16442);
xor U16529 (N_16529,N_16043,N_16390);
nor U16530 (N_16530,N_16485,N_16040);
nor U16531 (N_16531,N_16368,N_16144);
and U16532 (N_16532,N_16111,N_16414);
nor U16533 (N_16533,N_16407,N_16114);
nand U16534 (N_16534,N_16171,N_16476);
or U16535 (N_16535,N_16341,N_16488);
nor U16536 (N_16536,N_16091,N_16228);
nor U16537 (N_16537,N_16187,N_16376);
nor U16538 (N_16538,N_16138,N_16234);
nand U16539 (N_16539,N_16191,N_16205);
or U16540 (N_16540,N_16217,N_16375);
nor U16541 (N_16541,N_16105,N_16035);
and U16542 (N_16542,N_16340,N_16327);
or U16543 (N_16543,N_16347,N_16042);
or U16544 (N_16544,N_16329,N_16367);
nand U16545 (N_16545,N_16394,N_16317);
nor U16546 (N_16546,N_16370,N_16381);
or U16547 (N_16547,N_16478,N_16308);
or U16548 (N_16548,N_16117,N_16365);
and U16549 (N_16549,N_16307,N_16448);
nand U16550 (N_16550,N_16148,N_16299);
nor U16551 (N_16551,N_16262,N_16361);
or U16552 (N_16552,N_16493,N_16158);
and U16553 (N_16553,N_16238,N_16230);
xor U16554 (N_16554,N_16385,N_16441);
nand U16555 (N_16555,N_16349,N_16480);
xor U16556 (N_16556,N_16196,N_16427);
and U16557 (N_16557,N_16173,N_16292);
xnor U16558 (N_16558,N_16188,N_16344);
and U16559 (N_16559,N_16444,N_16312);
nand U16560 (N_16560,N_16486,N_16103);
or U16561 (N_16561,N_16082,N_16006);
xnor U16562 (N_16562,N_16302,N_16495);
xor U16563 (N_16563,N_16146,N_16240);
xor U16564 (N_16564,N_16076,N_16152);
or U16565 (N_16565,N_16156,N_16039);
xnor U16566 (N_16566,N_16363,N_16120);
nand U16567 (N_16567,N_16099,N_16342);
nand U16568 (N_16568,N_16023,N_16213);
or U16569 (N_16569,N_16216,N_16219);
xor U16570 (N_16570,N_16428,N_16295);
nand U16571 (N_16571,N_16372,N_16499);
or U16572 (N_16572,N_16101,N_16435);
xnor U16573 (N_16573,N_16463,N_16352);
and U16574 (N_16574,N_16189,N_16025);
nor U16575 (N_16575,N_16019,N_16041);
nor U16576 (N_16576,N_16182,N_16471);
or U16577 (N_16577,N_16440,N_16197);
or U16578 (N_16578,N_16069,N_16377);
or U16579 (N_16579,N_16297,N_16250);
and U16580 (N_16580,N_16249,N_16464);
nand U16581 (N_16581,N_16010,N_16033);
nand U16582 (N_16582,N_16183,N_16003);
nand U16583 (N_16583,N_16242,N_16174);
nand U16584 (N_16584,N_16017,N_16357);
xnor U16585 (N_16585,N_16130,N_16301);
nand U16586 (N_16586,N_16271,N_16348);
xnor U16587 (N_16587,N_16439,N_16294);
and U16588 (N_16588,N_16167,N_16026);
or U16589 (N_16589,N_16207,N_16395);
or U16590 (N_16590,N_16212,N_16413);
and U16591 (N_16591,N_16085,N_16354);
nor U16592 (N_16592,N_16009,N_16432);
xor U16593 (N_16593,N_16326,N_16371);
or U16594 (N_16594,N_16036,N_16362);
or U16595 (N_16595,N_16131,N_16402);
and U16596 (N_16596,N_16084,N_16489);
and U16597 (N_16597,N_16477,N_16151);
nor U16598 (N_16598,N_16123,N_16110);
or U16599 (N_16599,N_16481,N_16129);
and U16600 (N_16600,N_16396,N_16383);
nor U16601 (N_16601,N_16143,N_16264);
or U16602 (N_16602,N_16202,N_16350);
nand U16603 (N_16603,N_16054,N_16140);
nor U16604 (N_16604,N_16051,N_16425);
and U16605 (N_16605,N_16459,N_16200);
xor U16606 (N_16606,N_16384,N_16412);
nand U16607 (N_16607,N_16000,N_16479);
or U16608 (N_16608,N_16165,N_16155);
nand U16609 (N_16609,N_16388,N_16235);
nand U16610 (N_16610,N_16094,N_16223);
nand U16611 (N_16611,N_16373,N_16424);
nor U16612 (N_16612,N_16239,N_16136);
nor U16613 (N_16613,N_16285,N_16322);
nand U16614 (N_16614,N_16090,N_16355);
nor U16615 (N_16615,N_16303,N_16268);
and U16616 (N_16616,N_16360,N_16309);
and U16617 (N_16617,N_16072,N_16055);
nand U16618 (N_16618,N_16293,N_16184);
or U16619 (N_16619,N_16159,N_16345);
and U16620 (N_16620,N_16453,N_16139);
and U16621 (N_16621,N_16258,N_16289);
nand U16622 (N_16622,N_16192,N_16119);
nor U16623 (N_16623,N_16460,N_16245);
and U16624 (N_16624,N_16321,N_16106);
xnor U16625 (N_16625,N_16469,N_16150);
nand U16626 (N_16626,N_16014,N_16333);
xnor U16627 (N_16627,N_16487,N_16225);
or U16628 (N_16628,N_16020,N_16109);
nor U16629 (N_16629,N_16031,N_16443);
or U16630 (N_16630,N_16075,N_16267);
and U16631 (N_16631,N_16180,N_16121);
and U16632 (N_16632,N_16276,N_16113);
nor U16633 (N_16633,N_16287,N_16233);
nand U16634 (N_16634,N_16491,N_16338);
or U16635 (N_16635,N_16472,N_16204);
or U16636 (N_16636,N_16056,N_16430);
or U16637 (N_16637,N_16128,N_16405);
and U16638 (N_16638,N_16208,N_16122);
or U16639 (N_16639,N_16265,N_16497);
and U16640 (N_16640,N_16351,N_16005);
or U16641 (N_16641,N_16016,N_16408);
xnor U16642 (N_16642,N_16421,N_16401);
or U16643 (N_16643,N_16420,N_16203);
nor U16644 (N_16644,N_16236,N_16132);
nand U16645 (N_16645,N_16466,N_16314);
nor U16646 (N_16646,N_16305,N_16393);
nor U16647 (N_16647,N_16484,N_16324);
or U16648 (N_16648,N_16279,N_16241);
or U16649 (N_16649,N_16079,N_16380);
xnor U16650 (N_16650,N_16115,N_16112);
nor U16651 (N_16651,N_16013,N_16454);
and U16652 (N_16652,N_16283,N_16116);
nand U16653 (N_16653,N_16399,N_16290);
or U16654 (N_16654,N_16429,N_16356);
nor U16655 (N_16655,N_16398,N_16319);
nor U16656 (N_16656,N_16059,N_16474);
nor U16657 (N_16657,N_16296,N_16147);
and U16658 (N_16658,N_16073,N_16145);
xnor U16659 (N_16659,N_16181,N_16237);
and U16660 (N_16660,N_16462,N_16104);
or U16661 (N_16661,N_16157,N_16446);
xor U16662 (N_16662,N_16346,N_16142);
and U16663 (N_16663,N_16227,N_16369);
nand U16664 (N_16664,N_16437,N_16135);
nor U16665 (N_16665,N_16280,N_16176);
and U16666 (N_16666,N_16045,N_16275);
nand U16667 (N_16667,N_16201,N_16281);
xnor U16668 (N_16668,N_16323,N_16374);
or U16669 (N_16669,N_16364,N_16418);
nor U16670 (N_16670,N_16273,N_16387);
and U16671 (N_16671,N_16214,N_16198);
nand U16672 (N_16672,N_16067,N_16063);
nand U16673 (N_16673,N_16492,N_16331);
nand U16674 (N_16674,N_16263,N_16178);
xnor U16675 (N_16675,N_16298,N_16186);
xor U16676 (N_16676,N_16193,N_16087);
nand U16677 (N_16677,N_16272,N_16080);
or U16678 (N_16678,N_16461,N_16458);
or U16679 (N_16679,N_16053,N_16068);
nand U16680 (N_16680,N_16248,N_16391);
or U16681 (N_16681,N_16226,N_16259);
nor U16682 (N_16682,N_16411,N_16124);
and U16683 (N_16683,N_16447,N_16185);
xnor U16684 (N_16684,N_16027,N_16436);
nand U16685 (N_16685,N_16266,N_16433);
and U16686 (N_16686,N_16475,N_16282);
and U16687 (N_16687,N_16175,N_16086);
and U16688 (N_16688,N_16300,N_16277);
and U16689 (N_16689,N_16163,N_16048);
xnor U16690 (N_16690,N_16002,N_16215);
or U16691 (N_16691,N_16423,N_16335);
nor U16692 (N_16692,N_16199,N_16445);
nand U16693 (N_16693,N_16070,N_16452);
or U16694 (N_16694,N_16337,N_16030);
and U16695 (N_16695,N_16416,N_16247);
or U16696 (N_16696,N_16456,N_16389);
and U16697 (N_16697,N_16494,N_16270);
xor U16698 (N_16698,N_16194,N_16286);
or U16699 (N_16699,N_16470,N_16438);
or U16700 (N_16700,N_16320,N_16221);
and U16701 (N_16701,N_16037,N_16457);
or U16702 (N_16702,N_16089,N_16060);
nor U16703 (N_16703,N_16336,N_16229);
nor U16704 (N_16704,N_16310,N_16083);
nor U16705 (N_16705,N_16022,N_16318);
xor U16706 (N_16706,N_16392,N_16095);
and U16707 (N_16707,N_16256,N_16243);
nor U16708 (N_16708,N_16450,N_16251);
xor U16709 (N_16709,N_16004,N_16141);
xnor U16710 (N_16710,N_16096,N_16231);
or U16711 (N_16711,N_16137,N_16278);
nand U16712 (N_16712,N_16170,N_16021);
or U16713 (N_16713,N_16038,N_16451);
nor U16714 (N_16714,N_16306,N_16313);
and U16715 (N_16715,N_16066,N_16160);
nand U16716 (N_16716,N_16078,N_16001);
xnor U16717 (N_16717,N_16255,N_16422);
nor U16718 (N_16718,N_16100,N_16465);
or U16719 (N_16719,N_16269,N_16400);
xnor U16720 (N_16720,N_16149,N_16126);
nand U16721 (N_16721,N_16222,N_16483);
and U16722 (N_16722,N_16052,N_16209);
nand U16723 (N_16723,N_16403,N_16007);
xnor U16724 (N_16724,N_16029,N_16102);
xnor U16725 (N_16725,N_16012,N_16107);
nor U16726 (N_16726,N_16134,N_16127);
xnor U16727 (N_16727,N_16498,N_16426);
nand U16728 (N_16728,N_16164,N_16366);
nor U16729 (N_16729,N_16097,N_16334);
and U16730 (N_16730,N_16179,N_16092);
nand U16731 (N_16731,N_16049,N_16257);
nor U16732 (N_16732,N_16449,N_16496);
or U16733 (N_16733,N_16125,N_16252);
nand U16734 (N_16734,N_16406,N_16071);
and U16735 (N_16735,N_16133,N_16260);
xor U16736 (N_16736,N_16011,N_16254);
and U16737 (N_16737,N_16246,N_16058);
nor U16738 (N_16738,N_16098,N_16417);
xnor U16739 (N_16739,N_16244,N_16153);
xnor U16740 (N_16740,N_16093,N_16468);
xnor U16741 (N_16741,N_16467,N_16074);
nor U16742 (N_16742,N_16168,N_16044);
or U16743 (N_16743,N_16008,N_16118);
nor U16744 (N_16744,N_16166,N_16379);
nand U16745 (N_16745,N_16434,N_16415);
or U16746 (N_16746,N_16482,N_16065);
nand U16747 (N_16747,N_16378,N_16419);
and U16748 (N_16748,N_16218,N_16032);
and U16749 (N_16749,N_16409,N_16088);
nand U16750 (N_16750,N_16354,N_16291);
nor U16751 (N_16751,N_16380,N_16188);
nor U16752 (N_16752,N_16060,N_16094);
nand U16753 (N_16753,N_16316,N_16334);
and U16754 (N_16754,N_16294,N_16313);
nor U16755 (N_16755,N_16035,N_16001);
and U16756 (N_16756,N_16131,N_16000);
nand U16757 (N_16757,N_16239,N_16008);
and U16758 (N_16758,N_16454,N_16167);
nor U16759 (N_16759,N_16142,N_16351);
and U16760 (N_16760,N_16458,N_16454);
nor U16761 (N_16761,N_16435,N_16071);
or U16762 (N_16762,N_16403,N_16378);
nor U16763 (N_16763,N_16240,N_16175);
nand U16764 (N_16764,N_16447,N_16123);
nand U16765 (N_16765,N_16247,N_16154);
nand U16766 (N_16766,N_16302,N_16301);
nor U16767 (N_16767,N_16248,N_16174);
nand U16768 (N_16768,N_16156,N_16473);
or U16769 (N_16769,N_16230,N_16315);
nor U16770 (N_16770,N_16194,N_16404);
nand U16771 (N_16771,N_16414,N_16469);
xnor U16772 (N_16772,N_16148,N_16281);
xor U16773 (N_16773,N_16223,N_16220);
nor U16774 (N_16774,N_16039,N_16078);
and U16775 (N_16775,N_16002,N_16160);
and U16776 (N_16776,N_16395,N_16108);
and U16777 (N_16777,N_16499,N_16219);
or U16778 (N_16778,N_16413,N_16323);
nor U16779 (N_16779,N_16311,N_16007);
nor U16780 (N_16780,N_16478,N_16262);
or U16781 (N_16781,N_16157,N_16113);
or U16782 (N_16782,N_16026,N_16321);
and U16783 (N_16783,N_16071,N_16096);
and U16784 (N_16784,N_16137,N_16078);
and U16785 (N_16785,N_16000,N_16308);
nand U16786 (N_16786,N_16424,N_16286);
and U16787 (N_16787,N_16341,N_16277);
nand U16788 (N_16788,N_16005,N_16159);
nor U16789 (N_16789,N_16133,N_16348);
and U16790 (N_16790,N_16307,N_16186);
nor U16791 (N_16791,N_16432,N_16211);
xor U16792 (N_16792,N_16256,N_16332);
or U16793 (N_16793,N_16467,N_16314);
xnor U16794 (N_16794,N_16121,N_16475);
nand U16795 (N_16795,N_16238,N_16470);
xnor U16796 (N_16796,N_16438,N_16047);
xnor U16797 (N_16797,N_16392,N_16200);
xor U16798 (N_16798,N_16198,N_16217);
nand U16799 (N_16799,N_16137,N_16190);
nor U16800 (N_16800,N_16266,N_16328);
xor U16801 (N_16801,N_16406,N_16489);
nand U16802 (N_16802,N_16047,N_16280);
or U16803 (N_16803,N_16325,N_16388);
nand U16804 (N_16804,N_16146,N_16246);
and U16805 (N_16805,N_16363,N_16271);
nand U16806 (N_16806,N_16089,N_16404);
and U16807 (N_16807,N_16032,N_16244);
nor U16808 (N_16808,N_16376,N_16470);
nor U16809 (N_16809,N_16073,N_16007);
nand U16810 (N_16810,N_16040,N_16278);
nor U16811 (N_16811,N_16280,N_16140);
nor U16812 (N_16812,N_16030,N_16110);
xnor U16813 (N_16813,N_16057,N_16387);
or U16814 (N_16814,N_16387,N_16082);
and U16815 (N_16815,N_16109,N_16119);
nor U16816 (N_16816,N_16289,N_16410);
xor U16817 (N_16817,N_16227,N_16295);
nor U16818 (N_16818,N_16238,N_16403);
and U16819 (N_16819,N_16018,N_16087);
or U16820 (N_16820,N_16040,N_16086);
nor U16821 (N_16821,N_16273,N_16482);
nand U16822 (N_16822,N_16482,N_16227);
nor U16823 (N_16823,N_16339,N_16348);
xnor U16824 (N_16824,N_16200,N_16004);
nor U16825 (N_16825,N_16224,N_16302);
nand U16826 (N_16826,N_16349,N_16226);
nand U16827 (N_16827,N_16017,N_16432);
nor U16828 (N_16828,N_16229,N_16370);
nor U16829 (N_16829,N_16463,N_16167);
xnor U16830 (N_16830,N_16387,N_16462);
xor U16831 (N_16831,N_16221,N_16277);
or U16832 (N_16832,N_16196,N_16112);
and U16833 (N_16833,N_16032,N_16014);
and U16834 (N_16834,N_16020,N_16498);
nand U16835 (N_16835,N_16327,N_16212);
xor U16836 (N_16836,N_16412,N_16061);
xnor U16837 (N_16837,N_16078,N_16254);
or U16838 (N_16838,N_16336,N_16057);
nand U16839 (N_16839,N_16367,N_16074);
nor U16840 (N_16840,N_16428,N_16169);
and U16841 (N_16841,N_16206,N_16417);
nand U16842 (N_16842,N_16427,N_16136);
or U16843 (N_16843,N_16486,N_16412);
and U16844 (N_16844,N_16195,N_16033);
xor U16845 (N_16845,N_16292,N_16128);
and U16846 (N_16846,N_16338,N_16216);
and U16847 (N_16847,N_16423,N_16322);
nand U16848 (N_16848,N_16396,N_16053);
nand U16849 (N_16849,N_16371,N_16164);
nor U16850 (N_16850,N_16061,N_16005);
xnor U16851 (N_16851,N_16017,N_16459);
nor U16852 (N_16852,N_16264,N_16201);
nand U16853 (N_16853,N_16420,N_16294);
or U16854 (N_16854,N_16146,N_16124);
nand U16855 (N_16855,N_16181,N_16030);
or U16856 (N_16856,N_16379,N_16269);
xor U16857 (N_16857,N_16148,N_16314);
and U16858 (N_16858,N_16497,N_16499);
xor U16859 (N_16859,N_16049,N_16083);
nand U16860 (N_16860,N_16378,N_16157);
xor U16861 (N_16861,N_16011,N_16266);
xnor U16862 (N_16862,N_16388,N_16120);
nor U16863 (N_16863,N_16425,N_16328);
or U16864 (N_16864,N_16358,N_16153);
xor U16865 (N_16865,N_16134,N_16276);
and U16866 (N_16866,N_16173,N_16448);
xnor U16867 (N_16867,N_16328,N_16398);
or U16868 (N_16868,N_16443,N_16414);
nand U16869 (N_16869,N_16402,N_16250);
nor U16870 (N_16870,N_16041,N_16369);
nand U16871 (N_16871,N_16150,N_16087);
and U16872 (N_16872,N_16272,N_16147);
or U16873 (N_16873,N_16089,N_16474);
xor U16874 (N_16874,N_16367,N_16089);
xnor U16875 (N_16875,N_16487,N_16407);
nor U16876 (N_16876,N_16184,N_16313);
and U16877 (N_16877,N_16035,N_16116);
xnor U16878 (N_16878,N_16032,N_16361);
nand U16879 (N_16879,N_16193,N_16402);
and U16880 (N_16880,N_16438,N_16482);
or U16881 (N_16881,N_16227,N_16496);
and U16882 (N_16882,N_16300,N_16245);
xor U16883 (N_16883,N_16330,N_16187);
xnor U16884 (N_16884,N_16092,N_16182);
nor U16885 (N_16885,N_16209,N_16000);
nor U16886 (N_16886,N_16098,N_16471);
xnor U16887 (N_16887,N_16345,N_16265);
nand U16888 (N_16888,N_16236,N_16015);
or U16889 (N_16889,N_16123,N_16036);
xor U16890 (N_16890,N_16457,N_16298);
xor U16891 (N_16891,N_16233,N_16215);
xor U16892 (N_16892,N_16238,N_16474);
nor U16893 (N_16893,N_16226,N_16445);
and U16894 (N_16894,N_16464,N_16156);
or U16895 (N_16895,N_16472,N_16216);
xor U16896 (N_16896,N_16284,N_16212);
or U16897 (N_16897,N_16373,N_16341);
or U16898 (N_16898,N_16342,N_16392);
xor U16899 (N_16899,N_16021,N_16136);
or U16900 (N_16900,N_16216,N_16129);
xnor U16901 (N_16901,N_16186,N_16258);
xnor U16902 (N_16902,N_16065,N_16223);
or U16903 (N_16903,N_16227,N_16411);
nor U16904 (N_16904,N_16239,N_16462);
and U16905 (N_16905,N_16346,N_16184);
nor U16906 (N_16906,N_16116,N_16249);
xor U16907 (N_16907,N_16364,N_16068);
nand U16908 (N_16908,N_16268,N_16021);
nand U16909 (N_16909,N_16372,N_16349);
nor U16910 (N_16910,N_16450,N_16151);
xnor U16911 (N_16911,N_16274,N_16288);
xor U16912 (N_16912,N_16307,N_16195);
nand U16913 (N_16913,N_16084,N_16419);
xnor U16914 (N_16914,N_16161,N_16272);
nand U16915 (N_16915,N_16214,N_16066);
and U16916 (N_16916,N_16297,N_16038);
or U16917 (N_16917,N_16334,N_16286);
nor U16918 (N_16918,N_16340,N_16065);
or U16919 (N_16919,N_16271,N_16408);
nand U16920 (N_16920,N_16004,N_16026);
xor U16921 (N_16921,N_16347,N_16406);
or U16922 (N_16922,N_16160,N_16051);
nor U16923 (N_16923,N_16303,N_16230);
xnor U16924 (N_16924,N_16407,N_16337);
or U16925 (N_16925,N_16289,N_16182);
nand U16926 (N_16926,N_16071,N_16462);
nor U16927 (N_16927,N_16295,N_16189);
or U16928 (N_16928,N_16277,N_16373);
and U16929 (N_16929,N_16107,N_16324);
nor U16930 (N_16930,N_16488,N_16354);
and U16931 (N_16931,N_16154,N_16258);
or U16932 (N_16932,N_16429,N_16269);
nand U16933 (N_16933,N_16453,N_16492);
xor U16934 (N_16934,N_16277,N_16432);
nor U16935 (N_16935,N_16341,N_16257);
and U16936 (N_16936,N_16143,N_16218);
or U16937 (N_16937,N_16032,N_16321);
nand U16938 (N_16938,N_16315,N_16072);
and U16939 (N_16939,N_16238,N_16292);
xnor U16940 (N_16940,N_16313,N_16305);
or U16941 (N_16941,N_16203,N_16136);
xor U16942 (N_16942,N_16308,N_16241);
nor U16943 (N_16943,N_16394,N_16045);
nor U16944 (N_16944,N_16329,N_16211);
nor U16945 (N_16945,N_16066,N_16410);
nor U16946 (N_16946,N_16294,N_16343);
xnor U16947 (N_16947,N_16187,N_16063);
nor U16948 (N_16948,N_16286,N_16111);
nor U16949 (N_16949,N_16004,N_16082);
nand U16950 (N_16950,N_16210,N_16399);
xor U16951 (N_16951,N_16403,N_16492);
or U16952 (N_16952,N_16487,N_16426);
or U16953 (N_16953,N_16065,N_16177);
nand U16954 (N_16954,N_16452,N_16375);
and U16955 (N_16955,N_16248,N_16461);
nand U16956 (N_16956,N_16212,N_16142);
or U16957 (N_16957,N_16143,N_16035);
xnor U16958 (N_16958,N_16467,N_16393);
xnor U16959 (N_16959,N_16215,N_16112);
nand U16960 (N_16960,N_16416,N_16422);
nor U16961 (N_16961,N_16263,N_16019);
xnor U16962 (N_16962,N_16366,N_16058);
nand U16963 (N_16963,N_16190,N_16483);
nor U16964 (N_16964,N_16166,N_16236);
xor U16965 (N_16965,N_16457,N_16145);
or U16966 (N_16966,N_16373,N_16180);
nand U16967 (N_16967,N_16353,N_16413);
xnor U16968 (N_16968,N_16154,N_16302);
nand U16969 (N_16969,N_16158,N_16215);
nor U16970 (N_16970,N_16479,N_16260);
xor U16971 (N_16971,N_16272,N_16235);
nor U16972 (N_16972,N_16006,N_16255);
nand U16973 (N_16973,N_16195,N_16474);
or U16974 (N_16974,N_16399,N_16136);
nor U16975 (N_16975,N_16056,N_16095);
nor U16976 (N_16976,N_16262,N_16203);
nor U16977 (N_16977,N_16069,N_16395);
xnor U16978 (N_16978,N_16067,N_16333);
and U16979 (N_16979,N_16183,N_16238);
nor U16980 (N_16980,N_16457,N_16092);
nor U16981 (N_16981,N_16109,N_16390);
nand U16982 (N_16982,N_16494,N_16089);
nor U16983 (N_16983,N_16427,N_16244);
and U16984 (N_16984,N_16432,N_16041);
nand U16985 (N_16985,N_16155,N_16431);
and U16986 (N_16986,N_16140,N_16301);
or U16987 (N_16987,N_16323,N_16248);
nand U16988 (N_16988,N_16015,N_16195);
nor U16989 (N_16989,N_16239,N_16168);
xnor U16990 (N_16990,N_16369,N_16247);
nor U16991 (N_16991,N_16132,N_16215);
or U16992 (N_16992,N_16166,N_16089);
and U16993 (N_16993,N_16490,N_16466);
and U16994 (N_16994,N_16411,N_16053);
and U16995 (N_16995,N_16073,N_16224);
xnor U16996 (N_16996,N_16191,N_16274);
nand U16997 (N_16997,N_16354,N_16312);
nor U16998 (N_16998,N_16323,N_16353);
and U16999 (N_16999,N_16362,N_16377);
nand U17000 (N_17000,N_16519,N_16510);
and U17001 (N_17001,N_16918,N_16976);
nor U17002 (N_17002,N_16779,N_16514);
and U17003 (N_17003,N_16993,N_16921);
nor U17004 (N_17004,N_16875,N_16681);
xnor U17005 (N_17005,N_16694,N_16782);
or U17006 (N_17006,N_16788,N_16702);
xnor U17007 (N_17007,N_16617,N_16530);
nor U17008 (N_17008,N_16877,N_16748);
nor U17009 (N_17009,N_16879,N_16847);
xnor U17010 (N_17010,N_16715,N_16883);
and U17011 (N_17011,N_16683,N_16611);
or U17012 (N_17012,N_16943,N_16502);
nand U17013 (N_17013,N_16790,N_16718);
nor U17014 (N_17014,N_16789,N_16516);
and U17015 (N_17015,N_16769,N_16795);
nor U17016 (N_17016,N_16590,N_16658);
or U17017 (N_17017,N_16953,N_16816);
nand U17018 (N_17018,N_16619,N_16900);
nor U17019 (N_17019,N_16648,N_16717);
nand U17020 (N_17020,N_16886,N_16987);
nor U17021 (N_17021,N_16614,N_16928);
and U17022 (N_17022,N_16935,N_16692);
nand U17023 (N_17023,N_16913,N_16642);
or U17024 (N_17024,N_16861,N_16863);
xor U17025 (N_17025,N_16930,N_16624);
and U17026 (N_17026,N_16696,N_16950);
xor U17027 (N_17027,N_16641,N_16963);
nor U17028 (N_17028,N_16738,N_16830);
nand U17029 (N_17029,N_16966,N_16739);
nand U17030 (N_17030,N_16610,N_16821);
and U17031 (N_17031,N_16616,N_16629);
nor U17032 (N_17032,N_16815,N_16531);
xor U17033 (N_17033,N_16526,N_16991);
and U17034 (N_17034,N_16688,N_16547);
and U17035 (N_17035,N_16955,N_16798);
xor U17036 (N_17036,N_16994,N_16832);
and U17037 (N_17037,N_16975,N_16850);
xor U17038 (N_17038,N_16705,N_16727);
xor U17039 (N_17039,N_16587,N_16577);
nand U17040 (N_17040,N_16764,N_16890);
nand U17041 (N_17041,N_16562,N_16603);
and U17042 (N_17042,N_16982,N_16908);
and U17043 (N_17043,N_16527,N_16843);
nor U17044 (N_17044,N_16649,N_16778);
nand U17045 (N_17045,N_16689,N_16969);
nand U17046 (N_17046,N_16709,N_16541);
nor U17047 (N_17047,N_16672,N_16523);
nor U17048 (N_17048,N_16907,N_16631);
nand U17049 (N_17049,N_16786,N_16645);
and U17050 (N_17050,N_16671,N_16811);
nand U17051 (N_17051,N_16747,N_16916);
nor U17052 (N_17052,N_16989,N_16840);
nand U17053 (N_17053,N_16557,N_16712);
or U17054 (N_17054,N_16854,N_16568);
nor U17055 (N_17055,N_16653,N_16754);
nand U17056 (N_17056,N_16597,N_16549);
nand U17057 (N_17057,N_16996,N_16920);
or U17058 (N_17058,N_16759,N_16942);
and U17059 (N_17059,N_16765,N_16901);
and U17060 (N_17060,N_16538,N_16984);
xnor U17061 (N_17061,N_16876,N_16652);
nor U17062 (N_17062,N_16520,N_16539);
nor U17063 (N_17063,N_16882,N_16505);
xor U17064 (N_17064,N_16693,N_16885);
nand U17065 (N_17065,N_16753,N_16731);
nor U17066 (N_17066,N_16599,N_16501);
and U17067 (N_17067,N_16728,N_16504);
nor U17068 (N_17068,N_16826,N_16902);
nor U17069 (N_17069,N_16823,N_16615);
or U17070 (N_17070,N_16690,N_16936);
nand U17071 (N_17071,N_16896,N_16714);
and U17072 (N_17072,N_16824,N_16536);
or U17073 (N_17073,N_16721,N_16726);
and U17074 (N_17074,N_16851,N_16667);
and U17075 (N_17075,N_16745,N_16944);
and U17076 (N_17076,N_16707,N_16849);
nor U17077 (N_17077,N_16656,N_16810);
or U17078 (N_17078,N_16654,N_16762);
nor U17079 (N_17079,N_16939,N_16743);
nand U17080 (N_17080,N_16684,N_16595);
or U17081 (N_17081,N_16540,N_16682);
xor U17082 (N_17082,N_16749,N_16899);
xor U17083 (N_17083,N_16912,N_16589);
or U17084 (N_17084,N_16873,N_16904);
or U17085 (N_17085,N_16618,N_16639);
nor U17086 (N_17086,N_16767,N_16601);
nor U17087 (N_17087,N_16981,N_16632);
nand U17088 (N_17088,N_16646,N_16805);
nor U17089 (N_17089,N_16897,N_16914);
nand U17090 (N_17090,N_16970,N_16915);
or U17091 (N_17091,N_16543,N_16793);
or U17092 (N_17092,N_16723,N_16535);
nor U17093 (N_17093,N_16691,N_16609);
xor U17094 (N_17094,N_16522,N_16933);
nor U17095 (N_17095,N_16867,N_16881);
nand U17096 (N_17096,N_16623,N_16665);
nor U17097 (N_17097,N_16529,N_16818);
and U17098 (N_17098,N_16860,N_16679);
nor U17099 (N_17099,N_16554,N_16932);
or U17100 (N_17100,N_16750,N_16852);
or U17101 (N_17101,N_16704,N_16697);
nor U17102 (N_17102,N_16663,N_16725);
nor U17103 (N_17103,N_16834,N_16643);
nor U17104 (N_17104,N_16986,N_16708);
nor U17105 (N_17105,N_16760,N_16698);
or U17106 (N_17106,N_16768,N_16898);
nand U17107 (N_17107,N_16862,N_16870);
or U17108 (N_17108,N_16507,N_16559);
nand U17109 (N_17109,N_16751,N_16657);
nand U17110 (N_17110,N_16829,N_16763);
or U17111 (N_17111,N_16509,N_16736);
and U17112 (N_17112,N_16974,N_16819);
nor U17113 (N_17113,N_16513,N_16758);
or U17114 (N_17114,N_16700,N_16952);
nand U17115 (N_17115,N_16905,N_16940);
nand U17116 (N_17116,N_16521,N_16500);
xnor U17117 (N_17117,N_16638,N_16868);
xor U17118 (N_17118,N_16732,N_16848);
nand U17119 (N_17119,N_16670,N_16550);
xor U17120 (N_17120,N_16808,N_16894);
and U17121 (N_17121,N_16719,N_16836);
and U17122 (N_17122,N_16729,N_16580);
and U17123 (N_17123,N_16796,N_16792);
nor U17124 (N_17124,N_16674,N_16591);
xor U17125 (N_17125,N_16865,N_16605);
and U17126 (N_17126,N_16978,N_16911);
nor U17127 (N_17127,N_16613,N_16560);
nand U17128 (N_17128,N_16677,N_16695);
nor U17129 (N_17129,N_16666,N_16569);
xor U17130 (N_17130,N_16831,N_16737);
nand U17131 (N_17131,N_16553,N_16735);
nand U17132 (N_17132,N_16872,N_16888);
or U17133 (N_17133,N_16716,N_16965);
and U17134 (N_17134,N_16518,N_16977);
or U17135 (N_17135,N_16673,N_16630);
nand U17136 (N_17136,N_16581,N_16701);
or U17137 (N_17137,N_16551,N_16926);
or U17138 (N_17138,N_16946,N_16909);
xnor U17139 (N_17139,N_16724,N_16884);
nand U17140 (N_17140,N_16892,N_16676);
xnor U17141 (N_17141,N_16534,N_16962);
nor U17142 (N_17142,N_16576,N_16917);
nor U17143 (N_17143,N_16506,N_16703);
nor U17144 (N_17144,N_16803,N_16903);
or U17145 (N_17145,N_16659,N_16644);
and U17146 (N_17146,N_16746,N_16878);
xnor U17147 (N_17147,N_16864,N_16895);
and U17148 (N_17148,N_16572,N_16838);
xor U17149 (N_17149,N_16957,N_16844);
or U17150 (N_17150,N_16621,N_16660);
and U17151 (N_17151,N_16801,N_16706);
or U17152 (N_17152,N_16710,N_16687);
nor U17153 (N_17153,N_16937,N_16797);
and U17154 (N_17154,N_16855,N_16919);
or U17155 (N_17155,N_16794,N_16612);
nand U17156 (N_17156,N_16575,N_16999);
or U17157 (N_17157,N_16842,N_16800);
and U17158 (N_17158,N_16961,N_16563);
or U17159 (N_17159,N_16556,N_16635);
xnor U17160 (N_17160,N_16958,N_16813);
or U17161 (N_17161,N_16592,N_16925);
or U17162 (N_17162,N_16713,N_16776);
and U17163 (N_17163,N_16806,N_16584);
xnor U17164 (N_17164,N_16812,N_16809);
xor U17165 (N_17165,N_16734,N_16585);
or U17166 (N_17166,N_16625,N_16668);
nand U17167 (N_17167,N_16835,N_16633);
nor U17168 (N_17168,N_16814,N_16608);
nand U17169 (N_17169,N_16985,N_16561);
nor U17170 (N_17170,N_16740,N_16906);
nor U17171 (N_17171,N_16512,N_16941);
nand U17172 (N_17172,N_16678,N_16774);
or U17173 (N_17173,N_16775,N_16564);
or U17174 (N_17174,N_16664,N_16945);
nor U17175 (N_17175,N_16777,N_16533);
or U17176 (N_17176,N_16755,N_16785);
xnor U17177 (N_17177,N_16711,N_16511);
or U17178 (N_17178,N_16545,N_16983);
xor U17179 (N_17179,N_16650,N_16820);
xnor U17180 (N_17180,N_16596,N_16634);
xor U17181 (N_17181,N_16922,N_16787);
xor U17182 (N_17182,N_16620,N_16802);
xor U17183 (N_17183,N_16604,N_16600);
or U17184 (N_17184,N_16686,N_16532);
nand U17185 (N_17185,N_16756,N_16579);
or U17186 (N_17186,N_16742,N_16980);
nor U17187 (N_17187,N_16781,N_16567);
or U17188 (N_17188,N_16964,N_16929);
and U17189 (N_17189,N_16626,N_16992);
and U17190 (N_17190,N_16927,N_16997);
xor U17191 (N_17191,N_16967,N_16990);
nand U17192 (N_17192,N_16761,N_16858);
nand U17193 (N_17193,N_16524,N_16766);
or U17194 (N_17194,N_16947,N_16893);
or U17195 (N_17195,N_16948,N_16807);
nand U17196 (N_17196,N_16733,N_16949);
xnor U17197 (N_17197,N_16770,N_16588);
nand U17198 (N_17198,N_16586,N_16924);
xnor U17199 (N_17199,N_16871,N_16574);
xor U17200 (N_17200,N_16637,N_16817);
or U17201 (N_17201,N_16791,N_16773);
nand U17202 (N_17202,N_16972,N_16566);
nor U17203 (N_17203,N_16661,N_16573);
nand U17204 (N_17204,N_16874,N_16784);
nand U17205 (N_17205,N_16602,N_16910);
or U17206 (N_17206,N_16675,N_16833);
xor U17207 (N_17207,N_16845,N_16846);
and U17208 (N_17208,N_16598,N_16866);
nor U17209 (N_17209,N_16960,N_16627);
nor U17210 (N_17210,N_16571,N_16889);
and U17211 (N_17211,N_16951,N_16869);
or U17212 (N_17212,N_16954,N_16685);
nor U17213 (N_17213,N_16828,N_16772);
and U17214 (N_17214,N_16655,N_16544);
and U17215 (N_17215,N_16923,N_16730);
xor U17216 (N_17216,N_16517,N_16622);
or U17217 (N_17217,N_16570,N_16503);
nand U17218 (N_17218,N_16578,N_16565);
nand U17219 (N_17219,N_16979,N_16752);
nand U17220 (N_17220,N_16555,N_16841);
xnor U17221 (N_17221,N_16822,N_16891);
nor U17222 (N_17222,N_16548,N_16537);
nand U17223 (N_17223,N_16827,N_16780);
xnor U17224 (N_17224,N_16528,N_16931);
nand U17225 (N_17225,N_16662,N_16856);
and U17226 (N_17226,N_16998,N_16959);
or U17227 (N_17227,N_16783,N_16722);
and U17228 (N_17228,N_16825,N_16583);
and U17229 (N_17229,N_16651,N_16525);
or U17230 (N_17230,N_16552,N_16515);
xnor U17231 (N_17231,N_16973,N_16938);
xor U17232 (N_17232,N_16680,N_16593);
nor U17233 (N_17233,N_16988,N_16647);
or U17234 (N_17234,N_16607,N_16546);
nor U17235 (N_17235,N_16628,N_16640);
nor U17236 (N_17236,N_16636,N_16669);
and U17237 (N_17237,N_16857,N_16744);
nor U17238 (N_17238,N_16968,N_16799);
xnor U17239 (N_17239,N_16771,N_16956);
xor U17240 (N_17240,N_16839,N_16558);
and U17241 (N_17241,N_16594,N_16508);
xor U17242 (N_17242,N_16887,N_16757);
and U17243 (N_17243,N_16582,N_16804);
or U17244 (N_17244,N_16934,N_16699);
or U17245 (N_17245,N_16859,N_16720);
xor U17246 (N_17246,N_16542,N_16995);
nand U17247 (N_17247,N_16741,N_16853);
nor U17248 (N_17248,N_16971,N_16837);
nor U17249 (N_17249,N_16880,N_16606);
nand U17250 (N_17250,N_16921,N_16810);
or U17251 (N_17251,N_16663,N_16977);
nor U17252 (N_17252,N_16814,N_16807);
nor U17253 (N_17253,N_16570,N_16830);
or U17254 (N_17254,N_16693,N_16906);
or U17255 (N_17255,N_16793,N_16907);
nor U17256 (N_17256,N_16970,N_16986);
nand U17257 (N_17257,N_16627,N_16683);
xor U17258 (N_17258,N_16655,N_16914);
nor U17259 (N_17259,N_16804,N_16677);
nand U17260 (N_17260,N_16757,N_16860);
or U17261 (N_17261,N_16708,N_16614);
and U17262 (N_17262,N_16598,N_16573);
or U17263 (N_17263,N_16575,N_16976);
nand U17264 (N_17264,N_16595,N_16983);
xor U17265 (N_17265,N_16835,N_16808);
nor U17266 (N_17266,N_16836,N_16985);
xnor U17267 (N_17267,N_16802,N_16977);
nor U17268 (N_17268,N_16836,N_16587);
and U17269 (N_17269,N_16678,N_16879);
xor U17270 (N_17270,N_16971,N_16810);
nor U17271 (N_17271,N_16676,N_16838);
nand U17272 (N_17272,N_16764,N_16554);
xor U17273 (N_17273,N_16755,N_16542);
or U17274 (N_17274,N_16764,N_16695);
or U17275 (N_17275,N_16578,N_16795);
and U17276 (N_17276,N_16913,N_16986);
and U17277 (N_17277,N_16546,N_16536);
or U17278 (N_17278,N_16805,N_16924);
or U17279 (N_17279,N_16776,N_16835);
nor U17280 (N_17280,N_16519,N_16794);
xnor U17281 (N_17281,N_16771,N_16895);
nor U17282 (N_17282,N_16738,N_16539);
or U17283 (N_17283,N_16855,N_16583);
nand U17284 (N_17284,N_16822,N_16576);
nand U17285 (N_17285,N_16842,N_16557);
nor U17286 (N_17286,N_16721,N_16600);
nor U17287 (N_17287,N_16642,N_16732);
nor U17288 (N_17288,N_16731,N_16531);
or U17289 (N_17289,N_16600,N_16582);
nor U17290 (N_17290,N_16585,N_16746);
nor U17291 (N_17291,N_16641,N_16648);
nor U17292 (N_17292,N_16824,N_16906);
xor U17293 (N_17293,N_16753,N_16868);
xnor U17294 (N_17294,N_16698,N_16539);
nand U17295 (N_17295,N_16656,N_16702);
xnor U17296 (N_17296,N_16880,N_16598);
or U17297 (N_17297,N_16588,N_16907);
nand U17298 (N_17298,N_16514,N_16529);
and U17299 (N_17299,N_16542,N_16614);
and U17300 (N_17300,N_16512,N_16550);
xnor U17301 (N_17301,N_16870,N_16520);
or U17302 (N_17302,N_16707,N_16997);
or U17303 (N_17303,N_16648,N_16931);
nor U17304 (N_17304,N_16535,N_16737);
nor U17305 (N_17305,N_16983,N_16934);
xnor U17306 (N_17306,N_16837,N_16518);
or U17307 (N_17307,N_16654,N_16527);
xnor U17308 (N_17308,N_16668,N_16945);
nor U17309 (N_17309,N_16984,N_16587);
nor U17310 (N_17310,N_16831,N_16610);
xor U17311 (N_17311,N_16507,N_16862);
and U17312 (N_17312,N_16891,N_16881);
or U17313 (N_17313,N_16814,N_16848);
xnor U17314 (N_17314,N_16653,N_16854);
nand U17315 (N_17315,N_16832,N_16511);
and U17316 (N_17316,N_16720,N_16928);
xor U17317 (N_17317,N_16730,N_16716);
xnor U17318 (N_17318,N_16895,N_16713);
xnor U17319 (N_17319,N_16922,N_16861);
nand U17320 (N_17320,N_16876,N_16703);
nand U17321 (N_17321,N_16547,N_16685);
xnor U17322 (N_17322,N_16892,N_16927);
nand U17323 (N_17323,N_16625,N_16577);
or U17324 (N_17324,N_16982,N_16822);
nor U17325 (N_17325,N_16733,N_16903);
xor U17326 (N_17326,N_16509,N_16693);
nor U17327 (N_17327,N_16942,N_16638);
xnor U17328 (N_17328,N_16654,N_16546);
nor U17329 (N_17329,N_16627,N_16535);
or U17330 (N_17330,N_16829,N_16597);
or U17331 (N_17331,N_16965,N_16892);
nor U17332 (N_17332,N_16742,N_16505);
nor U17333 (N_17333,N_16656,N_16866);
nor U17334 (N_17334,N_16958,N_16636);
nand U17335 (N_17335,N_16538,N_16688);
nand U17336 (N_17336,N_16933,N_16916);
nand U17337 (N_17337,N_16661,N_16613);
xnor U17338 (N_17338,N_16966,N_16533);
nand U17339 (N_17339,N_16597,N_16691);
or U17340 (N_17340,N_16711,N_16538);
nor U17341 (N_17341,N_16510,N_16926);
xor U17342 (N_17342,N_16949,N_16577);
nand U17343 (N_17343,N_16638,N_16708);
and U17344 (N_17344,N_16946,N_16760);
or U17345 (N_17345,N_16636,N_16963);
and U17346 (N_17346,N_16535,N_16503);
and U17347 (N_17347,N_16703,N_16700);
or U17348 (N_17348,N_16860,N_16623);
xor U17349 (N_17349,N_16961,N_16996);
or U17350 (N_17350,N_16979,N_16538);
nand U17351 (N_17351,N_16854,N_16942);
nor U17352 (N_17352,N_16995,N_16569);
or U17353 (N_17353,N_16964,N_16975);
or U17354 (N_17354,N_16895,N_16997);
xor U17355 (N_17355,N_16936,N_16823);
or U17356 (N_17356,N_16989,N_16854);
nor U17357 (N_17357,N_16740,N_16774);
nand U17358 (N_17358,N_16600,N_16993);
nand U17359 (N_17359,N_16715,N_16779);
nor U17360 (N_17360,N_16580,N_16795);
xor U17361 (N_17361,N_16572,N_16754);
and U17362 (N_17362,N_16795,N_16529);
nand U17363 (N_17363,N_16938,N_16763);
or U17364 (N_17364,N_16629,N_16652);
nor U17365 (N_17365,N_16548,N_16767);
or U17366 (N_17366,N_16697,N_16588);
or U17367 (N_17367,N_16695,N_16744);
nand U17368 (N_17368,N_16681,N_16608);
or U17369 (N_17369,N_16742,N_16786);
nand U17370 (N_17370,N_16817,N_16926);
nor U17371 (N_17371,N_16590,N_16500);
and U17372 (N_17372,N_16995,N_16950);
xnor U17373 (N_17373,N_16658,N_16708);
and U17374 (N_17374,N_16919,N_16688);
xnor U17375 (N_17375,N_16652,N_16722);
xnor U17376 (N_17376,N_16572,N_16643);
and U17377 (N_17377,N_16793,N_16742);
nor U17378 (N_17378,N_16683,N_16591);
xor U17379 (N_17379,N_16823,N_16609);
nor U17380 (N_17380,N_16644,N_16797);
and U17381 (N_17381,N_16537,N_16738);
nor U17382 (N_17382,N_16852,N_16533);
xor U17383 (N_17383,N_16588,N_16526);
xor U17384 (N_17384,N_16757,N_16679);
nand U17385 (N_17385,N_16854,N_16606);
and U17386 (N_17386,N_16667,N_16608);
xnor U17387 (N_17387,N_16714,N_16599);
and U17388 (N_17388,N_16834,N_16551);
or U17389 (N_17389,N_16705,N_16564);
and U17390 (N_17390,N_16992,N_16933);
nor U17391 (N_17391,N_16962,N_16564);
xor U17392 (N_17392,N_16814,N_16899);
or U17393 (N_17393,N_16710,N_16891);
nand U17394 (N_17394,N_16551,N_16630);
nand U17395 (N_17395,N_16976,N_16532);
and U17396 (N_17396,N_16624,N_16570);
nor U17397 (N_17397,N_16945,N_16554);
xor U17398 (N_17398,N_16894,N_16690);
nor U17399 (N_17399,N_16683,N_16861);
xnor U17400 (N_17400,N_16875,N_16640);
and U17401 (N_17401,N_16871,N_16924);
and U17402 (N_17402,N_16715,N_16961);
or U17403 (N_17403,N_16721,N_16911);
xnor U17404 (N_17404,N_16757,N_16756);
nand U17405 (N_17405,N_16995,N_16917);
nand U17406 (N_17406,N_16993,N_16817);
xnor U17407 (N_17407,N_16557,N_16727);
xor U17408 (N_17408,N_16824,N_16953);
or U17409 (N_17409,N_16590,N_16747);
nand U17410 (N_17410,N_16634,N_16500);
and U17411 (N_17411,N_16997,N_16741);
and U17412 (N_17412,N_16930,N_16853);
xor U17413 (N_17413,N_16804,N_16545);
or U17414 (N_17414,N_16953,N_16950);
or U17415 (N_17415,N_16572,N_16533);
nand U17416 (N_17416,N_16731,N_16871);
and U17417 (N_17417,N_16882,N_16616);
nor U17418 (N_17418,N_16762,N_16822);
nand U17419 (N_17419,N_16748,N_16923);
nor U17420 (N_17420,N_16751,N_16699);
or U17421 (N_17421,N_16597,N_16948);
nand U17422 (N_17422,N_16719,N_16528);
xnor U17423 (N_17423,N_16802,N_16749);
nand U17424 (N_17424,N_16505,N_16678);
xor U17425 (N_17425,N_16689,N_16805);
or U17426 (N_17426,N_16937,N_16786);
nor U17427 (N_17427,N_16747,N_16978);
or U17428 (N_17428,N_16833,N_16625);
and U17429 (N_17429,N_16790,N_16633);
or U17430 (N_17430,N_16874,N_16805);
nor U17431 (N_17431,N_16730,N_16786);
nor U17432 (N_17432,N_16757,N_16924);
and U17433 (N_17433,N_16963,N_16631);
nand U17434 (N_17434,N_16537,N_16927);
nor U17435 (N_17435,N_16587,N_16739);
xnor U17436 (N_17436,N_16668,N_16626);
xor U17437 (N_17437,N_16891,N_16690);
nor U17438 (N_17438,N_16597,N_16919);
and U17439 (N_17439,N_16692,N_16540);
and U17440 (N_17440,N_16830,N_16795);
or U17441 (N_17441,N_16506,N_16537);
xnor U17442 (N_17442,N_16740,N_16762);
or U17443 (N_17443,N_16795,N_16772);
and U17444 (N_17444,N_16858,N_16880);
or U17445 (N_17445,N_16602,N_16542);
and U17446 (N_17446,N_16820,N_16785);
nor U17447 (N_17447,N_16684,N_16669);
nand U17448 (N_17448,N_16926,N_16891);
nor U17449 (N_17449,N_16912,N_16913);
xor U17450 (N_17450,N_16754,N_16694);
nor U17451 (N_17451,N_16724,N_16915);
nand U17452 (N_17452,N_16996,N_16846);
and U17453 (N_17453,N_16983,N_16574);
nor U17454 (N_17454,N_16641,N_16987);
or U17455 (N_17455,N_16777,N_16808);
or U17456 (N_17456,N_16825,N_16878);
or U17457 (N_17457,N_16637,N_16908);
or U17458 (N_17458,N_16976,N_16931);
and U17459 (N_17459,N_16666,N_16550);
and U17460 (N_17460,N_16735,N_16636);
xnor U17461 (N_17461,N_16613,N_16911);
xor U17462 (N_17462,N_16764,N_16945);
nor U17463 (N_17463,N_16942,N_16687);
or U17464 (N_17464,N_16864,N_16584);
and U17465 (N_17465,N_16989,N_16742);
nand U17466 (N_17466,N_16668,N_16679);
xor U17467 (N_17467,N_16580,N_16771);
or U17468 (N_17468,N_16907,N_16676);
or U17469 (N_17469,N_16875,N_16861);
nand U17470 (N_17470,N_16757,N_16532);
or U17471 (N_17471,N_16539,N_16670);
nor U17472 (N_17472,N_16553,N_16709);
nor U17473 (N_17473,N_16637,N_16645);
xnor U17474 (N_17474,N_16912,N_16836);
nor U17475 (N_17475,N_16636,N_16773);
or U17476 (N_17476,N_16532,N_16578);
nand U17477 (N_17477,N_16776,N_16621);
nor U17478 (N_17478,N_16868,N_16899);
or U17479 (N_17479,N_16926,N_16810);
and U17480 (N_17480,N_16894,N_16701);
or U17481 (N_17481,N_16894,N_16655);
nand U17482 (N_17482,N_16886,N_16521);
nand U17483 (N_17483,N_16920,N_16985);
and U17484 (N_17484,N_16614,N_16797);
nor U17485 (N_17485,N_16925,N_16526);
nand U17486 (N_17486,N_16957,N_16579);
xor U17487 (N_17487,N_16769,N_16843);
nand U17488 (N_17488,N_16823,N_16952);
and U17489 (N_17489,N_16683,N_16606);
xnor U17490 (N_17490,N_16986,N_16783);
and U17491 (N_17491,N_16718,N_16762);
nand U17492 (N_17492,N_16700,N_16801);
and U17493 (N_17493,N_16940,N_16578);
nor U17494 (N_17494,N_16943,N_16638);
nor U17495 (N_17495,N_16900,N_16638);
or U17496 (N_17496,N_16620,N_16503);
xnor U17497 (N_17497,N_16788,N_16648);
nand U17498 (N_17498,N_16988,N_16562);
or U17499 (N_17499,N_16861,N_16900);
nand U17500 (N_17500,N_17481,N_17443);
and U17501 (N_17501,N_17151,N_17104);
xnor U17502 (N_17502,N_17262,N_17438);
nor U17503 (N_17503,N_17233,N_17274);
and U17504 (N_17504,N_17480,N_17075);
nor U17505 (N_17505,N_17276,N_17291);
nor U17506 (N_17506,N_17257,N_17137);
xnor U17507 (N_17507,N_17147,N_17367);
nand U17508 (N_17508,N_17413,N_17471);
xnor U17509 (N_17509,N_17298,N_17074);
or U17510 (N_17510,N_17103,N_17477);
and U17511 (N_17511,N_17199,N_17008);
nand U17512 (N_17512,N_17178,N_17204);
and U17513 (N_17513,N_17122,N_17430);
and U17514 (N_17514,N_17183,N_17111);
and U17515 (N_17515,N_17217,N_17045);
xor U17516 (N_17516,N_17282,N_17088);
or U17517 (N_17517,N_17302,N_17351);
and U17518 (N_17518,N_17231,N_17492);
nand U17519 (N_17519,N_17190,N_17416);
nand U17520 (N_17520,N_17304,N_17154);
nand U17521 (N_17521,N_17335,N_17308);
xor U17522 (N_17522,N_17398,N_17431);
or U17523 (N_17523,N_17358,N_17319);
xnor U17524 (N_17524,N_17401,N_17148);
xor U17525 (N_17525,N_17346,N_17166);
xor U17526 (N_17526,N_17489,N_17258);
or U17527 (N_17527,N_17391,N_17465);
or U17528 (N_17528,N_17460,N_17037);
and U17529 (N_17529,N_17420,N_17429);
nand U17530 (N_17530,N_17264,N_17110);
xnor U17531 (N_17531,N_17113,N_17141);
or U17532 (N_17532,N_17452,N_17249);
or U17533 (N_17533,N_17330,N_17458);
xnor U17534 (N_17534,N_17027,N_17377);
nor U17535 (N_17535,N_17168,N_17162);
and U17536 (N_17536,N_17035,N_17055);
nand U17537 (N_17537,N_17207,N_17225);
or U17538 (N_17538,N_17371,N_17094);
xnor U17539 (N_17539,N_17373,N_17004);
xor U17540 (N_17540,N_17397,N_17063);
nand U17541 (N_17541,N_17089,N_17140);
nand U17542 (N_17542,N_17428,N_17191);
nor U17543 (N_17543,N_17261,N_17100);
and U17544 (N_17544,N_17213,N_17488);
and U17545 (N_17545,N_17219,N_17405);
nand U17546 (N_17546,N_17131,N_17186);
xnor U17547 (N_17547,N_17201,N_17378);
nor U17548 (N_17548,N_17365,N_17222);
nor U17549 (N_17549,N_17357,N_17423);
nand U17550 (N_17550,N_17019,N_17467);
xor U17551 (N_17551,N_17279,N_17014);
or U17552 (N_17552,N_17386,N_17145);
or U17553 (N_17553,N_17206,N_17172);
nand U17554 (N_17554,N_17252,N_17155);
nand U17555 (N_17555,N_17384,N_17390);
nand U17556 (N_17556,N_17067,N_17447);
nor U17557 (N_17557,N_17498,N_17192);
xor U17558 (N_17558,N_17434,N_17046);
or U17559 (N_17559,N_17372,N_17494);
and U17560 (N_17560,N_17181,N_17404);
xnor U17561 (N_17561,N_17226,N_17294);
or U17562 (N_17562,N_17086,N_17189);
xnor U17563 (N_17563,N_17196,N_17093);
and U17564 (N_17564,N_17385,N_17193);
xnor U17565 (N_17565,N_17180,N_17101);
nor U17566 (N_17566,N_17028,N_17096);
xor U17567 (N_17567,N_17248,N_17472);
xor U17568 (N_17568,N_17476,N_17057);
and U17569 (N_17569,N_17305,N_17059);
xnor U17570 (N_17570,N_17126,N_17129);
and U17571 (N_17571,N_17116,N_17095);
and U17572 (N_17572,N_17068,N_17102);
nor U17573 (N_17573,N_17177,N_17278);
xor U17574 (N_17574,N_17353,N_17070);
xor U17575 (N_17575,N_17297,N_17215);
xor U17576 (N_17576,N_17444,N_17237);
nand U17577 (N_17577,N_17013,N_17083);
xor U17578 (N_17578,N_17127,N_17295);
and U17579 (N_17579,N_17345,N_17221);
or U17580 (N_17580,N_17311,N_17451);
nand U17581 (N_17581,N_17486,N_17018);
nor U17582 (N_17582,N_17149,N_17240);
nand U17583 (N_17583,N_17034,N_17023);
and U17584 (N_17584,N_17200,N_17253);
or U17585 (N_17585,N_17119,N_17422);
nand U17586 (N_17586,N_17016,N_17382);
nor U17587 (N_17587,N_17009,N_17256);
nand U17588 (N_17588,N_17331,N_17164);
nand U17589 (N_17589,N_17203,N_17156);
nor U17590 (N_17590,N_17383,N_17473);
and U17591 (N_17591,N_17033,N_17343);
nor U17592 (N_17592,N_17024,N_17188);
xor U17593 (N_17593,N_17315,N_17107);
or U17594 (N_17594,N_17159,N_17364);
xnor U17595 (N_17595,N_17267,N_17321);
or U17596 (N_17596,N_17130,N_17006);
and U17597 (N_17597,N_17493,N_17121);
and U17598 (N_17598,N_17388,N_17112);
or U17599 (N_17599,N_17133,N_17146);
nand U17600 (N_17600,N_17449,N_17454);
and U17601 (N_17601,N_17029,N_17326);
xor U17602 (N_17602,N_17069,N_17436);
xor U17603 (N_17603,N_17470,N_17314);
nor U17604 (N_17604,N_17407,N_17427);
or U17605 (N_17605,N_17300,N_17051);
and U17606 (N_17606,N_17469,N_17475);
and U17607 (N_17607,N_17496,N_17411);
and U17608 (N_17608,N_17117,N_17079);
nor U17609 (N_17609,N_17169,N_17468);
nand U17610 (N_17610,N_17393,N_17165);
or U17611 (N_17611,N_17138,N_17446);
and U17612 (N_17612,N_17344,N_17058);
or U17613 (N_17613,N_17123,N_17182);
nor U17614 (N_17614,N_17439,N_17150);
or U17615 (N_17615,N_17032,N_17241);
or U17616 (N_17616,N_17339,N_17340);
or U17617 (N_17617,N_17318,N_17323);
or U17618 (N_17618,N_17433,N_17195);
and U17619 (N_17619,N_17002,N_17060);
and U17620 (N_17620,N_17224,N_17084);
or U17621 (N_17621,N_17463,N_17479);
or U17622 (N_17622,N_17399,N_17010);
nor U17623 (N_17623,N_17332,N_17462);
or U17624 (N_17624,N_17238,N_17409);
xnor U17625 (N_17625,N_17160,N_17026);
nor U17626 (N_17626,N_17350,N_17174);
or U17627 (N_17627,N_17142,N_17324);
nand U17628 (N_17628,N_17355,N_17333);
nor U17629 (N_17629,N_17485,N_17242);
xnor U17630 (N_17630,N_17025,N_17374);
nand U17631 (N_17631,N_17260,N_17320);
nor U17632 (N_17632,N_17263,N_17270);
nor U17633 (N_17633,N_17495,N_17266);
and U17634 (N_17634,N_17289,N_17005);
or U17635 (N_17635,N_17301,N_17272);
nor U17636 (N_17636,N_17359,N_17061);
nor U17637 (N_17637,N_17049,N_17212);
xnor U17638 (N_17638,N_17312,N_17209);
nand U17639 (N_17639,N_17342,N_17497);
and U17640 (N_17640,N_17456,N_17062);
or U17641 (N_17641,N_17361,N_17073);
nand U17642 (N_17642,N_17232,N_17487);
nand U17643 (N_17643,N_17031,N_17329);
nand U17644 (N_17644,N_17293,N_17236);
xnor U17645 (N_17645,N_17021,N_17442);
xnor U17646 (N_17646,N_17082,N_17464);
or U17647 (N_17647,N_17490,N_17072);
nor U17648 (N_17648,N_17099,N_17402);
nor U17649 (N_17649,N_17098,N_17280);
or U17650 (N_17650,N_17426,N_17482);
and U17651 (N_17651,N_17039,N_17296);
and U17652 (N_17652,N_17003,N_17017);
nand U17653 (N_17653,N_17125,N_17341);
nor U17654 (N_17654,N_17153,N_17227);
and U17655 (N_17655,N_17457,N_17408);
and U17656 (N_17656,N_17114,N_17375);
nor U17657 (N_17657,N_17175,N_17400);
and U17658 (N_17658,N_17491,N_17415);
nand U17659 (N_17659,N_17106,N_17327);
nor U17660 (N_17660,N_17223,N_17396);
nand U17661 (N_17661,N_17136,N_17229);
and U17662 (N_17662,N_17307,N_17007);
nor U17663 (N_17663,N_17414,N_17239);
nor U17664 (N_17664,N_17303,N_17387);
nand U17665 (N_17665,N_17380,N_17313);
nor U17666 (N_17666,N_17370,N_17265);
xnor U17667 (N_17667,N_17243,N_17379);
xor U17668 (N_17668,N_17255,N_17424);
xnor U17669 (N_17669,N_17080,N_17432);
xor U17670 (N_17670,N_17078,N_17115);
xnor U17671 (N_17671,N_17064,N_17211);
nand U17672 (N_17672,N_17336,N_17254);
nand U17673 (N_17673,N_17179,N_17418);
nand U17674 (N_17674,N_17288,N_17198);
xor U17675 (N_17675,N_17216,N_17050);
or U17676 (N_17676,N_17246,N_17362);
or U17677 (N_17677,N_17325,N_17389);
and U17678 (N_17678,N_17085,N_17269);
or U17679 (N_17679,N_17417,N_17478);
xor U17680 (N_17680,N_17283,N_17205);
and U17681 (N_17681,N_17077,N_17020);
and U17682 (N_17682,N_17306,N_17425);
and U17683 (N_17683,N_17435,N_17310);
xnor U17684 (N_17684,N_17048,N_17437);
nor U17685 (N_17685,N_17286,N_17381);
and U17686 (N_17686,N_17419,N_17171);
and U17687 (N_17687,N_17087,N_17030);
or U17688 (N_17688,N_17152,N_17356);
nor U17689 (N_17689,N_17292,N_17337);
or U17690 (N_17690,N_17392,N_17052);
and U17691 (N_17691,N_17076,N_17163);
and U17692 (N_17692,N_17316,N_17139);
nor U17693 (N_17693,N_17036,N_17053);
and U17694 (N_17694,N_17474,N_17167);
xor U17695 (N_17695,N_17285,N_17144);
and U17696 (N_17696,N_17124,N_17228);
xnor U17697 (N_17697,N_17054,N_17170);
xor U17698 (N_17698,N_17368,N_17208);
xor U17699 (N_17699,N_17275,N_17176);
nand U17700 (N_17700,N_17247,N_17056);
nand U17701 (N_17701,N_17230,N_17015);
nor U17702 (N_17702,N_17044,N_17348);
or U17703 (N_17703,N_17347,N_17218);
and U17704 (N_17704,N_17455,N_17338);
and U17705 (N_17705,N_17309,N_17065);
nor U17706 (N_17706,N_17042,N_17376);
xnor U17707 (N_17707,N_17459,N_17290);
xnor U17708 (N_17708,N_17421,N_17011);
and U17709 (N_17709,N_17081,N_17499);
and U17710 (N_17710,N_17202,N_17299);
and U17711 (N_17711,N_17360,N_17484);
or U17712 (N_17712,N_17038,N_17041);
and U17713 (N_17713,N_17363,N_17128);
and U17714 (N_17714,N_17047,N_17105);
xor U17715 (N_17715,N_17109,N_17092);
nor U17716 (N_17716,N_17161,N_17354);
nor U17717 (N_17717,N_17284,N_17158);
or U17718 (N_17718,N_17194,N_17322);
and U17719 (N_17719,N_17235,N_17157);
nand U17720 (N_17720,N_17453,N_17268);
xor U17721 (N_17721,N_17250,N_17234);
and U17722 (N_17722,N_17097,N_17173);
nand U17723 (N_17723,N_17352,N_17001);
nand U17724 (N_17724,N_17412,N_17184);
xor U17725 (N_17725,N_17394,N_17108);
nor U17726 (N_17726,N_17187,N_17328);
nand U17727 (N_17727,N_17271,N_17210);
nor U17728 (N_17728,N_17118,N_17040);
or U17729 (N_17729,N_17448,N_17369);
nor U17730 (N_17730,N_17012,N_17132);
and U17731 (N_17731,N_17244,N_17277);
nor U17732 (N_17732,N_17466,N_17134);
or U17733 (N_17733,N_17441,N_17273);
nand U17734 (N_17734,N_17483,N_17251);
nor U17735 (N_17735,N_17022,N_17066);
nor U17736 (N_17736,N_17445,N_17281);
nor U17737 (N_17737,N_17185,N_17000);
nor U17738 (N_17738,N_17287,N_17403);
nand U17739 (N_17739,N_17259,N_17450);
xor U17740 (N_17740,N_17090,N_17440);
or U17741 (N_17741,N_17406,N_17120);
and U17742 (N_17742,N_17091,N_17143);
or U17743 (N_17743,N_17395,N_17349);
or U17744 (N_17744,N_17317,N_17410);
nor U17745 (N_17745,N_17220,N_17043);
nand U17746 (N_17746,N_17366,N_17245);
or U17747 (N_17747,N_17461,N_17214);
and U17748 (N_17748,N_17135,N_17334);
or U17749 (N_17749,N_17197,N_17071);
xor U17750 (N_17750,N_17124,N_17494);
nand U17751 (N_17751,N_17201,N_17298);
and U17752 (N_17752,N_17098,N_17130);
or U17753 (N_17753,N_17405,N_17307);
xor U17754 (N_17754,N_17415,N_17100);
xor U17755 (N_17755,N_17436,N_17402);
nand U17756 (N_17756,N_17481,N_17270);
or U17757 (N_17757,N_17430,N_17296);
nor U17758 (N_17758,N_17372,N_17317);
or U17759 (N_17759,N_17194,N_17331);
and U17760 (N_17760,N_17373,N_17007);
nor U17761 (N_17761,N_17140,N_17003);
xor U17762 (N_17762,N_17243,N_17112);
xnor U17763 (N_17763,N_17098,N_17228);
nand U17764 (N_17764,N_17170,N_17033);
nor U17765 (N_17765,N_17007,N_17305);
nor U17766 (N_17766,N_17361,N_17013);
nor U17767 (N_17767,N_17064,N_17282);
or U17768 (N_17768,N_17311,N_17126);
nor U17769 (N_17769,N_17281,N_17315);
xnor U17770 (N_17770,N_17477,N_17381);
xor U17771 (N_17771,N_17033,N_17236);
xor U17772 (N_17772,N_17430,N_17102);
nand U17773 (N_17773,N_17145,N_17186);
or U17774 (N_17774,N_17052,N_17025);
and U17775 (N_17775,N_17428,N_17427);
and U17776 (N_17776,N_17227,N_17231);
xor U17777 (N_17777,N_17027,N_17182);
xor U17778 (N_17778,N_17253,N_17149);
and U17779 (N_17779,N_17472,N_17214);
or U17780 (N_17780,N_17249,N_17114);
or U17781 (N_17781,N_17049,N_17170);
or U17782 (N_17782,N_17196,N_17065);
nor U17783 (N_17783,N_17335,N_17068);
xnor U17784 (N_17784,N_17437,N_17447);
nor U17785 (N_17785,N_17308,N_17314);
xnor U17786 (N_17786,N_17216,N_17447);
or U17787 (N_17787,N_17043,N_17335);
or U17788 (N_17788,N_17355,N_17074);
nand U17789 (N_17789,N_17223,N_17020);
and U17790 (N_17790,N_17410,N_17395);
xor U17791 (N_17791,N_17359,N_17204);
and U17792 (N_17792,N_17246,N_17226);
or U17793 (N_17793,N_17179,N_17493);
and U17794 (N_17794,N_17108,N_17068);
nor U17795 (N_17795,N_17384,N_17240);
and U17796 (N_17796,N_17324,N_17179);
or U17797 (N_17797,N_17148,N_17384);
xnor U17798 (N_17798,N_17477,N_17438);
xor U17799 (N_17799,N_17254,N_17228);
and U17800 (N_17800,N_17494,N_17362);
or U17801 (N_17801,N_17305,N_17123);
xor U17802 (N_17802,N_17474,N_17312);
nor U17803 (N_17803,N_17290,N_17055);
xor U17804 (N_17804,N_17087,N_17375);
xnor U17805 (N_17805,N_17205,N_17219);
xor U17806 (N_17806,N_17001,N_17155);
or U17807 (N_17807,N_17448,N_17370);
nor U17808 (N_17808,N_17120,N_17133);
or U17809 (N_17809,N_17413,N_17445);
nor U17810 (N_17810,N_17195,N_17036);
nand U17811 (N_17811,N_17193,N_17128);
or U17812 (N_17812,N_17256,N_17260);
and U17813 (N_17813,N_17031,N_17387);
nor U17814 (N_17814,N_17202,N_17115);
nor U17815 (N_17815,N_17098,N_17033);
nand U17816 (N_17816,N_17221,N_17141);
nand U17817 (N_17817,N_17117,N_17445);
xnor U17818 (N_17818,N_17172,N_17280);
xnor U17819 (N_17819,N_17015,N_17009);
xnor U17820 (N_17820,N_17414,N_17270);
nand U17821 (N_17821,N_17414,N_17395);
or U17822 (N_17822,N_17307,N_17216);
nor U17823 (N_17823,N_17133,N_17491);
nor U17824 (N_17824,N_17066,N_17062);
and U17825 (N_17825,N_17395,N_17208);
nand U17826 (N_17826,N_17151,N_17001);
nand U17827 (N_17827,N_17483,N_17157);
or U17828 (N_17828,N_17040,N_17456);
xor U17829 (N_17829,N_17221,N_17200);
nor U17830 (N_17830,N_17311,N_17355);
xnor U17831 (N_17831,N_17315,N_17008);
or U17832 (N_17832,N_17450,N_17363);
nand U17833 (N_17833,N_17199,N_17091);
and U17834 (N_17834,N_17245,N_17140);
and U17835 (N_17835,N_17269,N_17152);
nand U17836 (N_17836,N_17399,N_17038);
and U17837 (N_17837,N_17220,N_17122);
xor U17838 (N_17838,N_17029,N_17090);
nand U17839 (N_17839,N_17459,N_17256);
nor U17840 (N_17840,N_17301,N_17056);
xnor U17841 (N_17841,N_17287,N_17272);
or U17842 (N_17842,N_17279,N_17254);
or U17843 (N_17843,N_17048,N_17486);
nand U17844 (N_17844,N_17306,N_17111);
nor U17845 (N_17845,N_17287,N_17362);
xor U17846 (N_17846,N_17077,N_17309);
and U17847 (N_17847,N_17358,N_17024);
and U17848 (N_17848,N_17067,N_17377);
xor U17849 (N_17849,N_17200,N_17070);
nor U17850 (N_17850,N_17378,N_17315);
nand U17851 (N_17851,N_17160,N_17046);
and U17852 (N_17852,N_17391,N_17151);
xnor U17853 (N_17853,N_17360,N_17351);
or U17854 (N_17854,N_17278,N_17246);
or U17855 (N_17855,N_17027,N_17491);
or U17856 (N_17856,N_17399,N_17476);
nor U17857 (N_17857,N_17421,N_17026);
xnor U17858 (N_17858,N_17376,N_17494);
or U17859 (N_17859,N_17123,N_17188);
or U17860 (N_17860,N_17177,N_17130);
xnor U17861 (N_17861,N_17024,N_17032);
nor U17862 (N_17862,N_17303,N_17238);
and U17863 (N_17863,N_17014,N_17182);
or U17864 (N_17864,N_17280,N_17194);
and U17865 (N_17865,N_17480,N_17490);
nor U17866 (N_17866,N_17469,N_17385);
or U17867 (N_17867,N_17152,N_17354);
xnor U17868 (N_17868,N_17127,N_17342);
xor U17869 (N_17869,N_17464,N_17332);
nor U17870 (N_17870,N_17259,N_17385);
xnor U17871 (N_17871,N_17269,N_17123);
or U17872 (N_17872,N_17288,N_17414);
nand U17873 (N_17873,N_17312,N_17236);
nand U17874 (N_17874,N_17073,N_17327);
nand U17875 (N_17875,N_17169,N_17321);
nand U17876 (N_17876,N_17321,N_17117);
xor U17877 (N_17877,N_17255,N_17137);
xor U17878 (N_17878,N_17344,N_17082);
xor U17879 (N_17879,N_17399,N_17344);
or U17880 (N_17880,N_17467,N_17126);
xnor U17881 (N_17881,N_17466,N_17188);
nor U17882 (N_17882,N_17247,N_17321);
or U17883 (N_17883,N_17254,N_17004);
and U17884 (N_17884,N_17062,N_17105);
nor U17885 (N_17885,N_17098,N_17066);
nor U17886 (N_17886,N_17359,N_17257);
or U17887 (N_17887,N_17390,N_17108);
or U17888 (N_17888,N_17267,N_17246);
xnor U17889 (N_17889,N_17353,N_17208);
xnor U17890 (N_17890,N_17171,N_17376);
and U17891 (N_17891,N_17453,N_17324);
and U17892 (N_17892,N_17485,N_17353);
or U17893 (N_17893,N_17461,N_17492);
or U17894 (N_17894,N_17390,N_17073);
and U17895 (N_17895,N_17155,N_17137);
nor U17896 (N_17896,N_17424,N_17452);
nand U17897 (N_17897,N_17374,N_17085);
or U17898 (N_17898,N_17414,N_17012);
or U17899 (N_17899,N_17020,N_17447);
xor U17900 (N_17900,N_17017,N_17214);
or U17901 (N_17901,N_17385,N_17415);
or U17902 (N_17902,N_17229,N_17470);
nor U17903 (N_17903,N_17096,N_17153);
or U17904 (N_17904,N_17373,N_17453);
or U17905 (N_17905,N_17155,N_17432);
nand U17906 (N_17906,N_17043,N_17222);
nor U17907 (N_17907,N_17138,N_17030);
xnor U17908 (N_17908,N_17194,N_17262);
nor U17909 (N_17909,N_17335,N_17054);
or U17910 (N_17910,N_17360,N_17100);
and U17911 (N_17911,N_17425,N_17011);
and U17912 (N_17912,N_17068,N_17306);
or U17913 (N_17913,N_17373,N_17496);
and U17914 (N_17914,N_17447,N_17038);
nor U17915 (N_17915,N_17220,N_17162);
xor U17916 (N_17916,N_17183,N_17458);
nand U17917 (N_17917,N_17248,N_17312);
and U17918 (N_17918,N_17253,N_17289);
and U17919 (N_17919,N_17493,N_17434);
xnor U17920 (N_17920,N_17401,N_17080);
or U17921 (N_17921,N_17473,N_17054);
or U17922 (N_17922,N_17435,N_17099);
nor U17923 (N_17923,N_17220,N_17225);
or U17924 (N_17924,N_17361,N_17024);
or U17925 (N_17925,N_17414,N_17312);
nor U17926 (N_17926,N_17109,N_17330);
xnor U17927 (N_17927,N_17416,N_17182);
and U17928 (N_17928,N_17304,N_17243);
or U17929 (N_17929,N_17137,N_17344);
nor U17930 (N_17930,N_17327,N_17090);
or U17931 (N_17931,N_17473,N_17093);
nand U17932 (N_17932,N_17290,N_17357);
xor U17933 (N_17933,N_17200,N_17056);
nor U17934 (N_17934,N_17253,N_17060);
nand U17935 (N_17935,N_17269,N_17405);
or U17936 (N_17936,N_17150,N_17129);
xor U17937 (N_17937,N_17117,N_17372);
nand U17938 (N_17938,N_17074,N_17454);
or U17939 (N_17939,N_17441,N_17247);
nand U17940 (N_17940,N_17367,N_17230);
and U17941 (N_17941,N_17070,N_17143);
or U17942 (N_17942,N_17355,N_17192);
xnor U17943 (N_17943,N_17288,N_17305);
and U17944 (N_17944,N_17052,N_17189);
nor U17945 (N_17945,N_17387,N_17007);
nor U17946 (N_17946,N_17288,N_17366);
nand U17947 (N_17947,N_17304,N_17351);
nand U17948 (N_17948,N_17032,N_17294);
xnor U17949 (N_17949,N_17280,N_17339);
nand U17950 (N_17950,N_17370,N_17407);
nand U17951 (N_17951,N_17272,N_17340);
and U17952 (N_17952,N_17431,N_17251);
nor U17953 (N_17953,N_17071,N_17431);
and U17954 (N_17954,N_17290,N_17020);
xor U17955 (N_17955,N_17004,N_17435);
or U17956 (N_17956,N_17318,N_17344);
nor U17957 (N_17957,N_17034,N_17485);
nor U17958 (N_17958,N_17121,N_17090);
xnor U17959 (N_17959,N_17321,N_17153);
or U17960 (N_17960,N_17454,N_17128);
nor U17961 (N_17961,N_17311,N_17204);
and U17962 (N_17962,N_17188,N_17491);
xnor U17963 (N_17963,N_17114,N_17284);
nor U17964 (N_17964,N_17160,N_17075);
and U17965 (N_17965,N_17051,N_17199);
or U17966 (N_17966,N_17000,N_17403);
nor U17967 (N_17967,N_17296,N_17467);
or U17968 (N_17968,N_17419,N_17360);
nor U17969 (N_17969,N_17350,N_17221);
and U17970 (N_17970,N_17325,N_17329);
or U17971 (N_17971,N_17243,N_17350);
nand U17972 (N_17972,N_17098,N_17387);
or U17973 (N_17973,N_17202,N_17024);
nor U17974 (N_17974,N_17432,N_17091);
nor U17975 (N_17975,N_17086,N_17152);
nand U17976 (N_17976,N_17311,N_17461);
nand U17977 (N_17977,N_17300,N_17329);
or U17978 (N_17978,N_17184,N_17352);
nor U17979 (N_17979,N_17450,N_17331);
and U17980 (N_17980,N_17487,N_17480);
or U17981 (N_17981,N_17248,N_17053);
xor U17982 (N_17982,N_17063,N_17303);
or U17983 (N_17983,N_17429,N_17168);
xnor U17984 (N_17984,N_17010,N_17385);
xnor U17985 (N_17985,N_17437,N_17191);
nand U17986 (N_17986,N_17486,N_17212);
nand U17987 (N_17987,N_17047,N_17336);
and U17988 (N_17988,N_17324,N_17410);
nor U17989 (N_17989,N_17052,N_17215);
nand U17990 (N_17990,N_17469,N_17190);
and U17991 (N_17991,N_17127,N_17260);
nor U17992 (N_17992,N_17156,N_17278);
and U17993 (N_17993,N_17201,N_17322);
nor U17994 (N_17994,N_17166,N_17193);
or U17995 (N_17995,N_17279,N_17087);
and U17996 (N_17996,N_17299,N_17137);
or U17997 (N_17997,N_17470,N_17359);
nor U17998 (N_17998,N_17268,N_17315);
or U17999 (N_17999,N_17276,N_17337);
and U18000 (N_18000,N_17894,N_17559);
and U18001 (N_18001,N_17917,N_17954);
nor U18002 (N_18002,N_17803,N_17527);
nand U18003 (N_18003,N_17617,N_17735);
xnor U18004 (N_18004,N_17883,N_17529);
and U18005 (N_18005,N_17530,N_17567);
nor U18006 (N_18006,N_17967,N_17950);
nor U18007 (N_18007,N_17522,N_17924);
and U18008 (N_18008,N_17711,N_17584);
xor U18009 (N_18009,N_17692,N_17948);
and U18010 (N_18010,N_17781,N_17551);
xor U18011 (N_18011,N_17818,N_17916);
nand U18012 (N_18012,N_17832,N_17969);
or U18013 (N_18013,N_17676,N_17675);
nor U18014 (N_18014,N_17784,N_17525);
or U18015 (N_18015,N_17820,N_17819);
nand U18016 (N_18016,N_17877,N_17626);
and U18017 (N_18017,N_17972,N_17662);
xor U18018 (N_18018,N_17956,N_17573);
xnor U18019 (N_18019,N_17758,N_17729);
nor U18020 (N_18020,N_17879,N_17629);
or U18021 (N_18021,N_17881,N_17787);
or U18022 (N_18022,N_17862,N_17989);
xnor U18023 (N_18023,N_17762,N_17724);
nand U18024 (N_18024,N_17851,N_17838);
and U18025 (N_18025,N_17607,N_17856);
nand U18026 (N_18026,N_17641,N_17586);
or U18027 (N_18027,N_17930,N_17760);
nand U18028 (N_18028,N_17911,N_17943);
and U18029 (N_18029,N_17857,N_17926);
nand U18030 (N_18030,N_17970,N_17783);
or U18031 (N_18031,N_17807,N_17557);
nand U18032 (N_18032,N_17562,N_17793);
xor U18033 (N_18033,N_17898,N_17827);
or U18034 (N_18034,N_17799,N_17550);
or U18035 (N_18035,N_17778,N_17652);
and U18036 (N_18036,N_17690,N_17825);
xnor U18037 (N_18037,N_17875,N_17891);
nor U18038 (N_18038,N_17951,N_17768);
and U18039 (N_18039,N_17661,N_17619);
nor U18040 (N_18040,N_17686,N_17983);
xor U18041 (N_18041,N_17854,N_17830);
xnor U18042 (N_18042,N_17625,N_17804);
nand U18043 (N_18043,N_17998,N_17543);
nor U18044 (N_18044,N_17897,N_17882);
or U18045 (N_18045,N_17821,N_17971);
nor U18046 (N_18046,N_17654,N_17893);
and U18047 (N_18047,N_17860,N_17791);
xor U18048 (N_18048,N_17955,N_17816);
xnor U18049 (N_18049,N_17975,N_17552);
nand U18050 (N_18050,N_17836,N_17513);
xor U18051 (N_18051,N_17831,N_17802);
and U18052 (N_18052,N_17865,N_17814);
nand U18053 (N_18053,N_17742,N_17558);
xnor U18054 (N_18054,N_17707,N_17623);
and U18055 (N_18055,N_17517,N_17611);
nor U18056 (N_18056,N_17702,N_17889);
nor U18057 (N_18057,N_17769,N_17963);
nand U18058 (N_18058,N_17608,N_17540);
xor U18059 (N_18059,N_17582,N_17642);
xor U18060 (N_18060,N_17866,N_17852);
nor U18061 (N_18061,N_17553,N_17904);
nand U18062 (N_18062,N_17655,N_17776);
nand U18063 (N_18063,N_17792,N_17789);
and U18064 (N_18064,N_17620,N_17964);
xor U18065 (N_18065,N_17687,N_17937);
and U18066 (N_18066,N_17940,N_17502);
xor U18067 (N_18067,N_17671,N_17660);
or U18068 (N_18068,N_17621,N_17603);
xnor U18069 (N_18069,N_17828,N_17706);
nand U18070 (N_18070,N_17849,N_17845);
nand U18071 (N_18071,N_17752,N_17941);
nand U18072 (N_18072,N_17563,N_17780);
nand U18073 (N_18073,N_17512,N_17679);
nor U18074 (N_18074,N_17734,N_17848);
nand U18075 (N_18075,N_17756,N_17506);
nor U18076 (N_18076,N_17744,N_17733);
or U18077 (N_18077,N_17839,N_17537);
and U18078 (N_18078,N_17986,N_17880);
nand U18079 (N_18079,N_17805,N_17531);
or U18080 (N_18080,N_17913,N_17561);
and U18081 (N_18081,N_17746,N_17566);
or U18082 (N_18082,N_17523,N_17764);
and U18083 (N_18083,N_17631,N_17919);
nor U18084 (N_18084,N_17666,N_17901);
nor U18085 (N_18085,N_17927,N_17934);
or U18086 (N_18086,N_17959,N_17598);
nand U18087 (N_18087,N_17507,N_17942);
and U18088 (N_18088,N_17736,N_17601);
nand U18089 (N_18089,N_17981,N_17922);
or U18090 (N_18090,N_17988,N_17790);
nand U18091 (N_18091,N_17578,N_17596);
or U18092 (N_18092,N_17520,N_17731);
nor U18093 (N_18093,N_17824,N_17571);
nor U18094 (N_18094,N_17508,N_17524);
nand U18095 (N_18095,N_17536,N_17696);
nor U18096 (N_18096,N_17976,N_17580);
and U18097 (N_18097,N_17777,N_17886);
nand U18098 (N_18098,N_17713,N_17750);
and U18099 (N_18099,N_17800,N_17723);
and U18100 (N_18100,N_17868,N_17797);
xor U18101 (N_18101,N_17811,N_17704);
or U18102 (N_18102,N_17929,N_17771);
nor U18103 (N_18103,N_17627,N_17590);
and U18104 (N_18104,N_17624,N_17946);
nor U18105 (N_18105,N_17863,N_17699);
or U18106 (N_18106,N_17535,N_17688);
and U18107 (N_18107,N_17812,N_17635);
nor U18108 (N_18108,N_17949,N_17726);
and U18109 (N_18109,N_17872,N_17546);
nand U18110 (N_18110,N_17966,N_17847);
and U18111 (N_18111,N_17589,N_17648);
nor U18112 (N_18112,N_17905,N_17766);
or U18113 (N_18113,N_17705,N_17544);
or U18114 (N_18114,N_17952,N_17869);
nor U18115 (N_18115,N_17759,N_17593);
nand U18116 (N_18116,N_17931,N_17606);
or U18117 (N_18117,N_17511,N_17521);
nand U18118 (N_18118,N_17801,N_17870);
and U18119 (N_18119,N_17815,N_17681);
and U18120 (N_18120,N_17638,N_17576);
nor U18121 (N_18121,N_17810,N_17984);
and U18122 (N_18122,N_17817,N_17616);
or U18123 (N_18123,N_17920,N_17565);
nor U18124 (N_18124,N_17747,N_17961);
and U18125 (N_18125,N_17906,N_17813);
nor U18126 (N_18126,N_17605,N_17604);
nor U18127 (N_18127,N_17665,N_17855);
xnor U18128 (N_18128,N_17575,N_17570);
nor U18129 (N_18129,N_17719,N_17829);
nor U18130 (N_18130,N_17910,N_17737);
nand U18131 (N_18131,N_17858,N_17700);
nand U18132 (N_18132,N_17718,N_17651);
or U18133 (N_18133,N_17895,N_17588);
nor U18134 (N_18134,N_17613,N_17569);
xor U18135 (N_18135,N_17892,N_17549);
or U18136 (N_18136,N_17915,N_17592);
xnor U18137 (N_18137,N_17936,N_17918);
xor U18138 (N_18138,N_17533,N_17809);
xor U18139 (N_18139,N_17614,N_17795);
xor U18140 (N_18140,N_17510,N_17646);
and U18141 (N_18141,N_17509,N_17663);
nor U18142 (N_18142,N_17987,N_17636);
and U18143 (N_18143,N_17712,N_17632);
and U18144 (N_18144,N_17767,N_17547);
nand U18145 (N_18145,N_17622,N_17977);
xor U18146 (N_18146,N_17722,N_17748);
nor U18147 (N_18147,N_17995,N_17628);
nand U18148 (N_18148,N_17779,N_17526);
xor U18149 (N_18149,N_17844,N_17841);
nand U18150 (N_18150,N_17907,N_17864);
xor U18151 (N_18151,N_17680,N_17554);
xnor U18152 (N_18152,N_17775,N_17720);
and U18153 (N_18153,N_17515,N_17861);
and U18154 (N_18154,N_17714,N_17504);
nand U18155 (N_18155,N_17965,N_17878);
xor U18156 (N_18156,N_17600,N_17501);
nand U18157 (N_18157,N_17572,N_17514);
nor U18158 (N_18158,N_17754,N_17739);
nand U18159 (N_18159,N_17698,N_17682);
and U18160 (N_18160,N_17826,N_17785);
and U18161 (N_18161,N_17822,N_17990);
or U18162 (N_18162,N_17677,N_17833);
xnor U18163 (N_18163,N_17564,N_17568);
nor U18164 (N_18164,N_17673,N_17903);
and U18165 (N_18165,N_17957,N_17656);
or U18166 (N_18166,N_17630,N_17500);
xor U18167 (N_18167,N_17843,N_17958);
or U18168 (N_18168,N_17867,N_17982);
xor U18169 (N_18169,N_17947,N_17659);
and U18170 (N_18170,N_17721,N_17953);
nor U18171 (N_18171,N_17850,N_17548);
xnor U18172 (N_18172,N_17710,N_17772);
xnor U18173 (N_18173,N_17798,N_17683);
xor U18174 (N_18174,N_17689,N_17727);
xor U18175 (N_18175,N_17939,N_17610);
and U18176 (N_18176,N_17658,N_17633);
xor U18177 (N_18177,N_17925,N_17770);
xnor U18178 (N_18178,N_17743,N_17871);
nand U18179 (N_18179,N_17973,N_17643);
nand U18180 (N_18180,N_17921,N_17539);
nor U18181 (N_18181,N_17577,N_17741);
nor U18182 (N_18182,N_17669,N_17896);
nor U18183 (N_18183,N_17932,N_17928);
and U18184 (N_18184,N_17962,N_17876);
xor U18185 (N_18185,N_17978,N_17516);
and U18186 (N_18186,N_17640,N_17745);
nand U18187 (N_18187,N_17703,N_17996);
or U18188 (N_18188,N_17587,N_17708);
xnor U18189 (N_18189,N_17837,N_17728);
nor U18190 (N_18190,N_17532,N_17579);
nand U18191 (N_18191,N_17796,N_17716);
or U18192 (N_18192,N_17755,N_17594);
nor U18193 (N_18193,N_17908,N_17823);
xnor U18194 (N_18194,N_17808,N_17538);
and U18195 (N_18195,N_17725,N_17935);
and U18196 (N_18196,N_17645,N_17709);
or U18197 (N_18197,N_17991,N_17597);
nor U18198 (N_18198,N_17674,N_17874);
xor U18199 (N_18199,N_17979,N_17732);
nor U18200 (N_18200,N_17693,N_17985);
or U18201 (N_18201,N_17999,N_17774);
nand U18202 (N_18202,N_17846,N_17794);
xnor U18203 (N_18203,N_17653,N_17644);
nand U18204 (N_18204,N_17761,N_17938);
xor U18205 (N_18205,N_17944,N_17585);
xor U18206 (N_18206,N_17884,N_17945);
nand U18207 (N_18207,N_17968,N_17583);
and U18208 (N_18208,N_17773,N_17888);
nand U18209 (N_18209,N_17560,N_17615);
nor U18210 (N_18210,N_17634,N_17909);
nor U18211 (N_18211,N_17618,N_17691);
nand U18212 (N_18212,N_17715,N_17694);
nor U18213 (N_18213,N_17599,N_17933);
nand U18214 (N_18214,N_17782,N_17859);
and U18215 (N_18215,N_17806,N_17649);
and U18216 (N_18216,N_17994,N_17612);
xnor U18217 (N_18217,N_17701,N_17835);
and U18218 (N_18218,N_17914,N_17697);
or U18219 (N_18219,N_17534,N_17528);
and U18220 (N_18220,N_17541,N_17503);
nand U18221 (N_18221,N_17555,N_17960);
nor U18222 (N_18222,N_17992,N_17738);
nand U18223 (N_18223,N_17834,N_17657);
xnor U18224 (N_18224,N_17647,N_17873);
or U18225 (N_18225,N_17902,N_17505);
and U18226 (N_18226,N_17602,N_17684);
and U18227 (N_18227,N_17591,N_17668);
and U18228 (N_18228,N_17730,N_17842);
nand U18229 (N_18229,N_17639,N_17980);
nor U18230 (N_18230,N_17519,N_17678);
nor U18231 (N_18231,N_17749,N_17664);
and U18232 (N_18232,N_17853,N_17923);
xnor U18233 (N_18233,N_17997,N_17887);
or U18234 (N_18234,N_17545,N_17751);
xnor U18235 (N_18235,N_17757,N_17788);
nor U18236 (N_18236,N_17890,N_17900);
xor U18237 (N_18237,N_17786,N_17753);
xor U18238 (N_18238,N_17695,N_17899);
nor U18239 (N_18239,N_17765,N_17717);
or U18240 (N_18240,N_17672,N_17542);
nor U18241 (N_18241,N_17912,N_17637);
xnor U18242 (N_18242,N_17670,N_17763);
nand U18243 (N_18243,N_17556,N_17581);
and U18244 (N_18244,N_17574,N_17993);
or U18245 (N_18245,N_17840,N_17885);
or U18246 (N_18246,N_17518,N_17595);
xor U18247 (N_18247,N_17650,N_17667);
and U18248 (N_18248,N_17609,N_17685);
xnor U18249 (N_18249,N_17974,N_17740);
and U18250 (N_18250,N_17559,N_17540);
nand U18251 (N_18251,N_17721,N_17631);
xor U18252 (N_18252,N_17967,N_17555);
and U18253 (N_18253,N_17523,N_17713);
nor U18254 (N_18254,N_17683,N_17710);
and U18255 (N_18255,N_17601,N_17917);
xor U18256 (N_18256,N_17541,N_17673);
and U18257 (N_18257,N_17880,N_17665);
or U18258 (N_18258,N_17884,N_17611);
nor U18259 (N_18259,N_17864,N_17857);
nor U18260 (N_18260,N_17530,N_17811);
or U18261 (N_18261,N_17997,N_17714);
xnor U18262 (N_18262,N_17925,N_17559);
nand U18263 (N_18263,N_17750,N_17654);
and U18264 (N_18264,N_17718,N_17654);
nor U18265 (N_18265,N_17618,N_17826);
nor U18266 (N_18266,N_17786,N_17525);
xnor U18267 (N_18267,N_17958,N_17971);
or U18268 (N_18268,N_17623,N_17562);
nand U18269 (N_18269,N_17623,N_17719);
and U18270 (N_18270,N_17814,N_17965);
or U18271 (N_18271,N_17676,N_17774);
and U18272 (N_18272,N_17565,N_17999);
xnor U18273 (N_18273,N_17769,N_17794);
nor U18274 (N_18274,N_17981,N_17692);
and U18275 (N_18275,N_17627,N_17949);
nand U18276 (N_18276,N_17889,N_17901);
xor U18277 (N_18277,N_17563,N_17612);
and U18278 (N_18278,N_17793,N_17987);
nor U18279 (N_18279,N_17921,N_17677);
and U18280 (N_18280,N_17625,N_17919);
xor U18281 (N_18281,N_17505,N_17909);
nor U18282 (N_18282,N_17987,N_17671);
nor U18283 (N_18283,N_17778,N_17659);
and U18284 (N_18284,N_17957,N_17627);
nand U18285 (N_18285,N_17750,N_17780);
nand U18286 (N_18286,N_17577,N_17604);
nand U18287 (N_18287,N_17790,N_17723);
and U18288 (N_18288,N_17973,N_17536);
xnor U18289 (N_18289,N_17515,N_17725);
nand U18290 (N_18290,N_17631,N_17515);
and U18291 (N_18291,N_17932,N_17766);
nand U18292 (N_18292,N_17511,N_17553);
and U18293 (N_18293,N_17550,N_17836);
xnor U18294 (N_18294,N_17877,N_17730);
or U18295 (N_18295,N_17945,N_17798);
nor U18296 (N_18296,N_17543,N_17701);
and U18297 (N_18297,N_17753,N_17819);
xor U18298 (N_18298,N_17589,N_17540);
and U18299 (N_18299,N_17839,N_17892);
nor U18300 (N_18300,N_17648,N_17791);
nand U18301 (N_18301,N_17839,N_17769);
xor U18302 (N_18302,N_17657,N_17909);
nor U18303 (N_18303,N_17871,N_17521);
and U18304 (N_18304,N_17883,N_17779);
nand U18305 (N_18305,N_17938,N_17500);
xnor U18306 (N_18306,N_17532,N_17726);
xnor U18307 (N_18307,N_17663,N_17982);
xnor U18308 (N_18308,N_17724,N_17738);
nor U18309 (N_18309,N_17671,N_17642);
nand U18310 (N_18310,N_17648,N_17513);
and U18311 (N_18311,N_17536,N_17905);
or U18312 (N_18312,N_17887,N_17500);
nor U18313 (N_18313,N_17836,N_17718);
nor U18314 (N_18314,N_17825,N_17721);
xnor U18315 (N_18315,N_17668,N_17797);
and U18316 (N_18316,N_17578,N_17660);
nor U18317 (N_18317,N_17579,N_17703);
xnor U18318 (N_18318,N_17622,N_17605);
xnor U18319 (N_18319,N_17524,N_17814);
or U18320 (N_18320,N_17861,N_17660);
xor U18321 (N_18321,N_17855,N_17800);
and U18322 (N_18322,N_17803,N_17566);
or U18323 (N_18323,N_17966,N_17636);
or U18324 (N_18324,N_17968,N_17653);
and U18325 (N_18325,N_17770,N_17786);
and U18326 (N_18326,N_17684,N_17504);
nor U18327 (N_18327,N_17557,N_17609);
or U18328 (N_18328,N_17860,N_17788);
or U18329 (N_18329,N_17893,N_17930);
nor U18330 (N_18330,N_17790,N_17629);
and U18331 (N_18331,N_17710,N_17724);
xor U18332 (N_18332,N_17634,N_17685);
nor U18333 (N_18333,N_17650,N_17974);
nand U18334 (N_18334,N_17839,N_17845);
or U18335 (N_18335,N_17732,N_17808);
xnor U18336 (N_18336,N_17688,N_17933);
nand U18337 (N_18337,N_17574,N_17800);
nand U18338 (N_18338,N_17836,N_17874);
nor U18339 (N_18339,N_17756,N_17552);
xnor U18340 (N_18340,N_17756,N_17795);
nand U18341 (N_18341,N_17872,N_17779);
nor U18342 (N_18342,N_17607,N_17722);
and U18343 (N_18343,N_17962,N_17991);
nor U18344 (N_18344,N_17631,N_17733);
and U18345 (N_18345,N_17818,N_17825);
and U18346 (N_18346,N_17543,N_17588);
xnor U18347 (N_18347,N_17526,N_17959);
nand U18348 (N_18348,N_17579,N_17666);
nor U18349 (N_18349,N_17946,N_17984);
or U18350 (N_18350,N_17813,N_17674);
nor U18351 (N_18351,N_17504,N_17865);
xor U18352 (N_18352,N_17536,N_17546);
and U18353 (N_18353,N_17968,N_17508);
xnor U18354 (N_18354,N_17957,N_17679);
nand U18355 (N_18355,N_17886,N_17644);
xor U18356 (N_18356,N_17968,N_17951);
and U18357 (N_18357,N_17505,N_17632);
or U18358 (N_18358,N_17992,N_17867);
and U18359 (N_18359,N_17953,N_17638);
nor U18360 (N_18360,N_17599,N_17972);
nor U18361 (N_18361,N_17615,N_17736);
or U18362 (N_18362,N_17736,N_17916);
nand U18363 (N_18363,N_17816,N_17556);
xnor U18364 (N_18364,N_17978,N_17835);
xor U18365 (N_18365,N_17673,N_17536);
xnor U18366 (N_18366,N_17503,N_17880);
nor U18367 (N_18367,N_17578,N_17919);
nor U18368 (N_18368,N_17816,N_17733);
or U18369 (N_18369,N_17844,N_17624);
and U18370 (N_18370,N_17503,N_17530);
nor U18371 (N_18371,N_17747,N_17779);
nand U18372 (N_18372,N_17720,N_17692);
nand U18373 (N_18373,N_17552,N_17523);
and U18374 (N_18374,N_17736,N_17626);
and U18375 (N_18375,N_17789,N_17956);
nor U18376 (N_18376,N_17664,N_17757);
nor U18377 (N_18377,N_17896,N_17928);
or U18378 (N_18378,N_17800,N_17608);
or U18379 (N_18379,N_17572,N_17744);
and U18380 (N_18380,N_17850,N_17871);
and U18381 (N_18381,N_17663,N_17848);
nor U18382 (N_18382,N_17698,N_17810);
or U18383 (N_18383,N_17823,N_17561);
nand U18384 (N_18384,N_17543,N_17717);
or U18385 (N_18385,N_17612,N_17535);
nor U18386 (N_18386,N_17559,N_17973);
and U18387 (N_18387,N_17515,N_17966);
and U18388 (N_18388,N_17713,N_17618);
xnor U18389 (N_18389,N_17837,N_17681);
or U18390 (N_18390,N_17978,N_17786);
nand U18391 (N_18391,N_17853,N_17535);
xnor U18392 (N_18392,N_17583,N_17922);
or U18393 (N_18393,N_17607,N_17685);
and U18394 (N_18394,N_17893,N_17655);
or U18395 (N_18395,N_17830,N_17742);
nor U18396 (N_18396,N_17974,N_17627);
nand U18397 (N_18397,N_17579,N_17874);
and U18398 (N_18398,N_17517,N_17866);
or U18399 (N_18399,N_17925,N_17887);
nor U18400 (N_18400,N_17887,N_17941);
nor U18401 (N_18401,N_17946,N_17556);
nor U18402 (N_18402,N_17943,N_17821);
and U18403 (N_18403,N_17988,N_17711);
and U18404 (N_18404,N_17536,N_17950);
nand U18405 (N_18405,N_17813,N_17581);
or U18406 (N_18406,N_17574,N_17665);
and U18407 (N_18407,N_17834,N_17763);
or U18408 (N_18408,N_17856,N_17950);
and U18409 (N_18409,N_17798,N_17561);
xor U18410 (N_18410,N_17512,N_17972);
nand U18411 (N_18411,N_17711,N_17789);
nand U18412 (N_18412,N_17540,N_17705);
xnor U18413 (N_18413,N_17924,N_17580);
and U18414 (N_18414,N_17921,N_17729);
nor U18415 (N_18415,N_17886,N_17827);
or U18416 (N_18416,N_17819,N_17766);
xnor U18417 (N_18417,N_17699,N_17730);
xnor U18418 (N_18418,N_17774,N_17685);
or U18419 (N_18419,N_17575,N_17671);
nor U18420 (N_18420,N_17803,N_17589);
or U18421 (N_18421,N_17675,N_17871);
nand U18422 (N_18422,N_17586,N_17766);
and U18423 (N_18423,N_17676,N_17783);
or U18424 (N_18424,N_17979,N_17619);
xor U18425 (N_18425,N_17781,N_17750);
and U18426 (N_18426,N_17736,N_17742);
and U18427 (N_18427,N_17716,N_17920);
or U18428 (N_18428,N_17812,N_17761);
and U18429 (N_18429,N_17868,N_17878);
xor U18430 (N_18430,N_17887,N_17630);
nor U18431 (N_18431,N_17528,N_17652);
nor U18432 (N_18432,N_17874,N_17840);
nand U18433 (N_18433,N_17961,N_17769);
and U18434 (N_18434,N_17725,N_17841);
or U18435 (N_18435,N_17891,N_17808);
or U18436 (N_18436,N_17846,N_17710);
xor U18437 (N_18437,N_17945,N_17558);
and U18438 (N_18438,N_17500,N_17861);
nor U18439 (N_18439,N_17794,N_17535);
nor U18440 (N_18440,N_17733,N_17616);
nor U18441 (N_18441,N_17642,N_17518);
nor U18442 (N_18442,N_17511,N_17650);
and U18443 (N_18443,N_17698,N_17666);
or U18444 (N_18444,N_17784,N_17849);
or U18445 (N_18445,N_17846,N_17923);
and U18446 (N_18446,N_17999,N_17892);
nor U18447 (N_18447,N_17621,N_17539);
nand U18448 (N_18448,N_17732,N_17830);
nand U18449 (N_18449,N_17793,N_17950);
nor U18450 (N_18450,N_17580,N_17710);
xor U18451 (N_18451,N_17838,N_17629);
nor U18452 (N_18452,N_17668,N_17908);
nor U18453 (N_18453,N_17882,N_17526);
nor U18454 (N_18454,N_17551,N_17566);
nor U18455 (N_18455,N_17646,N_17895);
nor U18456 (N_18456,N_17982,N_17956);
and U18457 (N_18457,N_17602,N_17972);
and U18458 (N_18458,N_17860,N_17680);
nand U18459 (N_18459,N_17786,N_17569);
nand U18460 (N_18460,N_17983,N_17903);
nand U18461 (N_18461,N_17633,N_17666);
xor U18462 (N_18462,N_17918,N_17838);
and U18463 (N_18463,N_17602,N_17513);
nor U18464 (N_18464,N_17938,N_17537);
and U18465 (N_18465,N_17871,N_17510);
and U18466 (N_18466,N_17658,N_17514);
nor U18467 (N_18467,N_17746,N_17681);
nand U18468 (N_18468,N_17764,N_17882);
xor U18469 (N_18469,N_17994,N_17985);
or U18470 (N_18470,N_17796,N_17795);
and U18471 (N_18471,N_17789,N_17730);
nor U18472 (N_18472,N_17749,N_17904);
or U18473 (N_18473,N_17873,N_17852);
nor U18474 (N_18474,N_17986,N_17803);
xnor U18475 (N_18475,N_17758,N_17928);
or U18476 (N_18476,N_17542,N_17832);
nand U18477 (N_18477,N_17943,N_17759);
or U18478 (N_18478,N_17801,N_17655);
nor U18479 (N_18479,N_17816,N_17893);
nand U18480 (N_18480,N_17937,N_17925);
nand U18481 (N_18481,N_17516,N_17598);
nor U18482 (N_18482,N_17993,N_17962);
and U18483 (N_18483,N_17706,N_17735);
xor U18484 (N_18484,N_17736,N_17720);
and U18485 (N_18485,N_17551,N_17812);
nor U18486 (N_18486,N_17800,N_17665);
and U18487 (N_18487,N_17846,N_17577);
nor U18488 (N_18488,N_17889,N_17642);
xnor U18489 (N_18489,N_17660,N_17692);
or U18490 (N_18490,N_17716,N_17668);
xor U18491 (N_18491,N_17545,N_17930);
nand U18492 (N_18492,N_17537,N_17928);
nand U18493 (N_18493,N_17823,N_17841);
nor U18494 (N_18494,N_17640,N_17998);
xnor U18495 (N_18495,N_17970,N_17607);
and U18496 (N_18496,N_17611,N_17551);
nand U18497 (N_18497,N_17652,N_17868);
and U18498 (N_18498,N_17538,N_17902);
nand U18499 (N_18499,N_17587,N_17999);
or U18500 (N_18500,N_18232,N_18120);
nor U18501 (N_18501,N_18019,N_18434);
nor U18502 (N_18502,N_18145,N_18275);
nor U18503 (N_18503,N_18318,N_18157);
and U18504 (N_18504,N_18316,N_18491);
nand U18505 (N_18505,N_18359,N_18304);
or U18506 (N_18506,N_18297,N_18403);
nor U18507 (N_18507,N_18184,N_18239);
xor U18508 (N_18508,N_18109,N_18039);
or U18509 (N_18509,N_18313,N_18223);
nand U18510 (N_18510,N_18284,N_18391);
xnor U18511 (N_18511,N_18212,N_18324);
and U18512 (N_18512,N_18083,N_18222);
xor U18513 (N_18513,N_18490,N_18398);
nand U18514 (N_18514,N_18066,N_18264);
nor U18515 (N_18515,N_18429,N_18333);
nor U18516 (N_18516,N_18044,N_18058);
or U18517 (N_18517,N_18390,N_18048);
nor U18518 (N_18518,N_18042,N_18213);
xor U18519 (N_18519,N_18111,N_18245);
xnor U18520 (N_18520,N_18260,N_18117);
and U18521 (N_18521,N_18495,N_18203);
nor U18522 (N_18522,N_18069,N_18104);
nor U18523 (N_18523,N_18010,N_18293);
and U18524 (N_18524,N_18431,N_18241);
nor U18525 (N_18525,N_18253,N_18279);
nor U18526 (N_18526,N_18497,N_18342);
nand U18527 (N_18527,N_18400,N_18000);
and U18528 (N_18528,N_18057,N_18452);
and U18529 (N_18529,N_18226,N_18075);
and U18530 (N_18530,N_18414,N_18063);
and U18531 (N_18531,N_18041,N_18012);
nor U18532 (N_18532,N_18233,N_18467);
nand U18533 (N_18533,N_18485,N_18221);
xnor U18534 (N_18534,N_18468,N_18220);
nand U18535 (N_18535,N_18072,N_18187);
nor U18536 (N_18536,N_18127,N_18248);
xor U18537 (N_18537,N_18102,N_18440);
nor U18538 (N_18538,N_18464,N_18166);
or U18539 (N_18539,N_18352,N_18374);
and U18540 (N_18540,N_18257,N_18116);
xor U18541 (N_18541,N_18475,N_18094);
nand U18542 (N_18542,N_18405,N_18422);
or U18543 (N_18543,N_18446,N_18056);
nand U18544 (N_18544,N_18165,N_18499);
nor U18545 (N_18545,N_18181,N_18219);
or U18546 (N_18546,N_18443,N_18473);
nand U18547 (N_18547,N_18394,N_18118);
nand U18548 (N_18548,N_18060,N_18035);
nand U18549 (N_18549,N_18050,N_18470);
or U18550 (N_18550,N_18110,N_18476);
nor U18551 (N_18551,N_18381,N_18065);
nand U18552 (N_18552,N_18216,N_18123);
xnor U18553 (N_18553,N_18457,N_18015);
or U18554 (N_18554,N_18283,N_18299);
xnor U18555 (N_18555,N_18023,N_18438);
and U18556 (N_18556,N_18054,N_18489);
or U18557 (N_18557,N_18462,N_18498);
and U18558 (N_18558,N_18418,N_18492);
and U18559 (N_18559,N_18406,N_18349);
nand U18560 (N_18560,N_18073,N_18142);
and U18561 (N_18561,N_18481,N_18001);
nor U18562 (N_18562,N_18286,N_18325);
and U18563 (N_18563,N_18100,N_18017);
nor U18564 (N_18564,N_18340,N_18049);
or U18565 (N_18565,N_18295,N_18122);
or U18566 (N_18566,N_18236,N_18266);
nand U18567 (N_18567,N_18327,N_18173);
and U18568 (N_18568,N_18303,N_18330);
nand U18569 (N_18569,N_18089,N_18254);
and U18570 (N_18570,N_18484,N_18027);
xnor U18571 (N_18571,N_18176,N_18441);
xnor U18572 (N_18572,N_18396,N_18105);
or U18573 (N_18573,N_18045,N_18119);
and U18574 (N_18574,N_18332,N_18336);
or U18575 (N_18575,N_18425,N_18315);
or U18576 (N_18576,N_18093,N_18435);
xor U18577 (N_18577,N_18183,N_18206);
or U18578 (N_18578,N_18387,N_18351);
xor U18579 (N_18579,N_18229,N_18258);
nand U18580 (N_18580,N_18404,N_18353);
and U18581 (N_18581,N_18141,N_18193);
nand U18582 (N_18582,N_18417,N_18259);
nand U18583 (N_18583,N_18186,N_18059);
nand U18584 (N_18584,N_18310,N_18494);
or U18585 (N_18585,N_18482,N_18433);
and U18586 (N_18586,N_18392,N_18150);
or U18587 (N_18587,N_18209,N_18004);
nor U18588 (N_18588,N_18134,N_18458);
xor U18589 (N_18589,N_18114,N_18115);
or U18590 (N_18590,N_18191,N_18098);
or U18591 (N_18591,N_18024,N_18029);
and U18592 (N_18592,N_18430,N_18235);
or U18593 (N_18593,N_18357,N_18133);
and U18594 (N_18594,N_18338,N_18179);
nand U18595 (N_18595,N_18466,N_18095);
nor U18596 (N_18596,N_18393,N_18486);
nand U18597 (N_18597,N_18265,N_18322);
nor U18598 (N_18598,N_18210,N_18269);
or U18599 (N_18599,N_18368,N_18106);
and U18600 (N_18600,N_18188,N_18159);
nand U18601 (N_18601,N_18345,N_18250);
and U18602 (N_18602,N_18428,N_18472);
nor U18603 (N_18603,N_18280,N_18361);
or U18604 (N_18604,N_18377,N_18407);
xnor U18605 (N_18605,N_18113,N_18389);
nand U18606 (N_18606,N_18447,N_18140);
xnor U18607 (N_18607,N_18294,N_18161);
nor U18608 (N_18608,N_18018,N_18085);
nor U18609 (N_18609,N_18300,N_18331);
xor U18610 (N_18610,N_18046,N_18070);
nor U18611 (N_18611,N_18323,N_18192);
or U18612 (N_18612,N_18397,N_18380);
or U18613 (N_18613,N_18419,N_18252);
nand U18614 (N_18614,N_18395,N_18432);
or U18615 (N_18615,N_18281,N_18454);
nand U18616 (N_18616,N_18308,N_18087);
nand U18617 (N_18617,N_18026,N_18347);
and U18618 (N_18618,N_18456,N_18080);
nand U18619 (N_18619,N_18341,N_18008);
nor U18620 (N_18620,N_18350,N_18167);
and U18621 (N_18621,N_18388,N_18137);
or U18622 (N_18622,N_18383,N_18180);
xnor U18623 (N_18623,N_18171,N_18092);
xnor U18624 (N_18624,N_18261,N_18288);
nand U18625 (N_18625,N_18439,N_18162);
nand U18626 (N_18626,N_18262,N_18363);
and U18627 (N_18627,N_18444,N_18423);
and U18628 (N_18628,N_18339,N_18047);
nand U18629 (N_18629,N_18243,N_18034);
nand U18630 (N_18630,N_18376,N_18409);
or U18631 (N_18631,N_18256,N_18451);
or U18632 (N_18632,N_18379,N_18202);
nor U18633 (N_18633,N_18449,N_18052);
or U18634 (N_18634,N_18346,N_18146);
and U18635 (N_18635,N_18354,N_18138);
nor U18636 (N_18636,N_18021,N_18125);
and U18637 (N_18637,N_18020,N_18465);
nor U18638 (N_18638,N_18459,N_18007);
xor U18639 (N_18639,N_18172,N_18311);
nand U18640 (N_18640,N_18287,N_18448);
nand U18641 (N_18641,N_18471,N_18025);
or U18642 (N_18642,N_18061,N_18282);
xor U18643 (N_18643,N_18121,N_18016);
nand U18644 (N_18644,N_18301,N_18153);
and U18645 (N_18645,N_18415,N_18372);
nand U18646 (N_18646,N_18413,N_18163);
nor U18647 (N_18647,N_18450,N_18129);
nor U18648 (N_18648,N_18197,N_18320);
xnor U18649 (N_18649,N_18211,N_18107);
and U18650 (N_18650,N_18190,N_18289);
nor U18651 (N_18651,N_18445,N_18096);
or U18652 (N_18652,N_18182,N_18329);
and U18653 (N_18653,N_18401,N_18097);
or U18654 (N_18654,N_18296,N_18399);
and U18655 (N_18655,N_18081,N_18128);
or U18656 (N_18656,N_18384,N_18437);
or U18657 (N_18657,N_18364,N_18463);
nor U18658 (N_18658,N_18496,N_18189);
xor U18659 (N_18659,N_18369,N_18426);
nand U18660 (N_18660,N_18231,N_18147);
nand U18661 (N_18661,N_18022,N_18263);
nor U18662 (N_18662,N_18319,N_18195);
and U18663 (N_18663,N_18074,N_18077);
nand U18664 (N_18664,N_18267,N_18099);
and U18665 (N_18665,N_18148,N_18108);
xor U18666 (N_18666,N_18086,N_18273);
or U18667 (N_18667,N_18224,N_18132);
xor U18668 (N_18668,N_18488,N_18237);
or U18669 (N_18669,N_18040,N_18208);
nor U18670 (N_18670,N_18360,N_18242);
nor U18671 (N_18671,N_18305,N_18067);
nor U18672 (N_18672,N_18402,N_18274);
nand U18673 (N_18673,N_18358,N_18234);
or U18674 (N_18674,N_18006,N_18317);
or U18675 (N_18675,N_18088,N_18478);
or U18676 (N_18676,N_18199,N_18314);
xor U18677 (N_18677,N_18386,N_18101);
nand U18678 (N_18678,N_18480,N_18469);
and U18679 (N_18679,N_18355,N_18170);
and U18680 (N_18680,N_18064,N_18068);
xnor U18681 (N_18681,N_18130,N_18453);
nand U18682 (N_18682,N_18156,N_18373);
nor U18683 (N_18683,N_18328,N_18420);
xnor U18684 (N_18684,N_18278,N_18144);
and U18685 (N_18685,N_18312,N_18168);
nor U18686 (N_18686,N_18427,N_18079);
or U18687 (N_18687,N_18178,N_18136);
or U18688 (N_18688,N_18043,N_18442);
nand U18689 (N_18689,N_18196,N_18071);
and U18690 (N_18690,N_18412,N_18230);
or U18691 (N_18691,N_18215,N_18032);
nor U18692 (N_18692,N_18014,N_18185);
xor U18693 (N_18693,N_18411,N_18307);
nor U18694 (N_18694,N_18177,N_18053);
xor U18695 (N_18695,N_18149,N_18285);
or U18696 (N_18696,N_18135,N_18362);
nor U18697 (N_18697,N_18055,N_18277);
xnor U18698 (N_18698,N_18348,N_18477);
xnor U18699 (N_18699,N_18218,N_18493);
nor U18700 (N_18700,N_18062,N_18337);
xnor U18701 (N_18701,N_18408,N_18483);
nor U18702 (N_18702,N_18272,N_18217);
nand U18703 (N_18703,N_18334,N_18090);
and U18704 (N_18704,N_18251,N_18051);
nor U18705 (N_18705,N_18028,N_18487);
or U18706 (N_18706,N_18091,N_18343);
or U18707 (N_18707,N_18201,N_18126);
and U18708 (N_18708,N_18082,N_18225);
nor U18709 (N_18709,N_18276,N_18474);
or U18710 (N_18710,N_18036,N_18292);
or U18711 (N_18711,N_18246,N_18461);
xnor U18712 (N_18712,N_18247,N_18255);
or U18713 (N_18713,N_18367,N_18321);
nor U18714 (N_18714,N_18356,N_18291);
and U18715 (N_18715,N_18227,N_18479);
nor U18716 (N_18716,N_18240,N_18326);
nand U18717 (N_18717,N_18037,N_18244);
and U18718 (N_18718,N_18460,N_18455);
xor U18719 (N_18719,N_18139,N_18424);
nor U18720 (N_18720,N_18436,N_18154);
nor U18721 (N_18721,N_18410,N_18152);
nand U18722 (N_18722,N_18155,N_18131);
and U18723 (N_18723,N_18084,N_18005);
xnor U18724 (N_18724,N_18112,N_18366);
or U18725 (N_18725,N_18009,N_18385);
or U18726 (N_18726,N_18271,N_18421);
xor U18727 (N_18727,N_18268,N_18011);
xnor U18728 (N_18728,N_18003,N_18198);
nor U18729 (N_18729,N_18002,N_18270);
nor U18730 (N_18730,N_18103,N_18344);
or U18731 (N_18731,N_18238,N_18174);
nor U18732 (N_18732,N_18031,N_18078);
and U18733 (N_18733,N_18335,N_18194);
or U18734 (N_18734,N_18169,N_18076);
or U18735 (N_18735,N_18298,N_18030);
and U18736 (N_18736,N_18124,N_18160);
or U18737 (N_18737,N_18214,N_18205);
nor U18738 (N_18738,N_18378,N_18143);
nand U18739 (N_18739,N_18204,N_18371);
nand U18740 (N_18740,N_18302,N_18151);
xor U18741 (N_18741,N_18416,N_18365);
nand U18742 (N_18742,N_18375,N_18207);
xnor U18743 (N_18743,N_18038,N_18200);
xor U18744 (N_18744,N_18033,N_18175);
or U18745 (N_18745,N_18249,N_18228);
nand U18746 (N_18746,N_18290,N_18013);
or U18747 (N_18747,N_18306,N_18158);
and U18748 (N_18748,N_18164,N_18309);
and U18749 (N_18749,N_18370,N_18382);
nand U18750 (N_18750,N_18482,N_18457);
xnor U18751 (N_18751,N_18097,N_18194);
or U18752 (N_18752,N_18153,N_18006);
nand U18753 (N_18753,N_18141,N_18462);
xor U18754 (N_18754,N_18393,N_18320);
nand U18755 (N_18755,N_18219,N_18269);
and U18756 (N_18756,N_18157,N_18434);
nor U18757 (N_18757,N_18332,N_18303);
xnor U18758 (N_18758,N_18013,N_18097);
and U18759 (N_18759,N_18084,N_18407);
xnor U18760 (N_18760,N_18203,N_18103);
or U18761 (N_18761,N_18013,N_18028);
nor U18762 (N_18762,N_18025,N_18146);
and U18763 (N_18763,N_18138,N_18399);
nand U18764 (N_18764,N_18200,N_18371);
nor U18765 (N_18765,N_18487,N_18168);
xnor U18766 (N_18766,N_18420,N_18353);
or U18767 (N_18767,N_18302,N_18125);
xor U18768 (N_18768,N_18254,N_18106);
nor U18769 (N_18769,N_18249,N_18185);
and U18770 (N_18770,N_18296,N_18087);
nand U18771 (N_18771,N_18220,N_18216);
nand U18772 (N_18772,N_18352,N_18459);
xnor U18773 (N_18773,N_18391,N_18396);
nand U18774 (N_18774,N_18395,N_18236);
xnor U18775 (N_18775,N_18263,N_18395);
nor U18776 (N_18776,N_18133,N_18137);
xnor U18777 (N_18777,N_18032,N_18430);
xor U18778 (N_18778,N_18478,N_18056);
and U18779 (N_18779,N_18284,N_18004);
or U18780 (N_18780,N_18415,N_18442);
and U18781 (N_18781,N_18116,N_18475);
nand U18782 (N_18782,N_18255,N_18316);
nand U18783 (N_18783,N_18266,N_18035);
or U18784 (N_18784,N_18423,N_18414);
and U18785 (N_18785,N_18195,N_18209);
xnor U18786 (N_18786,N_18116,N_18309);
and U18787 (N_18787,N_18052,N_18357);
xnor U18788 (N_18788,N_18056,N_18393);
nand U18789 (N_18789,N_18330,N_18307);
nand U18790 (N_18790,N_18167,N_18393);
and U18791 (N_18791,N_18174,N_18347);
nand U18792 (N_18792,N_18070,N_18090);
xnor U18793 (N_18793,N_18134,N_18484);
nor U18794 (N_18794,N_18464,N_18284);
nor U18795 (N_18795,N_18456,N_18326);
and U18796 (N_18796,N_18387,N_18384);
xnor U18797 (N_18797,N_18467,N_18041);
xor U18798 (N_18798,N_18401,N_18144);
or U18799 (N_18799,N_18485,N_18142);
nor U18800 (N_18800,N_18386,N_18496);
xor U18801 (N_18801,N_18426,N_18296);
nand U18802 (N_18802,N_18048,N_18482);
nand U18803 (N_18803,N_18360,N_18295);
nand U18804 (N_18804,N_18292,N_18331);
nand U18805 (N_18805,N_18036,N_18203);
xnor U18806 (N_18806,N_18078,N_18193);
and U18807 (N_18807,N_18159,N_18136);
or U18808 (N_18808,N_18170,N_18362);
nor U18809 (N_18809,N_18166,N_18294);
xor U18810 (N_18810,N_18385,N_18323);
or U18811 (N_18811,N_18010,N_18120);
and U18812 (N_18812,N_18327,N_18159);
xor U18813 (N_18813,N_18131,N_18228);
nor U18814 (N_18814,N_18375,N_18223);
nand U18815 (N_18815,N_18036,N_18200);
or U18816 (N_18816,N_18488,N_18312);
or U18817 (N_18817,N_18147,N_18449);
nand U18818 (N_18818,N_18430,N_18292);
and U18819 (N_18819,N_18133,N_18482);
or U18820 (N_18820,N_18263,N_18155);
and U18821 (N_18821,N_18330,N_18039);
or U18822 (N_18822,N_18460,N_18205);
and U18823 (N_18823,N_18086,N_18296);
nand U18824 (N_18824,N_18099,N_18462);
nand U18825 (N_18825,N_18002,N_18005);
nand U18826 (N_18826,N_18120,N_18221);
and U18827 (N_18827,N_18382,N_18246);
nor U18828 (N_18828,N_18446,N_18217);
xor U18829 (N_18829,N_18341,N_18198);
nand U18830 (N_18830,N_18084,N_18116);
xnor U18831 (N_18831,N_18387,N_18458);
nand U18832 (N_18832,N_18082,N_18361);
or U18833 (N_18833,N_18243,N_18326);
nand U18834 (N_18834,N_18497,N_18401);
and U18835 (N_18835,N_18280,N_18296);
and U18836 (N_18836,N_18105,N_18045);
xnor U18837 (N_18837,N_18489,N_18208);
xnor U18838 (N_18838,N_18148,N_18008);
and U18839 (N_18839,N_18346,N_18337);
or U18840 (N_18840,N_18177,N_18130);
nand U18841 (N_18841,N_18050,N_18278);
nor U18842 (N_18842,N_18233,N_18425);
nor U18843 (N_18843,N_18235,N_18364);
or U18844 (N_18844,N_18070,N_18198);
nand U18845 (N_18845,N_18102,N_18055);
and U18846 (N_18846,N_18113,N_18393);
and U18847 (N_18847,N_18160,N_18139);
and U18848 (N_18848,N_18415,N_18429);
and U18849 (N_18849,N_18125,N_18214);
or U18850 (N_18850,N_18134,N_18325);
nor U18851 (N_18851,N_18478,N_18298);
or U18852 (N_18852,N_18121,N_18266);
nor U18853 (N_18853,N_18078,N_18490);
nor U18854 (N_18854,N_18496,N_18362);
nor U18855 (N_18855,N_18117,N_18371);
or U18856 (N_18856,N_18299,N_18034);
nor U18857 (N_18857,N_18117,N_18121);
and U18858 (N_18858,N_18306,N_18437);
or U18859 (N_18859,N_18205,N_18327);
nand U18860 (N_18860,N_18104,N_18464);
and U18861 (N_18861,N_18426,N_18363);
nor U18862 (N_18862,N_18486,N_18386);
or U18863 (N_18863,N_18236,N_18293);
xor U18864 (N_18864,N_18368,N_18154);
nand U18865 (N_18865,N_18351,N_18030);
nor U18866 (N_18866,N_18200,N_18203);
nor U18867 (N_18867,N_18062,N_18076);
nand U18868 (N_18868,N_18448,N_18418);
xor U18869 (N_18869,N_18232,N_18149);
xor U18870 (N_18870,N_18055,N_18145);
and U18871 (N_18871,N_18075,N_18327);
or U18872 (N_18872,N_18135,N_18463);
and U18873 (N_18873,N_18444,N_18200);
and U18874 (N_18874,N_18362,N_18173);
xnor U18875 (N_18875,N_18279,N_18449);
xor U18876 (N_18876,N_18033,N_18076);
or U18877 (N_18877,N_18214,N_18340);
nor U18878 (N_18878,N_18487,N_18058);
and U18879 (N_18879,N_18008,N_18108);
or U18880 (N_18880,N_18004,N_18463);
and U18881 (N_18881,N_18004,N_18033);
nor U18882 (N_18882,N_18154,N_18216);
or U18883 (N_18883,N_18054,N_18492);
xnor U18884 (N_18884,N_18384,N_18112);
nand U18885 (N_18885,N_18248,N_18167);
nand U18886 (N_18886,N_18190,N_18463);
nor U18887 (N_18887,N_18453,N_18366);
xor U18888 (N_18888,N_18451,N_18110);
xor U18889 (N_18889,N_18427,N_18399);
or U18890 (N_18890,N_18344,N_18473);
nand U18891 (N_18891,N_18157,N_18016);
nand U18892 (N_18892,N_18482,N_18422);
or U18893 (N_18893,N_18320,N_18306);
and U18894 (N_18894,N_18135,N_18167);
nand U18895 (N_18895,N_18092,N_18295);
xnor U18896 (N_18896,N_18170,N_18077);
or U18897 (N_18897,N_18420,N_18019);
nor U18898 (N_18898,N_18343,N_18062);
nand U18899 (N_18899,N_18174,N_18459);
or U18900 (N_18900,N_18014,N_18481);
or U18901 (N_18901,N_18234,N_18413);
and U18902 (N_18902,N_18403,N_18155);
xor U18903 (N_18903,N_18264,N_18499);
nand U18904 (N_18904,N_18321,N_18388);
nand U18905 (N_18905,N_18428,N_18114);
or U18906 (N_18906,N_18251,N_18102);
or U18907 (N_18907,N_18220,N_18359);
nand U18908 (N_18908,N_18426,N_18441);
nor U18909 (N_18909,N_18076,N_18041);
or U18910 (N_18910,N_18250,N_18113);
or U18911 (N_18911,N_18197,N_18333);
xor U18912 (N_18912,N_18157,N_18046);
or U18913 (N_18913,N_18127,N_18101);
nor U18914 (N_18914,N_18179,N_18113);
or U18915 (N_18915,N_18344,N_18354);
or U18916 (N_18916,N_18212,N_18087);
xnor U18917 (N_18917,N_18091,N_18419);
and U18918 (N_18918,N_18296,N_18416);
nand U18919 (N_18919,N_18283,N_18061);
nor U18920 (N_18920,N_18217,N_18292);
nor U18921 (N_18921,N_18403,N_18440);
and U18922 (N_18922,N_18231,N_18027);
nand U18923 (N_18923,N_18465,N_18165);
and U18924 (N_18924,N_18101,N_18034);
xnor U18925 (N_18925,N_18409,N_18102);
nand U18926 (N_18926,N_18494,N_18363);
nand U18927 (N_18927,N_18432,N_18497);
nor U18928 (N_18928,N_18439,N_18249);
and U18929 (N_18929,N_18359,N_18019);
or U18930 (N_18930,N_18091,N_18328);
nand U18931 (N_18931,N_18131,N_18287);
nand U18932 (N_18932,N_18104,N_18081);
and U18933 (N_18933,N_18249,N_18161);
and U18934 (N_18934,N_18367,N_18065);
xnor U18935 (N_18935,N_18399,N_18280);
or U18936 (N_18936,N_18315,N_18489);
xnor U18937 (N_18937,N_18416,N_18079);
xnor U18938 (N_18938,N_18146,N_18065);
nor U18939 (N_18939,N_18264,N_18350);
nor U18940 (N_18940,N_18009,N_18335);
nor U18941 (N_18941,N_18185,N_18372);
and U18942 (N_18942,N_18332,N_18144);
xor U18943 (N_18943,N_18139,N_18029);
or U18944 (N_18944,N_18018,N_18431);
xnor U18945 (N_18945,N_18267,N_18001);
and U18946 (N_18946,N_18094,N_18279);
and U18947 (N_18947,N_18288,N_18408);
nand U18948 (N_18948,N_18452,N_18408);
nand U18949 (N_18949,N_18477,N_18021);
xnor U18950 (N_18950,N_18087,N_18256);
or U18951 (N_18951,N_18333,N_18423);
or U18952 (N_18952,N_18105,N_18087);
or U18953 (N_18953,N_18455,N_18201);
nand U18954 (N_18954,N_18237,N_18149);
and U18955 (N_18955,N_18132,N_18101);
nor U18956 (N_18956,N_18351,N_18000);
nor U18957 (N_18957,N_18189,N_18273);
nor U18958 (N_18958,N_18245,N_18064);
xnor U18959 (N_18959,N_18229,N_18071);
or U18960 (N_18960,N_18255,N_18478);
or U18961 (N_18961,N_18176,N_18248);
or U18962 (N_18962,N_18151,N_18076);
xnor U18963 (N_18963,N_18019,N_18249);
nor U18964 (N_18964,N_18402,N_18455);
or U18965 (N_18965,N_18160,N_18405);
nor U18966 (N_18966,N_18362,N_18331);
nor U18967 (N_18967,N_18158,N_18474);
and U18968 (N_18968,N_18465,N_18137);
nor U18969 (N_18969,N_18473,N_18350);
nand U18970 (N_18970,N_18253,N_18211);
nand U18971 (N_18971,N_18436,N_18217);
nor U18972 (N_18972,N_18270,N_18020);
nand U18973 (N_18973,N_18321,N_18104);
and U18974 (N_18974,N_18110,N_18262);
nand U18975 (N_18975,N_18439,N_18049);
and U18976 (N_18976,N_18075,N_18138);
and U18977 (N_18977,N_18319,N_18240);
or U18978 (N_18978,N_18303,N_18167);
or U18979 (N_18979,N_18047,N_18234);
xnor U18980 (N_18980,N_18040,N_18065);
or U18981 (N_18981,N_18151,N_18342);
nand U18982 (N_18982,N_18032,N_18425);
or U18983 (N_18983,N_18360,N_18225);
nor U18984 (N_18984,N_18388,N_18440);
or U18985 (N_18985,N_18127,N_18384);
or U18986 (N_18986,N_18169,N_18131);
nor U18987 (N_18987,N_18049,N_18006);
xnor U18988 (N_18988,N_18430,N_18377);
or U18989 (N_18989,N_18146,N_18302);
and U18990 (N_18990,N_18202,N_18395);
nand U18991 (N_18991,N_18303,N_18346);
and U18992 (N_18992,N_18051,N_18443);
or U18993 (N_18993,N_18196,N_18150);
xor U18994 (N_18994,N_18405,N_18209);
xnor U18995 (N_18995,N_18141,N_18342);
nand U18996 (N_18996,N_18172,N_18399);
nor U18997 (N_18997,N_18381,N_18075);
and U18998 (N_18998,N_18228,N_18483);
or U18999 (N_18999,N_18381,N_18238);
or U19000 (N_19000,N_18801,N_18802);
xnor U19001 (N_19001,N_18988,N_18654);
nor U19002 (N_19002,N_18666,N_18655);
nor U19003 (N_19003,N_18745,N_18785);
nor U19004 (N_19004,N_18888,N_18850);
and U19005 (N_19005,N_18670,N_18677);
nand U19006 (N_19006,N_18772,N_18693);
xor U19007 (N_19007,N_18832,N_18513);
or U19008 (N_19008,N_18936,N_18896);
nor U19009 (N_19009,N_18508,N_18731);
xnor U19010 (N_19010,N_18770,N_18911);
and U19011 (N_19011,N_18766,N_18605);
nand U19012 (N_19012,N_18705,N_18556);
or U19013 (N_19013,N_18930,N_18619);
nor U19014 (N_19014,N_18584,N_18664);
nand U19015 (N_19015,N_18918,N_18885);
or U19016 (N_19016,N_18637,N_18678);
or U19017 (N_19017,N_18505,N_18531);
nor U19018 (N_19018,N_18915,N_18815);
and U19019 (N_19019,N_18750,N_18681);
nand U19020 (N_19020,N_18868,N_18611);
nor U19021 (N_19021,N_18922,N_18582);
xor U19022 (N_19022,N_18916,N_18628);
or U19023 (N_19023,N_18763,N_18983);
xnor U19024 (N_19024,N_18842,N_18963);
and U19025 (N_19025,N_18536,N_18835);
or U19026 (N_19026,N_18703,N_18831);
nor U19027 (N_19027,N_18645,N_18525);
xnor U19028 (N_19028,N_18503,N_18547);
and U19029 (N_19029,N_18720,N_18601);
nor U19030 (N_19030,N_18587,N_18551);
or U19031 (N_19031,N_18585,N_18941);
xor U19032 (N_19032,N_18501,N_18775);
and U19033 (N_19033,N_18532,N_18638);
and U19034 (N_19034,N_18697,N_18538);
nor U19035 (N_19035,N_18722,N_18844);
xor U19036 (N_19036,N_18612,N_18728);
nand U19037 (N_19037,N_18984,N_18694);
xor U19038 (N_19038,N_18883,N_18928);
nand U19039 (N_19039,N_18620,N_18700);
or U19040 (N_19040,N_18895,N_18735);
nor U19041 (N_19041,N_18564,N_18784);
or U19042 (N_19042,N_18648,N_18644);
nand U19043 (N_19043,N_18980,N_18874);
and U19044 (N_19044,N_18956,N_18518);
or U19045 (N_19045,N_18991,N_18771);
or U19046 (N_19046,N_18899,N_18836);
and U19047 (N_19047,N_18864,N_18751);
or U19048 (N_19048,N_18816,N_18588);
xnor U19049 (N_19049,N_18867,N_18908);
nor U19050 (N_19050,N_18753,N_18553);
xnor U19051 (N_19051,N_18987,N_18923);
xor U19052 (N_19052,N_18990,N_18861);
nand U19053 (N_19053,N_18876,N_18892);
nand U19054 (N_19054,N_18934,N_18590);
and U19055 (N_19055,N_18760,N_18557);
and U19056 (N_19056,N_18546,N_18796);
or U19057 (N_19057,N_18737,N_18758);
nor U19058 (N_19058,N_18545,N_18625);
and U19059 (N_19059,N_18691,N_18597);
xor U19060 (N_19060,N_18929,N_18591);
xor U19061 (N_19061,N_18889,N_18920);
xor U19062 (N_19062,N_18897,N_18976);
xor U19063 (N_19063,N_18552,N_18849);
and U19064 (N_19064,N_18739,N_18989);
nor U19065 (N_19065,N_18807,N_18740);
nand U19066 (N_19066,N_18572,N_18790);
nor U19067 (N_19067,N_18841,N_18847);
or U19068 (N_19068,N_18643,N_18568);
and U19069 (N_19069,N_18774,N_18602);
and U19070 (N_19070,N_18819,N_18960);
nor U19071 (N_19071,N_18979,N_18875);
xnor U19072 (N_19072,N_18839,N_18732);
and U19073 (N_19073,N_18578,N_18729);
or U19074 (N_19074,N_18569,N_18893);
xor U19075 (N_19075,N_18562,N_18509);
or U19076 (N_19076,N_18792,N_18665);
and U19077 (N_19077,N_18629,N_18523);
nor U19078 (N_19078,N_18773,N_18887);
or U19079 (N_19079,N_18945,N_18527);
nor U19080 (N_19080,N_18676,N_18671);
nand U19081 (N_19081,N_18596,N_18610);
and U19082 (N_19082,N_18719,N_18811);
nand U19083 (N_19083,N_18827,N_18768);
xnor U19084 (N_19084,N_18798,N_18617);
or U19085 (N_19085,N_18971,N_18521);
nor U19086 (N_19086,N_18820,N_18723);
and U19087 (N_19087,N_18944,N_18765);
nor U19088 (N_19088,N_18573,N_18684);
or U19089 (N_19089,N_18948,N_18707);
xnor U19090 (N_19090,N_18913,N_18738);
nand U19091 (N_19091,N_18709,N_18794);
nor U19092 (N_19092,N_18608,N_18873);
or U19093 (N_19093,N_18789,N_18871);
nand U19094 (N_19094,N_18726,N_18517);
nand U19095 (N_19095,N_18717,N_18519);
nand U19096 (N_19096,N_18649,N_18878);
nand U19097 (N_19097,N_18622,N_18529);
xor U19098 (N_19098,N_18992,N_18997);
xor U19099 (N_19099,N_18621,N_18914);
and U19100 (N_19100,N_18969,N_18682);
or U19101 (N_19101,N_18797,N_18837);
nand U19102 (N_19102,N_18937,N_18506);
xor U19103 (N_19103,N_18688,N_18757);
nor U19104 (N_19104,N_18843,N_18769);
or U19105 (N_19105,N_18881,N_18882);
and U19106 (N_19106,N_18526,N_18539);
xnor U19107 (N_19107,N_18924,N_18860);
or U19108 (N_19108,N_18690,N_18884);
or U19109 (N_19109,N_18840,N_18639);
and U19110 (N_19110,N_18824,N_18950);
or U19111 (N_19111,N_18891,N_18764);
nor U19112 (N_19112,N_18942,N_18511);
nor U19113 (N_19113,N_18711,N_18958);
xnor U19114 (N_19114,N_18522,N_18533);
nand U19115 (N_19115,N_18626,N_18932);
or U19116 (N_19116,N_18579,N_18727);
and U19117 (N_19117,N_18927,N_18636);
xnor U19118 (N_19118,N_18669,N_18993);
and U19119 (N_19119,N_18662,N_18734);
nand U19120 (N_19120,N_18954,N_18982);
nor U19121 (N_19121,N_18633,N_18855);
nand U19122 (N_19122,N_18862,N_18951);
nor U19123 (N_19123,N_18904,N_18706);
or U19124 (N_19124,N_18800,N_18965);
and U19125 (N_19125,N_18656,N_18962);
nand U19126 (N_19126,N_18900,N_18968);
nand U19127 (N_19127,N_18859,N_18894);
nand U19128 (N_19128,N_18986,N_18692);
xor U19129 (N_19129,N_18685,N_18970);
nor U19130 (N_19130,N_18818,N_18675);
xnor U19131 (N_19131,N_18575,N_18780);
nand U19132 (N_19132,N_18615,N_18940);
nand U19133 (N_19133,N_18966,N_18632);
nor U19134 (N_19134,N_18565,N_18570);
nor U19135 (N_19135,N_18777,N_18826);
and U19136 (N_19136,N_18999,N_18592);
xnor U19137 (N_19137,N_18919,N_18761);
or U19138 (N_19138,N_18566,N_18890);
nor U19139 (N_19139,N_18528,N_18863);
nand U19140 (N_19140,N_18714,N_18679);
and U19141 (N_19141,N_18696,N_18985);
and U19142 (N_19142,N_18752,N_18994);
and U19143 (N_19143,N_18686,N_18939);
nor U19144 (N_19144,N_18530,N_18560);
nand U19145 (N_19145,N_18746,N_18917);
nand U19146 (N_19146,N_18550,N_18598);
or U19147 (N_19147,N_18870,N_18812);
and U19148 (N_19148,N_18846,N_18756);
nor U19149 (N_19149,N_18848,N_18957);
nor U19150 (N_19150,N_18786,N_18838);
or U19151 (N_19151,N_18907,N_18955);
or U19152 (N_19152,N_18886,N_18755);
and U19153 (N_19153,N_18667,N_18589);
and U19154 (N_19154,N_18754,N_18938);
nor U19155 (N_19155,N_18787,N_18724);
nand U19156 (N_19156,N_18658,N_18603);
or U19157 (N_19157,N_18708,N_18821);
or U19158 (N_19158,N_18563,N_18627);
or U19159 (N_19159,N_18555,N_18540);
xnor U19160 (N_19160,N_18743,N_18829);
or U19161 (N_19161,N_18793,N_18931);
nor U19162 (N_19162,N_18853,N_18520);
nand U19163 (N_19163,N_18813,N_18542);
and U19164 (N_19164,N_18715,N_18718);
xnor U19165 (N_19165,N_18759,N_18952);
xor U19166 (N_19166,N_18804,N_18834);
and U19167 (N_19167,N_18809,N_18594);
or U19168 (N_19168,N_18795,N_18537);
nor U19169 (N_19169,N_18504,N_18561);
xnor U19170 (N_19170,N_18652,N_18507);
and U19171 (N_19171,N_18781,N_18680);
and U19172 (N_19172,N_18609,N_18973);
or U19173 (N_19173,N_18803,N_18624);
nor U19174 (N_19174,N_18857,N_18817);
nand U19175 (N_19175,N_18613,N_18825);
nor U19176 (N_19176,N_18733,N_18600);
nand U19177 (N_19177,N_18869,N_18822);
or U19178 (N_19178,N_18500,N_18810);
nand U19179 (N_19179,N_18981,N_18704);
nand U19180 (N_19180,N_18959,N_18749);
and U19181 (N_19181,N_18748,N_18604);
nand U19182 (N_19182,N_18571,N_18783);
nand U19183 (N_19183,N_18935,N_18534);
xnor U19184 (N_19184,N_18701,N_18646);
nor U19185 (N_19185,N_18634,N_18630);
or U19186 (N_19186,N_18535,N_18668);
nor U19187 (N_19187,N_18713,N_18586);
nor U19188 (N_19188,N_18687,N_18660);
nor U19189 (N_19189,N_18702,N_18741);
xnor U19190 (N_19190,N_18607,N_18961);
or U19191 (N_19191,N_18880,N_18925);
xnor U19192 (N_19192,N_18788,N_18663);
and U19193 (N_19193,N_18974,N_18577);
or U19194 (N_19194,N_18830,N_18631);
nor U19195 (N_19195,N_18814,N_18618);
nand U19196 (N_19196,N_18799,N_18541);
nor U19197 (N_19197,N_18902,N_18779);
nor U19198 (N_19198,N_18910,N_18543);
nor U19199 (N_19199,N_18576,N_18548);
or U19200 (N_19200,N_18661,N_18653);
xnor U19201 (N_19201,N_18972,N_18964);
and U19202 (N_19202,N_18996,N_18512);
nor U19203 (N_19203,N_18549,N_18595);
and U19204 (N_19204,N_18642,N_18581);
nor U19205 (N_19205,N_18879,N_18901);
and U19206 (N_19206,N_18716,N_18730);
and U19207 (N_19207,N_18823,N_18791);
nand U19208 (N_19208,N_18593,N_18854);
xnor U19209 (N_19209,N_18683,N_18614);
nor U19210 (N_19210,N_18949,N_18657);
or U19211 (N_19211,N_18856,N_18712);
or U19212 (N_19212,N_18877,N_18742);
and U19213 (N_19213,N_18558,N_18544);
xor U19214 (N_19214,N_18721,N_18710);
nand U19215 (N_19215,N_18858,N_18574);
nand U19216 (N_19216,N_18674,N_18865);
nor U19217 (N_19217,N_18953,N_18998);
nand U19218 (N_19218,N_18806,N_18651);
or U19219 (N_19219,N_18909,N_18616);
or U19220 (N_19220,N_18623,N_18736);
or U19221 (N_19221,N_18967,N_18580);
and U19222 (N_19222,N_18872,N_18635);
nor U19223 (N_19223,N_18559,N_18510);
nand U19224 (N_19224,N_18946,N_18699);
or U19225 (N_19225,N_18672,N_18640);
nor U19226 (N_19226,N_18845,N_18502);
or U19227 (N_19227,N_18851,N_18599);
or U19228 (N_19228,N_18673,N_18921);
and U19229 (N_19229,N_18906,N_18698);
and U19230 (N_19230,N_18659,N_18943);
nand U19231 (N_19231,N_18975,N_18778);
nor U19232 (N_19232,N_18744,N_18762);
or U19233 (N_19233,N_18554,N_18524);
nand U19234 (N_19234,N_18695,N_18583);
nand U19235 (N_19235,N_18515,N_18805);
nand U19236 (N_19236,N_18933,N_18903);
nor U19237 (N_19237,N_18776,N_18978);
nor U19238 (N_19238,N_18852,N_18898);
nor U19239 (N_19239,N_18567,N_18725);
xor U19240 (N_19240,N_18767,N_18641);
nor U19241 (N_19241,N_18926,N_18947);
or U19242 (N_19242,N_18833,N_18514);
nand U19243 (N_19243,N_18782,N_18689);
and U19244 (N_19244,N_18647,N_18866);
or U19245 (N_19245,N_18828,N_18905);
nand U19246 (N_19246,N_18977,N_18995);
nor U19247 (N_19247,N_18912,N_18650);
and U19248 (N_19248,N_18808,N_18747);
or U19249 (N_19249,N_18516,N_18606);
and U19250 (N_19250,N_18980,N_18550);
nand U19251 (N_19251,N_18762,N_18544);
xnor U19252 (N_19252,N_18738,N_18709);
and U19253 (N_19253,N_18616,N_18529);
xor U19254 (N_19254,N_18897,N_18693);
or U19255 (N_19255,N_18595,N_18917);
and U19256 (N_19256,N_18911,N_18674);
nor U19257 (N_19257,N_18836,N_18802);
or U19258 (N_19258,N_18505,N_18697);
nand U19259 (N_19259,N_18795,N_18808);
nor U19260 (N_19260,N_18961,N_18895);
xnor U19261 (N_19261,N_18887,N_18816);
and U19262 (N_19262,N_18727,N_18916);
and U19263 (N_19263,N_18808,N_18859);
nor U19264 (N_19264,N_18655,N_18905);
xnor U19265 (N_19265,N_18800,N_18760);
and U19266 (N_19266,N_18706,N_18696);
xor U19267 (N_19267,N_18731,N_18813);
or U19268 (N_19268,N_18782,N_18711);
nand U19269 (N_19269,N_18706,N_18867);
nor U19270 (N_19270,N_18548,N_18666);
nand U19271 (N_19271,N_18661,N_18776);
and U19272 (N_19272,N_18747,N_18950);
and U19273 (N_19273,N_18951,N_18781);
xor U19274 (N_19274,N_18696,N_18866);
nand U19275 (N_19275,N_18811,N_18508);
nand U19276 (N_19276,N_18766,N_18673);
xnor U19277 (N_19277,N_18520,N_18979);
nor U19278 (N_19278,N_18866,N_18520);
xnor U19279 (N_19279,N_18592,N_18581);
nand U19280 (N_19280,N_18946,N_18795);
nand U19281 (N_19281,N_18555,N_18908);
or U19282 (N_19282,N_18554,N_18729);
nand U19283 (N_19283,N_18893,N_18944);
nand U19284 (N_19284,N_18926,N_18912);
and U19285 (N_19285,N_18905,N_18842);
xnor U19286 (N_19286,N_18544,N_18872);
nor U19287 (N_19287,N_18807,N_18833);
nor U19288 (N_19288,N_18859,N_18520);
xor U19289 (N_19289,N_18973,N_18869);
or U19290 (N_19290,N_18620,N_18993);
nand U19291 (N_19291,N_18702,N_18595);
or U19292 (N_19292,N_18904,N_18963);
nand U19293 (N_19293,N_18711,N_18974);
or U19294 (N_19294,N_18643,N_18716);
nand U19295 (N_19295,N_18517,N_18864);
or U19296 (N_19296,N_18830,N_18504);
or U19297 (N_19297,N_18988,N_18987);
nand U19298 (N_19298,N_18892,N_18924);
or U19299 (N_19299,N_18979,N_18600);
or U19300 (N_19300,N_18571,N_18888);
nand U19301 (N_19301,N_18707,N_18744);
or U19302 (N_19302,N_18877,N_18940);
xnor U19303 (N_19303,N_18575,N_18805);
and U19304 (N_19304,N_18633,N_18843);
and U19305 (N_19305,N_18751,N_18955);
nor U19306 (N_19306,N_18939,N_18935);
xnor U19307 (N_19307,N_18965,N_18765);
and U19308 (N_19308,N_18631,N_18619);
xnor U19309 (N_19309,N_18675,N_18792);
xnor U19310 (N_19310,N_18867,N_18668);
or U19311 (N_19311,N_18995,N_18602);
and U19312 (N_19312,N_18726,N_18521);
or U19313 (N_19313,N_18812,N_18659);
xnor U19314 (N_19314,N_18800,N_18804);
and U19315 (N_19315,N_18886,N_18602);
and U19316 (N_19316,N_18536,N_18586);
nor U19317 (N_19317,N_18607,N_18930);
nor U19318 (N_19318,N_18652,N_18687);
nor U19319 (N_19319,N_18624,N_18639);
or U19320 (N_19320,N_18674,N_18707);
xor U19321 (N_19321,N_18507,N_18799);
nand U19322 (N_19322,N_18714,N_18916);
or U19323 (N_19323,N_18772,N_18574);
nor U19324 (N_19324,N_18722,N_18823);
nand U19325 (N_19325,N_18988,N_18521);
xor U19326 (N_19326,N_18764,N_18973);
nor U19327 (N_19327,N_18753,N_18886);
nor U19328 (N_19328,N_18519,N_18714);
nand U19329 (N_19329,N_18874,N_18697);
and U19330 (N_19330,N_18803,N_18870);
xor U19331 (N_19331,N_18655,N_18507);
or U19332 (N_19332,N_18651,N_18776);
xor U19333 (N_19333,N_18970,N_18936);
nand U19334 (N_19334,N_18745,N_18755);
nand U19335 (N_19335,N_18964,N_18878);
and U19336 (N_19336,N_18564,N_18808);
xnor U19337 (N_19337,N_18797,N_18690);
and U19338 (N_19338,N_18832,N_18754);
nor U19339 (N_19339,N_18917,N_18554);
and U19340 (N_19340,N_18693,N_18738);
or U19341 (N_19341,N_18716,N_18604);
xor U19342 (N_19342,N_18920,N_18878);
nand U19343 (N_19343,N_18938,N_18682);
nor U19344 (N_19344,N_18561,N_18708);
nand U19345 (N_19345,N_18921,N_18742);
or U19346 (N_19346,N_18662,N_18595);
and U19347 (N_19347,N_18890,N_18610);
xnor U19348 (N_19348,N_18685,N_18739);
nor U19349 (N_19349,N_18620,N_18593);
xnor U19350 (N_19350,N_18599,N_18646);
nor U19351 (N_19351,N_18883,N_18820);
or U19352 (N_19352,N_18622,N_18515);
or U19353 (N_19353,N_18856,N_18616);
and U19354 (N_19354,N_18674,N_18628);
and U19355 (N_19355,N_18533,N_18905);
or U19356 (N_19356,N_18622,N_18502);
and U19357 (N_19357,N_18832,N_18981);
nand U19358 (N_19358,N_18715,N_18722);
nor U19359 (N_19359,N_18991,N_18512);
nand U19360 (N_19360,N_18750,N_18541);
nor U19361 (N_19361,N_18735,N_18777);
or U19362 (N_19362,N_18860,N_18541);
nand U19363 (N_19363,N_18674,N_18607);
xor U19364 (N_19364,N_18617,N_18826);
nor U19365 (N_19365,N_18847,N_18944);
or U19366 (N_19366,N_18548,N_18601);
or U19367 (N_19367,N_18704,N_18664);
nor U19368 (N_19368,N_18985,N_18663);
and U19369 (N_19369,N_18639,N_18815);
and U19370 (N_19370,N_18868,N_18508);
or U19371 (N_19371,N_18893,N_18618);
and U19372 (N_19372,N_18718,N_18716);
or U19373 (N_19373,N_18511,N_18999);
or U19374 (N_19374,N_18926,N_18969);
xnor U19375 (N_19375,N_18622,N_18847);
nor U19376 (N_19376,N_18965,N_18662);
nand U19377 (N_19377,N_18608,N_18910);
nor U19378 (N_19378,N_18754,N_18828);
or U19379 (N_19379,N_18888,N_18988);
xor U19380 (N_19380,N_18683,N_18826);
nor U19381 (N_19381,N_18896,N_18731);
xor U19382 (N_19382,N_18784,N_18633);
or U19383 (N_19383,N_18685,N_18742);
or U19384 (N_19384,N_18882,N_18691);
xnor U19385 (N_19385,N_18680,N_18827);
and U19386 (N_19386,N_18860,N_18896);
xor U19387 (N_19387,N_18687,N_18773);
nor U19388 (N_19388,N_18977,N_18507);
xnor U19389 (N_19389,N_18501,N_18807);
and U19390 (N_19390,N_18995,N_18885);
xnor U19391 (N_19391,N_18848,N_18977);
or U19392 (N_19392,N_18754,N_18712);
or U19393 (N_19393,N_18729,N_18556);
nand U19394 (N_19394,N_18962,N_18561);
and U19395 (N_19395,N_18552,N_18556);
nand U19396 (N_19396,N_18584,N_18509);
xnor U19397 (N_19397,N_18903,N_18779);
nor U19398 (N_19398,N_18974,N_18786);
or U19399 (N_19399,N_18918,N_18624);
nor U19400 (N_19400,N_18766,N_18707);
or U19401 (N_19401,N_18946,N_18786);
nand U19402 (N_19402,N_18533,N_18917);
nor U19403 (N_19403,N_18677,N_18962);
nor U19404 (N_19404,N_18787,N_18755);
xnor U19405 (N_19405,N_18920,N_18881);
and U19406 (N_19406,N_18956,N_18589);
nand U19407 (N_19407,N_18656,N_18997);
nand U19408 (N_19408,N_18573,N_18568);
nor U19409 (N_19409,N_18731,N_18891);
xnor U19410 (N_19410,N_18563,N_18829);
or U19411 (N_19411,N_18596,N_18977);
or U19412 (N_19412,N_18849,N_18708);
and U19413 (N_19413,N_18578,N_18990);
or U19414 (N_19414,N_18755,N_18860);
or U19415 (N_19415,N_18777,N_18726);
xor U19416 (N_19416,N_18638,N_18592);
or U19417 (N_19417,N_18632,N_18697);
or U19418 (N_19418,N_18874,N_18987);
and U19419 (N_19419,N_18572,N_18776);
and U19420 (N_19420,N_18696,N_18555);
nand U19421 (N_19421,N_18967,N_18635);
and U19422 (N_19422,N_18558,N_18873);
or U19423 (N_19423,N_18710,N_18604);
nand U19424 (N_19424,N_18953,N_18825);
nand U19425 (N_19425,N_18669,N_18626);
nor U19426 (N_19426,N_18776,N_18806);
and U19427 (N_19427,N_18758,N_18975);
nand U19428 (N_19428,N_18838,N_18873);
xor U19429 (N_19429,N_18729,N_18598);
nand U19430 (N_19430,N_18647,N_18641);
nand U19431 (N_19431,N_18769,N_18674);
or U19432 (N_19432,N_18560,N_18545);
and U19433 (N_19433,N_18655,N_18868);
xor U19434 (N_19434,N_18874,N_18632);
xnor U19435 (N_19435,N_18787,N_18703);
and U19436 (N_19436,N_18609,N_18671);
or U19437 (N_19437,N_18632,N_18734);
nor U19438 (N_19438,N_18765,N_18552);
or U19439 (N_19439,N_18745,N_18666);
xnor U19440 (N_19440,N_18714,N_18819);
and U19441 (N_19441,N_18762,N_18873);
or U19442 (N_19442,N_18953,N_18968);
xnor U19443 (N_19443,N_18979,N_18664);
or U19444 (N_19444,N_18685,N_18794);
xnor U19445 (N_19445,N_18877,N_18552);
or U19446 (N_19446,N_18982,N_18804);
and U19447 (N_19447,N_18784,N_18723);
nand U19448 (N_19448,N_18710,N_18600);
nand U19449 (N_19449,N_18854,N_18642);
nor U19450 (N_19450,N_18997,N_18983);
and U19451 (N_19451,N_18765,N_18798);
nand U19452 (N_19452,N_18872,N_18936);
or U19453 (N_19453,N_18891,N_18569);
or U19454 (N_19454,N_18523,N_18857);
nor U19455 (N_19455,N_18715,N_18767);
nand U19456 (N_19456,N_18848,N_18602);
or U19457 (N_19457,N_18844,N_18867);
nand U19458 (N_19458,N_18838,N_18618);
nor U19459 (N_19459,N_18818,N_18697);
nor U19460 (N_19460,N_18731,N_18965);
and U19461 (N_19461,N_18957,N_18956);
nand U19462 (N_19462,N_18587,N_18722);
nand U19463 (N_19463,N_18720,N_18992);
or U19464 (N_19464,N_18634,N_18537);
and U19465 (N_19465,N_18994,N_18663);
nand U19466 (N_19466,N_18661,N_18538);
and U19467 (N_19467,N_18867,N_18625);
nor U19468 (N_19468,N_18655,N_18569);
nor U19469 (N_19469,N_18548,N_18787);
and U19470 (N_19470,N_18685,N_18868);
and U19471 (N_19471,N_18819,N_18716);
nand U19472 (N_19472,N_18588,N_18612);
and U19473 (N_19473,N_18792,N_18610);
and U19474 (N_19474,N_18853,N_18977);
nand U19475 (N_19475,N_18572,N_18576);
xor U19476 (N_19476,N_18882,N_18808);
and U19477 (N_19477,N_18719,N_18937);
and U19478 (N_19478,N_18584,N_18706);
nand U19479 (N_19479,N_18997,N_18786);
and U19480 (N_19480,N_18525,N_18615);
or U19481 (N_19481,N_18898,N_18910);
nand U19482 (N_19482,N_18540,N_18802);
nor U19483 (N_19483,N_18661,N_18782);
and U19484 (N_19484,N_18984,N_18558);
or U19485 (N_19485,N_18690,N_18900);
or U19486 (N_19486,N_18795,N_18534);
or U19487 (N_19487,N_18848,N_18698);
nand U19488 (N_19488,N_18804,N_18706);
nand U19489 (N_19489,N_18593,N_18877);
nor U19490 (N_19490,N_18629,N_18557);
or U19491 (N_19491,N_18684,N_18781);
nor U19492 (N_19492,N_18755,N_18560);
xor U19493 (N_19493,N_18686,N_18918);
nor U19494 (N_19494,N_18975,N_18984);
nand U19495 (N_19495,N_18980,N_18803);
nor U19496 (N_19496,N_18513,N_18746);
and U19497 (N_19497,N_18563,N_18666);
and U19498 (N_19498,N_18912,N_18622);
or U19499 (N_19499,N_18664,N_18829);
and U19500 (N_19500,N_19026,N_19323);
or U19501 (N_19501,N_19479,N_19311);
nor U19502 (N_19502,N_19252,N_19031);
xor U19503 (N_19503,N_19380,N_19240);
nor U19504 (N_19504,N_19467,N_19263);
nor U19505 (N_19505,N_19387,N_19146);
and U19506 (N_19506,N_19207,N_19312);
or U19507 (N_19507,N_19091,N_19435);
nor U19508 (N_19508,N_19158,N_19102);
xor U19509 (N_19509,N_19454,N_19266);
xnor U19510 (N_19510,N_19292,N_19147);
or U19511 (N_19511,N_19044,N_19217);
nor U19512 (N_19512,N_19249,N_19388);
or U19513 (N_19513,N_19237,N_19081);
nand U19514 (N_19514,N_19112,N_19144);
or U19515 (N_19515,N_19153,N_19104);
nor U19516 (N_19516,N_19012,N_19325);
or U19517 (N_19517,N_19185,N_19346);
nor U19518 (N_19518,N_19087,N_19481);
or U19519 (N_19519,N_19241,N_19462);
nor U19520 (N_19520,N_19072,N_19428);
and U19521 (N_19521,N_19291,N_19353);
nand U19522 (N_19522,N_19315,N_19403);
or U19523 (N_19523,N_19352,N_19086);
xnor U19524 (N_19524,N_19351,N_19334);
nor U19525 (N_19525,N_19420,N_19362);
xor U19526 (N_19526,N_19431,N_19290);
xor U19527 (N_19527,N_19494,N_19399);
xnor U19528 (N_19528,N_19423,N_19140);
nor U19529 (N_19529,N_19269,N_19160);
and U19530 (N_19530,N_19302,N_19294);
xor U19531 (N_19531,N_19247,N_19298);
or U19532 (N_19532,N_19386,N_19344);
and U19533 (N_19533,N_19177,N_19011);
and U19534 (N_19534,N_19119,N_19490);
or U19535 (N_19535,N_19131,N_19054);
and U19536 (N_19536,N_19201,N_19022);
xnor U19537 (N_19537,N_19114,N_19264);
and U19538 (N_19538,N_19464,N_19169);
xor U19539 (N_19539,N_19419,N_19200);
nand U19540 (N_19540,N_19330,N_19157);
nor U19541 (N_19541,N_19198,N_19239);
nor U19542 (N_19542,N_19125,N_19190);
nand U19543 (N_19543,N_19371,N_19337);
xor U19544 (N_19544,N_19191,N_19324);
xnor U19545 (N_19545,N_19405,N_19111);
and U19546 (N_19546,N_19331,N_19329);
xnor U19547 (N_19547,N_19159,N_19393);
nor U19548 (N_19548,N_19375,N_19484);
nand U19549 (N_19549,N_19354,N_19376);
and U19550 (N_19550,N_19345,N_19439);
nand U19551 (N_19551,N_19016,N_19128);
nand U19552 (N_19552,N_19360,N_19283);
or U19553 (N_19553,N_19332,N_19094);
or U19554 (N_19554,N_19361,N_19305);
xor U19555 (N_19555,N_19052,N_19426);
xnor U19556 (N_19556,N_19414,N_19219);
nand U19557 (N_19557,N_19412,N_19319);
and U19558 (N_19558,N_19055,N_19188);
nor U19559 (N_19559,N_19434,N_19476);
nor U19560 (N_19560,N_19355,N_19372);
and U19561 (N_19561,N_19316,N_19304);
or U19562 (N_19562,N_19127,N_19489);
xor U19563 (N_19563,N_19058,N_19042);
xor U19564 (N_19564,N_19411,N_19167);
nor U19565 (N_19565,N_19450,N_19232);
nand U19566 (N_19566,N_19041,N_19357);
or U19567 (N_19567,N_19129,N_19113);
nand U19568 (N_19568,N_19027,N_19152);
nor U19569 (N_19569,N_19203,N_19233);
or U19570 (N_19570,N_19416,N_19370);
nand U19571 (N_19571,N_19229,N_19069);
nand U19572 (N_19572,N_19262,N_19496);
and U19573 (N_19573,N_19101,N_19289);
nand U19574 (N_19574,N_19183,N_19024);
nor U19575 (N_19575,N_19451,N_19231);
and U19576 (N_19576,N_19075,N_19347);
nand U19577 (N_19577,N_19488,N_19400);
nand U19578 (N_19578,N_19299,N_19084);
or U19579 (N_19579,N_19422,N_19491);
xnor U19580 (N_19580,N_19452,N_19222);
nor U19581 (N_19581,N_19076,N_19130);
nor U19582 (N_19582,N_19401,N_19336);
nor U19583 (N_19583,N_19214,N_19463);
and U19584 (N_19584,N_19293,N_19477);
nor U19585 (N_19585,N_19327,N_19482);
and U19586 (N_19586,N_19342,N_19381);
nand U19587 (N_19587,N_19155,N_19339);
nand U19588 (N_19588,N_19060,N_19284);
xor U19589 (N_19589,N_19065,N_19341);
xnor U19590 (N_19590,N_19030,N_19040);
nand U19591 (N_19591,N_19097,N_19404);
and U19592 (N_19592,N_19449,N_19138);
or U19593 (N_19593,N_19338,N_19103);
xnor U19594 (N_19594,N_19215,N_19279);
xor U19595 (N_19595,N_19020,N_19132);
and U19596 (N_19596,N_19460,N_19322);
nor U19597 (N_19597,N_19088,N_19184);
xnor U19598 (N_19598,N_19124,N_19073);
and U19599 (N_19599,N_19048,N_19406);
nand U19600 (N_19600,N_19270,N_19303);
nand U19601 (N_19601,N_19106,N_19250);
nand U19602 (N_19602,N_19261,N_19164);
nand U19603 (N_19603,N_19213,N_19333);
or U19604 (N_19604,N_19095,N_19487);
xor U19605 (N_19605,N_19149,N_19037);
nand U19606 (N_19606,N_19377,N_19282);
or U19607 (N_19607,N_19390,N_19474);
nor U19608 (N_19608,N_19363,N_19443);
nor U19609 (N_19609,N_19246,N_19326);
xnor U19610 (N_19610,N_19179,N_19046);
xnor U19611 (N_19611,N_19335,N_19468);
and U19612 (N_19612,N_19078,N_19227);
nand U19613 (N_19613,N_19062,N_19135);
xnor U19614 (N_19614,N_19275,N_19458);
nor U19615 (N_19615,N_19225,N_19154);
and U19616 (N_19616,N_19015,N_19145);
xor U19617 (N_19617,N_19417,N_19243);
or U19618 (N_19618,N_19379,N_19456);
nor U19619 (N_19619,N_19409,N_19485);
xor U19620 (N_19620,N_19259,N_19083);
xor U19621 (N_19621,N_19441,N_19396);
or U19622 (N_19622,N_19483,N_19133);
nand U19623 (N_19623,N_19093,N_19358);
or U19624 (N_19624,N_19096,N_19067);
nand U19625 (N_19625,N_19457,N_19415);
and U19626 (N_19626,N_19170,N_19236);
nand U19627 (N_19627,N_19445,N_19018);
nor U19628 (N_19628,N_19123,N_19430);
or U19629 (N_19629,N_19189,N_19107);
nor U19630 (N_19630,N_19465,N_19121);
and U19631 (N_19631,N_19251,N_19308);
and U19632 (N_19632,N_19148,N_19005);
nand U19633 (N_19633,N_19221,N_19255);
xnor U19634 (N_19634,N_19173,N_19367);
xor U19635 (N_19635,N_19014,N_19118);
or U19636 (N_19636,N_19009,N_19265);
nor U19637 (N_19637,N_19176,N_19280);
xnor U19638 (N_19638,N_19180,N_19248);
nor U19639 (N_19639,N_19021,N_19023);
nand U19640 (N_19640,N_19134,N_19204);
nor U19641 (N_19641,N_19056,N_19318);
xnor U19642 (N_19642,N_19492,N_19074);
or U19643 (N_19643,N_19100,N_19090);
or U19644 (N_19644,N_19306,N_19359);
nor U19645 (N_19645,N_19080,N_19427);
nor U19646 (N_19646,N_19286,N_19410);
nand U19647 (N_19647,N_19394,N_19013);
xnor U19648 (N_19648,N_19071,N_19234);
nand U19649 (N_19649,N_19008,N_19116);
nor U19650 (N_19650,N_19475,N_19373);
or U19651 (N_19651,N_19493,N_19092);
nor U19652 (N_19652,N_19230,N_19307);
xor U19653 (N_19653,N_19003,N_19010);
and U19654 (N_19654,N_19182,N_19105);
xor U19655 (N_19655,N_19047,N_19421);
or U19656 (N_19656,N_19137,N_19235);
xnor U19657 (N_19657,N_19453,N_19288);
or U19658 (N_19658,N_19006,N_19274);
and U19659 (N_19659,N_19163,N_19385);
nor U19660 (N_19660,N_19068,N_19444);
nand U19661 (N_19661,N_19098,N_19099);
or U19662 (N_19662,N_19328,N_19079);
xor U19663 (N_19663,N_19195,N_19402);
and U19664 (N_19664,N_19199,N_19242);
or U19665 (N_19665,N_19271,N_19036);
or U19666 (N_19666,N_19254,N_19178);
and U19667 (N_19667,N_19424,N_19438);
or U19668 (N_19668,N_19001,N_19368);
nor U19669 (N_19669,N_19193,N_19117);
nand U19670 (N_19670,N_19181,N_19162);
nor U19671 (N_19671,N_19066,N_19126);
nand U19672 (N_19672,N_19343,N_19161);
nand U19673 (N_19673,N_19407,N_19077);
nor U19674 (N_19674,N_19122,N_19142);
and U19675 (N_19675,N_19209,N_19166);
xor U19676 (N_19676,N_19287,N_19448);
or U19677 (N_19677,N_19436,N_19043);
xnor U19678 (N_19678,N_19466,N_19057);
nor U19679 (N_19679,N_19150,N_19297);
nor U19680 (N_19680,N_19384,N_19143);
and U19681 (N_19681,N_19019,N_19267);
nor U19682 (N_19682,N_19413,N_19038);
nor U19683 (N_19683,N_19408,N_19309);
nand U19684 (N_19684,N_19473,N_19165);
nor U19685 (N_19685,N_19244,N_19320);
nor U19686 (N_19686,N_19418,N_19211);
or U19687 (N_19687,N_19224,N_19349);
xnor U19688 (N_19688,N_19389,N_19470);
or U19689 (N_19689,N_19273,N_19205);
xnor U19690 (N_19690,N_19366,N_19356);
xnor U19691 (N_19691,N_19397,N_19197);
or U19692 (N_19692,N_19029,N_19398);
or U19693 (N_19693,N_19223,N_19051);
nor U19694 (N_19694,N_19480,N_19070);
or U19695 (N_19695,N_19032,N_19059);
and U19696 (N_19696,N_19002,N_19378);
nand U19697 (N_19697,N_19382,N_19141);
nand U19698 (N_19698,N_19256,N_19218);
and U19699 (N_19699,N_19478,N_19278);
and U19700 (N_19700,N_19272,N_19472);
xnor U19701 (N_19701,N_19257,N_19260);
nand U19702 (N_19702,N_19296,N_19208);
xor U19703 (N_19703,N_19364,N_19447);
nand U19704 (N_19704,N_19391,N_19168);
nor U19705 (N_19705,N_19295,N_19455);
nand U19706 (N_19706,N_19108,N_19499);
nor U19707 (N_19707,N_19238,N_19471);
and U19708 (N_19708,N_19035,N_19365);
nor U19709 (N_19709,N_19245,N_19082);
or U19710 (N_19710,N_19025,N_19039);
or U19711 (N_19711,N_19063,N_19210);
xnor U19712 (N_19712,N_19432,N_19350);
or U19713 (N_19713,N_19253,N_19392);
xor U19714 (N_19714,N_19175,N_19301);
xor U19715 (N_19715,N_19212,N_19061);
nor U19716 (N_19716,N_19498,N_19045);
or U19717 (N_19717,N_19226,N_19429);
nor U19718 (N_19718,N_19276,N_19139);
xor U19719 (N_19719,N_19194,N_19192);
xnor U19720 (N_19720,N_19085,N_19425);
and U19721 (N_19721,N_19268,N_19136);
or U19722 (N_19722,N_19442,N_19050);
xnor U19723 (N_19723,N_19258,N_19053);
and U19724 (N_19724,N_19348,N_19433);
nor U19725 (N_19725,N_19300,N_19310);
or U19726 (N_19726,N_19115,N_19110);
xnor U19727 (N_19727,N_19196,N_19395);
xnor U19728 (N_19728,N_19109,N_19172);
xor U19729 (N_19729,N_19446,N_19277);
or U19730 (N_19730,N_19437,N_19187);
xor U19731 (N_19731,N_19033,N_19028);
or U19732 (N_19732,N_19461,N_19049);
xnor U19733 (N_19733,N_19034,N_19228);
nand U19734 (N_19734,N_19007,N_19000);
nor U19735 (N_19735,N_19314,N_19369);
or U19736 (N_19736,N_19216,N_19374);
nor U19737 (N_19737,N_19004,N_19340);
and U19738 (N_19738,N_19469,N_19151);
nand U19739 (N_19739,N_19440,N_19120);
xnor U19740 (N_19740,N_19486,N_19156);
and U19741 (N_19741,N_19202,N_19171);
nand U19742 (N_19742,N_19285,N_19206);
nand U19743 (N_19743,N_19495,N_19089);
xnor U19744 (N_19744,N_19186,N_19281);
nor U19745 (N_19745,N_19064,N_19317);
or U19746 (N_19746,N_19220,N_19383);
nor U19747 (N_19747,N_19017,N_19174);
xor U19748 (N_19748,N_19459,N_19321);
nand U19749 (N_19749,N_19313,N_19497);
nor U19750 (N_19750,N_19491,N_19448);
and U19751 (N_19751,N_19259,N_19160);
or U19752 (N_19752,N_19198,N_19191);
or U19753 (N_19753,N_19449,N_19156);
or U19754 (N_19754,N_19288,N_19172);
nor U19755 (N_19755,N_19464,N_19140);
or U19756 (N_19756,N_19172,N_19132);
or U19757 (N_19757,N_19054,N_19276);
nor U19758 (N_19758,N_19118,N_19162);
nand U19759 (N_19759,N_19125,N_19305);
nor U19760 (N_19760,N_19371,N_19481);
nand U19761 (N_19761,N_19479,N_19340);
nor U19762 (N_19762,N_19112,N_19432);
or U19763 (N_19763,N_19033,N_19389);
and U19764 (N_19764,N_19312,N_19372);
and U19765 (N_19765,N_19437,N_19181);
nand U19766 (N_19766,N_19456,N_19477);
or U19767 (N_19767,N_19384,N_19111);
or U19768 (N_19768,N_19074,N_19253);
nand U19769 (N_19769,N_19212,N_19022);
and U19770 (N_19770,N_19419,N_19124);
nor U19771 (N_19771,N_19004,N_19391);
xor U19772 (N_19772,N_19074,N_19183);
nand U19773 (N_19773,N_19170,N_19226);
xnor U19774 (N_19774,N_19259,N_19009);
nand U19775 (N_19775,N_19462,N_19037);
nand U19776 (N_19776,N_19386,N_19475);
or U19777 (N_19777,N_19302,N_19438);
or U19778 (N_19778,N_19454,N_19160);
and U19779 (N_19779,N_19125,N_19282);
or U19780 (N_19780,N_19302,N_19410);
or U19781 (N_19781,N_19034,N_19269);
nor U19782 (N_19782,N_19145,N_19016);
or U19783 (N_19783,N_19200,N_19235);
nor U19784 (N_19784,N_19189,N_19496);
nand U19785 (N_19785,N_19274,N_19339);
nor U19786 (N_19786,N_19352,N_19251);
or U19787 (N_19787,N_19316,N_19200);
or U19788 (N_19788,N_19422,N_19198);
xor U19789 (N_19789,N_19475,N_19454);
or U19790 (N_19790,N_19118,N_19087);
nor U19791 (N_19791,N_19342,N_19202);
and U19792 (N_19792,N_19313,N_19457);
nor U19793 (N_19793,N_19185,N_19383);
xnor U19794 (N_19794,N_19246,N_19070);
and U19795 (N_19795,N_19243,N_19396);
nor U19796 (N_19796,N_19423,N_19295);
nand U19797 (N_19797,N_19381,N_19450);
xnor U19798 (N_19798,N_19229,N_19152);
or U19799 (N_19799,N_19107,N_19269);
or U19800 (N_19800,N_19245,N_19372);
nor U19801 (N_19801,N_19314,N_19177);
xnor U19802 (N_19802,N_19309,N_19335);
nor U19803 (N_19803,N_19351,N_19312);
xnor U19804 (N_19804,N_19257,N_19005);
and U19805 (N_19805,N_19420,N_19450);
nor U19806 (N_19806,N_19339,N_19372);
nand U19807 (N_19807,N_19349,N_19157);
nand U19808 (N_19808,N_19151,N_19452);
xnor U19809 (N_19809,N_19142,N_19287);
or U19810 (N_19810,N_19115,N_19171);
and U19811 (N_19811,N_19042,N_19017);
nor U19812 (N_19812,N_19018,N_19120);
and U19813 (N_19813,N_19207,N_19319);
xor U19814 (N_19814,N_19417,N_19416);
xnor U19815 (N_19815,N_19498,N_19179);
or U19816 (N_19816,N_19458,N_19262);
nand U19817 (N_19817,N_19360,N_19325);
nand U19818 (N_19818,N_19112,N_19371);
or U19819 (N_19819,N_19145,N_19403);
xnor U19820 (N_19820,N_19073,N_19158);
xor U19821 (N_19821,N_19401,N_19145);
and U19822 (N_19822,N_19390,N_19035);
and U19823 (N_19823,N_19058,N_19056);
nor U19824 (N_19824,N_19118,N_19013);
xnor U19825 (N_19825,N_19449,N_19342);
xor U19826 (N_19826,N_19413,N_19495);
xnor U19827 (N_19827,N_19240,N_19330);
and U19828 (N_19828,N_19360,N_19234);
and U19829 (N_19829,N_19130,N_19430);
xnor U19830 (N_19830,N_19113,N_19311);
or U19831 (N_19831,N_19193,N_19203);
or U19832 (N_19832,N_19266,N_19245);
xnor U19833 (N_19833,N_19420,N_19065);
nand U19834 (N_19834,N_19042,N_19410);
xor U19835 (N_19835,N_19066,N_19282);
xnor U19836 (N_19836,N_19323,N_19445);
xnor U19837 (N_19837,N_19245,N_19278);
or U19838 (N_19838,N_19082,N_19290);
nor U19839 (N_19839,N_19134,N_19183);
nand U19840 (N_19840,N_19096,N_19175);
and U19841 (N_19841,N_19191,N_19090);
nand U19842 (N_19842,N_19308,N_19385);
nor U19843 (N_19843,N_19208,N_19212);
and U19844 (N_19844,N_19318,N_19417);
or U19845 (N_19845,N_19171,N_19481);
and U19846 (N_19846,N_19070,N_19148);
and U19847 (N_19847,N_19488,N_19474);
xnor U19848 (N_19848,N_19416,N_19356);
nand U19849 (N_19849,N_19148,N_19164);
nor U19850 (N_19850,N_19266,N_19384);
or U19851 (N_19851,N_19416,N_19151);
or U19852 (N_19852,N_19444,N_19063);
and U19853 (N_19853,N_19084,N_19200);
xor U19854 (N_19854,N_19291,N_19390);
xnor U19855 (N_19855,N_19021,N_19116);
nor U19856 (N_19856,N_19496,N_19245);
xor U19857 (N_19857,N_19178,N_19329);
nor U19858 (N_19858,N_19493,N_19174);
or U19859 (N_19859,N_19391,N_19082);
nor U19860 (N_19860,N_19475,N_19164);
nand U19861 (N_19861,N_19310,N_19012);
or U19862 (N_19862,N_19270,N_19460);
and U19863 (N_19863,N_19068,N_19399);
xor U19864 (N_19864,N_19138,N_19211);
xnor U19865 (N_19865,N_19192,N_19156);
nand U19866 (N_19866,N_19213,N_19327);
nor U19867 (N_19867,N_19454,N_19228);
nand U19868 (N_19868,N_19121,N_19199);
and U19869 (N_19869,N_19344,N_19339);
and U19870 (N_19870,N_19127,N_19047);
xnor U19871 (N_19871,N_19280,N_19278);
or U19872 (N_19872,N_19023,N_19493);
or U19873 (N_19873,N_19104,N_19428);
and U19874 (N_19874,N_19294,N_19355);
nor U19875 (N_19875,N_19184,N_19046);
nand U19876 (N_19876,N_19188,N_19271);
xnor U19877 (N_19877,N_19029,N_19022);
or U19878 (N_19878,N_19200,N_19379);
or U19879 (N_19879,N_19154,N_19291);
nor U19880 (N_19880,N_19492,N_19119);
or U19881 (N_19881,N_19306,N_19150);
or U19882 (N_19882,N_19226,N_19160);
nand U19883 (N_19883,N_19265,N_19324);
or U19884 (N_19884,N_19487,N_19107);
nor U19885 (N_19885,N_19368,N_19270);
nor U19886 (N_19886,N_19115,N_19037);
nand U19887 (N_19887,N_19424,N_19014);
nor U19888 (N_19888,N_19046,N_19228);
xnor U19889 (N_19889,N_19029,N_19323);
and U19890 (N_19890,N_19006,N_19304);
nand U19891 (N_19891,N_19457,N_19365);
xor U19892 (N_19892,N_19498,N_19008);
or U19893 (N_19893,N_19347,N_19171);
nand U19894 (N_19894,N_19335,N_19158);
or U19895 (N_19895,N_19040,N_19147);
nand U19896 (N_19896,N_19189,N_19173);
and U19897 (N_19897,N_19099,N_19302);
and U19898 (N_19898,N_19217,N_19116);
nor U19899 (N_19899,N_19123,N_19276);
xnor U19900 (N_19900,N_19204,N_19060);
nand U19901 (N_19901,N_19226,N_19126);
or U19902 (N_19902,N_19299,N_19356);
or U19903 (N_19903,N_19089,N_19058);
nor U19904 (N_19904,N_19176,N_19088);
nor U19905 (N_19905,N_19375,N_19158);
or U19906 (N_19906,N_19157,N_19256);
xor U19907 (N_19907,N_19175,N_19181);
nand U19908 (N_19908,N_19024,N_19058);
xnor U19909 (N_19909,N_19244,N_19055);
xor U19910 (N_19910,N_19386,N_19130);
nor U19911 (N_19911,N_19370,N_19016);
and U19912 (N_19912,N_19258,N_19314);
or U19913 (N_19913,N_19348,N_19403);
and U19914 (N_19914,N_19259,N_19168);
or U19915 (N_19915,N_19210,N_19049);
xor U19916 (N_19916,N_19436,N_19493);
xnor U19917 (N_19917,N_19370,N_19469);
or U19918 (N_19918,N_19041,N_19033);
nand U19919 (N_19919,N_19482,N_19324);
xnor U19920 (N_19920,N_19357,N_19196);
nor U19921 (N_19921,N_19100,N_19475);
or U19922 (N_19922,N_19048,N_19472);
and U19923 (N_19923,N_19061,N_19027);
nor U19924 (N_19924,N_19389,N_19320);
nor U19925 (N_19925,N_19497,N_19167);
nor U19926 (N_19926,N_19049,N_19307);
or U19927 (N_19927,N_19319,N_19084);
or U19928 (N_19928,N_19307,N_19207);
nand U19929 (N_19929,N_19005,N_19145);
nand U19930 (N_19930,N_19147,N_19054);
nand U19931 (N_19931,N_19148,N_19284);
nor U19932 (N_19932,N_19143,N_19387);
and U19933 (N_19933,N_19356,N_19072);
nor U19934 (N_19934,N_19110,N_19238);
nand U19935 (N_19935,N_19200,N_19227);
and U19936 (N_19936,N_19217,N_19335);
nor U19937 (N_19937,N_19475,N_19298);
or U19938 (N_19938,N_19437,N_19424);
xor U19939 (N_19939,N_19310,N_19363);
nand U19940 (N_19940,N_19453,N_19465);
xor U19941 (N_19941,N_19275,N_19153);
and U19942 (N_19942,N_19046,N_19318);
and U19943 (N_19943,N_19424,N_19000);
nor U19944 (N_19944,N_19100,N_19008);
and U19945 (N_19945,N_19190,N_19085);
nand U19946 (N_19946,N_19225,N_19398);
nor U19947 (N_19947,N_19276,N_19393);
xnor U19948 (N_19948,N_19102,N_19393);
nor U19949 (N_19949,N_19351,N_19484);
nand U19950 (N_19950,N_19039,N_19047);
and U19951 (N_19951,N_19483,N_19028);
nand U19952 (N_19952,N_19117,N_19374);
nand U19953 (N_19953,N_19410,N_19176);
nand U19954 (N_19954,N_19147,N_19216);
and U19955 (N_19955,N_19195,N_19465);
nor U19956 (N_19956,N_19074,N_19368);
xor U19957 (N_19957,N_19127,N_19110);
or U19958 (N_19958,N_19084,N_19263);
nor U19959 (N_19959,N_19050,N_19229);
or U19960 (N_19960,N_19041,N_19035);
nand U19961 (N_19961,N_19399,N_19225);
and U19962 (N_19962,N_19399,N_19431);
nor U19963 (N_19963,N_19190,N_19071);
xor U19964 (N_19964,N_19071,N_19481);
or U19965 (N_19965,N_19470,N_19355);
xor U19966 (N_19966,N_19432,N_19170);
nand U19967 (N_19967,N_19325,N_19477);
xnor U19968 (N_19968,N_19227,N_19002);
xnor U19969 (N_19969,N_19151,N_19027);
nor U19970 (N_19970,N_19207,N_19486);
or U19971 (N_19971,N_19428,N_19247);
nor U19972 (N_19972,N_19016,N_19088);
or U19973 (N_19973,N_19278,N_19160);
nand U19974 (N_19974,N_19046,N_19082);
or U19975 (N_19975,N_19390,N_19177);
xnor U19976 (N_19976,N_19297,N_19084);
xnor U19977 (N_19977,N_19025,N_19262);
xnor U19978 (N_19978,N_19392,N_19238);
xor U19979 (N_19979,N_19241,N_19409);
xor U19980 (N_19980,N_19259,N_19128);
nor U19981 (N_19981,N_19000,N_19356);
nand U19982 (N_19982,N_19126,N_19464);
and U19983 (N_19983,N_19458,N_19121);
nor U19984 (N_19984,N_19495,N_19048);
nor U19985 (N_19985,N_19396,N_19276);
xor U19986 (N_19986,N_19031,N_19416);
xor U19987 (N_19987,N_19055,N_19136);
nor U19988 (N_19988,N_19340,N_19484);
xnor U19989 (N_19989,N_19466,N_19290);
and U19990 (N_19990,N_19225,N_19262);
nor U19991 (N_19991,N_19484,N_19082);
or U19992 (N_19992,N_19430,N_19451);
nor U19993 (N_19993,N_19039,N_19447);
xor U19994 (N_19994,N_19104,N_19468);
nand U19995 (N_19995,N_19105,N_19236);
xor U19996 (N_19996,N_19330,N_19433);
nand U19997 (N_19997,N_19388,N_19434);
nand U19998 (N_19998,N_19149,N_19082);
nand U19999 (N_19999,N_19309,N_19356);
nand U20000 (N_20000,N_19734,N_19708);
and U20001 (N_20001,N_19595,N_19913);
and U20002 (N_20002,N_19728,N_19548);
or U20003 (N_20003,N_19550,N_19906);
nor U20004 (N_20004,N_19677,N_19912);
or U20005 (N_20005,N_19924,N_19710);
and U20006 (N_20006,N_19925,N_19732);
and U20007 (N_20007,N_19841,N_19524);
and U20008 (N_20008,N_19768,N_19500);
nand U20009 (N_20009,N_19773,N_19937);
or U20010 (N_20010,N_19558,N_19953);
nor U20011 (N_20011,N_19599,N_19598);
and U20012 (N_20012,N_19715,N_19613);
or U20013 (N_20013,N_19887,N_19752);
or U20014 (N_20014,N_19770,N_19765);
and U20015 (N_20015,N_19626,N_19895);
nor U20016 (N_20016,N_19898,N_19984);
xnor U20017 (N_20017,N_19956,N_19927);
or U20018 (N_20018,N_19657,N_19593);
and U20019 (N_20019,N_19608,N_19920);
and U20020 (N_20020,N_19838,N_19828);
xnor U20021 (N_20021,N_19746,N_19591);
and U20022 (N_20022,N_19871,N_19504);
and U20023 (N_20023,N_19645,N_19712);
or U20024 (N_20024,N_19809,N_19901);
and U20025 (N_20025,N_19823,N_19831);
xor U20026 (N_20026,N_19580,N_19826);
and U20027 (N_20027,N_19852,N_19982);
or U20028 (N_20028,N_19949,N_19606);
nor U20029 (N_20029,N_19569,N_19944);
or U20030 (N_20030,N_19618,N_19601);
xor U20031 (N_20031,N_19588,N_19857);
xor U20032 (N_20032,N_19989,N_19623);
xor U20033 (N_20033,N_19789,N_19876);
nand U20034 (N_20034,N_19691,N_19639);
nand U20035 (N_20035,N_19865,N_19885);
nand U20036 (N_20036,N_19836,N_19676);
and U20037 (N_20037,N_19635,N_19778);
xnor U20038 (N_20038,N_19573,N_19597);
nand U20039 (N_20039,N_19977,N_19519);
nand U20040 (N_20040,N_19510,N_19549);
xnor U20041 (N_20041,N_19681,N_19833);
and U20042 (N_20042,N_19614,N_19709);
xnor U20043 (N_20043,N_19941,N_19513);
nand U20044 (N_20044,N_19514,N_19859);
xnor U20045 (N_20045,N_19603,N_19667);
nor U20046 (N_20046,N_19653,N_19844);
xnor U20047 (N_20047,N_19747,N_19743);
nor U20048 (N_20048,N_19585,N_19769);
nand U20049 (N_20049,N_19738,N_19813);
nor U20050 (N_20050,N_19849,N_19629);
xnor U20051 (N_20051,N_19797,N_19783);
xor U20052 (N_20052,N_19867,N_19640);
xor U20053 (N_20053,N_19670,N_19915);
and U20054 (N_20054,N_19527,N_19731);
nand U20055 (N_20055,N_19707,N_19532);
or U20056 (N_20056,N_19794,N_19511);
xnor U20057 (N_20057,N_19586,N_19858);
nor U20058 (N_20058,N_19868,N_19897);
xnor U20059 (N_20059,N_19526,N_19753);
or U20060 (N_20060,N_19620,N_19754);
xnor U20061 (N_20061,N_19967,N_19525);
and U20062 (N_20062,N_19636,N_19922);
or U20063 (N_20063,N_19861,N_19911);
xnor U20064 (N_20064,N_19693,N_19520);
xnor U20065 (N_20065,N_19723,N_19751);
xnor U20066 (N_20066,N_19505,N_19733);
nand U20067 (N_20067,N_19624,N_19850);
xnor U20068 (N_20068,N_19604,N_19963);
nor U20069 (N_20069,N_19840,N_19980);
xor U20070 (N_20070,N_19530,N_19947);
and U20071 (N_20071,N_19725,N_19870);
xor U20072 (N_20072,N_19706,N_19909);
and U20073 (N_20073,N_19656,N_19946);
xor U20074 (N_20074,N_19684,N_19851);
and U20075 (N_20075,N_19966,N_19735);
nand U20076 (N_20076,N_19644,N_19687);
xnor U20077 (N_20077,N_19816,N_19805);
nand U20078 (N_20078,N_19843,N_19666);
or U20079 (N_20079,N_19531,N_19727);
xnor U20080 (N_20080,N_19631,N_19787);
nor U20081 (N_20081,N_19655,N_19560);
nand U20082 (N_20082,N_19506,N_19522);
nor U20083 (N_20083,N_19501,N_19570);
and U20084 (N_20084,N_19689,N_19641);
nor U20085 (N_20085,N_19786,N_19829);
or U20086 (N_20086,N_19943,N_19521);
xnor U20087 (N_20087,N_19772,N_19776);
xnor U20088 (N_20088,N_19929,N_19933);
nor U20089 (N_20089,N_19872,N_19975);
nand U20090 (N_20090,N_19779,N_19819);
nor U20091 (N_20091,N_19824,N_19875);
nor U20092 (N_20092,N_19996,N_19896);
nor U20093 (N_20093,N_19917,N_19874);
or U20094 (N_20094,N_19842,N_19811);
or U20095 (N_20095,N_19546,N_19716);
xor U20096 (N_20096,N_19694,N_19995);
nor U20097 (N_20097,N_19642,N_19860);
or U20098 (N_20098,N_19584,N_19916);
nand U20099 (N_20099,N_19942,N_19888);
or U20100 (N_20100,N_19990,N_19628);
xnor U20101 (N_20101,N_19955,N_19661);
or U20102 (N_20102,N_19638,N_19886);
nor U20103 (N_20103,N_19553,N_19780);
xor U20104 (N_20104,N_19965,N_19535);
nor U20105 (N_20105,N_19697,N_19722);
xnor U20106 (N_20106,N_19799,N_19685);
xor U20107 (N_20107,N_19616,N_19503);
nand U20108 (N_20108,N_19766,N_19853);
nor U20109 (N_20109,N_19533,N_19664);
xor U20110 (N_20110,N_19627,N_19758);
nand U20111 (N_20111,N_19700,N_19889);
nor U20112 (N_20112,N_19515,N_19630);
and U20113 (N_20113,N_19764,N_19663);
xnor U20114 (N_20114,N_19565,N_19847);
nand U20115 (N_20115,N_19930,N_19936);
or U20116 (N_20116,N_19914,N_19948);
or U20117 (N_20117,N_19686,N_19902);
nor U20118 (N_20118,N_19818,N_19576);
and U20119 (N_20119,N_19517,N_19976);
and U20120 (N_20120,N_19908,N_19781);
nor U20121 (N_20121,N_19969,N_19581);
and U20122 (N_20122,N_19881,N_19846);
nand U20123 (N_20123,N_19997,N_19647);
and U20124 (N_20124,N_19621,N_19964);
nor U20125 (N_20125,N_19607,N_19755);
xnor U20126 (N_20126,N_19537,N_19981);
and U20127 (N_20127,N_19737,N_19701);
nor U20128 (N_20128,N_19643,N_19695);
nand U20129 (N_20129,N_19609,N_19993);
and U20130 (N_20130,N_19646,N_19932);
or U20131 (N_20131,N_19910,N_19745);
or U20132 (N_20132,N_19659,N_19918);
and U20133 (N_20133,N_19574,N_19951);
and U20134 (N_20134,N_19815,N_19680);
xor U20135 (N_20135,N_19692,N_19790);
xnor U20136 (N_20136,N_19547,N_19705);
xnor U20137 (N_20137,N_19534,N_19567);
or U20138 (N_20138,N_19600,N_19834);
and U20139 (N_20139,N_19862,N_19602);
or U20140 (N_20140,N_19583,N_19763);
xor U20141 (N_20141,N_19883,N_19698);
xnor U20142 (N_20142,N_19983,N_19962);
nor U20143 (N_20143,N_19894,N_19675);
or U20144 (N_20144,N_19971,N_19672);
or U20145 (N_20145,N_19654,N_19612);
xnor U20146 (N_20146,N_19748,N_19589);
xor U20147 (N_20147,N_19714,N_19704);
nand U20148 (N_20148,N_19991,N_19900);
or U20149 (N_20149,N_19827,N_19987);
nand U20150 (N_20150,N_19682,N_19651);
nand U20151 (N_20151,N_19726,N_19554);
nor U20152 (N_20152,N_19662,N_19978);
or U20153 (N_20153,N_19637,N_19795);
and U20154 (N_20154,N_19974,N_19830);
and U20155 (N_20155,N_19566,N_19959);
nor U20156 (N_20156,N_19696,N_19904);
xnor U20157 (N_20157,N_19671,N_19791);
and U20158 (N_20158,N_19939,N_19543);
xnor U20159 (N_20159,N_19587,N_19572);
xnor U20160 (N_20160,N_19541,N_19919);
or U20161 (N_20161,N_19890,N_19571);
or U20162 (N_20162,N_19740,N_19719);
nor U20163 (N_20163,N_19864,N_19760);
nand U20164 (N_20164,N_19523,N_19812);
and U20165 (N_20165,N_19882,N_19563);
xnor U20166 (N_20166,N_19577,N_19739);
nand U20167 (N_20167,N_19788,N_19528);
xor U20168 (N_20168,N_19721,N_19665);
xor U20169 (N_20169,N_19968,N_19832);
nor U20170 (N_20170,N_19810,N_19994);
xor U20171 (N_20171,N_19625,N_19935);
nor U20172 (N_20172,N_19668,N_19539);
nand U20173 (N_20173,N_19877,N_19702);
xor U20174 (N_20174,N_19683,N_19742);
nor U20175 (N_20175,N_19750,N_19958);
nor U20176 (N_20176,N_19934,N_19544);
and U20177 (N_20177,N_19502,N_19899);
and U20178 (N_20178,N_19724,N_19512);
nor U20179 (N_20179,N_19660,N_19869);
and U20180 (N_20180,N_19806,N_19960);
or U20181 (N_20181,N_19973,N_19718);
or U20182 (N_20182,N_19777,N_19596);
nand U20183 (N_20183,N_19744,N_19803);
and U20184 (N_20184,N_19713,N_19673);
nand U20185 (N_20185,N_19928,N_19756);
or U20186 (N_20186,N_19931,N_19774);
nor U20187 (N_20187,N_19863,N_19730);
nor U20188 (N_20188,N_19907,N_19945);
and U20189 (N_20189,N_19678,N_19837);
xnor U20190 (N_20190,N_19759,N_19761);
or U20191 (N_20191,N_19741,N_19800);
and U20192 (N_20192,N_19822,N_19988);
or U20193 (N_20193,N_19892,N_19674);
or U20194 (N_20194,N_19711,N_19542);
xor U20195 (N_20195,N_19938,N_19552);
and U20196 (N_20196,N_19650,N_19749);
or U20197 (N_20197,N_19820,N_19845);
and U20198 (N_20198,N_19545,N_19632);
nand U20199 (N_20199,N_19669,N_19649);
xnor U20200 (N_20200,N_19561,N_19950);
nand U20201 (N_20201,N_19891,N_19592);
and U20202 (N_20202,N_19954,N_19835);
nor U20203 (N_20203,N_19648,N_19568);
nor U20204 (N_20204,N_19855,N_19880);
xor U20205 (N_20205,N_19796,N_19893);
or U20206 (N_20206,N_19856,N_19762);
xnor U20207 (N_20207,N_19848,N_19564);
nand U20208 (N_20208,N_19559,N_19736);
nor U20209 (N_20209,N_19905,N_19952);
or U20210 (N_20210,N_19516,N_19633);
nor U20211 (N_20211,N_19555,N_19757);
xor U20212 (N_20212,N_19508,N_19615);
xor U20213 (N_20213,N_19538,N_19873);
or U20214 (N_20214,N_19579,N_19961);
nor U20215 (N_20215,N_19957,N_19782);
xor U20216 (N_20216,N_19921,N_19575);
nand U20217 (N_20217,N_19801,N_19866);
and U20218 (N_20218,N_19556,N_19729);
and U20219 (N_20219,N_19940,N_19720);
and U20220 (N_20220,N_19926,N_19839);
or U20221 (N_20221,N_19622,N_19652);
or U20222 (N_20222,N_19825,N_19985);
xor U20223 (N_20223,N_19807,N_19775);
and U20224 (N_20224,N_19879,N_19923);
nand U20225 (N_20225,N_19518,N_19884);
nand U20226 (N_20226,N_19507,N_19979);
nor U20227 (N_20227,N_19610,N_19793);
xnor U20228 (N_20228,N_19854,N_19784);
nand U20229 (N_20229,N_19998,N_19992);
or U20230 (N_20230,N_19617,N_19878);
or U20231 (N_20231,N_19619,N_19903);
and U20232 (N_20232,N_19594,N_19821);
or U20233 (N_20233,N_19808,N_19802);
or U20234 (N_20234,N_19562,N_19551);
and U20235 (N_20235,N_19767,N_19792);
nand U20236 (N_20236,N_19529,N_19611);
xnor U20237 (N_20237,N_19970,N_19536);
nor U20238 (N_20238,N_19590,N_19578);
and U20239 (N_20239,N_19972,N_19634);
nand U20240 (N_20240,N_19785,N_19817);
nor U20241 (N_20241,N_19540,N_19814);
or U20242 (N_20242,N_19582,N_19703);
xor U20243 (N_20243,N_19679,N_19509);
nand U20244 (N_20244,N_19688,N_19717);
nor U20245 (N_20245,N_19771,N_19699);
nand U20246 (N_20246,N_19658,N_19804);
xor U20247 (N_20247,N_19557,N_19798);
or U20248 (N_20248,N_19690,N_19986);
or U20249 (N_20249,N_19999,N_19605);
nand U20250 (N_20250,N_19572,N_19594);
nand U20251 (N_20251,N_19740,N_19785);
nand U20252 (N_20252,N_19845,N_19795);
and U20253 (N_20253,N_19733,N_19957);
nor U20254 (N_20254,N_19635,N_19896);
xor U20255 (N_20255,N_19617,N_19721);
nor U20256 (N_20256,N_19634,N_19653);
or U20257 (N_20257,N_19775,N_19544);
or U20258 (N_20258,N_19573,N_19549);
and U20259 (N_20259,N_19688,N_19965);
or U20260 (N_20260,N_19602,N_19841);
or U20261 (N_20261,N_19514,N_19821);
nand U20262 (N_20262,N_19657,N_19784);
and U20263 (N_20263,N_19758,N_19818);
nor U20264 (N_20264,N_19663,N_19807);
or U20265 (N_20265,N_19535,N_19795);
and U20266 (N_20266,N_19766,N_19877);
and U20267 (N_20267,N_19983,N_19709);
or U20268 (N_20268,N_19524,N_19792);
or U20269 (N_20269,N_19699,N_19934);
nand U20270 (N_20270,N_19514,N_19915);
and U20271 (N_20271,N_19501,N_19773);
nand U20272 (N_20272,N_19665,N_19777);
nand U20273 (N_20273,N_19502,N_19690);
xor U20274 (N_20274,N_19745,N_19696);
and U20275 (N_20275,N_19655,N_19960);
nand U20276 (N_20276,N_19611,N_19809);
and U20277 (N_20277,N_19854,N_19890);
and U20278 (N_20278,N_19786,N_19963);
and U20279 (N_20279,N_19919,N_19533);
nor U20280 (N_20280,N_19501,N_19799);
xnor U20281 (N_20281,N_19772,N_19831);
and U20282 (N_20282,N_19954,N_19657);
nand U20283 (N_20283,N_19899,N_19569);
nor U20284 (N_20284,N_19650,N_19647);
nor U20285 (N_20285,N_19804,N_19881);
xnor U20286 (N_20286,N_19773,N_19898);
and U20287 (N_20287,N_19506,N_19689);
xnor U20288 (N_20288,N_19643,N_19778);
or U20289 (N_20289,N_19855,N_19968);
nor U20290 (N_20290,N_19825,N_19629);
or U20291 (N_20291,N_19976,N_19632);
or U20292 (N_20292,N_19635,N_19872);
or U20293 (N_20293,N_19930,N_19622);
xnor U20294 (N_20294,N_19582,N_19822);
xnor U20295 (N_20295,N_19625,N_19981);
nor U20296 (N_20296,N_19938,N_19903);
nand U20297 (N_20297,N_19684,N_19938);
nor U20298 (N_20298,N_19821,N_19542);
xnor U20299 (N_20299,N_19764,N_19670);
or U20300 (N_20300,N_19535,N_19762);
or U20301 (N_20301,N_19548,N_19828);
nor U20302 (N_20302,N_19869,N_19661);
xnor U20303 (N_20303,N_19960,N_19945);
or U20304 (N_20304,N_19595,N_19539);
nand U20305 (N_20305,N_19953,N_19924);
xor U20306 (N_20306,N_19621,N_19957);
nand U20307 (N_20307,N_19784,N_19870);
nor U20308 (N_20308,N_19742,N_19944);
xor U20309 (N_20309,N_19984,N_19862);
nand U20310 (N_20310,N_19625,N_19514);
nand U20311 (N_20311,N_19993,N_19851);
nor U20312 (N_20312,N_19799,N_19659);
nor U20313 (N_20313,N_19719,N_19695);
xnor U20314 (N_20314,N_19636,N_19698);
or U20315 (N_20315,N_19939,N_19652);
nor U20316 (N_20316,N_19871,N_19630);
nor U20317 (N_20317,N_19826,N_19815);
and U20318 (N_20318,N_19810,N_19702);
nor U20319 (N_20319,N_19536,N_19857);
and U20320 (N_20320,N_19750,N_19560);
and U20321 (N_20321,N_19650,N_19788);
or U20322 (N_20322,N_19692,N_19578);
nor U20323 (N_20323,N_19840,N_19841);
nor U20324 (N_20324,N_19935,N_19540);
xnor U20325 (N_20325,N_19702,N_19872);
nor U20326 (N_20326,N_19925,N_19964);
xnor U20327 (N_20327,N_19766,N_19960);
and U20328 (N_20328,N_19842,N_19660);
nor U20329 (N_20329,N_19543,N_19657);
nand U20330 (N_20330,N_19954,N_19785);
and U20331 (N_20331,N_19528,N_19871);
nand U20332 (N_20332,N_19599,N_19630);
xor U20333 (N_20333,N_19719,N_19784);
and U20334 (N_20334,N_19990,N_19943);
nor U20335 (N_20335,N_19803,N_19667);
nor U20336 (N_20336,N_19641,N_19833);
or U20337 (N_20337,N_19517,N_19754);
xnor U20338 (N_20338,N_19862,N_19682);
nand U20339 (N_20339,N_19544,N_19603);
or U20340 (N_20340,N_19733,N_19939);
and U20341 (N_20341,N_19945,N_19981);
nor U20342 (N_20342,N_19937,N_19926);
and U20343 (N_20343,N_19633,N_19875);
and U20344 (N_20344,N_19917,N_19642);
nor U20345 (N_20345,N_19836,N_19597);
nand U20346 (N_20346,N_19919,N_19926);
xnor U20347 (N_20347,N_19653,N_19614);
xor U20348 (N_20348,N_19808,N_19792);
and U20349 (N_20349,N_19680,N_19634);
xor U20350 (N_20350,N_19691,N_19859);
or U20351 (N_20351,N_19671,N_19744);
nand U20352 (N_20352,N_19807,N_19945);
nor U20353 (N_20353,N_19830,N_19549);
nand U20354 (N_20354,N_19710,N_19907);
and U20355 (N_20355,N_19871,N_19615);
nor U20356 (N_20356,N_19919,N_19790);
or U20357 (N_20357,N_19829,N_19732);
xor U20358 (N_20358,N_19662,N_19855);
nor U20359 (N_20359,N_19812,N_19958);
xnor U20360 (N_20360,N_19992,N_19831);
and U20361 (N_20361,N_19709,N_19643);
and U20362 (N_20362,N_19995,N_19899);
nor U20363 (N_20363,N_19571,N_19509);
nand U20364 (N_20364,N_19738,N_19958);
nor U20365 (N_20365,N_19827,N_19715);
nor U20366 (N_20366,N_19650,N_19842);
and U20367 (N_20367,N_19754,N_19674);
nor U20368 (N_20368,N_19860,N_19771);
nand U20369 (N_20369,N_19795,N_19929);
or U20370 (N_20370,N_19566,N_19830);
nor U20371 (N_20371,N_19848,N_19950);
xnor U20372 (N_20372,N_19946,N_19876);
and U20373 (N_20373,N_19745,N_19504);
xor U20374 (N_20374,N_19673,N_19792);
nor U20375 (N_20375,N_19718,N_19931);
nor U20376 (N_20376,N_19882,N_19632);
nor U20377 (N_20377,N_19656,N_19718);
nor U20378 (N_20378,N_19796,N_19769);
and U20379 (N_20379,N_19523,N_19924);
or U20380 (N_20380,N_19834,N_19814);
xor U20381 (N_20381,N_19564,N_19703);
nand U20382 (N_20382,N_19625,N_19649);
or U20383 (N_20383,N_19686,N_19729);
nor U20384 (N_20384,N_19554,N_19919);
nor U20385 (N_20385,N_19820,N_19812);
or U20386 (N_20386,N_19551,N_19682);
xnor U20387 (N_20387,N_19875,N_19846);
nand U20388 (N_20388,N_19752,N_19688);
nand U20389 (N_20389,N_19604,N_19755);
xor U20390 (N_20390,N_19970,N_19679);
xor U20391 (N_20391,N_19598,N_19819);
and U20392 (N_20392,N_19823,N_19634);
xnor U20393 (N_20393,N_19601,N_19875);
xor U20394 (N_20394,N_19745,N_19833);
nand U20395 (N_20395,N_19655,N_19579);
and U20396 (N_20396,N_19956,N_19990);
or U20397 (N_20397,N_19512,N_19545);
or U20398 (N_20398,N_19755,N_19616);
or U20399 (N_20399,N_19780,N_19615);
or U20400 (N_20400,N_19886,N_19563);
and U20401 (N_20401,N_19864,N_19811);
nor U20402 (N_20402,N_19645,N_19812);
and U20403 (N_20403,N_19538,N_19647);
nor U20404 (N_20404,N_19935,N_19819);
or U20405 (N_20405,N_19704,N_19959);
xnor U20406 (N_20406,N_19636,N_19909);
and U20407 (N_20407,N_19613,N_19522);
and U20408 (N_20408,N_19940,N_19910);
nand U20409 (N_20409,N_19980,N_19665);
or U20410 (N_20410,N_19668,N_19910);
or U20411 (N_20411,N_19728,N_19538);
nand U20412 (N_20412,N_19562,N_19543);
nand U20413 (N_20413,N_19801,N_19995);
nand U20414 (N_20414,N_19820,N_19823);
and U20415 (N_20415,N_19697,N_19510);
xnor U20416 (N_20416,N_19889,N_19938);
or U20417 (N_20417,N_19580,N_19801);
or U20418 (N_20418,N_19755,N_19596);
nand U20419 (N_20419,N_19906,N_19771);
xor U20420 (N_20420,N_19515,N_19719);
or U20421 (N_20421,N_19573,N_19545);
or U20422 (N_20422,N_19559,N_19892);
or U20423 (N_20423,N_19581,N_19906);
or U20424 (N_20424,N_19746,N_19829);
and U20425 (N_20425,N_19724,N_19935);
and U20426 (N_20426,N_19670,N_19585);
nor U20427 (N_20427,N_19952,N_19983);
nor U20428 (N_20428,N_19785,N_19894);
xnor U20429 (N_20429,N_19738,N_19579);
xor U20430 (N_20430,N_19519,N_19659);
nand U20431 (N_20431,N_19721,N_19791);
or U20432 (N_20432,N_19618,N_19541);
or U20433 (N_20433,N_19936,N_19635);
and U20434 (N_20434,N_19919,N_19708);
nor U20435 (N_20435,N_19737,N_19772);
nand U20436 (N_20436,N_19812,N_19637);
and U20437 (N_20437,N_19530,N_19701);
nor U20438 (N_20438,N_19750,N_19661);
xor U20439 (N_20439,N_19836,N_19637);
xor U20440 (N_20440,N_19621,N_19694);
nor U20441 (N_20441,N_19931,N_19616);
xnor U20442 (N_20442,N_19508,N_19596);
or U20443 (N_20443,N_19814,N_19767);
nand U20444 (N_20444,N_19920,N_19753);
nand U20445 (N_20445,N_19627,N_19889);
xor U20446 (N_20446,N_19950,N_19719);
nor U20447 (N_20447,N_19608,N_19540);
and U20448 (N_20448,N_19524,N_19595);
or U20449 (N_20449,N_19716,N_19808);
xor U20450 (N_20450,N_19826,N_19915);
nor U20451 (N_20451,N_19755,N_19925);
and U20452 (N_20452,N_19515,N_19816);
xnor U20453 (N_20453,N_19788,N_19665);
nor U20454 (N_20454,N_19998,N_19711);
nor U20455 (N_20455,N_19629,N_19898);
nor U20456 (N_20456,N_19865,N_19515);
or U20457 (N_20457,N_19720,N_19944);
nand U20458 (N_20458,N_19679,N_19830);
or U20459 (N_20459,N_19533,N_19581);
or U20460 (N_20460,N_19686,N_19622);
nor U20461 (N_20461,N_19720,N_19590);
nand U20462 (N_20462,N_19597,N_19563);
or U20463 (N_20463,N_19650,N_19999);
xnor U20464 (N_20464,N_19911,N_19887);
or U20465 (N_20465,N_19863,N_19678);
nor U20466 (N_20466,N_19559,N_19878);
and U20467 (N_20467,N_19794,N_19899);
and U20468 (N_20468,N_19875,N_19885);
or U20469 (N_20469,N_19850,N_19571);
nor U20470 (N_20470,N_19926,N_19502);
xor U20471 (N_20471,N_19855,N_19656);
nand U20472 (N_20472,N_19829,N_19550);
nand U20473 (N_20473,N_19552,N_19831);
and U20474 (N_20474,N_19726,N_19648);
nand U20475 (N_20475,N_19531,N_19547);
xnor U20476 (N_20476,N_19675,N_19723);
nand U20477 (N_20477,N_19955,N_19660);
nand U20478 (N_20478,N_19738,N_19780);
and U20479 (N_20479,N_19569,N_19665);
xnor U20480 (N_20480,N_19953,N_19967);
xor U20481 (N_20481,N_19969,N_19633);
nor U20482 (N_20482,N_19559,N_19796);
nand U20483 (N_20483,N_19926,N_19548);
and U20484 (N_20484,N_19726,N_19519);
nor U20485 (N_20485,N_19731,N_19843);
or U20486 (N_20486,N_19955,N_19707);
nand U20487 (N_20487,N_19702,N_19643);
xor U20488 (N_20488,N_19656,N_19533);
nand U20489 (N_20489,N_19718,N_19744);
and U20490 (N_20490,N_19609,N_19725);
nand U20491 (N_20491,N_19529,N_19628);
nand U20492 (N_20492,N_19718,N_19600);
nor U20493 (N_20493,N_19655,N_19689);
nand U20494 (N_20494,N_19625,N_19809);
and U20495 (N_20495,N_19834,N_19703);
or U20496 (N_20496,N_19604,N_19503);
xor U20497 (N_20497,N_19854,N_19533);
or U20498 (N_20498,N_19880,N_19825);
nand U20499 (N_20499,N_19920,N_19621);
and U20500 (N_20500,N_20455,N_20411);
nand U20501 (N_20501,N_20464,N_20169);
or U20502 (N_20502,N_20232,N_20325);
or U20503 (N_20503,N_20493,N_20272);
nand U20504 (N_20504,N_20171,N_20226);
and U20505 (N_20505,N_20223,N_20075);
and U20506 (N_20506,N_20191,N_20220);
and U20507 (N_20507,N_20076,N_20205);
or U20508 (N_20508,N_20065,N_20119);
or U20509 (N_20509,N_20011,N_20121);
and U20510 (N_20510,N_20380,N_20352);
nor U20511 (N_20511,N_20015,N_20229);
and U20512 (N_20512,N_20402,N_20478);
or U20513 (N_20513,N_20339,N_20370);
nand U20514 (N_20514,N_20388,N_20115);
nand U20515 (N_20515,N_20218,N_20072);
and U20516 (N_20516,N_20060,N_20270);
xnor U20517 (N_20517,N_20194,N_20278);
and U20518 (N_20518,N_20097,N_20179);
nor U20519 (N_20519,N_20190,N_20499);
nor U20520 (N_20520,N_20333,N_20209);
and U20521 (N_20521,N_20048,N_20012);
and U20522 (N_20522,N_20444,N_20373);
or U20523 (N_20523,N_20476,N_20026);
and U20524 (N_20524,N_20160,N_20424);
and U20525 (N_20525,N_20303,N_20112);
nand U20526 (N_20526,N_20035,N_20286);
and U20527 (N_20527,N_20050,N_20042);
or U20528 (N_20528,N_20393,N_20488);
nor U20529 (N_20529,N_20372,N_20255);
nor U20530 (N_20530,N_20474,N_20292);
or U20531 (N_20531,N_20300,N_20203);
or U20532 (N_20532,N_20345,N_20439);
nor U20533 (N_20533,N_20264,N_20240);
and U20534 (N_20534,N_20355,N_20460);
or U20535 (N_20535,N_20058,N_20224);
or U20536 (N_20536,N_20420,N_20214);
or U20537 (N_20537,N_20120,N_20188);
nor U20538 (N_20538,N_20162,N_20418);
and U20539 (N_20539,N_20144,N_20268);
and U20540 (N_20540,N_20117,N_20349);
nand U20541 (N_20541,N_20201,N_20276);
or U20542 (N_20542,N_20416,N_20181);
or U20543 (N_20543,N_20248,N_20311);
or U20544 (N_20544,N_20010,N_20275);
nand U20545 (N_20545,N_20138,N_20423);
nor U20546 (N_20546,N_20344,N_20463);
and U20547 (N_20547,N_20441,N_20004);
xnor U20548 (N_20548,N_20128,N_20412);
and U20549 (N_20549,N_20009,N_20341);
xnor U20550 (N_20550,N_20364,N_20404);
nor U20551 (N_20551,N_20083,N_20314);
and U20552 (N_20552,N_20013,N_20195);
xnor U20553 (N_20553,N_20396,N_20206);
and U20554 (N_20554,N_20100,N_20090);
xor U20555 (N_20555,N_20435,N_20002);
or U20556 (N_20556,N_20134,N_20459);
or U20557 (N_20557,N_20041,N_20158);
xnor U20558 (N_20558,N_20484,N_20461);
xnor U20559 (N_20559,N_20385,N_20225);
nor U20560 (N_20560,N_20148,N_20305);
and U20561 (N_20561,N_20362,N_20453);
nand U20562 (N_20562,N_20197,N_20448);
nor U20563 (N_20563,N_20492,N_20308);
xnor U20564 (N_20564,N_20290,N_20283);
or U20565 (N_20565,N_20284,N_20094);
xor U20566 (N_20566,N_20182,N_20217);
or U20567 (N_20567,N_20122,N_20318);
and U20568 (N_20568,N_20108,N_20295);
nor U20569 (N_20569,N_20323,N_20274);
nor U20570 (N_20570,N_20129,N_20415);
and U20571 (N_20571,N_20399,N_20443);
and U20572 (N_20572,N_20353,N_20447);
nor U20573 (N_20573,N_20340,N_20422);
or U20574 (N_20574,N_20307,N_20174);
or U20575 (N_20575,N_20095,N_20467);
xnor U20576 (N_20576,N_20376,N_20106);
nor U20577 (N_20577,N_20001,N_20277);
nand U20578 (N_20578,N_20334,N_20228);
or U20579 (N_20579,N_20077,N_20235);
nor U20580 (N_20580,N_20375,N_20253);
nand U20581 (N_20581,N_20085,N_20037);
nand U20582 (N_20582,N_20098,N_20452);
nand U20583 (N_20583,N_20212,N_20433);
nand U20584 (N_20584,N_20165,N_20254);
xor U20585 (N_20585,N_20348,N_20329);
nor U20586 (N_20586,N_20031,N_20335);
or U20587 (N_20587,N_20466,N_20167);
or U20588 (N_20588,N_20238,N_20469);
or U20589 (N_20589,N_20070,N_20062);
xnor U20590 (N_20590,N_20316,N_20304);
xnor U20591 (N_20591,N_20326,N_20265);
xor U20592 (N_20592,N_20092,N_20242);
or U20593 (N_20593,N_20025,N_20337);
and U20594 (N_20594,N_20343,N_20354);
xor U20595 (N_20595,N_20193,N_20241);
nor U20596 (N_20596,N_20003,N_20434);
xor U20597 (N_20597,N_20246,N_20266);
nand U20598 (N_20598,N_20321,N_20462);
nand U20599 (N_20599,N_20403,N_20080);
xnor U20600 (N_20600,N_20152,N_20280);
and U20601 (N_20601,N_20103,N_20142);
xnor U20602 (N_20602,N_20027,N_20159);
nor U20603 (N_20603,N_20131,N_20387);
or U20604 (N_20604,N_20495,N_20118);
nand U20605 (N_20605,N_20319,N_20101);
xor U20606 (N_20606,N_20084,N_20456);
nand U20607 (N_20607,N_20306,N_20073);
and U20608 (N_20608,N_20057,N_20397);
or U20609 (N_20609,N_20019,N_20030);
or U20610 (N_20610,N_20279,N_20436);
and U20611 (N_20611,N_20458,N_20136);
and U20612 (N_20612,N_20309,N_20202);
and U20613 (N_20613,N_20081,N_20363);
xnor U20614 (N_20614,N_20389,N_20330);
nand U20615 (N_20615,N_20192,N_20175);
nor U20616 (N_20616,N_20168,N_20043);
xor U20617 (N_20617,N_20033,N_20164);
nand U20618 (N_20618,N_20296,N_20251);
or U20619 (N_20619,N_20130,N_20189);
or U20620 (N_20620,N_20327,N_20360);
or U20621 (N_20621,N_20088,N_20102);
or U20622 (N_20622,N_20281,N_20262);
and U20623 (N_20623,N_20124,N_20170);
nand U20624 (N_20624,N_20064,N_20199);
nor U20625 (N_20625,N_20395,N_20028);
xor U20626 (N_20626,N_20237,N_20239);
and U20627 (N_20627,N_20358,N_20173);
nor U20628 (N_20628,N_20410,N_20384);
nand U20629 (N_20629,N_20252,N_20491);
or U20630 (N_20630,N_20113,N_20213);
or U20631 (N_20631,N_20126,N_20347);
xnor U20632 (N_20632,N_20486,N_20114);
nor U20633 (N_20633,N_20267,N_20079);
or U20634 (N_20634,N_20078,N_20222);
nand U20635 (N_20635,N_20116,N_20074);
xor U20636 (N_20636,N_20089,N_20315);
and U20637 (N_20637,N_20227,N_20000);
nor U20638 (N_20638,N_20157,N_20479);
nand U20639 (N_20639,N_20377,N_20407);
xnor U20640 (N_20640,N_20470,N_20244);
xor U20641 (N_20641,N_20298,N_20398);
xor U20642 (N_20642,N_20297,N_20016);
nor U20643 (N_20643,N_20473,N_20143);
nor U20644 (N_20644,N_20332,N_20245);
or U20645 (N_20645,N_20346,N_20258);
and U20646 (N_20646,N_20086,N_20490);
nor U20647 (N_20647,N_20287,N_20029);
nand U20648 (N_20648,N_20310,N_20155);
nand U20649 (N_20649,N_20123,N_20301);
xor U20650 (N_20650,N_20233,N_20361);
and U20651 (N_20651,N_20430,N_20392);
and U20652 (N_20652,N_20317,N_20082);
nor U20653 (N_20653,N_20405,N_20055);
xor U20654 (N_20654,N_20342,N_20487);
xnor U20655 (N_20655,N_20038,N_20215);
nor U20656 (N_20656,N_20482,N_20256);
nand U20657 (N_20657,N_20145,N_20259);
nand U20658 (N_20658,N_20485,N_20053);
nand U20659 (N_20659,N_20178,N_20451);
xnor U20660 (N_20660,N_20400,N_20440);
or U20661 (N_20661,N_20294,N_20066);
nor U20662 (N_20662,N_20183,N_20198);
xnor U20663 (N_20663,N_20261,N_20040);
xnor U20664 (N_20664,N_20137,N_20285);
nor U20665 (N_20665,N_20250,N_20302);
and U20666 (N_20666,N_20008,N_20204);
or U20667 (N_20667,N_20431,N_20417);
and U20668 (N_20668,N_20437,N_20336);
xor U20669 (N_20669,N_20328,N_20034);
xor U20670 (N_20670,N_20052,N_20269);
nor U20671 (N_20671,N_20185,N_20429);
nand U20672 (N_20672,N_20046,N_20338);
nand U20673 (N_20673,N_20149,N_20263);
nand U20674 (N_20674,N_20379,N_20312);
nand U20675 (N_20675,N_20150,N_20054);
nand U20676 (N_20676,N_20391,N_20104);
or U20677 (N_20677,N_20378,N_20390);
and U20678 (N_20678,N_20005,N_20018);
or U20679 (N_20679,N_20408,N_20442);
nand U20680 (N_20680,N_20401,N_20497);
or U20681 (N_20681,N_20071,N_20371);
xnor U20682 (N_20682,N_20471,N_20051);
and U20683 (N_20683,N_20483,N_20465);
and U20684 (N_20684,N_20282,N_20432);
and U20685 (N_20685,N_20383,N_20350);
or U20686 (N_20686,N_20324,N_20357);
or U20687 (N_20687,N_20409,N_20180);
nand U20688 (N_20688,N_20450,N_20125);
or U20689 (N_20689,N_20386,N_20036);
nor U20690 (N_20690,N_20049,N_20020);
and U20691 (N_20691,N_20427,N_20156);
xor U20692 (N_20692,N_20024,N_20359);
nor U20693 (N_20693,N_20096,N_20059);
nand U20694 (N_20694,N_20367,N_20151);
xor U20695 (N_20695,N_20176,N_20207);
nand U20696 (N_20696,N_20068,N_20454);
or U20697 (N_20697,N_20200,N_20369);
or U20698 (N_20698,N_20127,N_20313);
nand U20699 (N_20699,N_20111,N_20186);
nand U20700 (N_20700,N_20172,N_20381);
nor U20701 (N_20701,N_20091,N_20047);
and U20702 (N_20702,N_20243,N_20247);
or U20703 (N_20703,N_20234,N_20061);
nand U20704 (N_20704,N_20219,N_20039);
or U20705 (N_20705,N_20105,N_20477);
xor U20706 (N_20706,N_20480,N_20069);
xnor U20707 (N_20707,N_20449,N_20067);
or U20708 (N_20708,N_20140,N_20110);
or U20709 (N_20709,N_20299,N_20472);
nor U20710 (N_20710,N_20132,N_20230);
nand U20711 (N_20711,N_20063,N_20022);
nor U20712 (N_20712,N_20221,N_20468);
and U20713 (N_20713,N_20356,N_20146);
and U20714 (N_20714,N_20406,N_20161);
nand U20715 (N_20715,N_20288,N_20216);
xor U20716 (N_20716,N_20093,N_20496);
or U20717 (N_20717,N_20421,N_20257);
nand U20718 (N_20718,N_20006,N_20498);
nand U20719 (N_20719,N_20141,N_20196);
xor U20720 (N_20720,N_20249,N_20322);
nand U20721 (N_20721,N_20394,N_20014);
and U20722 (N_20722,N_20425,N_20419);
and U20723 (N_20723,N_20428,N_20289);
xor U20724 (N_20724,N_20007,N_20438);
xnor U20725 (N_20725,N_20481,N_20445);
or U20726 (N_20726,N_20210,N_20236);
nand U20727 (N_20727,N_20382,N_20293);
or U20728 (N_20728,N_20211,N_20208);
nor U20729 (N_20729,N_20426,N_20446);
nor U20730 (N_20730,N_20260,N_20366);
and U20731 (N_20731,N_20184,N_20135);
nor U20732 (N_20732,N_20291,N_20457);
nand U20733 (N_20733,N_20133,N_20231);
xnor U20734 (N_20734,N_20368,N_20017);
nand U20735 (N_20735,N_20023,N_20166);
nor U20736 (N_20736,N_20087,N_20187);
xnor U20737 (N_20737,N_20045,N_20177);
and U20738 (N_20738,N_20414,N_20273);
and U20739 (N_20739,N_20475,N_20032);
xor U20740 (N_20740,N_20154,N_20494);
and U20741 (N_20741,N_20147,N_20489);
or U20742 (N_20742,N_20044,N_20107);
nor U20743 (N_20743,N_20139,N_20153);
xnor U20744 (N_20744,N_20413,N_20163);
nand U20745 (N_20745,N_20109,N_20021);
or U20746 (N_20746,N_20351,N_20374);
xnor U20747 (N_20747,N_20331,N_20271);
or U20748 (N_20748,N_20320,N_20365);
nor U20749 (N_20749,N_20056,N_20099);
and U20750 (N_20750,N_20087,N_20184);
nand U20751 (N_20751,N_20494,N_20329);
xnor U20752 (N_20752,N_20332,N_20214);
or U20753 (N_20753,N_20486,N_20171);
nor U20754 (N_20754,N_20488,N_20347);
or U20755 (N_20755,N_20490,N_20463);
and U20756 (N_20756,N_20255,N_20180);
or U20757 (N_20757,N_20217,N_20188);
nand U20758 (N_20758,N_20404,N_20094);
and U20759 (N_20759,N_20209,N_20156);
nand U20760 (N_20760,N_20228,N_20076);
nand U20761 (N_20761,N_20133,N_20087);
or U20762 (N_20762,N_20099,N_20302);
nor U20763 (N_20763,N_20373,N_20237);
or U20764 (N_20764,N_20227,N_20033);
nor U20765 (N_20765,N_20281,N_20034);
nor U20766 (N_20766,N_20317,N_20191);
nor U20767 (N_20767,N_20230,N_20229);
and U20768 (N_20768,N_20134,N_20220);
nor U20769 (N_20769,N_20290,N_20061);
nor U20770 (N_20770,N_20242,N_20090);
xnor U20771 (N_20771,N_20102,N_20042);
or U20772 (N_20772,N_20483,N_20347);
or U20773 (N_20773,N_20366,N_20234);
xnor U20774 (N_20774,N_20050,N_20052);
xor U20775 (N_20775,N_20174,N_20202);
and U20776 (N_20776,N_20281,N_20385);
nand U20777 (N_20777,N_20359,N_20044);
and U20778 (N_20778,N_20314,N_20351);
xor U20779 (N_20779,N_20408,N_20269);
nand U20780 (N_20780,N_20391,N_20021);
xor U20781 (N_20781,N_20497,N_20218);
or U20782 (N_20782,N_20339,N_20479);
or U20783 (N_20783,N_20243,N_20167);
nand U20784 (N_20784,N_20400,N_20066);
nor U20785 (N_20785,N_20225,N_20038);
xor U20786 (N_20786,N_20287,N_20355);
nand U20787 (N_20787,N_20397,N_20233);
nand U20788 (N_20788,N_20384,N_20347);
and U20789 (N_20789,N_20246,N_20190);
nand U20790 (N_20790,N_20287,N_20248);
nor U20791 (N_20791,N_20459,N_20009);
and U20792 (N_20792,N_20108,N_20179);
and U20793 (N_20793,N_20282,N_20022);
xor U20794 (N_20794,N_20026,N_20444);
xor U20795 (N_20795,N_20435,N_20267);
nor U20796 (N_20796,N_20060,N_20306);
or U20797 (N_20797,N_20327,N_20449);
nor U20798 (N_20798,N_20427,N_20486);
or U20799 (N_20799,N_20096,N_20357);
xnor U20800 (N_20800,N_20487,N_20148);
and U20801 (N_20801,N_20231,N_20320);
and U20802 (N_20802,N_20462,N_20233);
or U20803 (N_20803,N_20472,N_20125);
nor U20804 (N_20804,N_20361,N_20008);
and U20805 (N_20805,N_20102,N_20456);
nor U20806 (N_20806,N_20206,N_20236);
xor U20807 (N_20807,N_20214,N_20430);
nand U20808 (N_20808,N_20471,N_20043);
and U20809 (N_20809,N_20215,N_20228);
xor U20810 (N_20810,N_20481,N_20050);
nand U20811 (N_20811,N_20340,N_20376);
and U20812 (N_20812,N_20485,N_20100);
nor U20813 (N_20813,N_20426,N_20050);
and U20814 (N_20814,N_20179,N_20383);
nand U20815 (N_20815,N_20457,N_20037);
and U20816 (N_20816,N_20365,N_20142);
nand U20817 (N_20817,N_20439,N_20343);
and U20818 (N_20818,N_20042,N_20255);
nand U20819 (N_20819,N_20261,N_20421);
xor U20820 (N_20820,N_20039,N_20162);
and U20821 (N_20821,N_20164,N_20024);
nor U20822 (N_20822,N_20387,N_20063);
or U20823 (N_20823,N_20293,N_20107);
or U20824 (N_20824,N_20414,N_20250);
and U20825 (N_20825,N_20174,N_20438);
nor U20826 (N_20826,N_20495,N_20254);
nor U20827 (N_20827,N_20016,N_20495);
and U20828 (N_20828,N_20211,N_20483);
nand U20829 (N_20829,N_20206,N_20119);
or U20830 (N_20830,N_20133,N_20363);
or U20831 (N_20831,N_20392,N_20064);
nor U20832 (N_20832,N_20111,N_20458);
nand U20833 (N_20833,N_20209,N_20094);
and U20834 (N_20834,N_20084,N_20125);
xnor U20835 (N_20835,N_20296,N_20452);
xor U20836 (N_20836,N_20067,N_20121);
nor U20837 (N_20837,N_20197,N_20377);
nand U20838 (N_20838,N_20275,N_20466);
and U20839 (N_20839,N_20051,N_20167);
nor U20840 (N_20840,N_20070,N_20007);
nand U20841 (N_20841,N_20107,N_20300);
and U20842 (N_20842,N_20190,N_20389);
xor U20843 (N_20843,N_20176,N_20185);
and U20844 (N_20844,N_20074,N_20345);
nand U20845 (N_20845,N_20301,N_20427);
or U20846 (N_20846,N_20346,N_20126);
nand U20847 (N_20847,N_20030,N_20429);
nand U20848 (N_20848,N_20317,N_20067);
nor U20849 (N_20849,N_20124,N_20279);
and U20850 (N_20850,N_20016,N_20088);
nor U20851 (N_20851,N_20209,N_20426);
xnor U20852 (N_20852,N_20162,N_20022);
xor U20853 (N_20853,N_20397,N_20246);
and U20854 (N_20854,N_20142,N_20220);
nor U20855 (N_20855,N_20092,N_20281);
and U20856 (N_20856,N_20098,N_20277);
or U20857 (N_20857,N_20326,N_20338);
and U20858 (N_20858,N_20263,N_20465);
or U20859 (N_20859,N_20399,N_20372);
or U20860 (N_20860,N_20288,N_20300);
nand U20861 (N_20861,N_20408,N_20390);
nand U20862 (N_20862,N_20235,N_20262);
and U20863 (N_20863,N_20053,N_20360);
and U20864 (N_20864,N_20478,N_20030);
nor U20865 (N_20865,N_20356,N_20161);
xnor U20866 (N_20866,N_20301,N_20085);
nand U20867 (N_20867,N_20322,N_20209);
nand U20868 (N_20868,N_20396,N_20158);
and U20869 (N_20869,N_20457,N_20202);
nand U20870 (N_20870,N_20115,N_20009);
or U20871 (N_20871,N_20224,N_20305);
nand U20872 (N_20872,N_20072,N_20363);
nor U20873 (N_20873,N_20170,N_20225);
xor U20874 (N_20874,N_20257,N_20091);
nor U20875 (N_20875,N_20213,N_20310);
xor U20876 (N_20876,N_20433,N_20326);
nand U20877 (N_20877,N_20256,N_20349);
and U20878 (N_20878,N_20470,N_20115);
nor U20879 (N_20879,N_20420,N_20108);
nor U20880 (N_20880,N_20345,N_20414);
and U20881 (N_20881,N_20327,N_20177);
xnor U20882 (N_20882,N_20203,N_20431);
nor U20883 (N_20883,N_20292,N_20102);
nor U20884 (N_20884,N_20460,N_20044);
nor U20885 (N_20885,N_20126,N_20307);
and U20886 (N_20886,N_20127,N_20282);
or U20887 (N_20887,N_20379,N_20109);
or U20888 (N_20888,N_20486,N_20149);
nand U20889 (N_20889,N_20083,N_20027);
xor U20890 (N_20890,N_20008,N_20053);
nand U20891 (N_20891,N_20011,N_20286);
xnor U20892 (N_20892,N_20407,N_20214);
or U20893 (N_20893,N_20254,N_20012);
xnor U20894 (N_20894,N_20169,N_20077);
nor U20895 (N_20895,N_20190,N_20015);
xnor U20896 (N_20896,N_20442,N_20458);
nand U20897 (N_20897,N_20185,N_20110);
and U20898 (N_20898,N_20492,N_20392);
nand U20899 (N_20899,N_20216,N_20071);
xnor U20900 (N_20900,N_20251,N_20385);
and U20901 (N_20901,N_20382,N_20475);
or U20902 (N_20902,N_20151,N_20232);
and U20903 (N_20903,N_20391,N_20321);
nor U20904 (N_20904,N_20350,N_20332);
nand U20905 (N_20905,N_20065,N_20189);
or U20906 (N_20906,N_20335,N_20360);
and U20907 (N_20907,N_20416,N_20246);
nor U20908 (N_20908,N_20477,N_20229);
nor U20909 (N_20909,N_20020,N_20444);
or U20910 (N_20910,N_20334,N_20296);
xor U20911 (N_20911,N_20033,N_20271);
xor U20912 (N_20912,N_20177,N_20382);
and U20913 (N_20913,N_20207,N_20440);
or U20914 (N_20914,N_20180,N_20319);
or U20915 (N_20915,N_20233,N_20292);
or U20916 (N_20916,N_20041,N_20195);
nor U20917 (N_20917,N_20141,N_20450);
xor U20918 (N_20918,N_20406,N_20053);
or U20919 (N_20919,N_20407,N_20116);
xnor U20920 (N_20920,N_20038,N_20445);
and U20921 (N_20921,N_20370,N_20259);
or U20922 (N_20922,N_20342,N_20448);
xor U20923 (N_20923,N_20046,N_20429);
or U20924 (N_20924,N_20413,N_20230);
or U20925 (N_20925,N_20189,N_20104);
nor U20926 (N_20926,N_20042,N_20048);
or U20927 (N_20927,N_20312,N_20062);
xor U20928 (N_20928,N_20241,N_20199);
or U20929 (N_20929,N_20473,N_20346);
and U20930 (N_20930,N_20273,N_20491);
or U20931 (N_20931,N_20445,N_20415);
nor U20932 (N_20932,N_20033,N_20070);
nand U20933 (N_20933,N_20173,N_20134);
nand U20934 (N_20934,N_20476,N_20037);
and U20935 (N_20935,N_20093,N_20446);
xnor U20936 (N_20936,N_20429,N_20167);
or U20937 (N_20937,N_20256,N_20388);
nand U20938 (N_20938,N_20437,N_20390);
nor U20939 (N_20939,N_20434,N_20338);
nand U20940 (N_20940,N_20484,N_20495);
or U20941 (N_20941,N_20169,N_20246);
nand U20942 (N_20942,N_20097,N_20379);
nor U20943 (N_20943,N_20199,N_20155);
and U20944 (N_20944,N_20088,N_20154);
or U20945 (N_20945,N_20406,N_20254);
and U20946 (N_20946,N_20135,N_20141);
and U20947 (N_20947,N_20404,N_20300);
nand U20948 (N_20948,N_20353,N_20060);
xor U20949 (N_20949,N_20111,N_20215);
and U20950 (N_20950,N_20262,N_20218);
or U20951 (N_20951,N_20271,N_20233);
nor U20952 (N_20952,N_20498,N_20189);
and U20953 (N_20953,N_20061,N_20362);
and U20954 (N_20954,N_20343,N_20328);
xnor U20955 (N_20955,N_20110,N_20143);
xor U20956 (N_20956,N_20207,N_20276);
nand U20957 (N_20957,N_20027,N_20144);
and U20958 (N_20958,N_20139,N_20369);
xnor U20959 (N_20959,N_20082,N_20311);
or U20960 (N_20960,N_20134,N_20161);
xnor U20961 (N_20961,N_20278,N_20143);
nor U20962 (N_20962,N_20274,N_20040);
nand U20963 (N_20963,N_20020,N_20247);
nand U20964 (N_20964,N_20484,N_20401);
nor U20965 (N_20965,N_20404,N_20135);
and U20966 (N_20966,N_20498,N_20364);
or U20967 (N_20967,N_20037,N_20211);
nor U20968 (N_20968,N_20038,N_20383);
or U20969 (N_20969,N_20494,N_20043);
xor U20970 (N_20970,N_20270,N_20391);
xnor U20971 (N_20971,N_20249,N_20026);
and U20972 (N_20972,N_20106,N_20095);
nand U20973 (N_20973,N_20047,N_20045);
or U20974 (N_20974,N_20419,N_20284);
nor U20975 (N_20975,N_20440,N_20295);
nor U20976 (N_20976,N_20433,N_20183);
or U20977 (N_20977,N_20270,N_20058);
nor U20978 (N_20978,N_20121,N_20117);
xnor U20979 (N_20979,N_20321,N_20336);
nor U20980 (N_20980,N_20051,N_20092);
xor U20981 (N_20981,N_20333,N_20102);
xor U20982 (N_20982,N_20040,N_20038);
nand U20983 (N_20983,N_20153,N_20469);
xnor U20984 (N_20984,N_20329,N_20008);
or U20985 (N_20985,N_20063,N_20241);
xor U20986 (N_20986,N_20029,N_20051);
xnor U20987 (N_20987,N_20348,N_20283);
or U20988 (N_20988,N_20018,N_20269);
and U20989 (N_20989,N_20435,N_20425);
or U20990 (N_20990,N_20423,N_20079);
or U20991 (N_20991,N_20069,N_20101);
nor U20992 (N_20992,N_20178,N_20296);
xnor U20993 (N_20993,N_20426,N_20009);
nor U20994 (N_20994,N_20092,N_20083);
xnor U20995 (N_20995,N_20042,N_20029);
xnor U20996 (N_20996,N_20080,N_20431);
xnor U20997 (N_20997,N_20426,N_20465);
nor U20998 (N_20998,N_20126,N_20264);
xnor U20999 (N_20999,N_20226,N_20394);
nand U21000 (N_21000,N_20624,N_20748);
and U21001 (N_21001,N_20711,N_20617);
nand U21002 (N_21002,N_20915,N_20811);
xor U21003 (N_21003,N_20528,N_20782);
xnor U21004 (N_21004,N_20610,N_20847);
nand U21005 (N_21005,N_20836,N_20804);
or U21006 (N_21006,N_20575,N_20983);
nor U21007 (N_21007,N_20840,N_20523);
and U21008 (N_21008,N_20879,N_20877);
nor U21009 (N_21009,N_20548,N_20839);
or U21010 (N_21010,N_20921,N_20855);
or U21011 (N_21011,N_20513,N_20612);
nand U21012 (N_21012,N_20936,N_20912);
xor U21013 (N_21013,N_20502,N_20919);
nand U21014 (N_21014,N_20850,N_20928);
nand U21015 (N_21015,N_20571,N_20860);
xnor U21016 (N_21016,N_20686,N_20690);
xor U21017 (N_21017,N_20941,N_20520);
and U21018 (N_21018,N_20957,N_20680);
and U21019 (N_21019,N_20542,N_20543);
nand U21020 (N_21020,N_20696,N_20723);
xnor U21021 (N_21021,N_20628,N_20675);
nand U21022 (N_21022,N_20508,N_20933);
nor U21023 (N_21023,N_20909,N_20634);
and U21024 (N_21024,N_20753,N_20925);
xor U21025 (N_21025,N_20578,N_20638);
xor U21026 (N_21026,N_20793,N_20526);
xnor U21027 (N_21027,N_20947,N_20780);
or U21028 (N_21028,N_20777,N_20990);
or U21029 (N_21029,N_20946,N_20545);
and U21030 (N_21030,N_20630,N_20791);
xor U21031 (N_21031,N_20958,N_20721);
and U21032 (N_21032,N_20601,N_20832);
and U21033 (N_21033,N_20885,N_20707);
nand U21034 (N_21034,N_20734,N_20755);
and U21035 (N_21035,N_20962,N_20917);
nand U21036 (N_21036,N_20593,N_20954);
nor U21037 (N_21037,N_20812,N_20798);
nand U21038 (N_21038,N_20834,N_20605);
xor U21039 (N_21039,N_20911,N_20521);
xor U21040 (N_21040,N_20944,N_20703);
or U21041 (N_21041,N_20854,N_20988);
xnor U21042 (N_21042,N_20599,N_20658);
or U21043 (N_21043,N_20895,N_20500);
nand U21044 (N_21044,N_20640,N_20616);
nor U21045 (N_21045,N_20910,N_20637);
xnor U21046 (N_21046,N_20923,N_20740);
or U21047 (N_21047,N_20705,N_20861);
nor U21048 (N_21048,N_20982,N_20905);
and U21049 (N_21049,N_20689,N_20600);
or U21050 (N_21050,N_20532,N_20701);
xor U21051 (N_21051,N_20639,N_20514);
xor U21052 (N_21052,N_20670,N_20559);
nor U21053 (N_21053,N_20567,N_20677);
xnor U21054 (N_21054,N_20953,N_20626);
nand U21055 (N_21055,N_20949,N_20709);
nor U21056 (N_21056,N_20841,N_20980);
xor U21057 (N_21057,N_20975,N_20906);
and U21058 (N_21058,N_20706,N_20880);
nor U21059 (N_21059,N_20851,N_20713);
nor U21060 (N_21060,N_20817,N_20746);
or U21061 (N_21061,N_20903,N_20785);
nor U21062 (N_21062,N_20747,N_20971);
xnor U21063 (N_21063,N_20504,N_20752);
nand U21064 (N_21064,N_20918,N_20563);
or U21065 (N_21065,N_20862,N_20550);
or U21066 (N_21066,N_20636,N_20995);
xnor U21067 (N_21067,N_20655,N_20955);
xnor U21068 (N_21068,N_20683,N_20932);
and U21069 (N_21069,N_20889,N_20856);
nand U21070 (N_21070,N_20989,N_20687);
nand U21071 (N_21071,N_20647,N_20725);
nand U21072 (N_21072,N_20552,N_20887);
xor U21073 (N_21073,N_20778,N_20758);
xnor U21074 (N_21074,N_20622,N_20580);
nor U21075 (N_21075,N_20822,N_20669);
nand U21076 (N_21076,N_20651,N_20769);
or U21077 (N_21077,N_20700,N_20979);
or U21078 (N_21078,N_20838,N_20896);
nand U21079 (N_21079,N_20695,N_20770);
and U21080 (N_21080,N_20524,N_20809);
xor U21081 (N_21081,N_20566,N_20779);
nor U21082 (N_21082,N_20792,N_20914);
nand U21083 (N_21083,N_20754,N_20898);
and U21084 (N_21084,N_20576,N_20541);
and U21085 (N_21085,N_20611,N_20835);
xor U21086 (N_21086,N_20731,N_20924);
and U21087 (N_21087,N_20901,N_20930);
nand U21088 (N_21088,N_20570,N_20787);
nor U21089 (N_21089,N_20773,N_20897);
xor U21090 (N_21090,N_20682,N_20509);
nor U21091 (N_21091,N_20872,N_20875);
or U21092 (N_21092,N_20587,N_20907);
and U21093 (N_21093,N_20582,N_20594);
and U21094 (N_21094,N_20842,N_20558);
or U21095 (N_21095,N_20503,N_20865);
and U21096 (N_21096,N_20603,N_20867);
or U21097 (N_21097,N_20814,N_20950);
and U21098 (N_21098,N_20660,N_20678);
nor U21099 (N_21099,N_20940,N_20920);
or U21100 (N_21100,N_20987,N_20871);
and U21101 (N_21101,N_20583,N_20556);
or U21102 (N_21102,N_20813,N_20531);
and U21103 (N_21103,N_20938,N_20884);
and U21104 (N_21104,N_20863,N_20715);
or U21105 (N_21105,N_20935,N_20961);
nor U21106 (N_21106,N_20676,N_20684);
and U21107 (N_21107,N_20697,N_20800);
or U21108 (N_21108,N_20790,N_20592);
or U21109 (N_21109,N_20573,N_20968);
nor U21110 (N_21110,N_20641,N_20536);
xor U21111 (N_21111,N_20878,N_20537);
nand U21112 (N_21112,N_20623,N_20653);
or U21113 (N_21113,N_20751,N_20663);
and U21114 (N_21114,N_20665,N_20621);
xnor U21115 (N_21115,N_20619,N_20607);
nand U21116 (N_21116,N_20631,N_20560);
nand U21117 (N_21117,N_20688,N_20507);
and U21118 (N_21118,N_20998,N_20891);
xnor U21119 (N_21119,N_20674,N_20627);
nand U21120 (N_21120,N_20673,N_20849);
nor U21121 (N_21121,N_20985,N_20538);
nand U21122 (N_21122,N_20976,N_20994);
nand U21123 (N_21123,N_20650,N_20816);
nand U21124 (N_21124,N_20931,N_20744);
xor U21125 (N_21125,N_20551,N_20679);
and U21126 (N_21126,N_20539,N_20899);
nand U21127 (N_21127,N_20590,N_20781);
and U21128 (N_21128,N_20760,N_20997);
and U21129 (N_21129,N_20876,N_20529);
xor U21130 (N_21130,N_20963,N_20694);
or U21131 (N_21131,N_20894,N_20717);
nand U21132 (N_21132,N_20945,N_20757);
nand U21133 (N_21133,N_20595,N_20766);
nand U21134 (N_21134,N_20741,N_20805);
nor U21135 (N_21135,N_20726,N_20737);
and U21136 (N_21136,N_20719,N_20765);
nor U21137 (N_21137,N_20803,N_20750);
or U21138 (N_21138,N_20667,N_20685);
nand U21139 (N_21139,N_20827,N_20828);
xor U21140 (N_21140,N_20977,N_20892);
nor U21141 (N_21141,N_20718,N_20959);
xor U21142 (N_21142,N_20549,N_20972);
and U21143 (N_21143,N_20943,N_20618);
or U21144 (N_21144,N_20661,N_20649);
nand U21145 (N_21145,N_20739,N_20795);
and U21146 (N_21146,N_20716,N_20738);
xnor U21147 (N_21147,N_20632,N_20714);
nor U21148 (N_21148,N_20749,N_20656);
nand U21149 (N_21149,N_20613,N_20984);
nor U21150 (N_21150,N_20608,N_20562);
or U21151 (N_21151,N_20642,N_20824);
nor U21152 (N_21152,N_20808,N_20633);
nand U21153 (N_21153,N_20857,N_20648);
or U21154 (N_21154,N_20659,N_20643);
nand U21155 (N_21155,N_20698,N_20646);
nor U21156 (N_21156,N_20645,N_20888);
nand U21157 (N_21157,N_20807,N_20515);
nor U21158 (N_21158,N_20829,N_20761);
nor U21159 (N_21159,N_20598,N_20967);
or U21160 (N_21160,N_20708,N_20966);
xnor U21161 (N_21161,N_20729,N_20519);
xor U21162 (N_21162,N_20710,N_20743);
xor U21163 (N_21163,N_20527,N_20873);
nor U21164 (N_21164,N_20693,N_20819);
nand U21165 (N_21165,N_20820,N_20704);
nor U21166 (N_21166,N_20886,N_20801);
xnor U21167 (N_21167,N_20702,N_20506);
nand U21168 (N_21168,N_20555,N_20732);
and U21169 (N_21169,N_20794,N_20952);
nand U21170 (N_21170,N_20728,N_20581);
xor U21171 (N_21171,N_20881,N_20799);
or U21172 (N_21172,N_20596,N_20991);
nor U21173 (N_21173,N_20522,N_20553);
and U21174 (N_21174,N_20783,N_20916);
nor U21175 (N_21175,N_20908,N_20831);
nor U21176 (N_21176,N_20974,N_20591);
nor U21177 (N_21177,N_20561,N_20845);
nor U21178 (N_21178,N_20870,N_20826);
xnor U21179 (N_21179,N_20858,N_20774);
nand U21180 (N_21180,N_20934,N_20992);
xor U21181 (N_21181,N_20501,N_20929);
xor U21182 (N_21182,N_20604,N_20652);
or U21183 (N_21183,N_20797,N_20525);
and U21184 (N_21184,N_20733,N_20775);
xnor U21185 (N_21185,N_20668,N_20505);
xor U21186 (N_21186,N_20986,N_20964);
and U21187 (N_21187,N_20544,N_20602);
and U21188 (N_21188,N_20554,N_20745);
nand U21189 (N_21189,N_20666,N_20564);
and U21190 (N_21190,N_20771,N_20534);
nand U21191 (N_21191,N_20588,N_20759);
xnor U21192 (N_21192,N_20927,N_20846);
nor U21193 (N_21193,N_20939,N_20736);
nand U21194 (N_21194,N_20902,N_20609);
and U21195 (N_21195,N_20510,N_20823);
nor U21196 (N_21196,N_20951,N_20833);
nand U21197 (N_21197,N_20913,N_20904);
and U21198 (N_21198,N_20776,N_20970);
nor U21199 (N_21199,N_20796,N_20993);
xnor U21200 (N_21200,N_20784,N_20893);
nand U21201 (N_21201,N_20786,N_20772);
nand U21202 (N_21202,N_20981,N_20657);
nor U21203 (N_21203,N_20672,N_20868);
nand U21204 (N_21204,N_20965,N_20585);
nor U21205 (N_21205,N_20830,N_20629);
nand U21206 (N_21206,N_20712,N_20722);
xnor U21207 (N_21207,N_20844,N_20724);
and U21208 (N_21208,N_20699,N_20568);
xnor U21209 (N_21209,N_20586,N_20691);
nand U21210 (N_21210,N_20763,N_20517);
or U21211 (N_21211,N_20843,N_20756);
nand U21212 (N_21212,N_20900,N_20978);
nand U21213 (N_21213,N_20615,N_20546);
and U21214 (N_21214,N_20735,N_20620);
nor U21215 (N_21215,N_20569,N_20720);
nor U21216 (N_21216,N_20671,N_20727);
nor U21217 (N_21217,N_20540,N_20853);
and U21218 (N_21218,N_20789,N_20584);
or U21219 (N_21219,N_20654,N_20557);
nand U21220 (N_21220,N_20874,N_20511);
or U21221 (N_21221,N_20730,N_20764);
or U21222 (N_21222,N_20664,N_20681);
and U21223 (N_21223,N_20960,N_20815);
nor U21224 (N_21224,N_20530,N_20942);
nor U21225 (N_21225,N_20973,N_20890);
nor U21226 (N_21226,N_20635,N_20589);
or U21227 (N_21227,N_20883,N_20577);
nor U21228 (N_21228,N_20518,N_20866);
xor U21229 (N_21229,N_20996,N_20597);
or U21230 (N_21230,N_20574,N_20512);
and U21231 (N_21231,N_20692,N_20864);
xor U21232 (N_21232,N_20606,N_20802);
nor U21233 (N_21233,N_20937,N_20882);
nor U21234 (N_21234,N_20625,N_20810);
nor U21235 (N_21235,N_20948,N_20644);
xor U21236 (N_21236,N_20533,N_20579);
xor U21237 (N_21237,N_20922,N_20572);
and U21238 (N_21238,N_20837,N_20535);
and U21239 (N_21239,N_20788,N_20547);
nand U21240 (N_21240,N_20565,N_20859);
or U21241 (N_21241,N_20516,N_20999);
nand U21242 (N_21242,N_20614,N_20825);
or U21243 (N_21243,N_20926,N_20821);
and U21244 (N_21244,N_20852,N_20762);
nor U21245 (N_21245,N_20848,N_20818);
nor U21246 (N_21246,N_20956,N_20767);
xnor U21247 (N_21247,N_20742,N_20869);
nor U21248 (N_21248,N_20806,N_20969);
nor U21249 (N_21249,N_20662,N_20768);
nand U21250 (N_21250,N_20675,N_20830);
nor U21251 (N_21251,N_20575,N_20899);
nor U21252 (N_21252,N_20998,N_20682);
or U21253 (N_21253,N_20694,N_20511);
nor U21254 (N_21254,N_20755,N_20544);
and U21255 (N_21255,N_20960,N_20800);
nand U21256 (N_21256,N_20884,N_20894);
nand U21257 (N_21257,N_20967,N_20512);
or U21258 (N_21258,N_20905,N_20544);
or U21259 (N_21259,N_20644,N_20993);
xnor U21260 (N_21260,N_20539,N_20902);
xnor U21261 (N_21261,N_20622,N_20800);
or U21262 (N_21262,N_20555,N_20553);
and U21263 (N_21263,N_20900,N_20704);
nand U21264 (N_21264,N_20942,N_20893);
or U21265 (N_21265,N_20811,N_20565);
nand U21266 (N_21266,N_20651,N_20692);
xnor U21267 (N_21267,N_20600,N_20816);
and U21268 (N_21268,N_20904,N_20737);
xor U21269 (N_21269,N_20599,N_20529);
nand U21270 (N_21270,N_20964,N_20705);
and U21271 (N_21271,N_20760,N_20969);
nand U21272 (N_21272,N_20859,N_20773);
nor U21273 (N_21273,N_20567,N_20997);
or U21274 (N_21274,N_20736,N_20644);
or U21275 (N_21275,N_20676,N_20984);
nor U21276 (N_21276,N_20624,N_20773);
nor U21277 (N_21277,N_20991,N_20750);
xnor U21278 (N_21278,N_20591,N_20920);
nor U21279 (N_21279,N_20833,N_20502);
xnor U21280 (N_21280,N_20684,N_20833);
nand U21281 (N_21281,N_20630,N_20599);
xnor U21282 (N_21282,N_20762,N_20804);
and U21283 (N_21283,N_20812,N_20915);
nand U21284 (N_21284,N_20818,N_20924);
xor U21285 (N_21285,N_20638,N_20747);
nand U21286 (N_21286,N_20513,N_20759);
nand U21287 (N_21287,N_20751,N_20818);
nand U21288 (N_21288,N_20668,N_20867);
or U21289 (N_21289,N_20856,N_20873);
xnor U21290 (N_21290,N_20888,N_20515);
xor U21291 (N_21291,N_20713,N_20709);
and U21292 (N_21292,N_20533,N_20770);
xor U21293 (N_21293,N_20630,N_20844);
nand U21294 (N_21294,N_20688,N_20842);
nand U21295 (N_21295,N_20905,N_20960);
or U21296 (N_21296,N_20884,N_20599);
nor U21297 (N_21297,N_20663,N_20917);
nand U21298 (N_21298,N_20920,N_20533);
or U21299 (N_21299,N_20745,N_20970);
or U21300 (N_21300,N_20978,N_20972);
and U21301 (N_21301,N_20711,N_20552);
nor U21302 (N_21302,N_20831,N_20521);
or U21303 (N_21303,N_20647,N_20549);
and U21304 (N_21304,N_20966,N_20519);
and U21305 (N_21305,N_20610,N_20579);
xor U21306 (N_21306,N_20908,N_20741);
and U21307 (N_21307,N_20684,N_20540);
or U21308 (N_21308,N_20801,N_20881);
and U21309 (N_21309,N_20783,N_20769);
and U21310 (N_21310,N_20877,N_20825);
nor U21311 (N_21311,N_20553,N_20669);
nor U21312 (N_21312,N_20959,N_20542);
xor U21313 (N_21313,N_20714,N_20643);
xnor U21314 (N_21314,N_20541,N_20994);
or U21315 (N_21315,N_20616,N_20807);
nor U21316 (N_21316,N_20726,N_20504);
nor U21317 (N_21317,N_20967,N_20618);
xor U21318 (N_21318,N_20523,N_20785);
xor U21319 (N_21319,N_20583,N_20893);
and U21320 (N_21320,N_20810,N_20997);
xnor U21321 (N_21321,N_20754,N_20504);
nand U21322 (N_21322,N_20792,N_20622);
nand U21323 (N_21323,N_20813,N_20826);
and U21324 (N_21324,N_20573,N_20606);
nand U21325 (N_21325,N_20977,N_20747);
or U21326 (N_21326,N_20706,N_20946);
nand U21327 (N_21327,N_20557,N_20780);
xnor U21328 (N_21328,N_20916,N_20740);
and U21329 (N_21329,N_20693,N_20663);
nor U21330 (N_21330,N_20776,N_20660);
or U21331 (N_21331,N_20588,N_20541);
nor U21332 (N_21332,N_20981,N_20601);
xnor U21333 (N_21333,N_20876,N_20574);
nand U21334 (N_21334,N_20854,N_20616);
xor U21335 (N_21335,N_20742,N_20660);
or U21336 (N_21336,N_20520,N_20810);
xor U21337 (N_21337,N_20890,N_20936);
and U21338 (N_21338,N_20922,N_20784);
nand U21339 (N_21339,N_20707,N_20735);
or U21340 (N_21340,N_20574,N_20898);
or U21341 (N_21341,N_20642,N_20887);
nor U21342 (N_21342,N_20820,N_20725);
nand U21343 (N_21343,N_20792,N_20911);
nand U21344 (N_21344,N_20966,N_20504);
or U21345 (N_21345,N_20733,N_20957);
nand U21346 (N_21346,N_20653,N_20649);
nand U21347 (N_21347,N_20657,N_20613);
or U21348 (N_21348,N_20987,N_20941);
or U21349 (N_21349,N_20755,N_20866);
xor U21350 (N_21350,N_20520,N_20689);
xnor U21351 (N_21351,N_20777,N_20866);
nand U21352 (N_21352,N_20672,N_20567);
and U21353 (N_21353,N_20789,N_20979);
nor U21354 (N_21354,N_20629,N_20551);
nand U21355 (N_21355,N_20754,N_20900);
nor U21356 (N_21356,N_20751,N_20836);
nor U21357 (N_21357,N_20546,N_20716);
xor U21358 (N_21358,N_20976,N_20692);
xnor U21359 (N_21359,N_20752,N_20723);
or U21360 (N_21360,N_20504,N_20876);
or U21361 (N_21361,N_20713,N_20965);
nor U21362 (N_21362,N_20554,N_20948);
nand U21363 (N_21363,N_20967,N_20852);
xnor U21364 (N_21364,N_20694,N_20803);
and U21365 (N_21365,N_20660,N_20803);
xnor U21366 (N_21366,N_20920,N_20805);
nor U21367 (N_21367,N_20547,N_20606);
or U21368 (N_21368,N_20761,N_20658);
xor U21369 (N_21369,N_20511,N_20684);
or U21370 (N_21370,N_20871,N_20612);
and U21371 (N_21371,N_20700,N_20689);
nor U21372 (N_21372,N_20717,N_20842);
nor U21373 (N_21373,N_20642,N_20898);
xor U21374 (N_21374,N_20680,N_20993);
or U21375 (N_21375,N_20853,N_20579);
or U21376 (N_21376,N_20653,N_20561);
nand U21377 (N_21377,N_20675,N_20646);
and U21378 (N_21378,N_20591,N_20592);
and U21379 (N_21379,N_20507,N_20773);
nand U21380 (N_21380,N_20920,N_20701);
nor U21381 (N_21381,N_20820,N_20844);
xor U21382 (N_21382,N_20966,N_20798);
or U21383 (N_21383,N_20609,N_20666);
or U21384 (N_21384,N_20829,N_20980);
and U21385 (N_21385,N_20846,N_20612);
nor U21386 (N_21386,N_20540,N_20850);
or U21387 (N_21387,N_20898,N_20691);
xnor U21388 (N_21388,N_20634,N_20539);
or U21389 (N_21389,N_20951,N_20796);
nand U21390 (N_21390,N_20639,N_20735);
xor U21391 (N_21391,N_20747,N_20660);
and U21392 (N_21392,N_20839,N_20740);
or U21393 (N_21393,N_20533,N_20729);
nor U21394 (N_21394,N_20740,N_20618);
and U21395 (N_21395,N_20689,N_20769);
and U21396 (N_21396,N_20643,N_20518);
and U21397 (N_21397,N_20569,N_20551);
xnor U21398 (N_21398,N_20964,N_20520);
or U21399 (N_21399,N_20679,N_20751);
xor U21400 (N_21400,N_20797,N_20883);
or U21401 (N_21401,N_20737,N_20888);
and U21402 (N_21402,N_20976,N_20933);
and U21403 (N_21403,N_20731,N_20859);
nand U21404 (N_21404,N_20709,N_20967);
nor U21405 (N_21405,N_20610,N_20510);
xnor U21406 (N_21406,N_20725,N_20657);
and U21407 (N_21407,N_20884,N_20640);
and U21408 (N_21408,N_20522,N_20767);
or U21409 (N_21409,N_20662,N_20577);
and U21410 (N_21410,N_20868,N_20843);
nand U21411 (N_21411,N_20611,N_20519);
and U21412 (N_21412,N_20687,N_20586);
xnor U21413 (N_21413,N_20980,N_20552);
nand U21414 (N_21414,N_20835,N_20585);
or U21415 (N_21415,N_20614,N_20683);
or U21416 (N_21416,N_20833,N_20660);
nor U21417 (N_21417,N_20695,N_20671);
and U21418 (N_21418,N_20877,N_20626);
and U21419 (N_21419,N_20921,N_20664);
nand U21420 (N_21420,N_20602,N_20854);
nor U21421 (N_21421,N_20811,N_20815);
nor U21422 (N_21422,N_20580,N_20949);
xor U21423 (N_21423,N_20755,N_20878);
or U21424 (N_21424,N_20926,N_20886);
and U21425 (N_21425,N_20631,N_20725);
nor U21426 (N_21426,N_20688,N_20869);
nand U21427 (N_21427,N_20767,N_20578);
or U21428 (N_21428,N_20704,N_20793);
nand U21429 (N_21429,N_20859,N_20583);
nor U21430 (N_21430,N_20878,N_20553);
or U21431 (N_21431,N_20753,N_20920);
or U21432 (N_21432,N_20513,N_20926);
nand U21433 (N_21433,N_20949,N_20870);
nand U21434 (N_21434,N_20788,N_20612);
or U21435 (N_21435,N_20950,N_20764);
or U21436 (N_21436,N_20946,N_20641);
xnor U21437 (N_21437,N_20861,N_20598);
and U21438 (N_21438,N_20906,N_20876);
nor U21439 (N_21439,N_20718,N_20919);
nand U21440 (N_21440,N_20811,N_20766);
xnor U21441 (N_21441,N_20745,N_20522);
and U21442 (N_21442,N_20785,N_20759);
nor U21443 (N_21443,N_20867,N_20576);
xor U21444 (N_21444,N_20598,N_20756);
nand U21445 (N_21445,N_20796,N_20660);
or U21446 (N_21446,N_20643,N_20969);
or U21447 (N_21447,N_20819,N_20995);
or U21448 (N_21448,N_20788,N_20620);
xor U21449 (N_21449,N_20881,N_20673);
xor U21450 (N_21450,N_20823,N_20679);
nor U21451 (N_21451,N_20929,N_20927);
nand U21452 (N_21452,N_20601,N_20594);
nor U21453 (N_21453,N_20685,N_20893);
xnor U21454 (N_21454,N_20524,N_20637);
nand U21455 (N_21455,N_20705,N_20769);
nor U21456 (N_21456,N_20636,N_20545);
and U21457 (N_21457,N_20857,N_20533);
nor U21458 (N_21458,N_20948,N_20684);
nand U21459 (N_21459,N_20764,N_20974);
xnor U21460 (N_21460,N_20809,N_20534);
or U21461 (N_21461,N_20764,N_20843);
xor U21462 (N_21462,N_20725,N_20979);
xor U21463 (N_21463,N_20760,N_20998);
nand U21464 (N_21464,N_20775,N_20633);
or U21465 (N_21465,N_20844,N_20727);
nand U21466 (N_21466,N_20596,N_20741);
and U21467 (N_21467,N_20952,N_20884);
xnor U21468 (N_21468,N_20592,N_20942);
xnor U21469 (N_21469,N_20628,N_20733);
and U21470 (N_21470,N_20797,N_20798);
and U21471 (N_21471,N_20872,N_20641);
or U21472 (N_21472,N_20869,N_20781);
nor U21473 (N_21473,N_20861,N_20756);
and U21474 (N_21474,N_20518,N_20604);
nand U21475 (N_21475,N_20753,N_20591);
xor U21476 (N_21476,N_20898,N_20906);
nand U21477 (N_21477,N_20774,N_20825);
xnor U21478 (N_21478,N_20845,N_20859);
nor U21479 (N_21479,N_20954,N_20909);
or U21480 (N_21480,N_20626,N_20593);
or U21481 (N_21481,N_20625,N_20883);
nand U21482 (N_21482,N_20533,N_20986);
xnor U21483 (N_21483,N_20726,N_20688);
or U21484 (N_21484,N_20812,N_20916);
xnor U21485 (N_21485,N_20775,N_20585);
nand U21486 (N_21486,N_20661,N_20969);
nor U21487 (N_21487,N_20848,N_20916);
and U21488 (N_21488,N_20999,N_20644);
nand U21489 (N_21489,N_20500,N_20803);
xor U21490 (N_21490,N_20937,N_20513);
and U21491 (N_21491,N_20980,N_20669);
and U21492 (N_21492,N_20580,N_20708);
or U21493 (N_21493,N_20952,N_20700);
and U21494 (N_21494,N_20591,N_20628);
nand U21495 (N_21495,N_20923,N_20982);
xnor U21496 (N_21496,N_20533,N_20693);
nand U21497 (N_21497,N_20956,N_20868);
nor U21498 (N_21498,N_20835,N_20656);
or U21499 (N_21499,N_20575,N_20813);
nand U21500 (N_21500,N_21443,N_21289);
or U21501 (N_21501,N_21403,N_21001);
and U21502 (N_21502,N_21149,N_21376);
nor U21503 (N_21503,N_21236,N_21250);
or U21504 (N_21504,N_21315,N_21094);
xor U21505 (N_21505,N_21468,N_21395);
nand U21506 (N_21506,N_21169,N_21168);
or U21507 (N_21507,N_21055,N_21155);
nand U21508 (N_21508,N_21404,N_21392);
or U21509 (N_21509,N_21400,N_21491);
or U21510 (N_21510,N_21344,N_21386);
or U21511 (N_21511,N_21434,N_21273);
or U21512 (N_21512,N_21073,N_21298);
xor U21513 (N_21513,N_21226,N_21045);
and U21514 (N_21514,N_21077,N_21488);
or U21515 (N_21515,N_21104,N_21293);
xnor U21516 (N_21516,N_21388,N_21409);
or U21517 (N_21517,N_21249,N_21260);
xnor U21518 (N_21518,N_21188,N_21397);
xnor U21519 (N_21519,N_21133,N_21474);
and U21520 (N_21520,N_21145,N_21438);
nor U21521 (N_21521,N_21335,N_21261);
nor U21522 (N_21522,N_21117,N_21020);
nand U21523 (N_21523,N_21369,N_21229);
nand U21524 (N_21524,N_21053,N_21174);
and U21525 (N_21525,N_21485,N_21348);
nor U21526 (N_21526,N_21043,N_21206);
or U21527 (N_21527,N_21089,N_21129);
xnor U21528 (N_21528,N_21457,N_21317);
or U21529 (N_21529,N_21461,N_21148);
and U21530 (N_21530,N_21182,N_21465);
xnor U21531 (N_21531,N_21187,N_21230);
and U21532 (N_21532,N_21285,N_21452);
nor U21533 (N_21533,N_21337,N_21479);
nand U21534 (N_21534,N_21030,N_21201);
or U21535 (N_21535,N_21200,N_21290);
xnor U21536 (N_21536,N_21470,N_21278);
nor U21537 (N_21537,N_21351,N_21262);
xor U21538 (N_21538,N_21462,N_21365);
nand U21539 (N_21539,N_21464,N_21436);
or U21540 (N_21540,N_21000,N_21143);
nor U21541 (N_21541,N_21090,N_21498);
nand U21542 (N_21542,N_21179,N_21469);
and U21543 (N_21543,N_21435,N_21081);
xnor U21544 (N_21544,N_21252,N_21038);
or U21545 (N_21545,N_21368,N_21170);
or U21546 (N_21546,N_21451,N_21328);
nand U21547 (N_21547,N_21467,N_21387);
xnor U21548 (N_21548,N_21455,N_21439);
nor U21549 (N_21549,N_21151,N_21420);
or U21550 (N_21550,N_21183,N_21204);
nand U21551 (N_21551,N_21265,N_21096);
xor U21552 (N_21552,N_21256,N_21429);
nand U21553 (N_21553,N_21222,N_21458);
or U21554 (N_21554,N_21453,N_21220);
nand U21555 (N_21555,N_21408,N_21460);
and U21556 (N_21556,N_21046,N_21352);
nor U21557 (N_21557,N_21325,N_21152);
and U21558 (N_21558,N_21269,N_21196);
xor U21559 (N_21559,N_21132,N_21427);
and U21560 (N_21560,N_21058,N_21146);
nor U21561 (N_21561,N_21340,N_21047);
nor U21562 (N_21562,N_21490,N_21032);
xnor U21563 (N_21563,N_21211,N_21015);
and U21564 (N_21564,N_21082,N_21326);
nor U21565 (N_21565,N_21124,N_21336);
xnor U21566 (N_21566,N_21011,N_21426);
and U21567 (N_21567,N_21306,N_21061);
nor U21568 (N_21568,N_21428,N_21473);
or U21569 (N_21569,N_21016,N_21140);
nand U21570 (N_21570,N_21121,N_21318);
nand U21571 (N_21571,N_21186,N_21416);
xnor U21572 (N_21572,N_21144,N_21245);
and U21573 (N_21573,N_21033,N_21311);
nor U21574 (N_21574,N_21051,N_21123);
and U21575 (N_21575,N_21209,N_21358);
nand U21576 (N_21576,N_21379,N_21297);
or U21577 (N_21577,N_21181,N_21065);
and U21578 (N_21578,N_21069,N_21257);
and U21579 (N_21579,N_21173,N_21165);
or U21580 (N_21580,N_21307,N_21216);
or U21581 (N_21581,N_21382,N_21158);
and U21582 (N_21582,N_21477,N_21277);
and U21583 (N_21583,N_21419,N_21238);
nor U21584 (N_21584,N_21034,N_21421);
nor U21585 (N_21585,N_21237,N_21338);
nor U21586 (N_21586,N_21396,N_21423);
nand U21587 (N_21587,N_21118,N_21483);
nand U21588 (N_21588,N_21398,N_21192);
xor U21589 (N_21589,N_21242,N_21098);
nand U21590 (N_21590,N_21282,N_21355);
nor U21591 (N_21591,N_21363,N_21160);
nand U21592 (N_21592,N_21074,N_21272);
nor U21593 (N_21593,N_21171,N_21251);
nand U21594 (N_21594,N_21223,N_21418);
nor U21595 (N_21595,N_21346,N_21362);
nand U21596 (N_21596,N_21371,N_21197);
xor U21597 (N_21597,N_21432,N_21018);
nand U21598 (N_21598,N_21157,N_21029);
or U21599 (N_21599,N_21316,N_21243);
nand U21600 (N_21600,N_21422,N_21357);
xnor U21601 (N_21601,N_21304,N_21142);
and U21602 (N_21602,N_21414,N_21294);
or U21603 (N_21603,N_21449,N_21323);
or U21604 (N_21604,N_21111,N_21131);
xnor U21605 (N_21605,N_21099,N_21049);
xnor U21606 (N_21606,N_21139,N_21218);
or U21607 (N_21607,N_21303,N_21399);
xnor U21608 (N_21608,N_21417,N_21066);
xor U21609 (N_21609,N_21288,N_21381);
xnor U21610 (N_21610,N_21258,N_21302);
nor U21611 (N_21611,N_21027,N_21014);
nand U21612 (N_21612,N_21083,N_21301);
nor U21613 (N_21613,N_21300,N_21359);
nand U21614 (N_21614,N_21022,N_21079);
or U21615 (N_21615,N_21207,N_21482);
nand U21616 (N_21616,N_21166,N_21281);
nand U21617 (N_21617,N_21107,N_21086);
nor U21618 (N_21618,N_21361,N_21271);
nand U21619 (N_21619,N_21017,N_21393);
nand U21620 (N_21620,N_21008,N_21405);
nand U21621 (N_21621,N_21092,N_21101);
and U21622 (N_21622,N_21003,N_21356);
nor U21623 (N_21623,N_21232,N_21406);
nand U21624 (N_21624,N_21377,N_21366);
and U21625 (N_21625,N_21026,N_21343);
nor U21626 (N_21626,N_21342,N_21441);
and U21627 (N_21627,N_21070,N_21445);
xor U21628 (N_21628,N_21494,N_21385);
nand U21629 (N_21629,N_21091,N_21134);
nor U21630 (N_21630,N_21009,N_21279);
nor U21631 (N_21631,N_21076,N_21035);
and U21632 (N_21632,N_21276,N_21137);
nand U21633 (N_21633,N_21063,N_21122);
and U21634 (N_21634,N_21402,N_21135);
or U21635 (N_21635,N_21172,N_21180);
nor U21636 (N_21636,N_21010,N_21259);
nor U21637 (N_21637,N_21446,N_21225);
and U21638 (N_21638,N_21202,N_21475);
or U21639 (N_21639,N_21138,N_21078);
or U21640 (N_21640,N_21407,N_21112);
xnor U21641 (N_21641,N_21253,N_21036);
xnor U21642 (N_21642,N_21433,N_21347);
or U21643 (N_21643,N_21095,N_21495);
xnor U21644 (N_21644,N_21044,N_21324);
nor U21645 (N_21645,N_21239,N_21189);
nor U21646 (N_21646,N_21484,N_21270);
nor U21647 (N_21647,N_21425,N_21330);
and U21648 (N_21648,N_21108,N_21314);
or U21649 (N_21649,N_21125,N_21203);
nor U21650 (N_21650,N_21113,N_21109);
and U21651 (N_21651,N_21350,N_21219);
nor U21652 (N_21652,N_21349,N_21057);
nand U21653 (N_21653,N_21296,N_21309);
nor U21654 (N_21654,N_21028,N_21481);
and U21655 (N_21655,N_21321,N_21221);
xor U21656 (N_21656,N_21041,N_21486);
xnor U21657 (N_21657,N_21198,N_21450);
nand U21658 (N_21658,N_21437,N_21161);
nor U21659 (N_21659,N_21048,N_21459);
xor U21660 (N_21660,N_21067,N_21075);
or U21661 (N_21661,N_21240,N_21430);
nor U21662 (N_21662,N_21291,N_21312);
nand U21663 (N_21663,N_21106,N_21412);
or U21664 (N_21664,N_21054,N_21228);
and U21665 (N_21665,N_21332,N_21084);
nand U21666 (N_21666,N_21360,N_21322);
or U21667 (N_21667,N_21004,N_21103);
nor U21668 (N_21668,N_21115,N_21411);
xor U21669 (N_21669,N_21333,N_21019);
nand U21670 (N_21670,N_21320,N_21097);
nor U21671 (N_21671,N_21214,N_21401);
or U21672 (N_21672,N_21339,N_21224);
nor U21673 (N_21673,N_21105,N_21246);
nand U21674 (N_21674,N_21319,N_21141);
nand U21675 (N_21675,N_21005,N_21213);
nor U21676 (N_21676,N_21353,N_21410);
nand U21677 (N_21677,N_21128,N_21413);
and U21678 (N_21678,N_21275,N_21334);
xnor U21679 (N_21679,N_21331,N_21060);
xnor U21680 (N_21680,N_21012,N_21231);
or U21681 (N_21681,N_21233,N_21178);
or U21682 (N_21682,N_21177,N_21191);
or U21683 (N_21683,N_21378,N_21391);
nor U21684 (N_21684,N_21247,N_21002);
nor U21685 (N_21685,N_21056,N_21274);
or U21686 (N_21686,N_21195,N_21080);
nand U21687 (N_21687,N_21466,N_21476);
nand U21688 (N_21688,N_21120,N_21190);
xnor U21689 (N_21689,N_21389,N_21327);
xnor U21690 (N_21690,N_21025,N_21127);
nor U21691 (N_21691,N_21364,N_21313);
and U21692 (N_21692,N_21354,N_21496);
nor U21693 (N_21693,N_21292,N_21167);
or U21694 (N_21694,N_21440,N_21235);
nor U21695 (N_21695,N_21383,N_21042);
nor U21696 (N_21696,N_21308,N_21163);
xnor U21697 (N_21697,N_21305,N_21471);
nand U21698 (N_21698,N_21072,N_21489);
and U21699 (N_21699,N_21266,N_21267);
xnor U21700 (N_21700,N_21264,N_21085);
and U21701 (N_21701,N_21394,N_21062);
xnor U21702 (N_21702,N_21241,N_21024);
and U21703 (N_21703,N_21487,N_21448);
nand U21704 (N_21704,N_21156,N_21286);
or U21705 (N_21705,N_21444,N_21244);
or U21706 (N_21706,N_21064,N_21114);
and U21707 (N_21707,N_21193,N_21147);
and U21708 (N_21708,N_21234,N_21329);
nor U21709 (N_21709,N_21210,N_21031);
nor U21710 (N_21710,N_21215,N_21341);
nor U21711 (N_21711,N_21110,N_21102);
nand U21712 (N_21712,N_21299,N_21254);
xor U21713 (N_21713,N_21100,N_21478);
or U21714 (N_21714,N_21050,N_21480);
nor U21715 (N_21715,N_21119,N_21071);
and U21716 (N_21716,N_21284,N_21447);
nand U21717 (N_21717,N_21208,N_21093);
or U21718 (N_21718,N_21088,N_21492);
or U21719 (N_21719,N_21367,N_21268);
nand U21720 (N_21720,N_21006,N_21153);
or U21721 (N_21721,N_21205,N_21380);
nand U21722 (N_21722,N_21164,N_21497);
and U21723 (N_21723,N_21185,N_21162);
or U21724 (N_21724,N_21472,N_21375);
nor U21725 (N_21725,N_21263,N_21415);
or U21726 (N_21726,N_21431,N_21280);
nand U21727 (N_21727,N_21217,N_21374);
nand U21728 (N_21728,N_21021,N_21373);
and U21729 (N_21729,N_21007,N_21087);
nor U21730 (N_21730,N_21116,N_21039);
nor U21731 (N_21731,N_21283,N_21442);
nor U21732 (N_21732,N_21248,N_21255);
xor U21733 (N_21733,N_21456,N_21023);
xor U21734 (N_21734,N_21150,N_21227);
nand U21735 (N_21735,N_21370,N_21059);
and U21736 (N_21736,N_21184,N_21424);
or U21737 (N_21737,N_21310,N_21176);
nor U21738 (N_21738,N_21136,N_21372);
nor U21739 (N_21739,N_21345,N_21013);
nor U21740 (N_21740,N_21454,N_21194);
and U21741 (N_21741,N_21390,N_21037);
nand U21742 (N_21742,N_21159,N_21154);
nand U21743 (N_21743,N_21126,N_21295);
nor U21744 (N_21744,N_21040,N_21499);
nand U21745 (N_21745,N_21212,N_21068);
xor U21746 (N_21746,N_21384,N_21052);
or U21747 (N_21747,N_21287,N_21130);
and U21748 (N_21748,N_21199,N_21175);
nand U21749 (N_21749,N_21493,N_21463);
and U21750 (N_21750,N_21487,N_21159);
and U21751 (N_21751,N_21043,N_21495);
xnor U21752 (N_21752,N_21399,N_21407);
or U21753 (N_21753,N_21223,N_21125);
nor U21754 (N_21754,N_21399,N_21492);
or U21755 (N_21755,N_21325,N_21290);
or U21756 (N_21756,N_21044,N_21286);
nor U21757 (N_21757,N_21236,N_21043);
nor U21758 (N_21758,N_21475,N_21291);
or U21759 (N_21759,N_21186,N_21404);
xnor U21760 (N_21760,N_21091,N_21089);
nand U21761 (N_21761,N_21493,N_21047);
xnor U21762 (N_21762,N_21154,N_21421);
nor U21763 (N_21763,N_21025,N_21102);
xor U21764 (N_21764,N_21342,N_21162);
nand U21765 (N_21765,N_21293,N_21054);
and U21766 (N_21766,N_21012,N_21124);
nand U21767 (N_21767,N_21360,N_21281);
xor U21768 (N_21768,N_21190,N_21083);
nor U21769 (N_21769,N_21304,N_21001);
nor U21770 (N_21770,N_21476,N_21448);
nand U21771 (N_21771,N_21140,N_21474);
and U21772 (N_21772,N_21346,N_21475);
xnor U21773 (N_21773,N_21350,N_21198);
nor U21774 (N_21774,N_21375,N_21053);
nor U21775 (N_21775,N_21254,N_21262);
nand U21776 (N_21776,N_21294,N_21401);
nand U21777 (N_21777,N_21024,N_21080);
nand U21778 (N_21778,N_21087,N_21237);
nor U21779 (N_21779,N_21247,N_21064);
xor U21780 (N_21780,N_21150,N_21312);
and U21781 (N_21781,N_21025,N_21064);
or U21782 (N_21782,N_21387,N_21187);
nand U21783 (N_21783,N_21080,N_21192);
xor U21784 (N_21784,N_21398,N_21150);
xor U21785 (N_21785,N_21307,N_21269);
xnor U21786 (N_21786,N_21210,N_21086);
or U21787 (N_21787,N_21249,N_21215);
and U21788 (N_21788,N_21301,N_21170);
nor U21789 (N_21789,N_21072,N_21039);
or U21790 (N_21790,N_21400,N_21406);
or U21791 (N_21791,N_21085,N_21028);
xor U21792 (N_21792,N_21162,N_21495);
and U21793 (N_21793,N_21247,N_21368);
or U21794 (N_21794,N_21104,N_21240);
xor U21795 (N_21795,N_21341,N_21167);
nand U21796 (N_21796,N_21487,N_21069);
nor U21797 (N_21797,N_21265,N_21150);
nor U21798 (N_21798,N_21442,N_21265);
nor U21799 (N_21799,N_21149,N_21044);
nand U21800 (N_21800,N_21212,N_21022);
and U21801 (N_21801,N_21443,N_21265);
nand U21802 (N_21802,N_21406,N_21384);
nor U21803 (N_21803,N_21382,N_21052);
nor U21804 (N_21804,N_21227,N_21313);
or U21805 (N_21805,N_21279,N_21435);
nand U21806 (N_21806,N_21499,N_21323);
xnor U21807 (N_21807,N_21495,N_21300);
or U21808 (N_21808,N_21353,N_21489);
and U21809 (N_21809,N_21004,N_21101);
xnor U21810 (N_21810,N_21210,N_21394);
or U21811 (N_21811,N_21379,N_21385);
nand U21812 (N_21812,N_21176,N_21097);
nor U21813 (N_21813,N_21454,N_21447);
and U21814 (N_21814,N_21311,N_21342);
xnor U21815 (N_21815,N_21201,N_21305);
nor U21816 (N_21816,N_21212,N_21025);
and U21817 (N_21817,N_21107,N_21069);
nand U21818 (N_21818,N_21410,N_21384);
xor U21819 (N_21819,N_21101,N_21174);
nor U21820 (N_21820,N_21123,N_21354);
or U21821 (N_21821,N_21053,N_21234);
or U21822 (N_21822,N_21303,N_21124);
nand U21823 (N_21823,N_21160,N_21135);
nand U21824 (N_21824,N_21446,N_21141);
and U21825 (N_21825,N_21213,N_21237);
nand U21826 (N_21826,N_21385,N_21303);
nand U21827 (N_21827,N_21407,N_21191);
xor U21828 (N_21828,N_21108,N_21170);
nand U21829 (N_21829,N_21080,N_21163);
or U21830 (N_21830,N_21015,N_21476);
nand U21831 (N_21831,N_21098,N_21095);
xnor U21832 (N_21832,N_21309,N_21251);
nor U21833 (N_21833,N_21406,N_21120);
or U21834 (N_21834,N_21175,N_21125);
nand U21835 (N_21835,N_21333,N_21165);
nand U21836 (N_21836,N_21303,N_21155);
nor U21837 (N_21837,N_21455,N_21140);
nand U21838 (N_21838,N_21435,N_21224);
or U21839 (N_21839,N_21305,N_21499);
nand U21840 (N_21840,N_21107,N_21179);
nand U21841 (N_21841,N_21395,N_21016);
nor U21842 (N_21842,N_21380,N_21371);
and U21843 (N_21843,N_21397,N_21466);
nand U21844 (N_21844,N_21009,N_21144);
nand U21845 (N_21845,N_21492,N_21196);
xnor U21846 (N_21846,N_21217,N_21298);
and U21847 (N_21847,N_21106,N_21177);
and U21848 (N_21848,N_21020,N_21268);
and U21849 (N_21849,N_21344,N_21346);
or U21850 (N_21850,N_21040,N_21478);
xor U21851 (N_21851,N_21384,N_21446);
nand U21852 (N_21852,N_21242,N_21116);
nand U21853 (N_21853,N_21428,N_21482);
and U21854 (N_21854,N_21485,N_21014);
xor U21855 (N_21855,N_21118,N_21258);
nand U21856 (N_21856,N_21401,N_21282);
and U21857 (N_21857,N_21403,N_21290);
or U21858 (N_21858,N_21085,N_21232);
nand U21859 (N_21859,N_21283,N_21425);
or U21860 (N_21860,N_21213,N_21230);
and U21861 (N_21861,N_21093,N_21181);
or U21862 (N_21862,N_21083,N_21126);
or U21863 (N_21863,N_21485,N_21013);
or U21864 (N_21864,N_21499,N_21042);
and U21865 (N_21865,N_21382,N_21280);
and U21866 (N_21866,N_21039,N_21152);
and U21867 (N_21867,N_21192,N_21228);
xor U21868 (N_21868,N_21025,N_21093);
nand U21869 (N_21869,N_21432,N_21085);
xor U21870 (N_21870,N_21306,N_21369);
xnor U21871 (N_21871,N_21145,N_21442);
nor U21872 (N_21872,N_21488,N_21081);
nand U21873 (N_21873,N_21098,N_21354);
and U21874 (N_21874,N_21001,N_21460);
nand U21875 (N_21875,N_21203,N_21023);
xor U21876 (N_21876,N_21072,N_21474);
xnor U21877 (N_21877,N_21222,N_21245);
nand U21878 (N_21878,N_21468,N_21034);
and U21879 (N_21879,N_21172,N_21281);
and U21880 (N_21880,N_21061,N_21041);
and U21881 (N_21881,N_21320,N_21324);
nand U21882 (N_21882,N_21260,N_21479);
or U21883 (N_21883,N_21108,N_21072);
nand U21884 (N_21884,N_21489,N_21288);
or U21885 (N_21885,N_21484,N_21148);
xor U21886 (N_21886,N_21402,N_21387);
nor U21887 (N_21887,N_21260,N_21135);
nand U21888 (N_21888,N_21342,N_21268);
and U21889 (N_21889,N_21194,N_21007);
nand U21890 (N_21890,N_21233,N_21040);
nor U21891 (N_21891,N_21116,N_21488);
nand U21892 (N_21892,N_21041,N_21267);
or U21893 (N_21893,N_21116,N_21233);
or U21894 (N_21894,N_21354,N_21361);
xnor U21895 (N_21895,N_21002,N_21080);
and U21896 (N_21896,N_21238,N_21427);
and U21897 (N_21897,N_21241,N_21298);
or U21898 (N_21898,N_21084,N_21039);
xnor U21899 (N_21899,N_21457,N_21446);
xor U21900 (N_21900,N_21253,N_21083);
xor U21901 (N_21901,N_21049,N_21327);
or U21902 (N_21902,N_21308,N_21499);
xnor U21903 (N_21903,N_21046,N_21492);
and U21904 (N_21904,N_21171,N_21338);
and U21905 (N_21905,N_21388,N_21166);
xnor U21906 (N_21906,N_21184,N_21090);
nand U21907 (N_21907,N_21149,N_21130);
nand U21908 (N_21908,N_21415,N_21359);
nand U21909 (N_21909,N_21166,N_21195);
xor U21910 (N_21910,N_21289,N_21007);
xnor U21911 (N_21911,N_21240,N_21413);
nor U21912 (N_21912,N_21202,N_21107);
and U21913 (N_21913,N_21232,N_21470);
nand U21914 (N_21914,N_21110,N_21443);
nand U21915 (N_21915,N_21410,N_21028);
nor U21916 (N_21916,N_21136,N_21260);
nor U21917 (N_21917,N_21354,N_21039);
xnor U21918 (N_21918,N_21273,N_21378);
nand U21919 (N_21919,N_21098,N_21185);
and U21920 (N_21920,N_21034,N_21233);
or U21921 (N_21921,N_21494,N_21345);
nor U21922 (N_21922,N_21408,N_21491);
xnor U21923 (N_21923,N_21263,N_21458);
nand U21924 (N_21924,N_21397,N_21078);
nand U21925 (N_21925,N_21057,N_21175);
nor U21926 (N_21926,N_21013,N_21161);
nand U21927 (N_21927,N_21351,N_21331);
or U21928 (N_21928,N_21410,N_21135);
and U21929 (N_21929,N_21003,N_21471);
or U21930 (N_21930,N_21112,N_21041);
xnor U21931 (N_21931,N_21480,N_21056);
nand U21932 (N_21932,N_21154,N_21020);
xnor U21933 (N_21933,N_21107,N_21281);
and U21934 (N_21934,N_21408,N_21152);
or U21935 (N_21935,N_21215,N_21338);
xor U21936 (N_21936,N_21447,N_21147);
xnor U21937 (N_21937,N_21270,N_21297);
or U21938 (N_21938,N_21378,N_21205);
and U21939 (N_21939,N_21340,N_21399);
or U21940 (N_21940,N_21066,N_21137);
xor U21941 (N_21941,N_21209,N_21465);
and U21942 (N_21942,N_21022,N_21000);
or U21943 (N_21943,N_21026,N_21420);
or U21944 (N_21944,N_21377,N_21475);
or U21945 (N_21945,N_21122,N_21149);
xor U21946 (N_21946,N_21477,N_21207);
xor U21947 (N_21947,N_21141,N_21140);
or U21948 (N_21948,N_21092,N_21164);
nand U21949 (N_21949,N_21045,N_21339);
or U21950 (N_21950,N_21425,N_21095);
or U21951 (N_21951,N_21235,N_21460);
nand U21952 (N_21952,N_21151,N_21302);
nor U21953 (N_21953,N_21427,N_21047);
xnor U21954 (N_21954,N_21259,N_21196);
nor U21955 (N_21955,N_21363,N_21370);
xnor U21956 (N_21956,N_21149,N_21003);
nand U21957 (N_21957,N_21352,N_21112);
xor U21958 (N_21958,N_21382,N_21377);
or U21959 (N_21959,N_21235,N_21195);
nand U21960 (N_21960,N_21351,N_21465);
or U21961 (N_21961,N_21380,N_21429);
and U21962 (N_21962,N_21109,N_21350);
and U21963 (N_21963,N_21430,N_21179);
xnor U21964 (N_21964,N_21297,N_21197);
and U21965 (N_21965,N_21453,N_21471);
nand U21966 (N_21966,N_21367,N_21147);
xor U21967 (N_21967,N_21126,N_21078);
nor U21968 (N_21968,N_21002,N_21497);
xor U21969 (N_21969,N_21153,N_21121);
xnor U21970 (N_21970,N_21068,N_21023);
xor U21971 (N_21971,N_21317,N_21205);
nand U21972 (N_21972,N_21124,N_21329);
nand U21973 (N_21973,N_21432,N_21461);
and U21974 (N_21974,N_21275,N_21218);
and U21975 (N_21975,N_21305,N_21323);
or U21976 (N_21976,N_21179,N_21404);
nand U21977 (N_21977,N_21457,N_21404);
or U21978 (N_21978,N_21379,N_21063);
xor U21979 (N_21979,N_21469,N_21481);
nor U21980 (N_21980,N_21141,N_21388);
nand U21981 (N_21981,N_21383,N_21447);
or U21982 (N_21982,N_21397,N_21062);
and U21983 (N_21983,N_21095,N_21060);
and U21984 (N_21984,N_21100,N_21331);
nor U21985 (N_21985,N_21250,N_21125);
or U21986 (N_21986,N_21030,N_21296);
and U21987 (N_21987,N_21406,N_21184);
or U21988 (N_21988,N_21024,N_21454);
nand U21989 (N_21989,N_21457,N_21313);
nand U21990 (N_21990,N_21231,N_21217);
nand U21991 (N_21991,N_21473,N_21206);
and U21992 (N_21992,N_21491,N_21348);
and U21993 (N_21993,N_21404,N_21102);
and U21994 (N_21994,N_21045,N_21481);
nor U21995 (N_21995,N_21398,N_21495);
xor U21996 (N_21996,N_21355,N_21415);
or U21997 (N_21997,N_21462,N_21136);
nor U21998 (N_21998,N_21313,N_21343);
and U21999 (N_21999,N_21321,N_21155);
or U22000 (N_22000,N_21638,N_21722);
xor U22001 (N_22001,N_21560,N_21959);
or U22002 (N_22002,N_21792,N_21681);
nand U22003 (N_22003,N_21639,N_21993);
and U22004 (N_22004,N_21575,N_21589);
xor U22005 (N_22005,N_21509,N_21964);
or U22006 (N_22006,N_21502,N_21545);
nand U22007 (N_22007,N_21776,N_21745);
xnor U22008 (N_22008,N_21716,N_21797);
nand U22009 (N_22009,N_21944,N_21724);
nor U22010 (N_22010,N_21862,N_21652);
xnor U22011 (N_22011,N_21637,N_21885);
or U22012 (N_22012,N_21860,N_21867);
nand U22013 (N_22013,N_21826,N_21678);
or U22014 (N_22014,N_21870,N_21999);
nor U22015 (N_22015,N_21978,N_21768);
nor U22016 (N_22016,N_21613,N_21742);
or U22017 (N_22017,N_21780,N_21778);
or U22018 (N_22018,N_21705,N_21680);
or U22019 (N_22019,N_21900,N_21510);
nor U22020 (N_22020,N_21536,N_21901);
xnor U22021 (N_22021,N_21968,N_21789);
or U22022 (N_22022,N_21715,N_21773);
or U22023 (N_22023,N_21838,N_21933);
xor U22024 (N_22024,N_21597,N_21812);
nor U22025 (N_22025,N_21730,N_21833);
xnor U22026 (N_22026,N_21774,N_21903);
nor U22027 (N_22027,N_21522,N_21965);
xnor U22028 (N_22028,N_21887,N_21857);
or U22029 (N_22029,N_21854,N_21863);
and U22030 (N_22030,N_21634,N_21525);
nand U22031 (N_22031,N_21615,N_21620);
nand U22032 (N_22032,N_21759,N_21696);
nor U22033 (N_22033,N_21523,N_21769);
and U22034 (N_22034,N_21878,N_21704);
nor U22035 (N_22035,N_21518,N_21626);
and U22036 (N_22036,N_21700,N_21853);
and U22037 (N_22037,N_21654,N_21579);
and U22038 (N_22038,N_21594,N_21707);
nand U22039 (N_22039,N_21967,N_21922);
nand U22040 (N_22040,N_21849,N_21586);
xnor U22041 (N_22041,N_21985,N_21843);
or U22042 (N_22042,N_21657,N_21517);
xnor U22043 (N_22043,N_21512,N_21767);
xor U22044 (N_22044,N_21658,N_21784);
or U22045 (N_22045,N_21976,N_21568);
xnor U22046 (N_22046,N_21754,N_21874);
xor U22047 (N_22047,N_21814,N_21952);
or U22048 (N_22048,N_21701,N_21848);
or U22049 (N_22049,N_21617,N_21932);
nand U22050 (N_22050,N_21749,N_21864);
and U22051 (N_22051,N_21669,N_21732);
nor U22052 (N_22052,N_21636,N_21635);
nand U22053 (N_22053,N_21840,N_21771);
and U22054 (N_22054,N_21547,N_21736);
nand U22055 (N_22055,N_21795,N_21529);
and U22056 (N_22056,N_21508,N_21740);
nor U22057 (N_22057,N_21832,N_21851);
nor U22058 (N_22058,N_21915,N_21621);
nand U22059 (N_22059,N_21850,N_21643);
nor U22060 (N_22060,N_21905,N_21939);
nor U22061 (N_22061,N_21896,N_21582);
xnor U22062 (N_22062,N_21817,N_21645);
and U22063 (N_22063,N_21604,N_21734);
and U22064 (N_22064,N_21917,N_21721);
xor U22065 (N_22065,N_21894,N_21835);
or U22066 (N_22066,N_21514,N_21892);
or U22067 (N_22067,N_21747,N_21852);
and U22068 (N_22068,N_21893,N_21899);
nand U22069 (N_22069,N_21682,N_21764);
and U22070 (N_22070,N_21672,N_21962);
nand U22071 (N_22071,N_21709,N_21982);
or U22072 (N_22072,N_21554,N_21569);
xor U22073 (N_22073,N_21543,N_21690);
nor U22074 (N_22074,N_21844,N_21880);
nor U22075 (N_22075,N_21738,N_21719);
or U22076 (N_22076,N_21983,N_21783);
and U22077 (N_22077,N_21760,N_21666);
xor U22078 (N_22078,N_21623,N_21895);
xor U22079 (N_22079,N_21971,N_21611);
and U22080 (N_22080,N_21875,N_21839);
xor U22081 (N_22081,N_21744,N_21630);
or U22082 (N_22082,N_21607,N_21649);
nand U22083 (N_22083,N_21600,N_21866);
and U22084 (N_22084,N_21520,N_21741);
or U22085 (N_22085,N_21691,N_21775);
xor U22086 (N_22086,N_21820,N_21912);
nor U22087 (N_22087,N_21961,N_21631);
nor U22088 (N_22088,N_21949,N_21616);
xnor U22089 (N_22089,N_21923,N_21541);
or U22090 (N_22090,N_21947,N_21818);
nand U22091 (N_22091,N_21661,N_21998);
nand U22092 (N_22092,N_21981,N_21929);
nor U22093 (N_22093,N_21539,N_21650);
or U22094 (N_22094,N_21931,N_21928);
xor U22095 (N_22095,N_21717,N_21606);
xnor U22096 (N_22096,N_21565,N_21934);
or U22097 (N_22097,N_21946,N_21772);
nor U22098 (N_22098,N_21549,N_21969);
xor U22099 (N_22099,N_21587,N_21625);
nand U22100 (N_22100,N_21511,N_21927);
or U22101 (N_22101,N_21557,N_21914);
nor U22102 (N_22102,N_21533,N_21556);
nor U22103 (N_22103,N_21897,N_21803);
xnor U22104 (N_22104,N_21561,N_21941);
nor U22105 (N_22105,N_21788,N_21632);
or U22106 (N_22106,N_21913,N_21642);
nand U22107 (N_22107,N_21656,N_21675);
nand U22108 (N_22108,N_21994,N_21618);
nand U22109 (N_22109,N_21530,N_21662);
nand U22110 (N_22110,N_21954,N_21564);
xor U22111 (N_22111,N_21770,N_21723);
nor U22112 (N_22112,N_21567,N_21603);
xor U22113 (N_22113,N_21550,N_21801);
and U22114 (N_22114,N_21920,N_21842);
nor U22115 (N_22115,N_21515,N_21610);
or U22116 (N_22116,N_21697,N_21679);
nor U22117 (N_22117,N_21940,N_21871);
and U22118 (N_22118,N_21753,N_21629);
nand U22119 (N_22119,N_21703,N_21677);
and U22120 (N_22120,N_21644,N_21980);
nor U22121 (N_22121,N_21825,N_21823);
and U22122 (N_22122,N_21943,N_21712);
or U22123 (N_22123,N_21816,N_21785);
and U22124 (N_22124,N_21937,N_21910);
xnor U22125 (N_22125,N_21811,N_21648);
nand U22126 (N_22126,N_21755,N_21601);
and U22127 (N_22127,N_21956,N_21879);
nor U22128 (N_22128,N_21845,N_21595);
or U22129 (N_22129,N_21687,N_21787);
nor U22130 (N_22130,N_21918,N_21651);
nor U22131 (N_22131,N_21655,N_21726);
or U22132 (N_22132,N_21641,N_21997);
and U22133 (N_22133,N_21670,N_21861);
and U22134 (N_22134,N_21868,N_21828);
nand U22135 (N_22135,N_21519,N_21751);
or U22136 (N_22136,N_21667,N_21537);
or U22137 (N_22137,N_21966,N_21542);
nor U22138 (N_22138,N_21668,N_21526);
and U22139 (N_22139,N_21673,N_21806);
nor U22140 (N_22140,N_21809,N_21951);
nor U22141 (N_22141,N_21781,N_21988);
xnor U22142 (N_22142,N_21873,N_21752);
xor U22143 (N_22143,N_21622,N_21794);
xor U22144 (N_22144,N_21846,N_21647);
xor U22145 (N_22145,N_21693,N_21889);
or U22146 (N_22146,N_21714,N_21970);
xor U22147 (N_22147,N_21907,N_21583);
or U22148 (N_22148,N_21612,N_21599);
and U22149 (N_22149,N_21653,N_21869);
nor U22150 (N_22150,N_21566,N_21945);
and U22151 (N_22151,N_21761,N_21763);
and U22152 (N_22152,N_21505,N_21501);
nor U22153 (N_22153,N_21614,N_21802);
and U22154 (N_22154,N_21608,N_21572);
and U22155 (N_22155,N_21528,N_21824);
and U22156 (N_22156,N_21663,N_21591);
or U22157 (N_22157,N_21674,N_21698);
nand U22158 (N_22158,N_21975,N_21735);
nor U22159 (N_22159,N_21727,N_21916);
nor U22160 (N_22160,N_21737,N_21890);
nand U22161 (N_22161,N_21718,N_21936);
nor U22162 (N_22162,N_21555,N_21577);
and U22163 (N_22163,N_21979,N_21757);
and U22164 (N_22164,N_21562,N_21986);
nand U22165 (N_22165,N_21713,N_21743);
xor U22166 (N_22166,N_21989,N_21746);
xor U22167 (N_22167,N_21688,N_21633);
or U22168 (N_22168,N_21960,N_21596);
or U22169 (N_22169,N_21881,N_21911);
nor U22170 (N_22170,N_21991,N_21884);
nor U22171 (N_22171,N_21909,N_21908);
nor U22172 (N_22172,N_21585,N_21559);
nor U22173 (N_22173,N_21563,N_21856);
or U22174 (N_22174,N_21777,N_21748);
or U22175 (N_22175,N_21827,N_21782);
nor U22176 (N_22176,N_21921,N_21521);
nor U22177 (N_22177,N_21858,N_21588);
nand U22178 (N_22178,N_21963,N_21686);
or U22179 (N_22179,N_21834,N_21977);
or U22180 (N_22180,N_21859,N_21796);
or U22181 (N_22181,N_21882,N_21695);
and U22182 (N_22182,N_21646,N_21847);
xnor U22183 (N_22183,N_21711,N_21804);
and U22184 (N_22184,N_21762,N_21888);
nor U22185 (N_22185,N_21807,N_21808);
nand U22186 (N_22186,N_21831,N_21791);
xnor U22187 (N_22187,N_21948,N_21584);
and U22188 (N_22188,N_21731,N_21957);
nor U22189 (N_22189,N_21725,N_21955);
nor U22190 (N_22190,N_21904,N_21500);
nor U22191 (N_22191,N_21995,N_21671);
and U22192 (N_22192,N_21942,N_21627);
nand U22193 (N_22193,N_21786,N_21974);
nor U22194 (N_22194,N_21972,N_21506);
nor U22195 (N_22195,N_21544,N_21930);
nand U22196 (N_22196,N_21739,N_21513);
or U22197 (N_22197,N_21779,N_21938);
nand U22198 (N_22198,N_21609,N_21571);
nor U22199 (N_22199,N_21699,N_21958);
nand U22200 (N_22200,N_21593,N_21576);
and U22201 (N_22201,N_21619,N_21822);
xor U22202 (N_22202,N_21659,N_21935);
or U22203 (N_22203,N_21628,N_21708);
or U22204 (N_22204,N_21602,N_21837);
and U22205 (N_22205,N_21919,N_21685);
nor U22206 (N_22206,N_21992,N_21706);
or U22207 (N_22207,N_21953,N_21819);
nor U22208 (N_22208,N_21877,N_21507);
nor U22209 (N_22209,N_21660,N_21684);
nand U22210 (N_22210,N_21558,N_21527);
xor U22211 (N_22211,N_21876,N_21702);
and U22212 (N_22212,N_21570,N_21765);
nand U22213 (N_22213,N_21973,N_21640);
xnor U22214 (N_22214,N_21793,N_21798);
and U22215 (N_22215,N_21624,N_21590);
nor U22216 (N_22216,N_21720,N_21598);
nor U22217 (N_22217,N_21872,N_21551);
and U22218 (N_22218,N_21710,N_21950);
xor U22219 (N_22219,N_21924,N_21813);
nand U22220 (N_22220,N_21578,N_21580);
and U22221 (N_22221,N_21548,N_21503);
xor U22222 (N_22222,N_21592,N_21524);
nand U22223 (N_22223,N_21664,N_21552);
xnor U22224 (N_22224,N_21553,N_21865);
nand U22225 (N_22225,N_21540,N_21676);
nor U22226 (N_22226,N_21689,N_21830);
nand U22227 (N_22227,N_21574,N_21836);
and U22228 (N_22228,N_21504,N_21926);
and U22229 (N_22229,N_21534,N_21692);
nand U22230 (N_22230,N_21799,N_21573);
and U22231 (N_22231,N_21516,N_21750);
nor U22232 (N_22232,N_21886,N_21758);
xnor U22233 (N_22233,N_21902,N_21841);
nor U22234 (N_22234,N_21532,N_21683);
nor U22235 (N_22235,N_21800,N_21906);
or U22236 (N_22236,N_21766,N_21898);
nor U22237 (N_22237,N_21984,N_21815);
xor U22238 (N_22238,N_21821,N_21729);
or U22239 (N_22239,N_21790,N_21756);
xnor U22240 (N_22240,N_21996,N_21535);
nand U22241 (N_22241,N_21694,N_21987);
xnor U22242 (N_22242,N_21733,N_21531);
and U22243 (N_22243,N_21810,N_21829);
or U22244 (N_22244,N_21805,N_21665);
xor U22245 (N_22245,N_21581,N_21925);
xnor U22246 (N_22246,N_21990,N_21546);
or U22247 (N_22247,N_21891,N_21605);
or U22248 (N_22248,N_21728,N_21883);
nand U22249 (N_22249,N_21855,N_21538);
xnor U22250 (N_22250,N_21773,N_21781);
and U22251 (N_22251,N_21597,N_21971);
or U22252 (N_22252,N_21512,N_21837);
xor U22253 (N_22253,N_21787,N_21605);
and U22254 (N_22254,N_21544,N_21732);
nand U22255 (N_22255,N_21944,N_21891);
and U22256 (N_22256,N_21883,N_21774);
or U22257 (N_22257,N_21676,N_21986);
nand U22258 (N_22258,N_21835,N_21725);
and U22259 (N_22259,N_21564,N_21808);
nand U22260 (N_22260,N_21502,N_21784);
or U22261 (N_22261,N_21523,N_21849);
or U22262 (N_22262,N_21829,N_21903);
nand U22263 (N_22263,N_21867,N_21896);
xnor U22264 (N_22264,N_21835,N_21680);
nand U22265 (N_22265,N_21972,N_21847);
xnor U22266 (N_22266,N_21710,N_21658);
xor U22267 (N_22267,N_21932,N_21538);
nor U22268 (N_22268,N_21800,N_21718);
or U22269 (N_22269,N_21796,N_21906);
or U22270 (N_22270,N_21728,N_21658);
or U22271 (N_22271,N_21664,N_21790);
or U22272 (N_22272,N_21529,N_21839);
and U22273 (N_22273,N_21662,N_21978);
and U22274 (N_22274,N_21513,N_21900);
or U22275 (N_22275,N_21583,N_21761);
nor U22276 (N_22276,N_21678,N_21842);
and U22277 (N_22277,N_21575,N_21905);
or U22278 (N_22278,N_21594,N_21776);
and U22279 (N_22279,N_21617,N_21614);
or U22280 (N_22280,N_21616,N_21956);
xor U22281 (N_22281,N_21606,N_21990);
xor U22282 (N_22282,N_21812,N_21963);
xnor U22283 (N_22283,N_21772,N_21562);
xor U22284 (N_22284,N_21712,N_21703);
and U22285 (N_22285,N_21563,N_21661);
and U22286 (N_22286,N_21780,N_21632);
nand U22287 (N_22287,N_21815,N_21606);
or U22288 (N_22288,N_21809,N_21698);
nand U22289 (N_22289,N_21588,N_21799);
xor U22290 (N_22290,N_21757,N_21707);
nand U22291 (N_22291,N_21824,N_21742);
xnor U22292 (N_22292,N_21864,N_21924);
nand U22293 (N_22293,N_21745,N_21777);
or U22294 (N_22294,N_21668,N_21920);
xor U22295 (N_22295,N_21948,N_21731);
xor U22296 (N_22296,N_21508,N_21857);
xor U22297 (N_22297,N_21521,N_21874);
nand U22298 (N_22298,N_21556,N_21955);
nand U22299 (N_22299,N_21520,N_21771);
nand U22300 (N_22300,N_21818,N_21968);
xor U22301 (N_22301,N_21930,N_21630);
and U22302 (N_22302,N_21638,N_21648);
nand U22303 (N_22303,N_21856,N_21637);
xor U22304 (N_22304,N_21655,N_21748);
nand U22305 (N_22305,N_21961,N_21823);
xor U22306 (N_22306,N_21847,N_21833);
nor U22307 (N_22307,N_21705,N_21732);
or U22308 (N_22308,N_21693,N_21625);
nor U22309 (N_22309,N_21934,N_21764);
nor U22310 (N_22310,N_21731,N_21576);
and U22311 (N_22311,N_21887,N_21778);
nor U22312 (N_22312,N_21515,N_21602);
and U22313 (N_22313,N_21581,N_21513);
xnor U22314 (N_22314,N_21817,N_21770);
nor U22315 (N_22315,N_21539,N_21814);
nand U22316 (N_22316,N_21634,N_21645);
nor U22317 (N_22317,N_21739,N_21723);
or U22318 (N_22318,N_21885,N_21692);
nand U22319 (N_22319,N_21699,N_21661);
xnor U22320 (N_22320,N_21940,N_21727);
nor U22321 (N_22321,N_21609,N_21729);
nor U22322 (N_22322,N_21696,N_21666);
and U22323 (N_22323,N_21969,N_21945);
or U22324 (N_22324,N_21610,N_21884);
or U22325 (N_22325,N_21637,N_21987);
or U22326 (N_22326,N_21692,N_21586);
or U22327 (N_22327,N_21649,N_21763);
or U22328 (N_22328,N_21820,N_21793);
and U22329 (N_22329,N_21906,N_21678);
nor U22330 (N_22330,N_21946,N_21776);
and U22331 (N_22331,N_21769,N_21891);
nor U22332 (N_22332,N_21842,N_21982);
nand U22333 (N_22333,N_21577,N_21689);
xor U22334 (N_22334,N_21532,N_21767);
or U22335 (N_22335,N_21710,N_21851);
xnor U22336 (N_22336,N_21770,N_21740);
and U22337 (N_22337,N_21915,N_21706);
and U22338 (N_22338,N_21717,N_21602);
xor U22339 (N_22339,N_21953,N_21607);
and U22340 (N_22340,N_21685,N_21873);
xor U22341 (N_22341,N_21578,N_21689);
and U22342 (N_22342,N_21537,N_21693);
xnor U22343 (N_22343,N_21646,N_21750);
nand U22344 (N_22344,N_21620,N_21519);
and U22345 (N_22345,N_21986,N_21846);
and U22346 (N_22346,N_21565,N_21824);
nor U22347 (N_22347,N_21796,N_21974);
xor U22348 (N_22348,N_21963,N_21848);
nand U22349 (N_22349,N_21769,N_21568);
or U22350 (N_22350,N_21865,N_21566);
nor U22351 (N_22351,N_21658,N_21749);
or U22352 (N_22352,N_21747,N_21578);
nor U22353 (N_22353,N_21592,N_21614);
nor U22354 (N_22354,N_21560,N_21739);
nor U22355 (N_22355,N_21718,N_21656);
and U22356 (N_22356,N_21722,N_21634);
nor U22357 (N_22357,N_21764,N_21611);
nor U22358 (N_22358,N_21542,N_21936);
xnor U22359 (N_22359,N_21597,N_21963);
xnor U22360 (N_22360,N_21682,N_21833);
xor U22361 (N_22361,N_21584,N_21873);
nand U22362 (N_22362,N_21854,N_21652);
and U22363 (N_22363,N_21953,N_21717);
and U22364 (N_22364,N_21932,N_21560);
and U22365 (N_22365,N_21525,N_21937);
or U22366 (N_22366,N_21602,N_21826);
xor U22367 (N_22367,N_21792,N_21970);
nand U22368 (N_22368,N_21683,N_21988);
and U22369 (N_22369,N_21654,N_21732);
xnor U22370 (N_22370,N_21737,N_21503);
nor U22371 (N_22371,N_21779,N_21506);
or U22372 (N_22372,N_21613,N_21909);
and U22373 (N_22373,N_21769,N_21824);
and U22374 (N_22374,N_21734,N_21808);
nor U22375 (N_22375,N_21504,N_21931);
xnor U22376 (N_22376,N_21829,N_21553);
nor U22377 (N_22377,N_21515,N_21642);
or U22378 (N_22378,N_21954,N_21999);
or U22379 (N_22379,N_21538,N_21933);
xnor U22380 (N_22380,N_21815,N_21931);
or U22381 (N_22381,N_21969,N_21980);
xnor U22382 (N_22382,N_21974,N_21709);
or U22383 (N_22383,N_21670,N_21749);
nor U22384 (N_22384,N_21638,N_21652);
nand U22385 (N_22385,N_21687,N_21786);
and U22386 (N_22386,N_21504,N_21962);
nand U22387 (N_22387,N_21646,N_21706);
or U22388 (N_22388,N_21514,N_21880);
nor U22389 (N_22389,N_21993,N_21691);
nor U22390 (N_22390,N_21708,N_21937);
nor U22391 (N_22391,N_21599,N_21752);
nand U22392 (N_22392,N_21570,N_21783);
and U22393 (N_22393,N_21880,N_21851);
and U22394 (N_22394,N_21618,N_21811);
and U22395 (N_22395,N_21636,N_21943);
and U22396 (N_22396,N_21953,N_21713);
nand U22397 (N_22397,N_21681,N_21741);
xor U22398 (N_22398,N_21913,N_21504);
nor U22399 (N_22399,N_21552,N_21853);
or U22400 (N_22400,N_21946,N_21856);
nor U22401 (N_22401,N_21898,N_21961);
xor U22402 (N_22402,N_21804,N_21910);
nand U22403 (N_22403,N_21958,N_21779);
nand U22404 (N_22404,N_21641,N_21608);
or U22405 (N_22405,N_21662,N_21751);
nor U22406 (N_22406,N_21883,N_21585);
xor U22407 (N_22407,N_21881,N_21678);
nor U22408 (N_22408,N_21965,N_21783);
nor U22409 (N_22409,N_21665,N_21687);
nand U22410 (N_22410,N_21940,N_21634);
or U22411 (N_22411,N_21613,N_21589);
or U22412 (N_22412,N_21700,N_21670);
nor U22413 (N_22413,N_21608,N_21532);
and U22414 (N_22414,N_21694,N_21775);
and U22415 (N_22415,N_21898,N_21644);
and U22416 (N_22416,N_21780,N_21758);
or U22417 (N_22417,N_21813,N_21734);
or U22418 (N_22418,N_21919,N_21879);
and U22419 (N_22419,N_21609,N_21615);
nand U22420 (N_22420,N_21694,N_21791);
xor U22421 (N_22421,N_21600,N_21931);
xnor U22422 (N_22422,N_21737,N_21629);
xnor U22423 (N_22423,N_21974,N_21928);
xor U22424 (N_22424,N_21697,N_21754);
nor U22425 (N_22425,N_21834,N_21547);
nor U22426 (N_22426,N_21591,N_21707);
and U22427 (N_22427,N_21736,N_21616);
xor U22428 (N_22428,N_21870,N_21881);
and U22429 (N_22429,N_21904,N_21995);
nand U22430 (N_22430,N_21566,N_21930);
nor U22431 (N_22431,N_21573,N_21777);
nor U22432 (N_22432,N_21947,N_21871);
or U22433 (N_22433,N_21813,N_21654);
nor U22434 (N_22434,N_21709,N_21789);
nor U22435 (N_22435,N_21701,N_21674);
nand U22436 (N_22436,N_21563,N_21914);
or U22437 (N_22437,N_21866,N_21991);
xor U22438 (N_22438,N_21928,N_21805);
and U22439 (N_22439,N_21907,N_21765);
or U22440 (N_22440,N_21920,N_21951);
xor U22441 (N_22441,N_21827,N_21664);
nor U22442 (N_22442,N_21860,N_21783);
nand U22443 (N_22443,N_21540,N_21980);
nand U22444 (N_22444,N_21896,N_21801);
and U22445 (N_22445,N_21883,N_21896);
or U22446 (N_22446,N_21847,N_21517);
and U22447 (N_22447,N_21861,N_21572);
or U22448 (N_22448,N_21861,N_21527);
nand U22449 (N_22449,N_21830,N_21796);
xnor U22450 (N_22450,N_21820,N_21825);
nand U22451 (N_22451,N_21879,N_21993);
xnor U22452 (N_22452,N_21630,N_21835);
or U22453 (N_22453,N_21545,N_21940);
nand U22454 (N_22454,N_21816,N_21671);
or U22455 (N_22455,N_21696,N_21551);
xor U22456 (N_22456,N_21920,N_21538);
nand U22457 (N_22457,N_21915,N_21955);
or U22458 (N_22458,N_21758,N_21579);
nand U22459 (N_22459,N_21589,N_21648);
or U22460 (N_22460,N_21996,N_21932);
and U22461 (N_22461,N_21762,N_21918);
or U22462 (N_22462,N_21675,N_21500);
nand U22463 (N_22463,N_21825,N_21615);
nor U22464 (N_22464,N_21699,N_21847);
or U22465 (N_22465,N_21797,N_21695);
or U22466 (N_22466,N_21743,N_21942);
xnor U22467 (N_22467,N_21925,N_21966);
and U22468 (N_22468,N_21766,N_21580);
nor U22469 (N_22469,N_21879,N_21510);
or U22470 (N_22470,N_21905,N_21729);
and U22471 (N_22471,N_21716,N_21670);
xnor U22472 (N_22472,N_21842,N_21752);
nand U22473 (N_22473,N_21678,N_21782);
xnor U22474 (N_22474,N_21972,N_21832);
nor U22475 (N_22475,N_21561,N_21878);
or U22476 (N_22476,N_21780,N_21935);
or U22477 (N_22477,N_21518,N_21660);
and U22478 (N_22478,N_21507,N_21674);
xor U22479 (N_22479,N_21745,N_21990);
xor U22480 (N_22480,N_21626,N_21796);
or U22481 (N_22481,N_21897,N_21543);
nand U22482 (N_22482,N_21695,N_21731);
nor U22483 (N_22483,N_21976,N_21804);
or U22484 (N_22484,N_21822,N_21687);
or U22485 (N_22485,N_21853,N_21787);
xor U22486 (N_22486,N_21646,N_21661);
nor U22487 (N_22487,N_21637,N_21561);
xnor U22488 (N_22488,N_21900,N_21835);
xor U22489 (N_22489,N_21810,N_21889);
xnor U22490 (N_22490,N_21879,N_21815);
or U22491 (N_22491,N_21549,N_21739);
nor U22492 (N_22492,N_21577,N_21736);
xnor U22493 (N_22493,N_21530,N_21632);
xor U22494 (N_22494,N_21868,N_21871);
xor U22495 (N_22495,N_21593,N_21712);
nor U22496 (N_22496,N_21959,N_21603);
and U22497 (N_22497,N_21588,N_21976);
xor U22498 (N_22498,N_21690,N_21616);
or U22499 (N_22499,N_21612,N_21897);
xnor U22500 (N_22500,N_22396,N_22363);
or U22501 (N_22501,N_22357,N_22092);
nor U22502 (N_22502,N_22351,N_22206);
nand U22503 (N_22503,N_22065,N_22313);
nor U22504 (N_22504,N_22484,N_22094);
or U22505 (N_22505,N_22200,N_22441);
xnor U22506 (N_22506,N_22430,N_22075);
nand U22507 (N_22507,N_22290,N_22390);
xor U22508 (N_22508,N_22063,N_22186);
and U22509 (N_22509,N_22150,N_22174);
or U22510 (N_22510,N_22382,N_22018);
or U22511 (N_22511,N_22487,N_22283);
nor U22512 (N_22512,N_22127,N_22253);
xor U22513 (N_22513,N_22029,N_22259);
or U22514 (N_22514,N_22019,N_22496);
and U22515 (N_22515,N_22248,N_22458);
xor U22516 (N_22516,N_22422,N_22234);
xnor U22517 (N_22517,N_22109,N_22434);
or U22518 (N_22518,N_22268,N_22057);
nand U22519 (N_22519,N_22444,N_22446);
and U22520 (N_22520,N_22328,N_22260);
nor U22521 (N_22521,N_22231,N_22373);
and U22522 (N_22522,N_22452,N_22372);
nor U22523 (N_22523,N_22129,N_22433);
nand U22524 (N_22524,N_22130,N_22359);
or U22525 (N_22525,N_22355,N_22192);
and U22526 (N_22526,N_22404,N_22197);
or U22527 (N_22527,N_22407,N_22347);
or U22528 (N_22528,N_22442,N_22403);
xor U22529 (N_22529,N_22478,N_22324);
and U22530 (N_22530,N_22074,N_22326);
xnor U22531 (N_22531,N_22295,N_22199);
nand U22532 (N_22532,N_22047,N_22131);
and U22533 (N_22533,N_22070,N_22432);
or U22534 (N_22534,N_22447,N_22170);
nand U22535 (N_22535,N_22336,N_22195);
and U22536 (N_22536,N_22204,N_22414);
xor U22537 (N_22537,N_22165,N_22482);
and U22538 (N_22538,N_22083,N_22286);
or U22539 (N_22539,N_22015,N_22448);
or U22540 (N_22540,N_22191,N_22292);
or U22541 (N_22541,N_22171,N_22217);
xnor U22542 (N_22542,N_22300,N_22315);
xnor U22543 (N_22543,N_22456,N_22340);
and U22544 (N_22544,N_22269,N_22306);
nor U22545 (N_22545,N_22335,N_22319);
nor U22546 (N_22546,N_22180,N_22416);
or U22547 (N_22547,N_22054,N_22285);
nand U22548 (N_22548,N_22467,N_22473);
nor U22549 (N_22549,N_22461,N_22046);
xnor U22550 (N_22550,N_22077,N_22214);
nand U22551 (N_22551,N_22005,N_22250);
and U22552 (N_22552,N_22360,N_22021);
and U22553 (N_22553,N_22158,N_22037);
xor U22554 (N_22554,N_22270,N_22481);
or U22555 (N_22555,N_22266,N_22242);
and U22556 (N_22556,N_22145,N_22321);
and U22557 (N_22557,N_22072,N_22495);
and U22558 (N_22558,N_22398,N_22026);
xnor U22559 (N_22559,N_22344,N_22227);
and U22560 (N_22560,N_22207,N_22469);
nand U22561 (N_22561,N_22133,N_22451);
and U22562 (N_22562,N_22025,N_22004);
nand U22563 (N_22563,N_22142,N_22154);
and U22564 (N_22564,N_22464,N_22423);
nor U22565 (N_22565,N_22203,N_22213);
and U22566 (N_22566,N_22140,N_22041);
nand U22567 (N_22567,N_22125,N_22272);
or U22568 (N_22568,N_22366,N_22421);
nor U22569 (N_22569,N_22163,N_22440);
and U22570 (N_22570,N_22086,N_22405);
xnor U22571 (N_22571,N_22287,N_22182);
or U22572 (N_22572,N_22238,N_22349);
or U22573 (N_22573,N_22271,N_22159);
nand U22574 (N_22574,N_22190,N_22153);
or U22575 (N_22575,N_22168,N_22483);
nor U22576 (N_22576,N_22104,N_22329);
or U22577 (N_22577,N_22024,N_22330);
xor U22578 (N_22578,N_22308,N_22480);
and U22579 (N_22579,N_22090,N_22362);
nand U22580 (N_22580,N_22311,N_22001);
nor U22581 (N_22581,N_22252,N_22060);
and U22582 (N_22582,N_22393,N_22208);
nor U22583 (N_22583,N_22491,N_22143);
nand U22584 (N_22584,N_22034,N_22113);
or U22585 (N_22585,N_22101,N_22371);
or U22586 (N_22586,N_22148,N_22465);
and U22587 (N_22587,N_22114,N_22323);
nand U22588 (N_22588,N_22115,N_22350);
or U22589 (N_22589,N_22460,N_22410);
nor U22590 (N_22590,N_22341,N_22144);
xor U22591 (N_22591,N_22424,N_22388);
or U22592 (N_22592,N_22202,N_22157);
xnor U22593 (N_22593,N_22188,N_22009);
xor U22594 (N_22594,N_22408,N_22139);
nand U22595 (N_22595,N_22392,N_22080);
nand U22596 (N_22596,N_22189,N_22036);
xor U22597 (N_22597,N_22304,N_22184);
and U22598 (N_22598,N_22098,N_22117);
nor U22599 (N_22599,N_22365,N_22084);
or U22600 (N_22600,N_22087,N_22399);
and U22601 (N_22601,N_22278,N_22235);
or U22602 (N_22602,N_22042,N_22097);
xor U22603 (N_22603,N_22417,N_22370);
and U22604 (N_22604,N_22386,N_22221);
nand U22605 (N_22605,N_22239,N_22152);
xnor U22606 (N_22606,N_22010,N_22337);
or U22607 (N_22607,N_22339,N_22438);
and U22608 (N_22608,N_22008,N_22274);
xnor U22609 (N_22609,N_22056,N_22120);
nand U22610 (N_22610,N_22012,N_22361);
nor U22611 (N_22611,N_22474,N_22147);
nand U22612 (N_22612,N_22497,N_22003);
or U22613 (N_22613,N_22176,N_22429);
xnor U22614 (N_22614,N_22291,N_22126);
xor U22615 (N_22615,N_22400,N_22185);
xnor U22616 (N_22616,N_22151,N_22119);
xor U22617 (N_22617,N_22251,N_22215);
nor U22618 (N_22618,N_22111,N_22236);
nand U22619 (N_22619,N_22394,N_22121);
or U22620 (N_22620,N_22052,N_22379);
nor U22621 (N_22621,N_22102,N_22210);
nor U22622 (N_22622,N_22256,N_22307);
or U22623 (N_22623,N_22418,N_22476);
or U22624 (N_22624,N_22387,N_22020);
nand U22625 (N_22625,N_22228,N_22419);
xor U22626 (N_22626,N_22293,N_22017);
xor U22627 (N_22627,N_22116,N_22000);
xnor U22628 (N_22628,N_22312,N_22345);
nor U22629 (N_22629,N_22156,N_22318);
xor U22630 (N_22630,N_22289,N_22230);
or U22631 (N_22631,N_22078,N_22411);
nor U22632 (N_22632,N_22205,N_22169);
nand U22633 (N_22633,N_22279,N_22310);
xnor U22634 (N_22634,N_22317,N_22406);
xnor U22635 (N_22635,N_22367,N_22402);
xor U22636 (N_22636,N_22472,N_22016);
xor U22637 (N_22637,N_22437,N_22178);
xor U22638 (N_22638,N_22164,N_22489);
nand U22639 (N_22639,N_22353,N_22455);
xnor U22640 (N_22640,N_22082,N_22209);
nor U22641 (N_22641,N_22059,N_22332);
or U22642 (N_22642,N_22490,N_22175);
or U22643 (N_22643,N_22294,N_22492);
nand U22644 (N_22644,N_22105,N_22346);
xor U22645 (N_22645,N_22284,N_22305);
xnor U22646 (N_22646,N_22343,N_22425);
nand U22647 (N_22647,N_22118,N_22463);
nand U22648 (N_22648,N_22241,N_22462);
or U22649 (N_22649,N_22194,N_22179);
nor U22650 (N_22650,N_22006,N_22378);
nor U22651 (N_22651,N_22031,N_22401);
or U22652 (N_22652,N_22369,N_22161);
xnor U22653 (N_22653,N_22089,N_22229);
nor U22654 (N_22654,N_22428,N_22439);
or U22655 (N_22655,N_22348,N_22479);
xnor U22656 (N_22656,N_22245,N_22223);
and U22657 (N_22657,N_22043,N_22391);
xor U22658 (N_22658,N_22368,N_22028);
nand U22659 (N_22659,N_22040,N_22053);
nand U22660 (N_22660,N_22389,N_22415);
or U22661 (N_22661,N_22263,N_22322);
nand U22662 (N_22662,N_22013,N_22273);
and U22663 (N_22663,N_22201,N_22342);
and U22664 (N_22664,N_22264,N_22333);
xnor U22665 (N_22665,N_22212,N_22298);
xnor U22666 (N_22666,N_22240,N_22062);
nand U22667 (N_22667,N_22233,N_22088);
or U22668 (N_22668,N_22218,N_22067);
nor U22669 (N_22669,N_22011,N_22309);
nor U22670 (N_22670,N_22093,N_22470);
xor U22671 (N_22671,N_22220,N_22107);
nor U22672 (N_22672,N_22222,N_22356);
xor U22673 (N_22673,N_22475,N_22280);
or U22674 (N_22674,N_22299,N_22498);
or U22675 (N_22675,N_22219,N_22039);
and U22676 (N_22676,N_22395,N_22160);
nand U22677 (N_22677,N_22354,N_22376);
nor U22678 (N_22678,N_22499,N_22316);
nor U22679 (N_22679,N_22380,N_22466);
and U22680 (N_22680,N_22051,N_22486);
xor U22681 (N_22681,N_22431,N_22196);
xnor U22682 (N_22682,N_22471,N_22358);
nand U22683 (N_22683,N_22172,N_22288);
nand U22684 (N_22684,N_22030,N_22296);
nand U22685 (N_22685,N_22488,N_22050);
xor U22686 (N_22686,N_22038,N_22162);
nor U22687 (N_22687,N_22064,N_22257);
nor U22688 (N_22688,N_22187,N_22033);
and U22689 (N_22689,N_22173,N_22331);
nor U22690 (N_22690,N_22124,N_22211);
xnor U22691 (N_22691,N_22110,N_22081);
nand U22692 (N_22692,N_22058,N_22413);
and U22693 (N_22693,N_22375,N_22225);
nand U22694 (N_22694,N_22352,N_22303);
or U22695 (N_22695,N_22224,N_22327);
or U22696 (N_22696,N_22325,N_22091);
nor U22697 (N_22697,N_22485,N_22155);
and U22698 (N_22698,N_22141,N_22079);
nand U22699 (N_22699,N_22146,N_22071);
nand U22700 (N_22700,N_22426,N_22181);
and U22701 (N_22701,N_22061,N_22237);
nor U22702 (N_22702,N_22138,N_22377);
nor U22703 (N_22703,N_22108,N_22149);
nor U22704 (N_22704,N_22255,N_22445);
nor U22705 (N_22705,N_22122,N_22277);
nor U22706 (N_22706,N_22249,N_22383);
and U22707 (N_22707,N_22099,N_22243);
or U22708 (N_22708,N_22226,N_22297);
or U22709 (N_22709,N_22281,N_22014);
or U22710 (N_22710,N_22106,N_22302);
or U22711 (N_22711,N_22459,N_22477);
nor U22712 (N_22712,N_22069,N_22258);
nand U22713 (N_22713,N_22254,N_22420);
or U22714 (N_22714,N_22384,N_22457);
nor U22715 (N_22715,N_22049,N_22301);
nor U22716 (N_22716,N_22048,N_22449);
and U22717 (N_22717,N_22128,N_22103);
and U22718 (N_22718,N_22320,N_22007);
and U22719 (N_22719,N_22137,N_22454);
nor U22720 (N_22720,N_22374,N_22044);
xnor U22721 (N_22721,N_22436,N_22435);
nor U22722 (N_22722,N_22123,N_22045);
nand U22723 (N_22723,N_22450,N_22100);
and U22724 (N_22724,N_22132,N_22412);
nor U22725 (N_22725,N_22055,N_22468);
and U22726 (N_22726,N_22261,N_22246);
nand U22727 (N_22727,N_22216,N_22232);
nor U22728 (N_22728,N_22167,N_22032);
xor U22729 (N_22729,N_22334,N_22135);
or U22730 (N_22730,N_22076,N_22183);
or U22731 (N_22731,N_22381,N_22493);
nor U22732 (N_22732,N_22314,N_22409);
xnor U22733 (N_22733,N_22275,N_22177);
xor U22734 (N_22734,N_22276,N_22096);
nor U22735 (N_22735,N_22265,N_22027);
or U22736 (N_22736,N_22244,N_22068);
nor U22737 (N_22737,N_22385,N_22338);
nand U22738 (N_22738,N_22166,N_22066);
nand U22739 (N_22739,N_22095,N_22085);
and U22740 (N_22740,N_22022,N_22002);
xor U22741 (N_22741,N_22136,N_22453);
nand U22742 (N_22742,N_22112,N_22247);
xnor U22743 (N_22743,N_22262,N_22035);
xnor U22744 (N_22744,N_22397,N_22494);
xnor U22745 (N_22745,N_22443,N_22427);
xor U22746 (N_22746,N_22267,N_22023);
and U22747 (N_22747,N_22193,N_22282);
nand U22748 (N_22748,N_22364,N_22134);
xnor U22749 (N_22749,N_22198,N_22073);
nand U22750 (N_22750,N_22319,N_22119);
nand U22751 (N_22751,N_22428,N_22238);
or U22752 (N_22752,N_22052,N_22130);
nor U22753 (N_22753,N_22051,N_22056);
nand U22754 (N_22754,N_22042,N_22279);
and U22755 (N_22755,N_22253,N_22055);
and U22756 (N_22756,N_22101,N_22399);
nor U22757 (N_22757,N_22497,N_22118);
or U22758 (N_22758,N_22437,N_22193);
xor U22759 (N_22759,N_22074,N_22105);
or U22760 (N_22760,N_22467,N_22012);
nor U22761 (N_22761,N_22230,N_22472);
nand U22762 (N_22762,N_22165,N_22057);
nor U22763 (N_22763,N_22024,N_22163);
and U22764 (N_22764,N_22004,N_22473);
nor U22765 (N_22765,N_22387,N_22198);
nand U22766 (N_22766,N_22362,N_22427);
xnor U22767 (N_22767,N_22301,N_22462);
nand U22768 (N_22768,N_22409,N_22068);
and U22769 (N_22769,N_22176,N_22264);
or U22770 (N_22770,N_22148,N_22379);
nand U22771 (N_22771,N_22362,N_22409);
nor U22772 (N_22772,N_22447,N_22125);
and U22773 (N_22773,N_22306,N_22427);
xor U22774 (N_22774,N_22422,N_22472);
nand U22775 (N_22775,N_22371,N_22389);
and U22776 (N_22776,N_22146,N_22022);
nand U22777 (N_22777,N_22163,N_22332);
xnor U22778 (N_22778,N_22384,N_22314);
nand U22779 (N_22779,N_22439,N_22393);
and U22780 (N_22780,N_22029,N_22221);
nor U22781 (N_22781,N_22199,N_22438);
nor U22782 (N_22782,N_22089,N_22473);
or U22783 (N_22783,N_22153,N_22287);
and U22784 (N_22784,N_22219,N_22397);
nand U22785 (N_22785,N_22497,N_22147);
or U22786 (N_22786,N_22481,N_22345);
nor U22787 (N_22787,N_22015,N_22119);
or U22788 (N_22788,N_22184,N_22129);
nor U22789 (N_22789,N_22045,N_22210);
nand U22790 (N_22790,N_22040,N_22101);
and U22791 (N_22791,N_22213,N_22429);
or U22792 (N_22792,N_22103,N_22097);
or U22793 (N_22793,N_22253,N_22479);
and U22794 (N_22794,N_22155,N_22286);
and U22795 (N_22795,N_22011,N_22047);
and U22796 (N_22796,N_22114,N_22248);
nor U22797 (N_22797,N_22016,N_22386);
or U22798 (N_22798,N_22373,N_22478);
and U22799 (N_22799,N_22432,N_22039);
xnor U22800 (N_22800,N_22017,N_22011);
nor U22801 (N_22801,N_22430,N_22498);
and U22802 (N_22802,N_22042,N_22273);
and U22803 (N_22803,N_22397,N_22435);
and U22804 (N_22804,N_22202,N_22152);
nand U22805 (N_22805,N_22279,N_22242);
nor U22806 (N_22806,N_22469,N_22010);
nand U22807 (N_22807,N_22176,N_22188);
and U22808 (N_22808,N_22314,N_22195);
and U22809 (N_22809,N_22343,N_22273);
nand U22810 (N_22810,N_22211,N_22257);
nand U22811 (N_22811,N_22107,N_22100);
nor U22812 (N_22812,N_22494,N_22357);
and U22813 (N_22813,N_22016,N_22175);
or U22814 (N_22814,N_22265,N_22131);
nand U22815 (N_22815,N_22370,N_22127);
and U22816 (N_22816,N_22100,N_22301);
xor U22817 (N_22817,N_22338,N_22227);
and U22818 (N_22818,N_22264,N_22349);
nand U22819 (N_22819,N_22199,N_22436);
nor U22820 (N_22820,N_22170,N_22209);
nand U22821 (N_22821,N_22481,N_22172);
and U22822 (N_22822,N_22228,N_22092);
or U22823 (N_22823,N_22148,N_22364);
xnor U22824 (N_22824,N_22308,N_22394);
and U22825 (N_22825,N_22136,N_22492);
or U22826 (N_22826,N_22263,N_22355);
nand U22827 (N_22827,N_22408,N_22387);
nor U22828 (N_22828,N_22013,N_22309);
nand U22829 (N_22829,N_22257,N_22011);
and U22830 (N_22830,N_22447,N_22117);
or U22831 (N_22831,N_22176,N_22295);
nor U22832 (N_22832,N_22459,N_22183);
or U22833 (N_22833,N_22385,N_22220);
and U22834 (N_22834,N_22478,N_22155);
and U22835 (N_22835,N_22477,N_22100);
xor U22836 (N_22836,N_22301,N_22477);
xnor U22837 (N_22837,N_22167,N_22172);
nand U22838 (N_22838,N_22006,N_22132);
nand U22839 (N_22839,N_22211,N_22096);
nand U22840 (N_22840,N_22033,N_22199);
and U22841 (N_22841,N_22213,N_22015);
nand U22842 (N_22842,N_22354,N_22198);
or U22843 (N_22843,N_22241,N_22036);
nor U22844 (N_22844,N_22176,N_22377);
and U22845 (N_22845,N_22429,N_22265);
or U22846 (N_22846,N_22208,N_22338);
or U22847 (N_22847,N_22076,N_22383);
xnor U22848 (N_22848,N_22041,N_22077);
or U22849 (N_22849,N_22245,N_22437);
or U22850 (N_22850,N_22433,N_22066);
or U22851 (N_22851,N_22331,N_22437);
xor U22852 (N_22852,N_22250,N_22075);
nor U22853 (N_22853,N_22244,N_22288);
and U22854 (N_22854,N_22428,N_22208);
and U22855 (N_22855,N_22405,N_22362);
xor U22856 (N_22856,N_22233,N_22373);
xor U22857 (N_22857,N_22187,N_22186);
xor U22858 (N_22858,N_22120,N_22199);
nand U22859 (N_22859,N_22280,N_22192);
nand U22860 (N_22860,N_22107,N_22067);
and U22861 (N_22861,N_22393,N_22341);
nand U22862 (N_22862,N_22325,N_22098);
and U22863 (N_22863,N_22400,N_22098);
or U22864 (N_22864,N_22243,N_22222);
nand U22865 (N_22865,N_22075,N_22234);
xnor U22866 (N_22866,N_22316,N_22191);
and U22867 (N_22867,N_22073,N_22333);
and U22868 (N_22868,N_22254,N_22432);
nor U22869 (N_22869,N_22357,N_22355);
nand U22870 (N_22870,N_22388,N_22116);
or U22871 (N_22871,N_22293,N_22196);
and U22872 (N_22872,N_22436,N_22414);
and U22873 (N_22873,N_22456,N_22236);
xnor U22874 (N_22874,N_22123,N_22070);
and U22875 (N_22875,N_22440,N_22353);
nor U22876 (N_22876,N_22224,N_22024);
nand U22877 (N_22877,N_22338,N_22062);
nor U22878 (N_22878,N_22401,N_22395);
or U22879 (N_22879,N_22178,N_22390);
nor U22880 (N_22880,N_22486,N_22481);
or U22881 (N_22881,N_22441,N_22017);
or U22882 (N_22882,N_22275,N_22270);
xor U22883 (N_22883,N_22250,N_22168);
and U22884 (N_22884,N_22416,N_22395);
and U22885 (N_22885,N_22276,N_22195);
nand U22886 (N_22886,N_22154,N_22029);
or U22887 (N_22887,N_22014,N_22145);
nor U22888 (N_22888,N_22364,N_22224);
xnor U22889 (N_22889,N_22470,N_22306);
nand U22890 (N_22890,N_22360,N_22427);
and U22891 (N_22891,N_22437,N_22356);
xnor U22892 (N_22892,N_22335,N_22032);
xnor U22893 (N_22893,N_22350,N_22059);
and U22894 (N_22894,N_22085,N_22405);
nand U22895 (N_22895,N_22208,N_22469);
nand U22896 (N_22896,N_22297,N_22468);
xnor U22897 (N_22897,N_22087,N_22030);
and U22898 (N_22898,N_22112,N_22065);
xor U22899 (N_22899,N_22254,N_22073);
and U22900 (N_22900,N_22398,N_22473);
xnor U22901 (N_22901,N_22277,N_22375);
nand U22902 (N_22902,N_22394,N_22061);
nand U22903 (N_22903,N_22447,N_22395);
nor U22904 (N_22904,N_22183,N_22475);
nand U22905 (N_22905,N_22053,N_22275);
and U22906 (N_22906,N_22105,N_22357);
nor U22907 (N_22907,N_22456,N_22227);
xnor U22908 (N_22908,N_22271,N_22251);
xnor U22909 (N_22909,N_22490,N_22057);
and U22910 (N_22910,N_22282,N_22355);
nand U22911 (N_22911,N_22212,N_22104);
xor U22912 (N_22912,N_22073,N_22457);
and U22913 (N_22913,N_22099,N_22049);
nand U22914 (N_22914,N_22303,N_22485);
nor U22915 (N_22915,N_22284,N_22143);
xnor U22916 (N_22916,N_22394,N_22379);
xor U22917 (N_22917,N_22153,N_22478);
or U22918 (N_22918,N_22133,N_22140);
or U22919 (N_22919,N_22328,N_22154);
nor U22920 (N_22920,N_22293,N_22446);
xor U22921 (N_22921,N_22265,N_22443);
nand U22922 (N_22922,N_22399,N_22223);
nor U22923 (N_22923,N_22494,N_22323);
nand U22924 (N_22924,N_22203,N_22124);
or U22925 (N_22925,N_22139,N_22364);
xnor U22926 (N_22926,N_22007,N_22262);
xor U22927 (N_22927,N_22265,N_22376);
and U22928 (N_22928,N_22155,N_22214);
and U22929 (N_22929,N_22179,N_22373);
or U22930 (N_22930,N_22221,N_22476);
or U22931 (N_22931,N_22167,N_22131);
and U22932 (N_22932,N_22378,N_22267);
xor U22933 (N_22933,N_22174,N_22396);
nor U22934 (N_22934,N_22428,N_22435);
and U22935 (N_22935,N_22056,N_22084);
or U22936 (N_22936,N_22205,N_22066);
and U22937 (N_22937,N_22041,N_22444);
xnor U22938 (N_22938,N_22490,N_22136);
nand U22939 (N_22939,N_22490,N_22273);
or U22940 (N_22940,N_22357,N_22169);
and U22941 (N_22941,N_22394,N_22270);
and U22942 (N_22942,N_22047,N_22362);
xor U22943 (N_22943,N_22281,N_22273);
xor U22944 (N_22944,N_22051,N_22215);
and U22945 (N_22945,N_22147,N_22235);
xnor U22946 (N_22946,N_22330,N_22013);
nor U22947 (N_22947,N_22178,N_22269);
and U22948 (N_22948,N_22102,N_22079);
xnor U22949 (N_22949,N_22017,N_22389);
xor U22950 (N_22950,N_22457,N_22094);
or U22951 (N_22951,N_22399,N_22332);
and U22952 (N_22952,N_22468,N_22205);
or U22953 (N_22953,N_22089,N_22254);
and U22954 (N_22954,N_22219,N_22438);
nand U22955 (N_22955,N_22016,N_22489);
nor U22956 (N_22956,N_22049,N_22242);
nand U22957 (N_22957,N_22428,N_22214);
xor U22958 (N_22958,N_22441,N_22440);
or U22959 (N_22959,N_22111,N_22089);
xor U22960 (N_22960,N_22310,N_22061);
or U22961 (N_22961,N_22379,N_22230);
and U22962 (N_22962,N_22270,N_22264);
and U22963 (N_22963,N_22059,N_22278);
xnor U22964 (N_22964,N_22145,N_22395);
or U22965 (N_22965,N_22237,N_22236);
nor U22966 (N_22966,N_22469,N_22319);
xor U22967 (N_22967,N_22197,N_22451);
xnor U22968 (N_22968,N_22425,N_22041);
and U22969 (N_22969,N_22432,N_22400);
and U22970 (N_22970,N_22001,N_22238);
nor U22971 (N_22971,N_22116,N_22234);
nand U22972 (N_22972,N_22311,N_22425);
xor U22973 (N_22973,N_22300,N_22075);
and U22974 (N_22974,N_22452,N_22022);
xor U22975 (N_22975,N_22422,N_22016);
nand U22976 (N_22976,N_22334,N_22439);
nand U22977 (N_22977,N_22158,N_22191);
nand U22978 (N_22978,N_22411,N_22434);
xnor U22979 (N_22979,N_22403,N_22099);
or U22980 (N_22980,N_22237,N_22257);
and U22981 (N_22981,N_22280,N_22277);
nand U22982 (N_22982,N_22285,N_22016);
or U22983 (N_22983,N_22176,N_22103);
nor U22984 (N_22984,N_22239,N_22412);
and U22985 (N_22985,N_22295,N_22073);
or U22986 (N_22986,N_22173,N_22119);
nor U22987 (N_22987,N_22119,N_22226);
nor U22988 (N_22988,N_22305,N_22118);
nand U22989 (N_22989,N_22312,N_22202);
or U22990 (N_22990,N_22295,N_22194);
xor U22991 (N_22991,N_22033,N_22381);
nand U22992 (N_22992,N_22478,N_22434);
nand U22993 (N_22993,N_22353,N_22492);
and U22994 (N_22994,N_22116,N_22481);
or U22995 (N_22995,N_22348,N_22044);
nor U22996 (N_22996,N_22188,N_22374);
and U22997 (N_22997,N_22366,N_22166);
nand U22998 (N_22998,N_22138,N_22109);
xnor U22999 (N_22999,N_22336,N_22439);
or U23000 (N_23000,N_22870,N_22788);
nor U23001 (N_23001,N_22934,N_22645);
or U23002 (N_23002,N_22927,N_22694);
or U23003 (N_23003,N_22749,N_22562);
nand U23004 (N_23004,N_22973,N_22970);
xnor U23005 (N_23005,N_22708,N_22631);
or U23006 (N_23006,N_22961,N_22637);
nor U23007 (N_23007,N_22818,N_22502);
nand U23008 (N_23008,N_22619,N_22628);
nor U23009 (N_23009,N_22550,N_22807);
xor U23010 (N_23010,N_22994,N_22744);
or U23011 (N_23011,N_22852,N_22872);
nor U23012 (N_23012,N_22922,N_22769);
nor U23013 (N_23013,N_22907,N_22564);
nand U23014 (N_23014,N_22699,N_22756);
or U23015 (N_23015,N_22767,N_22919);
nor U23016 (N_23016,N_22596,N_22660);
xor U23017 (N_23017,N_22544,N_22833);
nand U23018 (N_23018,N_22946,N_22542);
and U23019 (N_23019,N_22939,N_22691);
or U23020 (N_23020,N_22832,N_22516);
or U23021 (N_23021,N_22803,N_22674);
or U23022 (N_23022,N_22552,N_22588);
nand U23023 (N_23023,N_22871,N_22903);
or U23024 (N_23024,N_22639,N_22658);
nand U23025 (N_23025,N_22992,N_22742);
or U23026 (N_23026,N_22666,N_22524);
xor U23027 (N_23027,N_22776,N_22789);
or U23028 (N_23028,N_22740,N_22572);
xor U23029 (N_23029,N_22600,N_22513);
xnor U23030 (N_23030,N_22997,N_22986);
xnor U23031 (N_23031,N_22816,N_22711);
or U23032 (N_23032,N_22610,N_22838);
nand U23033 (N_23033,N_22830,N_22541);
nand U23034 (N_23034,N_22608,N_22553);
nor U23035 (N_23035,N_22535,N_22844);
or U23036 (N_23036,N_22831,N_22501);
xor U23037 (N_23037,N_22839,N_22665);
or U23038 (N_23038,N_22612,N_22792);
nand U23039 (N_23039,N_22827,N_22587);
or U23040 (N_23040,N_22508,N_22719);
or U23041 (N_23041,N_22787,N_22681);
nor U23042 (N_23042,N_22851,N_22885);
nand U23043 (N_23043,N_22644,N_22743);
or U23044 (N_23044,N_22837,N_22960);
or U23045 (N_23045,N_22825,N_22783);
nand U23046 (N_23046,N_22504,N_22935);
nand U23047 (N_23047,N_22741,N_22649);
nand U23048 (N_23048,N_22656,N_22866);
and U23049 (N_23049,N_22750,N_22623);
and U23050 (N_23050,N_22926,N_22714);
nand U23051 (N_23051,N_22657,N_22916);
and U23052 (N_23052,N_22696,N_22579);
or U23053 (N_23053,N_22597,N_22526);
or U23054 (N_23054,N_22875,N_22510);
xnor U23055 (N_23055,N_22966,N_22672);
nand U23056 (N_23056,N_22748,N_22736);
nor U23057 (N_23057,N_22778,N_22601);
nand U23058 (N_23058,N_22642,N_22991);
or U23059 (N_23059,N_22799,N_22954);
xor U23060 (N_23060,N_22758,N_22928);
xnor U23061 (N_23061,N_22898,N_22828);
nand U23062 (N_23062,N_22841,N_22785);
or U23063 (N_23063,N_22591,N_22503);
or U23064 (N_23064,N_22583,N_22824);
nand U23065 (N_23065,N_22958,N_22811);
xnor U23066 (N_23066,N_22584,N_22709);
or U23067 (N_23067,N_22899,N_22774);
nand U23068 (N_23068,N_22707,N_22655);
nand U23069 (N_23069,N_22805,N_22646);
or U23070 (N_23070,N_22540,N_22904);
nor U23071 (N_23071,N_22887,N_22638);
nor U23072 (N_23072,N_22772,N_22545);
or U23073 (N_23073,N_22560,N_22819);
nor U23074 (N_23074,N_22940,N_22693);
nand U23075 (N_23075,N_22618,N_22640);
nor U23076 (N_23076,N_22864,N_22555);
nand U23077 (N_23077,N_22975,N_22520);
nand U23078 (N_23078,N_22697,N_22942);
nor U23079 (N_23079,N_22995,N_22802);
nand U23080 (N_23080,N_22775,N_22845);
nor U23081 (N_23081,N_22514,N_22941);
and U23082 (N_23082,N_22617,N_22790);
and U23083 (N_23083,N_22575,N_22533);
nor U23084 (N_23084,N_22668,N_22724);
and U23085 (N_23085,N_22972,N_22568);
nor U23086 (N_23086,N_22880,N_22673);
and U23087 (N_23087,N_22554,N_22761);
nor U23088 (N_23088,N_22705,N_22985);
xor U23089 (N_23089,N_22959,N_22721);
and U23090 (N_23090,N_22894,N_22730);
or U23091 (N_23091,N_22725,N_22731);
or U23092 (N_23092,N_22846,N_22506);
nor U23093 (N_23093,N_22951,N_22733);
nand U23094 (N_23094,N_22949,N_22808);
and U23095 (N_23095,N_22678,N_22703);
nor U23096 (N_23096,N_22902,N_22988);
nand U23097 (N_23097,N_22770,N_22868);
nor U23098 (N_23098,N_22751,N_22990);
and U23099 (N_23099,N_22918,N_22569);
nor U23100 (N_23100,N_22627,N_22576);
nand U23101 (N_23101,N_22689,N_22710);
xor U23102 (N_23102,N_22848,N_22684);
xor U23103 (N_23103,N_22909,N_22823);
xor U23104 (N_23104,N_22635,N_22806);
nor U23105 (N_23105,N_22862,N_22857);
nand U23106 (N_23106,N_22747,N_22980);
nand U23107 (N_23107,N_22944,N_22661);
nand U23108 (N_23108,N_22680,N_22715);
nor U23109 (N_23109,N_22523,N_22936);
and U23110 (N_23110,N_22893,N_22891);
or U23111 (N_23111,N_22763,N_22931);
xnor U23112 (N_23112,N_22701,N_22984);
and U23113 (N_23113,N_22964,N_22755);
xnor U23114 (N_23114,N_22873,N_22614);
and U23115 (N_23115,N_22539,N_22534);
and U23116 (N_23116,N_22571,N_22509);
nand U23117 (N_23117,N_22804,N_22598);
nand U23118 (N_23118,N_22877,N_22669);
nor U23119 (N_23119,N_22888,N_22515);
xor U23120 (N_23120,N_22739,N_22956);
nor U23121 (N_23121,N_22822,N_22521);
or U23122 (N_23122,N_22971,N_22621);
xor U23123 (N_23123,N_22757,N_22625);
nor U23124 (N_23124,N_22798,N_22817);
nor U23125 (N_23125,N_22737,N_22826);
or U23126 (N_23126,N_22895,N_22633);
nor U23127 (N_23127,N_22842,N_22905);
or U23128 (N_23128,N_22974,N_22603);
xnor U23129 (N_23129,N_22505,N_22652);
and U23130 (N_23130,N_22727,N_22595);
or U23131 (N_23131,N_22734,N_22843);
xnor U23132 (N_23132,N_22653,N_22886);
nand U23133 (N_23133,N_22728,N_22722);
or U23134 (N_23134,N_22917,N_22948);
nor U23135 (N_23135,N_22592,N_22593);
xor U23136 (N_23136,N_22930,N_22518);
xor U23137 (N_23137,N_22695,N_22978);
nor U23138 (N_23138,N_22671,N_22813);
nand U23139 (N_23139,N_22522,N_22585);
xor U23140 (N_23140,N_22746,N_22908);
nand U23141 (N_23141,N_22996,N_22795);
xor U23142 (N_23142,N_22869,N_22878);
nand U23143 (N_23143,N_22754,N_22613);
or U23144 (N_23144,N_22892,N_22912);
nand U23145 (N_23145,N_22753,N_22624);
xnor U23146 (N_23146,N_22945,N_22605);
or U23147 (N_23147,N_22791,N_22796);
nand U23148 (N_23148,N_22559,N_22543);
xor U23149 (N_23149,N_22814,N_22626);
xor U23150 (N_23150,N_22764,N_22580);
nor U23151 (N_23151,N_22692,N_22987);
nor U23152 (N_23152,N_22538,N_22937);
nand U23153 (N_23153,N_22519,N_22781);
nand U23154 (N_23154,N_22924,N_22570);
xnor U23155 (N_23155,N_22670,N_22664);
and U23156 (N_23156,N_22729,N_22890);
or U23157 (N_23157,N_22698,N_22933);
xnor U23158 (N_23158,N_22556,N_22815);
nor U23159 (N_23159,N_22820,N_22723);
nand U23160 (N_23160,N_22738,N_22551);
nand U23161 (N_23161,N_22547,N_22929);
nor U23162 (N_23162,N_22998,N_22906);
or U23163 (N_23163,N_22879,N_22786);
or U23164 (N_23164,N_22915,N_22910);
and U23165 (N_23165,N_22977,N_22889);
xor U23166 (N_23166,N_22962,N_22760);
or U23167 (N_23167,N_22511,N_22812);
and U23168 (N_23168,N_22525,N_22901);
nor U23169 (N_23169,N_22616,N_22943);
and U23170 (N_23170,N_22683,N_22688);
nor U23171 (N_23171,N_22810,N_22607);
nor U23172 (N_23172,N_22745,N_22548);
or U23173 (N_23173,N_22881,N_22549);
nor U23174 (N_23174,N_22883,N_22911);
nor U23175 (N_23175,N_22993,N_22953);
nand U23176 (N_23176,N_22771,N_22999);
nand U23177 (N_23177,N_22780,N_22573);
and U23178 (N_23178,N_22854,N_22720);
or U23179 (N_23179,N_22967,N_22766);
and U23180 (N_23180,N_22950,N_22858);
nor U23181 (N_23181,N_22923,N_22957);
and U23182 (N_23182,N_22622,N_22793);
and U23183 (N_23183,N_22982,N_22606);
and U23184 (N_23184,N_22650,N_22836);
or U23185 (N_23185,N_22884,N_22677);
xnor U23186 (N_23186,N_22863,N_22938);
or U23187 (N_23187,N_22609,N_22630);
nand U23188 (N_23188,N_22682,N_22578);
nor U23189 (N_23189,N_22762,N_22955);
nand U23190 (N_23190,N_22641,N_22735);
xor U23191 (N_23191,N_22849,N_22563);
xnor U23192 (N_23192,N_22794,N_22537);
or U23193 (N_23193,N_22651,N_22590);
xor U23194 (N_23194,N_22732,N_22856);
and U23195 (N_23195,N_22586,N_22861);
nand U23196 (N_23196,N_22685,N_22874);
nor U23197 (N_23197,N_22782,N_22765);
and U23198 (N_23198,N_22768,N_22500);
or U23199 (N_23199,N_22702,N_22557);
nor U23200 (N_23200,N_22835,N_22679);
or U23201 (N_23201,N_22700,N_22663);
or U23202 (N_23202,N_22636,N_22779);
nor U23203 (N_23203,N_22865,N_22920);
nand U23204 (N_23204,N_22634,N_22647);
or U23205 (N_23205,N_22876,N_22752);
or U23206 (N_23206,N_22611,N_22643);
nor U23207 (N_23207,N_22981,N_22581);
nor U23208 (N_23208,N_22594,N_22914);
or U23209 (N_23209,N_22577,N_22687);
nand U23210 (N_23210,N_22706,N_22952);
or U23211 (N_23211,N_22821,N_22712);
and U23212 (N_23212,N_22654,N_22983);
nand U23213 (N_23213,N_22602,N_22897);
and U23214 (N_23214,N_22773,N_22599);
xor U23215 (N_23215,N_22718,N_22530);
and U23216 (N_23216,N_22932,N_22859);
nand U23217 (N_23217,N_22512,N_22528);
nand U23218 (N_23218,N_22784,N_22809);
nor U23219 (N_23219,N_22531,N_22561);
or U23220 (N_23220,N_22834,N_22604);
nor U23221 (N_23221,N_22853,N_22759);
nand U23222 (N_23222,N_22867,N_22558);
xnor U23223 (N_23223,N_22567,N_22662);
xnor U23224 (N_23224,N_22517,N_22726);
nor U23225 (N_23225,N_22921,N_22797);
and U23226 (N_23226,N_22847,N_22913);
nor U23227 (N_23227,N_22690,N_22589);
or U23228 (N_23228,N_22565,N_22716);
nor U23229 (N_23229,N_22800,N_22829);
nor U23230 (N_23230,N_22546,N_22667);
and U23231 (N_23231,N_22704,N_22675);
nor U23232 (N_23232,N_22686,N_22629);
xor U23233 (N_23233,N_22777,N_22566);
nand U23234 (N_23234,N_22850,N_22963);
or U23235 (N_23235,N_22620,N_22968);
and U23236 (N_23236,N_22860,N_22574);
or U23237 (N_23237,N_22840,N_22713);
nor U23238 (N_23238,N_22615,N_22965);
nor U23239 (N_23239,N_22969,N_22979);
nor U23240 (N_23240,N_22582,N_22900);
nand U23241 (N_23241,N_22717,N_22801);
xor U23242 (N_23242,N_22896,N_22989);
nor U23243 (N_23243,N_22529,N_22532);
xnor U23244 (N_23244,N_22882,N_22855);
xor U23245 (N_23245,N_22976,N_22527);
and U23246 (N_23246,N_22648,N_22676);
or U23247 (N_23247,N_22947,N_22632);
or U23248 (N_23248,N_22925,N_22659);
nor U23249 (N_23249,N_22536,N_22507);
xor U23250 (N_23250,N_22581,N_22752);
nand U23251 (N_23251,N_22853,N_22597);
nor U23252 (N_23252,N_22862,N_22593);
and U23253 (N_23253,N_22865,N_22941);
nand U23254 (N_23254,N_22577,N_22653);
nand U23255 (N_23255,N_22975,N_22854);
and U23256 (N_23256,N_22534,N_22605);
nand U23257 (N_23257,N_22803,N_22691);
or U23258 (N_23258,N_22544,N_22567);
xor U23259 (N_23259,N_22951,N_22668);
nor U23260 (N_23260,N_22870,N_22686);
and U23261 (N_23261,N_22572,N_22663);
or U23262 (N_23262,N_22540,N_22791);
xnor U23263 (N_23263,N_22610,N_22913);
and U23264 (N_23264,N_22930,N_22941);
nand U23265 (N_23265,N_22547,N_22920);
nor U23266 (N_23266,N_22663,N_22931);
xnor U23267 (N_23267,N_22820,N_22642);
nand U23268 (N_23268,N_22919,N_22763);
or U23269 (N_23269,N_22684,N_22886);
and U23270 (N_23270,N_22805,N_22990);
xor U23271 (N_23271,N_22714,N_22923);
nand U23272 (N_23272,N_22939,N_22961);
nand U23273 (N_23273,N_22530,N_22539);
and U23274 (N_23274,N_22997,N_22860);
nor U23275 (N_23275,N_22509,N_22816);
nor U23276 (N_23276,N_22628,N_22945);
and U23277 (N_23277,N_22740,N_22652);
nand U23278 (N_23278,N_22746,N_22735);
nand U23279 (N_23279,N_22798,N_22543);
nor U23280 (N_23280,N_22695,N_22771);
xor U23281 (N_23281,N_22900,N_22522);
nor U23282 (N_23282,N_22533,N_22586);
or U23283 (N_23283,N_22972,N_22902);
nor U23284 (N_23284,N_22958,N_22920);
nor U23285 (N_23285,N_22659,N_22642);
xnor U23286 (N_23286,N_22910,N_22899);
and U23287 (N_23287,N_22623,N_22737);
or U23288 (N_23288,N_22921,N_22635);
xnor U23289 (N_23289,N_22919,N_22805);
xnor U23290 (N_23290,N_22712,N_22556);
and U23291 (N_23291,N_22502,N_22549);
xor U23292 (N_23292,N_22571,N_22942);
or U23293 (N_23293,N_22709,N_22618);
and U23294 (N_23294,N_22719,N_22684);
xor U23295 (N_23295,N_22794,N_22912);
nor U23296 (N_23296,N_22515,N_22747);
nor U23297 (N_23297,N_22968,N_22678);
xnor U23298 (N_23298,N_22961,N_22874);
nor U23299 (N_23299,N_22531,N_22619);
nor U23300 (N_23300,N_22612,N_22922);
and U23301 (N_23301,N_22655,N_22548);
nand U23302 (N_23302,N_22817,N_22587);
and U23303 (N_23303,N_22771,N_22654);
or U23304 (N_23304,N_22664,N_22831);
or U23305 (N_23305,N_22776,N_22507);
nor U23306 (N_23306,N_22712,N_22825);
and U23307 (N_23307,N_22805,N_22707);
nor U23308 (N_23308,N_22775,N_22638);
nand U23309 (N_23309,N_22945,N_22753);
nor U23310 (N_23310,N_22642,N_22583);
nand U23311 (N_23311,N_22870,N_22751);
nand U23312 (N_23312,N_22760,N_22781);
nand U23313 (N_23313,N_22870,N_22712);
and U23314 (N_23314,N_22911,N_22788);
and U23315 (N_23315,N_22847,N_22724);
or U23316 (N_23316,N_22733,N_22510);
nand U23317 (N_23317,N_22672,N_22500);
xnor U23318 (N_23318,N_22604,N_22777);
and U23319 (N_23319,N_22526,N_22585);
or U23320 (N_23320,N_22883,N_22923);
nand U23321 (N_23321,N_22675,N_22835);
and U23322 (N_23322,N_22634,N_22767);
nand U23323 (N_23323,N_22683,N_22873);
nand U23324 (N_23324,N_22980,N_22535);
and U23325 (N_23325,N_22810,N_22681);
nand U23326 (N_23326,N_22582,N_22937);
or U23327 (N_23327,N_22594,N_22932);
and U23328 (N_23328,N_22719,N_22611);
and U23329 (N_23329,N_22753,N_22517);
or U23330 (N_23330,N_22854,N_22766);
xnor U23331 (N_23331,N_22897,N_22974);
nor U23332 (N_23332,N_22967,N_22730);
or U23333 (N_23333,N_22604,N_22900);
or U23334 (N_23334,N_22811,N_22598);
and U23335 (N_23335,N_22759,N_22606);
or U23336 (N_23336,N_22660,N_22970);
or U23337 (N_23337,N_22788,N_22871);
and U23338 (N_23338,N_22575,N_22792);
nand U23339 (N_23339,N_22769,N_22544);
or U23340 (N_23340,N_22570,N_22845);
or U23341 (N_23341,N_22875,N_22980);
or U23342 (N_23342,N_22567,N_22910);
or U23343 (N_23343,N_22701,N_22683);
xor U23344 (N_23344,N_22604,N_22591);
nor U23345 (N_23345,N_22997,N_22927);
and U23346 (N_23346,N_22545,N_22541);
xor U23347 (N_23347,N_22672,N_22725);
nand U23348 (N_23348,N_22600,N_22642);
nor U23349 (N_23349,N_22755,N_22722);
or U23350 (N_23350,N_22622,N_22672);
and U23351 (N_23351,N_22694,N_22545);
nand U23352 (N_23352,N_22813,N_22643);
nand U23353 (N_23353,N_22606,N_22717);
nand U23354 (N_23354,N_22808,N_22543);
nor U23355 (N_23355,N_22563,N_22512);
nor U23356 (N_23356,N_22796,N_22651);
nand U23357 (N_23357,N_22711,N_22994);
or U23358 (N_23358,N_22688,N_22818);
or U23359 (N_23359,N_22751,N_22888);
nor U23360 (N_23360,N_22574,N_22993);
nor U23361 (N_23361,N_22813,N_22828);
and U23362 (N_23362,N_22745,N_22929);
or U23363 (N_23363,N_22561,N_22876);
nand U23364 (N_23364,N_22735,N_22829);
xnor U23365 (N_23365,N_22837,N_22710);
and U23366 (N_23366,N_22586,N_22976);
nand U23367 (N_23367,N_22600,N_22855);
nand U23368 (N_23368,N_22968,N_22528);
nor U23369 (N_23369,N_22976,N_22599);
nand U23370 (N_23370,N_22766,N_22975);
or U23371 (N_23371,N_22751,N_22713);
nand U23372 (N_23372,N_22883,N_22549);
nor U23373 (N_23373,N_22754,N_22709);
nand U23374 (N_23374,N_22631,N_22676);
nand U23375 (N_23375,N_22888,N_22860);
or U23376 (N_23376,N_22556,N_22659);
nor U23377 (N_23377,N_22773,N_22978);
nand U23378 (N_23378,N_22503,N_22752);
or U23379 (N_23379,N_22540,N_22655);
and U23380 (N_23380,N_22578,N_22997);
nand U23381 (N_23381,N_22985,N_22584);
and U23382 (N_23382,N_22516,N_22959);
nand U23383 (N_23383,N_22740,N_22566);
nor U23384 (N_23384,N_22876,N_22662);
nor U23385 (N_23385,N_22671,N_22683);
or U23386 (N_23386,N_22750,N_22817);
nand U23387 (N_23387,N_22743,N_22709);
and U23388 (N_23388,N_22952,N_22872);
xnor U23389 (N_23389,N_22638,N_22809);
nand U23390 (N_23390,N_22993,N_22591);
nand U23391 (N_23391,N_22569,N_22931);
or U23392 (N_23392,N_22833,N_22639);
or U23393 (N_23393,N_22639,N_22533);
xor U23394 (N_23394,N_22645,N_22538);
xnor U23395 (N_23395,N_22958,N_22624);
and U23396 (N_23396,N_22633,N_22914);
xor U23397 (N_23397,N_22752,N_22544);
or U23398 (N_23398,N_22851,N_22913);
nor U23399 (N_23399,N_22670,N_22651);
and U23400 (N_23400,N_22925,N_22516);
nand U23401 (N_23401,N_22702,N_22865);
nand U23402 (N_23402,N_22889,N_22749);
and U23403 (N_23403,N_22890,N_22553);
or U23404 (N_23404,N_22930,N_22566);
or U23405 (N_23405,N_22959,N_22676);
and U23406 (N_23406,N_22565,N_22560);
and U23407 (N_23407,N_22658,N_22729);
and U23408 (N_23408,N_22785,N_22965);
and U23409 (N_23409,N_22578,N_22663);
nor U23410 (N_23410,N_22957,N_22668);
xnor U23411 (N_23411,N_22865,N_22759);
xnor U23412 (N_23412,N_22983,N_22959);
nor U23413 (N_23413,N_22512,N_22715);
and U23414 (N_23414,N_22997,N_22869);
nand U23415 (N_23415,N_22554,N_22895);
nor U23416 (N_23416,N_22569,N_22750);
xor U23417 (N_23417,N_22573,N_22504);
xnor U23418 (N_23418,N_22516,N_22979);
or U23419 (N_23419,N_22738,N_22596);
or U23420 (N_23420,N_22815,N_22614);
nor U23421 (N_23421,N_22787,N_22894);
nor U23422 (N_23422,N_22643,N_22947);
or U23423 (N_23423,N_22529,N_22967);
nand U23424 (N_23424,N_22502,N_22593);
xor U23425 (N_23425,N_22980,N_22810);
or U23426 (N_23426,N_22996,N_22610);
and U23427 (N_23427,N_22773,N_22705);
nor U23428 (N_23428,N_22635,N_22984);
xor U23429 (N_23429,N_22940,N_22525);
xor U23430 (N_23430,N_22605,N_22559);
nand U23431 (N_23431,N_22947,N_22675);
or U23432 (N_23432,N_22734,N_22559);
nand U23433 (N_23433,N_22925,N_22976);
nand U23434 (N_23434,N_22568,N_22621);
xor U23435 (N_23435,N_22643,N_22566);
xnor U23436 (N_23436,N_22650,N_22507);
or U23437 (N_23437,N_22600,N_22802);
and U23438 (N_23438,N_22661,N_22771);
nor U23439 (N_23439,N_22591,N_22647);
nor U23440 (N_23440,N_22684,N_22987);
nor U23441 (N_23441,N_22756,N_22559);
and U23442 (N_23442,N_22741,N_22622);
and U23443 (N_23443,N_22752,N_22819);
xor U23444 (N_23444,N_22900,N_22873);
nand U23445 (N_23445,N_22753,N_22503);
and U23446 (N_23446,N_22880,N_22993);
xnor U23447 (N_23447,N_22887,N_22865);
nand U23448 (N_23448,N_22541,N_22647);
nor U23449 (N_23449,N_22785,N_22507);
nor U23450 (N_23450,N_22530,N_22647);
and U23451 (N_23451,N_22832,N_22505);
and U23452 (N_23452,N_22833,N_22991);
nor U23453 (N_23453,N_22525,N_22797);
and U23454 (N_23454,N_22567,N_22559);
xor U23455 (N_23455,N_22826,N_22526);
xnor U23456 (N_23456,N_22552,N_22762);
nor U23457 (N_23457,N_22944,N_22805);
nand U23458 (N_23458,N_22881,N_22824);
or U23459 (N_23459,N_22689,N_22736);
nor U23460 (N_23460,N_22731,N_22594);
nand U23461 (N_23461,N_22813,N_22706);
nor U23462 (N_23462,N_22936,N_22838);
and U23463 (N_23463,N_22658,N_22825);
or U23464 (N_23464,N_22997,N_22629);
nand U23465 (N_23465,N_22990,N_22852);
nand U23466 (N_23466,N_22844,N_22746);
xor U23467 (N_23467,N_22886,N_22698);
and U23468 (N_23468,N_22723,N_22824);
xnor U23469 (N_23469,N_22857,N_22569);
or U23470 (N_23470,N_22861,N_22628);
nor U23471 (N_23471,N_22900,N_22842);
or U23472 (N_23472,N_22624,N_22822);
nand U23473 (N_23473,N_22684,N_22888);
nand U23474 (N_23474,N_22671,N_22655);
or U23475 (N_23475,N_22972,N_22866);
nor U23476 (N_23476,N_22853,N_22885);
and U23477 (N_23477,N_22939,N_22710);
or U23478 (N_23478,N_22977,N_22981);
nor U23479 (N_23479,N_22862,N_22902);
nand U23480 (N_23480,N_22580,N_22817);
or U23481 (N_23481,N_22643,N_22720);
and U23482 (N_23482,N_22964,N_22983);
nor U23483 (N_23483,N_22586,N_22535);
or U23484 (N_23484,N_22639,N_22788);
nand U23485 (N_23485,N_22849,N_22719);
and U23486 (N_23486,N_22625,N_22722);
xor U23487 (N_23487,N_22799,N_22965);
nand U23488 (N_23488,N_22909,N_22570);
xnor U23489 (N_23489,N_22749,N_22540);
and U23490 (N_23490,N_22893,N_22521);
nor U23491 (N_23491,N_22578,N_22535);
and U23492 (N_23492,N_22647,N_22747);
xor U23493 (N_23493,N_22611,N_22860);
xnor U23494 (N_23494,N_22718,N_22624);
nor U23495 (N_23495,N_22665,N_22836);
nand U23496 (N_23496,N_22720,N_22609);
and U23497 (N_23497,N_22839,N_22518);
or U23498 (N_23498,N_22805,N_22994);
xor U23499 (N_23499,N_22594,N_22921);
and U23500 (N_23500,N_23268,N_23282);
or U23501 (N_23501,N_23201,N_23060);
nor U23502 (N_23502,N_23102,N_23182);
xnor U23503 (N_23503,N_23464,N_23442);
and U23504 (N_23504,N_23259,N_23325);
nand U23505 (N_23505,N_23183,N_23237);
or U23506 (N_23506,N_23430,N_23370);
nand U23507 (N_23507,N_23067,N_23088);
and U23508 (N_23508,N_23189,N_23145);
nand U23509 (N_23509,N_23125,N_23106);
or U23510 (N_23510,N_23200,N_23034);
xnor U23511 (N_23511,N_23077,N_23167);
nand U23512 (N_23512,N_23441,N_23160);
xnor U23513 (N_23513,N_23405,N_23298);
xor U23514 (N_23514,N_23236,N_23131);
nor U23515 (N_23515,N_23101,N_23312);
nand U23516 (N_23516,N_23350,N_23238);
xnor U23517 (N_23517,N_23164,N_23072);
nand U23518 (N_23518,N_23388,N_23460);
nor U23519 (N_23519,N_23425,N_23346);
nor U23520 (N_23520,N_23038,N_23165);
nand U23521 (N_23521,N_23279,N_23477);
or U23522 (N_23522,N_23311,N_23111);
xor U23523 (N_23523,N_23066,N_23152);
or U23524 (N_23524,N_23428,N_23222);
and U23525 (N_23525,N_23175,N_23407);
and U23526 (N_23526,N_23071,N_23126);
and U23527 (N_23527,N_23026,N_23417);
xnor U23528 (N_23528,N_23296,N_23031);
and U23529 (N_23529,N_23456,N_23098);
nor U23530 (N_23530,N_23452,N_23399);
xor U23531 (N_23531,N_23377,N_23040);
or U23532 (N_23532,N_23321,N_23406);
or U23533 (N_23533,N_23448,N_23254);
and U23534 (N_23534,N_23342,N_23157);
nor U23535 (N_23535,N_23260,N_23062);
nor U23536 (N_23536,N_23378,N_23356);
nand U23537 (N_23537,N_23443,N_23246);
nor U23538 (N_23538,N_23241,N_23371);
nor U23539 (N_23539,N_23057,N_23382);
or U23540 (N_23540,N_23297,N_23394);
nor U23541 (N_23541,N_23334,N_23366);
nor U23542 (N_23542,N_23413,N_23333);
xor U23543 (N_23543,N_23480,N_23411);
and U23544 (N_23544,N_23251,N_23243);
or U23545 (N_23545,N_23095,N_23229);
and U23546 (N_23546,N_23043,N_23089);
or U23547 (N_23547,N_23014,N_23016);
or U23548 (N_23548,N_23093,N_23338);
or U23549 (N_23549,N_23384,N_23219);
nand U23550 (N_23550,N_23252,N_23248);
nand U23551 (N_23551,N_23113,N_23196);
nor U23552 (N_23552,N_23436,N_23262);
xor U23553 (N_23553,N_23439,N_23315);
nor U23554 (N_23554,N_23212,N_23054);
nand U23555 (N_23555,N_23288,N_23128);
nor U23556 (N_23556,N_23115,N_23341);
nor U23557 (N_23557,N_23397,N_23322);
nor U23558 (N_23558,N_23037,N_23472);
nand U23559 (N_23559,N_23231,N_23427);
nor U23560 (N_23560,N_23142,N_23324);
xnor U23561 (N_23561,N_23150,N_23310);
xnor U23562 (N_23562,N_23025,N_23061);
and U23563 (N_23563,N_23485,N_23454);
xor U23564 (N_23564,N_23203,N_23151);
xnor U23565 (N_23565,N_23110,N_23055);
nand U23566 (N_23566,N_23455,N_23301);
xnor U23567 (N_23567,N_23249,N_23008);
or U23568 (N_23568,N_23476,N_23440);
nor U23569 (N_23569,N_23206,N_23159);
nand U23570 (N_23570,N_23372,N_23258);
or U23571 (N_23571,N_23363,N_23392);
and U23572 (N_23572,N_23359,N_23148);
nor U23573 (N_23573,N_23261,N_23404);
or U23574 (N_23574,N_23463,N_23272);
and U23575 (N_23575,N_23239,N_23070);
nand U23576 (N_23576,N_23433,N_23122);
and U23577 (N_23577,N_23143,N_23467);
nand U23578 (N_23578,N_23327,N_23461);
xor U23579 (N_23579,N_23494,N_23051);
nand U23580 (N_23580,N_23094,N_23220);
nor U23581 (N_23581,N_23158,N_23217);
and U23582 (N_23582,N_23257,N_23186);
and U23583 (N_23583,N_23487,N_23007);
nor U23584 (N_23584,N_23317,N_23409);
or U23585 (N_23585,N_23275,N_23303);
nor U23586 (N_23586,N_23277,N_23387);
nor U23587 (N_23587,N_23457,N_23365);
nand U23588 (N_23588,N_23465,N_23451);
xnor U23589 (N_23589,N_23116,N_23453);
and U23590 (N_23590,N_23065,N_23123);
or U23591 (N_23591,N_23245,N_23347);
xor U23592 (N_23592,N_23422,N_23362);
nand U23593 (N_23593,N_23000,N_23117);
nor U23594 (N_23594,N_23028,N_23069);
nand U23595 (N_23595,N_23432,N_23408);
nor U23596 (N_23596,N_23191,N_23267);
or U23597 (N_23597,N_23355,N_23400);
xor U23598 (N_23598,N_23082,N_23018);
and U23599 (N_23599,N_23002,N_23187);
nor U23600 (N_23600,N_23364,N_23214);
and U23601 (N_23601,N_23172,N_23368);
or U23602 (N_23602,N_23289,N_23367);
and U23603 (N_23603,N_23184,N_23147);
nor U23604 (N_23604,N_23188,N_23009);
xor U23605 (N_23605,N_23444,N_23438);
and U23606 (N_23606,N_23027,N_23195);
nor U23607 (N_23607,N_23086,N_23316);
and U23608 (N_23608,N_23129,N_23011);
nor U23609 (N_23609,N_23483,N_23389);
and U23610 (N_23610,N_23287,N_23215);
or U23611 (N_23611,N_23486,N_23264);
nand U23612 (N_23612,N_23462,N_23358);
xnor U23613 (N_23613,N_23210,N_23041);
xnor U23614 (N_23614,N_23280,N_23181);
and U23615 (N_23615,N_23420,N_23308);
xnor U23616 (N_23616,N_23180,N_23473);
or U23617 (N_23617,N_23445,N_23266);
or U23618 (N_23618,N_23235,N_23360);
and U23619 (N_23619,N_23058,N_23391);
nor U23620 (N_23620,N_23403,N_23044);
nand U23621 (N_23621,N_23369,N_23216);
and U23622 (N_23622,N_23307,N_23474);
xor U23623 (N_23623,N_23499,N_23139);
or U23624 (N_23624,N_23240,N_23396);
nor U23625 (N_23625,N_23039,N_23010);
nand U23626 (N_23626,N_23305,N_23414);
and U23627 (N_23627,N_23218,N_23050);
nand U23628 (N_23628,N_23336,N_23109);
xnor U23629 (N_23629,N_23173,N_23424);
nor U23630 (N_23630,N_23450,N_23381);
nand U23631 (N_23631,N_23100,N_23170);
xor U23632 (N_23632,N_23169,N_23437);
nor U23633 (N_23633,N_23299,N_23097);
nand U23634 (N_23634,N_23198,N_23314);
nand U23635 (N_23635,N_23223,N_23144);
and U23636 (N_23636,N_23036,N_23353);
nand U23637 (N_23637,N_23003,N_23030);
nand U23638 (N_23638,N_23373,N_23045);
nor U23639 (N_23639,N_23205,N_23114);
xnor U23640 (N_23640,N_23337,N_23343);
or U23641 (N_23641,N_23162,N_23185);
and U23642 (N_23642,N_23357,N_23471);
or U23643 (N_23643,N_23335,N_23118);
and U23644 (N_23644,N_23177,N_23402);
nand U23645 (N_23645,N_23211,N_23049);
nor U23646 (N_23646,N_23421,N_23291);
nand U23647 (N_23647,N_23141,N_23386);
nor U23648 (N_23648,N_23283,N_23458);
nand U23649 (N_23649,N_23419,N_23361);
nand U23650 (N_23650,N_23163,N_23161);
nor U23651 (N_23651,N_23006,N_23328);
nor U23652 (N_23652,N_23330,N_23395);
nor U23653 (N_23653,N_23446,N_23478);
or U23654 (N_23654,N_23119,N_23285);
xnor U23655 (N_23655,N_23107,N_23146);
or U23656 (N_23656,N_23329,N_23265);
nor U23657 (N_23657,N_23412,N_23497);
nand U23658 (N_23658,N_23326,N_23103);
xor U23659 (N_23659,N_23074,N_23004);
nand U23660 (N_23660,N_23256,N_23416);
or U23661 (N_23661,N_23208,N_23304);
nor U23662 (N_23662,N_23276,N_23390);
nor U23663 (N_23663,N_23255,N_23022);
or U23664 (N_23664,N_23012,N_23140);
nor U23665 (N_23665,N_23383,N_23380);
nor U23666 (N_23666,N_23230,N_23490);
xor U23667 (N_23667,N_23434,N_23349);
nand U23668 (N_23668,N_23099,N_23024);
nand U23669 (N_23669,N_23495,N_23019);
xor U23670 (N_23670,N_23052,N_23112);
or U23671 (N_23671,N_23127,N_23344);
xor U23672 (N_23672,N_23470,N_23042);
xnor U23673 (N_23673,N_23475,N_23084);
or U23674 (N_23674,N_23253,N_23247);
nor U23675 (N_23675,N_23429,N_23447);
nand U23676 (N_23676,N_23137,N_23068);
nand U23677 (N_23677,N_23393,N_23401);
or U23678 (N_23678,N_23435,N_23059);
or U23679 (N_23679,N_23138,N_23385);
nor U23680 (N_23680,N_23023,N_23064);
xnor U23681 (N_23681,N_23281,N_23076);
or U23682 (N_23682,N_23313,N_23479);
and U23683 (N_23683,N_23080,N_23284);
or U23684 (N_23684,N_23302,N_23331);
nor U23685 (N_23685,N_23431,N_23375);
or U23686 (N_23686,N_23073,N_23192);
xnor U23687 (N_23687,N_23482,N_23199);
nor U23688 (N_23688,N_23228,N_23046);
nand U23689 (N_23689,N_23345,N_23202);
or U23690 (N_23690,N_23318,N_23354);
or U23691 (N_23691,N_23493,N_23130);
or U23692 (N_23692,N_23092,N_23295);
and U23693 (N_23693,N_23048,N_23290);
nand U23694 (N_23694,N_23244,N_23468);
or U23695 (N_23695,N_23017,N_23149);
xor U23696 (N_23696,N_23204,N_23029);
nand U23697 (N_23697,N_23032,N_23124);
nor U23698 (N_23698,N_23174,N_23286);
nand U23699 (N_23699,N_23085,N_23020);
nor U23700 (N_23700,N_23178,N_23156);
nand U23701 (N_23701,N_23221,N_23423);
or U23702 (N_23702,N_23083,N_23047);
nor U23703 (N_23703,N_23090,N_23108);
and U23704 (N_23704,N_23352,N_23379);
nand U23705 (N_23705,N_23348,N_23035);
and U23706 (N_23706,N_23306,N_23274);
xor U23707 (N_23707,N_23376,N_23001);
xor U23708 (N_23708,N_23227,N_23294);
nor U23709 (N_23709,N_23418,N_23469);
nor U23710 (N_23710,N_23056,N_23233);
nand U23711 (N_23711,N_23120,N_23075);
or U23712 (N_23712,N_23351,N_23155);
or U23713 (N_23713,N_23320,N_23096);
and U23714 (N_23714,N_23105,N_23053);
nor U23715 (N_23715,N_23087,N_23153);
or U23716 (N_23716,N_23340,N_23484);
and U23717 (N_23717,N_23207,N_23224);
xnor U23718 (N_23718,N_23278,N_23300);
xor U23719 (N_23719,N_23190,N_23234);
nor U23720 (N_23720,N_23021,N_23063);
xor U23721 (N_23721,N_23332,N_23496);
or U23722 (N_23722,N_23339,N_23489);
and U23723 (N_23723,N_23133,N_23193);
or U23724 (N_23724,N_23498,N_23374);
or U23725 (N_23725,N_23319,N_23213);
or U23726 (N_23726,N_23079,N_23481);
and U23727 (N_23727,N_23132,N_23225);
and U23728 (N_23728,N_23121,N_23271);
nand U23729 (N_23729,N_23104,N_23323);
nor U23730 (N_23730,N_23242,N_23488);
nor U23731 (N_23731,N_23449,N_23263);
nor U23732 (N_23732,N_23171,N_23309);
or U23733 (N_23733,N_23209,N_23292);
nor U23734 (N_23734,N_23154,N_23293);
and U23735 (N_23735,N_23078,N_23273);
nand U23736 (N_23736,N_23270,N_23081);
or U23737 (N_23737,N_23091,N_23250);
nor U23738 (N_23738,N_23179,N_23013);
or U23739 (N_23739,N_23459,N_23426);
xnor U23740 (N_23740,N_23166,N_23194);
nor U23741 (N_23741,N_23136,N_23466);
and U23742 (N_23742,N_23226,N_23491);
nand U23743 (N_23743,N_23176,N_23232);
nand U23744 (N_23744,N_23005,N_23134);
xnor U23745 (N_23745,N_23269,N_23492);
or U23746 (N_23746,N_23015,N_23033);
xor U23747 (N_23747,N_23168,N_23410);
and U23748 (N_23748,N_23415,N_23197);
xor U23749 (N_23749,N_23135,N_23398);
or U23750 (N_23750,N_23091,N_23386);
and U23751 (N_23751,N_23226,N_23052);
or U23752 (N_23752,N_23460,N_23374);
nor U23753 (N_23753,N_23436,N_23429);
nand U23754 (N_23754,N_23442,N_23348);
nor U23755 (N_23755,N_23463,N_23353);
and U23756 (N_23756,N_23492,N_23249);
or U23757 (N_23757,N_23386,N_23050);
xor U23758 (N_23758,N_23456,N_23160);
xor U23759 (N_23759,N_23221,N_23368);
or U23760 (N_23760,N_23392,N_23354);
and U23761 (N_23761,N_23243,N_23405);
or U23762 (N_23762,N_23150,N_23176);
and U23763 (N_23763,N_23257,N_23234);
and U23764 (N_23764,N_23433,N_23231);
xor U23765 (N_23765,N_23274,N_23286);
and U23766 (N_23766,N_23491,N_23238);
and U23767 (N_23767,N_23318,N_23092);
nand U23768 (N_23768,N_23431,N_23031);
and U23769 (N_23769,N_23145,N_23004);
and U23770 (N_23770,N_23498,N_23373);
nand U23771 (N_23771,N_23274,N_23392);
nand U23772 (N_23772,N_23293,N_23217);
and U23773 (N_23773,N_23294,N_23263);
or U23774 (N_23774,N_23405,N_23380);
or U23775 (N_23775,N_23320,N_23495);
nand U23776 (N_23776,N_23400,N_23166);
and U23777 (N_23777,N_23359,N_23100);
nor U23778 (N_23778,N_23316,N_23067);
and U23779 (N_23779,N_23389,N_23178);
nand U23780 (N_23780,N_23408,N_23365);
nor U23781 (N_23781,N_23027,N_23441);
xor U23782 (N_23782,N_23111,N_23334);
or U23783 (N_23783,N_23339,N_23165);
nor U23784 (N_23784,N_23200,N_23152);
xnor U23785 (N_23785,N_23430,N_23396);
nor U23786 (N_23786,N_23174,N_23343);
nand U23787 (N_23787,N_23381,N_23326);
or U23788 (N_23788,N_23307,N_23410);
xnor U23789 (N_23789,N_23247,N_23334);
or U23790 (N_23790,N_23261,N_23019);
xnor U23791 (N_23791,N_23291,N_23134);
and U23792 (N_23792,N_23188,N_23317);
nand U23793 (N_23793,N_23068,N_23231);
and U23794 (N_23794,N_23162,N_23368);
xor U23795 (N_23795,N_23093,N_23117);
or U23796 (N_23796,N_23319,N_23464);
nor U23797 (N_23797,N_23427,N_23340);
and U23798 (N_23798,N_23069,N_23228);
nand U23799 (N_23799,N_23326,N_23362);
and U23800 (N_23800,N_23448,N_23333);
and U23801 (N_23801,N_23197,N_23202);
nand U23802 (N_23802,N_23063,N_23054);
or U23803 (N_23803,N_23110,N_23270);
nand U23804 (N_23804,N_23431,N_23058);
and U23805 (N_23805,N_23121,N_23295);
and U23806 (N_23806,N_23148,N_23275);
and U23807 (N_23807,N_23065,N_23358);
or U23808 (N_23808,N_23496,N_23477);
xor U23809 (N_23809,N_23260,N_23420);
and U23810 (N_23810,N_23121,N_23013);
nand U23811 (N_23811,N_23235,N_23349);
xor U23812 (N_23812,N_23218,N_23343);
xor U23813 (N_23813,N_23045,N_23250);
nor U23814 (N_23814,N_23438,N_23499);
xor U23815 (N_23815,N_23391,N_23067);
or U23816 (N_23816,N_23154,N_23374);
or U23817 (N_23817,N_23202,N_23337);
xor U23818 (N_23818,N_23219,N_23388);
nor U23819 (N_23819,N_23414,N_23464);
xnor U23820 (N_23820,N_23010,N_23452);
nor U23821 (N_23821,N_23326,N_23150);
nor U23822 (N_23822,N_23380,N_23213);
nand U23823 (N_23823,N_23080,N_23373);
nand U23824 (N_23824,N_23353,N_23019);
or U23825 (N_23825,N_23401,N_23426);
xor U23826 (N_23826,N_23164,N_23338);
nor U23827 (N_23827,N_23339,N_23352);
nor U23828 (N_23828,N_23249,N_23212);
nor U23829 (N_23829,N_23248,N_23475);
xor U23830 (N_23830,N_23211,N_23479);
xnor U23831 (N_23831,N_23380,N_23165);
nor U23832 (N_23832,N_23047,N_23162);
or U23833 (N_23833,N_23233,N_23373);
nor U23834 (N_23834,N_23013,N_23364);
nand U23835 (N_23835,N_23398,N_23122);
nand U23836 (N_23836,N_23411,N_23118);
or U23837 (N_23837,N_23176,N_23470);
or U23838 (N_23838,N_23390,N_23200);
or U23839 (N_23839,N_23424,N_23405);
or U23840 (N_23840,N_23122,N_23070);
nor U23841 (N_23841,N_23415,N_23382);
xnor U23842 (N_23842,N_23099,N_23110);
nand U23843 (N_23843,N_23203,N_23210);
xor U23844 (N_23844,N_23256,N_23358);
xnor U23845 (N_23845,N_23452,N_23233);
xor U23846 (N_23846,N_23064,N_23419);
or U23847 (N_23847,N_23141,N_23055);
nand U23848 (N_23848,N_23284,N_23380);
and U23849 (N_23849,N_23190,N_23104);
and U23850 (N_23850,N_23244,N_23243);
and U23851 (N_23851,N_23333,N_23163);
nand U23852 (N_23852,N_23186,N_23419);
xor U23853 (N_23853,N_23276,N_23163);
and U23854 (N_23854,N_23474,N_23402);
xor U23855 (N_23855,N_23275,N_23408);
and U23856 (N_23856,N_23469,N_23386);
xnor U23857 (N_23857,N_23119,N_23358);
xnor U23858 (N_23858,N_23347,N_23259);
or U23859 (N_23859,N_23436,N_23164);
and U23860 (N_23860,N_23357,N_23044);
and U23861 (N_23861,N_23225,N_23254);
nor U23862 (N_23862,N_23140,N_23402);
nor U23863 (N_23863,N_23104,N_23211);
nand U23864 (N_23864,N_23098,N_23110);
nor U23865 (N_23865,N_23370,N_23004);
nor U23866 (N_23866,N_23478,N_23483);
nand U23867 (N_23867,N_23399,N_23285);
xnor U23868 (N_23868,N_23024,N_23031);
nor U23869 (N_23869,N_23188,N_23224);
and U23870 (N_23870,N_23121,N_23079);
and U23871 (N_23871,N_23298,N_23052);
and U23872 (N_23872,N_23139,N_23470);
nor U23873 (N_23873,N_23255,N_23262);
nand U23874 (N_23874,N_23090,N_23244);
nor U23875 (N_23875,N_23398,N_23276);
and U23876 (N_23876,N_23149,N_23459);
nand U23877 (N_23877,N_23323,N_23006);
nand U23878 (N_23878,N_23123,N_23351);
and U23879 (N_23879,N_23336,N_23258);
and U23880 (N_23880,N_23032,N_23272);
xnor U23881 (N_23881,N_23177,N_23213);
nor U23882 (N_23882,N_23429,N_23012);
xor U23883 (N_23883,N_23075,N_23295);
or U23884 (N_23884,N_23483,N_23408);
nor U23885 (N_23885,N_23160,N_23245);
and U23886 (N_23886,N_23185,N_23458);
or U23887 (N_23887,N_23454,N_23071);
xor U23888 (N_23888,N_23149,N_23101);
or U23889 (N_23889,N_23130,N_23123);
xnor U23890 (N_23890,N_23385,N_23063);
and U23891 (N_23891,N_23228,N_23019);
nand U23892 (N_23892,N_23444,N_23334);
and U23893 (N_23893,N_23005,N_23251);
or U23894 (N_23894,N_23370,N_23036);
nor U23895 (N_23895,N_23018,N_23090);
xor U23896 (N_23896,N_23298,N_23373);
or U23897 (N_23897,N_23173,N_23019);
nand U23898 (N_23898,N_23359,N_23062);
and U23899 (N_23899,N_23237,N_23165);
nand U23900 (N_23900,N_23220,N_23293);
and U23901 (N_23901,N_23429,N_23420);
and U23902 (N_23902,N_23329,N_23079);
xor U23903 (N_23903,N_23304,N_23486);
or U23904 (N_23904,N_23476,N_23333);
xor U23905 (N_23905,N_23112,N_23465);
nor U23906 (N_23906,N_23225,N_23239);
xor U23907 (N_23907,N_23172,N_23339);
or U23908 (N_23908,N_23009,N_23135);
nor U23909 (N_23909,N_23478,N_23467);
or U23910 (N_23910,N_23339,N_23364);
nor U23911 (N_23911,N_23473,N_23348);
xor U23912 (N_23912,N_23098,N_23164);
or U23913 (N_23913,N_23188,N_23155);
and U23914 (N_23914,N_23366,N_23229);
xor U23915 (N_23915,N_23247,N_23259);
nor U23916 (N_23916,N_23449,N_23218);
xnor U23917 (N_23917,N_23065,N_23284);
or U23918 (N_23918,N_23441,N_23011);
nand U23919 (N_23919,N_23340,N_23047);
xor U23920 (N_23920,N_23229,N_23161);
nor U23921 (N_23921,N_23045,N_23469);
and U23922 (N_23922,N_23231,N_23025);
nand U23923 (N_23923,N_23317,N_23303);
and U23924 (N_23924,N_23270,N_23210);
or U23925 (N_23925,N_23191,N_23011);
nand U23926 (N_23926,N_23157,N_23189);
xnor U23927 (N_23927,N_23208,N_23172);
xor U23928 (N_23928,N_23346,N_23416);
and U23929 (N_23929,N_23212,N_23348);
nand U23930 (N_23930,N_23040,N_23372);
nand U23931 (N_23931,N_23249,N_23400);
nor U23932 (N_23932,N_23172,N_23422);
nand U23933 (N_23933,N_23064,N_23099);
nand U23934 (N_23934,N_23209,N_23169);
nor U23935 (N_23935,N_23220,N_23281);
xnor U23936 (N_23936,N_23435,N_23041);
or U23937 (N_23937,N_23149,N_23391);
nor U23938 (N_23938,N_23177,N_23362);
and U23939 (N_23939,N_23351,N_23431);
nand U23940 (N_23940,N_23394,N_23030);
xnor U23941 (N_23941,N_23319,N_23070);
xnor U23942 (N_23942,N_23287,N_23471);
nor U23943 (N_23943,N_23263,N_23497);
or U23944 (N_23944,N_23078,N_23359);
and U23945 (N_23945,N_23248,N_23040);
and U23946 (N_23946,N_23441,N_23470);
and U23947 (N_23947,N_23371,N_23007);
nor U23948 (N_23948,N_23499,N_23095);
nor U23949 (N_23949,N_23474,N_23163);
xnor U23950 (N_23950,N_23150,N_23076);
or U23951 (N_23951,N_23118,N_23228);
or U23952 (N_23952,N_23205,N_23217);
nor U23953 (N_23953,N_23065,N_23302);
nand U23954 (N_23954,N_23449,N_23017);
nor U23955 (N_23955,N_23059,N_23461);
or U23956 (N_23956,N_23317,N_23098);
xnor U23957 (N_23957,N_23296,N_23218);
xnor U23958 (N_23958,N_23218,N_23240);
and U23959 (N_23959,N_23164,N_23396);
nor U23960 (N_23960,N_23292,N_23114);
or U23961 (N_23961,N_23043,N_23031);
nand U23962 (N_23962,N_23040,N_23011);
or U23963 (N_23963,N_23329,N_23400);
nor U23964 (N_23964,N_23258,N_23251);
nor U23965 (N_23965,N_23006,N_23367);
nor U23966 (N_23966,N_23130,N_23435);
nor U23967 (N_23967,N_23306,N_23468);
nor U23968 (N_23968,N_23453,N_23459);
nor U23969 (N_23969,N_23397,N_23257);
nor U23970 (N_23970,N_23457,N_23035);
or U23971 (N_23971,N_23024,N_23222);
or U23972 (N_23972,N_23151,N_23142);
or U23973 (N_23973,N_23123,N_23275);
and U23974 (N_23974,N_23282,N_23182);
or U23975 (N_23975,N_23153,N_23053);
xnor U23976 (N_23976,N_23408,N_23498);
nand U23977 (N_23977,N_23352,N_23161);
xnor U23978 (N_23978,N_23399,N_23466);
nand U23979 (N_23979,N_23148,N_23110);
nor U23980 (N_23980,N_23302,N_23329);
or U23981 (N_23981,N_23335,N_23483);
and U23982 (N_23982,N_23244,N_23348);
nor U23983 (N_23983,N_23025,N_23139);
and U23984 (N_23984,N_23113,N_23109);
and U23985 (N_23985,N_23182,N_23076);
nand U23986 (N_23986,N_23445,N_23468);
nor U23987 (N_23987,N_23238,N_23475);
nand U23988 (N_23988,N_23474,N_23147);
and U23989 (N_23989,N_23298,N_23499);
and U23990 (N_23990,N_23410,N_23339);
or U23991 (N_23991,N_23112,N_23244);
or U23992 (N_23992,N_23340,N_23222);
or U23993 (N_23993,N_23451,N_23051);
or U23994 (N_23994,N_23354,N_23221);
nand U23995 (N_23995,N_23265,N_23482);
xor U23996 (N_23996,N_23269,N_23158);
xnor U23997 (N_23997,N_23001,N_23053);
nor U23998 (N_23998,N_23342,N_23316);
and U23999 (N_23999,N_23425,N_23301);
and U24000 (N_24000,N_23621,N_23807);
and U24001 (N_24001,N_23801,N_23638);
xor U24002 (N_24002,N_23646,N_23853);
xnor U24003 (N_24003,N_23787,N_23924);
xnor U24004 (N_24004,N_23572,N_23984);
xnor U24005 (N_24005,N_23901,N_23673);
nor U24006 (N_24006,N_23722,N_23653);
xor U24007 (N_24007,N_23980,N_23618);
nand U24008 (N_24008,N_23566,N_23660);
nand U24009 (N_24009,N_23734,N_23711);
nor U24010 (N_24010,N_23727,N_23669);
nand U24011 (N_24011,N_23602,N_23592);
or U24012 (N_24012,N_23679,N_23874);
nand U24013 (N_24013,N_23622,N_23681);
xnor U24014 (N_24014,N_23830,N_23696);
and U24015 (N_24015,N_23538,N_23838);
and U24016 (N_24016,N_23887,N_23897);
and U24017 (N_24017,N_23839,N_23820);
nor U24018 (N_24018,N_23857,N_23970);
nor U24019 (N_24019,N_23541,N_23919);
nand U24020 (N_24020,N_23684,N_23790);
or U24021 (N_24021,N_23674,N_23561);
nor U24022 (N_24022,N_23615,N_23862);
nor U24023 (N_24023,N_23803,N_23524);
nor U24024 (N_24024,N_23872,N_23962);
and U24025 (N_24025,N_23658,N_23979);
xnor U24026 (N_24026,N_23912,N_23822);
and U24027 (N_24027,N_23706,N_23865);
xor U24028 (N_24028,N_23695,N_23636);
xor U24029 (N_24029,N_23714,N_23604);
nor U24030 (N_24030,N_23914,N_23998);
nor U24031 (N_24031,N_23767,N_23743);
xor U24032 (N_24032,N_23725,N_23516);
nor U24033 (N_24033,N_23890,N_23596);
or U24034 (N_24034,N_23805,N_23661);
or U24035 (N_24035,N_23859,N_23748);
nand U24036 (N_24036,N_23502,N_23546);
nand U24037 (N_24037,N_23554,N_23573);
xnor U24038 (N_24038,N_23772,N_23928);
nor U24039 (N_24039,N_23730,N_23578);
xnor U24040 (N_24040,N_23946,N_23882);
nor U24041 (N_24041,N_23631,N_23733);
or U24042 (N_24042,N_23855,N_23771);
and U24043 (N_24043,N_23826,N_23934);
nand U24044 (N_24044,N_23782,N_23676);
nand U24045 (N_24045,N_23655,N_23964);
xor U24046 (N_24046,N_23837,N_23833);
or U24047 (N_24047,N_23836,N_23993);
xor U24048 (N_24048,N_23535,N_23614);
and U24049 (N_24049,N_23528,N_23827);
and U24050 (N_24050,N_23880,N_23608);
xnor U24051 (N_24051,N_23779,N_23944);
nor U24052 (N_24052,N_23851,N_23824);
and U24053 (N_24053,N_23550,N_23823);
nor U24054 (N_24054,N_23774,N_23809);
xnor U24055 (N_24055,N_23759,N_23635);
or U24056 (N_24056,N_23918,N_23935);
nor U24057 (N_24057,N_23847,N_23559);
and U24058 (N_24058,N_23586,N_23870);
xor U24059 (N_24059,N_23972,N_23783);
xor U24060 (N_24060,N_23540,N_23991);
or U24061 (N_24061,N_23907,N_23581);
and U24062 (N_24062,N_23504,N_23973);
and U24063 (N_24063,N_23902,N_23739);
nand U24064 (N_24064,N_23850,N_23988);
and U24065 (N_24065,N_23828,N_23603);
nand U24066 (N_24066,N_23571,N_23761);
nor U24067 (N_24067,N_23742,N_23952);
or U24068 (N_24068,N_23915,N_23968);
xnor U24069 (N_24069,N_23560,N_23792);
nand U24070 (N_24070,N_23536,N_23808);
xor U24071 (N_24071,N_23613,N_23508);
xor U24072 (N_24072,N_23665,N_23594);
xor U24073 (N_24073,N_23549,N_23703);
xnor U24074 (N_24074,N_23651,N_23694);
nand U24075 (N_24075,N_23738,N_23818);
xnor U24076 (N_24076,N_23943,N_23930);
or U24077 (N_24077,N_23806,N_23831);
nand U24078 (N_24078,N_23909,N_23843);
and U24079 (N_24079,N_23926,N_23815);
and U24080 (N_24080,N_23707,N_23971);
nand U24081 (N_24081,N_23987,N_23704);
and U24082 (N_24082,N_23526,N_23639);
and U24083 (N_24083,N_23741,N_23657);
xnor U24084 (N_24084,N_23796,N_23705);
nor U24085 (N_24085,N_23520,N_23537);
xnor U24086 (N_24086,N_23768,N_23766);
or U24087 (N_24087,N_23922,N_23997);
or U24088 (N_24088,N_23953,N_23794);
or U24089 (N_24089,N_23558,N_23640);
nand U24090 (N_24090,N_23903,N_23648);
xnor U24091 (N_24091,N_23925,N_23607);
and U24092 (N_24092,N_23686,N_23555);
nand U24093 (N_24093,N_23976,N_23598);
or U24094 (N_24094,N_23529,N_23793);
nand U24095 (N_24095,N_23515,N_23533);
nand U24096 (N_24096,N_23810,N_23729);
nand U24097 (N_24097,N_23990,N_23948);
nand U24098 (N_24098,N_23710,N_23947);
nor U24099 (N_24099,N_23685,N_23749);
xor U24100 (N_24100,N_23860,N_23888);
nor U24101 (N_24101,N_23652,N_23835);
nand U24102 (N_24102,N_23552,N_23786);
xor U24103 (N_24103,N_23871,N_23940);
or U24104 (N_24104,N_23737,N_23643);
or U24105 (N_24105,N_23965,N_23906);
nor U24106 (N_24106,N_23518,N_23975);
or U24107 (N_24107,N_23553,N_23777);
nor U24108 (N_24108,N_23866,N_23778);
nand U24109 (N_24109,N_23556,N_23671);
nand U24110 (N_24110,N_23693,N_23933);
or U24111 (N_24111,N_23878,N_23617);
nand U24112 (N_24112,N_23910,N_23637);
and U24113 (N_24113,N_23886,N_23644);
nand U24114 (N_24114,N_23896,N_23688);
xnor U24115 (N_24115,N_23534,N_23736);
nand U24116 (N_24116,N_23977,N_23717);
nand U24117 (N_24117,N_23869,N_23905);
nand U24118 (N_24118,N_23626,N_23891);
and U24119 (N_24119,N_23666,N_23601);
nand U24120 (N_24120,N_23858,N_23583);
and U24121 (N_24121,N_23620,N_23591);
or U24122 (N_24122,N_23670,N_23687);
nor U24123 (N_24123,N_23625,N_23623);
or U24124 (N_24124,N_23799,N_23931);
nand U24125 (N_24125,N_23868,N_23776);
nor U24126 (N_24126,N_23856,N_23764);
nand U24127 (N_24127,N_23852,N_23957);
xor U24128 (N_24128,N_23894,N_23753);
and U24129 (N_24129,N_23612,N_23732);
or U24130 (N_24130,N_23849,N_23718);
or U24131 (N_24131,N_23762,N_23974);
nand U24132 (N_24132,N_23932,N_23692);
and U24133 (N_24133,N_23819,N_23900);
nor U24134 (N_24134,N_23610,N_23570);
xnor U24135 (N_24135,N_23750,N_23611);
or U24136 (N_24136,N_23923,N_23659);
nand U24137 (N_24137,N_23527,N_23756);
nor U24138 (N_24138,N_23927,N_23667);
or U24139 (N_24139,N_23512,N_23689);
and U24140 (N_24140,N_23992,N_23713);
nand U24141 (N_24141,N_23816,N_23950);
nand U24142 (N_24142,N_23951,N_23548);
and U24143 (N_24143,N_23963,N_23812);
and U24144 (N_24144,N_23978,N_23728);
or U24145 (N_24145,N_23642,N_23916);
xor U24146 (N_24146,N_23697,N_23875);
or U24147 (N_24147,N_23629,N_23547);
and U24148 (N_24148,N_23510,N_23788);
and U24149 (N_24149,N_23543,N_23641);
nand U24150 (N_24150,N_23588,N_23532);
nor U24151 (N_24151,N_23752,N_23513);
and U24152 (N_24152,N_23505,N_23966);
xnor U24153 (N_24153,N_23584,N_23832);
and U24154 (N_24154,N_23892,N_23797);
and U24155 (N_24155,N_23921,N_23745);
nand U24156 (N_24156,N_23758,N_23521);
and U24157 (N_24157,N_23740,N_23677);
xnor U24158 (N_24158,N_23577,N_23829);
nand U24159 (N_24159,N_23895,N_23506);
nor U24160 (N_24160,N_23723,N_23715);
nor U24161 (N_24161,N_23763,N_23746);
and U24162 (N_24162,N_23985,N_23785);
nand U24163 (N_24163,N_23811,N_23877);
and U24164 (N_24164,N_23814,N_23841);
nor U24165 (N_24165,N_23663,N_23600);
and U24166 (N_24166,N_23873,N_23568);
xnor U24167 (N_24167,N_23567,N_23595);
xnor U24168 (N_24168,N_23509,N_23904);
nand U24169 (N_24169,N_23760,N_23709);
and U24170 (N_24170,N_23662,N_23589);
nor U24171 (N_24171,N_23956,N_23773);
nor U24172 (N_24172,N_23969,N_23542);
nand U24173 (N_24173,N_23525,N_23634);
xnor U24174 (N_24174,N_23755,N_23958);
xnor U24175 (N_24175,N_23562,N_23645);
xor U24176 (N_24176,N_23569,N_23938);
xnor U24177 (N_24177,N_23698,N_23883);
xnor U24178 (N_24178,N_23557,N_23587);
and U24179 (N_24179,N_23654,N_23664);
or U24180 (N_24180,N_23744,N_23937);
and U24181 (N_24181,N_23675,N_23593);
and U24182 (N_24182,N_23996,N_23702);
nand U24183 (N_24183,N_23920,N_23507);
or U24184 (N_24184,N_23834,N_23981);
and U24185 (N_24185,N_23983,N_23582);
or U24186 (N_24186,N_23735,N_23544);
or U24187 (N_24187,N_23795,N_23563);
xnor U24188 (N_24188,N_23845,N_23649);
and U24189 (N_24189,N_23501,N_23798);
nor U24190 (N_24190,N_23913,N_23959);
xnor U24191 (N_24191,N_23726,N_23672);
nand U24192 (N_24192,N_23719,N_23564);
and U24193 (N_24193,N_23628,N_23627);
nor U24194 (N_24194,N_23917,N_23580);
nand U24195 (N_24195,N_23844,N_23911);
nor U24196 (N_24196,N_23678,N_23683);
xor U24197 (N_24197,N_23864,N_23656);
xor U24198 (N_24198,N_23551,N_23701);
or U24199 (N_24199,N_23967,N_23863);
or U24200 (N_24200,N_23889,N_23605);
xor U24201 (N_24201,N_23765,N_23939);
xor U24202 (N_24202,N_23942,N_23775);
or U24203 (N_24203,N_23590,N_23517);
nand U24204 (N_24204,N_23708,N_23780);
nand U24205 (N_24205,N_23757,N_23961);
or U24206 (N_24206,N_23840,N_23690);
xnor U24207 (N_24207,N_23754,N_23781);
nor U24208 (N_24208,N_23522,N_23721);
or U24209 (N_24209,N_23955,N_23879);
nand U24210 (N_24210,N_23539,N_23867);
nand U24211 (N_24211,N_23576,N_23802);
or U24212 (N_24212,N_23954,N_23929);
or U24213 (N_24213,N_23500,N_23881);
and U24214 (N_24214,N_23530,N_23784);
and U24215 (N_24215,N_23609,N_23519);
xor U24216 (N_24216,N_23770,N_23616);
xnor U24217 (N_24217,N_23747,N_23574);
xor U24218 (N_24218,N_23791,N_23960);
and U24219 (N_24219,N_23597,N_23650);
or U24220 (N_24220,N_23619,N_23712);
nor U24221 (N_24221,N_23825,N_23821);
nor U24222 (N_24222,N_23514,N_23579);
nand U24223 (N_24223,N_23885,N_23699);
nor U24224 (N_24224,N_23769,N_23884);
nand U24225 (N_24225,N_23630,N_23949);
and U24226 (N_24226,N_23800,N_23632);
nand U24227 (N_24227,N_23982,N_23813);
and U24228 (N_24228,N_23545,N_23817);
nor U24229 (N_24229,N_23876,N_23503);
and U24230 (N_24230,N_23898,N_23846);
nand U24231 (N_24231,N_23680,N_23986);
xnor U24232 (N_24232,N_23848,N_23804);
and U24233 (N_24233,N_23624,N_23691);
nand U24234 (N_24234,N_23599,N_23531);
nor U24235 (N_24235,N_23751,N_23731);
xor U24236 (N_24236,N_23523,N_23716);
nand U24237 (N_24237,N_23647,N_23575);
nand U24238 (N_24238,N_23854,N_23565);
and U24239 (N_24239,N_23724,N_23682);
nand U24240 (N_24240,N_23720,N_23994);
and U24241 (N_24241,N_23941,N_23945);
or U24242 (N_24242,N_23633,N_23842);
nor U24243 (N_24243,N_23893,N_23861);
nor U24244 (N_24244,N_23995,N_23511);
xnor U24245 (N_24245,N_23908,N_23585);
and U24246 (N_24246,N_23999,N_23899);
and U24247 (N_24247,N_23989,N_23606);
xnor U24248 (N_24248,N_23668,N_23789);
and U24249 (N_24249,N_23936,N_23700);
xnor U24250 (N_24250,N_23610,N_23504);
and U24251 (N_24251,N_23988,N_23751);
and U24252 (N_24252,N_23826,N_23739);
xor U24253 (N_24253,N_23719,N_23611);
nand U24254 (N_24254,N_23600,N_23513);
nand U24255 (N_24255,N_23531,N_23986);
and U24256 (N_24256,N_23869,N_23669);
xor U24257 (N_24257,N_23537,N_23864);
or U24258 (N_24258,N_23746,N_23905);
nand U24259 (N_24259,N_23820,N_23715);
xnor U24260 (N_24260,N_23688,N_23559);
and U24261 (N_24261,N_23784,N_23801);
nand U24262 (N_24262,N_23867,N_23607);
and U24263 (N_24263,N_23514,N_23758);
xor U24264 (N_24264,N_23570,N_23711);
nor U24265 (N_24265,N_23933,N_23763);
xor U24266 (N_24266,N_23622,N_23835);
and U24267 (N_24267,N_23668,N_23931);
nand U24268 (N_24268,N_23916,N_23684);
nand U24269 (N_24269,N_23868,N_23840);
xnor U24270 (N_24270,N_23620,N_23571);
nor U24271 (N_24271,N_23768,N_23952);
or U24272 (N_24272,N_23638,N_23695);
and U24273 (N_24273,N_23834,N_23711);
or U24274 (N_24274,N_23883,N_23798);
xnor U24275 (N_24275,N_23613,N_23533);
nor U24276 (N_24276,N_23756,N_23872);
and U24277 (N_24277,N_23537,N_23919);
or U24278 (N_24278,N_23652,N_23796);
and U24279 (N_24279,N_23623,N_23707);
xnor U24280 (N_24280,N_23805,N_23999);
and U24281 (N_24281,N_23822,N_23694);
nand U24282 (N_24282,N_23606,N_23701);
and U24283 (N_24283,N_23526,N_23597);
xor U24284 (N_24284,N_23651,N_23744);
nand U24285 (N_24285,N_23994,N_23917);
or U24286 (N_24286,N_23690,N_23774);
or U24287 (N_24287,N_23593,N_23592);
xor U24288 (N_24288,N_23747,N_23536);
and U24289 (N_24289,N_23805,N_23539);
and U24290 (N_24290,N_23956,N_23550);
or U24291 (N_24291,N_23823,N_23929);
xnor U24292 (N_24292,N_23914,N_23884);
nor U24293 (N_24293,N_23767,N_23625);
xnor U24294 (N_24294,N_23910,N_23887);
xor U24295 (N_24295,N_23861,N_23652);
xor U24296 (N_24296,N_23832,N_23820);
nand U24297 (N_24297,N_23533,N_23939);
nand U24298 (N_24298,N_23970,N_23543);
and U24299 (N_24299,N_23660,N_23532);
and U24300 (N_24300,N_23692,N_23589);
or U24301 (N_24301,N_23992,N_23835);
and U24302 (N_24302,N_23622,N_23978);
and U24303 (N_24303,N_23845,N_23828);
nor U24304 (N_24304,N_23825,N_23694);
xnor U24305 (N_24305,N_23984,N_23566);
nor U24306 (N_24306,N_23526,N_23798);
xor U24307 (N_24307,N_23985,N_23583);
or U24308 (N_24308,N_23878,N_23514);
or U24309 (N_24309,N_23821,N_23758);
or U24310 (N_24310,N_23516,N_23987);
nor U24311 (N_24311,N_23680,N_23930);
and U24312 (N_24312,N_23509,N_23535);
and U24313 (N_24313,N_23562,N_23949);
xnor U24314 (N_24314,N_23878,N_23707);
nor U24315 (N_24315,N_23962,N_23884);
nand U24316 (N_24316,N_23769,N_23987);
or U24317 (N_24317,N_23556,N_23565);
nand U24318 (N_24318,N_23838,N_23572);
xor U24319 (N_24319,N_23758,N_23725);
or U24320 (N_24320,N_23632,N_23891);
nand U24321 (N_24321,N_23687,N_23581);
nor U24322 (N_24322,N_23650,N_23678);
nand U24323 (N_24323,N_23835,N_23535);
and U24324 (N_24324,N_23952,N_23924);
and U24325 (N_24325,N_23510,N_23839);
nor U24326 (N_24326,N_23667,N_23648);
or U24327 (N_24327,N_23796,N_23539);
nor U24328 (N_24328,N_23873,N_23867);
nand U24329 (N_24329,N_23905,N_23559);
nor U24330 (N_24330,N_23930,N_23532);
nor U24331 (N_24331,N_23950,N_23614);
and U24332 (N_24332,N_23659,N_23736);
nor U24333 (N_24333,N_23536,N_23844);
nand U24334 (N_24334,N_23832,N_23767);
and U24335 (N_24335,N_23983,N_23858);
nand U24336 (N_24336,N_23583,N_23694);
nand U24337 (N_24337,N_23623,N_23898);
xor U24338 (N_24338,N_23978,N_23892);
nor U24339 (N_24339,N_23574,N_23538);
nor U24340 (N_24340,N_23874,N_23899);
and U24341 (N_24341,N_23523,N_23951);
or U24342 (N_24342,N_23546,N_23613);
xnor U24343 (N_24343,N_23736,N_23723);
or U24344 (N_24344,N_23930,N_23805);
xnor U24345 (N_24345,N_23632,N_23660);
nand U24346 (N_24346,N_23964,N_23723);
nor U24347 (N_24347,N_23546,N_23606);
nor U24348 (N_24348,N_23671,N_23870);
xnor U24349 (N_24349,N_23727,N_23584);
and U24350 (N_24350,N_23802,N_23782);
and U24351 (N_24351,N_23846,N_23963);
xor U24352 (N_24352,N_23624,N_23792);
nand U24353 (N_24353,N_23986,N_23767);
nor U24354 (N_24354,N_23665,N_23763);
nor U24355 (N_24355,N_23752,N_23680);
nand U24356 (N_24356,N_23742,N_23861);
nor U24357 (N_24357,N_23641,N_23843);
nand U24358 (N_24358,N_23869,N_23765);
and U24359 (N_24359,N_23840,N_23560);
nand U24360 (N_24360,N_23587,N_23687);
nand U24361 (N_24361,N_23822,N_23994);
and U24362 (N_24362,N_23598,N_23921);
nor U24363 (N_24363,N_23505,N_23799);
and U24364 (N_24364,N_23993,N_23573);
and U24365 (N_24365,N_23562,N_23998);
and U24366 (N_24366,N_23773,N_23865);
or U24367 (N_24367,N_23861,N_23985);
or U24368 (N_24368,N_23817,N_23888);
or U24369 (N_24369,N_23742,N_23840);
and U24370 (N_24370,N_23796,N_23776);
nor U24371 (N_24371,N_23568,N_23603);
nand U24372 (N_24372,N_23916,N_23729);
nor U24373 (N_24373,N_23910,N_23963);
and U24374 (N_24374,N_23988,N_23642);
xor U24375 (N_24375,N_23577,N_23862);
nor U24376 (N_24376,N_23621,N_23607);
xnor U24377 (N_24377,N_23752,N_23800);
nand U24378 (N_24378,N_23638,N_23681);
nand U24379 (N_24379,N_23771,N_23510);
and U24380 (N_24380,N_23837,N_23577);
and U24381 (N_24381,N_23712,N_23885);
nor U24382 (N_24382,N_23834,N_23853);
or U24383 (N_24383,N_23924,N_23975);
nand U24384 (N_24384,N_23875,N_23859);
nand U24385 (N_24385,N_23565,N_23835);
and U24386 (N_24386,N_23516,N_23949);
or U24387 (N_24387,N_23755,N_23786);
xor U24388 (N_24388,N_23826,N_23644);
nand U24389 (N_24389,N_23518,N_23843);
and U24390 (N_24390,N_23761,N_23691);
nand U24391 (N_24391,N_23847,N_23797);
nand U24392 (N_24392,N_23817,N_23763);
nor U24393 (N_24393,N_23963,N_23819);
xor U24394 (N_24394,N_23967,N_23809);
or U24395 (N_24395,N_23513,N_23885);
or U24396 (N_24396,N_23506,N_23560);
or U24397 (N_24397,N_23650,N_23700);
and U24398 (N_24398,N_23742,N_23778);
or U24399 (N_24399,N_23910,N_23848);
or U24400 (N_24400,N_23776,N_23678);
or U24401 (N_24401,N_23943,N_23680);
xor U24402 (N_24402,N_23758,N_23732);
nor U24403 (N_24403,N_23798,N_23709);
and U24404 (N_24404,N_23836,N_23705);
or U24405 (N_24405,N_23977,N_23616);
nor U24406 (N_24406,N_23691,N_23781);
or U24407 (N_24407,N_23748,N_23704);
nand U24408 (N_24408,N_23508,N_23867);
nand U24409 (N_24409,N_23609,N_23534);
or U24410 (N_24410,N_23773,N_23809);
nor U24411 (N_24411,N_23739,N_23522);
xor U24412 (N_24412,N_23629,N_23786);
nor U24413 (N_24413,N_23792,N_23971);
and U24414 (N_24414,N_23686,N_23723);
or U24415 (N_24415,N_23783,N_23915);
and U24416 (N_24416,N_23799,N_23609);
xnor U24417 (N_24417,N_23779,N_23932);
nand U24418 (N_24418,N_23677,N_23981);
or U24419 (N_24419,N_23762,N_23700);
nand U24420 (N_24420,N_23667,N_23779);
xnor U24421 (N_24421,N_23809,N_23877);
xnor U24422 (N_24422,N_23789,N_23748);
and U24423 (N_24423,N_23585,N_23834);
xnor U24424 (N_24424,N_23837,N_23838);
nand U24425 (N_24425,N_23888,N_23799);
or U24426 (N_24426,N_23810,N_23636);
and U24427 (N_24427,N_23630,N_23646);
xnor U24428 (N_24428,N_23508,N_23565);
nand U24429 (N_24429,N_23905,N_23839);
nand U24430 (N_24430,N_23708,N_23876);
and U24431 (N_24431,N_23710,N_23527);
and U24432 (N_24432,N_23685,N_23572);
nand U24433 (N_24433,N_23525,N_23849);
nand U24434 (N_24434,N_23617,N_23502);
or U24435 (N_24435,N_23645,N_23558);
or U24436 (N_24436,N_23836,N_23571);
or U24437 (N_24437,N_23557,N_23581);
or U24438 (N_24438,N_23683,N_23613);
xnor U24439 (N_24439,N_23959,N_23752);
and U24440 (N_24440,N_23961,N_23672);
nor U24441 (N_24441,N_23919,N_23522);
xnor U24442 (N_24442,N_23540,N_23777);
and U24443 (N_24443,N_23927,N_23662);
and U24444 (N_24444,N_23813,N_23904);
and U24445 (N_24445,N_23953,N_23597);
and U24446 (N_24446,N_23622,N_23513);
or U24447 (N_24447,N_23606,N_23836);
nor U24448 (N_24448,N_23829,N_23592);
xnor U24449 (N_24449,N_23895,N_23695);
or U24450 (N_24450,N_23765,N_23790);
nand U24451 (N_24451,N_23834,N_23530);
or U24452 (N_24452,N_23623,N_23894);
or U24453 (N_24453,N_23630,N_23918);
nor U24454 (N_24454,N_23559,N_23505);
nor U24455 (N_24455,N_23736,N_23633);
nor U24456 (N_24456,N_23786,N_23782);
nor U24457 (N_24457,N_23766,N_23809);
xor U24458 (N_24458,N_23777,N_23892);
xnor U24459 (N_24459,N_23537,N_23905);
nand U24460 (N_24460,N_23864,N_23827);
xor U24461 (N_24461,N_23605,N_23975);
or U24462 (N_24462,N_23600,N_23712);
and U24463 (N_24463,N_23654,N_23621);
xnor U24464 (N_24464,N_23608,N_23793);
nand U24465 (N_24465,N_23937,N_23606);
and U24466 (N_24466,N_23644,N_23534);
and U24467 (N_24467,N_23773,N_23615);
nand U24468 (N_24468,N_23613,N_23980);
or U24469 (N_24469,N_23670,N_23672);
nand U24470 (N_24470,N_23855,N_23723);
or U24471 (N_24471,N_23830,N_23560);
xnor U24472 (N_24472,N_23983,N_23878);
nand U24473 (N_24473,N_23986,N_23966);
nand U24474 (N_24474,N_23780,N_23958);
or U24475 (N_24475,N_23780,N_23998);
nand U24476 (N_24476,N_23972,N_23667);
xnor U24477 (N_24477,N_23868,N_23689);
xor U24478 (N_24478,N_23553,N_23606);
or U24479 (N_24479,N_23852,N_23634);
nand U24480 (N_24480,N_23518,N_23835);
nand U24481 (N_24481,N_23727,N_23563);
and U24482 (N_24482,N_23716,N_23538);
nor U24483 (N_24483,N_23939,N_23722);
or U24484 (N_24484,N_23961,N_23507);
or U24485 (N_24485,N_23824,N_23599);
xnor U24486 (N_24486,N_23747,N_23822);
and U24487 (N_24487,N_23501,N_23710);
xor U24488 (N_24488,N_23857,N_23532);
nor U24489 (N_24489,N_23998,N_23526);
and U24490 (N_24490,N_23831,N_23674);
and U24491 (N_24491,N_23695,N_23899);
nand U24492 (N_24492,N_23801,N_23660);
and U24493 (N_24493,N_23706,N_23725);
nand U24494 (N_24494,N_23671,N_23837);
xor U24495 (N_24495,N_23618,N_23994);
and U24496 (N_24496,N_23540,N_23758);
nor U24497 (N_24497,N_23530,N_23683);
or U24498 (N_24498,N_23977,N_23505);
and U24499 (N_24499,N_23693,N_23601);
xor U24500 (N_24500,N_24240,N_24300);
or U24501 (N_24501,N_24451,N_24465);
and U24502 (N_24502,N_24442,N_24452);
nor U24503 (N_24503,N_24414,N_24255);
or U24504 (N_24504,N_24381,N_24496);
and U24505 (N_24505,N_24412,N_24060);
xnor U24506 (N_24506,N_24078,N_24369);
or U24507 (N_24507,N_24119,N_24396);
nand U24508 (N_24508,N_24021,N_24413);
and U24509 (N_24509,N_24242,N_24064);
nor U24510 (N_24510,N_24327,N_24473);
and U24511 (N_24511,N_24074,N_24354);
xor U24512 (N_24512,N_24339,N_24207);
and U24513 (N_24513,N_24007,N_24243);
or U24514 (N_24514,N_24206,N_24309);
nor U24515 (N_24515,N_24170,N_24357);
nand U24516 (N_24516,N_24211,N_24186);
or U24517 (N_24517,N_24422,N_24154);
or U24518 (N_24518,N_24398,N_24425);
and U24519 (N_24519,N_24157,N_24025);
nand U24520 (N_24520,N_24326,N_24185);
nor U24521 (N_24521,N_24387,N_24277);
and U24522 (N_24522,N_24023,N_24490);
and U24523 (N_24523,N_24230,N_24441);
nor U24524 (N_24524,N_24036,N_24378);
and U24525 (N_24525,N_24201,N_24343);
nor U24526 (N_24526,N_24337,N_24098);
and U24527 (N_24527,N_24139,N_24444);
nand U24528 (N_24528,N_24388,N_24426);
nand U24529 (N_24529,N_24392,N_24034);
xor U24530 (N_24530,N_24095,N_24006);
nor U24531 (N_24531,N_24436,N_24298);
xnor U24532 (N_24532,N_24429,N_24122);
or U24533 (N_24533,N_24279,N_24372);
or U24534 (N_24534,N_24477,N_24271);
xnor U24535 (N_24535,N_24345,N_24299);
or U24536 (N_24536,N_24248,N_24367);
or U24537 (N_24537,N_24432,N_24190);
xnor U24538 (N_24538,N_24333,N_24218);
or U24539 (N_24539,N_24081,N_24424);
nand U24540 (N_24540,N_24223,N_24180);
xor U24541 (N_24541,N_24056,N_24014);
and U24542 (N_24542,N_24137,N_24253);
and U24543 (N_24543,N_24498,N_24368);
nand U24544 (N_24544,N_24165,N_24022);
and U24545 (N_24545,N_24259,N_24316);
nand U24546 (N_24546,N_24152,N_24308);
xnor U24547 (N_24547,N_24177,N_24136);
nand U24548 (N_24548,N_24457,N_24312);
or U24549 (N_24549,N_24285,N_24251);
or U24550 (N_24550,N_24287,N_24407);
nand U24551 (N_24551,N_24408,N_24013);
nor U24552 (N_24552,N_24385,N_24335);
xnor U24553 (N_24553,N_24262,N_24289);
or U24554 (N_24554,N_24447,N_24020);
nor U24555 (N_24555,N_24075,N_24171);
and U24556 (N_24556,N_24461,N_24401);
xnor U24557 (N_24557,N_24043,N_24403);
and U24558 (N_24558,N_24062,N_24159);
nor U24559 (N_24559,N_24110,N_24116);
and U24560 (N_24560,N_24489,N_24303);
nor U24561 (N_24561,N_24449,N_24069);
nor U24562 (N_24562,N_24115,N_24295);
xnor U24563 (N_24563,N_24487,N_24358);
nand U24564 (N_24564,N_24213,N_24497);
or U24565 (N_24565,N_24435,N_24134);
nor U24566 (N_24566,N_24191,N_24376);
or U24567 (N_24567,N_24140,N_24146);
or U24568 (N_24568,N_24238,N_24061);
nor U24569 (N_24569,N_24224,N_24270);
or U24570 (N_24570,N_24173,N_24029);
and U24571 (N_24571,N_24433,N_24032);
xnor U24572 (N_24572,N_24313,N_24349);
nand U24573 (N_24573,N_24202,N_24492);
and U24574 (N_24574,N_24374,N_24305);
xnor U24575 (N_24575,N_24331,N_24482);
nor U24576 (N_24576,N_24417,N_24453);
nor U24577 (N_24577,N_24379,N_24252);
nand U24578 (N_24578,N_24005,N_24151);
nand U24579 (N_24579,N_24450,N_24306);
nand U24580 (N_24580,N_24200,N_24480);
or U24581 (N_24581,N_24082,N_24434);
or U24582 (N_24582,N_24012,N_24104);
xnor U24583 (N_24583,N_24227,N_24208);
or U24584 (N_24584,N_24281,N_24391);
nand U24585 (N_24585,N_24323,N_24090);
and U24586 (N_24586,N_24050,N_24419);
xor U24587 (N_24587,N_24024,N_24383);
nand U24588 (N_24588,N_24446,N_24045);
nand U24589 (N_24589,N_24468,N_24404);
and U24590 (N_24590,N_24031,N_24214);
xnor U24591 (N_24591,N_24059,N_24197);
xor U24592 (N_24592,N_24467,N_24189);
xnor U24593 (N_24593,N_24027,N_24149);
nor U24594 (N_24594,N_24071,N_24127);
and U24595 (N_24595,N_24117,N_24294);
or U24596 (N_24596,N_24340,N_24384);
xor U24597 (N_24597,N_24302,N_24263);
xor U24598 (N_24598,N_24073,N_24103);
and U24599 (N_24599,N_24125,N_24394);
or U24600 (N_24600,N_24009,N_24100);
xnor U24601 (N_24601,N_24113,N_24269);
and U24602 (N_24602,N_24229,N_24494);
and U24603 (N_24603,N_24355,N_24324);
nand U24604 (N_24604,N_24107,N_24237);
nand U24605 (N_24605,N_24373,N_24286);
xnor U24606 (N_24606,N_24430,N_24072);
and U24607 (N_24607,N_24364,N_24053);
nand U24608 (N_24608,N_24042,N_24019);
and U24609 (N_24609,N_24225,N_24123);
nor U24610 (N_24610,N_24063,N_24448);
and U24611 (N_24611,N_24011,N_24228);
xor U24612 (N_24612,N_24148,N_24096);
nand U24613 (N_24613,N_24194,N_24080);
or U24614 (N_24614,N_24344,N_24038);
or U24615 (N_24615,N_24010,N_24155);
xnor U24616 (N_24616,N_24455,N_24209);
nor U24617 (N_24617,N_24445,N_24280);
xor U24618 (N_24618,N_24421,N_24035);
nand U24619 (N_24619,N_24131,N_24239);
nor U24620 (N_24620,N_24484,N_24438);
nand U24621 (N_24621,N_24476,N_24472);
xor U24622 (N_24622,N_24405,N_24290);
nand U24623 (N_24623,N_24363,N_24478);
nor U24624 (N_24624,N_24321,N_24085);
xor U24625 (N_24625,N_24217,N_24052);
or U24626 (N_24626,N_24320,N_24192);
or U24627 (N_24627,N_24274,N_24030);
nand U24628 (N_24628,N_24334,N_24397);
nor U24629 (N_24629,N_24284,N_24348);
xnor U24630 (N_24630,N_24181,N_24215);
and U24631 (N_24631,N_24486,N_24428);
nor U24632 (N_24632,N_24283,N_24479);
nor U24633 (N_24633,N_24093,N_24493);
and U24634 (N_24634,N_24016,N_24301);
or U24635 (N_24635,N_24481,N_24356);
nand U24636 (N_24636,N_24244,N_24065);
nand U24637 (N_24637,N_24172,N_24499);
or U24638 (N_24638,N_24443,N_24114);
or U24639 (N_24639,N_24267,N_24199);
nor U24640 (N_24640,N_24328,N_24120);
and U24641 (N_24641,N_24393,N_24091);
and U24642 (N_24642,N_24166,N_24488);
nor U24643 (N_24643,N_24179,N_24322);
xnor U24644 (N_24644,N_24314,N_24341);
nand U24645 (N_24645,N_24147,N_24008);
nor U24646 (N_24646,N_24420,N_24000);
xnor U24647 (N_24647,N_24132,N_24288);
or U24648 (N_24648,N_24133,N_24458);
nor U24649 (N_24649,N_24070,N_24153);
or U24650 (N_24650,N_24454,N_24168);
nor U24651 (N_24651,N_24203,N_24351);
nor U24652 (N_24652,N_24247,N_24026);
nand U24653 (N_24653,N_24210,N_24233);
or U24654 (N_24654,N_24054,N_24418);
and U24655 (N_24655,N_24411,N_24291);
or U24656 (N_24656,N_24221,N_24099);
and U24657 (N_24657,N_24226,N_24018);
xor U24658 (N_24658,N_24205,N_24184);
or U24659 (N_24659,N_24278,N_24264);
or U24660 (N_24660,N_24282,N_24161);
and U24661 (N_24661,N_24097,N_24041);
or U24662 (N_24662,N_24195,N_24483);
and U24663 (N_24663,N_24048,N_24386);
nor U24664 (N_24664,N_24272,N_24163);
or U24665 (N_24665,N_24089,N_24268);
nor U24666 (N_24666,N_24187,N_24307);
xor U24667 (N_24667,N_24475,N_24491);
xor U24668 (N_24668,N_24040,N_24315);
nor U24669 (N_24669,N_24440,N_24220);
nor U24670 (N_24670,N_24317,N_24033);
xor U24671 (N_24671,N_24296,N_24245);
and U24672 (N_24672,N_24362,N_24111);
or U24673 (N_24673,N_24382,N_24439);
nand U24674 (N_24674,N_24402,N_24216);
and U24675 (N_24675,N_24256,N_24222);
and U24676 (N_24676,N_24182,N_24234);
xor U24677 (N_24677,N_24463,N_24347);
nor U24678 (N_24678,N_24410,N_24193);
xor U24679 (N_24679,N_24415,N_24126);
nand U24680 (N_24680,N_24361,N_24265);
nor U24681 (N_24681,N_24329,N_24047);
and U24682 (N_24682,N_24336,N_24460);
and U24683 (N_24683,N_24370,N_24332);
or U24684 (N_24684,N_24400,N_24437);
xor U24685 (N_24685,N_24260,N_24198);
nor U24686 (N_24686,N_24092,N_24456);
nand U24687 (N_24687,N_24338,N_24350);
nor U24688 (N_24688,N_24108,N_24086);
or U24689 (N_24689,N_24325,N_24156);
or U24690 (N_24690,N_24143,N_24360);
and U24691 (N_24691,N_24076,N_24112);
nand U24692 (N_24692,N_24250,N_24196);
or U24693 (N_24693,N_24219,N_24088);
xor U24694 (N_24694,N_24352,N_24004);
nand U24695 (N_24695,N_24462,N_24049);
nor U24696 (N_24696,N_24318,N_24395);
nor U24697 (N_24697,N_24145,N_24068);
xnor U24698 (N_24698,N_24375,N_24160);
nor U24699 (N_24699,N_24067,N_24311);
xnor U24700 (N_24700,N_24423,N_24231);
or U24701 (N_24701,N_24469,N_24261);
nor U24702 (N_24702,N_24001,N_24292);
xor U24703 (N_24703,N_24471,N_24365);
nand U24704 (N_24704,N_24051,N_24246);
nand U24705 (N_24705,N_24359,N_24002);
xnor U24706 (N_24706,N_24101,N_24017);
nand U24707 (N_24707,N_24121,N_24144);
nand U24708 (N_24708,N_24212,N_24150);
nand U24709 (N_24709,N_24174,N_24135);
and U24710 (N_24710,N_24106,N_24066);
nor U24711 (N_24711,N_24431,N_24276);
xnor U24712 (N_24712,N_24459,N_24046);
xnor U24713 (N_24713,N_24409,N_24380);
and U24714 (N_24714,N_24377,N_24175);
or U24715 (N_24715,N_24083,N_24130);
nand U24716 (N_24716,N_24079,N_24044);
and U24717 (N_24717,N_24319,N_24474);
xor U24718 (N_24718,N_24495,N_24102);
or U24719 (N_24719,N_24466,N_24167);
or U24720 (N_24720,N_24003,N_24128);
nor U24721 (N_24721,N_24158,N_24310);
or U24722 (N_24722,N_24297,N_24204);
nand U24723 (N_24723,N_24266,N_24254);
and U24724 (N_24724,N_24273,N_24485);
nor U24725 (N_24725,N_24039,N_24109);
nand U24726 (N_24726,N_24164,N_24169);
or U24727 (N_24727,N_24258,N_24142);
nand U24728 (N_24728,N_24235,N_24176);
and U24729 (N_24729,N_24232,N_24406);
nand U24730 (N_24730,N_24342,N_24118);
nor U24731 (N_24731,N_24057,N_24094);
nor U24732 (N_24732,N_24183,N_24141);
and U24733 (N_24733,N_24330,N_24249);
or U24734 (N_24734,N_24236,N_24390);
xnor U24735 (N_24735,N_24015,N_24464);
xnor U24736 (N_24736,N_24399,N_24188);
nor U24737 (N_24737,N_24138,N_24275);
or U24738 (N_24738,N_24241,N_24124);
or U24739 (N_24739,N_24178,N_24304);
nand U24740 (N_24740,N_24346,N_24416);
nor U24741 (N_24741,N_24028,N_24087);
nor U24742 (N_24742,N_24084,N_24293);
or U24743 (N_24743,N_24257,N_24037);
nand U24744 (N_24744,N_24353,N_24055);
nor U24745 (N_24745,N_24077,N_24366);
xnor U24746 (N_24746,N_24427,N_24389);
and U24747 (N_24747,N_24105,N_24371);
nor U24748 (N_24748,N_24162,N_24129);
nor U24749 (N_24749,N_24470,N_24058);
xnor U24750 (N_24750,N_24451,N_24029);
nor U24751 (N_24751,N_24058,N_24443);
or U24752 (N_24752,N_24302,N_24410);
nand U24753 (N_24753,N_24343,N_24429);
nand U24754 (N_24754,N_24224,N_24459);
nand U24755 (N_24755,N_24420,N_24473);
and U24756 (N_24756,N_24279,N_24082);
nor U24757 (N_24757,N_24058,N_24290);
or U24758 (N_24758,N_24295,N_24007);
nor U24759 (N_24759,N_24017,N_24355);
nand U24760 (N_24760,N_24219,N_24291);
xnor U24761 (N_24761,N_24236,N_24454);
nand U24762 (N_24762,N_24461,N_24136);
nand U24763 (N_24763,N_24128,N_24310);
xor U24764 (N_24764,N_24420,N_24018);
or U24765 (N_24765,N_24361,N_24339);
or U24766 (N_24766,N_24224,N_24454);
nor U24767 (N_24767,N_24027,N_24371);
and U24768 (N_24768,N_24037,N_24438);
xnor U24769 (N_24769,N_24186,N_24497);
nand U24770 (N_24770,N_24158,N_24154);
and U24771 (N_24771,N_24212,N_24259);
and U24772 (N_24772,N_24347,N_24455);
nand U24773 (N_24773,N_24462,N_24222);
xor U24774 (N_24774,N_24041,N_24330);
nor U24775 (N_24775,N_24404,N_24398);
or U24776 (N_24776,N_24351,N_24080);
xnor U24777 (N_24777,N_24164,N_24222);
nand U24778 (N_24778,N_24186,N_24201);
nor U24779 (N_24779,N_24381,N_24310);
or U24780 (N_24780,N_24031,N_24133);
nor U24781 (N_24781,N_24278,N_24063);
nand U24782 (N_24782,N_24454,N_24363);
or U24783 (N_24783,N_24047,N_24136);
or U24784 (N_24784,N_24039,N_24095);
and U24785 (N_24785,N_24193,N_24315);
nand U24786 (N_24786,N_24105,N_24418);
nor U24787 (N_24787,N_24248,N_24116);
nor U24788 (N_24788,N_24365,N_24087);
and U24789 (N_24789,N_24009,N_24001);
nor U24790 (N_24790,N_24423,N_24061);
xor U24791 (N_24791,N_24122,N_24164);
nand U24792 (N_24792,N_24013,N_24311);
or U24793 (N_24793,N_24144,N_24420);
and U24794 (N_24794,N_24290,N_24377);
or U24795 (N_24795,N_24067,N_24421);
nor U24796 (N_24796,N_24264,N_24415);
nand U24797 (N_24797,N_24199,N_24281);
nand U24798 (N_24798,N_24344,N_24124);
xor U24799 (N_24799,N_24320,N_24397);
nand U24800 (N_24800,N_24017,N_24406);
nand U24801 (N_24801,N_24312,N_24243);
or U24802 (N_24802,N_24498,N_24060);
or U24803 (N_24803,N_24132,N_24322);
and U24804 (N_24804,N_24312,N_24009);
nor U24805 (N_24805,N_24237,N_24193);
nand U24806 (N_24806,N_24421,N_24326);
xnor U24807 (N_24807,N_24096,N_24308);
and U24808 (N_24808,N_24068,N_24130);
nor U24809 (N_24809,N_24496,N_24190);
xor U24810 (N_24810,N_24391,N_24002);
xnor U24811 (N_24811,N_24148,N_24452);
nand U24812 (N_24812,N_24393,N_24375);
nor U24813 (N_24813,N_24329,N_24043);
nor U24814 (N_24814,N_24004,N_24302);
nand U24815 (N_24815,N_24136,N_24251);
xor U24816 (N_24816,N_24215,N_24083);
xnor U24817 (N_24817,N_24095,N_24062);
and U24818 (N_24818,N_24285,N_24286);
nor U24819 (N_24819,N_24047,N_24425);
and U24820 (N_24820,N_24373,N_24216);
nor U24821 (N_24821,N_24390,N_24149);
xnor U24822 (N_24822,N_24045,N_24397);
nand U24823 (N_24823,N_24453,N_24060);
xnor U24824 (N_24824,N_24423,N_24228);
nor U24825 (N_24825,N_24323,N_24132);
and U24826 (N_24826,N_24261,N_24295);
nand U24827 (N_24827,N_24081,N_24202);
nand U24828 (N_24828,N_24196,N_24307);
or U24829 (N_24829,N_24355,N_24082);
xor U24830 (N_24830,N_24117,N_24219);
nand U24831 (N_24831,N_24245,N_24375);
xor U24832 (N_24832,N_24229,N_24228);
nor U24833 (N_24833,N_24184,N_24023);
nor U24834 (N_24834,N_24152,N_24486);
or U24835 (N_24835,N_24047,N_24231);
nor U24836 (N_24836,N_24233,N_24372);
nor U24837 (N_24837,N_24248,N_24150);
and U24838 (N_24838,N_24085,N_24007);
nor U24839 (N_24839,N_24158,N_24185);
or U24840 (N_24840,N_24455,N_24322);
xor U24841 (N_24841,N_24482,N_24372);
xor U24842 (N_24842,N_24367,N_24316);
or U24843 (N_24843,N_24283,N_24358);
nand U24844 (N_24844,N_24421,N_24394);
or U24845 (N_24845,N_24240,N_24109);
xnor U24846 (N_24846,N_24489,N_24107);
nand U24847 (N_24847,N_24172,N_24396);
nor U24848 (N_24848,N_24380,N_24235);
nand U24849 (N_24849,N_24322,N_24081);
or U24850 (N_24850,N_24240,N_24289);
xor U24851 (N_24851,N_24291,N_24149);
xnor U24852 (N_24852,N_24241,N_24206);
xnor U24853 (N_24853,N_24298,N_24448);
nor U24854 (N_24854,N_24493,N_24304);
xor U24855 (N_24855,N_24422,N_24005);
xnor U24856 (N_24856,N_24158,N_24166);
and U24857 (N_24857,N_24168,N_24308);
or U24858 (N_24858,N_24112,N_24163);
nand U24859 (N_24859,N_24444,N_24102);
or U24860 (N_24860,N_24491,N_24156);
nand U24861 (N_24861,N_24118,N_24197);
or U24862 (N_24862,N_24429,N_24486);
nand U24863 (N_24863,N_24370,N_24482);
nand U24864 (N_24864,N_24132,N_24285);
nand U24865 (N_24865,N_24238,N_24112);
nor U24866 (N_24866,N_24359,N_24162);
and U24867 (N_24867,N_24414,N_24437);
or U24868 (N_24868,N_24283,N_24311);
and U24869 (N_24869,N_24236,N_24265);
nand U24870 (N_24870,N_24324,N_24198);
nor U24871 (N_24871,N_24030,N_24013);
nor U24872 (N_24872,N_24243,N_24152);
nor U24873 (N_24873,N_24222,N_24481);
nand U24874 (N_24874,N_24124,N_24020);
xnor U24875 (N_24875,N_24295,N_24027);
or U24876 (N_24876,N_24494,N_24262);
or U24877 (N_24877,N_24470,N_24021);
and U24878 (N_24878,N_24076,N_24022);
and U24879 (N_24879,N_24330,N_24088);
or U24880 (N_24880,N_24295,N_24209);
xor U24881 (N_24881,N_24279,N_24039);
and U24882 (N_24882,N_24272,N_24380);
or U24883 (N_24883,N_24385,N_24378);
and U24884 (N_24884,N_24435,N_24387);
xnor U24885 (N_24885,N_24443,N_24413);
and U24886 (N_24886,N_24289,N_24417);
xnor U24887 (N_24887,N_24409,N_24059);
xnor U24888 (N_24888,N_24272,N_24138);
xnor U24889 (N_24889,N_24148,N_24314);
and U24890 (N_24890,N_24357,N_24031);
or U24891 (N_24891,N_24411,N_24092);
nor U24892 (N_24892,N_24493,N_24497);
and U24893 (N_24893,N_24008,N_24180);
or U24894 (N_24894,N_24073,N_24164);
nand U24895 (N_24895,N_24299,N_24428);
or U24896 (N_24896,N_24198,N_24393);
nor U24897 (N_24897,N_24356,N_24186);
or U24898 (N_24898,N_24216,N_24022);
nand U24899 (N_24899,N_24120,N_24082);
or U24900 (N_24900,N_24098,N_24188);
or U24901 (N_24901,N_24391,N_24055);
xor U24902 (N_24902,N_24144,N_24088);
xor U24903 (N_24903,N_24162,N_24183);
xnor U24904 (N_24904,N_24084,N_24326);
nand U24905 (N_24905,N_24088,N_24382);
or U24906 (N_24906,N_24230,N_24180);
xnor U24907 (N_24907,N_24027,N_24209);
or U24908 (N_24908,N_24031,N_24348);
nand U24909 (N_24909,N_24193,N_24049);
nand U24910 (N_24910,N_24373,N_24301);
or U24911 (N_24911,N_24312,N_24319);
nand U24912 (N_24912,N_24292,N_24275);
nor U24913 (N_24913,N_24056,N_24420);
nand U24914 (N_24914,N_24019,N_24478);
nand U24915 (N_24915,N_24281,N_24409);
xnor U24916 (N_24916,N_24226,N_24256);
xor U24917 (N_24917,N_24069,N_24212);
nor U24918 (N_24918,N_24079,N_24251);
or U24919 (N_24919,N_24000,N_24402);
nand U24920 (N_24920,N_24259,N_24447);
or U24921 (N_24921,N_24026,N_24021);
or U24922 (N_24922,N_24108,N_24182);
or U24923 (N_24923,N_24455,N_24343);
nor U24924 (N_24924,N_24396,N_24472);
or U24925 (N_24925,N_24144,N_24142);
nor U24926 (N_24926,N_24477,N_24287);
and U24927 (N_24927,N_24447,N_24400);
and U24928 (N_24928,N_24323,N_24354);
nor U24929 (N_24929,N_24312,N_24220);
nand U24930 (N_24930,N_24317,N_24269);
and U24931 (N_24931,N_24236,N_24165);
or U24932 (N_24932,N_24109,N_24099);
nand U24933 (N_24933,N_24428,N_24295);
xnor U24934 (N_24934,N_24039,N_24336);
nand U24935 (N_24935,N_24459,N_24157);
and U24936 (N_24936,N_24367,N_24013);
or U24937 (N_24937,N_24461,N_24311);
or U24938 (N_24938,N_24281,N_24367);
nor U24939 (N_24939,N_24478,N_24026);
xor U24940 (N_24940,N_24316,N_24460);
and U24941 (N_24941,N_24284,N_24478);
xnor U24942 (N_24942,N_24226,N_24451);
xor U24943 (N_24943,N_24357,N_24019);
or U24944 (N_24944,N_24271,N_24274);
nor U24945 (N_24945,N_24039,N_24297);
or U24946 (N_24946,N_24032,N_24143);
nand U24947 (N_24947,N_24443,N_24110);
xnor U24948 (N_24948,N_24222,N_24055);
nand U24949 (N_24949,N_24089,N_24161);
nor U24950 (N_24950,N_24472,N_24059);
and U24951 (N_24951,N_24318,N_24057);
or U24952 (N_24952,N_24007,N_24463);
and U24953 (N_24953,N_24077,N_24076);
nor U24954 (N_24954,N_24315,N_24299);
nand U24955 (N_24955,N_24155,N_24408);
or U24956 (N_24956,N_24191,N_24114);
nand U24957 (N_24957,N_24145,N_24207);
xor U24958 (N_24958,N_24438,N_24361);
or U24959 (N_24959,N_24082,N_24447);
nand U24960 (N_24960,N_24163,N_24297);
nand U24961 (N_24961,N_24136,N_24159);
nor U24962 (N_24962,N_24339,N_24430);
nor U24963 (N_24963,N_24055,N_24269);
xor U24964 (N_24964,N_24039,N_24194);
or U24965 (N_24965,N_24486,N_24188);
and U24966 (N_24966,N_24336,N_24134);
nand U24967 (N_24967,N_24449,N_24345);
nand U24968 (N_24968,N_24387,N_24460);
nor U24969 (N_24969,N_24143,N_24379);
nand U24970 (N_24970,N_24234,N_24111);
nor U24971 (N_24971,N_24295,N_24165);
or U24972 (N_24972,N_24227,N_24147);
nand U24973 (N_24973,N_24461,N_24446);
nor U24974 (N_24974,N_24364,N_24270);
nand U24975 (N_24975,N_24044,N_24068);
or U24976 (N_24976,N_24468,N_24005);
or U24977 (N_24977,N_24064,N_24081);
nor U24978 (N_24978,N_24008,N_24268);
xnor U24979 (N_24979,N_24236,N_24078);
xor U24980 (N_24980,N_24406,N_24253);
xnor U24981 (N_24981,N_24497,N_24073);
or U24982 (N_24982,N_24031,N_24158);
xor U24983 (N_24983,N_24232,N_24157);
nand U24984 (N_24984,N_24042,N_24240);
nor U24985 (N_24985,N_24284,N_24137);
xor U24986 (N_24986,N_24253,N_24427);
nor U24987 (N_24987,N_24271,N_24471);
nor U24988 (N_24988,N_24031,N_24395);
or U24989 (N_24989,N_24208,N_24308);
xnor U24990 (N_24990,N_24499,N_24219);
or U24991 (N_24991,N_24265,N_24450);
and U24992 (N_24992,N_24341,N_24003);
xor U24993 (N_24993,N_24118,N_24463);
and U24994 (N_24994,N_24485,N_24241);
nand U24995 (N_24995,N_24189,N_24044);
and U24996 (N_24996,N_24253,N_24112);
nand U24997 (N_24997,N_24311,N_24202);
or U24998 (N_24998,N_24190,N_24087);
nand U24999 (N_24999,N_24025,N_24334);
or U25000 (N_25000,N_24691,N_24800);
nand U25001 (N_25001,N_24540,N_24585);
xnor U25002 (N_25002,N_24922,N_24698);
or U25003 (N_25003,N_24650,N_24633);
nor U25004 (N_25004,N_24736,N_24882);
and U25005 (N_25005,N_24911,N_24913);
or U25006 (N_25006,N_24660,N_24519);
or U25007 (N_25007,N_24915,N_24887);
nand U25008 (N_25008,N_24796,N_24825);
xor U25009 (N_25009,N_24646,N_24923);
and U25010 (N_25010,N_24728,N_24511);
and U25011 (N_25011,N_24997,N_24758);
xnor U25012 (N_25012,N_24544,N_24550);
and U25013 (N_25013,N_24600,N_24584);
and U25014 (N_25014,N_24576,N_24530);
nor U25015 (N_25015,N_24738,N_24756);
and U25016 (N_25016,N_24788,N_24675);
xor U25017 (N_25017,N_24921,N_24626);
and U25018 (N_25018,N_24851,N_24984);
or U25019 (N_25019,N_24569,N_24986);
or U25020 (N_25020,N_24876,N_24674);
and U25021 (N_25021,N_24558,N_24782);
nand U25022 (N_25022,N_24856,N_24898);
and U25023 (N_25023,N_24582,N_24652);
and U25024 (N_25024,N_24718,N_24719);
and U25025 (N_25025,N_24873,N_24501);
xnor U25026 (N_25026,N_24790,N_24505);
nor U25027 (N_25027,N_24679,N_24603);
nor U25028 (N_25028,N_24663,N_24656);
nand U25029 (N_25029,N_24586,N_24573);
xnor U25030 (N_25030,N_24725,N_24637);
or U25031 (N_25031,N_24744,N_24535);
xor U25032 (N_25032,N_24785,N_24534);
xnor U25033 (N_25033,N_24936,N_24602);
nor U25034 (N_25034,N_24754,N_24697);
nand U25035 (N_25035,N_24570,N_24543);
and U25036 (N_25036,N_24779,N_24716);
nand U25037 (N_25037,N_24925,N_24583);
nand U25038 (N_25038,N_24917,N_24651);
nand U25039 (N_25039,N_24566,N_24590);
xor U25040 (N_25040,N_24618,N_24761);
nor U25041 (N_25041,N_24955,N_24889);
nor U25042 (N_25042,N_24745,N_24737);
xor U25043 (N_25043,N_24730,N_24580);
nor U25044 (N_25044,N_24895,N_24561);
and U25045 (N_25045,N_24926,N_24962);
or U25046 (N_25046,N_24552,N_24639);
or U25047 (N_25047,N_24676,N_24808);
and U25048 (N_25048,N_24508,N_24980);
nor U25049 (N_25049,N_24933,N_24578);
and U25050 (N_25050,N_24733,N_24912);
nor U25051 (N_25051,N_24669,N_24806);
or U25052 (N_25052,N_24907,N_24867);
or U25053 (N_25053,N_24613,N_24765);
or U25054 (N_25054,N_24568,N_24598);
and U25055 (N_25055,N_24878,N_24666);
xnor U25056 (N_25056,N_24801,N_24546);
or U25057 (N_25057,N_24844,N_24963);
xnor U25058 (N_25058,N_24849,N_24942);
and U25059 (N_25059,N_24696,N_24909);
nor U25060 (N_25060,N_24644,N_24845);
or U25061 (N_25061,N_24727,N_24510);
or U25062 (N_25062,N_24563,N_24641);
and U25063 (N_25063,N_24930,N_24688);
xor U25064 (N_25064,N_24700,N_24556);
and U25065 (N_25065,N_24711,N_24871);
and U25066 (N_25066,N_24824,N_24720);
xnor U25067 (N_25067,N_24571,N_24807);
nand U25068 (N_25068,N_24786,N_24972);
nor U25069 (N_25069,N_24531,N_24662);
and U25070 (N_25070,N_24694,N_24717);
nor U25071 (N_25071,N_24577,N_24919);
or U25072 (N_25072,N_24755,N_24766);
nor U25073 (N_25073,N_24682,N_24635);
nand U25074 (N_25074,N_24702,N_24743);
xor U25075 (N_25075,N_24847,N_24502);
nor U25076 (N_25076,N_24701,N_24541);
xor U25077 (N_25077,N_24763,N_24833);
or U25078 (N_25078,N_24832,N_24950);
nand U25079 (N_25079,N_24593,N_24939);
nor U25080 (N_25080,N_24732,N_24841);
and U25081 (N_25081,N_24905,N_24750);
or U25082 (N_25082,N_24994,N_24523);
and U25083 (N_25083,N_24865,N_24961);
and U25084 (N_25084,N_24843,N_24545);
or U25085 (N_25085,N_24989,N_24695);
or U25086 (N_25086,N_24974,N_24802);
nor U25087 (N_25087,N_24692,N_24614);
nor U25088 (N_25088,N_24914,N_24529);
and U25089 (N_25089,N_24978,N_24524);
or U25090 (N_25090,N_24703,N_24596);
xnor U25091 (N_25091,N_24916,N_24854);
and U25092 (N_25092,N_24901,N_24612);
xnor U25093 (N_25093,N_24891,N_24855);
or U25094 (N_25094,N_24707,N_24734);
and U25095 (N_25095,N_24504,N_24789);
or U25096 (N_25096,N_24741,N_24759);
nor U25097 (N_25097,N_24599,N_24860);
nor U25098 (N_25098,N_24987,N_24776);
nor U25099 (N_25099,N_24653,N_24632);
or U25100 (N_25100,N_24668,N_24861);
and U25101 (N_25101,N_24944,N_24503);
nor U25102 (N_25102,N_24673,N_24588);
xor U25103 (N_25103,N_24814,N_24509);
xor U25104 (N_25104,N_24645,N_24817);
and U25105 (N_25105,N_24826,N_24623);
or U25106 (N_25106,N_24998,N_24985);
xor U25107 (N_25107,N_24611,N_24815);
nand U25108 (N_25108,N_24908,N_24553);
xor U25109 (N_25109,N_24559,N_24672);
nor U25110 (N_25110,N_24522,N_24798);
and U25111 (N_25111,N_24538,N_24627);
or U25112 (N_25112,N_24794,N_24670);
and U25113 (N_25113,N_24677,N_24533);
nor U25114 (N_25114,N_24512,N_24951);
nand U25115 (N_25115,N_24705,N_24838);
or U25116 (N_25116,N_24999,N_24591);
or U25117 (N_25117,N_24947,N_24760);
nand U25118 (N_25118,N_24771,N_24957);
and U25119 (N_25119,N_24729,N_24671);
xor U25120 (N_25120,N_24513,N_24858);
or U25121 (N_25121,N_24893,N_24875);
nand U25122 (N_25122,N_24708,N_24990);
or U25123 (N_25123,N_24956,N_24579);
and U25124 (N_25124,N_24954,N_24966);
or U25125 (N_25125,N_24795,N_24687);
xnor U25126 (N_25126,N_24879,N_24746);
xnor U25127 (N_25127,N_24629,N_24864);
nand U25128 (N_25128,N_24830,N_24622);
xnor U25129 (N_25129,N_24597,N_24965);
nor U25130 (N_25130,N_24836,N_24667);
and U25131 (N_25131,N_24935,N_24804);
nand U25132 (N_25132,N_24731,N_24615);
nand U25133 (N_25133,N_24967,N_24837);
and U25134 (N_25134,N_24564,N_24747);
xor U25135 (N_25135,N_24983,N_24781);
or U25136 (N_25136,N_24799,N_24778);
xor U25137 (N_25137,N_24740,N_24689);
or U25138 (N_25138,N_24940,N_24631);
nor U25139 (N_25139,N_24749,N_24772);
and U25140 (N_25140,N_24797,N_24938);
nor U25141 (N_25141,N_24880,N_24557);
and U25142 (N_25142,N_24681,N_24828);
nand U25143 (N_25143,N_24686,N_24555);
nand U25144 (N_25144,N_24767,N_24918);
nor U25145 (N_25145,N_24948,N_24812);
xor U25146 (N_25146,N_24848,N_24960);
nand U25147 (N_25147,N_24910,N_24636);
nor U25148 (N_25148,N_24827,N_24784);
nor U25149 (N_25149,N_24852,N_24520);
xor U25150 (N_25150,N_24969,N_24872);
nand U25151 (N_25151,N_24515,N_24621);
nand U25152 (N_25152,N_24565,N_24949);
nor U25153 (N_25153,N_24595,N_24774);
and U25154 (N_25154,N_24958,N_24775);
xor U25155 (N_25155,N_24979,N_24793);
or U25156 (N_25156,N_24589,N_24968);
nor U25157 (N_25157,N_24581,N_24693);
and U25158 (N_25158,N_24929,N_24721);
and U25159 (N_25159,N_24609,N_24946);
or U25160 (N_25160,N_24932,N_24710);
xor U25161 (N_25161,N_24560,N_24890);
or U25162 (N_25162,N_24587,N_24610);
and U25163 (N_25163,N_24648,N_24724);
nor U25164 (N_25164,N_24977,N_24823);
or U25165 (N_25165,N_24991,N_24988);
or U25166 (N_25166,N_24630,N_24964);
nor U25167 (N_25167,N_24869,N_24791);
or U25168 (N_25168,N_24619,N_24709);
nand U25169 (N_25169,N_24517,N_24680);
xor U25170 (N_25170,N_24769,N_24726);
or U25171 (N_25171,N_24715,N_24521);
nor U25172 (N_25172,N_24937,N_24883);
nand U25173 (N_25173,N_24748,N_24976);
xnor U25174 (N_25174,N_24518,N_24959);
and U25175 (N_25175,N_24699,N_24810);
xnor U25176 (N_25176,N_24846,N_24594);
nand U25177 (N_25177,N_24506,N_24567);
xor U25178 (N_25178,N_24712,N_24768);
and U25179 (N_25179,N_24548,N_24777);
nand U25180 (N_25180,N_24659,N_24975);
or U25181 (N_25181,N_24780,N_24894);
and U25182 (N_25182,N_24661,N_24642);
or U25183 (N_25183,N_24608,N_24886);
and U25184 (N_25184,N_24607,N_24752);
or U25185 (N_25185,N_24649,N_24742);
nand U25186 (N_25186,N_24902,N_24904);
and U25187 (N_25187,N_24866,N_24722);
xnor U25188 (N_25188,N_24616,N_24704);
xor U25189 (N_25189,N_24792,N_24945);
nand U25190 (N_25190,N_24970,N_24549);
and U25191 (N_25191,N_24850,N_24617);
xnor U25192 (N_25192,N_24992,N_24842);
xor U25193 (N_25193,N_24862,N_24877);
nor U25194 (N_25194,N_24857,N_24516);
or U25195 (N_25195,N_24996,N_24514);
or U25196 (N_25196,N_24829,N_24874);
nor U25197 (N_25197,N_24542,N_24931);
and U25198 (N_25198,N_24764,N_24820);
xnor U25199 (N_25199,N_24952,N_24606);
or U25200 (N_25200,N_24803,N_24625);
or U25201 (N_25201,N_24500,N_24863);
and U25202 (N_25202,N_24973,N_24928);
and U25203 (N_25203,N_24537,N_24624);
or U25204 (N_25204,N_24982,N_24528);
nor U25205 (N_25205,N_24525,N_24684);
nand U25206 (N_25206,N_24884,N_24575);
and U25207 (N_25207,N_24787,N_24547);
nand U25208 (N_25208,N_24536,N_24993);
nand U25209 (N_25209,N_24628,N_24818);
and U25210 (N_25210,N_24805,N_24507);
nand U25211 (N_25211,N_24643,N_24604);
or U25212 (N_25212,N_24574,N_24840);
xnor U25213 (N_25213,N_24813,N_24941);
xor U25214 (N_25214,N_24551,N_24739);
or U25215 (N_25215,N_24572,N_24757);
or U25216 (N_25216,N_24809,N_24562);
or U25217 (N_25217,N_24640,N_24834);
and U25218 (N_25218,N_24620,N_24527);
xnor U25219 (N_25219,N_24783,N_24920);
nand U25220 (N_25220,N_24835,N_24655);
or U25221 (N_25221,N_24816,N_24751);
nand U25222 (N_25222,N_24868,N_24735);
or U25223 (N_25223,N_24714,N_24554);
xnor U25224 (N_25224,N_24995,N_24683);
nand U25225 (N_25225,N_24927,N_24723);
xor U25226 (N_25226,N_24526,N_24870);
nor U25227 (N_25227,N_24831,N_24859);
xor U25228 (N_25228,N_24678,N_24888);
and U25229 (N_25229,N_24592,N_24657);
and U25230 (N_25230,N_24897,N_24971);
nand U25231 (N_25231,N_24881,N_24634);
or U25232 (N_25232,N_24839,N_24532);
nand U25233 (N_25233,N_24685,N_24899);
nand U25234 (N_25234,N_24690,N_24981);
nor U25235 (N_25235,N_24903,N_24906);
nand U25236 (N_25236,N_24853,N_24819);
xnor U25237 (N_25237,N_24539,N_24770);
or U25238 (N_25238,N_24601,N_24658);
nor U25239 (N_25239,N_24638,N_24811);
and U25240 (N_25240,N_24822,N_24892);
nor U25241 (N_25241,N_24762,N_24943);
xor U25242 (N_25242,N_24647,N_24706);
and U25243 (N_25243,N_24934,N_24953);
nor U25244 (N_25244,N_24665,N_24900);
xor U25245 (N_25245,N_24821,N_24664);
xnor U25246 (N_25246,N_24605,N_24885);
xnor U25247 (N_25247,N_24753,N_24713);
or U25248 (N_25248,N_24924,N_24896);
and U25249 (N_25249,N_24654,N_24773);
nor U25250 (N_25250,N_24500,N_24746);
or U25251 (N_25251,N_24795,N_24802);
nor U25252 (N_25252,N_24950,N_24852);
or U25253 (N_25253,N_24879,N_24686);
nand U25254 (N_25254,N_24667,N_24501);
or U25255 (N_25255,N_24678,N_24752);
xor U25256 (N_25256,N_24917,N_24830);
or U25257 (N_25257,N_24821,N_24639);
nand U25258 (N_25258,N_24540,N_24688);
nor U25259 (N_25259,N_24604,N_24764);
nand U25260 (N_25260,N_24670,N_24648);
nand U25261 (N_25261,N_24799,N_24853);
or U25262 (N_25262,N_24576,N_24647);
or U25263 (N_25263,N_24974,N_24551);
nand U25264 (N_25264,N_24991,N_24978);
nand U25265 (N_25265,N_24813,N_24773);
nor U25266 (N_25266,N_24735,N_24857);
xor U25267 (N_25267,N_24602,N_24820);
nor U25268 (N_25268,N_24904,N_24614);
nand U25269 (N_25269,N_24541,N_24879);
or U25270 (N_25270,N_24920,N_24939);
nor U25271 (N_25271,N_24843,N_24525);
nand U25272 (N_25272,N_24929,N_24621);
nor U25273 (N_25273,N_24667,N_24901);
nand U25274 (N_25274,N_24530,N_24995);
nor U25275 (N_25275,N_24618,N_24774);
nand U25276 (N_25276,N_24727,N_24526);
nand U25277 (N_25277,N_24579,N_24761);
and U25278 (N_25278,N_24927,N_24512);
and U25279 (N_25279,N_24693,N_24545);
and U25280 (N_25280,N_24861,N_24831);
or U25281 (N_25281,N_24938,N_24996);
or U25282 (N_25282,N_24535,N_24750);
nor U25283 (N_25283,N_24554,N_24944);
nand U25284 (N_25284,N_24744,N_24688);
or U25285 (N_25285,N_24701,N_24697);
nor U25286 (N_25286,N_24875,N_24889);
nor U25287 (N_25287,N_24687,N_24515);
nor U25288 (N_25288,N_24605,N_24964);
nor U25289 (N_25289,N_24977,N_24720);
nand U25290 (N_25290,N_24906,N_24530);
nand U25291 (N_25291,N_24722,N_24783);
or U25292 (N_25292,N_24942,N_24770);
nor U25293 (N_25293,N_24665,N_24510);
and U25294 (N_25294,N_24594,N_24901);
and U25295 (N_25295,N_24790,N_24561);
nor U25296 (N_25296,N_24578,N_24960);
nand U25297 (N_25297,N_24828,N_24838);
and U25298 (N_25298,N_24924,N_24639);
or U25299 (N_25299,N_24779,N_24621);
and U25300 (N_25300,N_24833,N_24707);
nand U25301 (N_25301,N_24991,N_24798);
or U25302 (N_25302,N_24748,N_24980);
nor U25303 (N_25303,N_24957,N_24703);
and U25304 (N_25304,N_24898,N_24929);
nand U25305 (N_25305,N_24573,N_24560);
nor U25306 (N_25306,N_24958,N_24518);
xor U25307 (N_25307,N_24928,N_24607);
nand U25308 (N_25308,N_24518,N_24689);
or U25309 (N_25309,N_24664,N_24987);
nor U25310 (N_25310,N_24552,N_24900);
nand U25311 (N_25311,N_24896,N_24686);
xor U25312 (N_25312,N_24810,N_24636);
xor U25313 (N_25313,N_24996,N_24979);
xor U25314 (N_25314,N_24701,N_24969);
xor U25315 (N_25315,N_24757,N_24718);
nor U25316 (N_25316,N_24821,N_24962);
and U25317 (N_25317,N_24645,N_24649);
xor U25318 (N_25318,N_24819,N_24908);
and U25319 (N_25319,N_24559,N_24938);
or U25320 (N_25320,N_24528,N_24590);
xor U25321 (N_25321,N_24520,N_24953);
nor U25322 (N_25322,N_24802,N_24831);
xnor U25323 (N_25323,N_24857,N_24952);
xor U25324 (N_25324,N_24932,N_24804);
nand U25325 (N_25325,N_24981,N_24818);
or U25326 (N_25326,N_24646,N_24611);
xor U25327 (N_25327,N_24887,N_24510);
nand U25328 (N_25328,N_24645,N_24979);
xor U25329 (N_25329,N_24622,N_24827);
nand U25330 (N_25330,N_24573,N_24864);
or U25331 (N_25331,N_24934,N_24597);
nor U25332 (N_25332,N_24769,N_24776);
nor U25333 (N_25333,N_24656,N_24818);
or U25334 (N_25334,N_24738,N_24963);
or U25335 (N_25335,N_24922,N_24542);
nor U25336 (N_25336,N_24554,N_24835);
xor U25337 (N_25337,N_24643,N_24704);
nand U25338 (N_25338,N_24934,N_24736);
nor U25339 (N_25339,N_24590,N_24973);
nor U25340 (N_25340,N_24891,N_24928);
or U25341 (N_25341,N_24624,N_24994);
nand U25342 (N_25342,N_24914,N_24892);
nand U25343 (N_25343,N_24605,N_24799);
or U25344 (N_25344,N_24720,N_24660);
xor U25345 (N_25345,N_24605,N_24523);
and U25346 (N_25346,N_24665,N_24702);
nand U25347 (N_25347,N_24525,N_24909);
and U25348 (N_25348,N_24907,N_24555);
or U25349 (N_25349,N_24526,N_24982);
xnor U25350 (N_25350,N_24936,N_24883);
nor U25351 (N_25351,N_24725,N_24693);
nor U25352 (N_25352,N_24699,N_24999);
and U25353 (N_25353,N_24577,N_24624);
or U25354 (N_25354,N_24517,N_24739);
xor U25355 (N_25355,N_24584,N_24872);
or U25356 (N_25356,N_24673,N_24627);
nand U25357 (N_25357,N_24736,N_24612);
nor U25358 (N_25358,N_24653,N_24507);
nor U25359 (N_25359,N_24829,N_24933);
nand U25360 (N_25360,N_24714,N_24838);
nand U25361 (N_25361,N_24848,N_24850);
or U25362 (N_25362,N_24625,N_24556);
or U25363 (N_25363,N_24554,N_24799);
or U25364 (N_25364,N_24915,N_24717);
or U25365 (N_25365,N_24843,N_24925);
nor U25366 (N_25366,N_24991,N_24678);
xnor U25367 (N_25367,N_24693,N_24801);
nor U25368 (N_25368,N_24691,N_24552);
xnor U25369 (N_25369,N_24874,N_24588);
and U25370 (N_25370,N_24751,N_24806);
and U25371 (N_25371,N_24649,N_24694);
xor U25372 (N_25372,N_24574,N_24661);
xor U25373 (N_25373,N_24996,N_24863);
xnor U25374 (N_25374,N_24624,N_24556);
or U25375 (N_25375,N_24518,N_24808);
and U25376 (N_25376,N_24576,N_24572);
nor U25377 (N_25377,N_24767,N_24733);
and U25378 (N_25378,N_24891,N_24987);
nand U25379 (N_25379,N_24744,N_24827);
xnor U25380 (N_25380,N_24977,N_24648);
or U25381 (N_25381,N_24808,N_24881);
xor U25382 (N_25382,N_24890,N_24742);
nand U25383 (N_25383,N_24938,N_24767);
xnor U25384 (N_25384,N_24707,N_24632);
nor U25385 (N_25385,N_24760,N_24502);
nand U25386 (N_25386,N_24545,N_24624);
or U25387 (N_25387,N_24672,N_24849);
nor U25388 (N_25388,N_24802,N_24562);
and U25389 (N_25389,N_24888,N_24977);
and U25390 (N_25390,N_24919,N_24634);
or U25391 (N_25391,N_24536,N_24634);
nand U25392 (N_25392,N_24873,N_24583);
nand U25393 (N_25393,N_24758,N_24952);
nor U25394 (N_25394,N_24689,N_24653);
nor U25395 (N_25395,N_24929,N_24638);
or U25396 (N_25396,N_24957,N_24676);
nor U25397 (N_25397,N_24814,N_24607);
or U25398 (N_25398,N_24875,N_24666);
and U25399 (N_25399,N_24772,N_24738);
xnor U25400 (N_25400,N_24966,N_24614);
or U25401 (N_25401,N_24844,N_24622);
nor U25402 (N_25402,N_24740,N_24707);
nand U25403 (N_25403,N_24752,N_24591);
nand U25404 (N_25404,N_24653,N_24761);
or U25405 (N_25405,N_24810,N_24551);
xor U25406 (N_25406,N_24911,N_24715);
nand U25407 (N_25407,N_24743,N_24625);
and U25408 (N_25408,N_24564,N_24865);
nor U25409 (N_25409,N_24550,N_24789);
xor U25410 (N_25410,N_24906,N_24780);
or U25411 (N_25411,N_24712,N_24709);
nor U25412 (N_25412,N_24978,N_24506);
or U25413 (N_25413,N_24634,N_24531);
nor U25414 (N_25414,N_24626,N_24541);
nand U25415 (N_25415,N_24627,N_24761);
or U25416 (N_25416,N_24614,N_24696);
xnor U25417 (N_25417,N_24697,N_24513);
xor U25418 (N_25418,N_24935,N_24551);
and U25419 (N_25419,N_24783,N_24570);
nand U25420 (N_25420,N_24994,N_24957);
nor U25421 (N_25421,N_24800,N_24812);
nand U25422 (N_25422,N_24798,N_24736);
xor U25423 (N_25423,N_24820,N_24897);
xnor U25424 (N_25424,N_24825,N_24847);
nor U25425 (N_25425,N_24802,N_24615);
nand U25426 (N_25426,N_24966,N_24643);
nor U25427 (N_25427,N_24572,N_24536);
and U25428 (N_25428,N_24817,N_24882);
xnor U25429 (N_25429,N_24889,N_24848);
nand U25430 (N_25430,N_24828,N_24680);
nand U25431 (N_25431,N_24726,N_24895);
and U25432 (N_25432,N_24940,N_24569);
and U25433 (N_25433,N_24856,N_24790);
nand U25434 (N_25434,N_24585,N_24989);
and U25435 (N_25435,N_24650,N_24894);
nand U25436 (N_25436,N_24566,N_24660);
nor U25437 (N_25437,N_24640,N_24750);
xnor U25438 (N_25438,N_24587,N_24832);
nand U25439 (N_25439,N_24523,N_24916);
nand U25440 (N_25440,N_24756,N_24590);
nor U25441 (N_25441,N_24732,N_24550);
xnor U25442 (N_25442,N_24823,N_24962);
nor U25443 (N_25443,N_24957,N_24893);
nor U25444 (N_25444,N_24530,N_24685);
and U25445 (N_25445,N_24806,N_24595);
xnor U25446 (N_25446,N_24674,N_24767);
nand U25447 (N_25447,N_24866,N_24648);
xnor U25448 (N_25448,N_24740,N_24659);
nor U25449 (N_25449,N_24866,N_24635);
or U25450 (N_25450,N_24699,N_24719);
nor U25451 (N_25451,N_24681,N_24848);
and U25452 (N_25452,N_24964,N_24931);
nand U25453 (N_25453,N_24653,N_24786);
nand U25454 (N_25454,N_24566,N_24883);
or U25455 (N_25455,N_24664,N_24786);
and U25456 (N_25456,N_24607,N_24846);
nor U25457 (N_25457,N_24559,N_24843);
or U25458 (N_25458,N_24644,N_24825);
or U25459 (N_25459,N_24935,N_24783);
xor U25460 (N_25460,N_24556,N_24867);
nor U25461 (N_25461,N_24680,N_24872);
nand U25462 (N_25462,N_24806,N_24858);
and U25463 (N_25463,N_24869,N_24958);
xor U25464 (N_25464,N_24720,N_24696);
or U25465 (N_25465,N_24743,N_24852);
nor U25466 (N_25466,N_24710,N_24904);
nand U25467 (N_25467,N_24600,N_24915);
xor U25468 (N_25468,N_24954,N_24717);
xor U25469 (N_25469,N_24781,N_24585);
xnor U25470 (N_25470,N_24548,N_24514);
nor U25471 (N_25471,N_24806,N_24813);
nand U25472 (N_25472,N_24803,N_24547);
or U25473 (N_25473,N_24793,N_24830);
nor U25474 (N_25474,N_24933,N_24559);
nand U25475 (N_25475,N_24805,N_24506);
xnor U25476 (N_25476,N_24876,N_24782);
nand U25477 (N_25477,N_24954,N_24550);
xor U25478 (N_25478,N_24692,N_24543);
xor U25479 (N_25479,N_24983,N_24798);
nor U25480 (N_25480,N_24999,N_24735);
xor U25481 (N_25481,N_24624,N_24714);
xor U25482 (N_25482,N_24646,N_24545);
or U25483 (N_25483,N_24934,N_24697);
nand U25484 (N_25484,N_24549,N_24858);
xnor U25485 (N_25485,N_24588,N_24880);
and U25486 (N_25486,N_24705,N_24620);
or U25487 (N_25487,N_24965,N_24515);
or U25488 (N_25488,N_24531,N_24670);
nand U25489 (N_25489,N_24739,N_24650);
and U25490 (N_25490,N_24652,N_24608);
nor U25491 (N_25491,N_24687,N_24692);
and U25492 (N_25492,N_24510,N_24856);
and U25493 (N_25493,N_24556,N_24529);
nor U25494 (N_25494,N_24556,N_24692);
nand U25495 (N_25495,N_24879,N_24930);
and U25496 (N_25496,N_24678,N_24941);
or U25497 (N_25497,N_24839,N_24692);
xnor U25498 (N_25498,N_24556,N_24672);
and U25499 (N_25499,N_24825,N_24633);
nand U25500 (N_25500,N_25490,N_25059);
xor U25501 (N_25501,N_25141,N_25224);
nor U25502 (N_25502,N_25152,N_25169);
nand U25503 (N_25503,N_25032,N_25303);
nor U25504 (N_25504,N_25351,N_25387);
xor U25505 (N_25505,N_25261,N_25321);
or U25506 (N_25506,N_25063,N_25019);
or U25507 (N_25507,N_25113,N_25349);
nor U25508 (N_25508,N_25455,N_25146);
nor U25509 (N_25509,N_25177,N_25083);
nor U25510 (N_25510,N_25134,N_25309);
nand U25511 (N_25511,N_25470,N_25363);
nor U25512 (N_25512,N_25244,N_25068);
xnor U25513 (N_25513,N_25208,N_25413);
or U25514 (N_25514,N_25373,N_25317);
or U25515 (N_25515,N_25442,N_25258);
nand U25516 (N_25516,N_25437,N_25415);
or U25517 (N_25517,N_25078,N_25478);
nand U25518 (N_25518,N_25306,N_25012);
nor U25519 (N_25519,N_25198,N_25411);
and U25520 (N_25520,N_25154,N_25376);
nand U25521 (N_25521,N_25060,N_25421);
xnor U25522 (N_25522,N_25372,N_25052);
nor U25523 (N_25523,N_25420,N_25294);
or U25524 (N_25524,N_25395,N_25170);
nor U25525 (N_25525,N_25162,N_25316);
or U25526 (N_25526,N_25220,N_25180);
or U25527 (N_25527,N_25089,N_25394);
and U25528 (N_25528,N_25211,N_25359);
or U25529 (N_25529,N_25353,N_25160);
nor U25530 (N_25530,N_25453,N_25048);
xor U25531 (N_25531,N_25054,N_25174);
nor U25532 (N_25532,N_25493,N_25179);
nand U25533 (N_25533,N_25219,N_25138);
nand U25534 (N_25534,N_25031,N_25489);
or U25535 (N_25535,N_25035,N_25272);
xor U25536 (N_25536,N_25188,N_25456);
and U25537 (N_25537,N_25221,N_25315);
xor U25538 (N_25538,N_25002,N_25466);
xnor U25539 (N_25539,N_25357,N_25304);
nor U25540 (N_25540,N_25235,N_25283);
xnor U25541 (N_25541,N_25055,N_25150);
and U25542 (N_25542,N_25229,N_25369);
or U25543 (N_25543,N_25405,N_25278);
or U25544 (N_25544,N_25013,N_25097);
xnor U25545 (N_25545,N_25492,N_25178);
xnor U25546 (N_25546,N_25117,N_25046);
xor U25547 (N_25547,N_25393,N_25092);
nor U25548 (N_25548,N_25151,N_25223);
and U25549 (N_25549,N_25191,N_25355);
or U25550 (N_25550,N_25389,N_25416);
nand U25551 (N_25551,N_25064,N_25039);
and U25552 (N_25552,N_25201,N_25287);
nand U25553 (N_25553,N_25047,N_25265);
xor U25554 (N_25554,N_25481,N_25105);
nor U25555 (N_25555,N_25330,N_25079);
xor U25556 (N_25556,N_25127,N_25368);
or U25557 (N_25557,N_25062,N_25307);
nor U25558 (N_25558,N_25488,N_25263);
and U25559 (N_25559,N_25271,N_25435);
and U25560 (N_25560,N_25439,N_25408);
nor U25561 (N_25561,N_25095,N_25377);
and U25562 (N_25562,N_25467,N_25018);
nor U25563 (N_25563,N_25218,N_25473);
nor U25564 (N_25564,N_25232,N_25338);
or U25565 (N_25565,N_25298,N_25014);
and U25566 (N_25566,N_25121,N_25257);
nor U25567 (N_25567,N_25238,N_25122);
and U25568 (N_25568,N_25192,N_25017);
or U25569 (N_25569,N_25418,N_25495);
and U25570 (N_25570,N_25143,N_25450);
nand U25571 (N_25571,N_25049,N_25277);
xor U25572 (N_25572,N_25427,N_25231);
xnor U25573 (N_25573,N_25148,N_25163);
xnor U25574 (N_25574,N_25248,N_25392);
and U25575 (N_25575,N_25390,N_25010);
or U25576 (N_25576,N_25431,N_25292);
or U25577 (N_25577,N_25157,N_25400);
xor U25578 (N_25578,N_25071,N_25254);
and U25579 (N_25579,N_25006,N_25274);
and U25580 (N_25580,N_25436,N_25434);
or U25581 (N_25581,N_25284,N_25098);
or U25582 (N_25582,N_25104,N_25356);
nand U25583 (N_25583,N_25381,N_25159);
and U25584 (N_25584,N_25275,N_25397);
nor U25585 (N_25585,N_25494,N_25202);
nor U25586 (N_25586,N_25074,N_25118);
xor U25587 (N_25587,N_25135,N_25056);
or U25588 (N_25588,N_25133,N_25332);
xnor U25589 (N_25589,N_25313,N_25172);
and U25590 (N_25590,N_25214,N_25227);
nor U25591 (N_25591,N_25026,N_25126);
and U25592 (N_25592,N_25086,N_25499);
and U25593 (N_25593,N_25199,N_25156);
nor U25594 (N_25594,N_25209,N_25008);
and U25595 (N_25595,N_25479,N_25354);
nand U25596 (N_25596,N_25385,N_25016);
or U25597 (N_25597,N_25144,N_25342);
and U25598 (N_25598,N_25419,N_25096);
nor U25599 (N_25599,N_25398,N_25058);
or U25600 (N_25600,N_25197,N_25324);
xor U25601 (N_25601,N_25230,N_25023);
xor U25602 (N_25602,N_25361,N_25477);
or U25603 (N_25603,N_25237,N_25391);
xor U25604 (N_25604,N_25430,N_25422);
and U25605 (N_25605,N_25036,N_25123);
xor U25606 (N_25606,N_25260,N_25399);
xnor U25607 (N_25607,N_25075,N_25102);
nor U25608 (N_25608,N_25358,N_25498);
nor U25609 (N_25609,N_25140,N_25320);
xnor U25610 (N_25610,N_25383,N_25417);
nor U25611 (N_25611,N_25034,N_25448);
and U25612 (N_25612,N_25491,N_25388);
xnor U25613 (N_25613,N_25094,N_25067);
nand U25614 (N_25614,N_25040,N_25299);
nor U25615 (N_25615,N_25020,N_25297);
nor U25616 (N_25616,N_25329,N_25279);
nand U25617 (N_25617,N_25291,N_25210);
or U25618 (N_25618,N_25186,N_25091);
and U25619 (N_25619,N_25382,N_25243);
xnor U25620 (N_25620,N_25264,N_25312);
nand U25621 (N_25621,N_25001,N_25241);
or U25622 (N_25622,N_25190,N_25166);
nor U25623 (N_25623,N_25308,N_25472);
nand U25624 (N_25624,N_25362,N_25222);
nand U25625 (N_25625,N_25195,N_25348);
or U25626 (N_25626,N_25167,N_25273);
nand U25627 (N_25627,N_25424,N_25480);
and U25628 (N_25628,N_25423,N_25245);
or U25629 (N_25629,N_25037,N_25249);
nor U25630 (N_25630,N_25425,N_25099);
nand U25631 (N_25631,N_25136,N_25027);
and U25632 (N_25632,N_25125,N_25289);
and U25633 (N_25633,N_25240,N_25438);
xor U25634 (N_25634,N_25485,N_25267);
or U25635 (N_25635,N_25404,N_25236);
or U25636 (N_25636,N_25280,N_25137);
or U25637 (N_25637,N_25459,N_25318);
and U25638 (N_25638,N_25295,N_25153);
xor U25639 (N_25639,N_25009,N_25203);
xor U25640 (N_25640,N_25290,N_25461);
or U25641 (N_25641,N_25270,N_25196);
nor U25642 (N_25642,N_25088,N_25446);
nor U25643 (N_25643,N_25449,N_25110);
xnor U25644 (N_25644,N_25452,N_25403);
nand U25645 (N_25645,N_25412,N_25084);
or U25646 (N_25646,N_25288,N_25454);
nand U25647 (N_25647,N_25407,N_25182);
xor U25648 (N_25648,N_25057,N_25004);
nand U25649 (N_25649,N_25130,N_25396);
or U25650 (N_25650,N_25073,N_25111);
nand U25651 (N_25651,N_25327,N_25352);
and U25652 (N_25652,N_25128,N_25380);
nor U25653 (N_25653,N_25370,N_25061);
or U25654 (N_25654,N_25041,N_25168);
nor U25655 (N_25655,N_25462,N_25410);
nand U25656 (N_25656,N_25319,N_25011);
or U25657 (N_25657,N_25256,N_25246);
nor U25658 (N_25658,N_25340,N_25124);
nor U25659 (N_25659,N_25255,N_25213);
nor U25660 (N_25660,N_25259,N_25486);
or U25661 (N_25661,N_25149,N_25193);
or U25662 (N_25662,N_25365,N_25028);
nor U25663 (N_25663,N_25326,N_25266);
or U25664 (N_25664,N_25476,N_25051);
and U25665 (N_25665,N_25253,N_25468);
and U25666 (N_25666,N_25482,N_25050);
xnor U25667 (N_25667,N_25072,N_25497);
and U25668 (N_25668,N_25090,N_25015);
and U25669 (N_25669,N_25234,N_25401);
nor U25670 (N_25670,N_25483,N_25311);
xor U25671 (N_25671,N_25005,N_25145);
nor U25672 (N_25672,N_25087,N_25030);
or U25673 (N_25673,N_25451,N_25206);
xor U25674 (N_25674,N_25331,N_25043);
nand U25675 (N_25675,N_25286,N_25333);
and U25676 (N_25676,N_25367,N_25189);
xnor U25677 (N_25677,N_25334,N_25469);
xor U25678 (N_25678,N_25100,N_25029);
nor U25679 (N_25679,N_25252,N_25108);
xor U25680 (N_25680,N_25250,N_25428);
nand U25681 (N_25681,N_25165,N_25360);
xnor U25682 (N_25682,N_25426,N_25239);
and U25683 (N_25683,N_25042,N_25132);
nand U25684 (N_25684,N_25336,N_25457);
xor U25685 (N_25685,N_25347,N_25185);
or U25686 (N_25686,N_25345,N_25033);
nor U25687 (N_25687,N_25021,N_25053);
nand U25688 (N_25688,N_25375,N_25378);
nor U25689 (N_25689,N_25080,N_25107);
nand U25690 (N_25690,N_25346,N_25475);
xor U25691 (N_25691,N_25215,N_25268);
or U25692 (N_25692,N_25205,N_25337);
or U25693 (N_25693,N_25176,N_25003);
and U25694 (N_25694,N_25296,N_25300);
nor U25695 (N_25695,N_25000,N_25460);
or U25696 (N_25696,N_25458,N_25322);
or U25697 (N_25697,N_25444,N_25226);
or U25698 (N_25698,N_25155,N_25301);
nand U25699 (N_25699,N_25386,N_25171);
xnor U25700 (N_25700,N_25371,N_25173);
xnor U25701 (N_25701,N_25487,N_25175);
nand U25702 (N_25702,N_25463,N_25164);
and U25703 (N_25703,N_25341,N_25474);
or U25704 (N_25704,N_25187,N_25207);
xor U25705 (N_25705,N_25120,N_25070);
or U25706 (N_25706,N_25409,N_25158);
and U25707 (N_25707,N_25082,N_25445);
nand U25708 (N_25708,N_25414,N_25093);
and U25709 (N_25709,N_25194,N_25429);
nand U25710 (N_25710,N_25496,N_25216);
nand U25711 (N_25711,N_25022,N_25465);
nor U25712 (N_25712,N_25247,N_25112);
nand U25713 (N_25713,N_25302,N_25106);
nor U25714 (N_25714,N_25262,N_25384);
xor U25715 (N_25715,N_25379,N_25116);
xor U25716 (N_25716,N_25131,N_25007);
and U25717 (N_25717,N_25184,N_25471);
xor U25718 (N_25718,N_25081,N_25103);
or U25719 (N_25719,N_25305,N_25077);
nand U25720 (N_25720,N_25281,N_25228);
nor U25721 (N_25721,N_25285,N_25441);
nor U25722 (N_25722,N_25310,N_25343);
nand U25723 (N_25723,N_25484,N_25119);
and U25724 (N_25724,N_25076,N_25366);
nor U25725 (N_25725,N_25025,N_25129);
nand U25726 (N_25726,N_25350,N_25440);
and U25727 (N_25727,N_25364,N_25045);
nor U25728 (N_25728,N_25325,N_25024);
xor U25729 (N_25729,N_25269,N_25443);
and U25730 (N_25730,N_25339,N_25161);
nor U25731 (N_25731,N_25464,N_25114);
xor U25732 (N_25732,N_25406,N_25044);
nand U25733 (N_25733,N_25276,N_25183);
xnor U25734 (N_25734,N_25323,N_25109);
or U25735 (N_25735,N_25242,N_25447);
xor U25736 (N_25736,N_25433,N_25225);
and U25737 (N_25737,N_25065,N_25217);
nand U25738 (N_25738,N_25432,N_25212);
nand U25739 (N_25739,N_25282,N_25115);
and U25740 (N_25740,N_25085,N_25374);
nor U25741 (N_25741,N_25038,N_25293);
nand U25742 (N_25742,N_25181,N_25251);
nand U25743 (N_25743,N_25344,N_25233);
or U25744 (N_25744,N_25147,N_25142);
nand U25745 (N_25745,N_25335,N_25066);
nor U25746 (N_25746,N_25101,N_25328);
and U25747 (N_25747,N_25069,N_25139);
or U25748 (N_25748,N_25314,N_25200);
nor U25749 (N_25749,N_25204,N_25402);
and U25750 (N_25750,N_25430,N_25398);
nand U25751 (N_25751,N_25341,N_25162);
xnor U25752 (N_25752,N_25375,N_25481);
or U25753 (N_25753,N_25305,N_25252);
nor U25754 (N_25754,N_25171,N_25132);
xnor U25755 (N_25755,N_25179,N_25337);
xnor U25756 (N_25756,N_25454,N_25270);
nand U25757 (N_25757,N_25342,N_25414);
xnor U25758 (N_25758,N_25276,N_25184);
or U25759 (N_25759,N_25041,N_25255);
xor U25760 (N_25760,N_25183,N_25158);
or U25761 (N_25761,N_25320,N_25231);
or U25762 (N_25762,N_25104,N_25347);
or U25763 (N_25763,N_25385,N_25366);
nand U25764 (N_25764,N_25232,N_25226);
and U25765 (N_25765,N_25238,N_25214);
and U25766 (N_25766,N_25414,N_25128);
or U25767 (N_25767,N_25037,N_25142);
xor U25768 (N_25768,N_25029,N_25431);
nand U25769 (N_25769,N_25260,N_25265);
xor U25770 (N_25770,N_25305,N_25232);
xnor U25771 (N_25771,N_25067,N_25032);
xor U25772 (N_25772,N_25380,N_25458);
and U25773 (N_25773,N_25238,N_25146);
nor U25774 (N_25774,N_25103,N_25349);
xor U25775 (N_25775,N_25130,N_25304);
or U25776 (N_25776,N_25382,N_25165);
or U25777 (N_25777,N_25161,N_25063);
nor U25778 (N_25778,N_25175,N_25280);
nand U25779 (N_25779,N_25286,N_25398);
xor U25780 (N_25780,N_25224,N_25468);
nand U25781 (N_25781,N_25247,N_25040);
nand U25782 (N_25782,N_25250,N_25238);
xnor U25783 (N_25783,N_25431,N_25389);
and U25784 (N_25784,N_25143,N_25150);
xor U25785 (N_25785,N_25161,N_25227);
nor U25786 (N_25786,N_25112,N_25012);
xnor U25787 (N_25787,N_25497,N_25309);
or U25788 (N_25788,N_25007,N_25397);
and U25789 (N_25789,N_25061,N_25011);
nand U25790 (N_25790,N_25302,N_25246);
xor U25791 (N_25791,N_25050,N_25332);
or U25792 (N_25792,N_25340,N_25157);
nand U25793 (N_25793,N_25213,N_25366);
nor U25794 (N_25794,N_25239,N_25386);
and U25795 (N_25795,N_25257,N_25324);
nor U25796 (N_25796,N_25002,N_25157);
nand U25797 (N_25797,N_25318,N_25089);
xnor U25798 (N_25798,N_25137,N_25368);
nor U25799 (N_25799,N_25169,N_25029);
nand U25800 (N_25800,N_25350,N_25267);
xnor U25801 (N_25801,N_25388,N_25438);
and U25802 (N_25802,N_25102,N_25223);
xnor U25803 (N_25803,N_25243,N_25472);
nand U25804 (N_25804,N_25357,N_25334);
and U25805 (N_25805,N_25478,N_25103);
xor U25806 (N_25806,N_25021,N_25246);
or U25807 (N_25807,N_25066,N_25065);
and U25808 (N_25808,N_25457,N_25305);
nor U25809 (N_25809,N_25129,N_25493);
nand U25810 (N_25810,N_25151,N_25056);
or U25811 (N_25811,N_25487,N_25252);
and U25812 (N_25812,N_25245,N_25405);
nor U25813 (N_25813,N_25073,N_25356);
or U25814 (N_25814,N_25364,N_25269);
xnor U25815 (N_25815,N_25330,N_25108);
nor U25816 (N_25816,N_25152,N_25025);
nor U25817 (N_25817,N_25067,N_25063);
and U25818 (N_25818,N_25339,N_25333);
nand U25819 (N_25819,N_25083,N_25432);
or U25820 (N_25820,N_25456,N_25242);
and U25821 (N_25821,N_25014,N_25459);
or U25822 (N_25822,N_25362,N_25406);
nor U25823 (N_25823,N_25431,N_25026);
and U25824 (N_25824,N_25142,N_25054);
or U25825 (N_25825,N_25160,N_25085);
nor U25826 (N_25826,N_25396,N_25252);
or U25827 (N_25827,N_25152,N_25058);
nand U25828 (N_25828,N_25177,N_25117);
xnor U25829 (N_25829,N_25220,N_25493);
nand U25830 (N_25830,N_25373,N_25078);
nor U25831 (N_25831,N_25005,N_25338);
xnor U25832 (N_25832,N_25286,N_25266);
and U25833 (N_25833,N_25089,N_25489);
nand U25834 (N_25834,N_25139,N_25010);
nand U25835 (N_25835,N_25186,N_25295);
nand U25836 (N_25836,N_25346,N_25255);
or U25837 (N_25837,N_25215,N_25211);
nor U25838 (N_25838,N_25172,N_25088);
nor U25839 (N_25839,N_25072,N_25154);
nand U25840 (N_25840,N_25375,N_25295);
or U25841 (N_25841,N_25080,N_25029);
and U25842 (N_25842,N_25257,N_25298);
or U25843 (N_25843,N_25461,N_25368);
and U25844 (N_25844,N_25329,N_25152);
and U25845 (N_25845,N_25459,N_25267);
xnor U25846 (N_25846,N_25253,N_25289);
xor U25847 (N_25847,N_25171,N_25362);
and U25848 (N_25848,N_25049,N_25342);
nand U25849 (N_25849,N_25051,N_25055);
or U25850 (N_25850,N_25270,N_25491);
or U25851 (N_25851,N_25001,N_25123);
or U25852 (N_25852,N_25062,N_25496);
nand U25853 (N_25853,N_25141,N_25388);
and U25854 (N_25854,N_25193,N_25109);
nor U25855 (N_25855,N_25424,N_25171);
xnor U25856 (N_25856,N_25304,N_25101);
nor U25857 (N_25857,N_25059,N_25376);
and U25858 (N_25858,N_25326,N_25053);
nor U25859 (N_25859,N_25057,N_25386);
xor U25860 (N_25860,N_25009,N_25394);
nor U25861 (N_25861,N_25094,N_25278);
nand U25862 (N_25862,N_25020,N_25003);
and U25863 (N_25863,N_25152,N_25097);
nor U25864 (N_25864,N_25452,N_25418);
nor U25865 (N_25865,N_25280,N_25325);
or U25866 (N_25866,N_25316,N_25154);
nor U25867 (N_25867,N_25141,N_25341);
and U25868 (N_25868,N_25184,N_25233);
and U25869 (N_25869,N_25338,N_25184);
or U25870 (N_25870,N_25357,N_25204);
nand U25871 (N_25871,N_25095,N_25435);
xor U25872 (N_25872,N_25172,N_25352);
nor U25873 (N_25873,N_25021,N_25206);
and U25874 (N_25874,N_25046,N_25080);
xor U25875 (N_25875,N_25171,N_25043);
and U25876 (N_25876,N_25465,N_25178);
and U25877 (N_25877,N_25356,N_25352);
nand U25878 (N_25878,N_25431,N_25359);
or U25879 (N_25879,N_25407,N_25012);
or U25880 (N_25880,N_25122,N_25357);
and U25881 (N_25881,N_25005,N_25464);
and U25882 (N_25882,N_25038,N_25481);
xor U25883 (N_25883,N_25124,N_25020);
and U25884 (N_25884,N_25145,N_25274);
and U25885 (N_25885,N_25304,N_25389);
or U25886 (N_25886,N_25075,N_25025);
or U25887 (N_25887,N_25497,N_25108);
nor U25888 (N_25888,N_25076,N_25104);
xnor U25889 (N_25889,N_25423,N_25163);
and U25890 (N_25890,N_25141,N_25175);
nand U25891 (N_25891,N_25245,N_25250);
or U25892 (N_25892,N_25103,N_25367);
xnor U25893 (N_25893,N_25405,N_25069);
or U25894 (N_25894,N_25098,N_25304);
nand U25895 (N_25895,N_25108,N_25220);
xor U25896 (N_25896,N_25497,N_25371);
and U25897 (N_25897,N_25083,N_25315);
or U25898 (N_25898,N_25011,N_25312);
xnor U25899 (N_25899,N_25310,N_25042);
and U25900 (N_25900,N_25115,N_25492);
or U25901 (N_25901,N_25354,N_25076);
and U25902 (N_25902,N_25185,N_25281);
xnor U25903 (N_25903,N_25178,N_25466);
xnor U25904 (N_25904,N_25316,N_25376);
nand U25905 (N_25905,N_25375,N_25416);
or U25906 (N_25906,N_25108,N_25119);
or U25907 (N_25907,N_25094,N_25429);
nand U25908 (N_25908,N_25401,N_25326);
nand U25909 (N_25909,N_25303,N_25287);
or U25910 (N_25910,N_25316,N_25482);
xnor U25911 (N_25911,N_25230,N_25337);
nand U25912 (N_25912,N_25362,N_25363);
and U25913 (N_25913,N_25098,N_25076);
and U25914 (N_25914,N_25271,N_25014);
or U25915 (N_25915,N_25166,N_25266);
xor U25916 (N_25916,N_25101,N_25400);
nand U25917 (N_25917,N_25493,N_25459);
or U25918 (N_25918,N_25360,N_25241);
xnor U25919 (N_25919,N_25083,N_25449);
nand U25920 (N_25920,N_25157,N_25067);
xnor U25921 (N_25921,N_25406,N_25483);
nor U25922 (N_25922,N_25167,N_25136);
nor U25923 (N_25923,N_25002,N_25478);
xor U25924 (N_25924,N_25363,N_25312);
nor U25925 (N_25925,N_25120,N_25128);
nor U25926 (N_25926,N_25179,N_25248);
xor U25927 (N_25927,N_25322,N_25095);
nand U25928 (N_25928,N_25431,N_25307);
and U25929 (N_25929,N_25165,N_25239);
nand U25930 (N_25930,N_25131,N_25265);
and U25931 (N_25931,N_25116,N_25246);
nand U25932 (N_25932,N_25443,N_25010);
nand U25933 (N_25933,N_25409,N_25273);
or U25934 (N_25934,N_25285,N_25357);
or U25935 (N_25935,N_25032,N_25157);
and U25936 (N_25936,N_25477,N_25335);
nor U25937 (N_25937,N_25153,N_25193);
nor U25938 (N_25938,N_25087,N_25052);
or U25939 (N_25939,N_25447,N_25213);
nor U25940 (N_25940,N_25090,N_25328);
nand U25941 (N_25941,N_25426,N_25268);
nand U25942 (N_25942,N_25458,N_25082);
nand U25943 (N_25943,N_25000,N_25280);
nand U25944 (N_25944,N_25361,N_25098);
and U25945 (N_25945,N_25001,N_25294);
nand U25946 (N_25946,N_25323,N_25217);
nand U25947 (N_25947,N_25353,N_25300);
nor U25948 (N_25948,N_25054,N_25186);
or U25949 (N_25949,N_25292,N_25236);
and U25950 (N_25950,N_25291,N_25112);
and U25951 (N_25951,N_25429,N_25087);
nor U25952 (N_25952,N_25293,N_25145);
or U25953 (N_25953,N_25327,N_25180);
xor U25954 (N_25954,N_25201,N_25133);
and U25955 (N_25955,N_25324,N_25006);
or U25956 (N_25956,N_25314,N_25309);
and U25957 (N_25957,N_25263,N_25272);
or U25958 (N_25958,N_25447,N_25156);
xnor U25959 (N_25959,N_25408,N_25425);
xnor U25960 (N_25960,N_25420,N_25256);
nor U25961 (N_25961,N_25037,N_25329);
nand U25962 (N_25962,N_25049,N_25098);
and U25963 (N_25963,N_25291,N_25168);
nor U25964 (N_25964,N_25442,N_25421);
nand U25965 (N_25965,N_25028,N_25368);
xnor U25966 (N_25966,N_25049,N_25033);
xnor U25967 (N_25967,N_25225,N_25073);
or U25968 (N_25968,N_25097,N_25398);
xor U25969 (N_25969,N_25219,N_25495);
nor U25970 (N_25970,N_25273,N_25473);
or U25971 (N_25971,N_25204,N_25441);
nand U25972 (N_25972,N_25393,N_25413);
and U25973 (N_25973,N_25302,N_25172);
nand U25974 (N_25974,N_25458,N_25176);
nor U25975 (N_25975,N_25365,N_25429);
nor U25976 (N_25976,N_25335,N_25177);
or U25977 (N_25977,N_25287,N_25143);
and U25978 (N_25978,N_25379,N_25305);
or U25979 (N_25979,N_25407,N_25242);
nand U25980 (N_25980,N_25119,N_25282);
or U25981 (N_25981,N_25264,N_25096);
and U25982 (N_25982,N_25095,N_25102);
nand U25983 (N_25983,N_25491,N_25463);
or U25984 (N_25984,N_25033,N_25118);
nand U25985 (N_25985,N_25458,N_25498);
nand U25986 (N_25986,N_25469,N_25432);
nor U25987 (N_25987,N_25211,N_25472);
xor U25988 (N_25988,N_25111,N_25018);
xnor U25989 (N_25989,N_25302,N_25364);
nand U25990 (N_25990,N_25411,N_25496);
nor U25991 (N_25991,N_25198,N_25306);
nand U25992 (N_25992,N_25374,N_25448);
nor U25993 (N_25993,N_25168,N_25351);
xor U25994 (N_25994,N_25363,N_25290);
or U25995 (N_25995,N_25359,N_25360);
and U25996 (N_25996,N_25010,N_25484);
and U25997 (N_25997,N_25136,N_25403);
nor U25998 (N_25998,N_25492,N_25453);
and U25999 (N_25999,N_25193,N_25431);
and U26000 (N_26000,N_25961,N_25805);
and U26001 (N_26001,N_25832,N_25515);
nor U26002 (N_26002,N_25762,N_25856);
and U26003 (N_26003,N_25924,N_25712);
xnor U26004 (N_26004,N_25703,N_25908);
nand U26005 (N_26005,N_25970,N_25543);
xnor U26006 (N_26006,N_25706,N_25842);
or U26007 (N_26007,N_25836,N_25707);
or U26008 (N_26008,N_25848,N_25877);
xor U26009 (N_26009,N_25993,N_25907);
or U26010 (N_26010,N_25768,N_25822);
nand U26011 (N_26011,N_25680,N_25992);
xor U26012 (N_26012,N_25675,N_25649);
and U26013 (N_26013,N_25687,N_25633);
or U26014 (N_26014,N_25904,N_25954);
or U26015 (N_26015,N_25879,N_25906);
or U26016 (N_26016,N_25532,N_25846);
or U26017 (N_26017,N_25779,N_25655);
nor U26018 (N_26018,N_25504,N_25670);
and U26019 (N_26019,N_25558,N_25641);
nand U26020 (N_26020,N_25819,N_25982);
or U26021 (N_26021,N_25895,N_25880);
nand U26022 (N_26022,N_25654,N_25894);
xor U26023 (N_26023,N_25913,N_25528);
nor U26024 (N_26024,N_25501,N_25890);
and U26025 (N_26025,N_25854,N_25696);
or U26026 (N_26026,N_25941,N_25588);
nor U26027 (N_26027,N_25682,N_25878);
xnor U26028 (N_26028,N_25853,N_25562);
nand U26029 (N_26029,N_25555,N_25778);
or U26030 (N_26030,N_25554,N_25512);
or U26031 (N_26031,N_25559,N_25591);
and U26032 (N_26032,N_25698,N_25661);
nand U26033 (N_26033,N_25803,N_25789);
xnor U26034 (N_26034,N_25615,N_25593);
xor U26035 (N_26035,N_25720,N_25817);
xor U26036 (N_26036,N_25694,N_25617);
nor U26037 (N_26037,N_25574,N_25598);
nand U26038 (N_26038,N_25724,N_25979);
or U26039 (N_26039,N_25688,N_25830);
nor U26040 (N_26040,N_25828,N_25564);
nand U26041 (N_26041,N_25807,N_25925);
nor U26042 (N_26042,N_25889,N_25810);
or U26043 (N_26043,N_25965,N_25918);
xor U26044 (N_26044,N_25699,N_25746);
and U26045 (N_26045,N_25963,N_25567);
xor U26046 (N_26046,N_25544,N_25763);
nand U26047 (N_26047,N_25530,N_25867);
xnor U26048 (N_26048,N_25935,N_25875);
xor U26049 (N_26049,N_25656,N_25891);
nor U26050 (N_26050,N_25843,N_25610);
and U26051 (N_26051,N_25708,N_25814);
or U26052 (N_26052,N_25604,N_25581);
or U26053 (N_26053,N_25785,N_25927);
xor U26054 (N_26054,N_25858,N_25769);
and U26055 (N_26055,N_25734,N_25948);
xnor U26056 (N_26056,N_25792,N_25933);
nand U26057 (N_26057,N_25804,N_25758);
nand U26058 (N_26058,N_25529,N_25825);
nand U26059 (N_26059,N_25565,N_25596);
or U26060 (N_26060,N_25851,N_25989);
nand U26061 (N_26061,N_25869,N_25956);
nor U26062 (N_26062,N_25795,N_25911);
and U26063 (N_26063,N_25909,N_25938);
nand U26064 (N_26064,N_25629,N_25626);
nor U26065 (N_26065,N_25930,N_25622);
and U26066 (N_26066,N_25630,N_25582);
nand U26067 (N_26067,N_25652,N_25981);
nor U26068 (N_26068,N_25648,N_25973);
nand U26069 (N_26069,N_25986,N_25943);
xnor U26070 (N_26070,N_25765,N_25619);
xnor U26071 (N_26071,N_25797,N_25577);
xor U26072 (N_26072,N_25841,N_25787);
xnor U26073 (N_26073,N_25600,N_25692);
nor U26074 (N_26074,N_25672,N_25944);
xor U26075 (N_26075,N_25829,N_25549);
nand U26076 (N_26076,N_25749,N_25645);
nor U26077 (N_26077,N_25627,N_25958);
and U26078 (N_26078,N_25540,N_25614);
nand U26079 (N_26079,N_25996,N_25953);
nor U26080 (N_26080,N_25662,N_25923);
and U26081 (N_26081,N_25820,N_25697);
nor U26082 (N_26082,N_25508,N_25998);
xor U26083 (N_26083,N_25527,N_25929);
or U26084 (N_26084,N_25945,N_25736);
or U26085 (N_26085,N_25994,N_25653);
or U26086 (N_26086,N_25862,N_25844);
nor U26087 (N_26087,N_25786,N_25603);
xnor U26088 (N_26088,N_25896,N_25566);
and U26089 (N_26089,N_25583,N_25521);
and U26090 (N_26090,N_25505,N_25885);
xor U26091 (N_26091,N_25545,N_25823);
nand U26092 (N_26092,N_25728,N_25731);
nand U26093 (N_26093,N_25886,N_25659);
and U26094 (N_26094,N_25678,N_25864);
and U26095 (N_26095,N_25818,N_25640);
or U26096 (N_26096,N_25753,N_25725);
nor U26097 (N_26097,N_25760,N_25937);
nand U26098 (N_26098,N_25606,N_25741);
nor U26099 (N_26099,N_25667,N_25560);
or U26100 (N_26100,N_25519,N_25681);
nand U26101 (N_26101,N_25892,N_25839);
nor U26102 (N_26102,N_25693,N_25899);
xnor U26103 (N_26103,N_25535,N_25815);
xor U26104 (N_26104,N_25538,N_25578);
nand U26105 (N_26105,N_25602,N_25548);
or U26106 (N_26106,N_25744,N_25928);
nor U26107 (N_26107,N_25557,N_25901);
and U26108 (N_26108,N_25643,N_25509);
xor U26109 (N_26109,N_25915,N_25526);
nor U26110 (N_26110,N_25638,N_25595);
and U26111 (N_26111,N_25684,N_25666);
or U26112 (N_26112,N_25912,N_25873);
and U26113 (N_26113,N_25585,N_25974);
or U26114 (N_26114,N_25639,N_25999);
and U26115 (N_26115,N_25754,N_25522);
and U26116 (N_26116,N_25533,N_25580);
and U26117 (N_26117,N_25919,N_25951);
nand U26118 (N_26118,N_25983,N_25761);
nand U26119 (N_26119,N_25556,N_25541);
or U26120 (N_26120,N_25801,N_25755);
and U26121 (N_26121,N_25613,N_25985);
or U26122 (N_26122,N_25671,N_25637);
and U26123 (N_26123,N_25914,N_25980);
nor U26124 (N_26124,N_25714,N_25863);
and U26125 (N_26125,N_25513,N_25766);
or U26126 (N_26126,N_25776,N_25686);
nor U26127 (N_26127,N_25618,N_25751);
xnor U26128 (N_26128,N_25866,N_25642);
nand U26129 (N_26129,N_25976,N_25503);
or U26130 (N_26130,N_25782,N_25722);
xnor U26131 (N_26131,N_25888,N_25920);
nand U26132 (N_26132,N_25690,N_25793);
and U26133 (N_26133,N_25516,N_25882);
or U26134 (N_26134,N_25995,N_25784);
nand U26135 (N_26135,N_25834,N_25808);
nand U26136 (N_26136,N_25546,N_25813);
xor U26137 (N_26137,N_25590,N_25972);
nand U26138 (N_26138,N_25571,N_25579);
and U26139 (N_26139,N_25936,N_25798);
xnor U26140 (N_26140,N_25931,N_25635);
nor U26141 (N_26141,N_25942,N_25676);
and U26142 (N_26142,N_25902,N_25800);
xnor U26143 (N_26143,N_25881,N_25733);
nor U26144 (N_26144,N_25838,N_25967);
nand U26145 (N_26145,N_25737,N_25771);
xnor U26146 (N_26146,N_25752,N_25791);
xnor U26147 (N_26147,N_25859,N_25732);
and U26148 (N_26148,N_25990,N_25774);
or U26149 (N_26149,N_25968,N_25845);
xnor U26150 (N_26150,N_25966,N_25991);
nor U26151 (N_26151,N_25865,N_25650);
xor U26152 (N_26152,N_25616,N_25917);
nand U26153 (N_26153,N_25940,N_25824);
nor U26154 (N_26154,N_25620,N_25647);
or U26155 (N_26155,N_25586,N_25860);
nor U26156 (N_26156,N_25644,N_25934);
nand U26157 (N_26157,N_25689,N_25589);
or U26158 (N_26158,N_25802,N_25592);
or U26159 (N_26159,N_25876,N_25921);
and U26160 (N_26160,N_25748,N_25777);
nor U26161 (N_26161,N_25975,N_25553);
and U26162 (N_26162,N_25511,N_25717);
or U26163 (N_26163,N_25947,N_25601);
nand U26164 (N_26164,N_25835,N_25514);
and U26165 (N_26165,N_25738,N_25520);
xnor U26166 (N_26166,N_25742,N_25857);
or U26167 (N_26167,N_25905,N_25796);
xor U26168 (N_26168,N_25716,N_25772);
or U26169 (N_26169,N_25922,N_25756);
nor U26170 (N_26170,N_25840,N_25628);
or U26171 (N_26171,N_25872,N_25576);
and U26172 (N_26172,N_25534,N_25887);
xnor U26173 (N_26173,N_25770,N_25568);
and U26174 (N_26174,N_25730,N_25827);
nand U26175 (N_26175,N_25539,N_25665);
and U26176 (N_26176,N_25570,N_25551);
nand U26177 (N_26177,N_25563,N_25683);
nor U26178 (N_26178,N_25898,N_25524);
nor U26179 (N_26179,N_25663,N_25855);
xnor U26180 (N_26180,N_25997,N_25542);
nand U26181 (N_26181,N_25783,N_25852);
nand U26182 (N_26182,N_25584,N_25757);
nor U26183 (N_26183,N_25893,N_25631);
xor U26184 (N_26184,N_25952,N_25646);
nand U26185 (N_26185,N_25988,N_25506);
xnor U26186 (N_26186,N_25870,N_25673);
xor U26187 (N_26187,N_25674,N_25547);
and U26188 (N_26188,N_25664,N_25572);
nand U26189 (N_26189,N_25811,N_25594);
or U26190 (N_26190,N_25525,N_25536);
nor U26191 (N_26191,N_25657,N_25704);
and U26192 (N_26192,N_25599,N_25969);
nand U26193 (N_26193,N_25719,N_25812);
xor U26194 (N_26194,N_25788,N_25569);
and U26195 (N_26195,N_25552,N_25874);
or U26196 (N_26196,N_25711,N_25621);
nor U26197 (N_26197,N_25861,N_25700);
xor U26198 (N_26198,N_25916,N_25910);
xor U26199 (N_26199,N_25971,N_25721);
nand U26200 (N_26200,N_25669,N_25850);
and U26201 (N_26201,N_25735,N_25587);
nand U26202 (N_26202,N_25960,N_25632);
nor U26203 (N_26203,N_25651,N_25950);
nor U26204 (N_26204,N_25932,N_25750);
nor U26205 (N_26205,N_25743,N_25957);
xor U26206 (N_26206,N_25561,N_25710);
nand U26207 (N_26207,N_25984,N_25691);
nand U26208 (N_26208,N_25764,N_25794);
nand U26209 (N_26209,N_25816,N_25790);
xnor U26210 (N_26210,N_25826,N_25883);
or U26211 (N_26211,N_25897,N_25962);
xnor U26212 (N_26212,N_25806,N_25668);
or U26213 (N_26213,N_25685,N_25926);
or U26214 (N_26214,N_25959,N_25903);
and U26215 (N_26215,N_25977,N_25821);
nor U26216 (N_26216,N_25660,N_25679);
nand U26217 (N_26217,N_25775,N_25739);
xor U26218 (N_26218,N_25833,N_25718);
and U26219 (N_26219,N_25726,N_25713);
and U26220 (N_26220,N_25809,N_25701);
and U26221 (N_26221,N_25955,N_25781);
nand U26222 (N_26222,N_25573,N_25518);
or U26223 (N_26223,N_25502,N_25500);
nand U26224 (N_26224,N_25507,N_25837);
or U26225 (N_26225,N_25517,N_25900);
nand U26226 (N_26226,N_25550,N_25939);
xnor U26227 (N_26227,N_25868,N_25799);
and U26228 (N_26228,N_25729,N_25624);
nor U26229 (N_26229,N_25702,N_25634);
and U26230 (N_26230,N_25597,N_25695);
xor U26231 (N_26231,N_25949,N_25523);
and U26232 (N_26232,N_25747,N_25575);
and U26233 (N_26233,N_25715,N_25607);
and U26234 (N_26234,N_25773,N_25531);
and U26235 (N_26235,N_25831,N_25964);
or U26236 (N_26236,N_25709,N_25978);
nand U26237 (N_26237,N_25608,N_25759);
or U26238 (N_26238,N_25611,N_25727);
xor U26239 (N_26239,N_25767,N_25987);
nor U26240 (N_26240,N_25946,N_25510);
nand U26241 (N_26241,N_25537,N_25723);
nand U26242 (N_26242,N_25612,N_25740);
nand U26243 (N_26243,N_25745,N_25871);
and U26244 (N_26244,N_25625,N_25658);
and U26245 (N_26245,N_25849,N_25605);
xnor U26246 (N_26246,N_25847,N_25884);
nand U26247 (N_26247,N_25780,N_25705);
or U26248 (N_26248,N_25636,N_25609);
or U26249 (N_26249,N_25623,N_25677);
and U26250 (N_26250,N_25766,N_25744);
nand U26251 (N_26251,N_25791,N_25820);
nand U26252 (N_26252,N_25603,N_25608);
or U26253 (N_26253,N_25916,N_25670);
or U26254 (N_26254,N_25824,N_25509);
or U26255 (N_26255,N_25925,N_25850);
xor U26256 (N_26256,N_25785,N_25964);
and U26257 (N_26257,N_25931,N_25662);
xnor U26258 (N_26258,N_25525,N_25760);
or U26259 (N_26259,N_25540,N_25531);
nand U26260 (N_26260,N_25591,N_25805);
nor U26261 (N_26261,N_25931,N_25598);
or U26262 (N_26262,N_25545,N_25942);
and U26263 (N_26263,N_25624,N_25732);
nor U26264 (N_26264,N_25855,N_25735);
xnor U26265 (N_26265,N_25613,N_25504);
xnor U26266 (N_26266,N_25504,N_25557);
or U26267 (N_26267,N_25950,N_25946);
or U26268 (N_26268,N_25552,N_25960);
xnor U26269 (N_26269,N_25993,N_25571);
nand U26270 (N_26270,N_25829,N_25852);
or U26271 (N_26271,N_25522,N_25944);
nand U26272 (N_26272,N_25857,N_25699);
nand U26273 (N_26273,N_25771,N_25749);
nor U26274 (N_26274,N_25778,N_25645);
or U26275 (N_26275,N_25707,N_25975);
nor U26276 (N_26276,N_25942,N_25556);
xnor U26277 (N_26277,N_25545,N_25513);
nand U26278 (N_26278,N_25895,N_25651);
xor U26279 (N_26279,N_25685,N_25553);
or U26280 (N_26280,N_25910,N_25698);
nand U26281 (N_26281,N_25780,N_25610);
or U26282 (N_26282,N_25882,N_25618);
and U26283 (N_26283,N_25757,N_25677);
nor U26284 (N_26284,N_25766,N_25763);
nand U26285 (N_26285,N_25691,N_25606);
nand U26286 (N_26286,N_25626,N_25789);
or U26287 (N_26287,N_25942,N_25869);
or U26288 (N_26288,N_25748,N_25687);
nand U26289 (N_26289,N_25527,N_25793);
nand U26290 (N_26290,N_25627,N_25845);
nand U26291 (N_26291,N_25528,N_25518);
nand U26292 (N_26292,N_25805,N_25546);
nor U26293 (N_26293,N_25856,N_25708);
xor U26294 (N_26294,N_25613,N_25589);
nand U26295 (N_26295,N_25875,N_25527);
nor U26296 (N_26296,N_25550,N_25675);
nand U26297 (N_26297,N_25530,N_25916);
or U26298 (N_26298,N_25627,N_25745);
xnor U26299 (N_26299,N_25747,N_25990);
nor U26300 (N_26300,N_25508,N_25525);
or U26301 (N_26301,N_25856,N_25728);
or U26302 (N_26302,N_25822,N_25715);
or U26303 (N_26303,N_25915,N_25765);
nor U26304 (N_26304,N_25847,N_25524);
xnor U26305 (N_26305,N_25978,N_25581);
nor U26306 (N_26306,N_25533,N_25853);
or U26307 (N_26307,N_25689,N_25606);
or U26308 (N_26308,N_25516,N_25755);
nand U26309 (N_26309,N_25545,N_25529);
or U26310 (N_26310,N_25908,N_25968);
and U26311 (N_26311,N_25885,N_25675);
nor U26312 (N_26312,N_25936,N_25826);
nor U26313 (N_26313,N_25763,N_25877);
nand U26314 (N_26314,N_25841,N_25542);
and U26315 (N_26315,N_25632,N_25834);
nand U26316 (N_26316,N_25575,N_25732);
nand U26317 (N_26317,N_25778,N_25617);
or U26318 (N_26318,N_25508,N_25952);
and U26319 (N_26319,N_25517,N_25693);
xnor U26320 (N_26320,N_25743,N_25986);
and U26321 (N_26321,N_25733,N_25702);
or U26322 (N_26322,N_25659,N_25606);
nand U26323 (N_26323,N_25667,N_25973);
nand U26324 (N_26324,N_25606,N_25904);
or U26325 (N_26325,N_25602,N_25635);
and U26326 (N_26326,N_25855,N_25620);
xor U26327 (N_26327,N_25996,N_25756);
nand U26328 (N_26328,N_25693,N_25959);
or U26329 (N_26329,N_25679,N_25942);
nor U26330 (N_26330,N_25731,N_25921);
nor U26331 (N_26331,N_25647,N_25619);
nor U26332 (N_26332,N_25561,N_25995);
and U26333 (N_26333,N_25861,N_25725);
xnor U26334 (N_26334,N_25879,N_25950);
and U26335 (N_26335,N_25691,N_25645);
and U26336 (N_26336,N_25930,N_25803);
xnor U26337 (N_26337,N_25772,N_25825);
xor U26338 (N_26338,N_25719,N_25947);
or U26339 (N_26339,N_25765,N_25879);
and U26340 (N_26340,N_25779,N_25770);
or U26341 (N_26341,N_25888,N_25696);
xor U26342 (N_26342,N_25605,N_25568);
and U26343 (N_26343,N_25793,N_25696);
and U26344 (N_26344,N_25918,N_25507);
xnor U26345 (N_26345,N_25834,N_25769);
nor U26346 (N_26346,N_25511,N_25551);
or U26347 (N_26347,N_25778,N_25877);
nand U26348 (N_26348,N_25978,N_25963);
nor U26349 (N_26349,N_25621,N_25544);
or U26350 (N_26350,N_25589,N_25855);
and U26351 (N_26351,N_25847,N_25709);
nand U26352 (N_26352,N_25704,N_25936);
or U26353 (N_26353,N_25762,N_25992);
nand U26354 (N_26354,N_25515,N_25716);
or U26355 (N_26355,N_25858,N_25703);
or U26356 (N_26356,N_25609,N_25698);
nor U26357 (N_26357,N_25899,N_25680);
nand U26358 (N_26358,N_25933,N_25670);
xor U26359 (N_26359,N_25563,N_25977);
nand U26360 (N_26360,N_25920,N_25604);
or U26361 (N_26361,N_25700,N_25830);
xnor U26362 (N_26362,N_25857,N_25991);
nor U26363 (N_26363,N_25734,N_25999);
or U26364 (N_26364,N_25634,N_25712);
nor U26365 (N_26365,N_25665,N_25994);
or U26366 (N_26366,N_25964,N_25554);
nand U26367 (N_26367,N_25638,N_25635);
nand U26368 (N_26368,N_25728,N_25582);
nor U26369 (N_26369,N_25890,N_25522);
or U26370 (N_26370,N_25796,N_25605);
nor U26371 (N_26371,N_25677,N_25938);
and U26372 (N_26372,N_25726,N_25661);
nand U26373 (N_26373,N_25790,N_25824);
or U26374 (N_26374,N_25634,N_25894);
or U26375 (N_26375,N_25860,N_25891);
xor U26376 (N_26376,N_25870,N_25862);
nor U26377 (N_26377,N_25732,N_25748);
or U26378 (N_26378,N_25830,N_25979);
and U26379 (N_26379,N_25762,N_25924);
or U26380 (N_26380,N_25638,N_25896);
nor U26381 (N_26381,N_25760,N_25576);
or U26382 (N_26382,N_25972,N_25994);
xnor U26383 (N_26383,N_25770,N_25820);
xnor U26384 (N_26384,N_25706,N_25671);
and U26385 (N_26385,N_25603,N_25650);
and U26386 (N_26386,N_25718,N_25952);
or U26387 (N_26387,N_25512,N_25750);
nand U26388 (N_26388,N_25988,N_25974);
nor U26389 (N_26389,N_25799,N_25962);
nand U26390 (N_26390,N_25861,N_25601);
and U26391 (N_26391,N_25718,N_25913);
or U26392 (N_26392,N_25869,N_25568);
and U26393 (N_26393,N_25996,N_25690);
xnor U26394 (N_26394,N_25857,N_25549);
or U26395 (N_26395,N_25740,N_25838);
nand U26396 (N_26396,N_25794,N_25598);
or U26397 (N_26397,N_25678,N_25906);
and U26398 (N_26398,N_25804,N_25898);
and U26399 (N_26399,N_25625,N_25767);
xnor U26400 (N_26400,N_25782,N_25839);
nor U26401 (N_26401,N_25601,N_25649);
xor U26402 (N_26402,N_25762,N_25504);
or U26403 (N_26403,N_25869,N_25801);
and U26404 (N_26404,N_25661,N_25851);
nor U26405 (N_26405,N_25882,N_25955);
and U26406 (N_26406,N_25785,N_25576);
or U26407 (N_26407,N_25728,N_25860);
xnor U26408 (N_26408,N_25919,N_25988);
nor U26409 (N_26409,N_25952,N_25630);
xnor U26410 (N_26410,N_25583,N_25810);
or U26411 (N_26411,N_25640,N_25783);
nor U26412 (N_26412,N_25719,N_25706);
nor U26413 (N_26413,N_25863,N_25740);
nor U26414 (N_26414,N_25813,N_25790);
and U26415 (N_26415,N_25815,N_25950);
nand U26416 (N_26416,N_25515,N_25960);
xnor U26417 (N_26417,N_25904,N_25882);
and U26418 (N_26418,N_25877,N_25874);
nor U26419 (N_26419,N_25862,N_25752);
nor U26420 (N_26420,N_25966,N_25525);
xor U26421 (N_26421,N_25807,N_25678);
nand U26422 (N_26422,N_25764,N_25976);
nand U26423 (N_26423,N_25992,N_25767);
nor U26424 (N_26424,N_25665,N_25770);
nor U26425 (N_26425,N_25831,N_25644);
nor U26426 (N_26426,N_25539,N_25832);
or U26427 (N_26427,N_25956,N_25827);
xor U26428 (N_26428,N_25831,N_25929);
or U26429 (N_26429,N_25844,N_25944);
nand U26430 (N_26430,N_25782,N_25720);
xor U26431 (N_26431,N_25915,N_25530);
or U26432 (N_26432,N_25956,N_25574);
and U26433 (N_26433,N_25642,N_25903);
nor U26434 (N_26434,N_25751,N_25536);
or U26435 (N_26435,N_25815,N_25600);
nor U26436 (N_26436,N_25736,N_25927);
and U26437 (N_26437,N_25871,N_25740);
or U26438 (N_26438,N_25961,N_25725);
xnor U26439 (N_26439,N_25564,N_25936);
xnor U26440 (N_26440,N_25574,N_25549);
nand U26441 (N_26441,N_25574,N_25954);
xnor U26442 (N_26442,N_25783,N_25907);
and U26443 (N_26443,N_25968,N_25780);
or U26444 (N_26444,N_25743,N_25917);
nor U26445 (N_26445,N_25822,N_25741);
or U26446 (N_26446,N_25856,N_25887);
and U26447 (N_26447,N_25754,N_25674);
nand U26448 (N_26448,N_25979,N_25840);
and U26449 (N_26449,N_25567,N_25843);
nor U26450 (N_26450,N_25792,N_25685);
and U26451 (N_26451,N_25582,N_25970);
nor U26452 (N_26452,N_25952,N_25773);
or U26453 (N_26453,N_25710,N_25685);
nor U26454 (N_26454,N_25747,N_25639);
xor U26455 (N_26455,N_25981,N_25856);
nand U26456 (N_26456,N_25823,N_25525);
or U26457 (N_26457,N_25861,N_25756);
or U26458 (N_26458,N_25788,N_25595);
and U26459 (N_26459,N_25851,N_25620);
nor U26460 (N_26460,N_25823,N_25704);
nor U26461 (N_26461,N_25659,N_25797);
nor U26462 (N_26462,N_25885,N_25891);
or U26463 (N_26463,N_25779,N_25901);
nor U26464 (N_26464,N_25797,N_25608);
xor U26465 (N_26465,N_25943,N_25533);
or U26466 (N_26466,N_25507,N_25597);
or U26467 (N_26467,N_25563,N_25688);
nand U26468 (N_26468,N_25790,N_25962);
nand U26469 (N_26469,N_25964,N_25647);
xor U26470 (N_26470,N_25533,N_25866);
nor U26471 (N_26471,N_25678,N_25614);
nand U26472 (N_26472,N_25740,N_25984);
and U26473 (N_26473,N_25896,N_25641);
or U26474 (N_26474,N_25560,N_25654);
and U26475 (N_26475,N_25621,N_25757);
nand U26476 (N_26476,N_25558,N_25506);
or U26477 (N_26477,N_25721,N_25743);
nand U26478 (N_26478,N_25624,N_25506);
or U26479 (N_26479,N_25906,N_25697);
nand U26480 (N_26480,N_25952,N_25665);
xnor U26481 (N_26481,N_25722,N_25824);
or U26482 (N_26482,N_25736,N_25826);
nor U26483 (N_26483,N_25718,N_25692);
nand U26484 (N_26484,N_25774,N_25747);
nand U26485 (N_26485,N_25626,N_25636);
nand U26486 (N_26486,N_25612,N_25909);
xnor U26487 (N_26487,N_25530,N_25999);
nor U26488 (N_26488,N_25690,N_25886);
nor U26489 (N_26489,N_25803,N_25938);
and U26490 (N_26490,N_25788,N_25670);
nand U26491 (N_26491,N_25564,N_25654);
nor U26492 (N_26492,N_25774,N_25717);
nor U26493 (N_26493,N_25502,N_25624);
xor U26494 (N_26494,N_25776,N_25964);
nor U26495 (N_26495,N_25757,N_25782);
nand U26496 (N_26496,N_25534,N_25676);
or U26497 (N_26497,N_25998,N_25510);
and U26498 (N_26498,N_25707,N_25671);
xor U26499 (N_26499,N_25532,N_25625);
nand U26500 (N_26500,N_26420,N_26229);
nor U26501 (N_26501,N_26172,N_26194);
and U26502 (N_26502,N_26016,N_26085);
nand U26503 (N_26503,N_26008,N_26313);
or U26504 (N_26504,N_26048,N_26222);
nor U26505 (N_26505,N_26156,N_26102);
xnor U26506 (N_26506,N_26025,N_26263);
xnor U26507 (N_26507,N_26493,N_26378);
xnor U26508 (N_26508,N_26496,N_26165);
xnor U26509 (N_26509,N_26004,N_26407);
xnor U26510 (N_26510,N_26461,N_26331);
xor U26511 (N_26511,N_26440,N_26240);
nor U26512 (N_26512,N_26435,N_26457);
or U26513 (N_26513,N_26284,N_26465);
and U26514 (N_26514,N_26302,N_26477);
nor U26515 (N_26515,N_26105,N_26178);
and U26516 (N_26516,N_26325,N_26315);
and U26517 (N_26517,N_26355,N_26221);
or U26518 (N_26518,N_26336,N_26065);
xor U26519 (N_26519,N_26140,N_26244);
nor U26520 (N_26520,N_26169,N_26013);
nand U26521 (N_26521,N_26344,N_26057);
nand U26522 (N_26522,N_26437,N_26304);
and U26523 (N_26523,N_26067,N_26359);
nor U26524 (N_26524,N_26324,N_26043);
and U26525 (N_26525,N_26494,N_26273);
and U26526 (N_26526,N_26414,N_26191);
nand U26527 (N_26527,N_26421,N_26093);
nor U26528 (N_26528,N_26342,N_26237);
nor U26529 (N_26529,N_26163,N_26151);
xor U26530 (N_26530,N_26101,N_26426);
nor U26531 (N_26531,N_26230,N_26103);
or U26532 (N_26532,N_26334,N_26022);
nand U26533 (N_26533,N_26187,N_26090);
nor U26534 (N_26534,N_26034,N_26193);
nor U26535 (N_26535,N_26285,N_26199);
xnor U26536 (N_26536,N_26363,N_26155);
nand U26537 (N_26537,N_26198,N_26417);
nand U26538 (N_26538,N_26291,N_26452);
or U26539 (N_26539,N_26394,N_26332);
nand U26540 (N_26540,N_26080,N_26039);
or U26541 (N_26541,N_26088,N_26147);
or U26542 (N_26542,N_26042,N_26097);
nor U26543 (N_26543,N_26442,N_26287);
and U26544 (N_26544,N_26021,N_26292);
xor U26545 (N_26545,N_26047,N_26033);
nor U26546 (N_26546,N_26145,N_26479);
and U26547 (N_26547,N_26390,N_26208);
nor U26548 (N_26548,N_26146,N_26252);
nor U26549 (N_26549,N_26449,N_26321);
nor U26550 (N_26550,N_26387,N_26020);
xnor U26551 (N_26551,N_26259,N_26430);
or U26552 (N_26552,N_26346,N_26214);
nor U26553 (N_26553,N_26408,N_26152);
xnor U26554 (N_26554,N_26185,N_26300);
nand U26555 (N_26555,N_26353,N_26003);
nand U26556 (N_26556,N_26403,N_26158);
nor U26557 (N_26557,N_26031,N_26148);
or U26558 (N_26558,N_26486,N_26074);
and U26559 (N_26559,N_26460,N_26436);
nor U26560 (N_26560,N_26100,N_26312);
nand U26561 (N_26561,N_26197,N_26226);
nor U26562 (N_26562,N_26162,N_26361);
or U26563 (N_26563,N_26371,N_26014);
xnor U26564 (N_26564,N_26175,N_26338);
and U26565 (N_26565,N_26410,N_26474);
or U26566 (N_26566,N_26200,N_26219);
nand U26567 (N_26567,N_26188,N_26419);
or U26568 (N_26568,N_26482,N_26468);
nand U26569 (N_26569,N_26379,N_26340);
nor U26570 (N_26570,N_26112,N_26428);
or U26571 (N_26571,N_26383,N_26083);
nor U26572 (N_26572,N_26395,N_26489);
or U26573 (N_26573,N_26012,N_26063);
and U26574 (N_26574,N_26377,N_26271);
xnor U26575 (N_26575,N_26201,N_26164);
and U26576 (N_26576,N_26433,N_26176);
nor U26577 (N_26577,N_26141,N_26231);
nand U26578 (N_26578,N_26220,N_26086);
xor U26579 (N_26579,N_26015,N_26011);
nor U26580 (N_26580,N_26356,N_26424);
or U26581 (N_26581,N_26352,N_26257);
and U26582 (N_26582,N_26351,N_26445);
or U26583 (N_26583,N_26216,N_26307);
xor U26584 (N_26584,N_26026,N_26143);
or U26585 (N_26585,N_26023,N_26217);
xnor U26586 (N_26586,N_26308,N_26125);
and U26587 (N_26587,N_26205,N_26478);
nand U26588 (N_26588,N_26471,N_26243);
nor U26589 (N_26589,N_26173,N_26157);
and U26590 (N_26590,N_26288,N_26397);
xnor U26591 (N_26591,N_26001,N_26116);
and U26592 (N_26592,N_26002,N_26398);
nor U26593 (N_26593,N_26073,N_26303);
xnor U26594 (N_26594,N_26429,N_26160);
and U26595 (N_26595,N_26076,N_26066);
nor U26596 (N_26596,N_26236,N_26062);
and U26597 (N_26597,N_26458,N_26498);
xor U26598 (N_26598,N_26211,N_26239);
and U26599 (N_26599,N_26427,N_26453);
or U26600 (N_26600,N_26079,N_26005);
xor U26601 (N_26601,N_26404,N_26225);
nor U26602 (N_26602,N_26215,N_26354);
xnor U26603 (N_26603,N_26118,N_26078);
xor U26604 (N_26604,N_26341,N_26044);
and U26605 (N_26605,N_26322,N_26451);
and U26606 (N_26606,N_26099,N_26382);
xnor U26607 (N_26607,N_26045,N_26087);
nand U26608 (N_26608,N_26444,N_26280);
xor U26609 (N_26609,N_26389,N_26174);
nand U26610 (N_26610,N_26349,N_26128);
or U26611 (N_26611,N_26446,N_26350);
and U26612 (N_26612,N_26281,N_26192);
or U26613 (N_26613,N_26159,N_26297);
nand U26614 (N_26614,N_26254,N_26117);
xnor U26615 (N_26615,N_26029,N_26268);
nand U26616 (N_26616,N_26035,N_26245);
or U26617 (N_26617,N_26272,N_26335);
xnor U26618 (N_26618,N_26058,N_26283);
nor U26619 (N_26619,N_26183,N_26372);
and U26620 (N_26620,N_26223,N_26234);
or U26621 (N_26621,N_26137,N_26463);
xor U26622 (N_26622,N_26380,N_26068);
and U26623 (N_26623,N_26092,N_26360);
nor U26624 (N_26624,N_26224,N_26119);
nand U26625 (N_26625,N_26274,N_26138);
or U26626 (N_26626,N_26434,N_26375);
or U26627 (N_26627,N_26030,N_26485);
and U26628 (N_26628,N_26111,N_26309);
nor U26629 (N_26629,N_26339,N_26399);
and U26630 (N_26630,N_26469,N_26053);
xnor U26631 (N_26631,N_26258,N_26209);
xnor U26632 (N_26632,N_26110,N_26054);
and U26633 (N_26633,N_26385,N_26497);
nand U26634 (N_26634,N_26368,N_26488);
or U26635 (N_26635,N_26282,N_26362);
and U26636 (N_26636,N_26171,N_26327);
and U26637 (N_26637,N_26052,N_26367);
nor U26638 (N_26638,N_26019,N_26075);
or U26639 (N_26639,N_26374,N_26227);
xnor U26640 (N_26640,N_26316,N_26267);
nand U26641 (N_26641,N_26050,N_26181);
and U26642 (N_26642,N_26213,N_26305);
and U26643 (N_26643,N_26406,N_26472);
xor U26644 (N_26644,N_26495,N_26310);
nor U26645 (N_26645,N_26328,N_26264);
and U26646 (N_26646,N_26006,N_26139);
and U26647 (N_26647,N_26409,N_26077);
or U26648 (N_26648,N_26195,N_26095);
or U26649 (N_26649,N_26207,N_26262);
and U26650 (N_26650,N_26246,N_26126);
nor U26651 (N_26651,N_26180,N_26476);
or U26652 (N_26652,N_26386,N_26412);
or U26653 (N_26653,N_26106,N_26010);
and U26654 (N_26654,N_26055,N_26484);
nand U26655 (N_26655,N_26134,N_26278);
nor U26656 (N_26656,N_26293,N_26130);
or U26657 (N_26657,N_26235,N_26337);
and U26658 (N_26658,N_26289,N_26317);
or U26659 (N_26659,N_26323,N_26464);
nor U26660 (N_26660,N_26402,N_26238);
xor U26661 (N_26661,N_26120,N_26135);
nand U26662 (N_26662,N_26483,N_26345);
nand U26663 (N_26663,N_26333,N_26091);
nor U26664 (N_26664,N_26329,N_26443);
nand U26665 (N_26665,N_26423,N_26467);
nor U26666 (N_26666,N_26277,N_26269);
and U26667 (N_26667,N_26122,N_26499);
nor U26668 (N_26668,N_26439,N_26115);
nor U26669 (N_26669,N_26186,N_26470);
xor U26670 (N_26670,N_26210,N_26069);
xor U26671 (N_26671,N_26425,N_26388);
nand U26672 (N_26672,N_26114,N_26203);
nor U26673 (N_26673,N_26487,N_26343);
nor U26674 (N_26674,N_26032,N_26438);
and U26675 (N_26675,N_26330,N_26036);
or U26676 (N_26676,N_26000,N_26142);
nand U26677 (N_26677,N_26275,N_26400);
nor U26678 (N_26678,N_26017,N_26204);
and U26679 (N_26679,N_26415,N_26318);
nor U26680 (N_26680,N_26391,N_26411);
xor U26681 (N_26681,N_26218,N_26276);
xor U26682 (N_26682,N_26326,N_26370);
nor U26683 (N_26683,N_26416,N_26179);
nor U26684 (N_26684,N_26247,N_26094);
nor U26685 (N_26685,N_26265,N_26369);
xnor U26686 (N_26686,N_26405,N_26061);
and U26687 (N_26687,N_26481,N_26384);
or U26688 (N_26688,N_26413,N_26466);
nand U26689 (N_26689,N_26441,N_26177);
or U26690 (N_26690,N_26396,N_26046);
or U26691 (N_26691,N_26168,N_26248);
and U26692 (N_26692,N_26459,N_26270);
and U26693 (N_26693,N_26249,N_26480);
nand U26694 (N_26694,N_26081,N_26206);
nand U26695 (N_26695,N_26071,N_26233);
and U26696 (N_26696,N_26051,N_26129);
nand U26697 (N_26697,N_26294,N_26127);
and U26698 (N_26698,N_26256,N_26311);
or U26699 (N_26699,N_26133,N_26348);
and U26700 (N_26700,N_26072,N_26266);
and U26701 (N_26701,N_26295,N_26376);
nand U26702 (N_26702,N_26364,N_26279);
nand U26703 (N_26703,N_26009,N_26286);
nor U26704 (N_26704,N_26123,N_26089);
and U26705 (N_26705,N_26491,N_26136);
and U26706 (N_26706,N_26298,N_26059);
xor U26707 (N_26707,N_26182,N_26365);
or U26708 (N_26708,N_26401,N_26018);
and U26709 (N_26709,N_26381,N_26166);
nand U26710 (N_26710,N_26455,N_26393);
nor U26711 (N_26711,N_26082,N_26260);
nor U26712 (N_26712,N_26228,N_26124);
xnor U26713 (N_26713,N_26450,N_26060);
xnor U26714 (N_26714,N_26358,N_26255);
nor U26715 (N_26715,N_26038,N_26056);
nor U26716 (N_26716,N_26306,N_26490);
nand U26717 (N_26717,N_26473,N_26261);
nand U26718 (N_26718,N_26121,N_26301);
or U26719 (N_26719,N_26153,N_26431);
or U26720 (N_26720,N_26492,N_26212);
nand U26721 (N_26721,N_26475,N_26041);
nor U26722 (N_26722,N_26454,N_26422);
nor U26723 (N_26723,N_26104,N_26250);
nor U26724 (N_26724,N_26241,N_26040);
or U26725 (N_26725,N_26150,N_26027);
nor U26726 (N_26726,N_26189,N_26296);
nand U26727 (N_26727,N_26373,N_26024);
nor U26728 (N_26728,N_26392,N_26184);
nor U26729 (N_26729,N_26202,N_26290);
xor U26730 (N_26730,N_26320,N_26037);
nor U26731 (N_26731,N_26299,N_26132);
xor U26732 (N_26732,N_26161,N_26190);
nand U26733 (N_26733,N_26131,N_26448);
nand U26734 (N_26734,N_26462,N_26347);
or U26735 (N_26735,N_26196,N_26144);
nand U26736 (N_26736,N_26070,N_26109);
and U26737 (N_26737,N_26108,N_26170);
xnor U26738 (N_26738,N_26232,N_26007);
nand U26739 (N_26739,N_26456,N_26447);
nand U26740 (N_26740,N_26096,N_26064);
xnor U26741 (N_26741,N_26314,N_26028);
or U26742 (N_26742,N_26418,N_26242);
nor U26743 (N_26743,N_26098,N_26049);
or U26744 (N_26744,N_26154,N_26149);
or U26745 (N_26745,N_26253,N_26251);
and U26746 (N_26746,N_26107,N_26167);
or U26747 (N_26747,N_26432,N_26357);
nand U26748 (N_26748,N_26084,N_26319);
nor U26749 (N_26749,N_26366,N_26113);
and U26750 (N_26750,N_26008,N_26495);
or U26751 (N_26751,N_26355,N_26172);
xor U26752 (N_26752,N_26495,N_26069);
xor U26753 (N_26753,N_26316,N_26362);
nand U26754 (N_26754,N_26411,N_26230);
and U26755 (N_26755,N_26236,N_26211);
xor U26756 (N_26756,N_26348,N_26090);
or U26757 (N_26757,N_26084,N_26249);
xnor U26758 (N_26758,N_26455,N_26477);
and U26759 (N_26759,N_26421,N_26470);
nand U26760 (N_26760,N_26026,N_26168);
nand U26761 (N_26761,N_26005,N_26151);
nand U26762 (N_26762,N_26337,N_26374);
and U26763 (N_26763,N_26067,N_26333);
nand U26764 (N_26764,N_26235,N_26279);
nor U26765 (N_26765,N_26112,N_26309);
nor U26766 (N_26766,N_26312,N_26450);
or U26767 (N_26767,N_26304,N_26431);
xor U26768 (N_26768,N_26315,N_26328);
nor U26769 (N_26769,N_26250,N_26026);
nand U26770 (N_26770,N_26069,N_26130);
and U26771 (N_26771,N_26008,N_26345);
xnor U26772 (N_26772,N_26054,N_26450);
nor U26773 (N_26773,N_26224,N_26411);
xor U26774 (N_26774,N_26433,N_26047);
nor U26775 (N_26775,N_26484,N_26366);
xnor U26776 (N_26776,N_26062,N_26267);
or U26777 (N_26777,N_26196,N_26250);
nand U26778 (N_26778,N_26262,N_26148);
and U26779 (N_26779,N_26425,N_26385);
or U26780 (N_26780,N_26357,N_26028);
nand U26781 (N_26781,N_26055,N_26307);
nor U26782 (N_26782,N_26448,N_26280);
or U26783 (N_26783,N_26008,N_26228);
xor U26784 (N_26784,N_26302,N_26049);
xor U26785 (N_26785,N_26262,N_26408);
or U26786 (N_26786,N_26088,N_26217);
xnor U26787 (N_26787,N_26217,N_26209);
xor U26788 (N_26788,N_26470,N_26031);
or U26789 (N_26789,N_26426,N_26037);
nor U26790 (N_26790,N_26163,N_26043);
or U26791 (N_26791,N_26421,N_26333);
and U26792 (N_26792,N_26165,N_26118);
or U26793 (N_26793,N_26404,N_26170);
nor U26794 (N_26794,N_26165,N_26292);
or U26795 (N_26795,N_26096,N_26482);
and U26796 (N_26796,N_26310,N_26114);
or U26797 (N_26797,N_26154,N_26066);
xnor U26798 (N_26798,N_26130,N_26459);
or U26799 (N_26799,N_26482,N_26261);
xnor U26800 (N_26800,N_26321,N_26477);
nand U26801 (N_26801,N_26316,N_26357);
nor U26802 (N_26802,N_26118,N_26137);
nor U26803 (N_26803,N_26103,N_26499);
nor U26804 (N_26804,N_26392,N_26268);
nand U26805 (N_26805,N_26033,N_26279);
nor U26806 (N_26806,N_26477,N_26298);
nor U26807 (N_26807,N_26046,N_26345);
nor U26808 (N_26808,N_26015,N_26007);
xor U26809 (N_26809,N_26239,N_26431);
or U26810 (N_26810,N_26443,N_26485);
and U26811 (N_26811,N_26320,N_26286);
xor U26812 (N_26812,N_26429,N_26441);
nand U26813 (N_26813,N_26043,N_26162);
nand U26814 (N_26814,N_26006,N_26027);
nor U26815 (N_26815,N_26233,N_26109);
nor U26816 (N_26816,N_26287,N_26113);
nor U26817 (N_26817,N_26217,N_26228);
nand U26818 (N_26818,N_26215,N_26469);
and U26819 (N_26819,N_26311,N_26061);
nor U26820 (N_26820,N_26311,N_26289);
nand U26821 (N_26821,N_26150,N_26340);
nand U26822 (N_26822,N_26121,N_26365);
nand U26823 (N_26823,N_26346,N_26218);
and U26824 (N_26824,N_26105,N_26174);
and U26825 (N_26825,N_26069,N_26382);
nor U26826 (N_26826,N_26332,N_26041);
nand U26827 (N_26827,N_26279,N_26318);
and U26828 (N_26828,N_26018,N_26354);
or U26829 (N_26829,N_26221,N_26414);
and U26830 (N_26830,N_26023,N_26176);
nor U26831 (N_26831,N_26310,N_26216);
and U26832 (N_26832,N_26288,N_26216);
nor U26833 (N_26833,N_26053,N_26493);
xnor U26834 (N_26834,N_26091,N_26490);
and U26835 (N_26835,N_26479,N_26344);
nor U26836 (N_26836,N_26203,N_26485);
xnor U26837 (N_26837,N_26279,N_26042);
or U26838 (N_26838,N_26043,N_26352);
nor U26839 (N_26839,N_26451,N_26143);
nor U26840 (N_26840,N_26210,N_26346);
or U26841 (N_26841,N_26457,N_26214);
or U26842 (N_26842,N_26069,N_26278);
xor U26843 (N_26843,N_26176,N_26311);
nand U26844 (N_26844,N_26382,N_26354);
and U26845 (N_26845,N_26310,N_26198);
xnor U26846 (N_26846,N_26112,N_26094);
nand U26847 (N_26847,N_26468,N_26499);
and U26848 (N_26848,N_26454,N_26235);
and U26849 (N_26849,N_26005,N_26191);
nand U26850 (N_26850,N_26195,N_26292);
nor U26851 (N_26851,N_26429,N_26126);
nand U26852 (N_26852,N_26089,N_26350);
and U26853 (N_26853,N_26072,N_26383);
xnor U26854 (N_26854,N_26018,N_26086);
or U26855 (N_26855,N_26352,N_26300);
xor U26856 (N_26856,N_26305,N_26490);
nand U26857 (N_26857,N_26287,N_26189);
xnor U26858 (N_26858,N_26203,N_26142);
xnor U26859 (N_26859,N_26389,N_26425);
xnor U26860 (N_26860,N_26024,N_26023);
nand U26861 (N_26861,N_26377,N_26088);
nand U26862 (N_26862,N_26173,N_26417);
and U26863 (N_26863,N_26189,N_26410);
and U26864 (N_26864,N_26389,N_26439);
or U26865 (N_26865,N_26113,N_26311);
nor U26866 (N_26866,N_26395,N_26495);
and U26867 (N_26867,N_26446,N_26467);
nand U26868 (N_26868,N_26040,N_26037);
xor U26869 (N_26869,N_26447,N_26040);
xnor U26870 (N_26870,N_26340,N_26118);
nor U26871 (N_26871,N_26384,N_26428);
xor U26872 (N_26872,N_26137,N_26155);
nor U26873 (N_26873,N_26236,N_26066);
nand U26874 (N_26874,N_26454,N_26249);
xor U26875 (N_26875,N_26297,N_26388);
and U26876 (N_26876,N_26288,N_26241);
nand U26877 (N_26877,N_26299,N_26201);
nor U26878 (N_26878,N_26120,N_26407);
xor U26879 (N_26879,N_26285,N_26157);
nand U26880 (N_26880,N_26460,N_26351);
and U26881 (N_26881,N_26149,N_26315);
and U26882 (N_26882,N_26371,N_26141);
xor U26883 (N_26883,N_26262,N_26307);
nand U26884 (N_26884,N_26442,N_26448);
nand U26885 (N_26885,N_26258,N_26148);
xnor U26886 (N_26886,N_26435,N_26307);
nor U26887 (N_26887,N_26236,N_26291);
xor U26888 (N_26888,N_26385,N_26110);
xor U26889 (N_26889,N_26258,N_26119);
or U26890 (N_26890,N_26253,N_26067);
and U26891 (N_26891,N_26402,N_26013);
nor U26892 (N_26892,N_26383,N_26275);
and U26893 (N_26893,N_26036,N_26426);
or U26894 (N_26894,N_26188,N_26127);
nand U26895 (N_26895,N_26151,N_26061);
or U26896 (N_26896,N_26308,N_26252);
nand U26897 (N_26897,N_26002,N_26084);
nor U26898 (N_26898,N_26263,N_26483);
nand U26899 (N_26899,N_26027,N_26437);
and U26900 (N_26900,N_26307,N_26401);
nand U26901 (N_26901,N_26259,N_26429);
xor U26902 (N_26902,N_26025,N_26072);
or U26903 (N_26903,N_26140,N_26488);
and U26904 (N_26904,N_26470,N_26370);
or U26905 (N_26905,N_26002,N_26206);
nor U26906 (N_26906,N_26312,N_26099);
and U26907 (N_26907,N_26097,N_26066);
nand U26908 (N_26908,N_26344,N_26270);
nand U26909 (N_26909,N_26175,N_26074);
nor U26910 (N_26910,N_26321,N_26207);
nor U26911 (N_26911,N_26375,N_26245);
nor U26912 (N_26912,N_26312,N_26282);
nor U26913 (N_26913,N_26094,N_26121);
nor U26914 (N_26914,N_26025,N_26107);
nand U26915 (N_26915,N_26482,N_26329);
nand U26916 (N_26916,N_26153,N_26146);
nand U26917 (N_26917,N_26046,N_26273);
nor U26918 (N_26918,N_26079,N_26068);
and U26919 (N_26919,N_26333,N_26158);
xor U26920 (N_26920,N_26282,N_26111);
nand U26921 (N_26921,N_26030,N_26193);
or U26922 (N_26922,N_26190,N_26153);
nand U26923 (N_26923,N_26452,N_26369);
xnor U26924 (N_26924,N_26036,N_26457);
and U26925 (N_26925,N_26126,N_26079);
or U26926 (N_26926,N_26048,N_26476);
xnor U26927 (N_26927,N_26273,N_26240);
nor U26928 (N_26928,N_26278,N_26262);
nor U26929 (N_26929,N_26223,N_26330);
and U26930 (N_26930,N_26243,N_26438);
or U26931 (N_26931,N_26291,N_26005);
nand U26932 (N_26932,N_26483,N_26324);
xnor U26933 (N_26933,N_26098,N_26366);
or U26934 (N_26934,N_26162,N_26121);
xor U26935 (N_26935,N_26295,N_26417);
xnor U26936 (N_26936,N_26149,N_26119);
and U26937 (N_26937,N_26135,N_26459);
or U26938 (N_26938,N_26367,N_26148);
and U26939 (N_26939,N_26281,N_26414);
nand U26940 (N_26940,N_26070,N_26195);
xnor U26941 (N_26941,N_26020,N_26424);
nand U26942 (N_26942,N_26276,N_26459);
xnor U26943 (N_26943,N_26060,N_26219);
nor U26944 (N_26944,N_26117,N_26438);
nor U26945 (N_26945,N_26302,N_26424);
and U26946 (N_26946,N_26483,N_26204);
nand U26947 (N_26947,N_26008,N_26287);
or U26948 (N_26948,N_26132,N_26263);
nor U26949 (N_26949,N_26173,N_26313);
nor U26950 (N_26950,N_26252,N_26040);
xnor U26951 (N_26951,N_26229,N_26345);
and U26952 (N_26952,N_26375,N_26421);
and U26953 (N_26953,N_26379,N_26245);
or U26954 (N_26954,N_26296,N_26052);
or U26955 (N_26955,N_26469,N_26447);
xor U26956 (N_26956,N_26145,N_26487);
xnor U26957 (N_26957,N_26280,N_26389);
or U26958 (N_26958,N_26296,N_26030);
xor U26959 (N_26959,N_26120,N_26345);
or U26960 (N_26960,N_26331,N_26038);
nor U26961 (N_26961,N_26413,N_26013);
xnor U26962 (N_26962,N_26149,N_26114);
xnor U26963 (N_26963,N_26437,N_26477);
nor U26964 (N_26964,N_26143,N_26285);
xor U26965 (N_26965,N_26146,N_26184);
nor U26966 (N_26966,N_26344,N_26333);
nor U26967 (N_26967,N_26107,N_26226);
and U26968 (N_26968,N_26227,N_26440);
or U26969 (N_26969,N_26319,N_26169);
and U26970 (N_26970,N_26102,N_26255);
and U26971 (N_26971,N_26389,N_26179);
nor U26972 (N_26972,N_26214,N_26454);
nand U26973 (N_26973,N_26216,N_26385);
nand U26974 (N_26974,N_26441,N_26100);
and U26975 (N_26975,N_26060,N_26132);
or U26976 (N_26976,N_26252,N_26357);
xnor U26977 (N_26977,N_26021,N_26297);
or U26978 (N_26978,N_26127,N_26123);
xor U26979 (N_26979,N_26479,N_26405);
nand U26980 (N_26980,N_26400,N_26294);
and U26981 (N_26981,N_26124,N_26266);
xor U26982 (N_26982,N_26044,N_26240);
nor U26983 (N_26983,N_26232,N_26083);
nor U26984 (N_26984,N_26239,N_26006);
nor U26985 (N_26985,N_26077,N_26417);
nor U26986 (N_26986,N_26393,N_26290);
and U26987 (N_26987,N_26145,N_26206);
or U26988 (N_26988,N_26343,N_26449);
and U26989 (N_26989,N_26340,N_26367);
nand U26990 (N_26990,N_26235,N_26180);
and U26991 (N_26991,N_26003,N_26188);
nor U26992 (N_26992,N_26427,N_26341);
xor U26993 (N_26993,N_26196,N_26413);
nor U26994 (N_26994,N_26013,N_26164);
nor U26995 (N_26995,N_26478,N_26150);
xnor U26996 (N_26996,N_26364,N_26362);
or U26997 (N_26997,N_26171,N_26121);
nand U26998 (N_26998,N_26031,N_26175);
and U26999 (N_26999,N_26014,N_26337);
and U27000 (N_27000,N_26915,N_26692);
nand U27001 (N_27001,N_26840,N_26554);
xor U27002 (N_27002,N_26894,N_26734);
nor U27003 (N_27003,N_26803,N_26611);
or U27004 (N_27004,N_26861,N_26826);
nand U27005 (N_27005,N_26910,N_26656);
nor U27006 (N_27006,N_26684,N_26811);
nor U27007 (N_27007,N_26975,N_26944);
and U27008 (N_27008,N_26675,N_26661);
nor U27009 (N_27009,N_26635,N_26839);
or U27010 (N_27010,N_26682,N_26818);
nand U27011 (N_27011,N_26738,N_26504);
xnor U27012 (N_27012,N_26770,N_26645);
or U27013 (N_27013,N_26882,N_26970);
or U27014 (N_27014,N_26771,N_26750);
or U27015 (N_27015,N_26763,N_26805);
nand U27016 (N_27016,N_26919,N_26776);
nand U27017 (N_27017,N_26769,N_26680);
nand U27018 (N_27018,N_26613,N_26922);
nand U27019 (N_27019,N_26817,N_26722);
or U27020 (N_27020,N_26916,N_26694);
xor U27021 (N_27021,N_26742,N_26555);
and U27022 (N_27022,N_26866,N_26996);
and U27023 (N_27023,N_26860,N_26604);
or U27024 (N_27024,N_26843,N_26991);
nand U27025 (N_27025,N_26886,N_26641);
nor U27026 (N_27026,N_26788,N_26774);
and U27027 (N_27027,N_26848,N_26507);
or U27028 (N_27028,N_26810,N_26527);
nand U27029 (N_27029,N_26535,N_26697);
or U27030 (N_27030,N_26683,N_26831);
nor U27031 (N_27031,N_26510,N_26726);
nand U27032 (N_27032,N_26727,N_26948);
xor U27033 (N_27033,N_26565,N_26812);
nand U27034 (N_27034,N_26949,N_26735);
xnor U27035 (N_27035,N_26652,N_26700);
and U27036 (N_27036,N_26506,N_26560);
and U27037 (N_27037,N_26723,N_26587);
nand U27038 (N_27038,N_26707,N_26868);
and U27039 (N_27039,N_26626,N_26962);
and U27040 (N_27040,N_26930,N_26779);
and U27041 (N_27041,N_26573,N_26899);
or U27042 (N_27042,N_26795,N_26855);
nor U27043 (N_27043,N_26595,N_26824);
and U27044 (N_27044,N_26950,N_26801);
xnor U27045 (N_27045,N_26925,N_26834);
nand U27046 (N_27046,N_26534,N_26719);
nor U27047 (N_27047,N_26516,N_26537);
and U27048 (N_27048,N_26714,N_26556);
and U27049 (N_27049,N_26711,N_26822);
or U27050 (N_27050,N_26836,N_26768);
and U27051 (N_27051,N_26663,N_26724);
nand U27052 (N_27052,N_26521,N_26924);
and U27053 (N_27053,N_26920,N_26881);
nor U27054 (N_27054,N_26851,N_26522);
nor U27055 (N_27055,N_26985,N_26783);
nor U27056 (N_27056,N_26935,N_26689);
or U27057 (N_27057,N_26998,N_26567);
nor U27058 (N_27058,N_26859,N_26501);
nor U27059 (N_27059,N_26829,N_26815);
or U27060 (N_27060,N_26885,N_26702);
and U27061 (N_27061,N_26664,N_26946);
and U27062 (N_27062,N_26736,N_26917);
or U27063 (N_27063,N_26942,N_26729);
nor U27064 (N_27064,N_26901,N_26845);
nand U27065 (N_27065,N_26814,N_26519);
or U27066 (N_27066,N_26819,N_26629);
or U27067 (N_27067,N_26508,N_26888);
and U27068 (N_27068,N_26832,N_26746);
xor U27069 (N_27069,N_26536,N_26932);
xor U27070 (N_27070,N_26551,N_26992);
nand U27071 (N_27071,N_26947,N_26878);
and U27072 (N_27072,N_26863,N_26909);
or U27073 (N_27073,N_26716,N_26647);
nand U27074 (N_27074,N_26913,N_26867);
nor U27075 (N_27075,N_26853,N_26908);
nand U27076 (N_27076,N_26575,N_26717);
nor U27077 (N_27077,N_26701,N_26679);
xor U27078 (N_27078,N_26571,N_26978);
or U27079 (N_27079,N_26790,N_26895);
or U27080 (N_27080,N_26879,N_26982);
xor U27081 (N_27081,N_26877,N_26509);
and U27082 (N_27082,N_26657,N_26753);
nor U27083 (N_27083,N_26951,N_26570);
xnor U27084 (N_27084,N_26512,N_26744);
nor U27085 (N_27085,N_26566,N_26606);
and U27086 (N_27086,N_26673,N_26983);
nand U27087 (N_27087,N_26614,N_26968);
or U27088 (N_27088,N_26852,N_26938);
nand U27089 (N_27089,N_26756,N_26806);
or U27090 (N_27090,N_26989,N_26796);
and U27091 (N_27091,N_26941,N_26772);
nor U27092 (N_27092,N_26609,N_26634);
and U27093 (N_27093,N_26691,N_26802);
nand U27094 (N_27094,N_26576,N_26775);
or U27095 (N_27095,N_26743,N_26637);
xnor U27096 (N_27096,N_26965,N_26631);
and U27097 (N_27097,N_26588,N_26876);
nand U27098 (N_27098,N_26705,N_26710);
nand U27099 (N_27099,N_26653,N_26869);
xnor U27100 (N_27100,N_26599,N_26612);
or U27101 (N_27101,N_26800,N_26593);
xnor U27102 (N_27102,N_26500,N_26754);
and U27103 (N_27103,N_26709,N_26695);
xor U27104 (N_27104,N_26532,N_26524);
and U27105 (N_27105,N_26986,N_26686);
and U27106 (N_27106,N_26579,N_26854);
nand U27107 (N_27107,N_26541,N_26973);
and U27108 (N_27108,N_26563,N_26830);
xnor U27109 (N_27109,N_26961,N_26513);
xor U27110 (N_27110,N_26720,N_26693);
xnor U27111 (N_27111,N_26933,N_26900);
nand U27112 (N_27112,N_26607,N_26601);
nor U27113 (N_27113,N_26622,N_26994);
xor U27114 (N_27114,N_26590,N_26557);
nor U27115 (N_27115,N_26548,N_26773);
and U27116 (N_27116,N_26542,N_26733);
and U27117 (N_27117,N_26666,N_26715);
nand U27118 (N_27118,N_26584,N_26993);
nand U27119 (N_27119,N_26999,N_26858);
and U27120 (N_27120,N_26823,N_26862);
and U27121 (N_27121,N_26791,N_26766);
nand U27122 (N_27122,N_26597,N_26728);
and U27123 (N_27123,N_26636,N_26990);
xnor U27124 (N_27124,N_26929,N_26530);
nand U27125 (N_27125,N_26887,N_26981);
xor U27126 (N_27126,N_26940,N_26850);
and U27127 (N_27127,N_26598,N_26934);
nor U27128 (N_27128,N_26794,N_26623);
xnor U27129 (N_27129,N_26897,N_26725);
or U27130 (N_27130,N_26875,N_26889);
and U27131 (N_27131,N_26677,N_26520);
nand U27132 (N_27132,N_26957,N_26552);
nor U27133 (N_27133,N_26540,N_26649);
nand U27134 (N_27134,N_26706,N_26748);
nand U27135 (N_27135,N_26837,N_26787);
or U27136 (N_27136,N_26997,N_26904);
and U27137 (N_27137,N_26966,N_26643);
nor U27138 (N_27138,N_26568,N_26730);
nand U27139 (N_27139,N_26971,N_26749);
xor U27140 (N_27140,N_26574,N_26610);
xnor U27141 (N_27141,N_26871,N_26865);
or U27142 (N_27142,N_26667,N_26760);
and U27143 (N_27143,N_26639,N_26918);
xnor U27144 (N_27144,N_26669,N_26620);
or U27145 (N_27145,N_26721,N_26870);
nor U27146 (N_27146,N_26959,N_26808);
xor U27147 (N_27147,N_26745,N_26905);
xor U27148 (N_27148,N_26928,N_26621);
or U27149 (N_27149,N_26618,N_26515);
nand U27150 (N_27150,N_26988,N_26931);
nor U27151 (N_27151,N_26615,N_26778);
nand U27152 (N_27152,N_26827,N_26529);
nand U27153 (N_27153,N_26681,N_26712);
xnor U27154 (N_27154,N_26646,N_26577);
nor U27155 (N_27155,N_26907,N_26873);
or U27156 (N_27156,N_26741,N_26650);
or U27157 (N_27157,N_26828,N_26703);
nand U27158 (N_27158,N_26671,N_26891);
nand U27159 (N_27159,N_26525,N_26580);
nor U27160 (N_27160,N_26651,N_26658);
and U27161 (N_27161,N_26953,N_26898);
nor U27162 (N_27162,N_26864,N_26648);
nand U27163 (N_27163,N_26505,N_26846);
or U27164 (N_27164,N_26572,N_26539);
xnor U27165 (N_27165,N_26708,N_26668);
xor U27166 (N_27166,N_26739,N_26676);
xor U27167 (N_27167,N_26856,N_26502);
nand U27168 (N_27168,N_26591,N_26893);
and U27169 (N_27169,N_26936,N_26632);
nor U27170 (N_27170,N_26628,N_26546);
xor U27171 (N_27171,N_26586,N_26782);
and U27172 (N_27172,N_26562,N_26758);
xnor U27173 (N_27173,N_26807,N_26678);
and U27174 (N_27174,N_26777,N_26955);
nor U27175 (N_27175,N_26841,N_26977);
or U27176 (N_27176,N_26964,N_26762);
nand U27177 (N_27177,N_26799,N_26761);
or U27178 (N_27178,N_26600,N_26872);
nor U27179 (N_27179,N_26644,N_26594);
or U27180 (N_27180,N_26857,N_26533);
and U27181 (N_27181,N_26627,N_26528);
or U27182 (N_27182,N_26624,N_26937);
xnor U27183 (N_27183,N_26902,N_26883);
xnor U27184 (N_27184,N_26583,N_26972);
nand U27185 (N_27185,N_26747,N_26820);
or U27186 (N_27186,N_26903,N_26764);
xor U27187 (N_27187,N_26561,N_26596);
or U27188 (N_27188,N_26699,N_26847);
nor U27189 (N_27189,N_26984,N_26798);
nor U27190 (N_27190,N_26813,N_26558);
and U27191 (N_27191,N_26617,N_26765);
or U27192 (N_27192,N_26665,N_26543);
or U27193 (N_27193,N_26655,N_26969);
or U27194 (N_27194,N_26732,N_26514);
xnor U27195 (N_27195,N_26792,N_26740);
xnor U27196 (N_27196,N_26526,N_26670);
xnor U27197 (N_27197,N_26659,N_26550);
xnor U27198 (N_27198,N_26995,N_26939);
nor U27199 (N_27199,N_26927,N_26906);
and U27200 (N_27200,N_26954,N_26833);
nand U27201 (N_27201,N_26688,N_26974);
or U27202 (N_27202,N_26980,N_26912);
nor U27203 (N_27203,N_26585,N_26967);
or U27204 (N_27204,N_26757,N_26958);
nand U27205 (N_27205,N_26625,N_26633);
or U27206 (N_27206,N_26896,N_26654);
and U27207 (N_27207,N_26698,N_26821);
or U27208 (N_27208,N_26638,N_26780);
and U27209 (N_27209,N_26553,N_26838);
or U27210 (N_27210,N_26549,N_26696);
xnor U27211 (N_27211,N_26713,N_26603);
nand U27212 (N_27212,N_26564,N_26503);
nor U27213 (N_27213,N_26874,N_26582);
or U27214 (N_27214,N_26602,N_26825);
or U27215 (N_27215,N_26616,N_26718);
xor U27216 (N_27216,N_26685,N_26605);
nor U27217 (N_27217,N_26786,N_26842);
and U27218 (N_27218,N_26731,N_26578);
nor U27219 (N_27219,N_26979,N_26785);
nand U27220 (N_27220,N_26662,N_26956);
xnor U27221 (N_27221,N_26789,N_26672);
nand U27222 (N_27222,N_26687,N_26926);
nor U27223 (N_27223,N_26531,N_26849);
and U27224 (N_27224,N_26884,N_26914);
xor U27225 (N_27225,N_26890,N_26518);
nor U27226 (N_27226,N_26911,N_26804);
and U27227 (N_27227,N_26538,N_26784);
nor U27228 (N_27228,N_26674,N_26511);
or U27229 (N_27229,N_26547,N_26960);
or U27230 (N_27230,N_26963,N_26809);
xnor U27231 (N_27231,N_26755,N_26545);
xnor U27232 (N_27232,N_26737,N_26976);
nand U27233 (N_27233,N_26816,N_26759);
and U27234 (N_27234,N_26952,N_26751);
or U27235 (N_27235,N_26523,N_26752);
xnor U27236 (N_27236,N_26844,N_26945);
xnor U27237 (N_27237,N_26517,N_26544);
and U27238 (N_27238,N_26569,N_26704);
nor U27239 (N_27239,N_26921,N_26767);
xnor U27240 (N_27240,N_26892,N_26619);
xnor U27241 (N_27241,N_26835,N_26660);
nor U27242 (N_27242,N_26793,N_26630);
and U27243 (N_27243,N_26781,N_26987);
xnor U27244 (N_27244,N_26559,N_26592);
or U27245 (N_27245,N_26640,N_26608);
nand U27246 (N_27246,N_26589,N_26797);
and U27247 (N_27247,N_26581,N_26943);
nand U27248 (N_27248,N_26642,N_26923);
and U27249 (N_27249,N_26690,N_26880);
xnor U27250 (N_27250,N_26915,N_26922);
nor U27251 (N_27251,N_26735,N_26521);
nand U27252 (N_27252,N_26670,N_26975);
xnor U27253 (N_27253,N_26556,N_26784);
and U27254 (N_27254,N_26795,N_26758);
nor U27255 (N_27255,N_26934,N_26752);
nor U27256 (N_27256,N_26990,N_26996);
nand U27257 (N_27257,N_26508,N_26670);
nand U27258 (N_27258,N_26614,N_26572);
or U27259 (N_27259,N_26986,N_26762);
nand U27260 (N_27260,N_26839,N_26847);
and U27261 (N_27261,N_26676,N_26893);
nand U27262 (N_27262,N_26719,N_26804);
xnor U27263 (N_27263,N_26861,N_26814);
nor U27264 (N_27264,N_26530,N_26996);
nor U27265 (N_27265,N_26884,N_26571);
and U27266 (N_27266,N_26811,N_26748);
or U27267 (N_27267,N_26693,N_26675);
xor U27268 (N_27268,N_26974,N_26754);
xor U27269 (N_27269,N_26794,N_26514);
nor U27270 (N_27270,N_26673,N_26580);
xnor U27271 (N_27271,N_26983,N_26705);
xnor U27272 (N_27272,N_26784,N_26798);
and U27273 (N_27273,N_26531,N_26921);
nand U27274 (N_27274,N_26619,N_26551);
xnor U27275 (N_27275,N_26611,N_26990);
or U27276 (N_27276,N_26556,N_26653);
nand U27277 (N_27277,N_26693,N_26721);
or U27278 (N_27278,N_26991,N_26778);
nand U27279 (N_27279,N_26962,N_26578);
or U27280 (N_27280,N_26910,N_26530);
and U27281 (N_27281,N_26865,N_26587);
nand U27282 (N_27282,N_26766,N_26747);
xnor U27283 (N_27283,N_26642,N_26900);
nand U27284 (N_27284,N_26520,N_26988);
or U27285 (N_27285,N_26606,N_26696);
and U27286 (N_27286,N_26849,N_26655);
or U27287 (N_27287,N_26758,N_26760);
xor U27288 (N_27288,N_26852,N_26547);
nor U27289 (N_27289,N_26883,N_26518);
and U27290 (N_27290,N_26664,N_26558);
nand U27291 (N_27291,N_26812,N_26967);
xor U27292 (N_27292,N_26803,N_26911);
xor U27293 (N_27293,N_26916,N_26653);
xnor U27294 (N_27294,N_26674,N_26500);
and U27295 (N_27295,N_26778,N_26883);
or U27296 (N_27296,N_26914,N_26931);
xor U27297 (N_27297,N_26721,N_26831);
or U27298 (N_27298,N_26544,N_26922);
xnor U27299 (N_27299,N_26775,N_26957);
or U27300 (N_27300,N_26760,N_26599);
and U27301 (N_27301,N_26814,N_26514);
nand U27302 (N_27302,N_26907,N_26609);
nand U27303 (N_27303,N_26513,N_26900);
or U27304 (N_27304,N_26938,N_26873);
xnor U27305 (N_27305,N_26502,N_26661);
nand U27306 (N_27306,N_26540,N_26788);
and U27307 (N_27307,N_26897,N_26875);
or U27308 (N_27308,N_26729,N_26673);
and U27309 (N_27309,N_26655,N_26536);
nand U27310 (N_27310,N_26737,N_26752);
nand U27311 (N_27311,N_26744,N_26906);
or U27312 (N_27312,N_26509,N_26687);
or U27313 (N_27313,N_26858,N_26784);
and U27314 (N_27314,N_26625,N_26713);
and U27315 (N_27315,N_26812,N_26995);
and U27316 (N_27316,N_26676,N_26714);
nand U27317 (N_27317,N_26508,N_26998);
or U27318 (N_27318,N_26941,N_26854);
nor U27319 (N_27319,N_26634,N_26642);
nand U27320 (N_27320,N_26564,N_26570);
and U27321 (N_27321,N_26726,N_26640);
and U27322 (N_27322,N_26615,N_26702);
nand U27323 (N_27323,N_26954,N_26532);
nor U27324 (N_27324,N_26543,N_26652);
nor U27325 (N_27325,N_26518,N_26766);
nor U27326 (N_27326,N_26955,N_26670);
nor U27327 (N_27327,N_26776,N_26691);
or U27328 (N_27328,N_26706,N_26965);
nand U27329 (N_27329,N_26557,N_26604);
nand U27330 (N_27330,N_26650,N_26782);
nand U27331 (N_27331,N_26634,N_26775);
nand U27332 (N_27332,N_26704,N_26636);
nor U27333 (N_27333,N_26511,N_26768);
or U27334 (N_27334,N_26904,N_26846);
and U27335 (N_27335,N_26796,N_26859);
nor U27336 (N_27336,N_26690,N_26771);
nor U27337 (N_27337,N_26802,N_26963);
nand U27338 (N_27338,N_26850,N_26778);
nor U27339 (N_27339,N_26596,N_26766);
and U27340 (N_27340,N_26754,N_26521);
nor U27341 (N_27341,N_26782,N_26996);
nor U27342 (N_27342,N_26883,N_26792);
nand U27343 (N_27343,N_26933,N_26567);
and U27344 (N_27344,N_26970,N_26872);
and U27345 (N_27345,N_26646,N_26890);
and U27346 (N_27346,N_26984,N_26928);
xnor U27347 (N_27347,N_26820,N_26614);
xor U27348 (N_27348,N_26824,N_26944);
xor U27349 (N_27349,N_26610,N_26937);
xnor U27350 (N_27350,N_26810,N_26979);
nor U27351 (N_27351,N_26747,N_26647);
xor U27352 (N_27352,N_26907,N_26567);
xor U27353 (N_27353,N_26785,N_26666);
or U27354 (N_27354,N_26740,N_26863);
xnor U27355 (N_27355,N_26731,N_26726);
nor U27356 (N_27356,N_26715,N_26537);
and U27357 (N_27357,N_26516,N_26929);
nand U27358 (N_27358,N_26755,N_26939);
nor U27359 (N_27359,N_26685,N_26580);
nand U27360 (N_27360,N_26577,N_26866);
nand U27361 (N_27361,N_26776,N_26654);
and U27362 (N_27362,N_26861,N_26666);
and U27363 (N_27363,N_26771,N_26683);
or U27364 (N_27364,N_26824,N_26841);
nand U27365 (N_27365,N_26853,N_26810);
and U27366 (N_27366,N_26596,N_26682);
or U27367 (N_27367,N_26746,N_26892);
and U27368 (N_27368,N_26519,N_26514);
xor U27369 (N_27369,N_26843,N_26887);
and U27370 (N_27370,N_26814,N_26987);
nand U27371 (N_27371,N_26663,N_26766);
or U27372 (N_27372,N_26723,N_26903);
xnor U27373 (N_27373,N_26810,N_26777);
and U27374 (N_27374,N_26865,N_26529);
nor U27375 (N_27375,N_26915,N_26955);
nand U27376 (N_27376,N_26823,N_26967);
or U27377 (N_27377,N_26701,N_26967);
and U27378 (N_27378,N_26972,N_26880);
nand U27379 (N_27379,N_26602,N_26517);
xnor U27380 (N_27380,N_26552,N_26682);
xor U27381 (N_27381,N_26694,N_26665);
xnor U27382 (N_27382,N_26796,N_26506);
and U27383 (N_27383,N_26869,N_26564);
and U27384 (N_27384,N_26928,N_26875);
and U27385 (N_27385,N_26701,N_26703);
and U27386 (N_27386,N_26566,N_26692);
xnor U27387 (N_27387,N_26581,N_26734);
nand U27388 (N_27388,N_26922,N_26876);
nand U27389 (N_27389,N_26656,N_26662);
or U27390 (N_27390,N_26807,N_26786);
or U27391 (N_27391,N_26976,N_26700);
xor U27392 (N_27392,N_26775,N_26503);
nand U27393 (N_27393,N_26524,N_26968);
nand U27394 (N_27394,N_26980,N_26826);
and U27395 (N_27395,N_26926,N_26613);
and U27396 (N_27396,N_26659,N_26630);
nor U27397 (N_27397,N_26929,N_26603);
nor U27398 (N_27398,N_26861,N_26513);
xor U27399 (N_27399,N_26522,N_26623);
or U27400 (N_27400,N_26672,N_26510);
nand U27401 (N_27401,N_26781,N_26651);
nor U27402 (N_27402,N_26804,N_26596);
nand U27403 (N_27403,N_26842,N_26568);
nand U27404 (N_27404,N_26906,N_26874);
or U27405 (N_27405,N_26903,N_26626);
or U27406 (N_27406,N_26547,N_26784);
nand U27407 (N_27407,N_26551,N_26589);
nor U27408 (N_27408,N_26913,N_26763);
and U27409 (N_27409,N_26724,N_26965);
nor U27410 (N_27410,N_26711,N_26839);
or U27411 (N_27411,N_26866,N_26814);
and U27412 (N_27412,N_26711,N_26557);
nor U27413 (N_27413,N_26539,N_26845);
xor U27414 (N_27414,N_26623,N_26669);
or U27415 (N_27415,N_26844,N_26707);
xnor U27416 (N_27416,N_26919,N_26872);
and U27417 (N_27417,N_26762,N_26949);
and U27418 (N_27418,N_26831,N_26918);
nand U27419 (N_27419,N_26633,N_26650);
xor U27420 (N_27420,N_26662,N_26528);
or U27421 (N_27421,N_26681,N_26994);
nor U27422 (N_27422,N_26871,N_26813);
or U27423 (N_27423,N_26929,N_26767);
and U27424 (N_27424,N_26806,N_26821);
xnor U27425 (N_27425,N_26872,N_26773);
and U27426 (N_27426,N_26802,N_26690);
or U27427 (N_27427,N_26803,N_26636);
and U27428 (N_27428,N_26959,N_26781);
xor U27429 (N_27429,N_26894,N_26711);
and U27430 (N_27430,N_26599,N_26856);
or U27431 (N_27431,N_26566,N_26670);
or U27432 (N_27432,N_26853,N_26675);
nand U27433 (N_27433,N_26523,N_26896);
xnor U27434 (N_27434,N_26545,N_26567);
nor U27435 (N_27435,N_26611,N_26927);
nor U27436 (N_27436,N_26979,N_26579);
nand U27437 (N_27437,N_26849,N_26854);
nor U27438 (N_27438,N_26588,N_26693);
or U27439 (N_27439,N_26856,N_26764);
or U27440 (N_27440,N_26551,N_26794);
xnor U27441 (N_27441,N_26593,N_26814);
nor U27442 (N_27442,N_26803,N_26591);
nand U27443 (N_27443,N_26985,N_26953);
nand U27444 (N_27444,N_26630,N_26818);
xnor U27445 (N_27445,N_26992,N_26804);
or U27446 (N_27446,N_26543,N_26894);
nand U27447 (N_27447,N_26721,N_26759);
nor U27448 (N_27448,N_26731,N_26602);
xor U27449 (N_27449,N_26647,N_26518);
xor U27450 (N_27450,N_26769,N_26598);
or U27451 (N_27451,N_26571,N_26863);
nor U27452 (N_27452,N_26635,N_26519);
nand U27453 (N_27453,N_26967,N_26626);
and U27454 (N_27454,N_26992,N_26622);
xnor U27455 (N_27455,N_26757,N_26682);
nand U27456 (N_27456,N_26752,N_26502);
xor U27457 (N_27457,N_26722,N_26585);
xor U27458 (N_27458,N_26745,N_26731);
nand U27459 (N_27459,N_26618,N_26907);
xnor U27460 (N_27460,N_26840,N_26555);
or U27461 (N_27461,N_26708,N_26709);
xor U27462 (N_27462,N_26697,N_26813);
nand U27463 (N_27463,N_26851,N_26707);
or U27464 (N_27464,N_26843,N_26574);
nand U27465 (N_27465,N_26572,N_26663);
xnor U27466 (N_27466,N_26792,N_26503);
nor U27467 (N_27467,N_26609,N_26633);
or U27468 (N_27468,N_26765,N_26579);
nor U27469 (N_27469,N_26757,N_26939);
and U27470 (N_27470,N_26749,N_26727);
and U27471 (N_27471,N_26548,N_26986);
and U27472 (N_27472,N_26944,N_26986);
or U27473 (N_27473,N_26623,N_26547);
and U27474 (N_27474,N_26802,N_26950);
nand U27475 (N_27475,N_26713,N_26710);
xnor U27476 (N_27476,N_26602,N_26767);
xor U27477 (N_27477,N_26734,N_26504);
xor U27478 (N_27478,N_26503,N_26689);
or U27479 (N_27479,N_26607,N_26741);
nor U27480 (N_27480,N_26651,N_26511);
or U27481 (N_27481,N_26660,N_26971);
nor U27482 (N_27482,N_26545,N_26611);
nand U27483 (N_27483,N_26957,N_26955);
and U27484 (N_27484,N_26546,N_26993);
or U27485 (N_27485,N_26689,N_26505);
nand U27486 (N_27486,N_26860,N_26544);
or U27487 (N_27487,N_26933,N_26606);
nand U27488 (N_27488,N_26573,N_26617);
and U27489 (N_27489,N_26713,N_26582);
nor U27490 (N_27490,N_26891,N_26887);
nor U27491 (N_27491,N_26616,N_26897);
nand U27492 (N_27492,N_26772,N_26657);
nand U27493 (N_27493,N_26622,N_26743);
and U27494 (N_27494,N_26580,N_26555);
nor U27495 (N_27495,N_26596,N_26563);
nand U27496 (N_27496,N_26809,N_26659);
nor U27497 (N_27497,N_26785,N_26724);
xnor U27498 (N_27498,N_26951,N_26760);
and U27499 (N_27499,N_26930,N_26973);
nand U27500 (N_27500,N_27343,N_27059);
nand U27501 (N_27501,N_27421,N_27222);
nand U27502 (N_27502,N_27102,N_27287);
nand U27503 (N_27503,N_27351,N_27472);
nor U27504 (N_27504,N_27228,N_27128);
xnor U27505 (N_27505,N_27290,N_27466);
xnor U27506 (N_27506,N_27104,N_27329);
or U27507 (N_27507,N_27109,N_27432);
and U27508 (N_27508,N_27181,N_27043);
xor U27509 (N_27509,N_27154,N_27010);
nand U27510 (N_27510,N_27251,N_27435);
nand U27511 (N_27511,N_27157,N_27315);
xor U27512 (N_27512,N_27121,N_27212);
xor U27513 (N_27513,N_27323,N_27230);
xor U27514 (N_27514,N_27373,N_27134);
xor U27515 (N_27515,N_27221,N_27397);
xnor U27516 (N_27516,N_27112,N_27022);
xnor U27517 (N_27517,N_27079,N_27327);
nor U27518 (N_27518,N_27250,N_27015);
nand U27519 (N_27519,N_27027,N_27114);
nand U27520 (N_27520,N_27280,N_27414);
or U27521 (N_27521,N_27139,N_27352);
or U27522 (N_27522,N_27493,N_27158);
nor U27523 (N_27523,N_27156,N_27370);
nand U27524 (N_27524,N_27462,N_27091);
xnor U27525 (N_27525,N_27021,N_27293);
nor U27526 (N_27526,N_27269,N_27305);
nor U27527 (N_27527,N_27444,N_27053);
or U27528 (N_27528,N_27190,N_27144);
or U27529 (N_27529,N_27403,N_27299);
and U27530 (N_27530,N_27488,N_27490);
nor U27531 (N_27531,N_27301,N_27012);
nand U27532 (N_27532,N_27252,N_27098);
and U27533 (N_27533,N_27185,N_27311);
xnor U27534 (N_27534,N_27032,N_27468);
nand U27535 (N_27535,N_27498,N_27197);
or U27536 (N_27536,N_27070,N_27087);
nor U27537 (N_27537,N_27470,N_27415);
xor U27538 (N_27538,N_27491,N_27233);
nand U27539 (N_27539,N_27424,N_27030);
xor U27540 (N_27540,N_27391,N_27120);
or U27541 (N_27541,N_27036,N_27009);
or U27542 (N_27542,N_27389,N_27013);
xnor U27543 (N_27543,N_27113,N_27001);
nand U27544 (N_27544,N_27225,N_27253);
nor U27545 (N_27545,N_27271,N_27122);
nand U27546 (N_27546,N_27038,N_27055);
or U27547 (N_27547,N_27460,N_27308);
or U27548 (N_27548,N_27071,N_27454);
nor U27549 (N_27549,N_27396,N_27292);
and U27550 (N_27550,N_27309,N_27367);
or U27551 (N_27551,N_27105,N_27473);
nand U27552 (N_27552,N_27196,N_27408);
nand U27553 (N_27553,N_27479,N_27474);
and U27554 (N_27554,N_27283,N_27060);
nor U27555 (N_27555,N_27320,N_27153);
xor U27556 (N_27556,N_27388,N_27118);
and U27557 (N_27557,N_27445,N_27406);
nand U27558 (N_27558,N_27205,N_27265);
and U27559 (N_27559,N_27215,N_27072);
nand U27560 (N_27560,N_27003,N_27483);
nor U27561 (N_27561,N_27363,N_27425);
nor U27562 (N_27562,N_27202,N_27167);
xnor U27563 (N_27563,N_27459,N_27078);
xnor U27564 (N_27564,N_27297,N_27235);
or U27565 (N_27565,N_27219,N_27260);
nor U27566 (N_27566,N_27180,N_27381);
or U27567 (N_27567,N_27400,N_27361);
nor U27568 (N_27568,N_27401,N_27116);
nand U27569 (N_27569,N_27130,N_27316);
nor U27570 (N_27570,N_27418,N_27177);
nor U27571 (N_27571,N_27140,N_27492);
nor U27572 (N_27572,N_27107,N_27188);
or U27573 (N_27573,N_27475,N_27049);
or U27574 (N_27574,N_27182,N_27249);
xnor U27575 (N_27575,N_27186,N_27448);
xnor U27576 (N_27576,N_27471,N_27321);
or U27577 (N_27577,N_27484,N_27168);
or U27578 (N_27578,N_27334,N_27127);
nand U27579 (N_27579,N_27467,N_27338);
xnor U27580 (N_27580,N_27437,N_27005);
or U27581 (N_27581,N_27183,N_27106);
xor U27582 (N_27582,N_27356,N_27075);
xnor U27583 (N_27583,N_27047,N_27399);
and U27584 (N_27584,N_27229,N_27199);
or U27585 (N_27585,N_27262,N_27068);
and U27586 (N_27586,N_27456,N_27014);
and U27587 (N_27587,N_27371,N_27236);
or U27588 (N_27588,N_27138,N_27482);
nand U27589 (N_27589,N_27463,N_27044);
xnor U27590 (N_27590,N_27023,N_27093);
and U27591 (N_27591,N_27423,N_27086);
nor U27592 (N_27592,N_27489,N_27045);
and U27593 (N_27593,N_27210,N_27089);
and U27594 (N_27594,N_27449,N_27458);
and U27595 (N_27595,N_27243,N_27357);
nor U27596 (N_27596,N_27244,N_27073);
xnor U27597 (N_27597,N_27439,N_27165);
and U27598 (N_27598,N_27436,N_27407);
xor U27599 (N_27599,N_27119,N_27246);
or U27600 (N_27600,N_27304,N_27175);
nand U27601 (N_27601,N_27143,N_27018);
and U27602 (N_27602,N_27149,N_27147);
nor U27603 (N_27603,N_27499,N_27056);
xnor U27604 (N_27604,N_27099,N_27275);
nand U27605 (N_27605,N_27189,N_27261);
or U27606 (N_27606,N_27000,N_27035);
nand U27607 (N_27607,N_27278,N_27477);
and U27608 (N_27608,N_27051,N_27485);
or U27609 (N_27609,N_27368,N_27455);
nor U27610 (N_27610,N_27402,N_27090);
or U27611 (N_27611,N_27211,N_27050);
nand U27612 (N_27612,N_27442,N_27220);
or U27613 (N_27613,N_27296,N_27240);
nor U27614 (N_27614,N_27163,N_27409);
and U27615 (N_27615,N_27344,N_27364);
nor U27616 (N_27616,N_27111,N_27312);
nand U27617 (N_27617,N_27065,N_27123);
or U27618 (N_27618,N_27339,N_27129);
nand U27619 (N_27619,N_27382,N_27310);
nand U27620 (N_27620,N_27386,N_27317);
nand U27621 (N_27621,N_27124,N_27410);
nand U27622 (N_27622,N_27446,N_27405);
nor U27623 (N_27623,N_27464,N_27080);
nor U27624 (N_27624,N_27259,N_27302);
nor U27625 (N_27625,N_27084,N_27207);
or U27626 (N_27626,N_27218,N_27092);
xor U27627 (N_27627,N_27313,N_27303);
or U27628 (N_27628,N_27480,N_27227);
and U27629 (N_27629,N_27335,N_27258);
nand U27630 (N_27630,N_27429,N_27179);
nor U27631 (N_27631,N_27209,N_27110);
or U27632 (N_27632,N_27340,N_27046);
xnor U27633 (N_27633,N_27039,N_27372);
nor U27634 (N_27634,N_27057,N_27216);
and U27635 (N_27635,N_27457,N_27172);
or U27636 (N_27636,N_27453,N_27132);
nor U27637 (N_27637,N_27131,N_27169);
and U27638 (N_27638,N_27257,N_27450);
and U27639 (N_27639,N_27101,N_27155);
and U27640 (N_27640,N_27268,N_27135);
nor U27641 (N_27641,N_27041,N_27150);
or U27642 (N_27642,N_27019,N_27413);
nand U27643 (N_27643,N_27193,N_27337);
and U27644 (N_27644,N_27162,N_27016);
xnor U27645 (N_27645,N_27034,N_27362);
nor U27646 (N_27646,N_27198,N_27224);
nand U27647 (N_27647,N_27497,N_27359);
xnor U27648 (N_27648,N_27024,N_27447);
nor U27649 (N_27649,N_27067,N_27342);
nor U27650 (N_27650,N_27360,N_27431);
and U27651 (N_27651,N_27237,N_27380);
nand U27652 (N_27652,N_27404,N_27349);
and U27653 (N_27653,N_27025,N_27208);
nor U27654 (N_27654,N_27213,N_27369);
nand U27655 (N_27655,N_27173,N_27200);
and U27656 (N_27656,N_27160,N_27322);
nand U27657 (N_27657,N_27494,N_27393);
or U27658 (N_27658,N_27384,N_27378);
nor U27659 (N_27659,N_27416,N_27478);
nand U27660 (N_27660,N_27146,N_27375);
xnor U27661 (N_27661,N_27203,N_27226);
or U27662 (N_27662,N_27097,N_27008);
or U27663 (N_27663,N_27277,N_27422);
nor U27664 (N_27664,N_27496,N_27379);
nor U27665 (N_27665,N_27486,N_27398);
nand U27666 (N_27666,N_27066,N_27242);
nand U27667 (N_27667,N_27083,N_27451);
nor U27668 (N_27668,N_27100,N_27232);
nor U27669 (N_27669,N_27347,N_27231);
nor U27670 (N_27670,N_27017,N_27255);
and U27671 (N_27671,N_27033,N_27108);
nor U27672 (N_27672,N_27440,N_27085);
or U27673 (N_27673,N_27161,N_27206);
or U27674 (N_27674,N_27095,N_27417);
nor U27675 (N_27675,N_27298,N_27088);
nor U27676 (N_27676,N_27286,N_27419);
or U27677 (N_27677,N_27054,N_27103);
nor U27678 (N_27678,N_27318,N_27319);
nor U27679 (N_27679,N_27267,N_27374);
xor U27680 (N_27680,N_27341,N_27052);
nor U27681 (N_27681,N_27285,N_27330);
nor U27682 (N_27682,N_27272,N_27064);
or U27683 (N_27683,N_27291,N_27062);
and U27684 (N_27684,N_27126,N_27133);
nor U27685 (N_27685,N_27238,N_27426);
and U27686 (N_27686,N_27331,N_27333);
nand U27687 (N_27687,N_27204,N_27411);
nand U27688 (N_27688,N_27171,N_27307);
nand U27689 (N_27689,N_27254,N_27420);
nor U27690 (N_27690,N_27273,N_27137);
or U27691 (N_27691,N_27314,N_27288);
nor U27692 (N_27692,N_27141,N_27366);
nand U27693 (N_27693,N_27069,N_27256);
and U27694 (N_27694,N_27270,N_27282);
xnor U27695 (N_27695,N_27148,N_27376);
nor U27696 (N_27696,N_27412,N_27248);
nand U27697 (N_27697,N_27040,N_27266);
nor U27698 (N_27698,N_27029,N_27026);
nor U27699 (N_27699,N_27145,N_27191);
or U27700 (N_27700,N_27115,N_27289);
xnor U27701 (N_27701,N_27395,N_27223);
or U27702 (N_27702,N_27387,N_27006);
and U27703 (N_27703,N_27495,N_27136);
xnor U27704 (N_27704,N_27170,N_27438);
nor U27705 (N_27705,N_27020,N_27394);
nor U27706 (N_27706,N_27377,N_27245);
nand U27707 (N_27707,N_27176,N_27194);
nor U27708 (N_27708,N_27263,N_27276);
or U27709 (N_27709,N_27241,N_27279);
or U27710 (N_27710,N_27452,N_27217);
and U27711 (N_27711,N_27355,N_27214);
or U27712 (N_27712,N_27332,N_27096);
or U27713 (N_27713,N_27348,N_27281);
nor U27714 (N_27714,N_27031,N_27002);
or U27715 (N_27715,N_27239,N_27325);
and U27716 (N_27716,N_27383,N_27336);
and U27717 (N_27717,N_27037,N_27063);
nand U27718 (N_27718,N_27433,N_27487);
or U27719 (N_27719,N_27094,N_27294);
nor U27720 (N_27720,N_27042,N_27082);
or U27721 (N_27721,N_27142,N_27187);
nor U27722 (N_27722,N_27178,N_27151);
nand U27723 (N_27723,N_27152,N_27306);
or U27724 (N_27724,N_27028,N_27365);
nor U27725 (N_27725,N_27443,N_27434);
nand U27726 (N_27726,N_27117,N_27166);
and U27727 (N_27727,N_27011,N_27295);
xor U27728 (N_27728,N_27076,N_27125);
xor U27729 (N_27729,N_27358,N_27048);
and U27730 (N_27730,N_27247,N_27346);
xnor U27731 (N_27731,N_27345,N_27184);
or U27732 (N_27732,N_27441,N_27234);
nor U27733 (N_27733,N_27164,N_27430);
nor U27734 (N_27734,N_27174,N_27007);
nor U27735 (N_27735,N_27081,N_27350);
or U27736 (N_27736,N_27353,N_27427);
xor U27737 (N_27737,N_27284,N_27300);
nand U27738 (N_27738,N_27159,N_27390);
xnor U27739 (N_27739,N_27392,N_27201);
nand U27740 (N_27740,N_27469,N_27074);
or U27741 (N_27741,N_27328,N_27274);
or U27742 (N_27742,N_27481,N_27476);
or U27743 (N_27743,N_27324,N_27264);
xor U27744 (N_27744,N_27385,N_27077);
xnor U27745 (N_27745,N_27061,N_27004);
and U27746 (N_27746,N_27354,N_27428);
or U27747 (N_27747,N_27058,N_27195);
and U27748 (N_27748,N_27192,N_27326);
nand U27749 (N_27749,N_27461,N_27465);
or U27750 (N_27750,N_27032,N_27432);
or U27751 (N_27751,N_27034,N_27485);
xnor U27752 (N_27752,N_27347,N_27128);
nand U27753 (N_27753,N_27010,N_27300);
nand U27754 (N_27754,N_27274,N_27449);
nor U27755 (N_27755,N_27247,N_27042);
nor U27756 (N_27756,N_27078,N_27254);
xor U27757 (N_27757,N_27388,N_27130);
nor U27758 (N_27758,N_27280,N_27069);
nand U27759 (N_27759,N_27367,N_27364);
xor U27760 (N_27760,N_27349,N_27337);
xor U27761 (N_27761,N_27462,N_27454);
xnor U27762 (N_27762,N_27428,N_27478);
nor U27763 (N_27763,N_27206,N_27191);
xor U27764 (N_27764,N_27032,N_27477);
nor U27765 (N_27765,N_27142,N_27280);
nand U27766 (N_27766,N_27413,N_27372);
xnor U27767 (N_27767,N_27350,N_27488);
and U27768 (N_27768,N_27040,N_27420);
and U27769 (N_27769,N_27443,N_27440);
nor U27770 (N_27770,N_27482,N_27483);
nor U27771 (N_27771,N_27135,N_27173);
nor U27772 (N_27772,N_27183,N_27246);
or U27773 (N_27773,N_27105,N_27065);
nand U27774 (N_27774,N_27262,N_27337);
nand U27775 (N_27775,N_27176,N_27096);
nor U27776 (N_27776,N_27360,N_27225);
and U27777 (N_27777,N_27391,N_27199);
xnor U27778 (N_27778,N_27312,N_27432);
nor U27779 (N_27779,N_27205,N_27211);
or U27780 (N_27780,N_27385,N_27166);
nor U27781 (N_27781,N_27460,N_27348);
or U27782 (N_27782,N_27160,N_27130);
or U27783 (N_27783,N_27099,N_27286);
nor U27784 (N_27784,N_27141,N_27028);
or U27785 (N_27785,N_27049,N_27366);
and U27786 (N_27786,N_27341,N_27372);
and U27787 (N_27787,N_27371,N_27169);
or U27788 (N_27788,N_27133,N_27189);
xnor U27789 (N_27789,N_27225,N_27252);
or U27790 (N_27790,N_27439,N_27032);
nand U27791 (N_27791,N_27255,N_27390);
and U27792 (N_27792,N_27138,N_27226);
nor U27793 (N_27793,N_27470,N_27302);
nor U27794 (N_27794,N_27250,N_27102);
and U27795 (N_27795,N_27247,N_27208);
and U27796 (N_27796,N_27267,N_27093);
xor U27797 (N_27797,N_27019,N_27361);
nor U27798 (N_27798,N_27271,N_27045);
and U27799 (N_27799,N_27067,N_27359);
xor U27800 (N_27800,N_27224,N_27048);
or U27801 (N_27801,N_27030,N_27091);
and U27802 (N_27802,N_27052,N_27277);
nand U27803 (N_27803,N_27366,N_27452);
nor U27804 (N_27804,N_27128,N_27305);
xor U27805 (N_27805,N_27288,N_27154);
nor U27806 (N_27806,N_27402,N_27144);
or U27807 (N_27807,N_27134,N_27170);
xor U27808 (N_27808,N_27101,N_27023);
nor U27809 (N_27809,N_27107,N_27346);
or U27810 (N_27810,N_27147,N_27167);
xnor U27811 (N_27811,N_27302,N_27069);
or U27812 (N_27812,N_27238,N_27395);
nor U27813 (N_27813,N_27156,N_27150);
nand U27814 (N_27814,N_27153,N_27023);
nand U27815 (N_27815,N_27143,N_27172);
xor U27816 (N_27816,N_27200,N_27245);
nand U27817 (N_27817,N_27254,N_27164);
and U27818 (N_27818,N_27135,N_27346);
xor U27819 (N_27819,N_27401,N_27246);
or U27820 (N_27820,N_27013,N_27145);
nand U27821 (N_27821,N_27027,N_27237);
nor U27822 (N_27822,N_27400,N_27119);
xnor U27823 (N_27823,N_27379,N_27053);
xnor U27824 (N_27824,N_27187,N_27305);
and U27825 (N_27825,N_27367,N_27053);
nor U27826 (N_27826,N_27032,N_27427);
or U27827 (N_27827,N_27408,N_27434);
or U27828 (N_27828,N_27306,N_27040);
nor U27829 (N_27829,N_27168,N_27448);
and U27830 (N_27830,N_27149,N_27166);
or U27831 (N_27831,N_27491,N_27087);
xnor U27832 (N_27832,N_27314,N_27079);
nand U27833 (N_27833,N_27333,N_27298);
and U27834 (N_27834,N_27488,N_27043);
nand U27835 (N_27835,N_27170,N_27492);
nor U27836 (N_27836,N_27160,N_27440);
xnor U27837 (N_27837,N_27369,N_27030);
xor U27838 (N_27838,N_27320,N_27095);
or U27839 (N_27839,N_27173,N_27300);
or U27840 (N_27840,N_27001,N_27178);
xnor U27841 (N_27841,N_27306,N_27012);
nand U27842 (N_27842,N_27331,N_27163);
nand U27843 (N_27843,N_27066,N_27074);
xor U27844 (N_27844,N_27108,N_27421);
nand U27845 (N_27845,N_27330,N_27273);
or U27846 (N_27846,N_27108,N_27455);
xnor U27847 (N_27847,N_27164,N_27077);
nand U27848 (N_27848,N_27315,N_27264);
or U27849 (N_27849,N_27415,N_27112);
and U27850 (N_27850,N_27087,N_27048);
and U27851 (N_27851,N_27035,N_27049);
nand U27852 (N_27852,N_27097,N_27115);
xnor U27853 (N_27853,N_27403,N_27474);
xor U27854 (N_27854,N_27131,N_27163);
nor U27855 (N_27855,N_27471,N_27172);
xor U27856 (N_27856,N_27333,N_27139);
xor U27857 (N_27857,N_27133,N_27111);
nor U27858 (N_27858,N_27242,N_27341);
xnor U27859 (N_27859,N_27083,N_27268);
nand U27860 (N_27860,N_27304,N_27270);
or U27861 (N_27861,N_27360,N_27018);
nor U27862 (N_27862,N_27226,N_27019);
nand U27863 (N_27863,N_27247,N_27037);
nor U27864 (N_27864,N_27117,N_27028);
or U27865 (N_27865,N_27376,N_27265);
nand U27866 (N_27866,N_27453,N_27335);
nor U27867 (N_27867,N_27054,N_27164);
nand U27868 (N_27868,N_27449,N_27172);
nor U27869 (N_27869,N_27364,N_27470);
nand U27870 (N_27870,N_27282,N_27344);
or U27871 (N_27871,N_27036,N_27047);
or U27872 (N_27872,N_27283,N_27348);
xor U27873 (N_27873,N_27434,N_27283);
nand U27874 (N_27874,N_27187,N_27424);
and U27875 (N_27875,N_27178,N_27090);
or U27876 (N_27876,N_27472,N_27197);
nand U27877 (N_27877,N_27362,N_27354);
xnor U27878 (N_27878,N_27297,N_27279);
and U27879 (N_27879,N_27268,N_27059);
xor U27880 (N_27880,N_27422,N_27197);
nor U27881 (N_27881,N_27245,N_27202);
or U27882 (N_27882,N_27285,N_27047);
or U27883 (N_27883,N_27285,N_27459);
nor U27884 (N_27884,N_27152,N_27199);
nand U27885 (N_27885,N_27228,N_27340);
nand U27886 (N_27886,N_27088,N_27177);
xnor U27887 (N_27887,N_27115,N_27426);
xnor U27888 (N_27888,N_27289,N_27181);
xnor U27889 (N_27889,N_27088,N_27059);
nor U27890 (N_27890,N_27091,N_27447);
nand U27891 (N_27891,N_27435,N_27466);
nor U27892 (N_27892,N_27156,N_27183);
xnor U27893 (N_27893,N_27204,N_27109);
nor U27894 (N_27894,N_27034,N_27432);
nand U27895 (N_27895,N_27381,N_27089);
xnor U27896 (N_27896,N_27484,N_27464);
or U27897 (N_27897,N_27498,N_27404);
nor U27898 (N_27898,N_27278,N_27249);
or U27899 (N_27899,N_27288,N_27067);
nand U27900 (N_27900,N_27096,N_27017);
xnor U27901 (N_27901,N_27402,N_27143);
and U27902 (N_27902,N_27054,N_27354);
nand U27903 (N_27903,N_27021,N_27244);
xor U27904 (N_27904,N_27410,N_27279);
and U27905 (N_27905,N_27219,N_27411);
nand U27906 (N_27906,N_27457,N_27003);
nor U27907 (N_27907,N_27331,N_27323);
or U27908 (N_27908,N_27392,N_27452);
and U27909 (N_27909,N_27198,N_27394);
xnor U27910 (N_27910,N_27426,N_27474);
and U27911 (N_27911,N_27343,N_27351);
nand U27912 (N_27912,N_27394,N_27288);
xor U27913 (N_27913,N_27113,N_27482);
and U27914 (N_27914,N_27114,N_27147);
nand U27915 (N_27915,N_27049,N_27030);
and U27916 (N_27916,N_27030,N_27276);
or U27917 (N_27917,N_27316,N_27064);
nand U27918 (N_27918,N_27213,N_27178);
xor U27919 (N_27919,N_27133,N_27068);
or U27920 (N_27920,N_27189,N_27497);
nor U27921 (N_27921,N_27011,N_27414);
or U27922 (N_27922,N_27047,N_27049);
or U27923 (N_27923,N_27393,N_27369);
xnor U27924 (N_27924,N_27394,N_27003);
xor U27925 (N_27925,N_27028,N_27423);
nand U27926 (N_27926,N_27167,N_27056);
nor U27927 (N_27927,N_27209,N_27249);
nand U27928 (N_27928,N_27082,N_27075);
xnor U27929 (N_27929,N_27153,N_27013);
nand U27930 (N_27930,N_27167,N_27008);
and U27931 (N_27931,N_27258,N_27293);
nand U27932 (N_27932,N_27409,N_27045);
or U27933 (N_27933,N_27108,N_27366);
or U27934 (N_27934,N_27229,N_27013);
xnor U27935 (N_27935,N_27347,N_27422);
and U27936 (N_27936,N_27498,N_27175);
or U27937 (N_27937,N_27335,N_27497);
nand U27938 (N_27938,N_27099,N_27070);
or U27939 (N_27939,N_27182,N_27421);
xnor U27940 (N_27940,N_27369,N_27288);
nand U27941 (N_27941,N_27312,N_27436);
nand U27942 (N_27942,N_27496,N_27463);
xor U27943 (N_27943,N_27414,N_27365);
and U27944 (N_27944,N_27321,N_27466);
and U27945 (N_27945,N_27260,N_27463);
xnor U27946 (N_27946,N_27470,N_27332);
or U27947 (N_27947,N_27191,N_27337);
and U27948 (N_27948,N_27191,N_27365);
or U27949 (N_27949,N_27423,N_27056);
xnor U27950 (N_27950,N_27454,N_27171);
and U27951 (N_27951,N_27215,N_27018);
xor U27952 (N_27952,N_27435,N_27392);
or U27953 (N_27953,N_27270,N_27307);
nor U27954 (N_27954,N_27415,N_27253);
nand U27955 (N_27955,N_27209,N_27365);
xnor U27956 (N_27956,N_27008,N_27180);
xnor U27957 (N_27957,N_27499,N_27002);
and U27958 (N_27958,N_27067,N_27072);
or U27959 (N_27959,N_27276,N_27400);
nand U27960 (N_27960,N_27237,N_27010);
xnor U27961 (N_27961,N_27250,N_27126);
nand U27962 (N_27962,N_27018,N_27430);
or U27963 (N_27963,N_27304,N_27384);
and U27964 (N_27964,N_27001,N_27038);
and U27965 (N_27965,N_27151,N_27284);
and U27966 (N_27966,N_27442,N_27007);
nand U27967 (N_27967,N_27319,N_27148);
xnor U27968 (N_27968,N_27264,N_27044);
nor U27969 (N_27969,N_27421,N_27432);
nand U27970 (N_27970,N_27122,N_27427);
or U27971 (N_27971,N_27219,N_27201);
xor U27972 (N_27972,N_27359,N_27419);
nor U27973 (N_27973,N_27194,N_27263);
or U27974 (N_27974,N_27185,N_27272);
xnor U27975 (N_27975,N_27445,N_27205);
nor U27976 (N_27976,N_27218,N_27320);
and U27977 (N_27977,N_27434,N_27070);
xor U27978 (N_27978,N_27429,N_27364);
and U27979 (N_27979,N_27260,N_27255);
xnor U27980 (N_27980,N_27028,N_27005);
nor U27981 (N_27981,N_27407,N_27499);
nand U27982 (N_27982,N_27152,N_27244);
nor U27983 (N_27983,N_27026,N_27225);
or U27984 (N_27984,N_27105,N_27015);
nor U27985 (N_27985,N_27436,N_27150);
or U27986 (N_27986,N_27163,N_27174);
or U27987 (N_27987,N_27061,N_27062);
or U27988 (N_27988,N_27435,N_27338);
nand U27989 (N_27989,N_27198,N_27253);
and U27990 (N_27990,N_27004,N_27357);
xor U27991 (N_27991,N_27155,N_27226);
nor U27992 (N_27992,N_27159,N_27116);
nor U27993 (N_27993,N_27258,N_27488);
or U27994 (N_27994,N_27310,N_27026);
nand U27995 (N_27995,N_27396,N_27191);
or U27996 (N_27996,N_27498,N_27148);
nand U27997 (N_27997,N_27413,N_27332);
or U27998 (N_27998,N_27313,N_27228);
and U27999 (N_27999,N_27123,N_27455);
nor U28000 (N_28000,N_27865,N_27772);
or U28001 (N_28001,N_27970,N_27948);
nor U28002 (N_28002,N_27935,N_27712);
nor U28003 (N_28003,N_27543,N_27907);
or U28004 (N_28004,N_27546,N_27963);
xor U28005 (N_28005,N_27657,N_27628);
or U28006 (N_28006,N_27651,N_27564);
xor U28007 (N_28007,N_27593,N_27547);
and U28008 (N_28008,N_27957,N_27888);
nor U28009 (N_28009,N_27811,N_27558);
or U28010 (N_28010,N_27678,N_27581);
or U28011 (N_28011,N_27579,N_27909);
nor U28012 (N_28012,N_27642,N_27713);
and U28013 (N_28013,N_27889,N_27655);
or U28014 (N_28014,N_27809,N_27896);
and U28015 (N_28015,N_27760,N_27727);
nor U28016 (N_28016,N_27683,N_27803);
and U28017 (N_28017,N_27956,N_27597);
and U28018 (N_28018,N_27568,N_27603);
nand U28019 (N_28019,N_27578,N_27753);
nand U28020 (N_28020,N_27658,N_27652);
nand U28021 (N_28021,N_27518,N_27924);
xor U28022 (N_28022,N_27976,N_27859);
xor U28023 (N_28023,N_27592,N_27737);
and U28024 (N_28024,N_27511,N_27993);
nor U28025 (N_28025,N_27696,N_27904);
and U28026 (N_28026,N_27875,N_27599);
or U28027 (N_28027,N_27750,N_27835);
xor U28028 (N_28028,N_27960,N_27653);
or U28029 (N_28029,N_27726,N_27707);
xnor U28030 (N_28030,N_27650,N_27685);
xnor U28031 (N_28031,N_27893,N_27885);
xnor U28032 (N_28032,N_27602,N_27919);
or U28033 (N_28033,N_27758,N_27596);
and U28034 (N_28034,N_27953,N_27998);
nand U28035 (N_28035,N_27855,N_27699);
and U28036 (N_28036,N_27669,N_27590);
or U28037 (N_28037,N_27792,N_27806);
nand U28038 (N_28038,N_27867,N_27580);
nor U28039 (N_28039,N_27979,N_27775);
or U28040 (N_28040,N_27744,N_27507);
or U28041 (N_28041,N_27981,N_27987);
xnor U28042 (N_28042,N_27673,N_27857);
nor U28043 (N_28043,N_27627,N_27873);
nand U28044 (N_28044,N_27980,N_27691);
nor U28045 (N_28045,N_27955,N_27954);
nand U28046 (N_28046,N_27519,N_27598);
nor U28047 (N_28047,N_27688,N_27938);
or U28048 (N_28048,N_27986,N_27572);
or U28049 (N_28049,N_27636,N_27648);
nand U28050 (N_28050,N_27508,N_27622);
nand U28051 (N_28051,N_27609,N_27585);
xnor U28052 (N_28052,N_27730,N_27894);
and U28053 (N_28053,N_27798,N_27520);
nand U28054 (N_28054,N_27757,N_27670);
nor U28055 (N_28055,N_27552,N_27567);
and U28056 (N_28056,N_27698,N_27640);
and U28057 (N_28057,N_27780,N_27969);
nand U28058 (N_28058,N_27706,N_27719);
or U28059 (N_28059,N_27765,N_27689);
or U28060 (N_28060,N_27529,N_27914);
xor U28061 (N_28061,N_27635,N_27851);
and U28062 (N_28062,N_27812,N_27883);
nand U28063 (N_28063,N_27509,N_27607);
nor U28064 (N_28064,N_27560,N_27790);
nor U28065 (N_28065,N_27756,N_27671);
nor U28066 (N_28066,N_27510,N_27537);
or U28067 (N_28067,N_27825,N_27837);
and U28068 (N_28068,N_27928,N_27664);
or U28069 (N_28069,N_27731,N_27800);
nand U28070 (N_28070,N_27831,N_27512);
xor U28071 (N_28071,N_27649,N_27668);
nand U28072 (N_28072,N_27697,N_27967);
nor U28073 (N_28073,N_27754,N_27677);
nor U28074 (N_28074,N_27912,N_27763);
nor U28075 (N_28075,N_27982,N_27899);
xnor U28076 (N_28076,N_27992,N_27538);
nand U28077 (N_28077,N_27715,N_27864);
nor U28078 (N_28078,N_27788,N_27524);
or U28079 (N_28079,N_27561,N_27815);
xor U28080 (N_28080,N_27556,N_27702);
nand U28081 (N_28081,N_27751,N_27946);
xor U28082 (N_28082,N_27692,N_27571);
nor U28083 (N_28083,N_27903,N_27900);
xnor U28084 (N_28084,N_27583,N_27791);
and U28085 (N_28085,N_27968,N_27921);
xnor U28086 (N_28086,N_27641,N_27724);
xnor U28087 (N_28087,N_27634,N_27600);
nor U28088 (N_28088,N_27879,N_27708);
nor U28089 (N_28089,N_27931,N_27770);
xnor U28090 (N_28090,N_27844,N_27858);
nand U28091 (N_28091,N_27725,N_27539);
or U28092 (N_28092,N_27728,N_27714);
and U28093 (N_28093,N_27872,N_27916);
nor U28094 (N_28094,N_27774,N_27762);
nand U28095 (N_28095,N_27802,N_27704);
nand U28096 (N_28096,N_27804,N_27613);
and U28097 (N_28097,N_27745,N_27974);
and U28098 (N_28098,N_27676,N_27828);
xor U28099 (N_28099,N_27794,N_27781);
nand U28100 (N_28100,N_27908,N_27682);
nand U28101 (N_28101,N_27755,N_27612);
nand U28102 (N_28102,N_27892,N_27942);
xnor U28103 (N_28103,N_27722,N_27782);
or U28104 (N_28104,N_27711,N_27742);
or U28105 (N_28105,N_27620,N_27686);
xor U28106 (N_28106,N_27501,N_27795);
xnor U28107 (N_28107,N_27608,N_27723);
and U28108 (N_28108,N_27523,N_27884);
xnor U28109 (N_28109,N_27965,N_27853);
nor U28110 (N_28110,N_27550,N_27710);
nand U28111 (N_28111,N_27674,N_27531);
nor U28112 (N_28112,N_27930,N_27721);
and U28113 (N_28113,N_27932,N_27882);
xnor U28114 (N_28114,N_27662,N_27874);
or U28115 (N_28115,N_27748,N_27623);
nand U28116 (N_28116,N_27517,N_27793);
nor U28117 (N_28117,N_27771,N_27820);
or U28118 (N_28118,N_27852,N_27766);
nor U28119 (N_28119,N_27565,N_27759);
nor U28120 (N_28120,N_27705,N_27933);
and U28121 (N_28121,N_27506,N_27513);
or U28122 (N_28122,N_27551,N_27749);
xor U28123 (N_28123,N_27500,N_27663);
nor U28124 (N_28124,N_27736,N_27557);
nor U28125 (N_28125,N_27923,N_27665);
nand U28126 (N_28126,N_27584,N_27962);
nor U28127 (N_28127,N_27569,N_27972);
xor U28128 (N_28128,N_27505,N_27562);
nand U28129 (N_28129,N_27880,N_27553);
and U28130 (N_28130,N_27514,N_27961);
or U28131 (N_28131,N_27783,N_27675);
xnor U28132 (N_28132,N_27667,N_27866);
nor U28133 (N_28133,N_27784,N_27843);
nand U28134 (N_28134,N_27776,N_27936);
or U28135 (N_28135,N_27536,N_27839);
and U28136 (N_28136,N_27822,N_27611);
nor U28137 (N_28137,N_27922,N_27545);
or U28138 (N_28138,N_27890,N_27847);
nor U28139 (N_28139,N_27540,N_27720);
or U28140 (N_28140,N_27973,N_27577);
or U28141 (N_28141,N_27595,N_27637);
or U28142 (N_28142,N_27827,N_27703);
xnor U28143 (N_28143,N_27548,N_27700);
nand U28144 (N_28144,N_27787,N_27824);
and U28145 (N_28145,N_27841,N_27810);
xor U28146 (N_28146,N_27639,N_27530);
nor U28147 (N_28147,N_27939,N_27582);
or U28148 (N_28148,N_27818,N_27575);
or U28149 (N_28149,N_27631,N_27937);
nand U28150 (N_28150,N_27990,N_27846);
xnor U28151 (N_28151,N_27918,N_27868);
or U28152 (N_28152,N_27528,N_27958);
xor U28153 (N_28153,N_27816,N_27616);
and U28154 (N_28154,N_27555,N_27945);
or U28155 (N_28155,N_27779,N_27615);
or U28156 (N_28156,N_27959,N_27944);
and U28157 (N_28157,N_27601,N_27949);
or U28158 (N_28158,N_27848,N_27834);
nor U28159 (N_28159,N_27638,N_27729);
xor U28160 (N_28160,N_27913,N_27854);
nand U28161 (N_28161,N_27629,N_27738);
or U28162 (N_28162,N_27764,N_27709);
xnor U28163 (N_28163,N_27610,N_27660);
nor U28164 (N_28164,N_27645,N_27680);
or U28165 (N_28165,N_27566,N_27805);
and U28166 (N_28166,N_27898,N_27984);
nor U28167 (N_28167,N_27503,N_27951);
and U28168 (N_28168,N_27814,N_27643);
nor U28169 (N_28169,N_27504,N_27886);
and U28170 (N_28170,N_27534,N_27861);
and U28171 (N_28171,N_27574,N_27617);
nor U28172 (N_28172,N_27717,N_27849);
nor U28173 (N_28173,N_27767,N_27606);
and U28174 (N_28174,N_27701,N_27694);
and U28175 (N_28175,N_27971,N_27807);
nor U28176 (N_28176,N_27785,N_27842);
nor U28177 (N_28177,N_27910,N_27777);
nor U28178 (N_28178,N_27752,N_27625);
and U28179 (N_28179,N_27789,N_27587);
nand U28180 (N_28180,N_27718,N_27915);
and U28181 (N_28181,N_27747,N_27860);
and U28182 (N_28182,N_27654,N_27521);
or U28183 (N_28183,N_27821,N_27619);
and U28184 (N_28184,N_27813,N_27988);
nor U28185 (N_28185,N_27515,N_27690);
nand U28186 (N_28186,N_27605,N_27687);
or U28187 (N_28187,N_27927,N_27527);
nand U28188 (N_28188,N_27659,N_27902);
xor U28189 (N_28189,N_27533,N_27934);
nand U28190 (N_28190,N_27773,N_27526);
and U28191 (N_28191,N_27950,N_27836);
xnor U28192 (N_28192,N_27502,N_27870);
nor U28193 (N_28193,N_27819,N_27863);
nor U28194 (N_28194,N_27850,N_27733);
nand U28195 (N_28195,N_27549,N_27830);
nor U28196 (N_28196,N_27522,N_27532);
or U28197 (N_28197,N_27646,N_27632);
nand U28198 (N_28198,N_27845,N_27877);
or U28199 (N_28199,N_27554,N_27693);
nor U28200 (N_28200,N_27621,N_27679);
nand U28201 (N_28201,N_27786,N_27768);
xor U28202 (N_28202,N_27977,N_27644);
or U28203 (N_28203,N_27535,N_27761);
and U28204 (N_28204,N_27618,N_27741);
nand U28205 (N_28205,N_27559,N_27797);
or U28206 (N_28206,N_27911,N_27684);
nand U28207 (N_28207,N_27833,N_27994);
and U28208 (N_28208,N_27801,N_27897);
or U28209 (N_28209,N_27591,N_27838);
or U28210 (N_28210,N_27589,N_27576);
or U28211 (N_28211,N_27695,N_27624);
and U28212 (N_28212,N_27808,N_27656);
nor U28213 (N_28213,N_27525,N_27862);
or U28214 (N_28214,N_27661,N_27563);
or U28215 (N_28215,N_27991,N_27743);
and U28216 (N_28216,N_27869,N_27966);
xor U28217 (N_28217,N_27633,N_27769);
and U28218 (N_28218,N_27666,N_27941);
or U28219 (N_28219,N_27626,N_27943);
and U28220 (N_28220,N_27732,N_27906);
and U28221 (N_28221,N_27735,N_27544);
xnor U28222 (N_28222,N_27878,N_27516);
xor U28223 (N_28223,N_27542,N_27856);
or U28224 (N_28224,N_27925,N_27995);
xor U28225 (N_28225,N_27840,N_27871);
or U28226 (N_28226,N_27876,N_27604);
xnor U28227 (N_28227,N_27778,N_27926);
nor U28228 (N_28228,N_27887,N_27929);
nand U28229 (N_28229,N_27826,N_27999);
nand U28230 (N_28230,N_27734,N_27978);
nor U28231 (N_28231,N_27829,N_27588);
nor U28232 (N_28232,N_27996,N_27630);
and U28233 (N_28233,N_27881,N_27672);
and U28234 (N_28234,N_27541,N_27964);
nor U28235 (N_28235,N_27570,N_27817);
xor U28236 (N_28236,N_27940,N_27799);
and U28237 (N_28237,N_27740,N_27614);
nor U28238 (N_28238,N_27989,N_27823);
xnor U28239 (N_28239,N_27891,N_27796);
nand U28240 (N_28240,N_27647,N_27952);
or U28241 (N_28241,N_27997,N_27716);
nand U28242 (N_28242,N_27901,N_27983);
and U28243 (N_28243,N_27739,N_27681);
nand U28244 (N_28244,N_27832,N_27985);
and U28245 (N_28245,N_27975,N_27905);
nor U28246 (N_28246,N_27594,N_27920);
or U28247 (N_28247,N_27746,N_27947);
and U28248 (N_28248,N_27573,N_27917);
and U28249 (N_28249,N_27895,N_27586);
or U28250 (N_28250,N_27570,N_27717);
nand U28251 (N_28251,N_27721,N_27851);
and U28252 (N_28252,N_27608,N_27955);
and U28253 (N_28253,N_27656,N_27676);
and U28254 (N_28254,N_27830,N_27960);
or U28255 (N_28255,N_27517,N_27999);
or U28256 (N_28256,N_27612,N_27505);
nor U28257 (N_28257,N_27541,N_27648);
nand U28258 (N_28258,N_27542,N_27502);
or U28259 (N_28259,N_27624,N_27767);
xor U28260 (N_28260,N_27804,N_27790);
nand U28261 (N_28261,N_27722,N_27743);
or U28262 (N_28262,N_27671,N_27943);
xnor U28263 (N_28263,N_27661,N_27643);
nand U28264 (N_28264,N_27829,N_27691);
nor U28265 (N_28265,N_27649,N_27930);
or U28266 (N_28266,N_27770,N_27711);
nor U28267 (N_28267,N_27956,N_27985);
nor U28268 (N_28268,N_27568,N_27616);
nor U28269 (N_28269,N_27795,N_27856);
xor U28270 (N_28270,N_27650,N_27621);
nand U28271 (N_28271,N_27526,N_27906);
and U28272 (N_28272,N_27839,N_27697);
nor U28273 (N_28273,N_27708,N_27817);
xnor U28274 (N_28274,N_27876,N_27906);
nor U28275 (N_28275,N_27540,N_27877);
or U28276 (N_28276,N_27775,N_27688);
nor U28277 (N_28277,N_27506,N_27993);
and U28278 (N_28278,N_27946,N_27776);
nand U28279 (N_28279,N_27518,N_27694);
and U28280 (N_28280,N_27806,N_27922);
and U28281 (N_28281,N_27766,N_27526);
or U28282 (N_28282,N_27532,N_27628);
and U28283 (N_28283,N_27501,N_27805);
nand U28284 (N_28284,N_27841,N_27700);
and U28285 (N_28285,N_27535,N_27541);
xor U28286 (N_28286,N_27810,N_27569);
nor U28287 (N_28287,N_27586,N_27808);
xnor U28288 (N_28288,N_27683,N_27917);
nand U28289 (N_28289,N_27922,N_27990);
nand U28290 (N_28290,N_27628,N_27826);
and U28291 (N_28291,N_27566,N_27533);
or U28292 (N_28292,N_27683,N_27698);
and U28293 (N_28293,N_27844,N_27871);
nor U28294 (N_28294,N_27926,N_27841);
or U28295 (N_28295,N_27725,N_27708);
nor U28296 (N_28296,N_27520,N_27825);
nor U28297 (N_28297,N_27986,N_27724);
and U28298 (N_28298,N_27988,N_27647);
nor U28299 (N_28299,N_27874,N_27608);
nand U28300 (N_28300,N_27950,N_27530);
xnor U28301 (N_28301,N_27628,N_27506);
nand U28302 (N_28302,N_27769,N_27568);
nand U28303 (N_28303,N_27808,N_27583);
nor U28304 (N_28304,N_27549,N_27878);
xnor U28305 (N_28305,N_27554,N_27606);
nand U28306 (N_28306,N_27621,N_27555);
xnor U28307 (N_28307,N_27844,N_27947);
or U28308 (N_28308,N_27591,N_27605);
nand U28309 (N_28309,N_27945,N_27999);
nor U28310 (N_28310,N_27555,N_27938);
or U28311 (N_28311,N_27897,N_27826);
nand U28312 (N_28312,N_27843,N_27501);
nor U28313 (N_28313,N_27707,N_27961);
nand U28314 (N_28314,N_27909,N_27710);
nand U28315 (N_28315,N_27641,N_27779);
or U28316 (N_28316,N_27508,N_27621);
xor U28317 (N_28317,N_27566,N_27898);
nand U28318 (N_28318,N_27873,N_27839);
xor U28319 (N_28319,N_27546,N_27939);
and U28320 (N_28320,N_27749,N_27947);
and U28321 (N_28321,N_27550,N_27853);
or U28322 (N_28322,N_27863,N_27977);
nand U28323 (N_28323,N_27750,N_27648);
and U28324 (N_28324,N_27546,N_27857);
nand U28325 (N_28325,N_27950,N_27703);
and U28326 (N_28326,N_27510,N_27526);
and U28327 (N_28327,N_27894,N_27650);
nor U28328 (N_28328,N_27697,N_27551);
or U28329 (N_28329,N_27577,N_27759);
nor U28330 (N_28330,N_27744,N_27954);
nand U28331 (N_28331,N_27665,N_27718);
nand U28332 (N_28332,N_27985,N_27522);
nor U28333 (N_28333,N_27568,N_27535);
or U28334 (N_28334,N_27671,N_27666);
and U28335 (N_28335,N_27862,N_27645);
xor U28336 (N_28336,N_27630,N_27668);
nor U28337 (N_28337,N_27585,N_27664);
or U28338 (N_28338,N_27802,N_27880);
and U28339 (N_28339,N_27800,N_27641);
nand U28340 (N_28340,N_27968,N_27590);
nand U28341 (N_28341,N_27861,N_27603);
and U28342 (N_28342,N_27626,N_27640);
nor U28343 (N_28343,N_27715,N_27722);
xor U28344 (N_28344,N_27637,N_27587);
nand U28345 (N_28345,N_27907,N_27601);
and U28346 (N_28346,N_27552,N_27518);
and U28347 (N_28347,N_27749,N_27761);
or U28348 (N_28348,N_27998,N_27665);
and U28349 (N_28349,N_27654,N_27869);
xor U28350 (N_28350,N_27823,N_27769);
nor U28351 (N_28351,N_27954,N_27541);
xnor U28352 (N_28352,N_27686,N_27822);
xor U28353 (N_28353,N_27645,N_27997);
xnor U28354 (N_28354,N_27697,N_27670);
nand U28355 (N_28355,N_27916,N_27902);
nor U28356 (N_28356,N_27914,N_27788);
nand U28357 (N_28357,N_27802,N_27763);
and U28358 (N_28358,N_27553,N_27709);
xor U28359 (N_28359,N_27796,N_27808);
nand U28360 (N_28360,N_27956,N_27521);
nor U28361 (N_28361,N_27719,N_27531);
nand U28362 (N_28362,N_27538,N_27808);
xor U28363 (N_28363,N_27925,N_27859);
nand U28364 (N_28364,N_27649,N_27690);
or U28365 (N_28365,N_27607,N_27869);
nand U28366 (N_28366,N_27994,N_27762);
or U28367 (N_28367,N_27933,N_27654);
nand U28368 (N_28368,N_27795,N_27983);
and U28369 (N_28369,N_27824,N_27773);
xnor U28370 (N_28370,N_27593,N_27573);
nand U28371 (N_28371,N_27601,N_27761);
xnor U28372 (N_28372,N_27888,N_27936);
xor U28373 (N_28373,N_27585,N_27741);
or U28374 (N_28374,N_27807,N_27505);
nor U28375 (N_28375,N_27625,N_27952);
xor U28376 (N_28376,N_27805,N_27896);
nor U28377 (N_28377,N_27983,N_27556);
and U28378 (N_28378,N_27848,N_27761);
and U28379 (N_28379,N_27684,N_27986);
nand U28380 (N_28380,N_27980,N_27534);
and U28381 (N_28381,N_27866,N_27979);
or U28382 (N_28382,N_27683,N_27522);
and U28383 (N_28383,N_27781,N_27688);
and U28384 (N_28384,N_27708,N_27537);
nand U28385 (N_28385,N_27629,N_27633);
or U28386 (N_28386,N_27773,N_27700);
nor U28387 (N_28387,N_27781,N_27665);
or U28388 (N_28388,N_27567,N_27622);
nor U28389 (N_28389,N_27970,N_27994);
nand U28390 (N_28390,N_27912,N_27684);
and U28391 (N_28391,N_27577,N_27669);
nand U28392 (N_28392,N_27973,N_27732);
and U28393 (N_28393,N_27603,N_27973);
xor U28394 (N_28394,N_27568,N_27820);
and U28395 (N_28395,N_27535,N_27739);
xnor U28396 (N_28396,N_27950,N_27962);
or U28397 (N_28397,N_27913,N_27511);
or U28398 (N_28398,N_27527,N_27650);
or U28399 (N_28399,N_27996,N_27916);
or U28400 (N_28400,N_27906,N_27787);
and U28401 (N_28401,N_27888,N_27945);
and U28402 (N_28402,N_27721,N_27526);
and U28403 (N_28403,N_27964,N_27707);
nor U28404 (N_28404,N_27650,N_27720);
and U28405 (N_28405,N_27882,N_27942);
nor U28406 (N_28406,N_27655,N_27991);
xnor U28407 (N_28407,N_27745,N_27643);
nand U28408 (N_28408,N_27745,N_27600);
nor U28409 (N_28409,N_27975,N_27925);
and U28410 (N_28410,N_27662,N_27883);
xnor U28411 (N_28411,N_27735,N_27800);
nand U28412 (N_28412,N_27641,N_27658);
nor U28413 (N_28413,N_27882,N_27651);
xor U28414 (N_28414,N_27710,N_27521);
or U28415 (N_28415,N_27714,N_27524);
nor U28416 (N_28416,N_27525,N_27763);
or U28417 (N_28417,N_27890,N_27966);
nand U28418 (N_28418,N_27844,N_27580);
or U28419 (N_28419,N_27918,N_27637);
or U28420 (N_28420,N_27527,N_27832);
xnor U28421 (N_28421,N_27760,N_27577);
and U28422 (N_28422,N_27506,N_27680);
nor U28423 (N_28423,N_27629,N_27639);
or U28424 (N_28424,N_27656,N_27549);
nor U28425 (N_28425,N_27928,N_27896);
and U28426 (N_28426,N_27885,N_27833);
and U28427 (N_28427,N_27812,N_27549);
nor U28428 (N_28428,N_27541,N_27922);
nor U28429 (N_28429,N_27603,N_27667);
nand U28430 (N_28430,N_27946,N_27899);
xor U28431 (N_28431,N_27582,N_27672);
and U28432 (N_28432,N_27706,N_27510);
nand U28433 (N_28433,N_27893,N_27602);
and U28434 (N_28434,N_27886,N_27915);
nand U28435 (N_28435,N_27741,N_27950);
or U28436 (N_28436,N_27622,N_27978);
xnor U28437 (N_28437,N_27790,N_27750);
nand U28438 (N_28438,N_27636,N_27671);
xnor U28439 (N_28439,N_27852,N_27549);
nand U28440 (N_28440,N_27806,N_27813);
nor U28441 (N_28441,N_27972,N_27540);
nor U28442 (N_28442,N_27930,N_27562);
or U28443 (N_28443,N_27595,N_27789);
xnor U28444 (N_28444,N_27785,N_27875);
or U28445 (N_28445,N_27736,N_27756);
or U28446 (N_28446,N_27614,N_27950);
nand U28447 (N_28447,N_27963,N_27969);
or U28448 (N_28448,N_27512,N_27821);
or U28449 (N_28449,N_27864,N_27663);
nor U28450 (N_28450,N_27748,N_27803);
and U28451 (N_28451,N_27880,N_27517);
and U28452 (N_28452,N_27578,N_27584);
or U28453 (N_28453,N_27780,N_27809);
or U28454 (N_28454,N_27768,N_27663);
nor U28455 (N_28455,N_27600,N_27885);
or U28456 (N_28456,N_27609,N_27752);
nor U28457 (N_28457,N_27790,N_27524);
nand U28458 (N_28458,N_27745,N_27911);
or U28459 (N_28459,N_27542,N_27533);
xnor U28460 (N_28460,N_27613,N_27746);
and U28461 (N_28461,N_27605,N_27840);
nor U28462 (N_28462,N_27926,N_27591);
nand U28463 (N_28463,N_27931,N_27698);
and U28464 (N_28464,N_27817,N_27739);
nand U28465 (N_28465,N_27579,N_27728);
xnor U28466 (N_28466,N_27995,N_27644);
or U28467 (N_28467,N_27629,N_27998);
nand U28468 (N_28468,N_27788,N_27545);
xnor U28469 (N_28469,N_27915,N_27984);
nor U28470 (N_28470,N_27768,N_27839);
xor U28471 (N_28471,N_27635,N_27775);
and U28472 (N_28472,N_27860,N_27744);
nor U28473 (N_28473,N_27900,N_27862);
xor U28474 (N_28474,N_27644,N_27534);
nor U28475 (N_28475,N_27677,N_27812);
and U28476 (N_28476,N_27656,N_27740);
or U28477 (N_28477,N_27543,N_27837);
nand U28478 (N_28478,N_27874,N_27791);
and U28479 (N_28479,N_27974,N_27747);
nand U28480 (N_28480,N_27821,N_27763);
nand U28481 (N_28481,N_27810,N_27908);
xor U28482 (N_28482,N_27610,N_27799);
and U28483 (N_28483,N_27862,N_27682);
or U28484 (N_28484,N_27736,N_27811);
nand U28485 (N_28485,N_27770,N_27893);
xnor U28486 (N_28486,N_27583,N_27699);
and U28487 (N_28487,N_27832,N_27908);
or U28488 (N_28488,N_27989,N_27748);
or U28489 (N_28489,N_27997,N_27849);
or U28490 (N_28490,N_27903,N_27627);
nand U28491 (N_28491,N_27972,N_27768);
or U28492 (N_28492,N_27599,N_27861);
nand U28493 (N_28493,N_27962,N_27628);
nor U28494 (N_28494,N_27928,N_27887);
nor U28495 (N_28495,N_27568,N_27691);
nand U28496 (N_28496,N_27941,N_27937);
or U28497 (N_28497,N_27768,N_27601);
nand U28498 (N_28498,N_27701,N_27921);
or U28499 (N_28499,N_27772,N_27726);
xnor U28500 (N_28500,N_28137,N_28089);
xnor U28501 (N_28501,N_28440,N_28378);
xnor U28502 (N_28502,N_28070,N_28004);
nor U28503 (N_28503,N_28125,N_28062);
nand U28504 (N_28504,N_28059,N_28422);
xor U28505 (N_28505,N_28131,N_28006);
xnor U28506 (N_28506,N_28161,N_28297);
xor U28507 (N_28507,N_28199,N_28118);
or U28508 (N_28508,N_28088,N_28415);
and U28509 (N_28509,N_28428,N_28323);
xnor U28510 (N_28510,N_28108,N_28110);
nand U28511 (N_28511,N_28265,N_28010);
and U28512 (N_28512,N_28171,N_28106);
nor U28513 (N_28513,N_28365,N_28429);
xnor U28514 (N_28514,N_28310,N_28348);
and U28515 (N_28515,N_28166,N_28233);
and U28516 (N_28516,N_28359,N_28256);
xor U28517 (N_28517,N_28068,N_28178);
nand U28518 (N_28518,N_28225,N_28040);
nor U28519 (N_28519,N_28017,N_28201);
xor U28520 (N_28520,N_28305,N_28212);
xnor U28521 (N_28521,N_28269,N_28044);
nand U28522 (N_28522,N_28342,N_28457);
nand U28523 (N_28523,N_28050,N_28200);
and U28524 (N_28524,N_28272,N_28350);
xor U28525 (N_28525,N_28172,N_28124);
nand U28526 (N_28526,N_28294,N_28151);
nor U28527 (N_28527,N_28009,N_28244);
or U28528 (N_28528,N_28379,N_28229);
or U28529 (N_28529,N_28005,N_28281);
nand U28530 (N_28530,N_28304,N_28283);
nor U28531 (N_28531,N_28038,N_28105);
nor U28532 (N_28532,N_28353,N_28218);
xor U28533 (N_28533,N_28288,N_28102);
and U28534 (N_28534,N_28339,N_28003);
or U28535 (N_28535,N_28321,N_28120);
nor U28536 (N_28536,N_28381,N_28421);
and U28537 (N_28537,N_28058,N_28332);
nor U28538 (N_28538,N_28008,N_28045);
xnor U28539 (N_28539,N_28356,N_28193);
nor U28540 (N_28540,N_28245,N_28352);
and U28541 (N_28541,N_28372,N_28338);
xnor U28542 (N_28542,N_28260,N_28111);
xor U28543 (N_28543,N_28441,N_28154);
xor U28544 (N_28544,N_28052,N_28483);
nand U28545 (N_28545,N_28484,N_28376);
nand U28546 (N_28546,N_28258,N_28046);
and U28547 (N_28547,N_28246,N_28217);
and U28548 (N_28548,N_28065,N_28159);
nor U28549 (N_28549,N_28398,N_28413);
or U28550 (N_28550,N_28150,N_28002);
nand U28551 (N_28551,N_28036,N_28481);
nor U28552 (N_28552,N_28165,N_28301);
nand U28553 (N_28553,N_28175,N_28148);
xnor U28554 (N_28554,N_28470,N_28486);
and U28555 (N_28555,N_28001,N_28435);
nor U28556 (N_28556,N_28396,N_28477);
and U28557 (N_28557,N_28267,N_28417);
nor U28558 (N_28558,N_28357,N_28029);
or U28559 (N_28559,N_28326,N_28063);
nor U28560 (N_28560,N_28375,N_28078);
or U28561 (N_28561,N_28087,N_28047);
or U28562 (N_28562,N_28264,N_28130);
or U28563 (N_28563,N_28182,N_28027);
xnor U28564 (N_28564,N_28026,N_28433);
xor U28565 (N_28565,N_28174,N_28257);
nand U28566 (N_28566,N_28259,N_28187);
nor U28567 (N_28567,N_28115,N_28176);
nand U28568 (N_28568,N_28416,N_28425);
and U28569 (N_28569,N_28117,N_28318);
nand U28570 (N_28570,N_28034,N_28266);
xnor U28571 (N_28571,N_28242,N_28162);
nand U28572 (N_28572,N_28292,N_28191);
or U28573 (N_28573,N_28168,N_28344);
or U28574 (N_28574,N_28449,N_28493);
and U28575 (N_28575,N_28018,N_28307);
xnor U28576 (N_28576,N_28138,N_28192);
nand U28577 (N_28577,N_28451,N_28313);
nand U28578 (N_28578,N_28430,N_28426);
or U28579 (N_28579,N_28136,N_28382);
nor U28580 (N_28580,N_28306,N_28055);
nand U28581 (N_28581,N_28360,N_28209);
nand U28582 (N_28582,N_28262,N_28494);
xor U28583 (N_28583,N_28400,N_28358);
nand U28584 (N_28584,N_28445,N_28465);
nor U28585 (N_28585,N_28143,N_28173);
and U28586 (N_28586,N_28189,N_28354);
nor U28587 (N_28587,N_28452,N_28127);
xnor U28588 (N_28588,N_28364,N_28412);
or U28589 (N_28589,N_28407,N_28196);
nand U28590 (N_28590,N_28028,N_28016);
nor U28591 (N_28591,N_28408,N_28346);
nor U28592 (N_28592,N_28496,N_28482);
xnor U28593 (N_28593,N_28324,N_28051);
or U28594 (N_28594,N_28167,N_28222);
nor U28595 (N_28595,N_28129,N_28438);
nand U28596 (N_28596,N_28156,N_28032);
nor U28597 (N_28597,N_28340,N_28456);
or U28598 (N_28598,N_28395,N_28023);
xnor U28599 (N_28599,N_28385,N_28128);
and U28600 (N_28600,N_28462,N_28060);
nor U28601 (N_28601,N_28049,N_28041);
or U28602 (N_28602,N_28231,N_28472);
xor U28603 (N_28603,N_28255,N_28077);
nand U28604 (N_28604,N_28071,N_28309);
and U28605 (N_28605,N_28424,N_28093);
nand U28606 (N_28606,N_28363,N_28180);
xnor U28607 (N_28607,N_28469,N_28160);
and U28608 (N_28608,N_28007,N_28139);
nor U28609 (N_28609,N_28302,N_28021);
nand U28610 (N_28610,N_28341,N_28223);
and U28611 (N_28611,N_28335,N_28277);
nor U28612 (N_28612,N_28019,N_28238);
and U28613 (N_28613,N_28022,N_28066);
xnor U28614 (N_28614,N_28183,N_28391);
and U28615 (N_28615,N_28237,N_28474);
nand U28616 (N_28616,N_28476,N_28099);
nor U28617 (N_28617,N_28351,N_28025);
xnor U28618 (N_28618,N_28250,N_28184);
nand U28619 (N_28619,N_28186,N_28000);
or U28620 (N_28620,N_28132,N_28431);
nor U28621 (N_28621,N_28056,N_28253);
or U28622 (N_28622,N_28295,N_28488);
nor U28623 (N_28623,N_28082,N_28075);
nand U28624 (N_28624,N_28163,N_28397);
nand U28625 (N_28625,N_28327,N_28444);
nor U28626 (N_28626,N_28399,N_28308);
nor U28627 (N_28627,N_28463,N_28155);
xnor U28628 (N_28628,N_28299,N_28211);
nor U28629 (N_28629,N_28454,N_28241);
or U28630 (N_28630,N_28461,N_28121);
nor U28631 (N_28631,N_28270,N_28053);
or U28632 (N_28632,N_28144,N_28490);
and U28633 (N_28633,N_28414,N_28406);
nor U28634 (N_28634,N_28458,N_28492);
and U28635 (N_28635,N_28337,N_28453);
and U28636 (N_28636,N_28142,N_28103);
nor U28637 (N_28637,N_28213,N_28020);
xnor U28638 (N_28638,N_28405,N_28202);
xnor U28639 (N_28639,N_28234,N_28439);
nor U28640 (N_28640,N_28328,N_28048);
nor U28641 (N_28641,N_28322,N_28164);
xor U28642 (N_28642,N_28073,N_28147);
nand U28643 (N_28643,N_28215,N_28355);
or U28644 (N_28644,N_28015,N_28320);
xor U28645 (N_28645,N_28325,N_28478);
nand U28646 (N_28646,N_28479,N_28276);
nand U28647 (N_28647,N_28409,N_28374);
nand U28648 (N_28648,N_28037,N_28498);
nor U28649 (N_28649,N_28370,N_28466);
nor U28650 (N_28650,N_28499,N_28081);
or U28651 (N_28651,N_28195,N_28141);
xnor U28652 (N_28652,N_28403,N_28094);
and U28653 (N_28653,N_28419,N_28236);
and U28654 (N_28654,N_28083,N_28442);
nor U28655 (N_28655,N_28248,N_28113);
or U28656 (N_28656,N_28158,N_28371);
and U28657 (N_28657,N_28384,N_28104);
nand U28658 (N_28658,N_28401,N_28092);
nand U28659 (N_28659,N_28079,N_28064);
nor U28660 (N_28660,N_28432,N_28135);
or U28661 (N_28661,N_28459,N_28254);
nor U28662 (N_28662,N_28411,N_28086);
nand U28663 (N_28663,N_28031,N_28315);
or U28664 (N_28664,N_28275,N_28054);
nand U28665 (N_28665,N_28091,N_28227);
nand U28666 (N_28666,N_28388,N_28263);
nand U28667 (N_28667,N_28467,N_28443);
or U28668 (N_28668,N_28284,N_28181);
nand U28669 (N_28669,N_28285,N_28373);
nand U28670 (N_28670,N_28291,N_28210);
nor U28671 (N_28671,N_28252,N_28273);
xor U28672 (N_28672,N_28293,N_28235);
and U28673 (N_28673,N_28024,N_28226);
nor U28674 (N_28674,N_28214,N_28423);
and U28675 (N_28675,N_28402,N_28289);
or U28676 (N_28676,N_28230,N_28393);
nor U28677 (N_28677,N_28146,N_28404);
nand U28678 (N_28678,N_28219,N_28035);
or U28679 (N_28679,N_28239,N_28311);
xnor U28680 (N_28680,N_28207,N_28336);
or U28681 (N_28681,N_28312,N_28446);
nand U28682 (N_28682,N_28437,N_28464);
xnor U28683 (N_28683,N_28487,N_28410);
nand U28684 (N_28684,N_28261,N_28434);
xnor U28685 (N_28685,N_28179,N_28185);
xnor U28686 (N_28686,N_28345,N_28491);
nand U28687 (N_28687,N_28190,N_28140);
and U28688 (N_28688,N_28169,N_28208);
nor U28689 (N_28689,N_28329,N_28122);
nand U28690 (N_28690,N_28387,N_28012);
nor U28691 (N_28691,N_28367,N_28224);
nor U28692 (N_28692,N_28468,N_28095);
nor U28693 (N_28693,N_28366,N_28380);
and U28694 (N_28694,N_28194,N_28177);
xor U28695 (N_28695,N_28039,N_28489);
and U28696 (N_28696,N_28427,N_28149);
xor U28697 (N_28697,N_28153,N_28447);
nand U28698 (N_28698,N_28377,N_28316);
xnor U28699 (N_28699,N_28203,N_28170);
or U28700 (N_28700,N_28290,N_28112);
nor U28701 (N_28701,N_28271,N_28330);
nor U28702 (N_28702,N_28084,N_28450);
nand U28703 (N_28703,N_28188,N_28247);
or U28704 (N_28704,N_28347,N_28300);
nor U28705 (N_28705,N_28033,N_28204);
xnor U28706 (N_28706,N_28298,N_28249);
nand U28707 (N_28707,N_28473,N_28333);
or U28708 (N_28708,N_28303,N_28296);
and U28709 (N_28709,N_28216,N_28317);
xor U28710 (N_28710,N_28042,N_28119);
nand U28711 (N_28711,N_28243,N_28485);
nor U28712 (N_28712,N_28030,N_28011);
and U28713 (N_28713,N_28343,N_28133);
xor U28714 (N_28714,N_28268,N_28278);
nor U28715 (N_28715,N_28436,N_28383);
nor U28716 (N_28716,N_28101,N_28471);
nor U28717 (N_28717,N_28134,N_28220);
nand U28718 (N_28718,N_28096,N_28090);
nor U28719 (N_28719,N_28349,N_28107);
or U28720 (N_28720,N_28098,N_28334);
or U28721 (N_28721,N_28221,N_28072);
xnor U28722 (N_28722,N_28206,N_28100);
and U28723 (N_28723,N_28069,N_28013);
and U28724 (N_28724,N_28455,N_28286);
xor U28725 (N_28725,N_28362,N_28361);
xor U28726 (N_28726,N_28240,N_28043);
xor U28727 (N_28727,N_28205,N_28420);
xnor U28728 (N_28728,N_28067,N_28394);
nand U28729 (N_28729,N_28197,N_28232);
nor U28730 (N_28730,N_28369,N_28123);
nor U28731 (N_28731,N_28460,N_28331);
xor U28732 (N_28732,N_28418,N_28114);
and U28733 (N_28733,N_28287,N_28152);
or U28734 (N_28734,N_28080,N_28085);
and U28735 (N_28735,N_28319,N_28280);
nand U28736 (N_28736,N_28274,N_28076);
or U28737 (N_28737,N_28057,N_28392);
and U28738 (N_28738,N_28495,N_28014);
or U28739 (N_28739,N_28390,N_28126);
xor U28740 (N_28740,N_28228,N_28314);
nand U28741 (N_28741,N_28116,N_28279);
nor U28742 (N_28742,N_28386,N_28282);
or U28743 (N_28743,N_28061,N_28251);
or U28744 (N_28744,N_28389,N_28480);
nor U28745 (N_28745,N_28497,N_28097);
nand U28746 (N_28746,N_28109,N_28368);
xnor U28747 (N_28747,N_28157,N_28198);
nand U28748 (N_28748,N_28448,N_28145);
nor U28749 (N_28749,N_28475,N_28074);
xnor U28750 (N_28750,N_28096,N_28328);
xor U28751 (N_28751,N_28384,N_28416);
or U28752 (N_28752,N_28287,N_28289);
nand U28753 (N_28753,N_28124,N_28431);
and U28754 (N_28754,N_28323,N_28257);
nor U28755 (N_28755,N_28050,N_28272);
xor U28756 (N_28756,N_28133,N_28197);
xnor U28757 (N_28757,N_28342,N_28361);
and U28758 (N_28758,N_28157,N_28032);
and U28759 (N_28759,N_28175,N_28072);
nand U28760 (N_28760,N_28443,N_28202);
nor U28761 (N_28761,N_28222,N_28344);
and U28762 (N_28762,N_28211,N_28445);
nand U28763 (N_28763,N_28298,N_28328);
or U28764 (N_28764,N_28191,N_28443);
nor U28765 (N_28765,N_28280,N_28359);
nor U28766 (N_28766,N_28012,N_28112);
xor U28767 (N_28767,N_28030,N_28450);
nor U28768 (N_28768,N_28465,N_28246);
and U28769 (N_28769,N_28042,N_28305);
and U28770 (N_28770,N_28255,N_28384);
nand U28771 (N_28771,N_28061,N_28351);
xor U28772 (N_28772,N_28459,N_28484);
and U28773 (N_28773,N_28399,N_28189);
or U28774 (N_28774,N_28199,N_28248);
nand U28775 (N_28775,N_28166,N_28197);
or U28776 (N_28776,N_28242,N_28020);
nand U28777 (N_28777,N_28221,N_28377);
or U28778 (N_28778,N_28407,N_28355);
nor U28779 (N_28779,N_28096,N_28067);
nand U28780 (N_28780,N_28310,N_28380);
and U28781 (N_28781,N_28277,N_28226);
nand U28782 (N_28782,N_28238,N_28476);
nor U28783 (N_28783,N_28380,N_28354);
nand U28784 (N_28784,N_28201,N_28476);
nand U28785 (N_28785,N_28183,N_28178);
xnor U28786 (N_28786,N_28189,N_28036);
or U28787 (N_28787,N_28285,N_28396);
nor U28788 (N_28788,N_28397,N_28297);
xor U28789 (N_28789,N_28491,N_28292);
xnor U28790 (N_28790,N_28483,N_28013);
and U28791 (N_28791,N_28243,N_28036);
and U28792 (N_28792,N_28040,N_28004);
nor U28793 (N_28793,N_28232,N_28411);
xnor U28794 (N_28794,N_28149,N_28412);
and U28795 (N_28795,N_28263,N_28236);
nand U28796 (N_28796,N_28380,N_28097);
and U28797 (N_28797,N_28035,N_28436);
and U28798 (N_28798,N_28298,N_28498);
and U28799 (N_28799,N_28159,N_28498);
or U28800 (N_28800,N_28140,N_28275);
nor U28801 (N_28801,N_28272,N_28478);
xor U28802 (N_28802,N_28286,N_28190);
and U28803 (N_28803,N_28307,N_28434);
or U28804 (N_28804,N_28369,N_28466);
or U28805 (N_28805,N_28487,N_28351);
or U28806 (N_28806,N_28361,N_28488);
or U28807 (N_28807,N_28292,N_28092);
and U28808 (N_28808,N_28438,N_28268);
nor U28809 (N_28809,N_28147,N_28472);
xnor U28810 (N_28810,N_28174,N_28222);
or U28811 (N_28811,N_28215,N_28200);
and U28812 (N_28812,N_28477,N_28079);
nor U28813 (N_28813,N_28093,N_28067);
nor U28814 (N_28814,N_28429,N_28444);
or U28815 (N_28815,N_28449,N_28463);
nor U28816 (N_28816,N_28129,N_28009);
nor U28817 (N_28817,N_28045,N_28363);
nor U28818 (N_28818,N_28228,N_28268);
and U28819 (N_28819,N_28140,N_28037);
xor U28820 (N_28820,N_28365,N_28115);
and U28821 (N_28821,N_28489,N_28367);
nand U28822 (N_28822,N_28425,N_28164);
or U28823 (N_28823,N_28220,N_28444);
nor U28824 (N_28824,N_28211,N_28318);
or U28825 (N_28825,N_28129,N_28198);
nor U28826 (N_28826,N_28285,N_28062);
nand U28827 (N_28827,N_28279,N_28113);
or U28828 (N_28828,N_28007,N_28118);
xnor U28829 (N_28829,N_28453,N_28496);
nand U28830 (N_28830,N_28055,N_28222);
and U28831 (N_28831,N_28417,N_28344);
xnor U28832 (N_28832,N_28087,N_28487);
nand U28833 (N_28833,N_28479,N_28487);
xnor U28834 (N_28834,N_28263,N_28489);
xnor U28835 (N_28835,N_28225,N_28152);
nand U28836 (N_28836,N_28311,N_28351);
nand U28837 (N_28837,N_28058,N_28462);
xnor U28838 (N_28838,N_28285,N_28237);
nand U28839 (N_28839,N_28133,N_28065);
nand U28840 (N_28840,N_28341,N_28167);
and U28841 (N_28841,N_28250,N_28127);
xor U28842 (N_28842,N_28423,N_28314);
or U28843 (N_28843,N_28455,N_28053);
nand U28844 (N_28844,N_28446,N_28428);
and U28845 (N_28845,N_28108,N_28109);
and U28846 (N_28846,N_28381,N_28274);
and U28847 (N_28847,N_28245,N_28196);
or U28848 (N_28848,N_28316,N_28374);
xnor U28849 (N_28849,N_28208,N_28344);
xnor U28850 (N_28850,N_28150,N_28072);
and U28851 (N_28851,N_28476,N_28265);
nand U28852 (N_28852,N_28316,N_28011);
xnor U28853 (N_28853,N_28388,N_28062);
xor U28854 (N_28854,N_28354,N_28114);
nor U28855 (N_28855,N_28018,N_28407);
xnor U28856 (N_28856,N_28430,N_28459);
and U28857 (N_28857,N_28253,N_28152);
and U28858 (N_28858,N_28060,N_28138);
or U28859 (N_28859,N_28178,N_28116);
xor U28860 (N_28860,N_28490,N_28306);
xnor U28861 (N_28861,N_28499,N_28305);
nand U28862 (N_28862,N_28466,N_28299);
or U28863 (N_28863,N_28141,N_28275);
xnor U28864 (N_28864,N_28120,N_28140);
nor U28865 (N_28865,N_28374,N_28216);
xor U28866 (N_28866,N_28121,N_28232);
xnor U28867 (N_28867,N_28142,N_28171);
and U28868 (N_28868,N_28307,N_28031);
nand U28869 (N_28869,N_28182,N_28458);
nor U28870 (N_28870,N_28234,N_28239);
nor U28871 (N_28871,N_28347,N_28120);
or U28872 (N_28872,N_28360,N_28362);
nand U28873 (N_28873,N_28074,N_28432);
xnor U28874 (N_28874,N_28341,N_28102);
and U28875 (N_28875,N_28136,N_28230);
nor U28876 (N_28876,N_28100,N_28074);
or U28877 (N_28877,N_28008,N_28369);
or U28878 (N_28878,N_28215,N_28167);
or U28879 (N_28879,N_28465,N_28481);
and U28880 (N_28880,N_28369,N_28252);
or U28881 (N_28881,N_28129,N_28364);
nor U28882 (N_28882,N_28397,N_28213);
or U28883 (N_28883,N_28333,N_28355);
xnor U28884 (N_28884,N_28443,N_28001);
and U28885 (N_28885,N_28426,N_28027);
nor U28886 (N_28886,N_28122,N_28388);
nor U28887 (N_28887,N_28231,N_28350);
nand U28888 (N_28888,N_28162,N_28152);
or U28889 (N_28889,N_28258,N_28067);
xor U28890 (N_28890,N_28213,N_28267);
nor U28891 (N_28891,N_28460,N_28442);
nor U28892 (N_28892,N_28147,N_28141);
or U28893 (N_28893,N_28498,N_28153);
xnor U28894 (N_28894,N_28466,N_28475);
xnor U28895 (N_28895,N_28430,N_28193);
xnor U28896 (N_28896,N_28238,N_28084);
and U28897 (N_28897,N_28141,N_28437);
and U28898 (N_28898,N_28274,N_28355);
xnor U28899 (N_28899,N_28103,N_28088);
xnor U28900 (N_28900,N_28327,N_28023);
or U28901 (N_28901,N_28116,N_28471);
nor U28902 (N_28902,N_28458,N_28455);
nand U28903 (N_28903,N_28493,N_28090);
or U28904 (N_28904,N_28267,N_28317);
xor U28905 (N_28905,N_28027,N_28454);
nand U28906 (N_28906,N_28321,N_28267);
nand U28907 (N_28907,N_28217,N_28059);
nand U28908 (N_28908,N_28450,N_28040);
nor U28909 (N_28909,N_28397,N_28338);
xnor U28910 (N_28910,N_28181,N_28076);
nand U28911 (N_28911,N_28468,N_28190);
nand U28912 (N_28912,N_28255,N_28139);
or U28913 (N_28913,N_28274,N_28074);
xor U28914 (N_28914,N_28016,N_28088);
and U28915 (N_28915,N_28066,N_28297);
and U28916 (N_28916,N_28103,N_28399);
and U28917 (N_28917,N_28061,N_28486);
and U28918 (N_28918,N_28052,N_28340);
and U28919 (N_28919,N_28383,N_28193);
and U28920 (N_28920,N_28431,N_28120);
and U28921 (N_28921,N_28481,N_28046);
nand U28922 (N_28922,N_28145,N_28065);
and U28923 (N_28923,N_28261,N_28013);
nor U28924 (N_28924,N_28289,N_28327);
xor U28925 (N_28925,N_28082,N_28436);
xnor U28926 (N_28926,N_28013,N_28018);
nor U28927 (N_28927,N_28090,N_28022);
nand U28928 (N_28928,N_28147,N_28477);
nor U28929 (N_28929,N_28121,N_28332);
or U28930 (N_28930,N_28475,N_28418);
or U28931 (N_28931,N_28491,N_28221);
xnor U28932 (N_28932,N_28351,N_28359);
nor U28933 (N_28933,N_28343,N_28235);
and U28934 (N_28934,N_28123,N_28021);
xor U28935 (N_28935,N_28362,N_28299);
xnor U28936 (N_28936,N_28050,N_28423);
xnor U28937 (N_28937,N_28440,N_28485);
nand U28938 (N_28938,N_28120,N_28044);
nand U28939 (N_28939,N_28234,N_28247);
nor U28940 (N_28940,N_28373,N_28341);
or U28941 (N_28941,N_28034,N_28028);
or U28942 (N_28942,N_28067,N_28408);
xnor U28943 (N_28943,N_28330,N_28006);
nand U28944 (N_28944,N_28206,N_28196);
nand U28945 (N_28945,N_28101,N_28474);
and U28946 (N_28946,N_28051,N_28372);
or U28947 (N_28947,N_28348,N_28451);
xor U28948 (N_28948,N_28430,N_28375);
and U28949 (N_28949,N_28447,N_28384);
nor U28950 (N_28950,N_28358,N_28102);
xnor U28951 (N_28951,N_28294,N_28324);
nand U28952 (N_28952,N_28177,N_28415);
or U28953 (N_28953,N_28032,N_28271);
nor U28954 (N_28954,N_28370,N_28285);
xor U28955 (N_28955,N_28085,N_28172);
and U28956 (N_28956,N_28041,N_28499);
or U28957 (N_28957,N_28228,N_28011);
xor U28958 (N_28958,N_28262,N_28401);
and U28959 (N_28959,N_28350,N_28095);
and U28960 (N_28960,N_28387,N_28313);
nand U28961 (N_28961,N_28124,N_28377);
nand U28962 (N_28962,N_28289,N_28308);
xnor U28963 (N_28963,N_28361,N_28487);
nand U28964 (N_28964,N_28423,N_28093);
nand U28965 (N_28965,N_28251,N_28036);
nor U28966 (N_28966,N_28397,N_28466);
or U28967 (N_28967,N_28300,N_28186);
or U28968 (N_28968,N_28264,N_28138);
nor U28969 (N_28969,N_28247,N_28289);
nor U28970 (N_28970,N_28318,N_28018);
xnor U28971 (N_28971,N_28362,N_28279);
nand U28972 (N_28972,N_28153,N_28228);
nand U28973 (N_28973,N_28379,N_28145);
nand U28974 (N_28974,N_28018,N_28163);
and U28975 (N_28975,N_28088,N_28004);
nand U28976 (N_28976,N_28441,N_28075);
and U28977 (N_28977,N_28412,N_28370);
and U28978 (N_28978,N_28226,N_28122);
nand U28979 (N_28979,N_28240,N_28378);
nand U28980 (N_28980,N_28322,N_28109);
or U28981 (N_28981,N_28094,N_28008);
xnor U28982 (N_28982,N_28241,N_28034);
nand U28983 (N_28983,N_28348,N_28092);
xor U28984 (N_28984,N_28121,N_28236);
nand U28985 (N_28985,N_28386,N_28432);
or U28986 (N_28986,N_28014,N_28102);
nand U28987 (N_28987,N_28305,N_28004);
nor U28988 (N_28988,N_28151,N_28097);
and U28989 (N_28989,N_28363,N_28177);
and U28990 (N_28990,N_28410,N_28343);
nor U28991 (N_28991,N_28182,N_28126);
nor U28992 (N_28992,N_28204,N_28381);
xor U28993 (N_28993,N_28166,N_28489);
xnor U28994 (N_28994,N_28431,N_28121);
xor U28995 (N_28995,N_28050,N_28472);
xnor U28996 (N_28996,N_28273,N_28404);
and U28997 (N_28997,N_28357,N_28286);
nand U28998 (N_28998,N_28174,N_28242);
nor U28999 (N_28999,N_28054,N_28274);
nand U29000 (N_29000,N_28536,N_28846);
and U29001 (N_29001,N_28887,N_28654);
and U29002 (N_29002,N_28738,N_28689);
nand U29003 (N_29003,N_28672,N_28911);
xnor U29004 (N_29004,N_28859,N_28816);
and U29005 (N_29005,N_28532,N_28899);
nand U29006 (N_29006,N_28783,N_28962);
nor U29007 (N_29007,N_28628,N_28798);
or U29008 (N_29008,N_28529,N_28773);
and U29009 (N_29009,N_28603,N_28568);
or U29010 (N_29010,N_28676,N_28582);
nand U29011 (N_29011,N_28758,N_28598);
or U29012 (N_29012,N_28700,N_28606);
and U29013 (N_29013,N_28727,N_28750);
and U29014 (N_29014,N_28819,N_28631);
nand U29015 (N_29015,N_28514,N_28537);
nor U29016 (N_29016,N_28611,N_28935);
and U29017 (N_29017,N_28993,N_28730);
nor U29018 (N_29018,N_28748,N_28665);
nor U29019 (N_29019,N_28726,N_28985);
nand U29020 (N_29020,N_28833,N_28566);
nand U29021 (N_29021,N_28921,N_28601);
or U29022 (N_29022,N_28704,N_28740);
and U29023 (N_29023,N_28602,N_28761);
nand U29024 (N_29024,N_28504,N_28973);
and U29025 (N_29025,N_28677,N_28904);
nand U29026 (N_29026,N_28570,N_28967);
nand U29027 (N_29027,N_28872,N_28511);
and U29028 (N_29028,N_28731,N_28818);
xor U29029 (N_29029,N_28564,N_28707);
nand U29030 (N_29030,N_28558,N_28926);
nor U29031 (N_29031,N_28950,N_28618);
xor U29032 (N_29032,N_28728,N_28625);
and U29033 (N_29033,N_28988,N_28938);
and U29034 (N_29034,N_28500,N_28678);
nand U29035 (N_29035,N_28538,N_28579);
nand U29036 (N_29036,N_28814,N_28745);
nand U29037 (N_29037,N_28876,N_28711);
nor U29038 (N_29038,N_28743,N_28643);
and U29039 (N_29039,N_28903,N_28615);
xnor U29040 (N_29040,N_28556,N_28512);
nand U29041 (N_29041,N_28778,N_28797);
or U29042 (N_29042,N_28834,N_28994);
nor U29043 (N_29043,N_28652,N_28679);
or U29044 (N_29044,N_28807,N_28775);
nand U29045 (N_29045,N_28546,N_28593);
or U29046 (N_29046,N_28729,N_28870);
and U29047 (N_29047,N_28976,N_28765);
or U29048 (N_29048,N_28604,N_28645);
and U29049 (N_29049,N_28609,N_28680);
nand U29050 (N_29050,N_28896,N_28649);
nor U29051 (N_29051,N_28684,N_28561);
xnor U29052 (N_29052,N_28721,N_28524);
or U29053 (N_29053,N_28811,N_28760);
nor U29054 (N_29054,N_28864,N_28724);
nor U29055 (N_29055,N_28660,N_28917);
nand U29056 (N_29056,N_28785,N_28505);
or U29057 (N_29057,N_28638,N_28966);
and U29058 (N_29058,N_28523,N_28709);
nand U29059 (N_29059,N_28632,N_28856);
nor U29060 (N_29060,N_28545,N_28795);
and U29061 (N_29061,N_28629,N_28883);
and U29062 (N_29062,N_28619,N_28626);
and U29063 (N_29063,N_28706,N_28831);
or U29064 (N_29064,N_28534,N_28793);
nand U29065 (N_29065,N_28884,N_28847);
xnor U29066 (N_29066,N_28995,N_28822);
nand U29067 (N_29067,N_28623,N_28923);
and U29068 (N_29068,N_28855,N_28553);
or U29069 (N_29069,N_28817,N_28624);
and U29070 (N_29070,N_28969,N_28812);
nor U29071 (N_29071,N_28640,N_28989);
and U29072 (N_29072,N_28791,N_28688);
or U29073 (N_29073,N_28563,N_28910);
nor U29074 (N_29074,N_28548,N_28501);
or U29075 (N_29075,N_28838,N_28908);
or U29076 (N_29076,N_28972,N_28755);
nor U29077 (N_29077,N_28861,N_28725);
nand U29078 (N_29078,N_28779,N_28737);
nand U29079 (N_29079,N_28590,N_28983);
and U29080 (N_29080,N_28658,N_28659);
nand U29081 (N_29081,N_28559,N_28999);
xnor U29082 (N_29082,N_28752,N_28915);
nor U29083 (N_29083,N_28844,N_28974);
nand U29084 (N_29084,N_28769,N_28881);
nand U29085 (N_29085,N_28698,N_28510);
xor U29086 (N_29086,N_28544,N_28875);
nor U29087 (N_29087,N_28820,N_28613);
or U29088 (N_29088,N_28521,N_28550);
nor U29089 (N_29089,N_28565,N_28719);
and U29090 (N_29090,N_28956,N_28502);
nand U29091 (N_29091,N_28703,N_28918);
nand U29092 (N_29092,N_28766,N_28979);
nor U29093 (N_29093,N_28694,N_28539);
and U29094 (N_29094,N_28897,N_28541);
xor U29095 (N_29095,N_28685,N_28647);
or U29096 (N_29096,N_28757,N_28549);
and U29097 (N_29097,N_28525,N_28715);
nand U29098 (N_29098,N_28936,N_28998);
nand U29099 (N_29099,N_28930,N_28691);
xor U29100 (N_29100,N_28746,N_28906);
nand U29101 (N_29101,N_28503,N_28800);
nor U29102 (N_29102,N_28522,N_28587);
xor U29103 (N_29103,N_28866,N_28806);
nand U29104 (N_29104,N_28599,N_28937);
nor U29105 (N_29105,N_28850,N_28986);
xnor U29106 (N_29106,N_28673,N_28944);
nand U29107 (N_29107,N_28576,N_28633);
and U29108 (N_29108,N_28916,N_28661);
xor U29109 (N_29109,N_28637,N_28718);
or U29110 (N_29110,N_28622,N_28580);
nand U29111 (N_29111,N_28687,N_28535);
or U29112 (N_29112,N_28581,N_28630);
nand U29113 (N_29113,N_28507,N_28843);
xnor U29114 (N_29114,N_28781,N_28853);
xnor U29115 (N_29115,N_28696,N_28981);
and U29116 (N_29116,N_28825,N_28509);
or U29117 (N_29117,N_28794,N_28931);
or U29118 (N_29118,N_28751,N_28686);
nand U29119 (N_29119,N_28965,N_28655);
or U29120 (N_29120,N_28513,N_28939);
nand U29121 (N_29121,N_28827,N_28701);
and U29122 (N_29122,N_28786,N_28877);
xor U29123 (N_29123,N_28805,N_28826);
or U29124 (N_29124,N_28552,N_28670);
nor U29125 (N_29125,N_28690,N_28878);
or U29126 (N_29126,N_28946,N_28753);
nand U29127 (N_29127,N_28955,N_28865);
and U29128 (N_29128,N_28650,N_28591);
nor U29129 (N_29129,N_28506,N_28790);
nand U29130 (N_29130,N_28767,N_28617);
xor U29131 (N_29131,N_28934,N_28895);
xor U29132 (N_29132,N_28953,N_28739);
nand U29133 (N_29133,N_28759,N_28968);
and U29134 (N_29134,N_28971,N_28662);
nand U29135 (N_29135,N_28891,N_28763);
xnor U29136 (N_29136,N_28666,N_28517);
nand U29137 (N_29137,N_28657,N_28848);
nand U29138 (N_29138,N_28792,N_28959);
nor U29139 (N_29139,N_28880,N_28720);
nand U29140 (N_29140,N_28656,N_28585);
xor U29141 (N_29141,N_28823,N_28924);
and U29142 (N_29142,N_28671,N_28799);
nand U29143 (N_29143,N_28642,N_28960);
or U29144 (N_29144,N_28929,N_28997);
nand U29145 (N_29145,N_28868,N_28577);
or U29146 (N_29146,N_28892,N_28970);
and U29147 (N_29147,N_28941,N_28902);
or U29148 (N_29148,N_28648,N_28554);
nand U29149 (N_29149,N_28942,N_28894);
nor U29150 (N_29150,N_28675,N_28832);
and U29151 (N_29151,N_28575,N_28519);
or U29152 (N_29152,N_28947,N_28889);
xor U29153 (N_29153,N_28515,N_28742);
nand U29154 (N_29154,N_28933,N_28734);
xor U29155 (N_29155,N_28695,N_28867);
nand U29156 (N_29156,N_28749,N_28957);
nor U29157 (N_29157,N_28574,N_28837);
and U29158 (N_29158,N_28569,N_28849);
and U29159 (N_29159,N_28716,N_28951);
nor U29160 (N_29160,N_28905,N_28900);
nand U29161 (N_29161,N_28871,N_28789);
xor U29162 (N_29162,N_28780,N_28772);
or U29163 (N_29163,N_28835,N_28879);
xnor U29164 (N_29164,N_28830,N_28768);
nand U29165 (N_29165,N_28901,N_28705);
or U29166 (N_29166,N_28620,N_28952);
nor U29167 (N_29167,N_28914,N_28782);
nand U29168 (N_29168,N_28940,N_28990);
nand U29169 (N_29169,N_28717,N_28949);
or U29170 (N_29170,N_28592,N_28610);
and U29171 (N_29171,N_28641,N_28635);
nor U29172 (N_29172,N_28646,N_28607);
xnor U29173 (N_29173,N_28943,N_28982);
and U29174 (N_29174,N_28810,N_28608);
xnor U29175 (N_29175,N_28653,N_28796);
or U29176 (N_29176,N_28714,N_28508);
nand U29177 (N_29177,N_28925,N_28595);
nor U29178 (N_29178,N_28913,N_28526);
nand U29179 (N_29179,N_28616,N_28770);
and U29180 (N_29180,N_28735,N_28804);
nor U29181 (N_29181,N_28784,N_28669);
nand U29182 (N_29182,N_28663,N_28862);
nand U29183 (N_29183,N_28588,N_28697);
and U29184 (N_29184,N_28928,N_28912);
nand U29185 (N_29185,N_28692,N_28774);
or U29186 (N_29186,N_28586,N_28845);
xnor U29187 (N_29187,N_28597,N_28828);
xnor U29188 (N_29188,N_28732,N_28922);
and U29189 (N_29189,N_28776,N_28991);
or U29190 (N_29190,N_28874,N_28614);
or U29191 (N_29191,N_28771,N_28762);
or U29192 (N_29192,N_28754,N_28621);
and U29193 (N_29193,N_28644,N_28898);
and U29194 (N_29194,N_28600,N_28664);
and U29195 (N_29195,N_28984,N_28975);
xnor U29196 (N_29196,N_28528,N_28747);
or U29197 (N_29197,N_28674,N_28699);
or U29198 (N_29198,N_28987,N_28605);
xnor U29199 (N_29199,N_28788,N_28869);
nand U29200 (N_29200,N_28516,N_28722);
xor U29201 (N_29201,N_28815,N_28557);
xnor U29202 (N_29202,N_28932,N_28945);
xor U29203 (N_29203,N_28713,N_28996);
nor U29204 (N_29204,N_28744,N_28840);
nand U29205 (N_29205,N_28992,N_28702);
xnor U29206 (N_29206,N_28839,N_28954);
xor U29207 (N_29207,N_28560,N_28741);
and U29208 (N_29208,N_28682,N_28777);
and U29209 (N_29209,N_28668,N_28683);
nor U29210 (N_29210,N_28961,N_28764);
nand U29211 (N_29211,N_28890,N_28723);
nor U29212 (N_29212,N_28882,N_28919);
and U29213 (N_29213,N_28578,N_28948);
or U29214 (N_29214,N_28873,N_28907);
nor U29215 (N_29215,N_28888,N_28543);
and U29216 (N_29216,N_28958,N_28808);
and U29217 (N_29217,N_28612,N_28567);
nor U29218 (N_29218,N_28885,N_28636);
and U29219 (N_29219,N_28571,N_28520);
nor U29220 (N_29220,N_28909,N_28710);
nand U29221 (N_29221,N_28634,N_28712);
xor U29222 (N_29222,N_28533,N_28803);
nand U29223 (N_29223,N_28572,N_28893);
or U29224 (N_29224,N_28540,N_28531);
nor U29225 (N_29225,N_28681,N_28736);
or U29226 (N_29226,N_28787,N_28756);
xnor U29227 (N_29227,N_28977,N_28978);
xor U29228 (N_29228,N_28927,N_28860);
and U29229 (N_29229,N_28821,N_28802);
xor U29230 (N_29230,N_28857,N_28963);
nor U29231 (N_29231,N_28858,N_28813);
nor U29232 (N_29232,N_28596,N_28627);
nand U29233 (N_29233,N_28801,N_28583);
nand U29234 (N_29234,N_28863,N_28542);
nand U29235 (N_29235,N_28573,N_28530);
nand U29236 (N_29236,N_28584,N_28562);
and U29237 (N_29237,N_28551,N_28667);
and U29238 (N_29238,N_28829,N_28733);
or U29239 (N_29239,N_28852,N_28809);
nand U29240 (N_29240,N_28886,N_28527);
or U29241 (N_29241,N_28708,N_28693);
nand U29242 (N_29242,N_28547,N_28594);
or U29243 (N_29243,N_28589,N_28518);
nor U29244 (N_29244,N_28836,N_28964);
xnor U29245 (N_29245,N_28854,N_28841);
nand U29246 (N_29246,N_28980,N_28651);
nand U29247 (N_29247,N_28824,N_28920);
nor U29248 (N_29248,N_28851,N_28639);
and U29249 (N_29249,N_28555,N_28842);
xor U29250 (N_29250,N_28615,N_28578);
or U29251 (N_29251,N_28643,N_28989);
and U29252 (N_29252,N_28536,N_28586);
nor U29253 (N_29253,N_28837,N_28789);
nor U29254 (N_29254,N_28975,N_28870);
and U29255 (N_29255,N_28565,N_28640);
and U29256 (N_29256,N_28570,N_28655);
xor U29257 (N_29257,N_28619,N_28525);
and U29258 (N_29258,N_28763,N_28997);
nor U29259 (N_29259,N_28804,N_28875);
xor U29260 (N_29260,N_28758,N_28947);
or U29261 (N_29261,N_28798,N_28684);
or U29262 (N_29262,N_28881,N_28571);
nor U29263 (N_29263,N_28799,N_28607);
or U29264 (N_29264,N_28538,N_28712);
nand U29265 (N_29265,N_28936,N_28658);
nor U29266 (N_29266,N_28554,N_28847);
nand U29267 (N_29267,N_28871,N_28540);
and U29268 (N_29268,N_28961,N_28598);
nor U29269 (N_29269,N_28764,N_28842);
or U29270 (N_29270,N_28809,N_28902);
xor U29271 (N_29271,N_28959,N_28870);
xnor U29272 (N_29272,N_28957,N_28919);
or U29273 (N_29273,N_28764,N_28537);
or U29274 (N_29274,N_28696,N_28649);
xor U29275 (N_29275,N_28913,N_28539);
nand U29276 (N_29276,N_28691,N_28995);
nor U29277 (N_29277,N_28714,N_28583);
or U29278 (N_29278,N_28915,N_28540);
xor U29279 (N_29279,N_28743,N_28974);
or U29280 (N_29280,N_28552,N_28739);
nor U29281 (N_29281,N_28551,N_28713);
and U29282 (N_29282,N_28944,N_28866);
xnor U29283 (N_29283,N_28947,N_28786);
nand U29284 (N_29284,N_28856,N_28816);
or U29285 (N_29285,N_28608,N_28553);
nand U29286 (N_29286,N_28588,N_28821);
nor U29287 (N_29287,N_28978,N_28926);
or U29288 (N_29288,N_28685,N_28642);
nand U29289 (N_29289,N_28721,N_28538);
nand U29290 (N_29290,N_28911,N_28622);
nor U29291 (N_29291,N_28541,N_28507);
and U29292 (N_29292,N_28541,N_28591);
xnor U29293 (N_29293,N_28941,N_28935);
nand U29294 (N_29294,N_28522,N_28753);
or U29295 (N_29295,N_28556,N_28675);
nor U29296 (N_29296,N_28728,N_28707);
and U29297 (N_29297,N_28593,N_28709);
nor U29298 (N_29298,N_28716,N_28585);
nand U29299 (N_29299,N_28575,N_28620);
and U29300 (N_29300,N_28740,N_28981);
nor U29301 (N_29301,N_28655,N_28526);
xnor U29302 (N_29302,N_28873,N_28944);
and U29303 (N_29303,N_28536,N_28693);
nor U29304 (N_29304,N_28925,N_28946);
and U29305 (N_29305,N_28670,N_28532);
nand U29306 (N_29306,N_28698,N_28585);
and U29307 (N_29307,N_28540,N_28984);
nor U29308 (N_29308,N_28892,N_28948);
and U29309 (N_29309,N_28869,N_28865);
xnor U29310 (N_29310,N_28625,N_28974);
nand U29311 (N_29311,N_28980,N_28818);
nor U29312 (N_29312,N_28556,N_28830);
xor U29313 (N_29313,N_28595,N_28957);
and U29314 (N_29314,N_28694,N_28824);
or U29315 (N_29315,N_28758,N_28826);
xnor U29316 (N_29316,N_28940,N_28922);
xor U29317 (N_29317,N_28553,N_28997);
nor U29318 (N_29318,N_28710,N_28539);
or U29319 (N_29319,N_28543,N_28739);
nand U29320 (N_29320,N_28657,N_28755);
or U29321 (N_29321,N_28972,N_28756);
xor U29322 (N_29322,N_28560,N_28959);
and U29323 (N_29323,N_28841,N_28780);
nor U29324 (N_29324,N_28580,N_28766);
xnor U29325 (N_29325,N_28888,N_28621);
or U29326 (N_29326,N_28599,N_28879);
xor U29327 (N_29327,N_28896,N_28786);
xnor U29328 (N_29328,N_28545,N_28891);
or U29329 (N_29329,N_28835,N_28659);
xor U29330 (N_29330,N_28976,N_28561);
nor U29331 (N_29331,N_28505,N_28720);
nor U29332 (N_29332,N_28614,N_28666);
nand U29333 (N_29333,N_28883,N_28966);
or U29334 (N_29334,N_28970,N_28859);
and U29335 (N_29335,N_28544,N_28988);
nor U29336 (N_29336,N_28844,N_28501);
nand U29337 (N_29337,N_28635,N_28758);
nor U29338 (N_29338,N_28707,N_28721);
nand U29339 (N_29339,N_28910,N_28614);
or U29340 (N_29340,N_28548,N_28985);
and U29341 (N_29341,N_28747,N_28787);
xor U29342 (N_29342,N_28833,N_28642);
nor U29343 (N_29343,N_28614,N_28683);
and U29344 (N_29344,N_28649,N_28984);
and U29345 (N_29345,N_28562,N_28941);
and U29346 (N_29346,N_28596,N_28663);
xor U29347 (N_29347,N_28811,N_28674);
and U29348 (N_29348,N_28843,N_28588);
and U29349 (N_29349,N_28604,N_28892);
and U29350 (N_29350,N_28996,N_28932);
nand U29351 (N_29351,N_28929,N_28773);
nand U29352 (N_29352,N_28892,N_28550);
nor U29353 (N_29353,N_28749,N_28602);
and U29354 (N_29354,N_28929,N_28697);
or U29355 (N_29355,N_28804,N_28525);
and U29356 (N_29356,N_28944,N_28738);
nand U29357 (N_29357,N_28998,N_28842);
nor U29358 (N_29358,N_28835,N_28523);
nand U29359 (N_29359,N_28524,N_28972);
nand U29360 (N_29360,N_28566,N_28606);
nor U29361 (N_29361,N_28960,N_28516);
or U29362 (N_29362,N_28750,N_28627);
nor U29363 (N_29363,N_28613,N_28651);
or U29364 (N_29364,N_28582,N_28736);
nor U29365 (N_29365,N_28506,N_28521);
nor U29366 (N_29366,N_28849,N_28555);
nor U29367 (N_29367,N_28811,N_28591);
nand U29368 (N_29368,N_28518,N_28955);
nand U29369 (N_29369,N_28735,N_28676);
and U29370 (N_29370,N_28801,N_28786);
or U29371 (N_29371,N_28891,N_28970);
xnor U29372 (N_29372,N_28891,N_28996);
or U29373 (N_29373,N_28908,N_28973);
nor U29374 (N_29374,N_28516,N_28680);
nor U29375 (N_29375,N_28566,N_28832);
nor U29376 (N_29376,N_28620,N_28684);
xor U29377 (N_29377,N_28667,N_28850);
xnor U29378 (N_29378,N_28581,N_28988);
nor U29379 (N_29379,N_28619,N_28526);
nand U29380 (N_29380,N_28801,N_28946);
nor U29381 (N_29381,N_28999,N_28847);
nand U29382 (N_29382,N_28806,N_28891);
nand U29383 (N_29383,N_28689,N_28691);
and U29384 (N_29384,N_28629,N_28931);
and U29385 (N_29385,N_28559,N_28513);
or U29386 (N_29386,N_28672,N_28664);
nand U29387 (N_29387,N_28651,N_28742);
or U29388 (N_29388,N_28637,N_28655);
and U29389 (N_29389,N_28845,N_28853);
nor U29390 (N_29390,N_28930,N_28662);
or U29391 (N_29391,N_28545,N_28667);
and U29392 (N_29392,N_28909,N_28508);
or U29393 (N_29393,N_28735,N_28890);
or U29394 (N_29394,N_28781,N_28898);
nand U29395 (N_29395,N_28904,N_28987);
nor U29396 (N_29396,N_28599,N_28541);
nand U29397 (N_29397,N_28699,N_28626);
and U29398 (N_29398,N_28538,N_28852);
or U29399 (N_29399,N_28985,N_28724);
xnor U29400 (N_29400,N_28862,N_28644);
and U29401 (N_29401,N_28631,N_28967);
nor U29402 (N_29402,N_28999,N_28504);
or U29403 (N_29403,N_28527,N_28721);
and U29404 (N_29404,N_28765,N_28829);
nand U29405 (N_29405,N_28772,N_28543);
or U29406 (N_29406,N_28744,N_28909);
xnor U29407 (N_29407,N_28731,N_28889);
xor U29408 (N_29408,N_28981,N_28903);
and U29409 (N_29409,N_28752,N_28908);
or U29410 (N_29410,N_28917,N_28830);
or U29411 (N_29411,N_28816,N_28642);
or U29412 (N_29412,N_28531,N_28808);
nand U29413 (N_29413,N_28886,N_28560);
nand U29414 (N_29414,N_28598,N_28564);
or U29415 (N_29415,N_28596,N_28801);
xnor U29416 (N_29416,N_28753,N_28921);
or U29417 (N_29417,N_28571,N_28674);
nor U29418 (N_29418,N_28642,N_28681);
nor U29419 (N_29419,N_28530,N_28880);
nor U29420 (N_29420,N_28765,N_28838);
and U29421 (N_29421,N_28771,N_28500);
or U29422 (N_29422,N_28805,N_28634);
nand U29423 (N_29423,N_28672,N_28620);
nor U29424 (N_29424,N_28735,N_28680);
xnor U29425 (N_29425,N_28743,N_28944);
nand U29426 (N_29426,N_28511,N_28664);
and U29427 (N_29427,N_28616,N_28840);
xor U29428 (N_29428,N_28783,N_28846);
and U29429 (N_29429,N_28500,N_28743);
xnor U29430 (N_29430,N_28665,N_28782);
xnor U29431 (N_29431,N_28728,N_28822);
and U29432 (N_29432,N_28868,N_28832);
nor U29433 (N_29433,N_28984,N_28769);
nand U29434 (N_29434,N_28661,N_28534);
or U29435 (N_29435,N_28585,N_28525);
nand U29436 (N_29436,N_28980,N_28875);
nor U29437 (N_29437,N_28523,N_28754);
or U29438 (N_29438,N_28622,N_28882);
or U29439 (N_29439,N_28740,N_28967);
or U29440 (N_29440,N_28829,N_28852);
and U29441 (N_29441,N_28578,N_28816);
nor U29442 (N_29442,N_28921,N_28534);
xor U29443 (N_29443,N_28776,N_28988);
and U29444 (N_29444,N_28567,N_28614);
nand U29445 (N_29445,N_28762,N_28661);
and U29446 (N_29446,N_28703,N_28904);
and U29447 (N_29447,N_28842,N_28800);
nor U29448 (N_29448,N_28863,N_28565);
or U29449 (N_29449,N_28838,N_28926);
nor U29450 (N_29450,N_28527,N_28702);
and U29451 (N_29451,N_28904,N_28505);
nor U29452 (N_29452,N_28672,N_28863);
xor U29453 (N_29453,N_28998,N_28879);
xor U29454 (N_29454,N_28912,N_28667);
xnor U29455 (N_29455,N_28625,N_28652);
nor U29456 (N_29456,N_28752,N_28843);
or U29457 (N_29457,N_28937,N_28701);
or U29458 (N_29458,N_28948,N_28634);
xor U29459 (N_29459,N_28640,N_28632);
nand U29460 (N_29460,N_28715,N_28955);
and U29461 (N_29461,N_28703,N_28568);
nor U29462 (N_29462,N_28704,N_28718);
nand U29463 (N_29463,N_28844,N_28629);
xor U29464 (N_29464,N_28659,N_28980);
nor U29465 (N_29465,N_28912,N_28954);
and U29466 (N_29466,N_28555,N_28509);
nand U29467 (N_29467,N_28544,N_28964);
nor U29468 (N_29468,N_28758,N_28642);
nor U29469 (N_29469,N_28629,N_28616);
xor U29470 (N_29470,N_28528,N_28720);
or U29471 (N_29471,N_28984,N_28829);
and U29472 (N_29472,N_28954,N_28945);
and U29473 (N_29473,N_28935,N_28948);
nand U29474 (N_29474,N_28551,N_28566);
nand U29475 (N_29475,N_28703,N_28716);
or U29476 (N_29476,N_28628,N_28960);
nand U29477 (N_29477,N_28955,N_28756);
nand U29478 (N_29478,N_28550,N_28744);
and U29479 (N_29479,N_28798,N_28904);
or U29480 (N_29480,N_28910,N_28500);
nor U29481 (N_29481,N_28603,N_28824);
or U29482 (N_29482,N_28969,N_28846);
and U29483 (N_29483,N_28816,N_28577);
nor U29484 (N_29484,N_28758,N_28753);
or U29485 (N_29485,N_28782,N_28890);
nor U29486 (N_29486,N_28587,N_28807);
and U29487 (N_29487,N_28591,N_28633);
nor U29488 (N_29488,N_28798,N_28528);
and U29489 (N_29489,N_28724,N_28837);
xor U29490 (N_29490,N_28744,N_28954);
nand U29491 (N_29491,N_28519,N_28929);
and U29492 (N_29492,N_28860,N_28954);
and U29493 (N_29493,N_28548,N_28588);
and U29494 (N_29494,N_28846,N_28719);
nor U29495 (N_29495,N_28694,N_28810);
xnor U29496 (N_29496,N_28698,N_28982);
xor U29497 (N_29497,N_28663,N_28737);
xor U29498 (N_29498,N_28989,N_28900);
xnor U29499 (N_29499,N_28691,N_28963);
nor U29500 (N_29500,N_29151,N_29390);
or U29501 (N_29501,N_29273,N_29185);
nand U29502 (N_29502,N_29055,N_29355);
or U29503 (N_29503,N_29478,N_29346);
nand U29504 (N_29504,N_29018,N_29286);
or U29505 (N_29505,N_29137,N_29143);
and U29506 (N_29506,N_29312,N_29259);
and U29507 (N_29507,N_29369,N_29230);
nand U29508 (N_29508,N_29232,N_29404);
or U29509 (N_29509,N_29172,N_29350);
or U29510 (N_29510,N_29285,N_29224);
xor U29511 (N_29511,N_29041,N_29288);
nor U29512 (N_29512,N_29376,N_29336);
nand U29513 (N_29513,N_29122,N_29193);
and U29514 (N_29514,N_29351,N_29457);
xor U29515 (N_29515,N_29294,N_29091);
or U29516 (N_29516,N_29121,N_29190);
nor U29517 (N_29517,N_29090,N_29277);
and U29518 (N_29518,N_29052,N_29204);
nor U29519 (N_29519,N_29059,N_29363);
or U29520 (N_29520,N_29313,N_29316);
and U29521 (N_29521,N_29419,N_29117);
nand U29522 (N_29522,N_29032,N_29399);
nand U29523 (N_29523,N_29485,N_29301);
and U29524 (N_29524,N_29183,N_29079);
nand U29525 (N_29525,N_29384,N_29153);
and U29526 (N_29526,N_29328,N_29378);
nand U29527 (N_29527,N_29407,N_29292);
xnor U29528 (N_29528,N_29207,N_29422);
nand U29529 (N_29529,N_29472,N_29278);
and U29530 (N_29530,N_29293,N_29499);
nor U29531 (N_29531,N_29130,N_29391);
nor U29532 (N_29532,N_29409,N_29198);
and U29533 (N_29533,N_29157,N_29231);
and U29534 (N_29534,N_29413,N_29053);
and U29535 (N_29535,N_29368,N_29467);
xor U29536 (N_29536,N_29327,N_29221);
or U29537 (N_29537,N_29490,N_29011);
xor U29538 (N_29538,N_29323,N_29210);
and U29539 (N_29539,N_29141,N_29333);
xor U29540 (N_29540,N_29297,N_29003);
or U29541 (N_29541,N_29038,N_29101);
nand U29542 (N_29542,N_29287,N_29021);
xor U29543 (N_29543,N_29206,N_29015);
xor U29544 (N_29544,N_29388,N_29106);
and U29545 (N_29545,N_29116,N_29072);
nand U29546 (N_29546,N_29402,N_29389);
nor U29547 (N_29547,N_29442,N_29337);
xnor U29548 (N_29548,N_29421,N_29353);
or U29549 (N_29549,N_29267,N_29274);
nand U29550 (N_29550,N_29234,N_29161);
nor U29551 (N_29551,N_29096,N_29061);
nand U29552 (N_29552,N_29475,N_29438);
xor U29553 (N_29553,N_29446,N_29058);
xor U29554 (N_29554,N_29086,N_29276);
nand U29555 (N_29555,N_29308,N_29420);
and U29556 (N_29556,N_29160,N_29163);
nor U29557 (N_29557,N_29436,N_29456);
nand U29558 (N_29558,N_29447,N_29361);
or U29559 (N_29559,N_29270,N_29074);
nand U29560 (N_29560,N_29034,N_29441);
xor U29561 (N_29561,N_29129,N_29089);
or U29562 (N_29562,N_29347,N_29497);
or U29563 (N_29563,N_29065,N_29386);
xnor U29564 (N_29564,N_29179,N_29482);
nor U29565 (N_29565,N_29462,N_29480);
xnor U29566 (N_29566,N_29318,N_29245);
and U29567 (N_29567,N_29127,N_29414);
nand U29568 (N_29568,N_29002,N_29178);
nor U29569 (N_29569,N_29395,N_29251);
nor U29570 (N_29570,N_29430,N_29097);
xnor U29571 (N_29571,N_29132,N_29374);
nor U29572 (N_29572,N_29162,N_29289);
and U29573 (N_29573,N_29315,N_29051);
nand U29574 (N_29574,N_29068,N_29281);
nand U29575 (N_29575,N_29334,N_29182);
nor U29576 (N_29576,N_29465,N_29008);
or U29577 (N_29577,N_29240,N_29118);
or U29578 (N_29578,N_29397,N_29254);
xnor U29579 (N_29579,N_29403,N_29145);
xor U29580 (N_29580,N_29266,N_29306);
nand U29581 (N_29581,N_29317,N_29147);
nor U29582 (N_29582,N_29261,N_29071);
and U29583 (N_29583,N_29037,N_29326);
and U29584 (N_29584,N_29426,N_29112);
and U29585 (N_29585,N_29126,N_29216);
nor U29586 (N_29586,N_29233,N_29241);
nor U29587 (N_29587,N_29452,N_29078);
or U29588 (N_29588,N_29335,N_29495);
nor U29589 (N_29589,N_29370,N_29082);
and U29590 (N_29590,N_29484,N_29498);
nand U29591 (N_29591,N_29170,N_29440);
nand U29592 (N_29592,N_29066,N_29060);
or U29593 (N_29593,N_29196,N_29385);
nor U29594 (N_29594,N_29155,N_29494);
or U29595 (N_29595,N_29049,N_29134);
nand U29596 (N_29596,N_29416,N_29022);
xnor U29597 (N_29597,N_29393,N_29105);
nor U29598 (N_29598,N_29464,N_29093);
or U29599 (N_29599,N_29237,N_29275);
and U29600 (N_29600,N_29036,N_29471);
xnor U29601 (N_29601,N_29146,N_29373);
or U29602 (N_29602,N_29283,N_29177);
and U29603 (N_29603,N_29257,N_29476);
xor U29604 (N_29604,N_29030,N_29017);
and U29605 (N_29605,N_29325,N_29213);
or U29606 (N_29606,N_29424,N_29372);
nor U29607 (N_29607,N_29050,N_29144);
and U29608 (N_29608,N_29228,N_29454);
xnor U29609 (N_29609,N_29290,N_29138);
nand U29610 (N_29610,N_29120,N_29453);
and U29611 (N_29611,N_29272,N_29455);
nand U29612 (N_29612,N_29473,N_29026);
nand U29613 (N_29613,N_29295,N_29152);
and U29614 (N_29614,N_29028,N_29062);
xnor U29615 (N_29615,N_29339,N_29045);
and U29616 (N_29616,N_29343,N_29492);
nand U29617 (N_29617,N_29340,N_29321);
nand U29618 (N_29618,N_29394,N_29107);
xor U29619 (N_29619,N_29268,N_29434);
nand U29620 (N_29620,N_29040,N_29262);
xnor U29621 (N_29621,N_29203,N_29165);
and U29622 (N_29622,N_29282,N_29135);
nor U29623 (N_29623,N_29223,N_29449);
nand U29624 (N_29624,N_29010,N_29463);
nor U29625 (N_29625,N_29004,N_29357);
xnor U29626 (N_29626,N_29020,N_29081);
or U29627 (N_29627,N_29077,N_29300);
nor U29628 (N_29628,N_29175,N_29171);
xnor U29629 (N_29629,N_29474,N_29252);
nand U29630 (N_29630,N_29070,N_29487);
or U29631 (N_29631,N_29253,N_29220);
nor U29632 (N_29632,N_29428,N_29481);
nor U29633 (N_29633,N_29310,N_29191);
and U29634 (N_29634,N_29131,N_29387);
or U29635 (N_29635,N_29125,N_29006);
nand U29636 (N_29636,N_29279,N_29298);
nand U29637 (N_29637,N_29095,N_29445);
nand U29638 (N_29638,N_29443,N_29205);
and U29639 (N_29639,N_29417,N_29271);
xnor U29640 (N_29640,N_29149,N_29469);
nor U29641 (N_29641,N_29103,N_29470);
and U29642 (N_29642,N_29007,N_29218);
and U29643 (N_29643,N_29344,N_29451);
or U29644 (N_29644,N_29083,N_29437);
nand U29645 (N_29645,N_29225,N_29263);
and U29646 (N_29646,N_29215,N_29012);
xnor U29647 (N_29647,N_29359,N_29201);
xnor U29648 (N_29648,N_29247,N_29219);
xnor U29649 (N_29649,N_29260,N_29075);
xor U29650 (N_29650,N_29119,N_29319);
or U29651 (N_29651,N_29305,N_29109);
nor U29652 (N_29652,N_29195,N_29330);
xnor U29653 (N_29653,N_29296,N_29444);
nand U29654 (N_29654,N_29354,N_29092);
nand U29655 (N_29655,N_29188,N_29069);
and U29656 (N_29656,N_29212,N_29450);
and U29657 (N_29657,N_29415,N_29358);
xnor U29658 (N_29658,N_29345,N_29189);
and U29659 (N_29659,N_29001,N_29236);
xnor U29660 (N_29660,N_29255,N_29084);
nor U29661 (N_29661,N_29202,N_29379);
nand U29662 (N_29662,N_29168,N_29488);
nor U29663 (N_29663,N_29331,N_29227);
xnor U29664 (N_29664,N_29104,N_29383);
nand U29665 (N_29665,N_29217,N_29375);
nor U29666 (N_29666,N_29024,N_29468);
xnor U29667 (N_29667,N_29329,N_29477);
nor U29668 (N_29668,N_29042,N_29418);
or U29669 (N_29669,N_29114,N_29088);
nand U29670 (N_29670,N_29133,N_29322);
nor U29671 (N_29671,N_29180,N_29159);
nand U29672 (N_29672,N_29029,N_29226);
nor U29673 (N_29673,N_29197,N_29239);
and U29674 (N_29674,N_29158,N_29192);
xnor U29675 (N_29675,N_29039,N_29176);
or U29676 (N_29676,N_29381,N_29269);
nand U29677 (N_29677,N_29238,N_29102);
nand U29678 (N_29678,N_29364,N_29479);
nor U29679 (N_29679,N_29256,N_29187);
nor U29680 (N_29680,N_29338,N_29398);
and U29681 (N_29681,N_29194,N_29087);
or U29682 (N_29682,N_29324,N_29244);
xor U29683 (N_29683,N_29023,N_29148);
xor U29684 (N_29684,N_29076,N_29461);
nor U29685 (N_29685,N_29491,N_29115);
or U29686 (N_29686,N_29320,N_29128);
and U29687 (N_29687,N_29064,N_29200);
or U29688 (N_29688,N_29044,N_29156);
nor U29689 (N_29689,N_29400,N_29307);
or U29690 (N_29690,N_29242,N_29229);
and U29691 (N_29691,N_29167,N_29031);
and U29692 (N_29692,N_29063,N_29164);
nand U29693 (N_29693,N_29166,N_29348);
or U29694 (N_29694,N_29009,N_29405);
nor U29695 (N_29695,N_29140,N_29291);
nor U29696 (N_29696,N_29136,N_29352);
nor U29697 (N_29697,N_29099,N_29408);
xnor U29698 (N_29698,N_29005,N_29433);
nor U29699 (N_29699,N_29284,N_29098);
nor U29700 (N_29700,N_29110,N_29342);
or U29701 (N_29701,N_29489,N_29458);
nand U29702 (N_29702,N_29214,N_29341);
and U29703 (N_29703,N_29332,N_29264);
nor U29704 (N_29704,N_29265,N_29067);
nor U29705 (N_29705,N_29249,N_29460);
xnor U29706 (N_29706,N_29448,N_29142);
xnor U29707 (N_29707,N_29435,N_29243);
nor U29708 (N_29708,N_29124,N_29173);
nor U29709 (N_29709,N_29432,N_29427);
or U29710 (N_29710,N_29056,N_29280);
nand U29711 (N_29711,N_29123,N_29033);
nor U29712 (N_29712,N_29392,N_29303);
xnor U29713 (N_29713,N_29365,N_29483);
nor U29714 (N_29714,N_29186,N_29043);
or U29715 (N_29715,N_29013,N_29396);
or U29716 (N_29716,N_29429,N_29139);
nor U29717 (N_29717,N_29169,N_29150);
xor U29718 (N_29718,N_29073,N_29154);
nor U29719 (N_29719,N_29356,N_29486);
nor U29720 (N_29720,N_29439,N_29094);
nand U29721 (N_29721,N_29360,N_29406);
nor U29722 (N_29722,N_29248,N_29367);
nor U29723 (N_29723,N_29035,N_29211);
or U29724 (N_29724,N_29493,N_29184);
xor U29725 (N_29725,N_29047,N_29208);
and U29726 (N_29726,N_29401,N_29246);
and U29727 (N_29727,N_29377,N_29431);
nor U29728 (N_29728,N_29100,N_29054);
nor U29729 (N_29729,N_29309,N_29411);
xor U29730 (N_29730,N_29025,N_29048);
or U29731 (N_29731,N_29250,N_29366);
nand U29732 (N_29732,N_29113,N_29371);
xnor U29733 (N_29733,N_29027,N_29019);
xnor U29734 (N_29734,N_29496,N_29199);
xnor U29735 (N_29735,N_29111,N_29174);
or U29736 (N_29736,N_29425,N_29080);
nor U29737 (N_29737,N_29382,N_29108);
and U29738 (N_29738,N_29046,N_29181);
nand U29739 (N_29739,N_29410,N_29209);
xor U29740 (N_29740,N_29459,N_29235);
nand U29741 (N_29741,N_29380,N_29014);
xnor U29742 (N_29742,N_29302,N_29016);
and U29743 (N_29743,N_29412,N_29222);
xnor U29744 (N_29744,N_29423,N_29258);
and U29745 (N_29745,N_29314,N_29311);
nand U29746 (N_29746,N_29057,N_29304);
nand U29747 (N_29747,N_29299,N_29466);
nand U29748 (N_29748,N_29000,N_29085);
xnor U29749 (N_29749,N_29349,N_29362);
xor U29750 (N_29750,N_29068,N_29149);
xnor U29751 (N_29751,N_29468,N_29354);
nand U29752 (N_29752,N_29188,N_29193);
xnor U29753 (N_29753,N_29189,N_29307);
nand U29754 (N_29754,N_29067,N_29300);
nand U29755 (N_29755,N_29214,N_29091);
xor U29756 (N_29756,N_29462,N_29254);
nor U29757 (N_29757,N_29481,N_29070);
nor U29758 (N_29758,N_29383,N_29043);
or U29759 (N_29759,N_29427,N_29228);
or U29760 (N_29760,N_29016,N_29116);
xnor U29761 (N_29761,N_29304,N_29176);
nor U29762 (N_29762,N_29004,N_29213);
nor U29763 (N_29763,N_29310,N_29002);
or U29764 (N_29764,N_29305,N_29067);
xnor U29765 (N_29765,N_29346,N_29019);
or U29766 (N_29766,N_29269,N_29095);
nand U29767 (N_29767,N_29475,N_29090);
or U29768 (N_29768,N_29437,N_29338);
or U29769 (N_29769,N_29385,N_29008);
nor U29770 (N_29770,N_29291,N_29340);
nand U29771 (N_29771,N_29422,N_29437);
xnor U29772 (N_29772,N_29392,N_29258);
xor U29773 (N_29773,N_29329,N_29103);
or U29774 (N_29774,N_29448,N_29447);
or U29775 (N_29775,N_29478,N_29372);
xor U29776 (N_29776,N_29112,N_29128);
nor U29777 (N_29777,N_29074,N_29202);
nand U29778 (N_29778,N_29193,N_29463);
and U29779 (N_29779,N_29068,N_29042);
nand U29780 (N_29780,N_29154,N_29408);
xnor U29781 (N_29781,N_29091,N_29171);
and U29782 (N_29782,N_29082,N_29291);
or U29783 (N_29783,N_29156,N_29356);
and U29784 (N_29784,N_29410,N_29048);
nand U29785 (N_29785,N_29356,N_29307);
nor U29786 (N_29786,N_29426,N_29340);
and U29787 (N_29787,N_29052,N_29224);
nand U29788 (N_29788,N_29431,N_29041);
and U29789 (N_29789,N_29050,N_29280);
xnor U29790 (N_29790,N_29304,N_29449);
or U29791 (N_29791,N_29430,N_29103);
nand U29792 (N_29792,N_29342,N_29251);
xor U29793 (N_29793,N_29330,N_29111);
nor U29794 (N_29794,N_29219,N_29288);
nor U29795 (N_29795,N_29266,N_29095);
nor U29796 (N_29796,N_29355,N_29173);
nand U29797 (N_29797,N_29365,N_29425);
or U29798 (N_29798,N_29015,N_29163);
xnor U29799 (N_29799,N_29103,N_29399);
xnor U29800 (N_29800,N_29167,N_29242);
nand U29801 (N_29801,N_29246,N_29231);
and U29802 (N_29802,N_29312,N_29081);
nor U29803 (N_29803,N_29394,N_29022);
or U29804 (N_29804,N_29388,N_29160);
or U29805 (N_29805,N_29349,N_29398);
nand U29806 (N_29806,N_29170,N_29328);
and U29807 (N_29807,N_29291,N_29165);
or U29808 (N_29808,N_29099,N_29385);
nand U29809 (N_29809,N_29040,N_29410);
and U29810 (N_29810,N_29478,N_29330);
xnor U29811 (N_29811,N_29083,N_29146);
nor U29812 (N_29812,N_29435,N_29255);
nand U29813 (N_29813,N_29008,N_29167);
or U29814 (N_29814,N_29190,N_29390);
and U29815 (N_29815,N_29467,N_29389);
nand U29816 (N_29816,N_29219,N_29416);
and U29817 (N_29817,N_29199,N_29418);
nor U29818 (N_29818,N_29339,N_29150);
and U29819 (N_29819,N_29006,N_29410);
or U29820 (N_29820,N_29362,N_29473);
nor U29821 (N_29821,N_29162,N_29209);
nand U29822 (N_29822,N_29416,N_29036);
or U29823 (N_29823,N_29077,N_29285);
and U29824 (N_29824,N_29294,N_29314);
or U29825 (N_29825,N_29250,N_29046);
or U29826 (N_29826,N_29356,N_29424);
xor U29827 (N_29827,N_29009,N_29312);
or U29828 (N_29828,N_29198,N_29290);
nor U29829 (N_29829,N_29024,N_29417);
nor U29830 (N_29830,N_29361,N_29355);
nand U29831 (N_29831,N_29084,N_29333);
or U29832 (N_29832,N_29335,N_29044);
nand U29833 (N_29833,N_29192,N_29150);
or U29834 (N_29834,N_29348,N_29032);
nor U29835 (N_29835,N_29130,N_29453);
nor U29836 (N_29836,N_29000,N_29314);
or U29837 (N_29837,N_29361,N_29453);
and U29838 (N_29838,N_29246,N_29422);
xnor U29839 (N_29839,N_29302,N_29445);
nor U29840 (N_29840,N_29261,N_29030);
nor U29841 (N_29841,N_29035,N_29451);
and U29842 (N_29842,N_29487,N_29190);
and U29843 (N_29843,N_29110,N_29433);
nor U29844 (N_29844,N_29351,N_29121);
or U29845 (N_29845,N_29371,N_29440);
nand U29846 (N_29846,N_29151,N_29316);
or U29847 (N_29847,N_29041,N_29091);
nor U29848 (N_29848,N_29057,N_29107);
nand U29849 (N_29849,N_29272,N_29090);
xnor U29850 (N_29850,N_29105,N_29042);
or U29851 (N_29851,N_29184,N_29105);
or U29852 (N_29852,N_29437,N_29056);
and U29853 (N_29853,N_29413,N_29464);
or U29854 (N_29854,N_29141,N_29210);
or U29855 (N_29855,N_29343,N_29334);
and U29856 (N_29856,N_29435,N_29298);
or U29857 (N_29857,N_29284,N_29291);
and U29858 (N_29858,N_29352,N_29089);
nand U29859 (N_29859,N_29481,N_29326);
xor U29860 (N_29860,N_29471,N_29158);
and U29861 (N_29861,N_29231,N_29270);
xnor U29862 (N_29862,N_29077,N_29450);
or U29863 (N_29863,N_29492,N_29337);
nand U29864 (N_29864,N_29272,N_29443);
nor U29865 (N_29865,N_29213,N_29314);
nand U29866 (N_29866,N_29011,N_29108);
nor U29867 (N_29867,N_29093,N_29289);
or U29868 (N_29868,N_29358,N_29077);
and U29869 (N_29869,N_29029,N_29033);
and U29870 (N_29870,N_29285,N_29164);
nand U29871 (N_29871,N_29420,N_29180);
and U29872 (N_29872,N_29410,N_29267);
or U29873 (N_29873,N_29156,N_29345);
nor U29874 (N_29874,N_29372,N_29233);
nand U29875 (N_29875,N_29254,N_29250);
xnor U29876 (N_29876,N_29268,N_29439);
nand U29877 (N_29877,N_29125,N_29136);
nor U29878 (N_29878,N_29101,N_29417);
or U29879 (N_29879,N_29152,N_29127);
or U29880 (N_29880,N_29130,N_29081);
nor U29881 (N_29881,N_29376,N_29374);
and U29882 (N_29882,N_29272,N_29171);
xnor U29883 (N_29883,N_29143,N_29056);
xor U29884 (N_29884,N_29339,N_29128);
xor U29885 (N_29885,N_29087,N_29137);
xnor U29886 (N_29886,N_29049,N_29117);
or U29887 (N_29887,N_29401,N_29055);
and U29888 (N_29888,N_29454,N_29003);
nand U29889 (N_29889,N_29301,N_29401);
xor U29890 (N_29890,N_29171,N_29212);
nand U29891 (N_29891,N_29397,N_29153);
nor U29892 (N_29892,N_29383,N_29018);
nand U29893 (N_29893,N_29012,N_29409);
nor U29894 (N_29894,N_29405,N_29387);
nor U29895 (N_29895,N_29174,N_29060);
or U29896 (N_29896,N_29379,N_29464);
or U29897 (N_29897,N_29065,N_29196);
xnor U29898 (N_29898,N_29063,N_29365);
nor U29899 (N_29899,N_29215,N_29037);
nor U29900 (N_29900,N_29249,N_29451);
or U29901 (N_29901,N_29063,N_29080);
nor U29902 (N_29902,N_29289,N_29029);
nor U29903 (N_29903,N_29356,N_29038);
nor U29904 (N_29904,N_29413,N_29216);
or U29905 (N_29905,N_29164,N_29186);
xnor U29906 (N_29906,N_29076,N_29426);
or U29907 (N_29907,N_29001,N_29454);
and U29908 (N_29908,N_29138,N_29187);
xnor U29909 (N_29909,N_29102,N_29434);
or U29910 (N_29910,N_29433,N_29009);
or U29911 (N_29911,N_29310,N_29307);
and U29912 (N_29912,N_29277,N_29271);
and U29913 (N_29913,N_29132,N_29428);
and U29914 (N_29914,N_29484,N_29263);
xor U29915 (N_29915,N_29476,N_29130);
xor U29916 (N_29916,N_29496,N_29495);
nand U29917 (N_29917,N_29464,N_29042);
or U29918 (N_29918,N_29022,N_29226);
nor U29919 (N_29919,N_29253,N_29373);
nor U29920 (N_29920,N_29051,N_29386);
nand U29921 (N_29921,N_29361,N_29226);
nand U29922 (N_29922,N_29271,N_29013);
nor U29923 (N_29923,N_29112,N_29121);
nand U29924 (N_29924,N_29306,N_29059);
or U29925 (N_29925,N_29406,N_29123);
or U29926 (N_29926,N_29243,N_29246);
or U29927 (N_29927,N_29462,N_29251);
and U29928 (N_29928,N_29240,N_29489);
and U29929 (N_29929,N_29000,N_29385);
or U29930 (N_29930,N_29080,N_29110);
xnor U29931 (N_29931,N_29106,N_29497);
and U29932 (N_29932,N_29254,N_29061);
or U29933 (N_29933,N_29238,N_29237);
or U29934 (N_29934,N_29154,N_29413);
and U29935 (N_29935,N_29023,N_29137);
nand U29936 (N_29936,N_29082,N_29060);
nor U29937 (N_29937,N_29308,N_29340);
xnor U29938 (N_29938,N_29459,N_29098);
xor U29939 (N_29939,N_29422,N_29283);
xnor U29940 (N_29940,N_29142,N_29096);
and U29941 (N_29941,N_29378,N_29465);
or U29942 (N_29942,N_29033,N_29269);
or U29943 (N_29943,N_29111,N_29006);
xnor U29944 (N_29944,N_29211,N_29131);
and U29945 (N_29945,N_29401,N_29380);
and U29946 (N_29946,N_29010,N_29122);
nor U29947 (N_29947,N_29494,N_29230);
nor U29948 (N_29948,N_29466,N_29008);
nand U29949 (N_29949,N_29149,N_29161);
nor U29950 (N_29950,N_29055,N_29329);
nor U29951 (N_29951,N_29395,N_29400);
nor U29952 (N_29952,N_29205,N_29364);
nand U29953 (N_29953,N_29062,N_29203);
nor U29954 (N_29954,N_29221,N_29249);
nand U29955 (N_29955,N_29382,N_29494);
nor U29956 (N_29956,N_29381,N_29400);
xor U29957 (N_29957,N_29218,N_29282);
or U29958 (N_29958,N_29484,N_29273);
xnor U29959 (N_29959,N_29310,N_29473);
nor U29960 (N_29960,N_29071,N_29341);
xnor U29961 (N_29961,N_29024,N_29485);
nand U29962 (N_29962,N_29222,N_29078);
xor U29963 (N_29963,N_29037,N_29078);
nor U29964 (N_29964,N_29460,N_29064);
and U29965 (N_29965,N_29307,N_29435);
and U29966 (N_29966,N_29040,N_29484);
xnor U29967 (N_29967,N_29238,N_29184);
nor U29968 (N_29968,N_29129,N_29030);
and U29969 (N_29969,N_29060,N_29439);
nand U29970 (N_29970,N_29288,N_29296);
nand U29971 (N_29971,N_29296,N_29147);
nand U29972 (N_29972,N_29384,N_29470);
xor U29973 (N_29973,N_29126,N_29061);
or U29974 (N_29974,N_29093,N_29388);
and U29975 (N_29975,N_29348,N_29401);
or U29976 (N_29976,N_29028,N_29358);
xnor U29977 (N_29977,N_29156,N_29205);
nand U29978 (N_29978,N_29279,N_29013);
xor U29979 (N_29979,N_29274,N_29194);
nand U29980 (N_29980,N_29121,N_29041);
xnor U29981 (N_29981,N_29315,N_29403);
or U29982 (N_29982,N_29187,N_29071);
or U29983 (N_29983,N_29264,N_29307);
nand U29984 (N_29984,N_29310,N_29217);
nor U29985 (N_29985,N_29175,N_29208);
nand U29986 (N_29986,N_29408,N_29364);
xor U29987 (N_29987,N_29231,N_29478);
nand U29988 (N_29988,N_29397,N_29474);
nor U29989 (N_29989,N_29146,N_29106);
and U29990 (N_29990,N_29118,N_29010);
nor U29991 (N_29991,N_29197,N_29115);
xor U29992 (N_29992,N_29493,N_29475);
or U29993 (N_29993,N_29079,N_29242);
xnor U29994 (N_29994,N_29185,N_29032);
or U29995 (N_29995,N_29394,N_29009);
nor U29996 (N_29996,N_29276,N_29310);
nor U29997 (N_29997,N_29421,N_29427);
and U29998 (N_29998,N_29171,N_29476);
xor U29999 (N_29999,N_29154,N_29354);
nor UO_0 (O_0,N_29598,N_29984);
nand UO_1 (O_1,N_29756,N_29736);
nor UO_2 (O_2,N_29986,N_29882);
xor UO_3 (O_3,N_29716,N_29715);
xor UO_4 (O_4,N_29798,N_29722);
nor UO_5 (O_5,N_29668,N_29837);
xor UO_6 (O_6,N_29849,N_29703);
and UO_7 (O_7,N_29966,N_29794);
xnor UO_8 (O_8,N_29556,N_29990);
or UO_9 (O_9,N_29602,N_29840);
and UO_10 (O_10,N_29777,N_29909);
xor UO_11 (O_11,N_29856,N_29779);
nand UO_12 (O_12,N_29510,N_29859);
and UO_13 (O_13,N_29573,N_29612);
nor UO_14 (O_14,N_29737,N_29910);
and UO_15 (O_15,N_29818,N_29525);
xnor UO_16 (O_16,N_29652,N_29620);
xnor UO_17 (O_17,N_29554,N_29877);
and UO_18 (O_18,N_29871,N_29797);
xnor UO_19 (O_19,N_29610,N_29952);
nand UO_20 (O_20,N_29985,N_29650);
and UO_21 (O_21,N_29613,N_29531);
nand UO_22 (O_22,N_29862,N_29567);
xor UO_23 (O_23,N_29561,N_29568);
and UO_24 (O_24,N_29635,N_29894);
nor UO_25 (O_25,N_29532,N_29653);
nor UO_26 (O_26,N_29796,N_29606);
nand UO_27 (O_27,N_29884,N_29900);
nand UO_28 (O_28,N_29754,N_29747);
nor UO_29 (O_29,N_29762,N_29964);
or UO_30 (O_30,N_29816,N_29608);
nand UO_31 (O_31,N_29979,N_29681);
and UO_32 (O_32,N_29908,N_29911);
nor UO_33 (O_33,N_29592,N_29898);
or UO_34 (O_34,N_29834,N_29727);
or UO_35 (O_35,N_29582,N_29508);
xnor UO_36 (O_36,N_29790,N_29746);
xnor UO_37 (O_37,N_29583,N_29999);
nor UO_38 (O_38,N_29698,N_29920);
and UO_39 (O_39,N_29804,N_29629);
nand UO_40 (O_40,N_29923,N_29850);
nand UO_41 (O_41,N_29551,N_29994);
nor UO_42 (O_42,N_29874,N_29899);
xnor UO_43 (O_43,N_29578,N_29667);
nand UO_44 (O_44,N_29671,N_29868);
xnor UO_45 (O_45,N_29648,N_29555);
nor UO_46 (O_46,N_29546,N_29872);
nor UO_47 (O_47,N_29824,N_29593);
xnor UO_48 (O_48,N_29757,N_29596);
and UO_49 (O_49,N_29765,N_29748);
xnor UO_50 (O_50,N_29811,N_29623);
xnor UO_51 (O_51,N_29883,N_29584);
or UO_52 (O_52,N_29530,N_29505);
nand UO_53 (O_53,N_29538,N_29970);
nand UO_54 (O_54,N_29625,N_29502);
nor UO_55 (O_55,N_29776,N_29692);
nor UO_56 (O_56,N_29517,N_29822);
nand UO_57 (O_57,N_29792,N_29574);
nor UO_58 (O_58,N_29861,N_29697);
nor UO_59 (O_59,N_29518,N_29627);
or UO_60 (O_60,N_29763,N_29604);
or UO_61 (O_61,N_29649,N_29809);
nand UO_62 (O_62,N_29702,N_29624);
nor UO_63 (O_63,N_29563,N_29634);
and UO_64 (O_64,N_29904,N_29944);
or UO_65 (O_65,N_29768,N_29988);
xnor UO_66 (O_66,N_29646,N_29553);
xnor UO_67 (O_67,N_29847,N_29549);
nor UO_68 (O_68,N_29934,N_29526);
nand UO_69 (O_69,N_29865,N_29921);
nand UO_70 (O_70,N_29742,N_29562);
xor UO_71 (O_71,N_29889,N_29577);
or UO_72 (O_72,N_29683,N_29838);
or UO_73 (O_73,N_29600,N_29548);
xnor UO_74 (O_74,N_29619,N_29954);
nor UO_75 (O_75,N_29951,N_29643);
and UO_76 (O_76,N_29689,N_29784);
and UO_77 (O_77,N_29786,N_29719);
nand UO_78 (O_78,N_29626,N_29977);
and UO_79 (O_79,N_29971,N_29879);
xor UO_80 (O_80,N_29841,N_29915);
or UO_81 (O_81,N_29739,N_29806);
xnor UO_82 (O_82,N_29559,N_29659);
xor UO_83 (O_83,N_29942,N_29672);
xnor UO_84 (O_84,N_29919,N_29521);
and UO_85 (O_85,N_29750,N_29789);
nor UO_86 (O_86,N_29867,N_29922);
xnor UO_87 (O_87,N_29654,N_29744);
and UO_88 (O_88,N_29876,N_29607);
and UO_89 (O_89,N_29983,N_29959);
and UO_90 (O_90,N_29647,N_29903);
nand UO_91 (O_91,N_29881,N_29886);
nand UO_92 (O_92,N_29938,N_29890);
and UO_93 (O_93,N_29718,N_29611);
and UO_94 (O_94,N_29957,N_29860);
and UO_95 (O_95,N_29699,N_29560);
nand UO_96 (O_96,N_29541,N_29972);
and UO_97 (O_97,N_29677,N_29975);
and UO_98 (O_98,N_29793,N_29773);
xnor UO_99 (O_99,N_29805,N_29543);
xor UO_100 (O_100,N_29520,N_29863);
nor UO_101 (O_101,N_29812,N_29946);
or UO_102 (O_102,N_29769,N_29925);
xor UO_103 (O_103,N_29767,N_29726);
or UO_104 (O_104,N_29760,N_29933);
and UO_105 (O_105,N_29707,N_29914);
or UO_106 (O_106,N_29992,N_29945);
nor UO_107 (O_107,N_29950,N_29527);
nand UO_108 (O_108,N_29766,N_29690);
xor UO_109 (O_109,N_29522,N_29993);
nor UO_110 (O_110,N_29755,N_29693);
and UO_111 (O_111,N_29571,N_29981);
nand UO_112 (O_112,N_29803,N_29953);
nor UO_113 (O_113,N_29674,N_29928);
and UO_114 (O_114,N_29982,N_29752);
or UO_115 (O_115,N_29775,N_29829);
xnor UO_116 (O_116,N_29733,N_29980);
nor UO_117 (O_117,N_29570,N_29597);
nor UO_118 (O_118,N_29545,N_29800);
or UO_119 (O_119,N_29708,N_29615);
and UO_120 (O_120,N_29580,N_29887);
and UO_121 (O_121,N_29529,N_29632);
or UO_122 (O_122,N_29636,N_29720);
xnor UO_123 (O_123,N_29851,N_29997);
nand UO_124 (O_124,N_29967,N_29658);
nand UO_125 (O_125,N_29761,N_29701);
nor UO_126 (O_126,N_29717,N_29565);
nor UO_127 (O_127,N_29687,N_29732);
or UO_128 (O_128,N_29869,N_29682);
nor UO_129 (O_129,N_29758,N_29873);
nor UO_130 (O_130,N_29936,N_29503);
and UO_131 (O_131,N_29519,N_29590);
nand UO_132 (O_132,N_29641,N_29864);
nor UO_133 (O_133,N_29855,N_29723);
xnor UO_134 (O_134,N_29947,N_29644);
nand UO_135 (O_135,N_29956,N_29588);
xor UO_136 (O_136,N_29516,N_29845);
xnor UO_137 (O_137,N_29704,N_29601);
or UO_138 (O_138,N_29738,N_29891);
or UO_139 (O_139,N_29963,N_29534);
and UO_140 (O_140,N_29536,N_29791);
or UO_141 (O_141,N_29528,N_29509);
nor UO_142 (O_142,N_29948,N_29506);
and UO_143 (O_143,N_29991,N_29848);
nor UO_144 (O_144,N_29550,N_29637);
nand UO_145 (O_145,N_29655,N_29617);
or UO_146 (O_146,N_29741,N_29788);
and UO_147 (O_147,N_29735,N_29572);
and UO_148 (O_148,N_29638,N_29996);
nor UO_149 (O_149,N_29675,N_29815);
and UO_150 (O_150,N_29857,N_29616);
or UO_151 (O_151,N_29770,N_29622);
or UO_152 (O_152,N_29751,N_29599);
nand UO_153 (O_153,N_29853,N_29844);
nor UO_154 (O_154,N_29830,N_29673);
or UO_155 (O_155,N_29662,N_29783);
xor UO_156 (O_156,N_29621,N_29913);
xor UO_157 (O_157,N_29524,N_29594);
and UO_158 (O_158,N_29795,N_29749);
nand UO_159 (O_159,N_29579,N_29552);
nor UO_160 (O_160,N_29513,N_29817);
and UO_161 (O_161,N_29895,N_29709);
xor UO_162 (O_162,N_29745,N_29771);
xnor UO_163 (O_163,N_29680,N_29810);
xnor UO_164 (O_164,N_29962,N_29827);
xnor UO_165 (O_165,N_29927,N_29535);
nand UO_166 (O_166,N_29603,N_29631);
xor UO_167 (O_167,N_29888,N_29633);
nor UO_168 (O_168,N_29721,N_29614);
nor UO_169 (O_169,N_29686,N_29897);
and UO_170 (O_170,N_29696,N_29780);
and UO_171 (O_171,N_29778,N_29968);
nor UO_172 (O_172,N_29586,N_29918);
nand UO_173 (O_173,N_29842,N_29581);
xnor UO_174 (O_174,N_29670,N_29782);
nand UO_175 (O_175,N_29833,N_29669);
and UO_176 (O_176,N_29935,N_29866);
or UO_177 (O_177,N_29905,N_29896);
and UO_178 (O_178,N_29729,N_29640);
and UO_179 (O_179,N_29839,N_29825);
nor UO_180 (O_180,N_29685,N_29504);
or UO_181 (O_181,N_29916,N_29802);
nand UO_182 (O_182,N_29878,N_29743);
xnor UO_183 (O_183,N_29605,N_29835);
or UO_184 (O_184,N_29511,N_29700);
or UO_185 (O_185,N_29730,N_29679);
xnor UO_186 (O_186,N_29912,N_29892);
nand UO_187 (O_187,N_29514,N_29772);
and UO_188 (O_188,N_29901,N_29836);
or UO_189 (O_189,N_29706,N_29907);
and UO_190 (O_190,N_29846,N_29774);
nand UO_191 (O_191,N_29870,N_29808);
or UO_192 (O_192,N_29595,N_29820);
and UO_193 (O_193,N_29998,N_29566);
xor UO_194 (O_194,N_29712,N_29926);
or UO_195 (O_195,N_29710,N_29569);
xor UO_196 (O_196,N_29821,N_29585);
xor UO_197 (O_197,N_29929,N_29828);
or UO_198 (O_198,N_29759,N_29724);
nand UO_199 (O_199,N_29656,N_29941);
or UO_200 (O_200,N_29955,N_29533);
nor UO_201 (O_201,N_29875,N_29819);
and UO_202 (O_202,N_29695,N_29558);
nand UO_203 (O_203,N_29575,N_29960);
and UO_204 (O_204,N_29930,N_29725);
and UO_205 (O_205,N_29661,N_29691);
nand UO_206 (O_206,N_29801,N_29937);
nand UO_207 (O_207,N_29714,N_29501);
nand UO_208 (O_208,N_29740,N_29665);
or UO_209 (O_209,N_29978,N_29540);
xor UO_210 (O_210,N_29987,N_29932);
and UO_211 (O_211,N_29564,N_29523);
nand UO_212 (O_212,N_29630,N_29576);
xnor UO_213 (O_213,N_29547,N_29974);
xnor UO_214 (O_214,N_29807,N_29642);
and UO_215 (O_215,N_29678,N_29753);
and UO_216 (O_216,N_29591,N_29628);
or UO_217 (O_217,N_29666,N_29858);
and UO_218 (O_218,N_29813,N_29973);
xor UO_219 (O_219,N_29734,N_29684);
xnor UO_220 (O_220,N_29976,N_29969);
or UO_221 (O_221,N_29832,N_29852);
nand UO_222 (O_222,N_29949,N_29542);
xor UO_223 (O_223,N_29711,N_29557);
or UO_224 (O_224,N_29826,N_29544);
nand UO_225 (O_225,N_29799,N_29664);
nor UO_226 (O_226,N_29814,N_29943);
nor UO_227 (O_227,N_29764,N_29728);
nor UO_228 (O_228,N_29515,N_29589);
xor UO_229 (O_229,N_29939,N_29537);
nor UO_230 (O_230,N_29651,N_29781);
nor UO_231 (O_231,N_29843,N_29609);
nand UO_232 (O_232,N_29906,N_29639);
or UO_233 (O_233,N_29688,N_29995);
xor UO_234 (O_234,N_29940,N_29965);
nand UO_235 (O_235,N_29785,N_29660);
and UO_236 (O_236,N_29618,N_29587);
nor UO_237 (O_237,N_29961,N_29989);
and UO_238 (O_238,N_29500,N_29958);
or UO_239 (O_239,N_29507,N_29657);
and UO_240 (O_240,N_29885,N_29823);
or UO_241 (O_241,N_29917,N_29512);
and UO_242 (O_242,N_29663,N_29893);
nand UO_243 (O_243,N_29676,N_29924);
nor UO_244 (O_244,N_29787,N_29880);
and UO_245 (O_245,N_29854,N_29694);
nor UO_246 (O_246,N_29713,N_29645);
xnor UO_247 (O_247,N_29731,N_29931);
or UO_248 (O_248,N_29539,N_29705);
nor UO_249 (O_249,N_29831,N_29902);
nor UO_250 (O_250,N_29770,N_29816);
nor UO_251 (O_251,N_29746,N_29712);
nor UO_252 (O_252,N_29790,N_29533);
xnor UO_253 (O_253,N_29743,N_29791);
nor UO_254 (O_254,N_29542,N_29950);
nand UO_255 (O_255,N_29859,N_29567);
and UO_256 (O_256,N_29684,N_29940);
nand UO_257 (O_257,N_29608,N_29876);
and UO_258 (O_258,N_29638,N_29595);
or UO_259 (O_259,N_29795,N_29834);
xor UO_260 (O_260,N_29795,N_29915);
nand UO_261 (O_261,N_29738,N_29539);
nand UO_262 (O_262,N_29702,N_29524);
nor UO_263 (O_263,N_29769,N_29781);
xnor UO_264 (O_264,N_29602,N_29682);
nor UO_265 (O_265,N_29674,N_29564);
or UO_266 (O_266,N_29898,N_29590);
nand UO_267 (O_267,N_29651,N_29518);
nand UO_268 (O_268,N_29638,N_29849);
nor UO_269 (O_269,N_29525,N_29522);
nand UO_270 (O_270,N_29683,N_29908);
or UO_271 (O_271,N_29890,N_29967);
nor UO_272 (O_272,N_29909,N_29762);
nor UO_273 (O_273,N_29506,N_29743);
xnor UO_274 (O_274,N_29513,N_29833);
and UO_275 (O_275,N_29618,N_29832);
nand UO_276 (O_276,N_29619,N_29850);
nand UO_277 (O_277,N_29808,N_29731);
xor UO_278 (O_278,N_29544,N_29579);
xnor UO_279 (O_279,N_29710,N_29923);
xor UO_280 (O_280,N_29598,N_29664);
xor UO_281 (O_281,N_29785,N_29603);
and UO_282 (O_282,N_29673,N_29525);
and UO_283 (O_283,N_29837,N_29701);
nand UO_284 (O_284,N_29581,N_29851);
xor UO_285 (O_285,N_29572,N_29988);
nor UO_286 (O_286,N_29954,N_29650);
nor UO_287 (O_287,N_29797,N_29979);
nand UO_288 (O_288,N_29863,N_29782);
nor UO_289 (O_289,N_29837,N_29959);
nor UO_290 (O_290,N_29714,N_29724);
xnor UO_291 (O_291,N_29778,N_29501);
and UO_292 (O_292,N_29679,N_29531);
xor UO_293 (O_293,N_29991,N_29669);
nand UO_294 (O_294,N_29712,N_29642);
xnor UO_295 (O_295,N_29888,N_29716);
nor UO_296 (O_296,N_29723,N_29827);
or UO_297 (O_297,N_29589,N_29925);
nand UO_298 (O_298,N_29953,N_29610);
or UO_299 (O_299,N_29639,N_29955);
or UO_300 (O_300,N_29758,N_29501);
or UO_301 (O_301,N_29885,N_29899);
or UO_302 (O_302,N_29978,N_29523);
nor UO_303 (O_303,N_29562,N_29673);
or UO_304 (O_304,N_29572,N_29609);
or UO_305 (O_305,N_29525,N_29527);
or UO_306 (O_306,N_29764,N_29978);
or UO_307 (O_307,N_29610,N_29509);
nand UO_308 (O_308,N_29711,N_29797);
nor UO_309 (O_309,N_29857,N_29697);
xnor UO_310 (O_310,N_29935,N_29944);
nand UO_311 (O_311,N_29843,N_29765);
xor UO_312 (O_312,N_29613,N_29670);
and UO_313 (O_313,N_29992,N_29884);
or UO_314 (O_314,N_29977,N_29951);
or UO_315 (O_315,N_29905,N_29635);
and UO_316 (O_316,N_29676,N_29566);
nor UO_317 (O_317,N_29679,N_29753);
xor UO_318 (O_318,N_29552,N_29903);
nand UO_319 (O_319,N_29970,N_29829);
and UO_320 (O_320,N_29567,N_29999);
nor UO_321 (O_321,N_29725,N_29723);
nor UO_322 (O_322,N_29591,N_29747);
nor UO_323 (O_323,N_29855,N_29922);
xnor UO_324 (O_324,N_29851,N_29743);
or UO_325 (O_325,N_29614,N_29805);
or UO_326 (O_326,N_29993,N_29617);
nor UO_327 (O_327,N_29967,N_29642);
or UO_328 (O_328,N_29877,N_29625);
or UO_329 (O_329,N_29676,N_29734);
and UO_330 (O_330,N_29805,N_29943);
nor UO_331 (O_331,N_29801,N_29629);
and UO_332 (O_332,N_29889,N_29825);
nor UO_333 (O_333,N_29832,N_29538);
nor UO_334 (O_334,N_29615,N_29691);
and UO_335 (O_335,N_29770,N_29822);
or UO_336 (O_336,N_29688,N_29690);
xor UO_337 (O_337,N_29915,N_29734);
or UO_338 (O_338,N_29649,N_29783);
or UO_339 (O_339,N_29888,N_29829);
xnor UO_340 (O_340,N_29605,N_29614);
and UO_341 (O_341,N_29960,N_29945);
xnor UO_342 (O_342,N_29771,N_29917);
or UO_343 (O_343,N_29989,N_29580);
or UO_344 (O_344,N_29713,N_29519);
and UO_345 (O_345,N_29626,N_29993);
xnor UO_346 (O_346,N_29750,N_29844);
nor UO_347 (O_347,N_29682,N_29799);
or UO_348 (O_348,N_29778,N_29610);
xor UO_349 (O_349,N_29985,N_29906);
and UO_350 (O_350,N_29626,N_29583);
xnor UO_351 (O_351,N_29880,N_29614);
or UO_352 (O_352,N_29742,N_29869);
nand UO_353 (O_353,N_29688,N_29981);
nor UO_354 (O_354,N_29936,N_29683);
xor UO_355 (O_355,N_29964,N_29546);
nor UO_356 (O_356,N_29692,N_29588);
xnor UO_357 (O_357,N_29726,N_29984);
nand UO_358 (O_358,N_29671,N_29590);
and UO_359 (O_359,N_29528,N_29650);
xnor UO_360 (O_360,N_29880,N_29694);
xor UO_361 (O_361,N_29511,N_29695);
and UO_362 (O_362,N_29812,N_29545);
or UO_363 (O_363,N_29522,N_29628);
nor UO_364 (O_364,N_29987,N_29622);
and UO_365 (O_365,N_29684,N_29593);
or UO_366 (O_366,N_29708,N_29553);
and UO_367 (O_367,N_29504,N_29582);
nand UO_368 (O_368,N_29842,N_29725);
nor UO_369 (O_369,N_29622,N_29884);
or UO_370 (O_370,N_29579,N_29639);
or UO_371 (O_371,N_29531,N_29712);
and UO_372 (O_372,N_29628,N_29653);
or UO_373 (O_373,N_29647,N_29599);
nor UO_374 (O_374,N_29957,N_29772);
and UO_375 (O_375,N_29760,N_29834);
or UO_376 (O_376,N_29624,N_29771);
and UO_377 (O_377,N_29836,N_29845);
xnor UO_378 (O_378,N_29885,N_29902);
nor UO_379 (O_379,N_29622,N_29907);
or UO_380 (O_380,N_29825,N_29556);
xor UO_381 (O_381,N_29839,N_29924);
nand UO_382 (O_382,N_29546,N_29740);
nand UO_383 (O_383,N_29965,N_29509);
or UO_384 (O_384,N_29794,N_29571);
nand UO_385 (O_385,N_29509,N_29970);
nand UO_386 (O_386,N_29851,N_29578);
or UO_387 (O_387,N_29963,N_29703);
or UO_388 (O_388,N_29835,N_29560);
xnor UO_389 (O_389,N_29935,N_29876);
xnor UO_390 (O_390,N_29952,N_29753);
nor UO_391 (O_391,N_29998,N_29798);
xnor UO_392 (O_392,N_29911,N_29700);
or UO_393 (O_393,N_29761,N_29879);
xnor UO_394 (O_394,N_29836,N_29888);
nand UO_395 (O_395,N_29539,N_29600);
and UO_396 (O_396,N_29948,N_29510);
xor UO_397 (O_397,N_29688,N_29819);
nand UO_398 (O_398,N_29598,N_29982);
nand UO_399 (O_399,N_29652,N_29701);
or UO_400 (O_400,N_29707,N_29955);
nor UO_401 (O_401,N_29678,N_29966);
and UO_402 (O_402,N_29706,N_29687);
or UO_403 (O_403,N_29600,N_29728);
nand UO_404 (O_404,N_29990,N_29999);
nand UO_405 (O_405,N_29595,N_29631);
and UO_406 (O_406,N_29599,N_29741);
xnor UO_407 (O_407,N_29999,N_29770);
nand UO_408 (O_408,N_29814,N_29916);
nand UO_409 (O_409,N_29798,N_29607);
xor UO_410 (O_410,N_29804,N_29934);
xnor UO_411 (O_411,N_29942,N_29747);
or UO_412 (O_412,N_29610,N_29777);
or UO_413 (O_413,N_29910,N_29866);
xnor UO_414 (O_414,N_29756,N_29990);
xor UO_415 (O_415,N_29952,N_29797);
xor UO_416 (O_416,N_29986,N_29900);
and UO_417 (O_417,N_29759,N_29640);
nand UO_418 (O_418,N_29959,N_29509);
or UO_419 (O_419,N_29533,N_29868);
and UO_420 (O_420,N_29580,N_29539);
nand UO_421 (O_421,N_29577,N_29551);
and UO_422 (O_422,N_29857,N_29869);
and UO_423 (O_423,N_29683,N_29705);
nand UO_424 (O_424,N_29741,N_29773);
and UO_425 (O_425,N_29983,N_29836);
or UO_426 (O_426,N_29663,N_29869);
nor UO_427 (O_427,N_29702,N_29876);
or UO_428 (O_428,N_29956,N_29600);
nor UO_429 (O_429,N_29917,N_29601);
and UO_430 (O_430,N_29693,N_29928);
nor UO_431 (O_431,N_29971,N_29954);
nand UO_432 (O_432,N_29620,N_29633);
or UO_433 (O_433,N_29744,N_29580);
nand UO_434 (O_434,N_29512,N_29602);
xnor UO_435 (O_435,N_29692,N_29551);
xnor UO_436 (O_436,N_29983,N_29940);
or UO_437 (O_437,N_29996,N_29660);
and UO_438 (O_438,N_29652,N_29712);
and UO_439 (O_439,N_29987,N_29674);
and UO_440 (O_440,N_29774,N_29939);
xnor UO_441 (O_441,N_29726,N_29686);
nand UO_442 (O_442,N_29641,N_29890);
nor UO_443 (O_443,N_29938,N_29544);
and UO_444 (O_444,N_29945,N_29606);
or UO_445 (O_445,N_29517,N_29556);
or UO_446 (O_446,N_29536,N_29592);
and UO_447 (O_447,N_29879,N_29917);
and UO_448 (O_448,N_29924,N_29953);
and UO_449 (O_449,N_29796,N_29681);
and UO_450 (O_450,N_29528,N_29845);
nor UO_451 (O_451,N_29722,N_29667);
xnor UO_452 (O_452,N_29939,N_29517);
nor UO_453 (O_453,N_29825,N_29853);
or UO_454 (O_454,N_29649,N_29977);
and UO_455 (O_455,N_29921,N_29950);
and UO_456 (O_456,N_29716,N_29524);
xnor UO_457 (O_457,N_29500,N_29768);
or UO_458 (O_458,N_29799,N_29808);
xor UO_459 (O_459,N_29980,N_29504);
and UO_460 (O_460,N_29829,N_29704);
nor UO_461 (O_461,N_29663,N_29743);
or UO_462 (O_462,N_29753,N_29667);
and UO_463 (O_463,N_29671,N_29600);
nand UO_464 (O_464,N_29982,N_29795);
nor UO_465 (O_465,N_29723,N_29910);
and UO_466 (O_466,N_29973,N_29540);
nor UO_467 (O_467,N_29989,N_29672);
and UO_468 (O_468,N_29795,N_29677);
nand UO_469 (O_469,N_29778,N_29783);
and UO_470 (O_470,N_29870,N_29571);
nand UO_471 (O_471,N_29872,N_29894);
nor UO_472 (O_472,N_29942,N_29792);
and UO_473 (O_473,N_29840,N_29558);
or UO_474 (O_474,N_29916,N_29887);
and UO_475 (O_475,N_29969,N_29828);
nand UO_476 (O_476,N_29728,N_29817);
xor UO_477 (O_477,N_29740,N_29943);
or UO_478 (O_478,N_29508,N_29557);
and UO_479 (O_479,N_29759,N_29625);
xnor UO_480 (O_480,N_29571,N_29862);
or UO_481 (O_481,N_29504,N_29981);
or UO_482 (O_482,N_29807,N_29668);
or UO_483 (O_483,N_29515,N_29635);
and UO_484 (O_484,N_29737,N_29714);
nor UO_485 (O_485,N_29510,N_29667);
or UO_486 (O_486,N_29755,N_29632);
nor UO_487 (O_487,N_29665,N_29809);
xor UO_488 (O_488,N_29619,N_29559);
xnor UO_489 (O_489,N_29886,N_29505);
or UO_490 (O_490,N_29914,N_29676);
or UO_491 (O_491,N_29855,N_29838);
and UO_492 (O_492,N_29785,N_29962);
or UO_493 (O_493,N_29857,N_29590);
or UO_494 (O_494,N_29810,N_29588);
or UO_495 (O_495,N_29619,N_29665);
or UO_496 (O_496,N_29886,N_29975);
nand UO_497 (O_497,N_29697,N_29612);
nand UO_498 (O_498,N_29545,N_29515);
xor UO_499 (O_499,N_29661,N_29773);
and UO_500 (O_500,N_29527,N_29868);
or UO_501 (O_501,N_29571,N_29739);
and UO_502 (O_502,N_29529,N_29876);
nor UO_503 (O_503,N_29502,N_29767);
or UO_504 (O_504,N_29984,N_29800);
nor UO_505 (O_505,N_29521,N_29599);
nor UO_506 (O_506,N_29899,N_29895);
and UO_507 (O_507,N_29966,N_29975);
and UO_508 (O_508,N_29589,N_29631);
and UO_509 (O_509,N_29665,N_29864);
xnor UO_510 (O_510,N_29802,N_29610);
nand UO_511 (O_511,N_29767,N_29709);
nor UO_512 (O_512,N_29597,N_29666);
xor UO_513 (O_513,N_29822,N_29782);
xor UO_514 (O_514,N_29729,N_29661);
nand UO_515 (O_515,N_29952,N_29780);
and UO_516 (O_516,N_29948,N_29655);
xor UO_517 (O_517,N_29705,N_29811);
and UO_518 (O_518,N_29645,N_29665);
nand UO_519 (O_519,N_29963,N_29653);
nand UO_520 (O_520,N_29887,N_29567);
nand UO_521 (O_521,N_29924,N_29793);
nor UO_522 (O_522,N_29606,N_29645);
nand UO_523 (O_523,N_29761,N_29650);
or UO_524 (O_524,N_29969,N_29734);
nor UO_525 (O_525,N_29644,N_29841);
nand UO_526 (O_526,N_29571,N_29693);
nand UO_527 (O_527,N_29614,N_29960);
nor UO_528 (O_528,N_29501,N_29824);
xnor UO_529 (O_529,N_29749,N_29568);
nand UO_530 (O_530,N_29680,N_29738);
and UO_531 (O_531,N_29622,N_29936);
nand UO_532 (O_532,N_29768,N_29780);
xnor UO_533 (O_533,N_29947,N_29929);
or UO_534 (O_534,N_29801,N_29855);
nor UO_535 (O_535,N_29809,N_29938);
and UO_536 (O_536,N_29971,N_29901);
xor UO_537 (O_537,N_29604,N_29658);
or UO_538 (O_538,N_29855,N_29740);
or UO_539 (O_539,N_29716,N_29538);
and UO_540 (O_540,N_29830,N_29751);
nand UO_541 (O_541,N_29645,N_29556);
and UO_542 (O_542,N_29521,N_29505);
nor UO_543 (O_543,N_29899,N_29708);
or UO_544 (O_544,N_29936,N_29883);
nand UO_545 (O_545,N_29835,N_29683);
nand UO_546 (O_546,N_29804,N_29643);
and UO_547 (O_547,N_29790,N_29614);
xor UO_548 (O_548,N_29893,N_29954);
and UO_549 (O_549,N_29936,N_29869);
xor UO_550 (O_550,N_29505,N_29743);
nand UO_551 (O_551,N_29835,N_29601);
and UO_552 (O_552,N_29704,N_29659);
nand UO_553 (O_553,N_29619,N_29648);
and UO_554 (O_554,N_29538,N_29874);
nor UO_555 (O_555,N_29719,N_29904);
xnor UO_556 (O_556,N_29940,N_29923);
xnor UO_557 (O_557,N_29708,N_29874);
or UO_558 (O_558,N_29908,N_29804);
xor UO_559 (O_559,N_29892,N_29544);
nand UO_560 (O_560,N_29618,N_29730);
xor UO_561 (O_561,N_29628,N_29657);
nand UO_562 (O_562,N_29807,N_29880);
or UO_563 (O_563,N_29940,N_29795);
nand UO_564 (O_564,N_29876,N_29945);
nor UO_565 (O_565,N_29736,N_29579);
xnor UO_566 (O_566,N_29873,N_29877);
and UO_567 (O_567,N_29883,N_29614);
or UO_568 (O_568,N_29950,N_29801);
or UO_569 (O_569,N_29648,N_29584);
and UO_570 (O_570,N_29909,N_29990);
xnor UO_571 (O_571,N_29761,N_29579);
nand UO_572 (O_572,N_29859,N_29704);
nand UO_573 (O_573,N_29906,N_29669);
xnor UO_574 (O_574,N_29920,N_29700);
and UO_575 (O_575,N_29925,N_29546);
nand UO_576 (O_576,N_29707,N_29696);
and UO_577 (O_577,N_29751,N_29793);
or UO_578 (O_578,N_29963,N_29661);
and UO_579 (O_579,N_29578,N_29796);
or UO_580 (O_580,N_29895,N_29945);
xor UO_581 (O_581,N_29539,N_29568);
nor UO_582 (O_582,N_29631,N_29582);
nand UO_583 (O_583,N_29611,N_29522);
or UO_584 (O_584,N_29800,N_29994);
or UO_585 (O_585,N_29565,N_29699);
nand UO_586 (O_586,N_29784,N_29566);
xor UO_587 (O_587,N_29995,N_29676);
nor UO_588 (O_588,N_29978,N_29743);
nor UO_589 (O_589,N_29985,N_29618);
nor UO_590 (O_590,N_29652,N_29966);
nor UO_591 (O_591,N_29809,N_29811);
xor UO_592 (O_592,N_29943,N_29853);
and UO_593 (O_593,N_29594,N_29902);
xnor UO_594 (O_594,N_29697,N_29526);
or UO_595 (O_595,N_29511,N_29653);
nand UO_596 (O_596,N_29543,N_29786);
xnor UO_597 (O_597,N_29820,N_29923);
nand UO_598 (O_598,N_29860,N_29746);
or UO_599 (O_599,N_29896,N_29700);
nor UO_600 (O_600,N_29875,N_29602);
and UO_601 (O_601,N_29875,N_29501);
and UO_602 (O_602,N_29941,N_29547);
or UO_603 (O_603,N_29846,N_29962);
nor UO_604 (O_604,N_29961,N_29761);
nand UO_605 (O_605,N_29649,N_29535);
and UO_606 (O_606,N_29738,N_29554);
xnor UO_607 (O_607,N_29684,N_29693);
or UO_608 (O_608,N_29998,N_29855);
nand UO_609 (O_609,N_29975,N_29942);
and UO_610 (O_610,N_29879,N_29628);
or UO_611 (O_611,N_29737,N_29715);
nor UO_612 (O_612,N_29860,N_29801);
nor UO_613 (O_613,N_29634,N_29879);
and UO_614 (O_614,N_29524,N_29734);
nand UO_615 (O_615,N_29972,N_29607);
xnor UO_616 (O_616,N_29821,N_29757);
nand UO_617 (O_617,N_29553,N_29956);
and UO_618 (O_618,N_29853,N_29968);
and UO_619 (O_619,N_29657,N_29557);
and UO_620 (O_620,N_29562,N_29575);
nand UO_621 (O_621,N_29963,N_29722);
nor UO_622 (O_622,N_29581,N_29598);
nor UO_623 (O_623,N_29828,N_29986);
and UO_624 (O_624,N_29804,N_29969);
and UO_625 (O_625,N_29985,N_29582);
xor UO_626 (O_626,N_29980,N_29868);
and UO_627 (O_627,N_29977,N_29933);
and UO_628 (O_628,N_29611,N_29903);
or UO_629 (O_629,N_29868,N_29975);
xor UO_630 (O_630,N_29748,N_29529);
or UO_631 (O_631,N_29559,N_29517);
and UO_632 (O_632,N_29951,N_29833);
nand UO_633 (O_633,N_29567,N_29689);
and UO_634 (O_634,N_29502,N_29953);
or UO_635 (O_635,N_29985,N_29962);
and UO_636 (O_636,N_29676,N_29820);
nor UO_637 (O_637,N_29851,N_29904);
nand UO_638 (O_638,N_29959,N_29876);
xor UO_639 (O_639,N_29797,N_29687);
xnor UO_640 (O_640,N_29521,N_29957);
nand UO_641 (O_641,N_29547,N_29608);
or UO_642 (O_642,N_29696,N_29548);
xor UO_643 (O_643,N_29846,N_29658);
xnor UO_644 (O_644,N_29721,N_29676);
nand UO_645 (O_645,N_29695,N_29680);
nor UO_646 (O_646,N_29634,N_29593);
nor UO_647 (O_647,N_29861,N_29929);
nor UO_648 (O_648,N_29865,N_29777);
nor UO_649 (O_649,N_29684,N_29772);
nand UO_650 (O_650,N_29628,N_29687);
xnor UO_651 (O_651,N_29937,N_29522);
nand UO_652 (O_652,N_29630,N_29801);
nor UO_653 (O_653,N_29923,N_29681);
nor UO_654 (O_654,N_29582,N_29646);
or UO_655 (O_655,N_29978,N_29864);
nor UO_656 (O_656,N_29950,N_29749);
xnor UO_657 (O_657,N_29553,N_29755);
nor UO_658 (O_658,N_29571,N_29940);
xor UO_659 (O_659,N_29952,N_29577);
and UO_660 (O_660,N_29838,N_29641);
or UO_661 (O_661,N_29902,N_29713);
xor UO_662 (O_662,N_29821,N_29572);
xor UO_663 (O_663,N_29513,N_29701);
nand UO_664 (O_664,N_29770,N_29669);
and UO_665 (O_665,N_29527,N_29891);
nand UO_666 (O_666,N_29582,N_29887);
xor UO_667 (O_667,N_29513,N_29674);
and UO_668 (O_668,N_29516,N_29843);
xor UO_669 (O_669,N_29969,N_29550);
nor UO_670 (O_670,N_29545,N_29594);
nor UO_671 (O_671,N_29733,N_29842);
or UO_672 (O_672,N_29759,N_29537);
xor UO_673 (O_673,N_29908,N_29915);
nand UO_674 (O_674,N_29817,N_29671);
or UO_675 (O_675,N_29781,N_29668);
nor UO_676 (O_676,N_29974,N_29524);
xnor UO_677 (O_677,N_29922,N_29983);
xnor UO_678 (O_678,N_29947,N_29510);
nand UO_679 (O_679,N_29543,N_29661);
and UO_680 (O_680,N_29621,N_29648);
xnor UO_681 (O_681,N_29817,N_29768);
and UO_682 (O_682,N_29819,N_29545);
xnor UO_683 (O_683,N_29826,N_29816);
xnor UO_684 (O_684,N_29820,N_29534);
and UO_685 (O_685,N_29629,N_29536);
and UO_686 (O_686,N_29663,N_29946);
or UO_687 (O_687,N_29594,N_29966);
nor UO_688 (O_688,N_29923,N_29585);
nor UO_689 (O_689,N_29956,N_29546);
or UO_690 (O_690,N_29909,N_29632);
or UO_691 (O_691,N_29990,N_29571);
xor UO_692 (O_692,N_29610,N_29575);
xor UO_693 (O_693,N_29836,N_29976);
and UO_694 (O_694,N_29953,N_29699);
and UO_695 (O_695,N_29710,N_29665);
or UO_696 (O_696,N_29581,N_29667);
and UO_697 (O_697,N_29527,N_29979);
nand UO_698 (O_698,N_29634,N_29937);
and UO_699 (O_699,N_29550,N_29617);
nand UO_700 (O_700,N_29960,N_29610);
nor UO_701 (O_701,N_29773,N_29552);
nor UO_702 (O_702,N_29780,N_29688);
nor UO_703 (O_703,N_29776,N_29713);
nand UO_704 (O_704,N_29820,N_29693);
nand UO_705 (O_705,N_29952,N_29874);
xor UO_706 (O_706,N_29798,N_29588);
nor UO_707 (O_707,N_29850,N_29836);
xor UO_708 (O_708,N_29655,N_29977);
or UO_709 (O_709,N_29591,N_29567);
or UO_710 (O_710,N_29576,N_29824);
or UO_711 (O_711,N_29706,N_29982);
xor UO_712 (O_712,N_29869,N_29952);
nand UO_713 (O_713,N_29561,N_29647);
and UO_714 (O_714,N_29812,N_29763);
or UO_715 (O_715,N_29988,N_29554);
and UO_716 (O_716,N_29857,N_29714);
and UO_717 (O_717,N_29950,N_29879);
nand UO_718 (O_718,N_29516,N_29796);
nand UO_719 (O_719,N_29535,N_29871);
nand UO_720 (O_720,N_29526,N_29684);
or UO_721 (O_721,N_29614,N_29897);
and UO_722 (O_722,N_29591,N_29671);
nor UO_723 (O_723,N_29648,N_29597);
and UO_724 (O_724,N_29589,N_29683);
nand UO_725 (O_725,N_29896,N_29689);
or UO_726 (O_726,N_29882,N_29972);
nor UO_727 (O_727,N_29857,N_29758);
nand UO_728 (O_728,N_29755,N_29532);
or UO_729 (O_729,N_29783,N_29775);
nand UO_730 (O_730,N_29774,N_29899);
nor UO_731 (O_731,N_29840,N_29874);
nor UO_732 (O_732,N_29767,N_29845);
nor UO_733 (O_733,N_29973,N_29700);
or UO_734 (O_734,N_29586,N_29597);
nand UO_735 (O_735,N_29932,N_29625);
or UO_736 (O_736,N_29957,N_29612);
nand UO_737 (O_737,N_29947,N_29761);
nor UO_738 (O_738,N_29866,N_29843);
nor UO_739 (O_739,N_29907,N_29827);
or UO_740 (O_740,N_29928,N_29962);
nor UO_741 (O_741,N_29804,N_29684);
xnor UO_742 (O_742,N_29501,N_29504);
or UO_743 (O_743,N_29521,N_29836);
nor UO_744 (O_744,N_29682,N_29674);
xnor UO_745 (O_745,N_29870,N_29662);
and UO_746 (O_746,N_29953,N_29604);
or UO_747 (O_747,N_29904,N_29947);
xnor UO_748 (O_748,N_29951,N_29947);
nor UO_749 (O_749,N_29708,N_29665);
and UO_750 (O_750,N_29996,N_29580);
nor UO_751 (O_751,N_29902,N_29812);
nor UO_752 (O_752,N_29673,N_29630);
xor UO_753 (O_753,N_29658,N_29951);
or UO_754 (O_754,N_29939,N_29974);
xnor UO_755 (O_755,N_29588,N_29534);
nand UO_756 (O_756,N_29933,N_29596);
xor UO_757 (O_757,N_29619,N_29613);
nand UO_758 (O_758,N_29516,N_29560);
xor UO_759 (O_759,N_29883,N_29811);
nor UO_760 (O_760,N_29539,N_29938);
or UO_761 (O_761,N_29546,N_29563);
or UO_762 (O_762,N_29538,N_29906);
nand UO_763 (O_763,N_29668,N_29869);
or UO_764 (O_764,N_29863,N_29996);
nand UO_765 (O_765,N_29928,N_29771);
xnor UO_766 (O_766,N_29605,N_29933);
nor UO_767 (O_767,N_29513,N_29733);
xnor UO_768 (O_768,N_29902,N_29726);
or UO_769 (O_769,N_29853,N_29937);
or UO_770 (O_770,N_29516,N_29901);
nor UO_771 (O_771,N_29500,N_29831);
nand UO_772 (O_772,N_29864,N_29780);
xor UO_773 (O_773,N_29523,N_29741);
nor UO_774 (O_774,N_29925,N_29540);
and UO_775 (O_775,N_29906,N_29796);
nand UO_776 (O_776,N_29861,N_29650);
or UO_777 (O_777,N_29537,N_29560);
xor UO_778 (O_778,N_29906,N_29843);
xnor UO_779 (O_779,N_29711,N_29740);
or UO_780 (O_780,N_29942,N_29765);
xnor UO_781 (O_781,N_29712,N_29803);
nor UO_782 (O_782,N_29534,N_29639);
nand UO_783 (O_783,N_29623,N_29596);
nand UO_784 (O_784,N_29531,N_29899);
xnor UO_785 (O_785,N_29547,N_29537);
xor UO_786 (O_786,N_29773,N_29780);
nor UO_787 (O_787,N_29688,N_29929);
xor UO_788 (O_788,N_29946,N_29928);
nand UO_789 (O_789,N_29752,N_29888);
nor UO_790 (O_790,N_29827,N_29918);
nor UO_791 (O_791,N_29584,N_29632);
or UO_792 (O_792,N_29825,N_29900);
nand UO_793 (O_793,N_29733,N_29765);
nand UO_794 (O_794,N_29950,N_29892);
and UO_795 (O_795,N_29679,N_29674);
and UO_796 (O_796,N_29973,N_29861);
nand UO_797 (O_797,N_29535,N_29882);
nor UO_798 (O_798,N_29550,N_29612);
and UO_799 (O_799,N_29807,N_29868);
xor UO_800 (O_800,N_29509,N_29785);
or UO_801 (O_801,N_29936,N_29706);
xnor UO_802 (O_802,N_29571,N_29737);
xnor UO_803 (O_803,N_29917,N_29685);
and UO_804 (O_804,N_29985,N_29802);
nand UO_805 (O_805,N_29618,N_29694);
nand UO_806 (O_806,N_29946,N_29818);
nor UO_807 (O_807,N_29726,N_29587);
nor UO_808 (O_808,N_29561,N_29901);
or UO_809 (O_809,N_29914,N_29752);
nor UO_810 (O_810,N_29886,N_29990);
nand UO_811 (O_811,N_29517,N_29789);
nor UO_812 (O_812,N_29533,N_29565);
and UO_813 (O_813,N_29982,N_29793);
xor UO_814 (O_814,N_29883,N_29738);
or UO_815 (O_815,N_29609,N_29851);
nand UO_816 (O_816,N_29704,N_29746);
and UO_817 (O_817,N_29832,N_29760);
and UO_818 (O_818,N_29503,N_29773);
or UO_819 (O_819,N_29563,N_29679);
nor UO_820 (O_820,N_29690,N_29517);
nand UO_821 (O_821,N_29985,N_29772);
nor UO_822 (O_822,N_29684,N_29638);
or UO_823 (O_823,N_29720,N_29772);
or UO_824 (O_824,N_29642,N_29711);
xor UO_825 (O_825,N_29841,N_29748);
nor UO_826 (O_826,N_29968,N_29523);
xnor UO_827 (O_827,N_29582,N_29808);
and UO_828 (O_828,N_29912,N_29724);
nand UO_829 (O_829,N_29629,N_29606);
nand UO_830 (O_830,N_29554,N_29656);
xnor UO_831 (O_831,N_29707,N_29746);
nand UO_832 (O_832,N_29677,N_29778);
or UO_833 (O_833,N_29834,N_29690);
xnor UO_834 (O_834,N_29542,N_29772);
nor UO_835 (O_835,N_29689,N_29571);
xnor UO_836 (O_836,N_29717,N_29861);
and UO_837 (O_837,N_29765,N_29652);
xnor UO_838 (O_838,N_29588,N_29690);
or UO_839 (O_839,N_29751,N_29501);
xor UO_840 (O_840,N_29801,N_29636);
and UO_841 (O_841,N_29864,N_29670);
nor UO_842 (O_842,N_29681,N_29891);
xor UO_843 (O_843,N_29968,N_29534);
xor UO_844 (O_844,N_29840,N_29640);
nand UO_845 (O_845,N_29941,N_29866);
nand UO_846 (O_846,N_29631,N_29856);
nor UO_847 (O_847,N_29986,N_29798);
nand UO_848 (O_848,N_29868,N_29987);
or UO_849 (O_849,N_29990,N_29962);
nand UO_850 (O_850,N_29550,N_29880);
or UO_851 (O_851,N_29931,N_29690);
or UO_852 (O_852,N_29684,N_29903);
and UO_853 (O_853,N_29787,N_29784);
and UO_854 (O_854,N_29790,N_29675);
nand UO_855 (O_855,N_29846,N_29806);
xnor UO_856 (O_856,N_29621,N_29587);
and UO_857 (O_857,N_29714,N_29745);
nand UO_858 (O_858,N_29524,N_29689);
and UO_859 (O_859,N_29872,N_29711);
and UO_860 (O_860,N_29798,N_29580);
and UO_861 (O_861,N_29605,N_29587);
nand UO_862 (O_862,N_29750,N_29697);
nor UO_863 (O_863,N_29961,N_29637);
xor UO_864 (O_864,N_29803,N_29806);
nor UO_865 (O_865,N_29960,N_29832);
xor UO_866 (O_866,N_29909,N_29847);
xnor UO_867 (O_867,N_29764,N_29610);
xor UO_868 (O_868,N_29940,N_29987);
xnor UO_869 (O_869,N_29803,N_29779);
nand UO_870 (O_870,N_29668,N_29851);
nand UO_871 (O_871,N_29547,N_29659);
nor UO_872 (O_872,N_29718,N_29531);
or UO_873 (O_873,N_29941,N_29791);
nor UO_874 (O_874,N_29703,N_29674);
and UO_875 (O_875,N_29939,N_29634);
nor UO_876 (O_876,N_29736,N_29811);
nand UO_877 (O_877,N_29667,N_29742);
or UO_878 (O_878,N_29890,N_29683);
nand UO_879 (O_879,N_29626,N_29833);
or UO_880 (O_880,N_29608,N_29974);
and UO_881 (O_881,N_29573,N_29847);
xor UO_882 (O_882,N_29647,N_29780);
or UO_883 (O_883,N_29749,N_29843);
or UO_884 (O_884,N_29535,N_29988);
or UO_885 (O_885,N_29994,N_29566);
nand UO_886 (O_886,N_29703,N_29917);
and UO_887 (O_887,N_29868,N_29804);
or UO_888 (O_888,N_29687,N_29982);
xor UO_889 (O_889,N_29990,N_29685);
nor UO_890 (O_890,N_29990,N_29919);
or UO_891 (O_891,N_29688,N_29911);
or UO_892 (O_892,N_29657,N_29659);
and UO_893 (O_893,N_29814,N_29705);
xnor UO_894 (O_894,N_29652,N_29790);
nand UO_895 (O_895,N_29890,N_29933);
xnor UO_896 (O_896,N_29928,N_29923);
xnor UO_897 (O_897,N_29630,N_29623);
or UO_898 (O_898,N_29795,N_29914);
nor UO_899 (O_899,N_29590,N_29868);
and UO_900 (O_900,N_29820,N_29548);
xor UO_901 (O_901,N_29833,N_29915);
or UO_902 (O_902,N_29894,N_29774);
nor UO_903 (O_903,N_29691,N_29887);
or UO_904 (O_904,N_29523,N_29889);
and UO_905 (O_905,N_29621,N_29726);
nand UO_906 (O_906,N_29704,N_29821);
nand UO_907 (O_907,N_29898,N_29990);
nor UO_908 (O_908,N_29841,N_29658);
xor UO_909 (O_909,N_29553,N_29552);
or UO_910 (O_910,N_29693,N_29912);
or UO_911 (O_911,N_29983,N_29581);
nand UO_912 (O_912,N_29654,N_29835);
xor UO_913 (O_913,N_29579,N_29964);
xnor UO_914 (O_914,N_29756,N_29556);
or UO_915 (O_915,N_29690,N_29543);
nand UO_916 (O_916,N_29934,N_29984);
and UO_917 (O_917,N_29973,N_29560);
or UO_918 (O_918,N_29844,N_29611);
and UO_919 (O_919,N_29580,N_29960);
nand UO_920 (O_920,N_29934,N_29684);
or UO_921 (O_921,N_29833,N_29566);
nor UO_922 (O_922,N_29584,N_29929);
nor UO_923 (O_923,N_29600,N_29578);
xor UO_924 (O_924,N_29971,N_29705);
xor UO_925 (O_925,N_29639,N_29936);
or UO_926 (O_926,N_29584,N_29661);
nand UO_927 (O_927,N_29923,N_29595);
nand UO_928 (O_928,N_29746,N_29758);
nor UO_929 (O_929,N_29753,N_29711);
xor UO_930 (O_930,N_29602,N_29891);
nor UO_931 (O_931,N_29914,N_29796);
xor UO_932 (O_932,N_29943,N_29677);
nor UO_933 (O_933,N_29712,N_29954);
or UO_934 (O_934,N_29910,N_29735);
nor UO_935 (O_935,N_29560,N_29773);
or UO_936 (O_936,N_29897,N_29999);
nand UO_937 (O_937,N_29907,N_29839);
nand UO_938 (O_938,N_29621,N_29965);
nand UO_939 (O_939,N_29903,N_29802);
nand UO_940 (O_940,N_29842,N_29520);
nor UO_941 (O_941,N_29685,N_29821);
xor UO_942 (O_942,N_29717,N_29737);
nor UO_943 (O_943,N_29813,N_29899);
nor UO_944 (O_944,N_29702,N_29651);
nand UO_945 (O_945,N_29644,N_29763);
nor UO_946 (O_946,N_29975,N_29835);
or UO_947 (O_947,N_29604,N_29552);
xnor UO_948 (O_948,N_29967,N_29757);
and UO_949 (O_949,N_29547,N_29994);
xor UO_950 (O_950,N_29875,N_29917);
and UO_951 (O_951,N_29939,N_29941);
nor UO_952 (O_952,N_29892,N_29696);
or UO_953 (O_953,N_29995,N_29925);
or UO_954 (O_954,N_29569,N_29527);
or UO_955 (O_955,N_29720,N_29625);
xnor UO_956 (O_956,N_29627,N_29646);
xnor UO_957 (O_957,N_29975,N_29742);
or UO_958 (O_958,N_29578,N_29619);
xnor UO_959 (O_959,N_29981,N_29985);
xnor UO_960 (O_960,N_29849,N_29524);
or UO_961 (O_961,N_29639,N_29864);
and UO_962 (O_962,N_29612,N_29692);
nand UO_963 (O_963,N_29759,N_29539);
or UO_964 (O_964,N_29788,N_29594);
nand UO_965 (O_965,N_29970,N_29751);
nor UO_966 (O_966,N_29948,N_29809);
nand UO_967 (O_967,N_29799,N_29939);
or UO_968 (O_968,N_29694,N_29645);
xnor UO_969 (O_969,N_29978,N_29995);
xor UO_970 (O_970,N_29573,N_29531);
xnor UO_971 (O_971,N_29775,N_29878);
nor UO_972 (O_972,N_29931,N_29906);
or UO_973 (O_973,N_29686,N_29581);
xor UO_974 (O_974,N_29768,N_29519);
or UO_975 (O_975,N_29780,N_29500);
or UO_976 (O_976,N_29968,N_29810);
and UO_977 (O_977,N_29980,N_29942);
or UO_978 (O_978,N_29820,N_29857);
and UO_979 (O_979,N_29717,N_29960);
nand UO_980 (O_980,N_29616,N_29889);
nor UO_981 (O_981,N_29556,N_29886);
and UO_982 (O_982,N_29715,N_29516);
or UO_983 (O_983,N_29879,N_29682);
and UO_984 (O_984,N_29880,N_29842);
or UO_985 (O_985,N_29678,N_29759);
or UO_986 (O_986,N_29912,N_29536);
nor UO_987 (O_987,N_29882,N_29824);
and UO_988 (O_988,N_29835,N_29644);
or UO_989 (O_989,N_29561,N_29895);
nand UO_990 (O_990,N_29650,N_29796);
nand UO_991 (O_991,N_29551,N_29922);
or UO_992 (O_992,N_29762,N_29750);
xor UO_993 (O_993,N_29980,N_29649);
xnor UO_994 (O_994,N_29945,N_29523);
and UO_995 (O_995,N_29883,N_29707);
xnor UO_996 (O_996,N_29967,N_29772);
nand UO_997 (O_997,N_29623,N_29894);
or UO_998 (O_998,N_29845,N_29860);
nor UO_999 (O_999,N_29910,N_29937);
xnor UO_1000 (O_1000,N_29809,N_29917);
nand UO_1001 (O_1001,N_29708,N_29683);
and UO_1002 (O_1002,N_29506,N_29582);
xor UO_1003 (O_1003,N_29551,N_29531);
nand UO_1004 (O_1004,N_29905,N_29718);
and UO_1005 (O_1005,N_29846,N_29754);
nor UO_1006 (O_1006,N_29979,N_29627);
nand UO_1007 (O_1007,N_29661,N_29967);
nand UO_1008 (O_1008,N_29778,N_29628);
and UO_1009 (O_1009,N_29979,N_29555);
nor UO_1010 (O_1010,N_29675,N_29695);
xor UO_1011 (O_1011,N_29793,N_29958);
and UO_1012 (O_1012,N_29849,N_29804);
nor UO_1013 (O_1013,N_29554,N_29575);
or UO_1014 (O_1014,N_29798,N_29538);
nand UO_1015 (O_1015,N_29765,N_29893);
nor UO_1016 (O_1016,N_29701,N_29817);
or UO_1017 (O_1017,N_29606,N_29627);
or UO_1018 (O_1018,N_29846,N_29515);
and UO_1019 (O_1019,N_29864,N_29601);
nand UO_1020 (O_1020,N_29617,N_29782);
nor UO_1021 (O_1021,N_29573,N_29578);
nor UO_1022 (O_1022,N_29785,N_29748);
nand UO_1023 (O_1023,N_29978,N_29575);
nor UO_1024 (O_1024,N_29536,N_29620);
xor UO_1025 (O_1025,N_29579,N_29925);
nand UO_1026 (O_1026,N_29778,N_29799);
xor UO_1027 (O_1027,N_29984,N_29786);
xor UO_1028 (O_1028,N_29969,N_29557);
or UO_1029 (O_1029,N_29640,N_29934);
nand UO_1030 (O_1030,N_29724,N_29767);
and UO_1031 (O_1031,N_29752,N_29638);
xor UO_1032 (O_1032,N_29916,N_29845);
nand UO_1033 (O_1033,N_29675,N_29558);
nor UO_1034 (O_1034,N_29875,N_29564);
or UO_1035 (O_1035,N_29912,N_29930);
and UO_1036 (O_1036,N_29977,N_29823);
xor UO_1037 (O_1037,N_29991,N_29722);
xor UO_1038 (O_1038,N_29846,N_29948);
nor UO_1039 (O_1039,N_29680,N_29664);
xnor UO_1040 (O_1040,N_29920,N_29515);
or UO_1041 (O_1041,N_29654,N_29559);
and UO_1042 (O_1042,N_29814,N_29778);
nand UO_1043 (O_1043,N_29597,N_29717);
or UO_1044 (O_1044,N_29939,N_29958);
or UO_1045 (O_1045,N_29995,N_29538);
nand UO_1046 (O_1046,N_29851,N_29605);
nand UO_1047 (O_1047,N_29606,N_29673);
nand UO_1048 (O_1048,N_29651,N_29787);
nor UO_1049 (O_1049,N_29665,N_29813);
or UO_1050 (O_1050,N_29751,N_29790);
or UO_1051 (O_1051,N_29563,N_29503);
nand UO_1052 (O_1052,N_29540,N_29791);
nand UO_1053 (O_1053,N_29658,N_29784);
xor UO_1054 (O_1054,N_29818,N_29926);
nand UO_1055 (O_1055,N_29917,N_29926);
or UO_1056 (O_1056,N_29981,N_29513);
and UO_1057 (O_1057,N_29836,N_29501);
xor UO_1058 (O_1058,N_29983,N_29653);
and UO_1059 (O_1059,N_29678,N_29732);
nand UO_1060 (O_1060,N_29935,N_29711);
or UO_1061 (O_1061,N_29732,N_29870);
nor UO_1062 (O_1062,N_29713,N_29792);
nand UO_1063 (O_1063,N_29862,N_29921);
xor UO_1064 (O_1064,N_29924,N_29702);
nand UO_1065 (O_1065,N_29761,N_29571);
or UO_1066 (O_1066,N_29820,N_29513);
and UO_1067 (O_1067,N_29714,N_29899);
or UO_1068 (O_1068,N_29502,N_29895);
or UO_1069 (O_1069,N_29749,N_29814);
and UO_1070 (O_1070,N_29800,N_29607);
nor UO_1071 (O_1071,N_29983,N_29744);
nand UO_1072 (O_1072,N_29967,N_29857);
or UO_1073 (O_1073,N_29878,N_29647);
nor UO_1074 (O_1074,N_29923,N_29658);
or UO_1075 (O_1075,N_29504,N_29564);
nand UO_1076 (O_1076,N_29895,N_29907);
and UO_1077 (O_1077,N_29557,N_29528);
xnor UO_1078 (O_1078,N_29541,N_29562);
nand UO_1079 (O_1079,N_29826,N_29512);
nand UO_1080 (O_1080,N_29687,N_29815);
nor UO_1081 (O_1081,N_29932,N_29623);
nor UO_1082 (O_1082,N_29946,N_29586);
nand UO_1083 (O_1083,N_29832,N_29999);
and UO_1084 (O_1084,N_29724,N_29909);
nor UO_1085 (O_1085,N_29839,N_29859);
xnor UO_1086 (O_1086,N_29897,N_29512);
xnor UO_1087 (O_1087,N_29713,N_29613);
nor UO_1088 (O_1088,N_29613,N_29593);
nor UO_1089 (O_1089,N_29792,N_29523);
nand UO_1090 (O_1090,N_29533,N_29679);
nand UO_1091 (O_1091,N_29873,N_29760);
nor UO_1092 (O_1092,N_29889,N_29702);
nor UO_1093 (O_1093,N_29528,N_29853);
xnor UO_1094 (O_1094,N_29896,N_29929);
nor UO_1095 (O_1095,N_29723,N_29717);
xnor UO_1096 (O_1096,N_29953,N_29866);
nor UO_1097 (O_1097,N_29776,N_29849);
or UO_1098 (O_1098,N_29717,N_29871);
and UO_1099 (O_1099,N_29708,N_29631);
and UO_1100 (O_1100,N_29806,N_29575);
xnor UO_1101 (O_1101,N_29507,N_29635);
xor UO_1102 (O_1102,N_29590,N_29565);
nor UO_1103 (O_1103,N_29869,N_29629);
nor UO_1104 (O_1104,N_29952,N_29768);
xor UO_1105 (O_1105,N_29993,N_29637);
nand UO_1106 (O_1106,N_29975,N_29789);
xor UO_1107 (O_1107,N_29725,N_29906);
nand UO_1108 (O_1108,N_29821,N_29872);
or UO_1109 (O_1109,N_29712,N_29548);
and UO_1110 (O_1110,N_29641,N_29675);
xnor UO_1111 (O_1111,N_29521,N_29937);
nand UO_1112 (O_1112,N_29917,N_29737);
xor UO_1113 (O_1113,N_29722,N_29651);
and UO_1114 (O_1114,N_29524,N_29786);
nor UO_1115 (O_1115,N_29815,N_29683);
and UO_1116 (O_1116,N_29789,N_29620);
nand UO_1117 (O_1117,N_29635,N_29987);
or UO_1118 (O_1118,N_29961,N_29901);
or UO_1119 (O_1119,N_29752,N_29791);
xor UO_1120 (O_1120,N_29830,N_29813);
or UO_1121 (O_1121,N_29523,N_29852);
nand UO_1122 (O_1122,N_29524,N_29730);
nand UO_1123 (O_1123,N_29599,N_29602);
nand UO_1124 (O_1124,N_29704,N_29631);
nor UO_1125 (O_1125,N_29726,N_29970);
xnor UO_1126 (O_1126,N_29646,N_29958);
or UO_1127 (O_1127,N_29805,N_29606);
xor UO_1128 (O_1128,N_29660,N_29656);
and UO_1129 (O_1129,N_29913,N_29741);
nor UO_1130 (O_1130,N_29760,N_29862);
xor UO_1131 (O_1131,N_29701,N_29635);
nor UO_1132 (O_1132,N_29559,N_29920);
nand UO_1133 (O_1133,N_29586,N_29702);
nor UO_1134 (O_1134,N_29746,N_29987);
nand UO_1135 (O_1135,N_29551,N_29877);
or UO_1136 (O_1136,N_29699,N_29583);
and UO_1137 (O_1137,N_29543,N_29686);
xor UO_1138 (O_1138,N_29667,N_29794);
nand UO_1139 (O_1139,N_29805,N_29721);
nand UO_1140 (O_1140,N_29835,N_29522);
or UO_1141 (O_1141,N_29982,N_29691);
nand UO_1142 (O_1142,N_29519,N_29850);
and UO_1143 (O_1143,N_29654,N_29763);
nor UO_1144 (O_1144,N_29578,N_29892);
nand UO_1145 (O_1145,N_29865,N_29846);
nand UO_1146 (O_1146,N_29898,N_29770);
nand UO_1147 (O_1147,N_29785,N_29697);
and UO_1148 (O_1148,N_29819,N_29581);
xnor UO_1149 (O_1149,N_29954,N_29700);
or UO_1150 (O_1150,N_29745,N_29639);
and UO_1151 (O_1151,N_29861,N_29939);
nor UO_1152 (O_1152,N_29777,N_29826);
or UO_1153 (O_1153,N_29525,N_29638);
or UO_1154 (O_1154,N_29565,N_29783);
and UO_1155 (O_1155,N_29868,N_29720);
nand UO_1156 (O_1156,N_29927,N_29866);
or UO_1157 (O_1157,N_29937,N_29729);
nor UO_1158 (O_1158,N_29837,N_29789);
and UO_1159 (O_1159,N_29883,N_29708);
nand UO_1160 (O_1160,N_29560,N_29660);
xor UO_1161 (O_1161,N_29901,N_29976);
nor UO_1162 (O_1162,N_29885,N_29637);
nand UO_1163 (O_1163,N_29529,N_29943);
xnor UO_1164 (O_1164,N_29701,N_29997);
xor UO_1165 (O_1165,N_29794,N_29960);
nor UO_1166 (O_1166,N_29692,N_29624);
xor UO_1167 (O_1167,N_29932,N_29887);
or UO_1168 (O_1168,N_29873,N_29854);
xor UO_1169 (O_1169,N_29872,N_29653);
and UO_1170 (O_1170,N_29731,N_29547);
or UO_1171 (O_1171,N_29587,N_29790);
nor UO_1172 (O_1172,N_29517,N_29943);
and UO_1173 (O_1173,N_29783,N_29725);
or UO_1174 (O_1174,N_29514,N_29577);
and UO_1175 (O_1175,N_29905,N_29638);
or UO_1176 (O_1176,N_29892,N_29758);
nand UO_1177 (O_1177,N_29974,N_29792);
nor UO_1178 (O_1178,N_29542,N_29781);
nand UO_1179 (O_1179,N_29724,N_29984);
and UO_1180 (O_1180,N_29540,N_29659);
nor UO_1181 (O_1181,N_29533,N_29905);
nand UO_1182 (O_1182,N_29793,N_29523);
nor UO_1183 (O_1183,N_29864,N_29668);
or UO_1184 (O_1184,N_29727,N_29611);
xnor UO_1185 (O_1185,N_29985,N_29834);
and UO_1186 (O_1186,N_29709,N_29857);
xor UO_1187 (O_1187,N_29648,N_29755);
nand UO_1188 (O_1188,N_29922,N_29732);
nor UO_1189 (O_1189,N_29521,N_29681);
or UO_1190 (O_1190,N_29799,N_29575);
and UO_1191 (O_1191,N_29966,N_29974);
xnor UO_1192 (O_1192,N_29757,N_29922);
xnor UO_1193 (O_1193,N_29846,N_29668);
nand UO_1194 (O_1194,N_29782,N_29749);
xor UO_1195 (O_1195,N_29840,N_29990);
nor UO_1196 (O_1196,N_29660,N_29970);
and UO_1197 (O_1197,N_29781,N_29707);
nand UO_1198 (O_1198,N_29657,N_29966);
or UO_1199 (O_1199,N_29756,N_29667);
nand UO_1200 (O_1200,N_29878,N_29799);
or UO_1201 (O_1201,N_29801,N_29936);
and UO_1202 (O_1202,N_29599,N_29549);
nand UO_1203 (O_1203,N_29604,N_29887);
nor UO_1204 (O_1204,N_29759,N_29819);
nor UO_1205 (O_1205,N_29891,N_29760);
xnor UO_1206 (O_1206,N_29700,N_29656);
nand UO_1207 (O_1207,N_29617,N_29983);
xnor UO_1208 (O_1208,N_29575,N_29706);
nand UO_1209 (O_1209,N_29787,N_29734);
nand UO_1210 (O_1210,N_29842,N_29525);
and UO_1211 (O_1211,N_29518,N_29743);
xor UO_1212 (O_1212,N_29575,N_29680);
or UO_1213 (O_1213,N_29941,N_29761);
nand UO_1214 (O_1214,N_29787,N_29856);
or UO_1215 (O_1215,N_29654,N_29774);
xor UO_1216 (O_1216,N_29557,N_29906);
and UO_1217 (O_1217,N_29891,N_29616);
or UO_1218 (O_1218,N_29763,N_29597);
xnor UO_1219 (O_1219,N_29722,N_29894);
nor UO_1220 (O_1220,N_29609,N_29933);
nor UO_1221 (O_1221,N_29596,N_29982);
nor UO_1222 (O_1222,N_29663,N_29591);
nand UO_1223 (O_1223,N_29694,N_29934);
nor UO_1224 (O_1224,N_29662,N_29964);
xnor UO_1225 (O_1225,N_29991,N_29684);
or UO_1226 (O_1226,N_29523,N_29547);
nand UO_1227 (O_1227,N_29523,N_29538);
and UO_1228 (O_1228,N_29837,N_29530);
and UO_1229 (O_1229,N_29663,N_29805);
nand UO_1230 (O_1230,N_29978,N_29704);
and UO_1231 (O_1231,N_29506,N_29551);
and UO_1232 (O_1232,N_29516,N_29780);
or UO_1233 (O_1233,N_29939,N_29622);
or UO_1234 (O_1234,N_29977,N_29999);
xor UO_1235 (O_1235,N_29999,N_29659);
nand UO_1236 (O_1236,N_29726,N_29534);
nand UO_1237 (O_1237,N_29808,N_29958);
nor UO_1238 (O_1238,N_29708,N_29950);
and UO_1239 (O_1239,N_29819,N_29973);
and UO_1240 (O_1240,N_29707,N_29911);
xor UO_1241 (O_1241,N_29597,N_29521);
nor UO_1242 (O_1242,N_29704,N_29764);
and UO_1243 (O_1243,N_29996,N_29975);
xnor UO_1244 (O_1244,N_29870,N_29700);
xnor UO_1245 (O_1245,N_29503,N_29629);
nand UO_1246 (O_1246,N_29524,N_29810);
and UO_1247 (O_1247,N_29591,N_29510);
nor UO_1248 (O_1248,N_29894,N_29912);
and UO_1249 (O_1249,N_29792,N_29916);
and UO_1250 (O_1250,N_29634,N_29915);
and UO_1251 (O_1251,N_29899,N_29509);
nand UO_1252 (O_1252,N_29953,N_29865);
nand UO_1253 (O_1253,N_29862,N_29889);
and UO_1254 (O_1254,N_29579,N_29591);
nand UO_1255 (O_1255,N_29510,N_29767);
nor UO_1256 (O_1256,N_29717,N_29505);
nand UO_1257 (O_1257,N_29948,N_29824);
xnor UO_1258 (O_1258,N_29724,N_29606);
and UO_1259 (O_1259,N_29672,N_29940);
nand UO_1260 (O_1260,N_29529,N_29879);
nand UO_1261 (O_1261,N_29736,N_29575);
xnor UO_1262 (O_1262,N_29774,N_29842);
or UO_1263 (O_1263,N_29764,N_29957);
and UO_1264 (O_1264,N_29907,N_29861);
nand UO_1265 (O_1265,N_29572,N_29832);
nor UO_1266 (O_1266,N_29599,N_29706);
and UO_1267 (O_1267,N_29700,N_29856);
xnor UO_1268 (O_1268,N_29547,N_29642);
xor UO_1269 (O_1269,N_29969,N_29918);
or UO_1270 (O_1270,N_29549,N_29804);
nand UO_1271 (O_1271,N_29612,N_29749);
nor UO_1272 (O_1272,N_29796,N_29539);
nand UO_1273 (O_1273,N_29848,N_29726);
nor UO_1274 (O_1274,N_29919,N_29719);
nor UO_1275 (O_1275,N_29576,N_29574);
nor UO_1276 (O_1276,N_29942,N_29584);
or UO_1277 (O_1277,N_29650,N_29937);
xnor UO_1278 (O_1278,N_29504,N_29964);
nand UO_1279 (O_1279,N_29548,N_29683);
nand UO_1280 (O_1280,N_29897,N_29555);
or UO_1281 (O_1281,N_29945,N_29520);
or UO_1282 (O_1282,N_29547,N_29992);
nand UO_1283 (O_1283,N_29806,N_29804);
nor UO_1284 (O_1284,N_29865,N_29720);
or UO_1285 (O_1285,N_29934,N_29932);
nor UO_1286 (O_1286,N_29500,N_29826);
or UO_1287 (O_1287,N_29666,N_29701);
nand UO_1288 (O_1288,N_29780,N_29621);
and UO_1289 (O_1289,N_29956,N_29979);
and UO_1290 (O_1290,N_29775,N_29636);
and UO_1291 (O_1291,N_29907,N_29818);
nand UO_1292 (O_1292,N_29578,N_29863);
nor UO_1293 (O_1293,N_29834,N_29921);
nand UO_1294 (O_1294,N_29660,N_29760);
nand UO_1295 (O_1295,N_29756,N_29717);
and UO_1296 (O_1296,N_29744,N_29878);
or UO_1297 (O_1297,N_29673,N_29925);
nor UO_1298 (O_1298,N_29612,N_29799);
and UO_1299 (O_1299,N_29567,N_29721);
nor UO_1300 (O_1300,N_29933,N_29579);
or UO_1301 (O_1301,N_29939,N_29519);
or UO_1302 (O_1302,N_29605,N_29615);
or UO_1303 (O_1303,N_29816,N_29722);
and UO_1304 (O_1304,N_29848,N_29869);
nand UO_1305 (O_1305,N_29810,N_29932);
xnor UO_1306 (O_1306,N_29536,N_29742);
nand UO_1307 (O_1307,N_29614,N_29679);
xnor UO_1308 (O_1308,N_29670,N_29828);
xnor UO_1309 (O_1309,N_29602,N_29553);
xnor UO_1310 (O_1310,N_29867,N_29542);
nor UO_1311 (O_1311,N_29778,N_29999);
nor UO_1312 (O_1312,N_29710,N_29655);
xor UO_1313 (O_1313,N_29839,N_29669);
xor UO_1314 (O_1314,N_29743,N_29947);
xor UO_1315 (O_1315,N_29744,N_29883);
xnor UO_1316 (O_1316,N_29732,N_29917);
nor UO_1317 (O_1317,N_29655,N_29957);
and UO_1318 (O_1318,N_29597,N_29649);
nor UO_1319 (O_1319,N_29804,N_29745);
and UO_1320 (O_1320,N_29876,N_29537);
and UO_1321 (O_1321,N_29913,N_29676);
or UO_1322 (O_1322,N_29505,N_29800);
nand UO_1323 (O_1323,N_29679,N_29557);
nand UO_1324 (O_1324,N_29680,N_29699);
or UO_1325 (O_1325,N_29599,N_29992);
nor UO_1326 (O_1326,N_29876,N_29504);
or UO_1327 (O_1327,N_29715,N_29757);
xor UO_1328 (O_1328,N_29776,N_29809);
xnor UO_1329 (O_1329,N_29982,N_29508);
or UO_1330 (O_1330,N_29681,N_29976);
or UO_1331 (O_1331,N_29835,N_29849);
and UO_1332 (O_1332,N_29617,N_29960);
xor UO_1333 (O_1333,N_29833,N_29557);
or UO_1334 (O_1334,N_29914,N_29849);
and UO_1335 (O_1335,N_29925,N_29886);
xnor UO_1336 (O_1336,N_29641,N_29865);
or UO_1337 (O_1337,N_29858,N_29883);
nand UO_1338 (O_1338,N_29557,N_29556);
xnor UO_1339 (O_1339,N_29995,N_29861);
nand UO_1340 (O_1340,N_29602,N_29676);
xnor UO_1341 (O_1341,N_29924,N_29971);
xor UO_1342 (O_1342,N_29828,N_29741);
nand UO_1343 (O_1343,N_29624,N_29980);
xnor UO_1344 (O_1344,N_29818,N_29504);
nand UO_1345 (O_1345,N_29666,N_29868);
xnor UO_1346 (O_1346,N_29824,N_29561);
nand UO_1347 (O_1347,N_29900,N_29649);
xnor UO_1348 (O_1348,N_29819,N_29829);
nand UO_1349 (O_1349,N_29707,N_29888);
nand UO_1350 (O_1350,N_29968,N_29689);
nand UO_1351 (O_1351,N_29998,N_29852);
nand UO_1352 (O_1352,N_29572,N_29916);
nand UO_1353 (O_1353,N_29865,N_29957);
nor UO_1354 (O_1354,N_29501,N_29554);
xor UO_1355 (O_1355,N_29592,N_29688);
and UO_1356 (O_1356,N_29816,N_29900);
xor UO_1357 (O_1357,N_29677,N_29527);
xor UO_1358 (O_1358,N_29553,N_29735);
nand UO_1359 (O_1359,N_29848,N_29687);
nand UO_1360 (O_1360,N_29639,N_29654);
and UO_1361 (O_1361,N_29999,N_29577);
nand UO_1362 (O_1362,N_29705,N_29697);
or UO_1363 (O_1363,N_29864,N_29983);
nand UO_1364 (O_1364,N_29706,N_29921);
nor UO_1365 (O_1365,N_29576,N_29639);
xor UO_1366 (O_1366,N_29604,N_29500);
xor UO_1367 (O_1367,N_29840,N_29971);
xnor UO_1368 (O_1368,N_29688,N_29737);
nand UO_1369 (O_1369,N_29937,N_29760);
nand UO_1370 (O_1370,N_29602,N_29705);
or UO_1371 (O_1371,N_29568,N_29911);
xor UO_1372 (O_1372,N_29672,N_29894);
nor UO_1373 (O_1373,N_29922,N_29850);
nor UO_1374 (O_1374,N_29595,N_29816);
xor UO_1375 (O_1375,N_29909,N_29655);
and UO_1376 (O_1376,N_29601,N_29863);
nor UO_1377 (O_1377,N_29581,N_29679);
and UO_1378 (O_1378,N_29856,N_29610);
xnor UO_1379 (O_1379,N_29987,N_29655);
and UO_1380 (O_1380,N_29733,N_29632);
and UO_1381 (O_1381,N_29505,N_29629);
nor UO_1382 (O_1382,N_29823,N_29793);
xnor UO_1383 (O_1383,N_29684,N_29651);
and UO_1384 (O_1384,N_29810,N_29755);
or UO_1385 (O_1385,N_29966,N_29762);
xor UO_1386 (O_1386,N_29946,N_29905);
nor UO_1387 (O_1387,N_29800,N_29824);
nand UO_1388 (O_1388,N_29679,N_29595);
and UO_1389 (O_1389,N_29861,N_29548);
or UO_1390 (O_1390,N_29540,N_29841);
nor UO_1391 (O_1391,N_29707,N_29719);
nand UO_1392 (O_1392,N_29858,N_29998);
xnor UO_1393 (O_1393,N_29710,N_29838);
nor UO_1394 (O_1394,N_29747,N_29704);
nor UO_1395 (O_1395,N_29587,N_29653);
nor UO_1396 (O_1396,N_29617,N_29630);
and UO_1397 (O_1397,N_29936,N_29751);
nand UO_1398 (O_1398,N_29681,N_29852);
xnor UO_1399 (O_1399,N_29635,N_29557);
or UO_1400 (O_1400,N_29610,N_29615);
and UO_1401 (O_1401,N_29506,N_29847);
nand UO_1402 (O_1402,N_29515,N_29601);
xor UO_1403 (O_1403,N_29592,N_29910);
nor UO_1404 (O_1404,N_29827,N_29633);
nor UO_1405 (O_1405,N_29906,N_29594);
xor UO_1406 (O_1406,N_29835,N_29832);
and UO_1407 (O_1407,N_29623,N_29830);
nor UO_1408 (O_1408,N_29706,N_29526);
and UO_1409 (O_1409,N_29987,N_29501);
or UO_1410 (O_1410,N_29875,N_29892);
xor UO_1411 (O_1411,N_29996,N_29509);
or UO_1412 (O_1412,N_29885,N_29691);
nor UO_1413 (O_1413,N_29655,N_29613);
nand UO_1414 (O_1414,N_29731,N_29730);
nand UO_1415 (O_1415,N_29514,N_29673);
or UO_1416 (O_1416,N_29609,N_29689);
nor UO_1417 (O_1417,N_29525,N_29606);
xor UO_1418 (O_1418,N_29808,N_29553);
nor UO_1419 (O_1419,N_29824,N_29724);
and UO_1420 (O_1420,N_29825,N_29647);
nor UO_1421 (O_1421,N_29510,N_29731);
xnor UO_1422 (O_1422,N_29897,N_29616);
and UO_1423 (O_1423,N_29811,N_29512);
nand UO_1424 (O_1424,N_29502,N_29944);
and UO_1425 (O_1425,N_29671,N_29642);
and UO_1426 (O_1426,N_29594,N_29817);
xnor UO_1427 (O_1427,N_29502,N_29546);
xnor UO_1428 (O_1428,N_29680,N_29782);
nand UO_1429 (O_1429,N_29569,N_29504);
nand UO_1430 (O_1430,N_29616,N_29735);
or UO_1431 (O_1431,N_29805,N_29563);
and UO_1432 (O_1432,N_29598,N_29888);
and UO_1433 (O_1433,N_29716,N_29864);
nor UO_1434 (O_1434,N_29638,N_29686);
nor UO_1435 (O_1435,N_29777,N_29748);
nor UO_1436 (O_1436,N_29759,N_29701);
nand UO_1437 (O_1437,N_29854,N_29835);
xnor UO_1438 (O_1438,N_29782,N_29615);
nor UO_1439 (O_1439,N_29533,N_29849);
xnor UO_1440 (O_1440,N_29921,N_29840);
xnor UO_1441 (O_1441,N_29740,N_29783);
xnor UO_1442 (O_1442,N_29991,N_29674);
and UO_1443 (O_1443,N_29629,N_29728);
nand UO_1444 (O_1444,N_29916,N_29567);
or UO_1445 (O_1445,N_29547,N_29565);
or UO_1446 (O_1446,N_29913,N_29963);
nand UO_1447 (O_1447,N_29662,N_29746);
xor UO_1448 (O_1448,N_29629,N_29833);
and UO_1449 (O_1449,N_29621,N_29657);
and UO_1450 (O_1450,N_29755,N_29574);
and UO_1451 (O_1451,N_29696,N_29541);
or UO_1452 (O_1452,N_29690,N_29722);
xnor UO_1453 (O_1453,N_29927,N_29936);
or UO_1454 (O_1454,N_29529,N_29613);
and UO_1455 (O_1455,N_29717,N_29620);
and UO_1456 (O_1456,N_29805,N_29648);
nor UO_1457 (O_1457,N_29851,N_29702);
xnor UO_1458 (O_1458,N_29702,N_29608);
nor UO_1459 (O_1459,N_29952,N_29598);
or UO_1460 (O_1460,N_29953,N_29589);
or UO_1461 (O_1461,N_29570,N_29505);
or UO_1462 (O_1462,N_29921,N_29643);
nor UO_1463 (O_1463,N_29751,N_29938);
nand UO_1464 (O_1464,N_29844,N_29762);
nand UO_1465 (O_1465,N_29800,N_29507);
nand UO_1466 (O_1466,N_29881,N_29763);
or UO_1467 (O_1467,N_29599,N_29761);
nor UO_1468 (O_1468,N_29836,N_29561);
and UO_1469 (O_1469,N_29801,N_29960);
nand UO_1470 (O_1470,N_29702,N_29883);
xor UO_1471 (O_1471,N_29949,N_29891);
or UO_1472 (O_1472,N_29789,N_29678);
xnor UO_1473 (O_1473,N_29975,N_29913);
nand UO_1474 (O_1474,N_29956,N_29914);
nand UO_1475 (O_1475,N_29957,N_29558);
nor UO_1476 (O_1476,N_29561,N_29660);
xor UO_1477 (O_1477,N_29626,N_29660);
and UO_1478 (O_1478,N_29641,N_29730);
nand UO_1479 (O_1479,N_29803,N_29626);
nor UO_1480 (O_1480,N_29961,N_29715);
nor UO_1481 (O_1481,N_29605,N_29932);
or UO_1482 (O_1482,N_29811,N_29587);
xnor UO_1483 (O_1483,N_29543,N_29501);
nand UO_1484 (O_1484,N_29776,N_29680);
nand UO_1485 (O_1485,N_29529,N_29952);
and UO_1486 (O_1486,N_29512,N_29645);
nand UO_1487 (O_1487,N_29964,N_29883);
nand UO_1488 (O_1488,N_29798,N_29545);
nand UO_1489 (O_1489,N_29571,N_29674);
or UO_1490 (O_1490,N_29584,N_29606);
nand UO_1491 (O_1491,N_29738,N_29525);
nor UO_1492 (O_1492,N_29701,N_29521);
nand UO_1493 (O_1493,N_29703,N_29972);
xnor UO_1494 (O_1494,N_29528,N_29868);
or UO_1495 (O_1495,N_29644,N_29833);
nor UO_1496 (O_1496,N_29629,N_29600);
xnor UO_1497 (O_1497,N_29658,N_29783);
and UO_1498 (O_1498,N_29865,N_29722);
or UO_1499 (O_1499,N_29658,N_29600);
and UO_1500 (O_1500,N_29895,N_29816);
nor UO_1501 (O_1501,N_29848,N_29710);
and UO_1502 (O_1502,N_29934,N_29542);
nand UO_1503 (O_1503,N_29941,N_29619);
or UO_1504 (O_1504,N_29757,N_29870);
nand UO_1505 (O_1505,N_29946,N_29691);
nor UO_1506 (O_1506,N_29760,N_29701);
nand UO_1507 (O_1507,N_29646,N_29931);
xor UO_1508 (O_1508,N_29553,N_29724);
or UO_1509 (O_1509,N_29680,N_29705);
xnor UO_1510 (O_1510,N_29686,N_29619);
and UO_1511 (O_1511,N_29763,N_29647);
xnor UO_1512 (O_1512,N_29889,N_29688);
nand UO_1513 (O_1513,N_29749,N_29956);
and UO_1514 (O_1514,N_29731,N_29880);
nand UO_1515 (O_1515,N_29730,N_29887);
nor UO_1516 (O_1516,N_29904,N_29630);
nand UO_1517 (O_1517,N_29683,N_29620);
or UO_1518 (O_1518,N_29681,N_29832);
xor UO_1519 (O_1519,N_29977,N_29948);
nor UO_1520 (O_1520,N_29796,N_29828);
or UO_1521 (O_1521,N_29894,N_29698);
and UO_1522 (O_1522,N_29530,N_29924);
nor UO_1523 (O_1523,N_29969,N_29749);
or UO_1524 (O_1524,N_29886,N_29510);
nand UO_1525 (O_1525,N_29794,N_29697);
and UO_1526 (O_1526,N_29554,N_29838);
and UO_1527 (O_1527,N_29824,N_29873);
nor UO_1528 (O_1528,N_29992,N_29558);
nand UO_1529 (O_1529,N_29608,N_29601);
and UO_1530 (O_1530,N_29839,N_29763);
and UO_1531 (O_1531,N_29684,N_29900);
or UO_1532 (O_1532,N_29689,N_29648);
and UO_1533 (O_1533,N_29798,N_29698);
xor UO_1534 (O_1534,N_29591,N_29531);
and UO_1535 (O_1535,N_29836,N_29815);
or UO_1536 (O_1536,N_29816,N_29607);
and UO_1537 (O_1537,N_29865,N_29712);
nand UO_1538 (O_1538,N_29798,N_29770);
nor UO_1539 (O_1539,N_29733,N_29546);
nand UO_1540 (O_1540,N_29784,N_29786);
xor UO_1541 (O_1541,N_29722,N_29718);
and UO_1542 (O_1542,N_29876,N_29591);
xnor UO_1543 (O_1543,N_29866,N_29895);
xnor UO_1544 (O_1544,N_29535,N_29875);
nand UO_1545 (O_1545,N_29666,N_29639);
xor UO_1546 (O_1546,N_29996,N_29644);
and UO_1547 (O_1547,N_29879,N_29932);
or UO_1548 (O_1548,N_29961,N_29798);
nand UO_1549 (O_1549,N_29762,N_29571);
nor UO_1550 (O_1550,N_29993,N_29600);
nor UO_1551 (O_1551,N_29880,N_29763);
and UO_1552 (O_1552,N_29903,N_29710);
nand UO_1553 (O_1553,N_29527,N_29793);
and UO_1554 (O_1554,N_29771,N_29591);
nor UO_1555 (O_1555,N_29683,N_29728);
nand UO_1556 (O_1556,N_29511,N_29759);
xor UO_1557 (O_1557,N_29987,N_29641);
and UO_1558 (O_1558,N_29617,N_29783);
or UO_1559 (O_1559,N_29629,N_29927);
xor UO_1560 (O_1560,N_29929,N_29679);
nand UO_1561 (O_1561,N_29528,N_29975);
and UO_1562 (O_1562,N_29646,N_29933);
and UO_1563 (O_1563,N_29699,N_29564);
nor UO_1564 (O_1564,N_29725,N_29597);
or UO_1565 (O_1565,N_29891,N_29578);
nor UO_1566 (O_1566,N_29575,N_29920);
nand UO_1567 (O_1567,N_29864,N_29543);
nand UO_1568 (O_1568,N_29934,N_29721);
or UO_1569 (O_1569,N_29734,N_29884);
or UO_1570 (O_1570,N_29947,N_29521);
and UO_1571 (O_1571,N_29503,N_29528);
nand UO_1572 (O_1572,N_29717,N_29558);
nor UO_1573 (O_1573,N_29598,N_29964);
xor UO_1574 (O_1574,N_29998,N_29875);
nand UO_1575 (O_1575,N_29816,N_29566);
nand UO_1576 (O_1576,N_29681,N_29887);
or UO_1577 (O_1577,N_29817,N_29700);
nor UO_1578 (O_1578,N_29965,N_29619);
xnor UO_1579 (O_1579,N_29647,N_29655);
and UO_1580 (O_1580,N_29998,N_29697);
and UO_1581 (O_1581,N_29802,N_29712);
xnor UO_1582 (O_1582,N_29762,N_29657);
nand UO_1583 (O_1583,N_29799,N_29903);
xor UO_1584 (O_1584,N_29948,N_29524);
xnor UO_1585 (O_1585,N_29626,N_29919);
xnor UO_1586 (O_1586,N_29626,N_29616);
nor UO_1587 (O_1587,N_29968,N_29979);
and UO_1588 (O_1588,N_29928,N_29720);
or UO_1589 (O_1589,N_29861,N_29853);
nand UO_1590 (O_1590,N_29997,N_29683);
and UO_1591 (O_1591,N_29912,N_29765);
nor UO_1592 (O_1592,N_29774,N_29653);
nor UO_1593 (O_1593,N_29993,N_29838);
nand UO_1594 (O_1594,N_29570,N_29986);
nor UO_1595 (O_1595,N_29820,N_29890);
xnor UO_1596 (O_1596,N_29919,N_29836);
and UO_1597 (O_1597,N_29508,N_29630);
and UO_1598 (O_1598,N_29775,N_29550);
or UO_1599 (O_1599,N_29774,N_29682);
and UO_1600 (O_1600,N_29630,N_29705);
nor UO_1601 (O_1601,N_29676,N_29741);
nand UO_1602 (O_1602,N_29957,N_29571);
nand UO_1603 (O_1603,N_29867,N_29976);
nor UO_1604 (O_1604,N_29960,N_29902);
and UO_1605 (O_1605,N_29991,N_29989);
and UO_1606 (O_1606,N_29987,N_29678);
or UO_1607 (O_1607,N_29626,N_29701);
xnor UO_1608 (O_1608,N_29886,N_29595);
xor UO_1609 (O_1609,N_29548,N_29620);
and UO_1610 (O_1610,N_29658,N_29503);
nand UO_1611 (O_1611,N_29836,N_29711);
or UO_1612 (O_1612,N_29918,N_29575);
and UO_1613 (O_1613,N_29541,N_29912);
nand UO_1614 (O_1614,N_29668,N_29972);
and UO_1615 (O_1615,N_29820,N_29550);
and UO_1616 (O_1616,N_29545,N_29544);
or UO_1617 (O_1617,N_29856,N_29936);
or UO_1618 (O_1618,N_29662,N_29732);
nor UO_1619 (O_1619,N_29725,N_29711);
nor UO_1620 (O_1620,N_29656,N_29824);
and UO_1621 (O_1621,N_29891,N_29868);
and UO_1622 (O_1622,N_29720,N_29812);
nor UO_1623 (O_1623,N_29879,N_29673);
and UO_1624 (O_1624,N_29508,N_29681);
nand UO_1625 (O_1625,N_29773,N_29918);
xnor UO_1626 (O_1626,N_29726,N_29608);
xnor UO_1627 (O_1627,N_29521,N_29829);
nand UO_1628 (O_1628,N_29767,N_29882);
and UO_1629 (O_1629,N_29915,N_29591);
xnor UO_1630 (O_1630,N_29724,N_29729);
nor UO_1631 (O_1631,N_29925,N_29913);
or UO_1632 (O_1632,N_29620,N_29770);
and UO_1633 (O_1633,N_29666,N_29774);
nand UO_1634 (O_1634,N_29897,N_29772);
nor UO_1635 (O_1635,N_29962,N_29616);
and UO_1636 (O_1636,N_29634,N_29929);
nand UO_1637 (O_1637,N_29728,N_29695);
nand UO_1638 (O_1638,N_29782,N_29886);
or UO_1639 (O_1639,N_29879,N_29639);
nor UO_1640 (O_1640,N_29750,N_29720);
and UO_1641 (O_1641,N_29848,N_29800);
nor UO_1642 (O_1642,N_29718,N_29671);
xnor UO_1643 (O_1643,N_29853,N_29885);
nand UO_1644 (O_1644,N_29532,N_29812);
and UO_1645 (O_1645,N_29884,N_29508);
nor UO_1646 (O_1646,N_29766,N_29826);
and UO_1647 (O_1647,N_29517,N_29578);
xnor UO_1648 (O_1648,N_29936,N_29756);
nor UO_1649 (O_1649,N_29922,N_29709);
nor UO_1650 (O_1650,N_29956,N_29765);
xnor UO_1651 (O_1651,N_29502,N_29946);
xor UO_1652 (O_1652,N_29946,N_29829);
nor UO_1653 (O_1653,N_29713,N_29548);
nand UO_1654 (O_1654,N_29700,N_29809);
and UO_1655 (O_1655,N_29954,N_29741);
xnor UO_1656 (O_1656,N_29984,N_29876);
xor UO_1657 (O_1657,N_29596,N_29534);
xnor UO_1658 (O_1658,N_29519,N_29979);
nand UO_1659 (O_1659,N_29882,N_29571);
xnor UO_1660 (O_1660,N_29758,N_29669);
nand UO_1661 (O_1661,N_29855,N_29537);
nand UO_1662 (O_1662,N_29510,N_29775);
xnor UO_1663 (O_1663,N_29910,N_29608);
and UO_1664 (O_1664,N_29506,N_29990);
and UO_1665 (O_1665,N_29791,N_29740);
or UO_1666 (O_1666,N_29786,N_29792);
xnor UO_1667 (O_1667,N_29849,N_29998);
nor UO_1668 (O_1668,N_29970,N_29634);
or UO_1669 (O_1669,N_29879,N_29979);
and UO_1670 (O_1670,N_29656,N_29752);
or UO_1671 (O_1671,N_29983,N_29962);
xor UO_1672 (O_1672,N_29692,N_29616);
nand UO_1673 (O_1673,N_29829,N_29812);
xor UO_1674 (O_1674,N_29745,N_29574);
xnor UO_1675 (O_1675,N_29795,N_29867);
nor UO_1676 (O_1676,N_29984,N_29939);
or UO_1677 (O_1677,N_29649,N_29715);
or UO_1678 (O_1678,N_29863,N_29761);
or UO_1679 (O_1679,N_29756,N_29589);
and UO_1680 (O_1680,N_29616,N_29805);
and UO_1681 (O_1681,N_29722,N_29948);
nor UO_1682 (O_1682,N_29665,N_29682);
nor UO_1683 (O_1683,N_29639,N_29593);
nand UO_1684 (O_1684,N_29839,N_29939);
nand UO_1685 (O_1685,N_29731,N_29718);
nand UO_1686 (O_1686,N_29561,N_29906);
or UO_1687 (O_1687,N_29694,N_29892);
and UO_1688 (O_1688,N_29777,N_29587);
or UO_1689 (O_1689,N_29736,N_29637);
xnor UO_1690 (O_1690,N_29888,N_29886);
xnor UO_1691 (O_1691,N_29939,N_29837);
or UO_1692 (O_1692,N_29845,N_29530);
and UO_1693 (O_1693,N_29802,N_29678);
or UO_1694 (O_1694,N_29689,N_29883);
xor UO_1695 (O_1695,N_29977,N_29884);
or UO_1696 (O_1696,N_29857,N_29803);
and UO_1697 (O_1697,N_29772,N_29569);
nor UO_1698 (O_1698,N_29599,N_29593);
xor UO_1699 (O_1699,N_29768,N_29513);
xnor UO_1700 (O_1700,N_29636,N_29943);
xor UO_1701 (O_1701,N_29854,N_29641);
nor UO_1702 (O_1702,N_29954,N_29642);
and UO_1703 (O_1703,N_29700,N_29509);
or UO_1704 (O_1704,N_29734,N_29925);
nor UO_1705 (O_1705,N_29830,N_29918);
nand UO_1706 (O_1706,N_29749,N_29665);
and UO_1707 (O_1707,N_29945,N_29863);
and UO_1708 (O_1708,N_29843,N_29998);
and UO_1709 (O_1709,N_29984,N_29973);
nand UO_1710 (O_1710,N_29924,N_29569);
or UO_1711 (O_1711,N_29674,N_29989);
nand UO_1712 (O_1712,N_29556,N_29616);
xor UO_1713 (O_1713,N_29658,N_29729);
nand UO_1714 (O_1714,N_29620,N_29784);
nand UO_1715 (O_1715,N_29709,N_29699);
and UO_1716 (O_1716,N_29700,N_29556);
and UO_1717 (O_1717,N_29951,N_29504);
xnor UO_1718 (O_1718,N_29948,N_29501);
or UO_1719 (O_1719,N_29759,N_29688);
nand UO_1720 (O_1720,N_29726,N_29644);
nor UO_1721 (O_1721,N_29580,N_29525);
nor UO_1722 (O_1722,N_29622,N_29912);
nand UO_1723 (O_1723,N_29730,N_29553);
nand UO_1724 (O_1724,N_29633,N_29526);
and UO_1725 (O_1725,N_29606,N_29713);
and UO_1726 (O_1726,N_29795,N_29539);
nand UO_1727 (O_1727,N_29670,N_29927);
nand UO_1728 (O_1728,N_29576,N_29812);
xnor UO_1729 (O_1729,N_29883,N_29734);
nand UO_1730 (O_1730,N_29784,N_29708);
nand UO_1731 (O_1731,N_29913,N_29699);
or UO_1732 (O_1732,N_29753,N_29887);
nor UO_1733 (O_1733,N_29976,N_29948);
nor UO_1734 (O_1734,N_29835,N_29756);
xnor UO_1735 (O_1735,N_29753,N_29716);
and UO_1736 (O_1736,N_29584,N_29682);
nand UO_1737 (O_1737,N_29591,N_29519);
nand UO_1738 (O_1738,N_29595,N_29845);
nor UO_1739 (O_1739,N_29666,N_29638);
xnor UO_1740 (O_1740,N_29940,N_29581);
xor UO_1741 (O_1741,N_29664,N_29520);
xnor UO_1742 (O_1742,N_29995,N_29756);
or UO_1743 (O_1743,N_29721,N_29615);
and UO_1744 (O_1744,N_29846,N_29931);
and UO_1745 (O_1745,N_29913,N_29737);
xor UO_1746 (O_1746,N_29808,N_29644);
nor UO_1747 (O_1747,N_29960,N_29904);
and UO_1748 (O_1748,N_29734,N_29950);
nor UO_1749 (O_1749,N_29828,N_29816);
and UO_1750 (O_1750,N_29659,N_29564);
nor UO_1751 (O_1751,N_29903,N_29658);
xor UO_1752 (O_1752,N_29677,N_29603);
xor UO_1753 (O_1753,N_29682,N_29588);
and UO_1754 (O_1754,N_29967,N_29861);
or UO_1755 (O_1755,N_29592,N_29743);
nor UO_1756 (O_1756,N_29700,N_29761);
and UO_1757 (O_1757,N_29979,N_29914);
and UO_1758 (O_1758,N_29848,N_29556);
xor UO_1759 (O_1759,N_29933,N_29791);
nor UO_1760 (O_1760,N_29729,N_29665);
and UO_1761 (O_1761,N_29765,N_29871);
xor UO_1762 (O_1762,N_29910,N_29625);
or UO_1763 (O_1763,N_29829,N_29637);
xor UO_1764 (O_1764,N_29698,N_29891);
nand UO_1765 (O_1765,N_29904,N_29708);
xnor UO_1766 (O_1766,N_29853,N_29782);
nand UO_1767 (O_1767,N_29869,N_29701);
nor UO_1768 (O_1768,N_29704,N_29540);
nand UO_1769 (O_1769,N_29997,N_29872);
or UO_1770 (O_1770,N_29533,N_29656);
xor UO_1771 (O_1771,N_29737,N_29599);
and UO_1772 (O_1772,N_29992,N_29854);
nand UO_1773 (O_1773,N_29842,N_29777);
or UO_1774 (O_1774,N_29765,N_29515);
xnor UO_1775 (O_1775,N_29802,N_29904);
nand UO_1776 (O_1776,N_29669,N_29775);
nand UO_1777 (O_1777,N_29963,N_29872);
nor UO_1778 (O_1778,N_29610,N_29902);
and UO_1779 (O_1779,N_29969,N_29861);
or UO_1780 (O_1780,N_29621,N_29822);
nor UO_1781 (O_1781,N_29940,N_29964);
and UO_1782 (O_1782,N_29765,N_29768);
xor UO_1783 (O_1783,N_29533,N_29709);
nand UO_1784 (O_1784,N_29904,N_29515);
nor UO_1785 (O_1785,N_29877,N_29985);
or UO_1786 (O_1786,N_29503,N_29919);
and UO_1787 (O_1787,N_29714,N_29554);
nor UO_1788 (O_1788,N_29671,N_29576);
xor UO_1789 (O_1789,N_29791,N_29744);
or UO_1790 (O_1790,N_29848,N_29592);
or UO_1791 (O_1791,N_29634,N_29714);
and UO_1792 (O_1792,N_29856,N_29981);
xor UO_1793 (O_1793,N_29822,N_29561);
xnor UO_1794 (O_1794,N_29885,N_29801);
nor UO_1795 (O_1795,N_29926,N_29534);
and UO_1796 (O_1796,N_29839,N_29829);
nor UO_1797 (O_1797,N_29946,N_29558);
nor UO_1798 (O_1798,N_29903,N_29758);
nor UO_1799 (O_1799,N_29778,N_29973);
xor UO_1800 (O_1800,N_29910,N_29598);
and UO_1801 (O_1801,N_29669,N_29601);
or UO_1802 (O_1802,N_29505,N_29801);
nand UO_1803 (O_1803,N_29625,N_29584);
xor UO_1804 (O_1804,N_29967,N_29991);
xnor UO_1805 (O_1805,N_29603,N_29503);
nand UO_1806 (O_1806,N_29682,N_29890);
nand UO_1807 (O_1807,N_29628,N_29545);
and UO_1808 (O_1808,N_29875,N_29707);
nor UO_1809 (O_1809,N_29737,N_29536);
nand UO_1810 (O_1810,N_29875,N_29634);
nand UO_1811 (O_1811,N_29845,N_29955);
nand UO_1812 (O_1812,N_29586,N_29764);
and UO_1813 (O_1813,N_29972,N_29732);
nand UO_1814 (O_1814,N_29508,N_29592);
or UO_1815 (O_1815,N_29816,N_29759);
and UO_1816 (O_1816,N_29667,N_29593);
or UO_1817 (O_1817,N_29972,N_29572);
xor UO_1818 (O_1818,N_29613,N_29949);
nand UO_1819 (O_1819,N_29556,N_29524);
nand UO_1820 (O_1820,N_29528,N_29998);
and UO_1821 (O_1821,N_29743,N_29557);
and UO_1822 (O_1822,N_29513,N_29976);
nand UO_1823 (O_1823,N_29837,N_29543);
nand UO_1824 (O_1824,N_29819,N_29800);
xnor UO_1825 (O_1825,N_29748,N_29991);
nand UO_1826 (O_1826,N_29647,N_29715);
xor UO_1827 (O_1827,N_29577,N_29521);
or UO_1828 (O_1828,N_29883,N_29898);
or UO_1829 (O_1829,N_29821,N_29681);
and UO_1830 (O_1830,N_29544,N_29772);
nor UO_1831 (O_1831,N_29800,N_29790);
and UO_1832 (O_1832,N_29824,N_29748);
nor UO_1833 (O_1833,N_29873,N_29519);
or UO_1834 (O_1834,N_29680,N_29797);
or UO_1835 (O_1835,N_29592,N_29796);
and UO_1836 (O_1836,N_29786,N_29938);
nand UO_1837 (O_1837,N_29722,N_29848);
nand UO_1838 (O_1838,N_29617,N_29966);
and UO_1839 (O_1839,N_29899,N_29545);
or UO_1840 (O_1840,N_29993,N_29596);
and UO_1841 (O_1841,N_29921,N_29732);
nor UO_1842 (O_1842,N_29657,N_29889);
or UO_1843 (O_1843,N_29827,N_29699);
nor UO_1844 (O_1844,N_29634,N_29539);
nor UO_1845 (O_1845,N_29875,N_29652);
or UO_1846 (O_1846,N_29551,N_29707);
or UO_1847 (O_1847,N_29667,N_29898);
and UO_1848 (O_1848,N_29932,N_29898);
nor UO_1849 (O_1849,N_29868,N_29945);
nor UO_1850 (O_1850,N_29888,N_29786);
nor UO_1851 (O_1851,N_29638,N_29846);
nor UO_1852 (O_1852,N_29926,N_29823);
and UO_1853 (O_1853,N_29685,N_29980);
nor UO_1854 (O_1854,N_29554,N_29814);
and UO_1855 (O_1855,N_29616,N_29598);
and UO_1856 (O_1856,N_29839,N_29876);
and UO_1857 (O_1857,N_29822,N_29944);
nor UO_1858 (O_1858,N_29680,N_29583);
and UO_1859 (O_1859,N_29533,N_29777);
nand UO_1860 (O_1860,N_29769,N_29843);
nor UO_1861 (O_1861,N_29656,N_29640);
and UO_1862 (O_1862,N_29896,N_29827);
and UO_1863 (O_1863,N_29952,N_29803);
xnor UO_1864 (O_1864,N_29998,N_29816);
nand UO_1865 (O_1865,N_29569,N_29873);
nand UO_1866 (O_1866,N_29622,N_29829);
nor UO_1867 (O_1867,N_29727,N_29860);
nand UO_1868 (O_1868,N_29799,N_29611);
or UO_1869 (O_1869,N_29718,N_29568);
and UO_1870 (O_1870,N_29829,N_29861);
nor UO_1871 (O_1871,N_29753,N_29780);
nor UO_1872 (O_1872,N_29701,N_29596);
nor UO_1873 (O_1873,N_29609,N_29698);
nor UO_1874 (O_1874,N_29735,N_29816);
xnor UO_1875 (O_1875,N_29950,N_29989);
nor UO_1876 (O_1876,N_29831,N_29786);
nand UO_1877 (O_1877,N_29937,N_29637);
and UO_1878 (O_1878,N_29562,N_29754);
nor UO_1879 (O_1879,N_29926,N_29573);
xor UO_1880 (O_1880,N_29618,N_29647);
or UO_1881 (O_1881,N_29821,N_29686);
nand UO_1882 (O_1882,N_29913,N_29810);
or UO_1883 (O_1883,N_29839,N_29711);
and UO_1884 (O_1884,N_29892,N_29818);
nand UO_1885 (O_1885,N_29503,N_29895);
or UO_1886 (O_1886,N_29668,N_29878);
and UO_1887 (O_1887,N_29895,N_29569);
nor UO_1888 (O_1888,N_29685,N_29662);
nor UO_1889 (O_1889,N_29765,N_29521);
and UO_1890 (O_1890,N_29703,N_29749);
xor UO_1891 (O_1891,N_29920,N_29810);
nor UO_1892 (O_1892,N_29708,N_29588);
or UO_1893 (O_1893,N_29661,N_29825);
and UO_1894 (O_1894,N_29719,N_29711);
or UO_1895 (O_1895,N_29685,N_29794);
nand UO_1896 (O_1896,N_29956,N_29882);
nor UO_1897 (O_1897,N_29711,N_29956);
xor UO_1898 (O_1898,N_29855,N_29644);
and UO_1899 (O_1899,N_29558,N_29995);
or UO_1900 (O_1900,N_29867,N_29839);
and UO_1901 (O_1901,N_29839,N_29789);
xor UO_1902 (O_1902,N_29559,N_29772);
nand UO_1903 (O_1903,N_29633,N_29826);
xor UO_1904 (O_1904,N_29777,N_29949);
or UO_1905 (O_1905,N_29958,N_29642);
nand UO_1906 (O_1906,N_29916,N_29925);
nand UO_1907 (O_1907,N_29693,N_29788);
nand UO_1908 (O_1908,N_29865,N_29622);
or UO_1909 (O_1909,N_29787,N_29820);
nor UO_1910 (O_1910,N_29805,N_29874);
and UO_1911 (O_1911,N_29811,N_29987);
nor UO_1912 (O_1912,N_29937,N_29881);
nand UO_1913 (O_1913,N_29712,N_29815);
nand UO_1914 (O_1914,N_29951,N_29522);
and UO_1915 (O_1915,N_29597,N_29878);
nand UO_1916 (O_1916,N_29597,N_29836);
and UO_1917 (O_1917,N_29957,N_29854);
nand UO_1918 (O_1918,N_29526,N_29544);
xnor UO_1919 (O_1919,N_29552,N_29502);
xnor UO_1920 (O_1920,N_29656,N_29697);
and UO_1921 (O_1921,N_29754,N_29744);
or UO_1922 (O_1922,N_29814,N_29613);
xor UO_1923 (O_1923,N_29635,N_29995);
nand UO_1924 (O_1924,N_29866,N_29584);
nor UO_1925 (O_1925,N_29917,N_29652);
and UO_1926 (O_1926,N_29687,N_29500);
and UO_1927 (O_1927,N_29612,N_29995);
nand UO_1928 (O_1928,N_29550,N_29703);
nor UO_1929 (O_1929,N_29743,N_29998);
nor UO_1930 (O_1930,N_29844,N_29699);
xor UO_1931 (O_1931,N_29994,N_29713);
xor UO_1932 (O_1932,N_29929,N_29773);
nand UO_1933 (O_1933,N_29736,N_29849);
nor UO_1934 (O_1934,N_29993,N_29750);
nand UO_1935 (O_1935,N_29871,N_29975);
or UO_1936 (O_1936,N_29594,N_29641);
nor UO_1937 (O_1937,N_29814,N_29617);
nor UO_1938 (O_1938,N_29700,N_29613);
nor UO_1939 (O_1939,N_29989,N_29981);
nand UO_1940 (O_1940,N_29744,N_29668);
nand UO_1941 (O_1941,N_29844,N_29698);
nor UO_1942 (O_1942,N_29780,N_29691);
or UO_1943 (O_1943,N_29709,N_29771);
and UO_1944 (O_1944,N_29902,N_29688);
or UO_1945 (O_1945,N_29730,N_29771);
nand UO_1946 (O_1946,N_29559,N_29886);
xor UO_1947 (O_1947,N_29810,N_29565);
and UO_1948 (O_1948,N_29841,N_29821);
nand UO_1949 (O_1949,N_29700,N_29985);
or UO_1950 (O_1950,N_29615,N_29736);
xnor UO_1951 (O_1951,N_29791,N_29799);
nor UO_1952 (O_1952,N_29843,N_29862);
nor UO_1953 (O_1953,N_29520,N_29703);
nand UO_1954 (O_1954,N_29897,N_29721);
nor UO_1955 (O_1955,N_29722,N_29946);
and UO_1956 (O_1956,N_29923,N_29763);
xnor UO_1957 (O_1957,N_29691,N_29916);
nor UO_1958 (O_1958,N_29755,N_29820);
and UO_1959 (O_1959,N_29569,N_29718);
xnor UO_1960 (O_1960,N_29815,N_29517);
or UO_1961 (O_1961,N_29865,N_29813);
nor UO_1962 (O_1962,N_29775,N_29724);
xnor UO_1963 (O_1963,N_29671,N_29800);
xor UO_1964 (O_1964,N_29598,N_29815);
nand UO_1965 (O_1965,N_29623,N_29609);
or UO_1966 (O_1966,N_29834,N_29711);
nor UO_1967 (O_1967,N_29862,N_29994);
nor UO_1968 (O_1968,N_29721,N_29620);
and UO_1969 (O_1969,N_29652,N_29825);
nand UO_1970 (O_1970,N_29785,N_29584);
nor UO_1971 (O_1971,N_29538,N_29881);
nand UO_1972 (O_1972,N_29866,N_29790);
or UO_1973 (O_1973,N_29640,N_29942);
nand UO_1974 (O_1974,N_29957,N_29856);
nor UO_1975 (O_1975,N_29914,N_29532);
or UO_1976 (O_1976,N_29985,N_29897);
nor UO_1977 (O_1977,N_29863,N_29662);
nor UO_1978 (O_1978,N_29841,N_29656);
or UO_1979 (O_1979,N_29861,N_29839);
xor UO_1980 (O_1980,N_29638,N_29694);
nor UO_1981 (O_1981,N_29863,N_29607);
or UO_1982 (O_1982,N_29932,N_29651);
nor UO_1983 (O_1983,N_29805,N_29957);
and UO_1984 (O_1984,N_29984,N_29527);
nand UO_1985 (O_1985,N_29591,N_29959);
or UO_1986 (O_1986,N_29752,N_29894);
or UO_1987 (O_1987,N_29679,N_29588);
nand UO_1988 (O_1988,N_29869,N_29625);
or UO_1989 (O_1989,N_29674,N_29824);
nand UO_1990 (O_1990,N_29906,N_29600);
nor UO_1991 (O_1991,N_29860,N_29690);
or UO_1992 (O_1992,N_29511,N_29679);
and UO_1993 (O_1993,N_29713,N_29582);
nor UO_1994 (O_1994,N_29748,N_29807);
or UO_1995 (O_1995,N_29918,N_29978);
xor UO_1996 (O_1996,N_29751,N_29633);
xnor UO_1997 (O_1997,N_29789,N_29759);
or UO_1998 (O_1998,N_29750,N_29883);
and UO_1999 (O_1999,N_29663,N_29519);
or UO_2000 (O_2000,N_29577,N_29661);
nor UO_2001 (O_2001,N_29714,N_29538);
xor UO_2002 (O_2002,N_29950,N_29767);
or UO_2003 (O_2003,N_29959,N_29685);
and UO_2004 (O_2004,N_29525,N_29571);
and UO_2005 (O_2005,N_29991,N_29896);
or UO_2006 (O_2006,N_29914,N_29517);
nand UO_2007 (O_2007,N_29956,N_29764);
xor UO_2008 (O_2008,N_29723,N_29517);
nor UO_2009 (O_2009,N_29542,N_29874);
nor UO_2010 (O_2010,N_29931,N_29787);
and UO_2011 (O_2011,N_29649,N_29678);
nor UO_2012 (O_2012,N_29507,N_29502);
nand UO_2013 (O_2013,N_29837,N_29561);
and UO_2014 (O_2014,N_29558,N_29605);
nand UO_2015 (O_2015,N_29701,N_29942);
or UO_2016 (O_2016,N_29514,N_29757);
nand UO_2017 (O_2017,N_29730,N_29542);
or UO_2018 (O_2018,N_29776,N_29814);
and UO_2019 (O_2019,N_29597,N_29891);
and UO_2020 (O_2020,N_29630,N_29598);
or UO_2021 (O_2021,N_29516,N_29972);
nor UO_2022 (O_2022,N_29606,N_29656);
or UO_2023 (O_2023,N_29709,N_29784);
and UO_2024 (O_2024,N_29503,N_29771);
or UO_2025 (O_2025,N_29998,N_29804);
and UO_2026 (O_2026,N_29943,N_29786);
and UO_2027 (O_2027,N_29882,N_29856);
nand UO_2028 (O_2028,N_29607,N_29724);
nor UO_2029 (O_2029,N_29657,N_29939);
nor UO_2030 (O_2030,N_29502,N_29511);
nor UO_2031 (O_2031,N_29929,N_29966);
and UO_2032 (O_2032,N_29633,N_29670);
nor UO_2033 (O_2033,N_29873,N_29549);
nor UO_2034 (O_2034,N_29934,N_29589);
and UO_2035 (O_2035,N_29782,N_29798);
and UO_2036 (O_2036,N_29599,N_29842);
and UO_2037 (O_2037,N_29756,N_29794);
xor UO_2038 (O_2038,N_29605,N_29737);
nand UO_2039 (O_2039,N_29510,N_29501);
nor UO_2040 (O_2040,N_29738,N_29947);
nor UO_2041 (O_2041,N_29818,N_29587);
nand UO_2042 (O_2042,N_29899,N_29562);
xor UO_2043 (O_2043,N_29892,N_29941);
xnor UO_2044 (O_2044,N_29888,N_29933);
nand UO_2045 (O_2045,N_29838,N_29567);
nor UO_2046 (O_2046,N_29573,N_29902);
xor UO_2047 (O_2047,N_29802,N_29919);
xor UO_2048 (O_2048,N_29695,N_29553);
nor UO_2049 (O_2049,N_29879,N_29566);
or UO_2050 (O_2050,N_29857,N_29850);
nand UO_2051 (O_2051,N_29931,N_29650);
nor UO_2052 (O_2052,N_29539,N_29888);
or UO_2053 (O_2053,N_29763,N_29669);
or UO_2054 (O_2054,N_29820,N_29888);
or UO_2055 (O_2055,N_29587,N_29638);
xnor UO_2056 (O_2056,N_29977,N_29826);
and UO_2057 (O_2057,N_29957,N_29677);
or UO_2058 (O_2058,N_29839,N_29877);
nand UO_2059 (O_2059,N_29861,N_29840);
or UO_2060 (O_2060,N_29639,N_29721);
nor UO_2061 (O_2061,N_29615,N_29686);
nor UO_2062 (O_2062,N_29620,N_29903);
nand UO_2063 (O_2063,N_29828,N_29515);
or UO_2064 (O_2064,N_29680,N_29618);
nand UO_2065 (O_2065,N_29564,N_29539);
nor UO_2066 (O_2066,N_29628,N_29933);
and UO_2067 (O_2067,N_29715,N_29730);
nor UO_2068 (O_2068,N_29987,N_29567);
and UO_2069 (O_2069,N_29670,N_29805);
and UO_2070 (O_2070,N_29538,N_29703);
nand UO_2071 (O_2071,N_29832,N_29520);
xnor UO_2072 (O_2072,N_29920,N_29762);
nand UO_2073 (O_2073,N_29651,N_29951);
xnor UO_2074 (O_2074,N_29643,N_29698);
and UO_2075 (O_2075,N_29930,N_29526);
nor UO_2076 (O_2076,N_29533,N_29883);
xor UO_2077 (O_2077,N_29948,N_29962);
nor UO_2078 (O_2078,N_29738,N_29690);
nor UO_2079 (O_2079,N_29821,N_29848);
nor UO_2080 (O_2080,N_29527,N_29973);
nor UO_2081 (O_2081,N_29826,N_29800);
and UO_2082 (O_2082,N_29886,N_29868);
nor UO_2083 (O_2083,N_29545,N_29762);
nand UO_2084 (O_2084,N_29909,N_29550);
or UO_2085 (O_2085,N_29676,N_29871);
xnor UO_2086 (O_2086,N_29681,N_29879);
xor UO_2087 (O_2087,N_29884,N_29778);
nand UO_2088 (O_2088,N_29682,N_29563);
or UO_2089 (O_2089,N_29931,N_29783);
xor UO_2090 (O_2090,N_29625,N_29645);
and UO_2091 (O_2091,N_29802,N_29501);
and UO_2092 (O_2092,N_29649,N_29679);
nor UO_2093 (O_2093,N_29802,N_29613);
nand UO_2094 (O_2094,N_29677,N_29905);
and UO_2095 (O_2095,N_29960,N_29741);
nor UO_2096 (O_2096,N_29732,N_29595);
and UO_2097 (O_2097,N_29761,N_29997);
xor UO_2098 (O_2098,N_29966,N_29952);
nand UO_2099 (O_2099,N_29659,N_29859);
and UO_2100 (O_2100,N_29905,N_29578);
nand UO_2101 (O_2101,N_29673,N_29913);
nor UO_2102 (O_2102,N_29666,N_29611);
nand UO_2103 (O_2103,N_29885,N_29844);
nor UO_2104 (O_2104,N_29860,N_29984);
or UO_2105 (O_2105,N_29501,N_29921);
nor UO_2106 (O_2106,N_29667,N_29632);
and UO_2107 (O_2107,N_29656,N_29876);
xor UO_2108 (O_2108,N_29617,N_29967);
or UO_2109 (O_2109,N_29512,N_29606);
nand UO_2110 (O_2110,N_29731,N_29521);
and UO_2111 (O_2111,N_29599,N_29742);
or UO_2112 (O_2112,N_29928,N_29533);
nand UO_2113 (O_2113,N_29813,N_29891);
nor UO_2114 (O_2114,N_29546,N_29748);
xor UO_2115 (O_2115,N_29724,N_29712);
or UO_2116 (O_2116,N_29717,N_29527);
nand UO_2117 (O_2117,N_29844,N_29641);
or UO_2118 (O_2118,N_29710,N_29920);
xnor UO_2119 (O_2119,N_29713,N_29509);
nand UO_2120 (O_2120,N_29976,N_29853);
and UO_2121 (O_2121,N_29739,N_29616);
nor UO_2122 (O_2122,N_29532,N_29651);
and UO_2123 (O_2123,N_29596,N_29787);
or UO_2124 (O_2124,N_29693,N_29530);
xor UO_2125 (O_2125,N_29677,N_29626);
nand UO_2126 (O_2126,N_29609,N_29665);
xnor UO_2127 (O_2127,N_29526,N_29584);
nor UO_2128 (O_2128,N_29538,N_29564);
xor UO_2129 (O_2129,N_29882,N_29754);
nor UO_2130 (O_2130,N_29829,N_29576);
and UO_2131 (O_2131,N_29996,N_29736);
and UO_2132 (O_2132,N_29789,N_29595);
nor UO_2133 (O_2133,N_29593,N_29827);
xor UO_2134 (O_2134,N_29542,N_29614);
nand UO_2135 (O_2135,N_29537,N_29598);
nand UO_2136 (O_2136,N_29999,N_29688);
nand UO_2137 (O_2137,N_29691,N_29969);
nor UO_2138 (O_2138,N_29712,N_29554);
or UO_2139 (O_2139,N_29579,N_29910);
and UO_2140 (O_2140,N_29604,N_29573);
and UO_2141 (O_2141,N_29659,N_29668);
nor UO_2142 (O_2142,N_29625,N_29641);
xnor UO_2143 (O_2143,N_29877,N_29688);
or UO_2144 (O_2144,N_29919,N_29623);
and UO_2145 (O_2145,N_29704,N_29726);
xnor UO_2146 (O_2146,N_29920,N_29862);
and UO_2147 (O_2147,N_29651,N_29547);
and UO_2148 (O_2148,N_29945,N_29905);
nand UO_2149 (O_2149,N_29600,N_29692);
nand UO_2150 (O_2150,N_29557,N_29862);
nand UO_2151 (O_2151,N_29784,N_29664);
nand UO_2152 (O_2152,N_29886,N_29876);
and UO_2153 (O_2153,N_29731,N_29991);
and UO_2154 (O_2154,N_29659,N_29770);
xnor UO_2155 (O_2155,N_29949,N_29875);
or UO_2156 (O_2156,N_29876,N_29685);
or UO_2157 (O_2157,N_29723,N_29602);
or UO_2158 (O_2158,N_29934,N_29649);
nand UO_2159 (O_2159,N_29757,N_29987);
nand UO_2160 (O_2160,N_29658,N_29706);
nor UO_2161 (O_2161,N_29878,N_29696);
or UO_2162 (O_2162,N_29657,N_29886);
nand UO_2163 (O_2163,N_29644,N_29787);
nor UO_2164 (O_2164,N_29977,N_29912);
nor UO_2165 (O_2165,N_29883,N_29931);
or UO_2166 (O_2166,N_29844,N_29548);
or UO_2167 (O_2167,N_29514,N_29912);
or UO_2168 (O_2168,N_29912,N_29814);
nand UO_2169 (O_2169,N_29848,N_29983);
xnor UO_2170 (O_2170,N_29515,N_29865);
xor UO_2171 (O_2171,N_29887,N_29797);
or UO_2172 (O_2172,N_29977,N_29598);
nor UO_2173 (O_2173,N_29531,N_29543);
or UO_2174 (O_2174,N_29794,N_29545);
nor UO_2175 (O_2175,N_29768,N_29917);
nor UO_2176 (O_2176,N_29744,N_29603);
and UO_2177 (O_2177,N_29793,N_29746);
and UO_2178 (O_2178,N_29797,N_29523);
nand UO_2179 (O_2179,N_29726,N_29595);
nor UO_2180 (O_2180,N_29522,N_29982);
nand UO_2181 (O_2181,N_29827,N_29792);
or UO_2182 (O_2182,N_29929,N_29649);
or UO_2183 (O_2183,N_29759,N_29835);
xor UO_2184 (O_2184,N_29827,N_29964);
or UO_2185 (O_2185,N_29655,N_29531);
and UO_2186 (O_2186,N_29978,N_29956);
nor UO_2187 (O_2187,N_29551,N_29915);
or UO_2188 (O_2188,N_29774,N_29999);
xor UO_2189 (O_2189,N_29839,N_29723);
nand UO_2190 (O_2190,N_29981,N_29622);
or UO_2191 (O_2191,N_29568,N_29859);
or UO_2192 (O_2192,N_29993,N_29985);
nor UO_2193 (O_2193,N_29742,N_29840);
and UO_2194 (O_2194,N_29826,N_29728);
nor UO_2195 (O_2195,N_29709,N_29736);
xnor UO_2196 (O_2196,N_29680,N_29969);
xnor UO_2197 (O_2197,N_29634,N_29997);
xnor UO_2198 (O_2198,N_29754,N_29785);
nor UO_2199 (O_2199,N_29842,N_29697);
or UO_2200 (O_2200,N_29929,N_29526);
nor UO_2201 (O_2201,N_29530,N_29701);
or UO_2202 (O_2202,N_29751,N_29632);
xnor UO_2203 (O_2203,N_29669,N_29696);
or UO_2204 (O_2204,N_29678,N_29584);
xnor UO_2205 (O_2205,N_29633,N_29940);
nor UO_2206 (O_2206,N_29867,N_29898);
nand UO_2207 (O_2207,N_29672,N_29534);
xnor UO_2208 (O_2208,N_29794,N_29517);
nor UO_2209 (O_2209,N_29740,N_29594);
nand UO_2210 (O_2210,N_29648,N_29844);
nand UO_2211 (O_2211,N_29752,N_29979);
nor UO_2212 (O_2212,N_29590,N_29945);
and UO_2213 (O_2213,N_29920,N_29520);
nor UO_2214 (O_2214,N_29514,N_29549);
or UO_2215 (O_2215,N_29706,N_29971);
nand UO_2216 (O_2216,N_29953,N_29890);
xor UO_2217 (O_2217,N_29803,N_29978);
and UO_2218 (O_2218,N_29940,N_29993);
xnor UO_2219 (O_2219,N_29895,N_29659);
nand UO_2220 (O_2220,N_29561,N_29910);
and UO_2221 (O_2221,N_29659,N_29574);
nor UO_2222 (O_2222,N_29642,N_29881);
nand UO_2223 (O_2223,N_29885,N_29811);
nor UO_2224 (O_2224,N_29911,N_29607);
nand UO_2225 (O_2225,N_29533,N_29557);
and UO_2226 (O_2226,N_29732,N_29993);
and UO_2227 (O_2227,N_29989,N_29779);
nor UO_2228 (O_2228,N_29695,N_29741);
xnor UO_2229 (O_2229,N_29638,N_29913);
xor UO_2230 (O_2230,N_29946,N_29800);
xnor UO_2231 (O_2231,N_29931,N_29586);
nor UO_2232 (O_2232,N_29588,N_29527);
or UO_2233 (O_2233,N_29911,N_29686);
xnor UO_2234 (O_2234,N_29866,N_29897);
xor UO_2235 (O_2235,N_29962,N_29600);
and UO_2236 (O_2236,N_29671,N_29709);
xor UO_2237 (O_2237,N_29725,N_29850);
and UO_2238 (O_2238,N_29920,N_29960);
or UO_2239 (O_2239,N_29645,N_29834);
nor UO_2240 (O_2240,N_29738,N_29535);
and UO_2241 (O_2241,N_29841,N_29937);
or UO_2242 (O_2242,N_29615,N_29879);
nor UO_2243 (O_2243,N_29816,N_29951);
nand UO_2244 (O_2244,N_29863,N_29538);
or UO_2245 (O_2245,N_29697,N_29587);
nor UO_2246 (O_2246,N_29738,N_29611);
and UO_2247 (O_2247,N_29785,N_29565);
xor UO_2248 (O_2248,N_29994,N_29953);
or UO_2249 (O_2249,N_29544,N_29628);
nor UO_2250 (O_2250,N_29589,N_29591);
or UO_2251 (O_2251,N_29753,N_29842);
or UO_2252 (O_2252,N_29837,N_29722);
xnor UO_2253 (O_2253,N_29733,N_29677);
nor UO_2254 (O_2254,N_29668,N_29904);
and UO_2255 (O_2255,N_29609,N_29578);
and UO_2256 (O_2256,N_29692,N_29910);
nor UO_2257 (O_2257,N_29906,N_29567);
xnor UO_2258 (O_2258,N_29976,N_29962);
xnor UO_2259 (O_2259,N_29921,N_29966);
xor UO_2260 (O_2260,N_29525,N_29685);
xnor UO_2261 (O_2261,N_29774,N_29992);
nor UO_2262 (O_2262,N_29992,N_29516);
nor UO_2263 (O_2263,N_29531,N_29555);
and UO_2264 (O_2264,N_29556,N_29687);
nor UO_2265 (O_2265,N_29843,N_29595);
nand UO_2266 (O_2266,N_29830,N_29763);
nor UO_2267 (O_2267,N_29645,N_29727);
and UO_2268 (O_2268,N_29556,N_29716);
xnor UO_2269 (O_2269,N_29854,N_29513);
nor UO_2270 (O_2270,N_29802,N_29553);
nand UO_2271 (O_2271,N_29873,N_29788);
nor UO_2272 (O_2272,N_29595,N_29642);
nor UO_2273 (O_2273,N_29650,N_29832);
or UO_2274 (O_2274,N_29908,N_29549);
and UO_2275 (O_2275,N_29931,N_29950);
nand UO_2276 (O_2276,N_29923,N_29826);
and UO_2277 (O_2277,N_29521,N_29867);
nor UO_2278 (O_2278,N_29911,N_29547);
or UO_2279 (O_2279,N_29945,N_29551);
or UO_2280 (O_2280,N_29642,N_29924);
nand UO_2281 (O_2281,N_29513,N_29875);
or UO_2282 (O_2282,N_29895,N_29966);
nand UO_2283 (O_2283,N_29598,N_29710);
xor UO_2284 (O_2284,N_29727,N_29525);
xor UO_2285 (O_2285,N_29889,N_29619);
xor UO_2286 (O_2286,N_29887,N_29934);
nand UO_2287 (O_2287,N_29619,N_29780);
and UO_2288 (O_2288,N_29748,N_29687);
nand UO_2289 (O_2289,N_29859,N_29928);
and UO_2290 (O_2290,N_29875,N_29935);
or UO_2291 (O_2291,N_29769,N_29995);
nor UO_2292 (O_2292,N_29715,N_29532);
nor UO_2293 (O_2293,N_29635,N_29794);
xor UO_2294 (O_2294,N_29698,N_29570);
xor UO_2295 (O_2295,N_29900,N_29640);
or UO_2296 (O_2296,N_29644,N_29587);
nor UO_2297 (O_2297,N_29843,N_29692);
and UO_2298 (O_2298,N_29544,N_29809);
nor UO_2299 (O_2299,N_29743,N_29906);
nand UO_2300 (O_2300,N_29970,N_29688);
and UO_2301 (O_2301,N_29663,N_29637);
or UO_2302 (O_2302,N_29756,N_29555);
nand UO_2303 (O_2303,N_29810,N_29623);
or UO_2304 (O_2304,N_29884,N_29932);
xnor UO_2305 (O_2305,N_29866,N_29923);
and UO_2306 (O_2306,N_29677,N_29841);
nand UO_2307 (O_2307,N_29766,N_29955);
xor UO_2308 (O_2308,N_29596,N_29656);
and UO_2309 (O_2309,N_29929,N_29969);
xor UO_2310 (O_2310,N_29784,N_29788);
xor UO_2311 (O_2311,N_29757,N_29741);
nand UO_2312 (O_2312,N_29528,N_29798);
nand UO_2313 (O_2313,N_29707,N_29547);
and UO_2314 (O_2314,N_29795,N_29853);
nor UO_2315 (O_2315,N_29836,N_29731);
or UO_2316 (O_2316,N_29724,N_29858);
xor UO_2317 (O_2317,N_29796,N_29844);
nand UO_2318 (O_2318,N_29526,N_29583);
and UO_2319 (O_2319,N_29928,N_29594);
or UO_2320 (O_2320,N_29762,N_29534);
nor UO_2321 (O_2321,N_29880,N_29688);
and UO_2322 (O_2322,N_29725,N_29727);
and UO_2323 (O_2323,N_29747,N_29505);
or UO_2324 (O_2324,N_29773,N_29979);
nand UO_2325 (O_2325,N_29843,N_29891);
and UO_2326 (O_2326,N_29868,N_29519);
nor UO_2327 (O_2327,N_29571,N_29676);
and UO_2328 (O_2328,N_29599,N_29675);
or UO_2329 (O_2329,N_29708,N_29639);
nand UO_2330 (O_2330,N_29897,N_29675);
xor UO_2331 (O_2331,N_29743,N_29857);
nor UO_2332 (O_2332,N_29526,N_29698);
and UO_2333 (O_2333,N_29762,N_29884);
xnor UO_2334 (O_2334,N_29727,N_29634);
xor UO_2335 (O_2335,N_29890,N_29666);
nand UO_2336 (O_2336,N_29632,N_29770);
and UO_2337 (O_2337,N_29575,N_29893);
nor UO_2338 (O_2338,N_29613,N_29888);
or UO_2339 (O_2339,N_29768,N_29924);
xnor UO_2340 (O_2340,N_29611,N_29927);
xnor UO_2341 (O_2341,N_29943,N_29829);
xor UO_2342 (O_2342,N_29779,N_29955);
or UO_2343 (O_2343,N_29957,N_29893);
or UO_2344 (O_2344,N_29917,N_29867);
nand UO_2345 (O_2345,N_29911,N_29821);
nand UO_2346 (O_2346,N_29787,N_29691);
or UO_2347 (O_2347,N_29718,N_29714);
xor UO_2348 (O_2348,N_29710,N_29799);
or UO_2349 (O_2349,N_29650,N_29924);
nor UO_2350 (O_2350,N_29892,N_29744);
or UO_2351 (O_2351,N_29783,N_29699);
xor UO_2352 (O_2352,N_29877,N_29624);
or UO_2353 (O_2353,N_29534,N_29749);
nor UO_2354 (O_2354,N_29611,N_29725);
and UO_2355 (O_2355,N_29708,N_29900);
or UO_2356 (O_2356,N_29782,N_29520);
nand UO_2357 (O_2357,N_29697,N_29871);
nand UO_2358 (O_2358,N_29863,N_29946);
and UO_2359 (O_2359,N_29845,N_29950);
nor UO_2360 (O_2360,N_29747,N_29928);
or UO_2361 (O_2361,N_29808,N_29752);
or UO_2362 (O_2362,N_29542,N_29799);
nand UO_2363 (O_2363,N_29881,N_29675);
and UO_2364 (O_2364,N_29785,N_29793);
and UO_2365 (O_2365,N_29730,N_29830);
xor UO_2366 (O_2366,N_29950,N_29592);
or UO_2367 (O_2367,N_29543,N_29910);
or UO_2368 (O_2368,N_29957,N_29826);
nand UO_2369 (O_2369,N_29651,N_29666);
nand UO_2370 (O_2370,N_29714,N_29778);
xnor UO_2371 (O_2371,N_29935,N_29835);
nor UO_2372 (O_2372,N_29701,N_29661);
nand UO_2373 (O_2373,N_29848,N_29512);
xnor UO_2374 (O_2374,N_29598,N_29887);
xnor UO_2375 (O_2375,N_29886,N_29890);
and UO_2376 (O_2376,N_29597,N_29969);
xor UO_2377 (O_2377,N_29735,N_29793);
or UO_2378 (O_2378,N_29924,N_29581);
or UO_2379 (O_2379,N_29777,N_29550);
xnor UO_2380 (O_2380,N_29649,N_29871);
and UO_2381 (O_2381,N_29697,N_29848);
nor UO_2382 (O_2382,N_29537,N_29591);
or UO_2383 (O_2383,N_29875,N_29980);
or UO_2384 (O_2384,N_29733,N_29845);
and UO_2385 (O_2385,N_29743,N_29741);
xor UO_2386 (O_2386,N_29860,N_29699);
xnor UO_2387 (O_2387,N_29685,N_29884);
and UO_2388 (O_2388,N_29853,N_29659);
xnor UO_2389 (O_2389,N_29843,N_29787);
nand UO_2390 (O_2390,N_29547,N_29691);
and UO_2391 (O_2391,N_29765,N_29754);
or UO_2392 (O_2392,N_29853,N_29532);
xor UO_2393 (O_2393,N_29903,N_29918);
and UO_2394 (O_2394,N_29816,N_29620);
nor UO_2395 (O_2395,N_29830,N_29863);
and UO_2396 (O_2396,N_29679,N_29846);
and UO_2397 (O_2397,N_29909,N_29967);
or UO_2398 (O_2398,N_29886,N_29803);
nor UO_2399 (O_2399,N_29918,N_29980);
nor UO_2400 (O_2400,N_29699,N_29670);
xor UO_2401 (O_2401,N_29844,N_29993);
or UO_2402 (O_2402,N_29864,N_29947);
or UO_2403 (O_2403,N_29921,N_29750);
nand UO_2404 (O_2404,N_29960,N_29628);
nand UO_2405 (O_2405,N_29994,N_29501);
and UO_2406 (O_2406,N_29704,N_29611);
nand UO_2407 (O_2407,N_29768,N_29628);
or UO_2408 (O_2408,N_29900,N_29719);
xnor UO_2409 (O_2409,N_29668,N_29561);
or UO_2410 (O_2410,N_29955,N_29544);
nor UO_2411 (O_2411,N_29559,N_29999);
xnor UO_2412 (O_2412,N_29774,N_29722);
nor UO_2413 (O_2413,N_29538,N_29894);
xor UO_2414 (O_2414,N_29762,N_29664);
or UO_2415 (O_2415,N_29881,N_29625);
nor UO_2416 (O_2416,N_29825,N_29856);
and UO_2417 (O_2417,N_29930,N_29918);
nand UO_2418 (O_2418,N_29670,N_29614);
and UO_2419 (O_2419,N_29861,N_29952);
or UO_2420 (O_2420,N_29728,N_29761);
or UO_2421 (O_2421,N_29659,N_29633);
xor UO_2422 (O_2422,N_29683,N_29840);
nand UO_2423 (O_2423,N_29795,N_29531);
nor UO_2424 (O_2424,N_29641,N_29832);
nand UO_2425 (O_2425,N_29674,N_29716);
nand UO_2426 (O_2426,N_29871,N_29657);
nor UO_2427 (O_2427,N_29970,N_29840);
xnor UO_2428 (O_2428,N_29810,N_29910);
nor UO_2429 (O_2429,N_29664,N_29628);
nor UO_2430 (O_2430,N_29905,N_29591);
or UO_2431 (O_2431,N_29736,N_29937);
nor UO_2432 (O_2432,N_29957,N_29698);
nor UO_2433 (O_2433,N_29925,N_29730);
or UO_2434 (O_2434,N_29916,N_29817);
xnor UO_2435 (O_2435,N_29770,N_29664);
xor UO_2436 (O_2436,N_29764,N_29581);
xnor UO_2437 (O_2437,N_29669,N_29672);
nand UO_2438 (O_2438,N_29795,N_29607);
xor UO_2439 (O_2439,N_29925,N_29774);
nor UO_2440 (O_2440,N_29505,N_29944);
xnor UO_2441 (O_2441,N_29858,N_29941);
xor UO_2442 (O_2442,N_29720,N_29896);
nand UO_2443 (O_2443,N_29619,N_29895);
xor UO_2444 (O_2444,N_29856,N_29672);
nor UO_2445 (O_2445,N_29500,N_29960);
xnor UO_2446 (O_2446,N_29657,N_29649);
or UO_2447 (O_2447,N_29784,N_29597);
or UO_2448 (O_2448,N_29508,N_29947);
and UO_2449 (O_2449,N_29706,N_29669);
or UO_2450 (O_2450,N_29710,N_29954);
nor UO_2451 (O_2451,N_29512,N_29732);
xor UO_2452 (O_2452,N_29902,N_29850);
and UO_2453 (O_2453,N_29799,N_29914);
nor UO_2454 (O_2454,N_29794,N_29528);
and UO_2455 (O_2455,N_29554,N_29904);
nand UO_2456 (O_2456,N_29867,N_29681);
nor UO_2457 (O_2457,N_29787,N_29624);
and UO_2458 (O_2458,N_29517,N_29824);
xnor UO_2459 (O_2459,N_29989,N_29829);
and UO_2460 (O_2460,N_29785,N_29856);
nor UO_2461 (O_2461,N_29614,N_29623);
nor UO_2462 (O_2462,N_29774,N_29826);
and UO_2463 (O_2463,N_29929,N_29696);
nor UO_2464 (O_2464,N_29539,N_29555);
or UO_2465 (O_2465,N_29728,N_29891);
nand UO_2466 (O_2466,N_29871,N_29981);
or UO_2467 (O_2467,N_29898,N_29690);
nand UO_2468 (O_2468,N_29867,N_29644);
and UO_2469 (O_2469,N_29785,N_29834);
and UO_2470 (O_2470,N_29577,N_29686);
and UO_2471 (O_2471,N_29733,N_29802);
nor UO_2472 (O_2472,N_29788,N_29584);
nor UO_2473 (O_2473,N_29702,N_29836);
xnor UO_2474 (O_2474,N_29780,N_29663);
nand UO_2475 (O_2475,N_29858,N_29920);
nand UO_2476 (O_2476,N_29869,N_29915);
xor UO_2477 (O_2477,N_29851,N_29892);
and UO_2478 (O_2478,N_29961,N_29920);
nor UO_2479 (O_2479,N_29718,N_29693);
and UO_2480 (O_2480,N_29647,N_29928);
nor UO_2481 (O_2481,N_29925,N_29583);
nor UO_2482 (O_2482,N_29803,N_29710);
or UO_2483 (O_2483,N_29928,N_29561);
nand UO_2484 (O_2484,N_29821,N_29692);
nand UO_2485 (O_2485,N_29659,N_29752);
or UO_2486 (O_2486,N_29647,N_29521);
nand UO_2487 (O_2487,N_29913,N_29522);
xnor UO_2488 (O_2488,N_29678,N_29750);
nand UO_2489 (O_2489,N_29845,N_29906);
nor UO_2490 (O_2490,N_29888,N_29569);
or UO_2491 (O_2491,N_29501,N_29705);
nor UO_2492 (O_2492,N_29799,N_29753);
and UO_2493 (O_2493,N_29966,N_29862);
or UO_2494 (O_2494,N_29960,N_29923);
nor UO_2495 (O_2495,N_29657,N_29879);
nor UO_2496 (O_2496,N_29741,N_29657);
nand UO_2497 (O_2497,N_29872,N_29611);
and UO_2498 (O_2498,N_29774,N_29797);
or UO_2499 (O_2499,N_29948,N_29859);
xnor UO_2500 (O_2500,N_29788,N_29910);
xor UO_2501 (O_2501,N_29892,N_29791);
xnor UO_2502 (O_2502,N_29640,N_29938);
xnor UO_2503 (O_2503,N_29640,N_29953);
nor UO_2504 (O_2504,N_29588,N_29616);
nor UO_2505 (O_2505,N_29563,N_29673);
and UO_2506 (O_2506,N_29828,N_29724);
nor UO_2507 (O_2507,N_29721,N_29835);
and UO_2508 (O_2508,N_29561,N_29766);
and UO_2509 (O_2509,N_29808,N_29883);
or UO_2510 (O_2510,N_29555,N_29915);
and UO_2511 (O_2511,N_29617,N_29649);
nor UO_2512 (O_2512,N_29681,N_29928);
or UO_2513 (O_2513,N_29944,N_29658);
and UO_2514 (O_2514,N_29745,N_29579);
nor UO_2515 (O_2515,N_29988,N_29910);
and UO_2516 (O_2516,N_29823,N_29631);
nor UO_2517 (O_2517,N_29742,N_29732);
nor UO_2518 (O_2518,N_29563,N_29833);
xor UO_2519 (O_2519,N_29570,N_29883);
nand UO_2520 (O_2520,N_29979,N_29556);
nor UO_2521 (O_2521,N_29795,N_29874);
xnor UO_2522 (O_2522,N_29800,N_29546);
nand UO_2523 (O_2523,N_29951,N_29632);
nand UO_2524 (O_2524,N_29683,N_29632);
nor UO_2525 (O_2525,N_29717,N_29838);
nor UO_2526 (O_2526,N_29972,N_29773);
xnor UO_2527 (O_2527,N_29892,N_29529);
nor UO_2528 (O_2528,N_29635,N_29551);
or UO_2529 (O_2529,N_29731,N_29933);
nand UO_2530 (O_2530,N_29894,N_29833);
xor UO_2531 (O_2531,N_29897,N_29931);
xor UO_2532 (O_2532,N_29981,N_29787);
nor UO_2533 (O_2533,N_29852,N_29740);
nand UO_2534 (O_2534,N_29817,N_29953);
nand UO_2535 (O_2535,N_29976,N_29865);
or UO_2536 (O_2536,N_29756,N_29829);
nor UO_2537 (O_2537,N_29914,N_29993);
nand UO_2538 (O_2538,N_29983,N_29955);
xnor UO_2539 (O_2539,N_29579,N_29787);
nand UO_2540 (O_2540,N_29774,N_29663);
and UO_2541 (O_2541,N_29967,N_29777);
xor UO_2542 (O_2542,N_29515,N_29650);
xor UO_2543 (O_2543,N_29560,N_29989);
and UO_2544 (O_2544,N_29968,N_29710);
and UO_2545 (O_2545,N_29542,N_29788);
or UO_2546 (O_2546,N_29855,N_29861);
and UO_2547 (O_2547,N_29708,N_29989);
nor UO_2548 (O_2548,N_29950,N_29690);
or UO_2549 (O_2549,N_29543,N_29691);
and UO_2550 (O_2550,N_29645,N_29912);
nor UO_2551 (O_2551,N_29954,N_29575);
nand UO_2552 (O_2552,N_29771,N_29690);
and UO_2553 (O_2553,N_29802,N_29770);
nor UO_2554 (O_2554,N_29636,N_29626);
nor UO_2555 (O_2555,N_29868,N_29695);
and UO_2556 (O_2556,N_29836,N_29877);
nand UO_2557 (O_2557,N_29972,N_29665);
or UO_2558 (O_2558,N_29886,N_29712);
xnor UO_2559 (O_2559,N_29876,N_29534);
xnor UO_2560 (O_2560,N_29917,N_29697);
and UO_2561 (O_2561,N_29909,N_29851);
nor UO_2562 (O_2562,N_29568,N_29882);
xor UO_2563 (O_2563,N_29941,N_29507);
nor UO_2564 (O_2564,N_29583,N_29534);
xnor UO_2565 (O_2565,N_29835,N_29822);
or UO_2566 (O_2566,N_29619,N_29956);
xnor UO_2567 (O_2567,N_29973,N_29754);
xor UO_2568 (O_2568,N_29853,N_29911);
nor UO_2569 (O_2569,N_29509,N_29710);
nor UO_2570 (O_2570,N_29540,N_29512);
xor UO_2571 (O_2571,N_29979,N_29780);
nand UO_2572 (O_2572,N_29616,N_29599);
nor UO_2573 (O_2573,N_29628,N_29567);
nand UO_2574 (O_2574,N_29692,N_29903);
nor UO_2575 (O_2575,N_29763,N_29636);
nor UO_2576 (O_2576,N_29918,N_29539);
nor UO_2577 (O_2577,N_29885,N_29523);
and UO_2578 (O_2578,N_29777,N_29944);
nor UO_2579 (O_2579,N_29513,N_29865);
or UO_2580 (O_2580,N_29891,N_29947);
and UO_2581 (O_2581,N_29673,N_29904);
xor UO_2582 (O_2582,N_29664,N_29865);
nor UO_2583 (O_2583,N_29869,N_29854);
nand UO_2584 (O_2584,N_29566,N_29553);
nor UO_2585 (O_2585,N_29777,N_29560);
or UO_2586 (O_2586,N_29848,N_29536);
nand UO_2587 (O_2587,N_29854,N_29672);
nand UO_2588 (O_2588,N_29915,N_29628);
and UO_2589 (O_2589,N_29545,N_29688);
and UO_2590 (O_2590,N_29881,N_29679);
xnor UO_2591 (O_2591,N_29629,N_29699);
xor UO_2592 (O_2592,N_29706,N_29830);
xnor UO_2593 (O_2593,N_29740,N_29645);
or UO_2594 (O_2594,N_29811,N_29720);
nand UO_2595 (O_2595,N_29880,N_29718);
nor UO_2596 (O_2596,N_29739,N_29912);
nand UO_2597 (O_2597,N_29886,N_29873);
nand UO_2598 (O_2598,N_29504,N_29594);
nand UO_2599 (O_2599,N_29927,N_29848);
or UO_2600 (O_2600,N_29898,N_29988);
nor UO_2601 (O_2601,N_29889,N_29665);
or UO_2602 (O_2602,N_29988,N_29573);
nor UO_2603 (O_2603,N_29786,N_29672);
nand UO_2604 (O_2604,N_29971,N_29928);
nor UO_2605 (O_2605,N_29816,N_29933);
or UO_2606 (O_2606,N_29736,N_29618);
or UO_2607 (O_2607,N_29558,N_29649);
nor UO_2608 (O_2608,N_29686,N_29850);
nand UO_2609 (O_2609,N_29516,N_29713);
and UO_2610 (O_2610,N_29700,N_29766);
xnor UO_2611 (O_2611,N_29646,N_29957);
nand UO_2612 (O_2612,N_29574,N_29957);
and UO_2613 (O_2613,N_29649,N_29943);
and UO_2614 (O_2614,N_29515,N_29717);
xnor UO_2615 (O_2615,N_29908,N_29873);
nor UO_2616 (O_2616,N_29900,N_29529);
and UO_2617 (O_2617,N_29657,N_29754);
or UO_2618 (O_2618,N_29985,N_29509);
or UO_2619 (O_2619,N_29658,N_29575);
or UO_2620 (O_2620,N_29738,N_29694);
or UO_2621 (O_2621,N_29859,N_29522);
xnor UO_2622 (O_2622,N_29554,N_29741);
nand UO_2623 (O_2623,N_29890,N_29756);
or UO_2624 (O_2624,N_29559,N_29636);
nand UO_2625 (O_2625,N_29933,N_29764);
nor UO_2626 (O_2626,N_29637,N_29700);
and UO_2627 (O_2627,N_29574,N_29876);
and UO_2628 (O_2628,N_29521,N_29646);
nor UO_2629 (O_2629,N_29922,N_29790);
nor UO_2630 (O_2630,N_29849,N_29818);
nor UO_2631 (O_2631,N_29801,N_29993);
xor UO_2632 (O_2632,N_29969,N_29971);
or UO_2633 (O_2633,N_29593,N_29537);
nor UO_2634 (O_2634,N_29948,N_29683);
xor UO_2635 (O_2635,N_29812,N_29569);
nor UO_2636 (O_2636,N_29737,N_29728);
nor UO_2637 (O_2637,N_29980,N_29708);
and UO_2638 (O_2638,N_29916,N_29641);
nand UO_2639 (O_2639,N_29853,N_29714);
nand UO_2640 (O_2640,N_29577,N_29537);
and UO_2641 (O_2641,N_29955,N_29504);
or UO_2642 (O_2642,N_29586,N_29757);
nor UO_2643 (O_2643,N_29825,N_29501);
and UO_2644 (O_2644,N_29710,N_29845);
xor UO_2645 (O_2645,N_29738,N_29733);
nor UO_2646 (O_2646,N_29916,N_29818);
or UO_2647 (O_2647,N_29991,N_29909);
and UO_2648 (O_2648,N_29621,N_29909);
and UO_2649 (O_2649,N_29649,N_29594);
nand UO_2650 (O_2650,N_29539,N_29526);
xnor UO_2651 (O_2651,N_29973,N_29812);
and UO_2652 (O_2652,N_29883,N_29525);
and UO_2653 (O_2653,N_29542,N_29749);
or UO_2654 (O_2654,N_29726,N_29979);
and UO_2655 (O_2655,N_29747,N_29669);
and UO_2656 (O_2656,N_29853,N_29678);
and UO_2657 (O_2657,N_29675,N_29754);
nand UO_2658 (O_2658,N_29916,N_29538);
nand UO_2659 (O_2659,N_29618,N_29902);
nand UO_2660 (O_2660,N_29606,N_29814);
or UO_2661 (O_2661,N_29649,N_29989);
nand UO_2662 (O_2662,N_29914,N_29699);
xnor UO_2663 (O_2663,N_29735,N_29557);
or UO_2664 (O_2664,N_29819,N_29670);
nor UO_2665 (O_2665,N_29800,N_29880);
nor UO_2666 (O_2666,N_29668,N_29984);
or UO_2667 (O_2667,N_29724,N_29609);
xnor UO_2668 (O_2668,N_29993,N_29988);
xor UO_2669 (O_2669,N_29839,N_29799);
nor UO_2670 (O_2670,N_29538,N_29727);
or UO_2671 (O_2671,N_29539,N_29639);
or UO_2672 (O_2672,N_29525,N_29804);
xor UO_2673 (O_2673,N_29719,N_29546);
nor UO_2674 (O_2674,N_29953,N_29711);
nand UO_2675 (O_2675,N_29698,N_29851);
nand UO_2676 (O_2676,N_29604,N_29746);
nand UO_2677 (O_2677,N_29951,N_29841);
or UO_2678 (O_2678,N_29933,N_29716);
or UO_2679 (O_2679,N_29860,N_29707);
and UO_2680 (O_2680,N_29611,N_29974);
xor UO_2681 (O_2681,N_29839,N_29990);
nand UO_2682 (O_2682,N_29794,N_29660);
or UO_2683 (O_2683,N_29850,N_29508);
nand UO_2684 (O_2684,N_29610,N_29824);
xnor UO_2685 (O_2685,N_29692,N_29815);
nor UO_2686 (O_2686,N_29784,N_29604);
nor UO_2687 (O_2687,N_29540,N_29645);
nand UO_2688 (O_2688,N_29943,N_29810);
or UO_2689 (O_2689,N_29773,N_29686);
and UO_2690 (O_2690,N_29740,N_29832);
nand UO_2691 (O_2691,N_29964,N_29922);
nand UO_2692 (O_2692,N_29828,N_29950);
or UO_2693 (O_2693,N_29652,N_29523);
nor UO_2694 (O_2694,N_29700,N_29802);
and UO_2695 (O_2695,N_29961,N_29621);
nor UO_2696 (O_2696,N_29644,N_29999);
xor UO_2697 (O_2697,N_29666,N_29563);
nand UO_2698 (O_2698,N_29904,N_29607);
or UO_2699 (O_2699,N_29622,N_29618);
nand UO_2700 (O_2700,N_29882,N_29783);
nand UO_2701 (O_2701,N_29789,N_29733);
or UO_2702 (O_2702,N_29527,N_29738);
or UO_2703 (O_2703,N_29629,N_29642);
or UO_2704 (O_2704,N_29927,N_29888);
or UO_2705 (O_2705,N_29794,N_29719);
nand UO_2706 (O_2706,N_29707,N_29985);
nand UO_2707 (O_2707,N_29773,N_29594);
or UO_2708 (O_2708,N_29898,N_29553);
nand UO_2709 (O_2709,N_29798,N_29724);
and UO_2710 (O_2710,N_29658,N_29759);
nor UO_2711 (O_2711,N_29863,N_29760);
nor UO_2712 (O_2712,N_29648,N_29772);
xor UO_2713 (O_2713,N_29534,N_29911);
nand UO_2714 (O_2714,N_29696,N_29599);
and UO_2715 (O_2715,N_29966,N_29679);
and UO_2716 (O_2716,N_29969,N_29917);
or UO_2717 (O_2717,N_29919,N_29914);
nand UO_2718 (O_2718,N_29684,N_29721);
xnor UO_2719 (O_2719,N_29746,N_29797);
and UO_2720 (O_2720,N_29694,N_29750);
or UO_2721 (O_2721,N_29782,N_29534);
nand UO_2722 (O_2722,N_29708,N_29823);
nand UO_2723 (O_2723,N_29791,N_29698);
nor UO_2724 (O_2724,N_29544,N_29733);
xor UO_2725 (O_2725,N_29545,N_29590);
and UO_2726 (O_2726,N_29732,N_29640);
or UO_2727 (O_2727,N_29926,N_29742);
or UO_2728 (O_2728,N_29959,N_29840);
nor UO_2729 (O_2729,N_29541,N_29900);
nand UO_2730 (O_2730,N_29672,N_29568);
nor UO_2731 (O_2731,N_29641,N_29737);
or UO_2732 (O_2732,N_29573,N_29939);
and UO_2733 (O_2733,N_29761,N_29506);
and UO_2734 (O_2734,N_29712,N_29745);
xnor UO_2735 (O_2735,N_29837,N_29930);
nand UO_2736 (O_2736,N_29649,N_29914);
or UO_2737 (O_2737,N_29730,N_29841);
or UO_2738 (O_2738,N_29732,N_29628);
or UO_2739 (O_2739,N_29750,N_29656);
nand UO_2740 (O_2740,N_29502,N_29964);
nand UO_2741 (O_2741,N_29900,N_29795);
nand UO_2742 (O_2742,N_29902,N_29937);
and UO_2743 (O_2743,N_29652,N_29619);
or UO_2744 (O_2744,N_29766,N_29717);
xnor UO_2745 (O_2745,N_29807,N_29606);
and UO_2746 (O_2746,N_29777,N_29902);
nand UO_2747 (O_2747,N_29663,N_29986);
nor UO_2748 (O_2748,N_29712,N_29837);
and UO_2749 (O_2749,N_29637,N_29628);
nor UO_2750 (O_2750,N_29592,N_29751);
nand UO_2751 (O_2751,N_29931,N_29849);
xnor UO_2752 (O_2752,N_29902,N_29892);
xor UO_2753 (O_2753,N_29793,N_29675);
xnor UO_2754 (O_2754,N_29688,N_29709);
and UO_2755 (O_2755,N_29554,N_29977);
nand UO_2756 (O_2756,N_29603,N_29537);
xnor UO_2757 (O_2757,N_29868,N_29558);
xor UO_2758 (O_2758,N_29921,N_29844);
nor UO_2759 (O_2759,N_29841,N_29755);
xnor UO_2760 (O_2760,N_29995,N_29795);
nand UO_2761 (O_2761,N_29976,N_29761);
and UO_2762 (O_2762,N_29972,N_29983);
nor UO_2763 (O_2763,N_29636,N_29711);
and UO_2764 (O_2764,N_29560,N_29529);
and UO_2765 (O_2765,N_29597,N_29644);
nand UO_2766 (O_2766,N_29852,N_29525);
or UO_2767 (O_2767,N_29779,N_29857);
nor UO_2768 (O_2768,N_29901,N_29545);
nor UO_2769 (O_2769,N_29749,N_29575);
and UO_2770 (O_2770,N_29831,N_29966);
or UO_2771 (O_2771,N_29636,N_29754);
or UO_2772 (O_2772,N_29617,N_29980);
and UO_2773 (O_2773,N_29985,N_29569);
xnor UO_2774 (O_2774,N_29873,N_29779);
and UO_2775 (O_2775,N_29804,N_29655);
nor UO_2776 (O_2776,N_29700,N_29906);
and UO_2777 (O_2777,N_29526,N_29524);
xor UO_2778 (O_2778,N_29517,N_29756);
xor UO_2779 (O_2779,N_29530,N_29775);
xor UO_2780 (O_2780,N_29656,N_29743);
nand UO_2781 (O_2781,N_29889,N_29850);
nand UO_2782 (O_2782,N_29957,N_29693);
nand UO_2783 (O_2783,N_29514,N_29830);
and UO_2784 (O_2784,N_29688,N_29867);
and UO_2785 (O_2785,N_29820,N_29772);
and UO_2786 (O_2786,N_29943,N_29694);
nand UO_2787 (O_2787,N_29783,N_29541);
and UO_2788 (O_2788,N_29750,N_29967);
or UO_2789 (O_2789,N_29632,N_29852);
or UO_2790 (O_2790,N_29885,N_29573);
nand UO_2791 (O_2791,N_29603,N_29577);
and UO_2792 (O_2792,N_29795,N_29791);
and UO_2793 (O_2793,N_29895,N_29814);
nor UO_2794 (O_2794,N_29814,N_29620);
nor UO_2795 (O_2795,N_29611,N_29547);
and UO_2796 (O_2796,N_29955,N_29826);
nand UO_2797 (O_2797,N_29686,N_29942);
and UO_2798 (O_2798,N_29789,N_29619);
and UO_2799 (O_2799,N_29878,N_29557);
nor UO_2800 (O_2800,N_29909,N_29879);
and UO_2801 (O_2801,N_29974,N_29522);
xor UO_2802 (O_2802,N_29542,N_29847);
nand UO_2803 (O_2803,N_29995,N_29541);
nand UO_2804 (O_2804,N_29719,N_29886);
xor UO_2805 (O_2805,N_29676,N_29930);
or UO_2806 (O_2806,N_29751,N_29583);
or UO_2807 (O_2807,N_29635,N_29799);
and UO_2808 (O_2808,N_29807,N_29690);
and UO_2809 (O_2809,N_29806,N_29576);
nand UO_2810 (O_2810,N_29923,N_29952);
and UO_2811 (O_2811,N_29756,N_29738);
or UO_2812 (O_2812,N_29799,N_29516);
xor UO_2813 (O_2813,N_29636,N_29528);
and UO_2814 (O_2814,N_29920,N_29964);
or UO_2815 (O_2815,N_29586,N_29596);
xor UO_2816 (O_2816,N_29826,N_29518);
nor UO_2817 (O_2817,N_29991,N_29813);
nand UO_2818 (O_2818,N_29645,N_29875);
nand UO_2819 (O_2819,N_29605,N_29816);
xor UO_2820 (O_2820,N_29820,N_29746);
and UO_2821 (O_2821,N_29761,N_29586);
nand UO_2822 (O_2822,N_29920,N_29790);
nor UO_2823 (O_2823,N_29818,N_29640);
nor UO_2824 (O_2824,N_29641,N_29835);
nor UO_2825 (O_2825,N_29680,N_29704);
nor UO_2826 (O_2826,N_29803,N_29938);
xor UO_2827 (O_2827,N_29621,N_29586);
and UO_2828 (O_2828,N_29776,N_29833);
and UO_2829 (O_2829,N_29720,N_29672);
or UO_2830 (O_2830,N_29731,N_29823);
and UO_2831 (O_2831,N_29694,N_29642);
nor UO_2832 (O_2832,N_29803,N_29724);
and UO_2833 (O_2833,N_29505,N_29864);
nor UO_2834 (O_2834,N_29780,N_29840);
xor UO_2835 (O_2835,N_29570,N_29795);
or UO_2836 (O_2836,N_29909,N_29985);
nor UO_2837 (O_2837,N_29545,N_29841);
nor UO_2838 (O_2838,N_29505,N_29769);
nand UO_2839 (O_2839,N_29991,N_29834);
or UO_2840 (O_2840,N_29644,N_29643);
or UO_2841 (O_2841,N_29635,N_29554);
and UO_2842 (O_2842,N_29510,N_29717);
xnor UO_2843 (O_2843,N_29791,N_29711);
or UO_2844 (O_2844,N_29897,N_29937);
and UO_2845 (O_2845,N_29672,N_29875);
xor UO_2846 (O_2846,N_29773,N_29576);
nand UO_2847 (O_2847,N_29659,N_29916);
xnor UO_2848 (O_2848,N_29605,N_29735);
nand UO_2849 (O_2849,N_29826,N_29992);
nand UO_2850 (O_2850,N_29964,N_29825);
xnor UO_2851 (O_2851,N_29759,N_29863);
or UO_2852 (O_2852,N_29865,N_29644);
xnor UO_2853 (O_2853,N_29982,N_29969);
and UO_2854 (O_2854,N_29976,N_29588);
xor UO_2855 (O_2855,N_29661,N_29907);
nor UO_2856 (O_2856,N_29662,N_29663);
and UO_2857 (O_2857,N_29548,N_29947);
nor UO_2858 (O_2858,N_29950,N_29746);
or UO_2859 (O_2859,N_29779,N_29625);
or UO_2860 (O_2860,N_29869,N_29733);
nand UO_2861 (O_2861,N_29808,N_29845);
nor UO_2862 (O_2862,N_29674,N_29661);
xnor UO_2863 (O_2863,N_29920,N_29590);
xnor UO_2864 (O_2864,N_29986,N_29667);
and UO_2865 (O_2865,N_29680,N_29526);
and UO_2866 (O_2866,N_29620,N_29600);
nor UO_2867 (O_2867,N_29521,N_29941);
xor UO_2868 (O_2868,N_29785,N_29838);
or UO_2869 (O_2869,N_29566,N_29774);
nand UO_2870 (O_2870,N_29878,N_29889);
and UO_2871 (O_2871,N_29973,N_29637);
or UO_2872 (O_2872,N_29681,N_29834);
nor UO_2873 (O_2873,N_29698,N_29721);
xnor UO_2874 (O_2874,N_29630,N_29972);
xnor UO_2875 (O_2875,N_29850,N_29528);
or UO_2876 (O_2876,N_29648,N_29993);
and UO_2877 (O_2877,N_29661,N_29685);
xor UO_2878 (O_2878,N_29932,N_29735);
nand UO_2879 (O_2879,N_29946,N_29654);
nor UO_2880 (O_2880,N_29616,N_29552);
and UO_2881 (O_2881,N_29901,N_29799);
nand UO_2882 (O_2882,N_29650,N_29741);
nand UO_2883 (O_2883,N_29981,N_29951);
nand UO_2884 (O_2884,N_29750,N_29699);
xor UO_2885 (O_2885,N_29618,N_29919);
xnor UO_2886 (O_2886,N_29760,N_29882);
xor UO_2887 (O_2887,N_29605,N_29685);
xor UO_2888 (O_2888,N_29730,N_29923);
nor UO_2889 (O_2889,N_29663,N_29911);
or UO_2890 (O_2890,N_29772,N_29963);
and UO_2891 (O_2891,N_29771,N_29746);
xnor UO_2892 (O_2892,N_29913,N_29752);
nor UO_2893 (O_2893,N_29942,N_29793);
or UO_2894 (O_2894,N_29959,N_29953);
nand UO_2895 (O_2895,N_29775,N_29747);
or UO_2896 (O_2896,N_29874,N_29547);
nand UO_2897 (O_2897,N_29666,N_29834);
nand UO_2898 (O_2898,N_29589,N_29507);
nand UO_2899 (O_2899,N_29806,N_29923);
and UO_2900 (O_2900,N_29594,N_29968);
and UO_2901 (O_2901,N_29878,N_29858);
nor UO_2902 (O_2902,N_29618,N_29527);
nand UO_2903 (O_2903,N_29677,N_29912);
nor UO_2904 (O_2904,N_29553,N_29933);
or UO_2905 (O_2905,N_29528,N_29598);
xnor UO_2906 (O_2906,N_29594,N_29765);
xor UO_2907 (O_2907,N_29541,N_29576);
or UO_2908 (O_2908,N_29782,N_29993);
and UO_2909 (O_2909,N_29596,N_29676);
or UO_2910 (O_2910,N_29605,N_29769);
nand UO_2911 (O_2911,N_29641,N_29839);
nand UO_2912 (O_2912,N_29801,N_29533);
xnor UO_2913 (O_2913,N_29555,N_29744);
nor UO_2914 (O_2914,N_29655,N_29637);
nand UO_2915 (O_2915,N_29691,N_29931);
xnor UO_2916 (O_2916,N_29532,N_29744);
nor UO_2917 (O_2917,N_29532,N_29711);
xnor UO_2918 (O_2918,N_29578,N_29636);
and UO_2919 (O_2919,N_29970,N_29636);
or UO_2920 (O_2920,N_29744,N_29953);
or UO_2921 (O_2921,N_29566,N_29962);
and UO_2922 (O_2922,N_29906,N_29752);
nor UO_2923 (O_2923,N_29501,N_29528);
nand UO_2924 (O_2924,N_29629,N_29607);
or UO_2925 (O_2925,N_29976,N_29997);
or UO_2926 (O_2926,N_29985,N_29516);
and UO_2927 (O_2927,N_29706,N_29620);
and UO_2928 (O_2928,N_29558,N_29627);
or UO_2929 (O_2929,N_29969,N_29904);
xor UO_2930 (O_2930,N_29787,N_29962);
xor UO_2931 (O_2931,N_29940,N_29726);
xor UO_2932 (O_2932,N_29971,N_29836);
xnor UO_2933 (O_2933,N_29913,N_29576);
and UO_2934 (O_2934,N_29503,N_29704);
xnor UO_2935 (O_2935,N_29918,N_29550);
xor UO_2936 (O_2936,N_29504,N_29745);
nand UO_2937 (O_2937,N_29867,N_29880);
nand UO_2938 (O_2938,N_29966,N_29704);
xor UO_2939 (O_2939,N_29676,N_29976);
nor UO_2940 (O_2940,N_29679,N_29706);
xor UO_2941 (O_2941,N_29839,N_29975);
or UO_2942 (O_2942,N_29863,N_29970);
or UO_2943 (O_2943,N_29877,N_29694);
and UO_2944 (O_2944,N_29651,N_29721);
or UO_2945 (O_2945,N_29701,N_29886);
or UO_2946 (O_2946,N_29818,N_29564);
nand UO_2947 (O_2947,N_29501,N_29556);
and UO_2948 (O_2948,N_29515,N_29860);
or UO_2949 (O_2949,N_29667,N_29644);
nand UO_2950 (O_2950,N_29656,N_29675);
nor UO_2951 (O_2951,N_29950,N_29664);
nand UO_2952 (O_2952,N_29989,N_29611);
or UO_2953 (O_2953,N_29959,N_29773);
or UO_2954 (O_2954,N_29509,N_29922);
xnor UO_2955 (O_2955,N_29989,N_29561);
nor UO_2956 (O_2956,N_29787,N_29963);
nor UO_2957 (O_2957,N_29700,N_29981);
nor UO_2958 (O_2958,N_29970,N_29928);
xor UO_2959 (O_2959,N_29939,N_29576);
nand UO_2960 (O_2960,N_29662,N_29715);
or UO_2961 (O_2961,N_29670,N_29682);
xor UO_2962 (O_2962,N_29706,N_29503);
and UO_2963 (O_2963,N_29763,N_29904);
xnor UO_2964 (O_2964,N_29541,N_29550);
nor UO_2965 (O_2965,N_29746,N_29693);
xor UO_2966 (O_2966,N_29989,N_29625);
and UO_2967 (O_2967,N_29792,N_29502);
or UO_2968 (O_2968,N_29702,N_29820);
xor UO_2969 (O_2969,N_29896,N_29933);
xnor UO_2970 (O_2970,N_29727,N_29574);
nand UO_2971 (O_2971,N_29518,N_29990);
nand UO_2972 (O_2972,N_29866,N_29947);
and UO_2973 (O_2973,N_29512,N_29586);
and UO_2974 (O_2974,N_29527,N_29924);
nor UO_2975 (O_2975,N_29708,N_29727);
xor UO_2976 (O_2976,N_29592,N_29711);
nor UO_2977 (O_2977,N_29852,N_29556);
xnor UO_2978 (O_2978,N_29696,N_29758);
and UO_2979 (O_2979,N_29881,N_29910);
and UO_2980 (O_2980,N_29574,N_29828);
nor UO_2981 (O_2981,N_29720,N_29799);
nand UO_2982 (O_2982,N_29575,N_29714);
xor UO_2983 (O_2983,N_29791,N_29776);
nor UO_2984 (O_2984,N_29810,N_29645);
and UO_2985 (O_2985,N_29584,N_29913);
nand UO_2986 (O_2986,N_29989,N_29916);
and UO_2987 (O_2987,N_29918,N_29809);
and UO_2988 (O_2988,N_29962,N_29771);
and UO_2989 (O_2989,N_29710,N_29684);
nand UO_2990 (O_2990,N_29595,N_29937);
or UO_2991 (O_2991,N_29667,N_29905);
or UO_2992 (O_2992,N_29809,N_29843);
and UO_2993 (O_2993,N_29616,N_29784);
nand UO_2994 (O_2994,N_29727,N_29717);
nor UO_2995 (O_2995,N_29922,N_29568);
nand UO_2996 (O_2996,N_29513,N_29767);
or UO_2997 (O_2997,N_29935,N_29517);
or UO_2998 (O_2998,N_29738,N_29600);
nor UO_2999 (O_2999,N_29665,N_29656);
nand UO_3000 (O_3000,N_29918,N_29887);
xor UO_3001 (O_3001,N_29869,N_29902);
xor UO_3002 (O_3002,N_29603,N_29591);
and UO_3003 (O_3003,N_29812,N_29653);
xnor UO_3004 (O_3004,N_29722,N_29574);
nand UO_3005 (O_3005,N_29689,N_29685);
nor UO_3006 (O_3006,N_29851,N_29754);
xor UO_3007 (O_3007,N_29502,N_29970);
nor UO_3008 (O_3008,N_29973,N_29614);
nand UO_3009 (O_3009,N_29759,N_29987);
nor UO_3010 (O_3010,N_29800,N_29663);
or UO_3011 (O_3011,N_29830,N_29809);
nand UO_3012 (O_3012,N_29993,N_29518);
nand UO_3013 (O_3013,N_29936,N_29838);
or UO_3014 (O_3014,N_29856,N_29908);
and UO_3015 (O_3015,N_29943,N_29847);
nor UO_3016 (O_3016,N_29667,N_29648);
xnor UO_3017 (O_3017,N_29736,N_29770);
and UO_3018 (O_3018,N_29701,N_29732);
nor UO_3019 (O_3019,N_29881,N_29842);
xor UO_3020 (O_3020,N_29854,N_29587);
or UO_3021 (O_3021,N_29934,N_29905);
xor UO_3022 (O_3022,N_29980,N_29778);
or UO_3023 (O_3023,N_29896,N_29986);
and UO_3024 (O_3024,N_29801,N_29785);
xnor UO_3025 (O_3025,N_29681,N_29528);
xnor UO_3026 (O_3026,N_29685,N_29744);
or UO_3027 (O_3027,N_29541,N_29516);
xor UO_3028 (O_3028,N_29998,N_29702);
or UO_3029 (O_3029,N_29696,N_29618);
or UO_3030 (O_3030,N_29737,N_29566);
and UO_3031 (O_3031,N_29526,N_29545);
nand UO_3032 (O_3032,N_29707,N_29515);
or UO_3033 (O_3033,N_29945,N_29838);
nand UO_3034 (O_3034,N_29819,N_29750);
xnor UO_3035 (O_3035,N_29647,N_29739);
nor UO_3036 (O_3036,N_29741,N_29524);
nand UO_3037 (O_3037,N_29754,N_29799);
nor UO_3038 (O_3038,N_29995,N_29762);
and UO_3039 (O_3039,N_29813,N_29924);
nand UO_3040 (O_3040,N_29599,N_29540);
and UO_3041 (O_3041,N_29538,N_29918);
and UO_3042 (O_3042,N_29538,N_29503);
or UO_3043 (O_3043,N_29780,N_29512);
nor UO_3044 (O_3044,N_29511,N_29570);
and UO_3045 (O_3045,N_29710,N_29615);
and UO_3046 (O_3046,N_29786,N_29823);
nand UO_3047 (O_3047,N_29504,N_29760);
xor UO_3048 (O_3048,N_29760,N_29768);
or UO_3049 (O_3049,N_29711,N_29527);
and UO_3050 (O_3050,N_29929,N_29648);
nand UO_3051 (O_3051,N_29963,N_29524);
or UO_3052 (O_3052,N_29613,N_29906);
xnor UO_3053 (O_3053,N_29697,N_29695);
or UO_3054 (O_3054,N_29937,N_29506);
nor UO_3055 (O_3055,N_29926,N_29852);
xnor UO_3056 (O_3056,N_29876,N_29937);
nand UO_3057 (O_3057,N_29687,N_29698);
nor UO_3058 (O_3058,N_29722,N_29684);
and UO_3059 (O_3059,N_29739,N_29993);
and UO_3060 (O_3060,N_29868,N_29832);
xnor UO_3061 (O_3061,N_29805,N_29862);
xnor UO_3062 (O_3062,N_29703,N_29721);
and UO_3063 (O_3063,N_29999,N_29540);
or UO_3064 (O_3064,N_29814,N_29592);
nor UO_3065 (O_3065,N_29688,N_29560);
and UO_3066 (O_3066,N_29762,N_29794);
and UO_3067 (O_3067,N_29738,N_29896);
xor UO_3068 (O_3068,N_29907,N_29569);
xor UO_3069 (O_3069,N_29739,N_29672);
xnor UO_3070 (O_3070,N_29944,N_29682);
nor UO_3071 (O_3071,N_29514,N_29643);
nor UO_3072 (O_3072,N_29627,N_29702);
or UO_3073 (O_3073,N_29835,N_29518);
nor UO_3074 (O_3074,N_29886,N_29716);
nor UO_3075 (O_3075,N_29637,N_29837);
or UO_3076 (O_3076,N_29926,N_29578);
xnor UO_3077 (O_3077,N_29973,N_29645);
nor UO_3078 (O_3078,N_29551,N_29670);
or UO_3079 (O_3079,N_29823,N_29812);
xnor UO_3080 (O_3080,N_29842,N_29566);
and UO_3081 (O_3081,N_29971,N_29739);
and UO_3082 (O_3082,N_29668,N_29935);
and UO_3083 (O_3083,N_29636,N_29886);
and UO_3084 (O_3084,N_29724,N_29540);
and UO_3085 (O_3085,N_29755,N_29950);
and UO_3086 (O_3086,N_29724,N_29642);
and UO_3087 (O_3087,N_29500,N_29887);
xnor UO_3088 (O_3088,N_29647,N_29792);
nor UO_3089 (O_3089,N_29736,N_29895);
nand UO_3090 (O_3090,N_29637,N_29917);
or UO_3091 (O_3091,N_29949,N_29566);
xor UO_3092 (O_3092,N_29614,N_29781);
and UO_3093 (O_3093,N_29558,N_29751);
and UO_3094 (O_3094,N_29957,N_29640);
nand UO_3095 (O_3095,N_29827,N_29726);
nand UO_3096 (O_3096,N_29755,N_29550);
or UO_3097 (O_3097,N_29963,N_29730);
or UO_3098 (O_3098,N_29679,N_29994);
xnor UO_3099 (O_3099,N_29750,N_29792);
xor UO_3100 (O_3100,N_29887,N_29564);
or UO_3101 (O_3101,N_29667,N_29557);
nand UO_3102 (O_3102,N_29923,N_29832);
nand UO_3103 (O_3103,N_29923,N_29872);
nand UO_3104 (O_3104,N_29602,N_29922);
or UO_3105 (O_3105,N_29946,N_29761);
nor UO_3106 (O_3106,N_29803,N_29502);
nor UO_3107 (O_3107,N_29655,N_29806);
xnor UO_3108 (O_3108,N_29523,N_29515);
xor UO_3109 (O_3109,N_29922,N_29705);
or UO_3110 (O_3110,N_29833,N_29880);
xnor UO_3111 (O_3111,N_29871,N_29576);
xnor UO_3112 (O_3112,N_29966,N_29682);
nand UO_3113 (O_3113,N_29772,N_29928);
or UO_3114 (O_3114,N_29862,N_29935);
and UO_3115 (O_3115,N_29597,N_29869);
xnor UO_3116 (O_3116,N_29915,N_29870);
or UO_3117 (O_3117,N_29563,N_29827);
and UO_3118 (O_3118,N_29871,N_29811);
or UO_3119 (O_3119,N_29878,N_29928);
and UO_3120 (O_3120,N_29529,N_29535);
xnor UO_3121 (O_3121,N_29967,N_29928);
nand UO_3122 (O_3122,N_29835,N_29875);
nor UO_3123 (O_3123,N_29580,N_29899);
nor UO_3124 (O_3124,N_29877,N_29763);
xnor UO_3125 (O_3125,N_29529,N_29964);
xnor UO_3126 (O_3126,N_29669,N_29909);
or UO_3127 (O_3127,N_29512,N_29576);
or UO_3128 (O_3128,N_29681,N_29973);
or UO_3129 (O_3129,N_29514,N_29980);
nor UO_3130 (O_3130,N_29865,N_29642);
nor UO_3131 (O_3131,N_29655,N_29607);
and UO_3132 (O_3132,N_29696,N_29595);
xnor UO_3133 (O_3133,N_29806,N_29636);
and UO_3134 (O_3134,N_29537,N_29699);
nand UO_3135 (O_3135,N_29589,N_29931);
nor UO_3136 (O_3136,N_29792,N_29763);
nand UO_3137 (O_3137,N_29923,N_29594);
nor UO_3138 (O_3138,N_29818,N_29553);
and UO_3139 (O_3139,N_29823,N_29500);
and UO_3140 (O_3140,N_29803,N_29904);
xor UO_3141 (O_3141,N_29886,N_29571);
nor UO_3142 (O_3142,N_29703,N_29841);
xnor UO_3143 (O_3143,N_29648,N_29777);
and UO_3144 (O_3144,N_29802,N_29728);
or UO_3145 (O_3145,N_29821,N_29666);
or UO_3146 (O_3146,N_29856,N_29567);
nor UO_3147 (O_3147,N_29892,N_29900);
or UO_3148 (O_3148,N_29647,N_29900);
xnor UO_3149 (O_3149,N_29992,N_29703);
xor UO_3150 (O_3150,N_29760,N_29971);
or UO_3151 (O_3151,N_29935,N_29978);
and UO_3152 (O_3152,N_29619,N_29697);
or UO_3153 (O_3153,N_29800,N_29737);
nand UO_3154 (O_3154,N_29517,N_29648);
xor UO_3155 (O_3155,N_29736,N_29688);
nand UO_3156 (O_3156,N_29779,N_29899);
or UO_3157 (O_3157,N_29659,N_29526);
or UO_3158 (O_3158,N_29518,N_29808);
xor UO_3159 (O_3159,N_29930,N_29546);
nand UO_3160 (O_3160,N_29802,N_29905);
nand UO_3161 (O_3161,N_29547,N_29972);
xor UO_3162 (O_3162,N_29544,N_29562);
xor UO_3163 (O_3163,N_29942,N_29825);
xnor UO_3164 (O_3164,N_29850,N_29958);
and UO_3165 (O_3165,N_29747,N_29626);
nor UO_3166 (O_3166,N_29695,N_29545);
or UO_3167 (O_3167,N_29624,N_29687);
xnor UO_3168 (O_3168,N_29832,N_29582);
and UO_3169 (O_3169,N_29528,N_29888);
nor UO_3170 (O_3170,N_29634,N_29973);
nand UO_3171 (O_3171,N_29689,N_29732);
xnor UO_3172 (O_3172,N_29663,N_29521);
nand UO_3173 (O_3173,N_29658,N_29621);
nand UO_3174 (O_3174,N_29687,N_29514);
nor UO_3175 (O_3175,N_29542,N_29504);
nand UO_3176 (O_3176,N_29788,N_29848);
xnor UO_3177 (O_3177,N_29720,N_29709);
nor UO_3178 (O_3178,N_29636,N_29516);
nand UO_3179 (O_3179,N_29819,N_29913);
xor UO_3180 (O_3180,N_29730,N_29533);
xor UO_3181 (O_3181,N_29730,N_29735);
and UO_3182 (O_3182,N_29509,N_29863);
nor UO_3183 (O_3183,N_29951,N_29649);
nand UO_3184 (O_3184,N_29647,N_29656);
xor UO_3185 (O_3185,N_29961,N_29560);
and UO_3186 (O_3186,N_29651,N_29583);
or UO_3187 (O_3187,N_29873,N_29587);
nor UO_3188 (O_3188,N_29589,N_29818);
nand UO_3189 (O_3189,N_29836,N_29760);
and UO_3190 (O_3190,N_29644,N_29547);
nor UO_3191 (O_3191,N_29984,N_29943);
nor UO_3192 (O_3192,N_29924,N_29708);
nand UO_3193 (O_3193,N_29671,N_29562);
xnor UO_3194 (O_3194,N_29544,N_29521);
and UO_3195 (O_3195,N_29782,N_29849);
or UO_3196 (O_3196,N_29780,N_29565);
nand UO_3197 (O_3197,N_29773,N_29980);
xnor UO_3198 (O_3198,N_29743,N_29507);
nand UO_3199 (O_3199,N_29752,N_29728);
nor UO_3200 (O_3200,N_29607,N_29909);
or UO_3201 (O_3201,N_29997,N_29712);
nand UO_3202 (O_3202,N_29950,N_29693);
xor UO_3203 (O_3203,N_29735,N_29996);
nor UO_3204 (O_3204,N_29885,N_29711);
xor UO_3205 (O_3205,N_29785,N_29649);
xnor UO_3206 (O_3206,N_29555,N_29573);
nand UO_3207 (O_3207,N_29585,N_29667);
nand UO_3208 (O_3208,N_29869,N_29575);
or UO_3209 (O_3209,N_29644,N_29562);
nand UO_3210 (O_3210,N_29964,N_29636);
xor UO_3211 (O_3211,N_29640,N_29567);
nor UO_3212 (O_3212,N_29860,N_29811);
xor UO_3213 (O_3213,N_29860,N_29575);
nand UO_3214 (O_3214,N_29666,N_29559);
xnor UO_3215 (O_3215,N_29718,N_29874);
xnor UO_3216 (O_3216,N_29864,N_29809);
nor UO_3217 (O_3217,N_29959,N_29779);
or UO_3218 (O_3218,N_29849,N_29666);
xor UO_3219 (O_3219,N_29749,N_29869);
nor UO_3220 (O_3220,N_29728,N_29995);
nand UO_3221 (O_3221,N_29936,N_29939);
xnor UO_3222 (O_3222,N_29987,N_29681);
xnor UO_3223 (O_3223,N_29748,N_29547);
nor UO_3224 (O_3224,N_29792,N_29894);
xor UO_3225 (O_3225,N_29901,N_29511);
xor UO_3226 (O_3226,N_29983,N_29945);
and UO_3227 (O_3227,N_29523,N_29781);
and UO_3228 (O_3228,N_29985,N_29631);
or UO_3229 (O_3229,N_29529,N_29815);
xnor UO_3230 (O_3230,N_29724,N_29971);
or UO_3231 (O_3231,N_29878,N_29896);
and UO_3232 (O_3232,N_29684,N_29803);
or UO_3233 (O_3233,N_29728,N_29875);
nand UO_3234 (O_3234,N_29614,N_29592);
and UO_3235 (O_3235,N_29938,N_29837);
nand UO_3236 (O_3236,N_29948,N_29893);
nor UO_3237 (O_3237,N_29749,N_29985);
nand UO_3238 (O_3238,N_29927,N_29756);
nand UO_3239 (O_3239,N_29719,N_29585);
or UO_3240 (O_3240,N_29621,N_29851);
and UO_3241 (O_3241,N_29570,N_29744);
nand UO_3242 (O_3242,N_29682,N_29601);
and UO_3243 (O_3243,N_29584,N_29552);
or UO_3244 (O_3244,N_29525,N_29897);
nand UO_3245 (O_3245,N_29682,N_29535);
and UO_3246 (O_3246,N_29963,N_29731);
nand UO_3247 (O_3247,N_29904,N_29559);
or UO_3248 (O_3248,N_29632,N_29847);
and UO_3249 (O_3249,N_29580,N_29804);
and UO_3250 (O_3250,N_29568,N_29767);
and UO_3251 (O_3251,N_29595,N_29877);
nor UO_3252 (O_3252,N_29933,N_29769);
xnor UO_3253 (O_3253,N_29745,N_29513);
or UO_3254 (O_3254,N_29599,N_29876);
nor UO_3255 (O_3255,N_29876,N_29767);
nor UO_3256 (O_3256,N_29809,N_29623);
nor UO_3257 (O_3257,N_29862,N_29856);
nor UO_3258 (O_3258,N_29734,N_29780);
nand UO_3259 (O_3259,N_29903,N_29969);
or UO_3260 (O_3260,N_29859,N_29828);
and UO_3261 (O_3261,N_29749,N_29947);
xnor UO_3262 (O_3262,N_29800,N_29664);
nor UO_3263 (O_3263,N_29515,N_29775);
nor UO_3264 (O_3264,N_29845,N_29597);
or UO_3265 (O_3265,N_29991,N_29752);
or UO_3266 (O_3266,N_29774,N_29642);
or UO_3267 (O_3267,N_29559,N_29775);
nand UO_3268 (O_3268,N_29952,N_29837);
xor UO_3269 (O_3269,N_29838,N_29503);
or UO_3270 (O_3270,N_29840,N_29895);
xor UO_3271 (O_3271,N_29583,N_29967);
or UO_3272 (O_3272,N_29865,N_29725);
nor UO_3273 (O_3273,N_29629,N_29704);
or UO_3274 (O_3274,N_29914,N_29753);
xor UO_3275 (O_3275,N_29819,N_29781);
or UO_3276 (O_3276,N_29502,N_29598);
xnor UO_3277 (O_3277,N_29545,N_29685);
xor UO_3278 (O_3278,N_29614,N_29585);
nand UO_3279 (O_3279,N_29741,N_29862);
and UO_3280 (O_3280,N_29938,N_29548);
and UO_3281 (O_3281,N_29743,N_29930);
xor UO_3282 (O_3282,N_29740,N_29760);
nor UO_3283 (O_3283,N_29535,N_29526);
or UO_3284 (O_3284,N_29692,N_29528);
and UO_3285 (O_3285,N_29893,N_29719);
nand UO_3286 (O_3286,N_29543,N_29935);
nand UO_3287 (O_3287,N_29662,N_29768);
xnor UO_3288 (O_3288,N_29968,N_29892);
nor UO_3289 (O_3289,N_29598,N_29980);
and UO_3290 (O_3290,N_29990,N_29776);
and UO_3291 (O_3291,N_29771,N_29689);
and UO_3292 (O_3292,N_29915,N_29862);
nand UO_3293 (O_3293,N_29675,N_29785);
and UO_3294 (O_3294,N_29696,N_29751);
and UO_3295 (O_3295,N_29974,N_29536);
or UO_3296 (O_3296,N_29801,N_29765);
or UO_3297 (O_3297,N_29837,N_29728);
xor UO_3298 (O_3298,N_29613,N_29580);
nor UO_3299 (O_3299,N_29782,N_29784);
xor UO_3300 (O_3300,N_29910,N_29966);
nor UO_3301 (O_3301,N_29879,N_29960);
or UO_3302 (O_3302,N_29940,N_29570);
or UO_3303 (O_3303,N_29668,N_29980);
nand UO_3304 (O_3304,N_29955,N_29720);
or UO_3305 (O_3305,N_29709,N_29677);
xor UO_3306 (O_3306,N_29622,N_29586);
xnor UO_3307 (O_3307,N_29882,N_29644);
and UO_3308 (O_3308,N_29840,N_29665);
or UO_3309 (O_3309,N_29831,N_29809);
nand UO_3310 (O_3310,N_29792,N_29517);
and UO_3311 (O_3311,N_29523,N_29915);
or UO_3312 (O_3312,N_29613,N_29742);
nor UO_3313 (O_3313,N_29644,N_29894);
xnor UO_3314 (O_3314,N_29925,N_29554);
xor UO_3315 (O_3315,N_29756,N_29812);
or UO_3316 (O_3316,N_29825,N_29991);
and UO_3317 (O_3317,N_29800,N_29944);
or UO_3318 (O_3318,N_29784,N_29893);
nand UO_3319 (O_3319,N_29766,N_29801);
and UO_3320 (O_3320,N_29716,N_29732);
nand UO_3321 (O_3321,N_29937,N_29659);
xnor UO_3322 (O_3322,N_29640,N_29591);
nand UO_3323 (O_3323,N_29881,N_29867);
or UO_3324 (O_3324,N_29732,N_29877);
nor UO_3325 (O_3325,N_29517,N_29993);
xor UO_3326 (O_3326,N_29826,N_29884);
nand UO_3327 (O_3327,N_29736,N_29700);
nand UO_3328 (O_3328,N_29507,N_29966);
and UO_3329 (O_3329,N_29568,N_29795);
and UO_3330 (O_3330,N_29713,N_29782);
xor UO_3331 (O_3331,N_29605,N_29784);
or UO_3332 (O_3332,N_29747,N_29511);
nand UO_3333 (O_3333,N_29545,N_29630);
xnor UO_3334 (O_3334,N_29663,N_29548);
and UO_3335 (O_3335,N_29766,N_29518);
xor UO_3336 (O_3336,N_29798,N_29885);
nor UO_3337 (O_3337,N_29583,N_29900);
xnor UO_3338 (O_3338,N_29946,N_29670);
nand UO_3339 (O_3339,N_29923,N_29865);
nand UO_3340 (O_3340,N_29800,N_29828);
nor UO_3341 (O_3341,N_29704,N_29738);
or UO_3342 (O_3342,N_29737,N_29844);
xnor UO_3343 (O_3343,N_29658,N_29538);
nand UO_3344 (O_3344,N_29732,N_29797);
xor UO_3345 (O_3345,N_29964,N_29786);
or UO_3346 (O_3346,N_29925,N_29803);
or UO_3347 (O_3347,N_29536,N_29701);
nor UO_3348 (O_3348,N_29662,N_29580);
nor UO_3349 (O_3349,N_29698,N_29741);
or UO_3350 (O_3350,N_29599,N_29703);
nand UO_3351 (O_3351,N_29540,N_29908);
xor UO_3352 (O_3352,N_29617,N_29553);
nand UO_3353 (O_3353,N_29797,N_29650);
and UO_3354 (O_3354,N_29803,N_29926);
xnor UO_3355 (O_3355,N_29607,N_29754);
xnor UO_3356 (O_3356,N_29557,N_29517);
and UO_3357 (O_3357,N_29672,N_29593);
and UO_3358 (O_3358,N_29684,N_29895);
nor UO_3359 (O_3359,N_29649,N_29505);
and UO_3360 (O_3360,N_29574,N_29596);
and UO_3361 (O_3361,N_29972,N_29636);
xor UO_3362 (O_3362,N_29556,N_29574);
or UO_3363 (O_3363,N_29667,N_29877);
or UO_3364 (O_3364,N_29866,N_29920);
xnor UO_3365 (O_3365,N_29857,N_29797);
nand UO_3366 (O_3366,N_29601,N_29820);
xnor UO_3367 (O_3367,N_29806,N_29957);
nor UO_3368 (O_3368,N_29607,N_29810);
and UO_3369 (O_3369,N_29763,N_29694);
nand UO_3370 (O_3370,N_29920,N_29634);
nor UO_3371 (O_3371,N_29673,N_29663);
nand UO_3372 (O_3372,N_29644,N_29905);
nand UO_3373 (O_3373,N_29853,N_29809);
xor UO_3374 (O_3374,N_29649,N_29996);
nor UO_3375 (O_3375,N_29974,N_29599);
nand UO_3376 (O_3376,N_29935,N_29912);
and UO_3377 (O_3377,N_29588,N_29918);
xnor UO_3378 (O_3378,N_29821,N_29930);
nand UO_3379 (O_3379,N_29852,N_29686);
and UO_3380 (O_3380,N_29635,N_29522);
and UO_3381 (O_3381,N_29742,N_29773);
or UO_3382 (O_3382,N_29639,N_29851);
or UO_3383 (O_3383,N_29619,N_29807);
xnor UO_3384 (O_3384,N_29943,N_29632);
and UO_3385 (O_3385,N_29622,N_29580);
or UO_3386 (O_3386,N_29765,N_29753);
nor UO_3387 (O_3387,N_29651,N_29726);
or UO_3388 (O_3388,N_29532,N_29736);
nor UO_3389 (O_3389,N_29941,N_29689);
and UO_3390 (O_3390,N_29667,N_29501);
nand UO_3391 (O_3391,N_29869,N_29580);
nor UO_3392 (O_3392,N_29512,N_29571);
xnor UO_3393 (O_3393,N_29925,N_29763);
or UO_3394 (O_3394,N_29981,N_29935);
xor UO_3395 (O_3395,N_29981,N_29558);
nor UO_3396 (O_3396,N_29860,N_29636);
xor UO_3397 (O_3397,N_29678,N_29964);
xor UO_3398 (O_3398,N_29989,N_29812);
nand UO_3399 (O_3399,N_29697,N_29919);
xor UO_3400 (O_3400,N_29648,N_29719);
xor UO_3401 (O_3401,N_29601,N_29766);
nor UO_3402 (O_3402,N_29828,N_29797);
xnor UO_3403 (O_3403,N_29841,N_29885);
nand UO_3404 (O_3404,N_29621,N_29885);
and UO_3405 (O_3405,N_29789,N_29740);
and UO_3406 (O_3406,N_29710,N_29716);
nor UO_3407 (O_3407,N_29564,N_29747);
or UO_3408 (O_3408,N_29911,N_29995);
nor UO_3409 (O_3409,N_29957,N_29625);
nor UO_3410 (O_3410,N_29909,N_29796);
or UO_3411 (O_3411,N_29915,N_29894);
nor UO_3412 (O_3412,N_29818,N_29820);
xor UO_3413 (O_3413,N_29559,N_29968);
or UO_3414 (O_3414,N_29500,N_29820);
xnor UO_3415 (O_3415,N_29779,N_29549);
nor UO_3416 (O_3416,N_29942,N_29817);
xnor UO_3417 (O_3417,N_29931,N_29663);
or UO_3418 (O_3418,N_29687,N_29664);
nand UO_3419 (O_3419,N_29572,N_29673);
or UO_3420 (O_3420,N_29756,N_29546);
and UO_3421 (O_3421,N_29586,N_29741);
xor UO_3422 (O_3422,N_29541,N_29819);
or UO_3423 (O_3423,N_29892,N_29828);
and UO_3424 (O_3424,N_29504,N_29735);
nand UO_3425 (O_3425,N_29941,N_29606);
and UO_3426 (O_3426,N_29776,N_29524);
xor UO_3427 (O_3427,N_29882,N_29554);
nand UO_3428 (O_3428,N_29865,N_29769);
or UO_3429 (O_3429,N_29547,N_29677);
xnor UO_3430 (O_3430,N_29684,N_29711);
xor UO_3431 (O_3431,N_29922,N_29552);
or UO_3432 (O_3432,N_29977,N_29850);
nor UO_3433 (O_3433,N_29817,N_29693);
or UO_3434 (O_3434,N_29950,N_29607);
or UO_3435 (O_3435,N_29948,N_29735);
or UO_3436 (O_3436,N_29661,N_29960);
nand UO_3437 (O_3437,N_29860,N_29967);
or UO_3438 (O_3438,N_29681,N_29620);
or UO_3439 (O_3439,N_29699,N_29649);
xnor UO_3440 (O_3440,N_29545,N_29635);
nand UO_3441 (O_3441,N_29819,N_29528);
or UO_3442 (O_3442,N_29785,N_29762);
nand UO_3443 (O_3443,N_29674,N_29653);
xnor UO_3444 (O_3444,N_29607,N_29960);
nand UO_3445 (O_3445,N_29611,N_29579);
nor UO_3446 (O_3446,N_29686,N_29659);
and UO_3447 (O_3447,N_29598,N_29960);
or UO_3448 (O_3448,N_29587,N_29872);
or UO_3449 (O_3449,N_29961,N_29549);
nand UO_3450 (O_3450,N_29808,N_29664);
xor UO_3451 (O_3451,N_29937,N_29927);
xnor UO_3452 (O_3452,N_29723,N_29870);
xor UO_3453 (O_3453,N_29864,N_29893);
or UO_3454 (O_3454,N_29581,N_29685);
and UO_3455 (O_3455,N_29855,N_29841);
nand UO_3456 (O_3456,N_29747,N_29627);
nand UO_3457 (O_3457,N_29881,N_29816);
and UO_3458 (O_3458,N_29734,N_29980);
nand UO_3459 (O_3459,N_29569,N_29659);
and UO_3460 (O_3460,N_29837,N_29736);
and UO_3461 (O_3461,N_29969,N_29838);
nand UO_3462 (O_3462,N_29840,N_29875);
xor UO_3463 (O_3463,N_29693,N_29600);
and UO_3464 (O_3464,N_29791,N_29748);
and UO_3465 (O_3465,N_29900,N_29761);
or UO_3466 (O_3466,N_29621,N_29603);
or UO_3467 (O_3467,N_29687,N_29852);
nand UO_3468 (O_3468,N_29924,N_29829);
nor UO_3469 (O_3469,N_29696,N_29584);
or UO_3470 (O_3470,N_29860,N_29578);
nand UO_3471 (O_3471,N_29649,N_29901);
or UO_3472 (O_3472,N_29811,N_29748);
nor UO_3473 (O_3473,N_29984,N_29896);
nand UO_3474 (O_3474,N_29664,N_29715);
or UO_3475 (O_3475,N_29646,N_29847);
and UO_3476 (O_3476,N_29906,N_29860);
nor UO_3477 (O_3477,N_29978,N_29567);
or UO_3478 (O_3478,N_29948,N_29644);
or UO_3479 (O_3479,N_29641,N_29553);
nand UO_3480 (O_3480,N_29903,N_29664);
and UO_3481 (O_3481,N_29766,N_29746);
xor UO_3482 (O_3482,N_29534,N_29805);
xor UO_3483 (O_3483,N_29737,N_29993);
xor UO_3484 (O_3484,N_29866,N_29664);
and UO_3485 (O_3485,N_29967,N_29771);
nand UO_3486 (O_3486,N_29924,N_29890);
xnor UO_3487 (O_3487,N_29858,N_29726);
nand UO_3488 (O_3488,N_29743,N_29708);
nor UO_3489 (O_3489,N_29621,N_29732);
nor UO_3490 (O_3490,N_29854,N_29853);
or UO_3491 (O_3491,N_29961,N_29762);
nand UO_3492 (O_3492,N_29709,N_29928);
nand UO_3493 (O_3493,N_29706,N_29811);
xor UO_3494 (O_3494,N_29620,N_29604);
and UO_3495 (O_3495,N_29815,N_29702);
nor UO_3496 (O_3496,N_29983,N_29870);
nand UO_3497 (O_3497,N_29747,N_29986);
nor UO_3498 (O_3498,N_29936,N_29551);
and UO_3499 (O_3499,N_29714,N_29978);
endmodule