module basic_1000_10000_1500_2_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5004,N_5006,N_5007,N_5008,N_5010,N_5011,N_5012,N_5017,N_5019,N_5022,N_5023,N_5024,N_5026,N_5029,N_5030,N_5031,N_5033,N_5034,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5047,N_5048,N_5049,N_5053,N_5054,N_5055,N_5056,N_5057,N_5059,N_5064,N_5065,N_5066,N_5069,N_5070,N_5071,N_5072,N_5074,N_5076,N_5077,N_5078,N_5080,N_5082,N_5083,N_5084,N_5086,N_5088,N_5090,N_5094,N_5095,N_5096,N_5097,N_5100,N_5101,N_5102,N_5103,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5113,N_5115,N_5117,N_5118,N_5119,N_5120,N_5122,N_5123,N_5124,N_5125,N_5127,N_5128,N_5130,N_5131,N_5133,N_5134,N_5136,N_5137,N_5139,N_5140,N_5143,N_5145,N_5146,N_5151,N_5153,N_5156,N_5157,N_5159,N_5162,N_5163,N_5164,N_5166,N_5167,N_5169,N_5173,N_5174,N_5175,N_5177,N_5178,N_5179,N_5182,N_5183,N_5184,N_5188,N_5189,N_5194,N_5195,N_5196,N_5198,N_5199,N_5201,N_5202,N_5203,N_5205,N_5207,N_5208,N_5210,N_5214,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5226,N_5228,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5240,N_5241,N_5242,N_5244,N_5246,N_5247,N_5248,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5259,N_5261,N_5262,N_5263,N_5266,N_5267,N_5268,N_5270,N_5271,N_5273,N_5274,N_5275,N_5280,N_5282,N_5284,N_5285,N_5286,N_5288,N_5291,N_5292,N_5294,N_5295,N_5298,N_5300,N_5302,N_5303,N_5304,N_5306,N_5307,N_5310,N_5311,N_5314,N_5316,N_5317,N_5318,N_5319,N_5320,N_5322,N_5323,N_5324,N_5325,N_5327,N_5329,N_5330,N_5331,N_5333,N_5335,N_5338,N_5339,N_5342,N_5344,N_5346,N_5349,N_5350,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5360,N_5363,N_5364,N_5367,N_5368,N_5370,N_5372,N_5373,N_5374,N_5376,N_5377,N_5378,N_5379,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5390,N_5392,N_5393,N_5394,N_5396,N_5397,N_5399,N_5401,N_5402,N_5403,N_5404,N_5409,N_5411,N_5414,N_5415,N_5417,N_5418,N_5421,N_5428,N_5429,N_5431,N_5434,N_5435,N_5436,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5445,N_5446,N_5448,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5458,N_5459,N_5464,N_5465,N_5466,N_5467,N_5470,N_5471,N_5472,N_5473,N_5474,N_5477,N_5480,N_5481,N_5484,N_5485,N_5486,N_5488,N_5491,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5500,N_5501,N_5502,N_5504,N_5505,N_5506,N_5507,N_5509,N_5512,N_5513,N_5514,N_5518,N_5519,N_5521,N_5522,N_5523,N_5525,N_5528,N_5530,N_5533,N_5534,N_5535,N_5536,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5546,N_5547,N_5548,N_5550,N_5551,N_5552,N_5555,N_5556,N_5557,N_5561,N_5562,N_5566,N_5567,N_5570,N_5571,N_5574,N_5576,N_5577,N_5581,N_5582,N_5583,N_5586,N_5587,N_5588,N_5589,N_5592,N_5594,N_5596,N_5600,N_5601,N_5604,N_5606,N_5610,N_5611,N_5612,N_5614,N_5616,N_5617,N_5618,N_5619,N_5621,N_5622,N_5625,N_5626,N_5628,N_5629,N_5630,N_5632,N_5633,N_5634,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5644,N_5645,N_5646,N_5651,N_5654,N_5655,N_5656,N_5658,N_5659,N_5660,N_5661,N_5664,N_5667,N_5669,N_5670,N_5671,N_5672,N_5675,N_5677,N_5681,N_5683,N_5684,N_5685,N_5687,N_5688,N_5691,N_5692,N_5693,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5705,N_5708,N_5710,N_5714,N_5715,N_5716,N_5718,N_5719,N_5721,N_5723,N_5725,N_5727,N_5729,N_5730,N_5733,N_5736,N_5737,N_5739,N_5740,N_5745,N_5746,N_5748,N_5749,N_5750,N_5753,N_5754,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5766,N_5767,N_5768,N_5770,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5782,N_5783,N_5784,N_5785,N_5790,N_5793,N_5794,N_5798,N_5801,N_5803,N_5807,N_5808,N_5809,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5819,N_5820,N_5821,N_5822,N_5825,N_5826,N_5829,N_5831,N_5832,N_5833,N_5834,N_5838,N_5839,N_5840,N_5842,N_5844,N_5846,N_5847,N_5848,N_5849,N_5853,N_5854,N_5855,N_5857,N_5858,N_5861,N_5863,N_5864,N_5865,N_5867,N_5868,N_5869,N_5870,N_5873,N_5874,N_5876,N_5877,N_5879,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5890,N_5891,N_5893,N_5894,N_5895,N_5900,N_5901,N_5902,N_5904,N_5905,N_5906,N_5907,N_5910,N_5912,N_5914,N_5915,N_5916,N_5917,N_5919,N_5922,N_5924,N_5925,N_5927,N_5928,N_5932,N_5933,N_5934,N_5937,N_5938,N_5941,N_5942,N_5944,N_5945,N_5946,N_5947,N_5948,N_5950,N_5953,N_5954,N_5956,N_5959,N_5960,N_5961,N_5962,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5972,N_5974,N_5975,N_5979,N_5981,N_5982,N_5983,N_5986,N_5987,N_5988,N_5990,N_5992,N_5993,N_5994,N_5997,N_5998,N_5999,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6014,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6027,N_6028,N_6030,N_6031,N_6032,N_6033,N_6035,N_6036,N_6040,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6053,N_6054,N_6055,N_6057,N_6058,N_6060,N_6061,N_6063,N_6065,N_6067,N_6071,N_6072,N_6076,N_6077,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6086,N_6089,N_6092,N_6093,N_6095,N_6097,N_6098,N_6101,N_6103,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6115,N_6116,N_6122,N_6123,N_6125,N_6126,N_6128,N_6130,N_6131,N_6132,N_6133,N_6135,N_6137,N_6139,N_6140,N_6143,N_6144,N_6145,N_6147,N_6148,N_6149,N_6151,N_6153,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6162,N_6166,N_6167,N_6168,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6178,N_6179,N_6182,N_6184,N_6185,N_6186,N_6187,N_6189,N_6190,N_6191,N_6194,N_6195,N_6196,N_6198,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6216,N_6217,N_6219,N_6220,N_6221,N_6223,N_6225,N_6227,N_6230,N_6231,N_6232,N_6233,N_6235,N_6237,N_6238,N_6240,N_6241,N_6242,N_6244,N_6248,N_6250,N_6251,N_6253,N_6254,N_6255,N_6257,N_6263,N_6265,N_6266,N_6268,N_6269,N_6273,N_6274,N_6275,N_6276,N_6277,N_6279,N_6280,N_6281,N_6283,N_6286,N_6287,N_6289,N_6291,N_6293,N_6294,N_6295,N_6296,N_6297,N_6301,N_6303,N_6304,N_6305,N_6306,N_6307,N_6309,N_6310,N_6312,N_6315,N_6316,N_6317,N_6318,N_6319,N_6321,N_6323,N_6324,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6334,N_6336,N_6338,N_6340,N_6342,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6352,N_6353,N_6355,N_6356,N_6357,N_6358,N_6359,N_6363,N_6364,N_6366,N_6367,N_6368,N_6371,N_6374,N_6375,N_6379,N_6383,N_6384,N_6387,N_6390,N_6391,N_6392,N_6394,N_6395,N_6396,N_6398,N_6399,N_6402,N_6405,N_6409,N_6410,N_6415,N_6418,N_6419,N_6420,N_6422,N_6424,N_6425,N_6426,N_6429,N_6430,N_6431,N_6433,N_6435,N_6438,N_6441,N_6442,N_6444,N_6445,N_6446,N_6447,N_6448,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6458,N_6461,N_6462,N_6464,N_6465,N_6466,N_6469,N_6472,N_6474,N_6477,N_6479,N_6483,N_6487,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6506,N_6508,N_6509,N_6510,N_6513,N_6514,N_6515,N_6517,N_6518,N_6519,N_6521,N_6522,N_6523,N_6524,N_6525,N_6527,N_6528,N_6529,N_6530,N_6531,N_6533,N_6535,N_6537,N_6538,N_6539,N_6540,N_6542,N_6544,N_6545,N_6546,N_6547,N_6548,N_6550,N_6551,N_6552,N_6557,N_6561,N_6562,N_6564,N_6568,N_6569,N_6573,N_6574,N_6576,N_6579,N_6580,N_6581,N_6583,N_6585,N_6586,N_6587,N_6589,N_6590,N_6591,N_6592,N_6593,N_6595,N_6596,N_6597,N_6598,N_6601,N_6603,N_6605,N_6607,N_6610,N_6611,N_6612,N_6617,N_6618,N_6619,N_6622,N_6624,N_6626,N_6628,N_6634,N_6636,N_6637,N_6638,N_6639,N_6641,N_6642,N_6644,N_6646,N_6647,N_6648,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6662,N_6665,N_6667,N_6668,N_6669,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6684,N_6688,N_6689,N_6690,N_6693,N_6694,N_6695,N_6696,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6721,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6731,N_6732,N_6733,N_6734,N_6739,N_6742,N_6743,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6756,N_6758,N_6760,N_6761,N_6763,N_6764,N_6765,N_6767,N_6768,N_6769,N_6770,N_6776,N_6777,N_6778,N_6780,N_6781,N_6782,N_6785,N_6786,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6801,N_6803,N_6805,N_6807,N_6809,N_6811,N_6812,N_6813,N_6815,N_6818,N_6822,N_6823,N_6824,N_6825,N_6827,N_6828,N_6829,N_6830,N_6832,N_6834,N_6836,N_6837,N_6838,N_6839,N_6840,N_6843,N_6845,N_6847,N_6849,N_6850,N_6852,N_6853,N_6854,N_6857,N_6858,N_6859,N_6860,N_6861,N_6866,N_6867,N_6868,N_6870,N_6872,N_6873,N_6874,N_6876,N_6878,N_6880,N_6881,N_6884,N_6885,N_6888,N_6891,N_6892,N_6893,N_6895,N_6896,N_6897,N_6898,N_6901,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6910,N_6912,N_6913,N_6914,N_6917,N_6918,N_6919,N_6920,N_6921,N_6923,N_6924,N_6925,N_6929,N_6934,N_6935,N_6936,N_6938,N_6940,N_6947,N_6948,N_6950,N_6952,N_6953,N_6954,N_6957,N_6958,N_6959,N_6961,N_6965,N_6967,N_6971,N_6972,N_6974,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6983,N_6984,N_6985,N_6987,N_6988,N_6989,N_6991,N_6995,N_6997,N_6998,N_7000,N_7002,N_7003,N_7004,N_7005,N_7007,N_7008,N_7009,N_7011,N_7013,N_7014,N_7015,N_7017,N_7019,N_7020,N_7022,N_7023,N_7024,N_7025,N_7028,N_7030,N_7031,N_7032,N_7033,N_7035,N_7036,N_7037,N_7041,N_7043,N_7044,N_7045,N_7046,N_7047,N_7049,N_7050,N_7051,N_7052,N_7054,N_7055,N_7056,N_7057,N_7059,N_7060,N_7061,N_7062,N_7063,N_7065,N_7066,N_7071,N_7072,N_7073,N_7077,N_7078,N_7079,N_7081,N_7083,N_7085,N_7087,N_7088,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7099,N_7100,N_7106,N_7108,N_7109,N_7110,N_7111,N_7112,N_7114,N_7115,N_7117,N_7119,N_7121,N_7122,N_7123,N_7125,N_7127,N_7129,N_7130,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7142,N_7143,N_7144,N_7146,N_7147,N_7148,N_7151,N_7156,N_7157,N_7161,N_7163,N_7165,N_7167,N_7168,N_7169,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7179,N_7180,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7203,N_7205,N_7207,N_7208,N_7211,N_7215,N_7216,N_7217,N_7218,N_7220,N_7221,N_7223,N_7224,N_7226,N_7227,N_7228,N_7229,N_7234,N_7235,N_7239,N_7240,N_7241,N_7245,N_7246,N_7247,N_7249,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7259,N_7260,N_7261,N_7267,N_7269,N_7270,N_7271,N_7273,N_7278,N_7279,N_7280,N_7281,N_7288,N_7289,N_7290,N_7291,N_7292,N_7297,N_7299,N_7300,N_7301,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7316,N_7318,N_7320,N_7323,N_7324,N_7326,N_7327,N_7328,N_7330,N_7331,N_7333,N_7336,N_7339,N_7340,N_7344,N_7345,N_7347,N_7350,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7362,N_7363,N_7365,N_7366,N_7367,N_7368,N_7369,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7382,N_7384,N_7389,N_7390,N_7394,N_7395,N_7396,N_7397,N_7398,N_7400,N_7401,N_7402,N_7403,N_7407,N_7409,N_7412,N_7413,N_7415,N_7417,N_7419,N_7420,N_7422,N_7423,N_7427,N_7433,N_7434,N_7435,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7455,N_7456,N_7458,N_7459,N_7460,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7470,N_7472,N_7474,N_7478,N_7479,N_7480,N_7483,N_7485,N_7486,N_7488,N_7492,N_7493,N_7494,N_7496,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7509,N_7510,N_7513,N_7514,N_7516,N_7517,N_7518,N_7519,N_7520,N_7523,N_7527,N_7528,N_7529,N_7530,N_7531,N_7533,N_7534,N_7537,N_7538,N_7540,N_7542,N_7543,N_7545,N_7548,N_7549,N_7550,N_7551,N_7552,N_7555,N_7557,N_7558,N_7560,N_7563,N_7564,N_7567,N_7568,N_7569,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7583,N_7585,N_7586,N_7588,N_7589,N_7590,N_7593,N_7597,N_7599,N_7600,N_7602,N_7603,N_7604,N_7606,N_7608,N_7610,N_7611,N_7612,N_7613,N_7615,N_7617,N_7619,N_7620,N_7622,N_7624,N_7625,N_7626,N_7628,N_7631,N_7634,N_7635,N_7636,N_7638,N_7639,N_7640,N_7641,N_7642,N_7644,N_7645,N_7646,N_7648,N_7649,N_7650,N_7653,N_7654,N_7655,N_7659,N_7660,N_7661,N_7663,N_7664,N_7665,N_7667,N_7668,N_7669,N_7670,N_7672,N_7675,N_7676,N_7677,N_7679,N_7681,N_7683,N_7684,N_7688,N_7689,N_7690,N_7694,N_7695,N_7696,N_7697,N_7698,N_7700,N_7701,N_7702,N_7703,N_7704,N_7706,N_7708,N_7709,N_7711,N_7715,N_7717,N_7718,N_7719,N_7720,N_7724,N_7725,N_7726,N_7728,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7739,N_7741,N_7742,N_7743,N_7744,N_7745,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7755,N_7756,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7768,N_7770,N_7771,N_7774,N_7775,N_7776,N_7778,N_7781,N_7782,N_7783,N_7784,N_7785,N_7787,N_7788,N_7789,N_7792,N_7794,N_7796,N_7797,N_7799,N_7800,N_7804,N_7805,N_7811,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7820,N_7821,N_7822,N_7823,N_7825,N_7826,N_7828,N_7831,N_7838,N_7839,N_7840,N_7842,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7852,N_7853,N_7857,N_7859,N_7860,N_7862,N_7864,N_7865,N_7867,N_7869,N_7870,N_7871,N_7873,N_7874,N_7875,N_7876,N_7878,N_7880,N_7884,N_7886,N_7887,N_7888,N_7891,N_7894,N_7896,N_7898,N_7900,N_7901,N_7903,N_7905,N_7907,N_7908,N_7909,N_7910,N_7911,N_7913,N_7915,N_7916,N_7918,N_7919,N_7920,N_7921,N_7924,N_7925,N_7926,N_7927,N_7929,N_7931,N_7932,N_7934,N_7935,N_7936,N_7937,N_7940,N_7941,N_7942,N_7943,N_7946,N_7950,N_7951,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7968,N_7969,N_7972,N_7973,N_7975,N_7980,N_7981,N_7982,N_7983,N_7984,N_7986,N_7988,N_7991,N_7992,N_7993,N_7995,N_7999,N_8000,N_8001,N_8002,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8012,N_8014,N_8016,N_8018,N_8019,N_8020,N_8021,N_8025,N_8026,N_8027,N_8029,N_8030,N_8032,N_8035,N_8036,N_8039,N_8041,N_8043,N_8044,N_8045,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8057,N_8060,N_8061,N_8062,N_8063,N_8069,N_8070,N_8071,N_8072,N_8074,N_8076,N_8079,N_8080,N_8081,N_8083,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8092,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8113,N_8114,N_8117,N_8118,N_8119,N_8121,N_8123,N_8125,N_8126,N_8127,N_8129,N_8130,N_8132,N_8133,N_8135,N_8136,N_8138,N_8139,N_8143,N_8144,N_8147,N_8148,N_8149,N_8150,N_8151,N_8159,N_8160,N_8163,N_8167,N_8169,N_8170,N_8174,N_8177,N_8178,N_8180,N_8181,N_8182,N_8183,N_8186,N_8189,N_8191,N_8192,N_8194,N_8196,N_8197,N_8198,N_8206,N_8209,N_8210,N_8211,N_8212,N_8214,N_8215,N_8217,N_8218,N_8219,N_8225,N_8228,N_8230,N_8231,N_8237,N_8239,N_8242,N_8243,N_8244,N_8245,N_8246,N_8251,N_8252,N_8254,N_8257,N_8258,N_8259,N_8260,N_8262,N_8263,N_8264,N_8265,N_8267,N_8269,N_8271,N_8272,N_8273,N_8274,N_8275,N_8278,N_8279,N_8280,N_8281,N_8282,N_8284,N_8288,N_8289,N_8291,N_8293,N_8294,N_8295,N_8298,N_8300,N_8304,N_8306,N_8307,N_8309,N_8311,N_8312,N_8316,N_8318,N_8320,N_8321,N_8323,N_8324,N_8325,N_8329,N_8330,N_8334,N_8335,N_8337,N_8338,N_8339,N_8340,N_8341,N_8345,N_8347,N_8348,N_8351,N_8352,N_8355,N_8356,N_8357,N_8358,N_8359,N_8362,N_8364,N_8365,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8374,N_8375,N_8376,N_8378,N_8379,N_8380,N_8383,N_8384,N_8385,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8400,N_8402,N_8403,N_8405,N_8406,N_8407,N_8408,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8422,N_8423,N_8424,N_8425,N_8426,N_8428,N_8430,N_8432,N_8433,N_8434,N_8438,N_8441,N_8444,N_8445,N_8450,N_8453,N_8455,N_8457,N_8458,N_8459,N_8460,N_8461,N_8463,N_8464,N_8465,N_8466,N_8467,N_8469,N_8470,N_8471,N_8472,N_8473,N_8475,N_8477,N_8478,N_8479,N_8480,N_8483,N_8484,N_8487,N_8488,N_8495,N_8496,N_8497,N_8498,N_8499,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8510,N_8512,N_8513,N_8515,N_8516,N_8517,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8534,N_8535,N_8536,N_8538,N_8542,N_8543,N_8544,N_8548,N_8552,N_8553,N_8554,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8564,N_8566,N_8569,N_8570,N_8571,N_8573,N_8574,N_8576,N_8578,N_8579,N_8580,N_8581,N_8584,N_8585,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8594,N_8595,N_8596,N_8597,N_8601,N_8602,N_8603,N_8604,N_8605,N_8607,N_8609,N_8610,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8619,N_8620,N_8622,N_8624,N_8626,N_8627,N_8628,N_8630,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8640,N_8642,N_8643,N_8645,N_8646,N_8648,N_8649,N_8650,N_8653,N_8658,N_8660,N_8661,N_8662,N_8663,N_8666,N_8667,N_8669,N_8670,N_8673,N_8674,N_8676,N_8678,N_8681,N_8682,N_8684,N_8685,N_8686,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8698,N_8701,N_8702,N_8704,N_8705,N_8706,N_8707,N_8708,N_8710,N_8711,N_8712,N_8713,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8722,N_8727,N_8728,N_8729,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8739,N_8740,N_8742,N_8743,N_8745,N_8748,N_8749,N_8750,N_8752,N_8754,N_8756,N_8758,N_8760,N_8761,N_8762,N_8763,N_8765,N_8767,N_8768,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8785,N_8786,N_8788,N_8791,N_8792,N_8793,N_8794,N_8795,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8816,N_8817,N_8818,N_8820,N_8825,N_8826,N_8827,N_8828,N_8829,N_8831,N_8832,N_8833,N_8836,N_8838,N_8839,N_8843,N_8846,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8857,N_8859,N_8860,N_8861,N_8862,N_8864,N_8865,N_8866,N_8868,N_8869,N_8870,N_8873,N_8875,N_8877,N_8879,N_8880,N_8881,N_8886,N_8892,N_8896,N_8897,N_8898,N_8899,N_8901,N_8902,N_8903,N_8905,N_8906,N_8907,N_8909,N_8910,N_8912,N_8913,N_8915,N_8916,N_8917,N_8918,N_8920,N_8923,N_8925,N_8927,N_8929,N_8931,N_8935,N_8937,N_8939,N_8940,N_8942,N_8944,N_8945,N_8946,N_8950,N_8951,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8965,N_8967,N_8968,N_8971,N_8975,N_8976,N_8977,N_8979,N_8983,N_8984,N_8985,N_8987,N_8988,N_8991,N_8993,N_8994,N_8995,N_8997,N_8998,N_9003,N_9004,N_9005,N_9006,N_9007,N_9009,N_9010,N_9014,N_9015,N_9016,N_9020,N_9021,N_9022,N_9023,N_9024,N_9026,N_9027,N_9030,N_9031,N_9032,N_9035,N_9036,N_9037,N_9040,N_9042,N_9044,N_9047,N_9049,N_9052,N_9053,N_9055,N_9057,N_9058,N_9065,N_9066,N_9067,N_9068,N_9069,N_9073,N_9075,N_9076,N_9077,N_9079,N_9080,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9090,N_9091,N_9092,N_9093,N_9096,N_9097,N_9102,N_9103,N_9105,N_9106,N_9110,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9122,N_9123,N_9124,N_9131,N_9132,N_9133,N_9134,N_9135,N_9137,N_9141,N_9142,N_9144,N_9146,N_9147,N_9149,N_9150,N_9151,N_9152,N_9153,N_9155,N_9156,N_9157,N_9158,N_9162,N_9165,N_9166,N_9167,N_9170,N_9171,N_9173,N_9176,N_9179,N_9181,N_9182,N_9183,N_9184,N_9186,N_9187,N_9190,N_9192,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9206,N_9207,N_9208,N_9210,N_9211,N_9212,N_9214,N_9216,N_9217,N_9219,N_9220,N_9222,N_9223,N_9224,N_9227,N_9228,N_9229,N_9230,N_9232,N_9233,N_9235,N_9236,N_9237,N_9238,N_9240,N_9242,N_9243,N_9244,N_9247,N_9248,N_9249,N_9250,N_9252,N_9254,N_9255,N_9257,N_9260,N_9263,N_9265,N_9268,N_9270,N_9271,N_9274,N_9275,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9293,N_9296,N_9297,N_9298,N_9299,N_9306,N_9307,N_9308,N_9310,N_9311,N_9312,N_9318,N_9319,N_9320,N_9321,N_9322,N_9326,N_9327,N_9329,N_9333,N_9336,N_9337,N_9339,N_9342,N_9343,N_9344,N_9346,N_9349,N_9350,N_9355,N_9357,N_9358,N_9361,N_9362,N_9363,N_9366,N_9367,N_9368,N_9369,N_9370,N_9372,N_9373,N_9375,N_9376,N_9377,N_9379,N_9380,N_9382,N_9384,N_9385,N_9387,N_9389,N_9390,N_9391,N_9392,N_9394,N_9395,N_9396,N_9399,N_9401,N_9402,N_9403,N_9404,N_9406,N_9407,N_9408,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9428,N_9429,N_9431,N_9434,N_9435,N_9439,N_9442,N_9444,N_9447,N_9448,N_9449,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9461,N_9463,N_9464,N_9467,N_9468,N_9470,N_9471,N_9473,N_9477,N_9479,N_9480,N_9484,N_9488,N_9491,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9502,N_9504,N_9505,N_9506,N_9507,N_9510,N_9511,N_9513,N_9514,N_9516,N_9517,N_9520,N_9523,N_9525,N_9526,N_9527,N_9531,N_9534,N_9538,N_9541,N_9543,N_9544,N_9545,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9558,N_9559,N_9565,N_9575,N_9576,N_9577,N_9580,N_9581,N_9582,N_9584,N_9585,N_9586,N_9589,N_9590,N_9593,N_9594,N_9600,N_9601,N_9602,N_9603,N_9604,N_9606,N_9608,N_9610,N_9611,N_9612,N_9614,N_9618,N_9620,N_9623,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9632,N_9633,N_9634,N_9635,N_9639,N_9641,N_9645,N_9646,N_9648,N_9649,N_9650,N_9652,N_9653,N_9654,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9668,N_9669,N_9671,N_9672,N_9674,N_9676,N_9678,N_9681,N_9682,N_9683,N_9686,N_9688,N_9690,N_9691,N_9692,N_9695,N_9699,N_9700,N_9701,N_9703,N_9705,N_9709,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9731,N_9733,N_9734,N_9735,N_9738,N_9739,N_9740,N_9741,N_9742,N_9745,N_9746,N_9747,N_9748,N_9750,N_9752,N_9753,N_9754,N_9756,N_9758,N_9760,N_9761,N_9762,N_9764,N_9765,N_9766,N_9767,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9778,N_9779,N_9781,N_9783,N_9784,N_9786,N_9790,N_9792,N_9793,N_9795,N_9796,N_9797,N_9798,N_9803,N_9804,N_9805,N_9807,N_9809,N_9812,N_9813,N_9817,N_9818,N_9820,N_9825,N_9826,N_9827,N_9828,N_9831,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9847,N_9850,N_9851,N_9852,N_9854,N_9855,N_9858,N_9859,N_9860,N_9861,N_9863,N_9864,N_9866,N_9868,N_9869,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9878,N_9879,N_9880,N_9882,N_9883,N_9884,N_9887,N_9892,N_9894,N_9895,N_9896,N_9897,N_9899,N_9900,N_9901,N_9906,N_9907,N_9910,N_9911,N_9912,N_9913,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9925,N_9927,N_9928,N_9935,N_9939,N_9940,N_9942,N_9946,N_9948,N_9949,N_9951,N_9955,N_9958,N_9960,N_9962,N_9963,N_9968,N_9973,N_9975,N_9976,N_9978,N_9979,N_9980,N_9981,N_9982,N_9986,N_9987,N_9988,N_9990,N_9991,N_9992,N_9993,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_233,In_76);
or U1 (N_1,In_188,In_213);
nand U2 (N_2,In_831,In_821);
and U3 (N_3,In_986,In_429);
nand U4 (N_4,In_192,In_604);
and U5 (N_5,In_5,In_806);
nand U6 (N_6,In_371,In_397);
nor U7 (N_7,In_288,In_648);
nor U8 (N_8,In_770,In_104);
nor U9 (N_9,In_535,In_217);
and U10 (N_10,In_202,In_178);
nor U11 (N_11,In_682,In_787);
xor U12 (N_12,In_426,In_654);
nor U13 (N_13,In_269,In_227);
and U14 (N_14,In_857,In_749);
nand U15 (N_15,In_897,In_574);
nor U16 (N_16,In_475,In_533);
or U17 (N_17,In_113,In_260);
xnor U18 (N_18,In_567,In_35);
nor U19 (N_19,In_268,In_655);
nand U20 (N_20,In_144,In_414);
and U21 (N_21,In_491,In_669);
or U22 (N_22,In_685,In_52);
and U23 (N_23,In_918,In_455);
nand U24 (N_24,In_273,In_605);
or U25 (N_25,In_622,In_582);
nand U26 (N_26,In_809,In_319);
nor U27 (N_27,In_481,In_150);
or U28 (N_28,In_644,In_106);
nand U29 (N_29,In_247,In_982);
and U30 (N_30,In_142,In_374);
nor U31 (N_31,In_692,In_703);
or U32 (N_32,In_314,In_381);
or U33 (N_33,In_662,In_744);
and U34 (N_34,In_148,In_863);
or U35 (N_35,In_927,In_282);
and U36 (N_36,In_651,In_814);
and U37 (N_37,In_23,In_454);
nor U38 (N_38,In_922,In_805);
nor U39 (N_39,In_80,In_796);
or U40 (N_40,In_496,In_509);
nand U41 (N_41,In_418,In_584);
nor U42 (N_42,In_248,In_717);
or U43 (N_43,In_862,In_577);
and U44 (N_44,In_38,In_867);
or U45 (N_45,In_553,In_262);
xor U46 (N_46,In_132,In_846);
nor U47 (N_47,In_930,In_981);
nor U48 (N_48,In_743,In_665);
and U49 (N_49,In_732,In_546);
nor U50 (N_50,In_524,In_684);
nor U51 (N_51,In_904,In_103);
nand U52 (N_52,In_112,In_708);
nor U53 (N_53,In_354,In_837);
and U54 (N_54,In_82,In_847);
xor U55 (N_55,In_102,In_543);
nor U56 (N_56,In_396,In_766);
xor U57 (N_57,In_780,In_72);
and U58 (N_58,In_125,In_841);
and U59 (N_59,In_915,In_842);
nor U60 (N_60,In_91,In_435);
and U61 (N_61,In_287,In_306);
or U62 (N_62,In_932,In_597);
nor U63 (N_63,In_490,In_758);
nand U64 (N_64,In_569,In_187);
xor U65 (N_65,In_962,In_660);
nand U66 (N_66,In_13,In_398);
or U67 (N_67,In_757,In_228);
nand U68 (N_68,In_512,In_377);
nand U69 (N_69,In_70,In_718);
or U70 (N_70,In_32,In_804);
nand U71 (N_71,In_312,In_39);
nor U72 (N_72,In_712,In_589);
xnor U73 (N_73,In_444,In_368);
nor U74 (N_74,In_898,In_781);
or U75 (N_75,In_741,In_204);
or U76 (N_76,In_189,In_297);
nor U77 (N_77,In_385,In_800);
nor U78 (N_78,In_812,In_552);
nand U79 (N_79,In_166,In_351);
or U80 (N_80,In_753,In_608);
nor U81 (N_81,In_532,In_353);
and U82 (N_82,In_77,In_807);
and U83 (N_83,In_497,In_564);
nand U84 (N_84,In_161,In_172);
nor U85 (N_85,In_924,In_340);
nand U86 (N_86,In_44,In_58);
nor U87 (N_87,In_405,In_246);
nor U88 (N_88,In_430,In_350);
nand U89 (N_89,In_295,In_754);
nand U90 (N_90,In_279,In_464);
and U91 (N_91,In_713,In_561);
or U92 (N_92,In_861,In_794);
nand U93 (N_93,In_699,In_487);
nor U94 (N_94,In_680,In_225);
nand U95 (N_95,In_126,In_85);
nand U96 (N_96,In_493,In_56);
or U97 (N_97,In_941,In_899);
nand U98 (N_98,In_120,In_571);
or U99 (N_99,In_737,In_894);
nor U100 (N_100,In_467,In_652);
nor U101 (N_101,In_394,In_49);
or U102 (N_102,In_24,In_290);
or U103 (N_103,In_688,In_357);
nor U104 (N_104,In_68,In_122);
nand U105 (N_105,In_283,In_214);
or U106 (N_106,In_566,In_829);
or U107 (N_107,In_191,In_154);
or U108 (N_108,In_928,In_627);
or U109 (N_109,In_591,In_105);
nor U110 (N_110,In_690,In_175);
or U111 (N_111,In_506,In_501);
nor U112 (N_112,In_598,In_380);
nor U113 (N_113,In_756,In_793);
nand U114 (N_114,In_453,In_10);
or U115 (N_115,In_60,In_366);
xnor U116 (N_116,In_560,In_65);
and U117 (N_117,In_693,In_205);
nand U118 (N_118,In_379,In_639);
or U119 (N_119,In_782,In_201);
and U120 (N_120,In_346,In_859);
or U121 (N_121,In_519,In_315);
and U122 (N_122,In_983,In_503);
nor U123 (N_123,In_722,In_724);
nand U124 (N_124,In_412,In_289);
and U125 (N_125,In_992,In_222);
nor U126 (N_126,In_152,In_539);
or U127 (N_127,In_638,In_551);
nor U128 (N_128,In_446,In_704);
or U129 (N_129,In_558,In_4);
or U130 (N_130,In_22,In_265);
xnor U131 (N_131,In_590,In_659);
xnor U132 (N_132,In_799,In_719);
or U133 (N_133,In_988,In_739);
nand U134 (N_134,In_0,In_107);
nor U135 (N_135,In_738,In_736);
nor U136 (N_136,In_452,In_447);
nor U137 (N_137,In_970,In_98);
and U138 (N_138,In_402,In_230);
or U139 (N_139,In_384,In_995);
nor U140 (N_140,In_925,In_697);
and U141 (N_141,In_840,In_514);
xor U142 (N_142,In_740,In_403);
nor U143 (N_143,In_733,In_136);
nor U144 (N_144,In_254,In_26);
and U145 (N_145,In_751,In_186);
xnor U146 (N_146,In_42,In_167);
nor U147 (N_147,In_518,In_727);
and U148 (N_148,In_957,In_969);
nor U149 (N_149,In_965,In_792);
or U150 (N_150,In_968,In_876);
nor U151 (N_151,In_536,In_668);
and U152 (N_152,In_728,In_183);
and U153 (N_153,In_801,In_6);
and U154 (N_154,In_270,In_275);
nor U155 (N_155,In_284,In_33);
nor U156 (N_156,In_845,In_411);
nand U157 (N_157,In_785,In_401);
xnor U158 (N_158,In_313,In_825);
nand U159 (N_159,In_675,In_303);
xor U160 (N_160,In_208,In_895);
xnor U161 (N_161,In_231,In_267);
and U162 (N_162,In_909,In_579);
nor U163 (N_163,In_523,In_238);
and U164 (N_164,In_600,In_343);
nor U165 (N_165,In_20,In_310);
nor U166 (N_166,In_413,In_917);
xnor U167 (N_167,In_308,In_159);
nor U168 (N_168,In_271,In_66);
or U169 (N_169,In_939,In_291);
and U170 (N_170,In_74,In_530);
or U171 (N_171,In_907,In_856);
xnor U172 (N_172,In_469,In_823);
nor U173 (N_173,In_694,In_153);
nand U174 (N_174,In_702,In_147);
and U175 (N_175,In_151,In_160);
nor U176 (N_176,In_892,In_991);
nor U177 (N_177,In_215,In_838);
xnor U178 (N_178,In_302,In_94);
and U179 (N_179,In_869,In_936);
nor U180 (N_180,In_14,In_257);
or U181 (N_181,In_48,In_145);
nor U182 (N_182,In_721,In_990);
nor U183 (N_183,In_468,In_725);
and U184 (N_184,In_677,In_365);
and U185 (N_185,In_210,In_93);
nor U186 (N_186,In_479,In_933);
xor U187 (N_187,In_250,In_813);
nor U188 (N_188,In_352,In_47);
nor U189 (N_189,In_701,In_667);
and U190 (N_190,In_849,In_855);
nor U191 (N_191,In_223,In_562);
nand U192 (N_192,In_602,In_92);
nor U193 (N_193,In_811,In_864);
nor U194 (N_194,In_948,In_937);
nand U195 (N_195,In_232,In_342);
or U196 (N_196,In_369,In_544);
nand U197 (N_197,In_179,In_383);
or U198 (N_198,In_996,In_321);
nor U199 (N_199,In_913,In_197);
or U200 (N_200,In_83,In_767);
and U201 (N_201,In_653,In_119);
and U202 (N_202,In_760,In_601);
or U203 (N_203,In_580,In_771);
or U204 (N_204,In_963,In_635);
or U205 (N_205,In_956,In_529);
and U206 (N_206,In_575,In_78);
xor U207 (N_207,In_173,In_362);
and U208 (N_208,In_244,In_537);
nor U209 (N_209,In_695,In_670);
xnor U210 (N_210,In_391,In_603);
nor U211 (N_211,In_619,In_410);
or U212 (N_212,In_599,In_972);
and U213 (N_213,In_372,In_860);
and U214 (N_214,In_696,In_243);
or U215 (N_215,In_209,In_124);
nor U216 (N_216,In_832,In_317);
nand U217 (N_217,In_111,In_616);
or U218 (N_218,In_320,In_489);
or U219 (N_219,In_824,In_43);
or U220 (N_220,In_367,In_613);
xnor U221 (N_221,In_185,In_253);
nor U222 (N_222,In_943,In_830);
nor U223 (N_223,In_504,In_871);
and U224 (N_224,In_8,In_775);
nand U225 (N_225,In_436,In_683);
xor U226 (N_226,In_181,In_798);
and U227 (N_227,In_643,In_339);
nor U228 (N_228,In_997,In_1);
nand U229 (N_229,In_822,In_576);
nor U230 (N_230,In_500,In_387);
nand U231 (N_231,In_108,In_517);
and U232 (N_232,In_345,In_581);
nor U233 (N_233,In_671,In_324);
and U234 (N_234,In_11,In_515);
nand U235 (N_235,In_180,In_707);
nand U236 (N_236,In_709,In_255);
nor U237 (N_237,In_890,In_772);
nand U238 (N_238,In_316,In_661);
nor U239 (N_239,In_274,In_51);
nor U240 (N_240,In_538,In_559);
nand U241 (N_241,In_207,In_585);
nand U242 (N_242,In_168,In_563);
or U243 (N_243,In_656,In_929);
nor U244 (N_244,In_934,In_139);
and U245 (N_245,In_820,In_184);
nor U246 (N_246,In_382,In_555);
and U247 (N_247,In_71,In_672);
xor U248 (N_248,In_110,In_466);
nand U249 (N_249,In_908,In_827);
nor U250 (N_250,In_964,In_980);
nor U251 (N_251,In_9,In_637);
nor U252 (N_252,In_606,In_90);
or U253 (N_253,In_818,In_331);
nor U254 (N_254,In_463,In_67);
nand U255 (N_255,In_901,In_762);
nand U256 (N_256,In_657,In_61);
nand U257 (N_257,In_165,In_25);
nand U258 (N_258,In_417,In_525);
and U259 (N_259,In_157,In_878);
or U260 (N_260,In_761,In_994);
or U261 (N_261,In_286,In_245);
and U262 (N_262,In_236,In_285);
nor U263 (N_263,In_221,In_596);
or U264 (N_264,In_587,In_53);
or U265 (N_265,In_905,In_508);
and U266 (N_266,In_307,In_681);
or U267 (N_267,In_141,In_549);
xor U268 (N_268,In_620,In_406);
nand U269 (N_269,In_358,In_868);
nand U270 (N_270,In_114,In_364);
nor U271 (N_271,In_164,In_41);
nor U272 (N_272,In_344,In_220);
and U273 (N_273,In_592,In_12);
or U274 (N_274,In_926,In_54);
nand U275 (N_275,In_768,In_495);
or U276 (N_276,In_121,In_974);
nor U277 (N_277,In_797,In_674);
xnor U278 (N_278,In_158,In_710);
nor U279 (N_279,In_931,In_477);
and U280 (N_280,In_663,In_541);
and U281 (N_281,In_570,In_547);
and U282 (N_282,In_631,In_568);
nand U283 (N_283,In_673,In_200);
xnor U284 (N_284,In_370,In_473);
nand U285 (N_285,In_872,In_773);
or U286 (N_286,In_296,In_935);
xnor U287 (N_287,In_629,In_609);
nand U288 (N_288,In_706,In_258);
nor U289 (N_289,In_949,In_646);
xnor U290 (N_290,In_816,In_920);
nor U291 (N_291,In_534,In_115);
nor U292 (N_292,In_218,In_338);
and U293 (N_293,In_624,In_947);
or U294 (N_294,In_887,In_755);
and U295 (N_295,In_206,In_439);
nand U296 (N_296,In_610,In_526);
or U297 (N_297,In_664,In_689);
xor U298 (N_298,In_86,In_276);
nand U299 (N_299,In_212,In_626);
nor U300 (N_300,In_263,In_131);
nor U301 (N_301,In_516,In_376);
and U302 (N_302,In_779,In_3);
nand U303 (N_303,In_21,In_774);
or U304 (N_304,In_615,In_415);
nor U305 (N_305,In_942,In_765);
nand U306 (N_306,In_910,In_416);
xnor U307 (N_307,In_557,In_19);
and U308 (N_308,In_998,In_99);
xor U309 (N_309,In_789,In_441);
nor U310 (N_310,In_731,In_146);
or U311 (N_311,In_640,In_836);
or U312 (N_312,In_261,In_171);
and U313 (N_313,In_450,In_828);
nor U314 (N_314,In_434,In_443);
or U315 (N_315,In_75,In_176);
nor U316 (N_316,In_726,In_88);
nand U317 (N_317,In_843,In_961);
nor U318 (N_318,In_449,In_323);
nand U319 (N_319,In_819,In_30);
or U320 (N_320,In_483,In_62);
nand U321 (N_321,In_459,In_746);
nor U322 (N_322,In_118,In_999);
or U323 (N_323,In_676,In_955);
nand U324 (N_324,In_240,In_437);
and U325 (N_325,In_833,In_853);
and U326 (N_326,In_747,In_850);
nand U327 (N_327,In_885,In_329);
or U328 (N_328,In_470,In_216);
nand U329 (N_329,In_226,In_916);
nand U330 (N_330,In_356,In_636);
nor U331 (N_331,In_486,In_896);
nand U332 (N_332,In_953,In_542);
nand U333 (N_333,In_304,In_198);
or U334 (N_334,In_633,In_866);
xnor U335 (N_335,In_548,In_137);
nor U336 (N_336,In_425,In_123);
nor U337 (N_337,In_127,In_128);
nand U338 (N_338,In_888,In_133);
and U339 (N_339,In_720,In_891);
nor U340 (N_340,In_595,In_742);
nor U341 (N_341,In_686,In_911);
or U342 (N_342,In_117,In_388);
or U343 (N_343,In_266,In_630);
nor U344 (N_344,In_634,In_752);
and U345 (N_345,In_883,In_759);
and U346 (N_346,In_815,In_978);
and U347 (N_347,In_714,In_618);
nor U348 (N_348,In_400,In_328);
and U349 (N_349,In_389,In_333);
nand U350 (N_350,In_984,In_241);
or U351 (N_351,In_723,In_407);
and U352 (N_352,In_912,In_427);
and U353 (N_353,In_521,In_392);
and U354 (N_354,In_193,In_36);
nor U355 (N_355,In_461,In_698);
xor U356 (N_356,In_420,In_211);
and U357 (N_357,In_881,In_488);
nand U358 (N_358,In_457,In_873);
nor U359 (N_359,In_802,In_31);
and U360 (N_360,In_919,In_527);
or U361 (N_361,In_734,In_393);
xnor U362 (N_362,In_572,In_777);
or U363 (N_363,In_55,In_554);
nor U364 (N_364,In_502,In_29);
nand U365 (N_365,In_390,In_858);
nand U366 (N_366,In_510,In_817);
xor U367 (N_367,In_373,In_237);
nand U368 (N_368,In_174,In_973);
or U369 (N_369,In_666,In_318);
or U370 (N_370,In_482,In_960);
nand U371 (N_371,In_348,In_292);
or U372 (N_372,In_795,In_810);
nor U373 (N_373,In_776,In_784);
nand U374 (N_374,In_79,In_195);
nor U375 (N_375,In_507,In_903);
nor U376 (N_376,In_251,In_623);
or U377 (N_377,In_900,In_874);
and U378 (N_378,In_880,In_945);
nor U379 (N_379,In_484,In_422);
nor U380 (N_380,In_182,In_641);
nand U381 (N_381,In_89,In_64);
xnor U382 (N_382,In_143,In_341);
xor U383 (N_383,In_647,In_149);
xnor U384 (N_384,In_378,In_330);
nor U385 (N_385,In_69,In_505);
and U386 (N_386,In_687,In_556);
xnor U387 (N_387,In_950,In_940);
and U388 (N_388,In_298,In_498);
or U389 (N_389,In_617,In_778);
nand U390 (N_390,In_478,In_471);
nand U391 (N_391,In_421,In_305);
nand U392 (N_392,In_229,In_395);
or U393 (N_393,In_852,In_844);
nor U394 (N_394,In_879,In_573);
and U395 (N_395,In_854,In_140);
nor U396 (N_396,In_419,In_848);
xnor U397 (N_397,In_116,In_224);
nand U398 (N_398,In_545,In_884);
and U399 (N_399,In_993,In_642);
nor U400 (N_400,In_632,In_336);
nand U401 (N_401,In_985,In_386);
nand U402 (N_402,In_650,In_451);
and U403 (N_403,In_95,In_327);
xnor U404 (N_404,In_485,In_97);
or U405 (N_405,In_729,In_163);
and U406 (N_406,In_989,In_399);
nor U407 (N_407,In_938,In_259);
nor U408 (N_408,In_281,In_235);
and U409 (N_409,In_870,In_875);
or U410 (N_410,In_790,In_886);
or U411 (N_411,In_611,In_404);
nand U412 (N_412,In_588,In_788);
xor U413 (N_413,In_256,In_700);
or U414 (N_414,In_480,In_906);
nand U415 (N_415,In_332,In_134);
xnor U416 (N_416,In_474,In_347);
and U417 (N_417,In_252,In_162);
nor U418 (N_418,In_431,In_277);
nand U419 (N_419,In_349,In_967);
and U420 (N_420,In_309,In_882);
or U421 (N_421,In_46,In_300);
and U422 (N_422,In_958,In_976);
nand U423 (N_423,In_944,In_522);
nor U424 (N_424,In_803,In_607);
or U425 (N_425,In_101,In_326);
or U426 (N_426,In_40,In_448);
and U427 (N_427,In_155,In_360);
or U428 (N_428,In_130,In_199);
nor U429 (N_429,In_791,In_966);
and U430 (N_430,In_359,In_835);
nand U431 (N_431,In_409,In_839);
xnor U432 (N_432,In_977,In_96);
nand U433 (N_433,In_15,In_280);
nand U434 (N_434,In_594,In_625);
or U435 (N_435,In_239,In_363);
or U436 (N_436,In_540,In_34);
nor U437 (N_437,In_196,In_921);
and U438 (N_438,In_954,In_764);
nand U439 (N_439,In_177,In_63);
nand U440 (N_440,In_783,In_628);
or U441 (N_441,In_135,In_442);
or U442 (N_442,In_494,In_293);
or U443 (N_443,In_2,In_614);
and U444 (N_444,In_649,In_465);
nand U445 (N_445,In_492,In_987);
nor U446 (N_446,In_902,In_45);
and U447 (N_447,In_129,In_299);
and U448 (N_448,In_971,In_445);
nand U449 (N_449,In_834,In_301);
nor U450 (N_450,In_578,In_550);
nor U451 (N_451,In_337,In_889);
nand U452 (N_452,In_264,In_57);
and U453 (N_453,In_786,In_423);
and U454 (N_454,In_375,In_745);
or U455 (N_455,In_511,In_750);
xnor U456 (N_456,In_335,In_460);
and U457 (N_457,In_769,In_826);
or U458 (N_458,In_433,In_658);
or U459 (N_459,In_249,In_715);
nor U460 (N_460,In_865,In_408);
or U461 (N_461,In_194,In_18);
and U462 (N_462,In_27,In_278);
and U463 (N_463,In_59,In_735);
and U464 (N_464,In_311,In_877);
xnor U465 (N_465,In_87,In_893);
or U466 (N_466,In_520,In_705);
and U467 (N_467,In_294,In_322);
or U468 (N_468,In_458,In_219);
nor U469 (N_469,In_432,In_361);
or U470 (N_470,In_959,In_583);
nand U471 (N_471,In_428,In_438);
nor U472 (N_472,In_170,In_424);
and U473 (N_473,In_951,In_472);
or U474 (N_474,In_190,In_81);
xnor U475 (N_475,In_28,In_242);
nor U476 (N_476,In_156,In_716);
nor U477 (N_477,In_440,In_16);
nand U478 (N_478,In_678,In_612);
and U479 (N_479,In_203,In_946);
nor U480 (N_480,In_586,In_763);
and U481 (N_481,In_17,In_851);
xnor U482 (N_482,In_528,In_979);
and U483 (N_483,In_914,In_691);
and U484 (N_484,In_234,In_808);
xnor U485 (N_485,In_499,In_565);
nand U486 (N_486,In_952,In_37);
nand U487 (N_487,In_531,In_100);
nand U488 (N_488,In_50,In_456);
or U489 (N_489,In_7,In_462);
and U490 (N_490,In_975,In_645);
nand U491 (N_491,In_476,In_334);
nor U492 (N_492,In_621,In_513);
nor U493 (N_493,In_355,In_84);
nand U494 (N_494,In_169,In_325);
and U495 (N_495,In_272,In_593);
nor U496 (N_496,In_73,In_923);
nand U497 (N_497,In_730,In_138);
nand U498 (N_498,In_711,In_748);
nand U499 (N_499,In_109,In_679);
or U500 (N_500,In_283,In_827);
nor U501 (N_501,In_184,In_619);
or U502 (N_502,In_206,In_108);
and U503 (N_503,In_596,In_462);
xnor U504 (N_504,In_183,In_409);
and U505 (N_505,In_302,In_590);
nand U506 (N_506,In_314,In_361);
xor U507 (N_507,In_919,In_360);
nor U508 (N_508,In_939,In_549);
nand U509 (N_509,In_847,In_200);
and U510 (N_510,In_961,In_940);
nand U511 (N_511,In_822,In_450);
or U512 (N_512,In_82,In_950);
xnor U513 (N_513,In_113,In_941);
and U514 (N_514,In_983,In_44);
nor U515 (N_515,In_320,In_917);
nor U516 (N_516,In_491,In_554);
or U517 (N_517,In_640,In_797);
xor U518 (N_518,In_354,In_5);
and U519 (N_519,In_976,In_914);
and U520 (N_520,In_647,In_69);
and U521 (N_521,In_769,In_922);
or U522 (N_522,In_872,In_125);
nor U523 (N_523,In_456,In_658);
nand U524 (N_524,In_400,In_851);
nor U525 (N_525,In_529,In_382);
nor U526 (N_526,In_864,In_594);
nor U527 (N_527,In_735,In_432);
or U528 (N_528,In_478,In_274);
nand U529 (N_529,In_561,In_555);
nand U530 (N_530,In_305,In_489);
nand U531 (N_531,In_762,In_658);
and U532 (N_532,In_390,In_535);
and U533 (N_533,In_398,In_480);
and U534 (N_534,In_435,In_331);
nand U535 (N_535,In_167,In_892);
and U536 (N_536,In_645,In_343);
and U537 (N_537,In_783,In_873);
xnor U538 (N_538,In_234,In_231);
or U539 (N_539,In_612,In_421);
nor U540 (N_540,In_48,In_890);
nand U541 (N_541,In_618,In_703);
or U542 (N_542,In_793,In_264);
nor U543 (N_543,In_297,In_813);
or U544 (N_544,In_881,In_857);
and U545 (N_545,In_647,In_158);
or U546 (N_546,In_873,In_14);
nor U547 (N_547,In_640,In_815);
and U548 (N_548,In_888,In_355);
xnor U549 (N_549,In_165,In_773);
and U550 (N_550,In_139,In_433);
or U551 (N_551,In_37,In_593);
or U552 (N_552,In_349,In_411);
or U553 (N_553,In_881,In_461);
and U554 (N_554,In_23,In_604);
nand U555 (N_555,In_413,In_964);
nor U556 (N_556,In_252,In_862);
nand U557 (N_557,In_282,In_416);
or U558 (N_558,In_341,In_967);
nand U559 (N_559,In_415,In_676);
nand U560 (N_560,In_299,In_420);
and U561 (N_561,In_364,In_122);
or U562 (N_562,In_943,In_743);
nand U563 (N_563,In_27,In_506);
nor U564 (N_564,In_845,In_151);
or U565 (N_565,In_369,In_316);
and U566 (N_566,In_626,In_862);
nor U567 (N_567,In_213,In_606);
and U568 (N_568,In_611,In_291);
xnor U569 (N_569,In_604,In_978);
or U570 (N_570,In_553,In_393);
nand U571 (N_571,In_452,In_704);
or U572 (N_572,In_124,In_154);
or U573 (N_573,In_810,In_127);
nand U574 (N_574,In_695,In_479);
or U575 (N_575,In_697,In_86);
or U576 (N_576,In_38,In_277);
nor U577 (N_577,In_256,In_747);
nand U578 (N_578,In_383,In_774);
nand U579 (N_579,In_837,In_69);
xor U580 (N_580,In_439,In_781);
or U581 (N_581,In_748,In_814);
or U582 (N_582,In_767,In_69);
and U583 (N_583,In_538,In_102);
or U584 (N_584,In_100,In_743);
or U585 (N_585,In_873,In_106);
nand U586 (N_586,In_613,In_433);
nand U587 (N_587,In_741,In_878);
and U588 (N_588,In_525,In_155);
xor U589 (N_589,In_532,In_813);
and U590 (N_590,In_961,In_239);
xnor U591 (N_591,In_279,In_759);
nor U592 (N_592,In_749,In_605);
nand U593 (N_593,In_466,In_478);
or U594 (N_594,In_88,In_486);
or U595 (N_595,In_690,In_44);
xnor U596 (N_596,In_195,In_924);
nand U597 (N_597,In_30,In_789);
or U598 (N_598,In_778,In_141);
nand U599 (N_599,In_630,In_15);
and U600 (N_600,In_396,In_638);
nor U601 (N_601,In_671,In_510);
or U602 (N_602,In_796,In_872);
xor U603 (N_603,In_925,In_394);
or U604 (N_604,In_656,In_948);
xor U605 (N_605,In_277,In_244);
nand U606 (N_606,In_381,In_857);
and U607 (N_607,In_912,In_749);
or U608 (N_608,In_944,In_292);
nor U609 (N_609,In_903,In_220);
xor U610 (N_610,In_678,In_600);
and U611 (N_611,In_990,In_261);
nor U612 (N_612,In_357,In_422);
and U613 (N_613,In_455,In_738);
xor U614 (N_614,In_899,In_812);
and U615 (N_615,In_531,In_261);
nor U616 (N_616,In_363,In_736);
or U617 (N_617,In_213,In_534);
or U618 (N_618,In_877,In_191);
and U619 (N_619,In_846,In_948);
nor U620 (N_620,In_107,In_945);
or U621 (N_621,In_621,In_882);
and U622 (N_622,In_516,In_540);
and U623 (N_623,In_443,In_150);
nand U624 (N_624,In_492,In_174);
and U625 (N_625,In_964,In_525);
nor U626 (N_626,In_943,In_915);
and U627 (N_627,In_565,In_827);
nor U628 (N_628,In_571,In_240);
or U629 (N_629,In_697,In_673);
and U630 (N_630,In_229,In_976);
and U631 (N_631,In_264,In_671);
and U632 (N_632,In_262,In_77);
nor U633 (N_633,In_738,In_908);
nor U634 (N_634,In_975,In_419);
nand U635 (N_635,In_165,In_180);
or U636 (N_636,In_496,In_350);
and U637 (N_637,In_580,In_406);
or U638 (N_638,In_75,In_872);
nand U639 (N_639,In_842,In_757);
and U640 (N_640,In_826,In_662);
nor U641 (N_641,In_414,In_353);
or U642 (N_642,In_449,In_93);
nor U643 (N_643,In_680,In_317);
and U644 (N_644,In_26,In_394);
or U645 (N_645,In_444,In_592);
nand U646 (N_646,In_510,In_14);
nor U647 (N_647,In_470,In_336);
xnor U648 (N_648,In_734,In_170);
nor U649 (N_649,In_450,In_419);
nor U650 (N_650,In_672,In_660);
or U651 (N_651,In_116,In_327);
and U652 (N_652,In_726,In_826);
nand U653 (N_653,In_89,In_699);
or U654 (N_654,In_703,In_349);
or U655 (N_655,In_80,In_748);
nand U656 (N_656,In_836,In_20);
xnor U657 (N_657,In_644,In_946);
and U658 (N_658,In_225,In_557);
nor U659 (N_659,In_685,In_63);
nor U660 (N_660,In_28,In_183);
nor U661 (N_661,In_664,In_753);
nor U662 (N_662,In_121,In_797);
xor U663 (N_663,In_215,In_426);
nor U664 (N_664,In_863,In_793);
nor U665 (N_665,In_598,In_808);
and U666 (N_666,In_194,In_419);
nand U667 (N_667,In_464,In_789);
nor U668 (N_668,In_488,In_614);
nor U669 (N_669,In_828,In_843);
and U670 (N_670,In_622,In_870);
xnor U671 (N_671,In_983,In_769);
xnor U672 (N_672,In_238,In_839);
and U673 (N_673,In_980,In_622);
and U674 (N_674,In_488,In_463);
xor U675 (N_675,In_820,In_498);
nand U676 (N_676,In_511,In_82);
or U677 (N_677,In_964,In_372);
nor U678 (N_678,In_345,In_998);
nand U679 (N_679,In_502,In_31);
and U680 (N_680,In_367,In_658);
nand U681 (N_681,In_973,In_840);
nor U682 (N_682,In_229,In_323);
or U683 (N_683,In_722,In_702);
nor U684 (N_684,In_304,In_176);
or U685 (N_685,In_327,In_100);
nand U686 (N_686,In_544,In_677);
and U687 (N_687,In_237,In_986);
nor U688 (N_688,In_789,In_921);
or U689 (N_689,In_140,In_722);
and U690 (N_690,In_766,In_869);
nor U691 (N_691,In_794,In_179);
nand U692 (N_692,In_719,In_801);
xor U693 (N_693,In_289,In_490);
or U694 (N_694,In_187,In_965);
xor U695 (N_695,In_158,In_670);
or U696 (N_696,In_876,In_795);
nand U697 (N_697,In_633,In_470);
xnor U698 (N_698,In_445,In_159);
xnor U699 (N_699,In_99,In_829);
and U700 (N_700,In_70,In_966);
or U701 (N_701,In_331,In_858);
nand U702 (N_702,In_695,In_774);
nor U703 (N_703,In_603,In_411);
or U704 (N_704,In_439,In_356);
nand U705 (N_705,In_71,In_866);
and U706 (N_706,In_613,In_936);
nand U707 (N_707,In_562,In_134);
nor U708 (N_708,In_380,In_843);
or U709 (N_709,In_1,In_305);
and U710 (N_710,In_968,In_723);
or U711 (N_711,In_199,In_359);
or U712 (N_712,In_569,In_145);
xnor U713 (N_713,In_329,In_956);
nand U714 (N_714,In_852,In_574);
xnor U715 (N_715,In_89,In_531);
xnor U716 (N_716,In_37,In_996);
or U717 (N_717,In_810,In_617);
or U718 (N_718,In_341,In_89);
and U719 (N_719,In_850,In_322);
nand U720 (N_720,In_353,In_300);
or U721 (N_721,In_215,In_815);
and U722 (N_722,In_721,In_629);
and U723 (N_723,In_801,In_466);
or U724 (N_724,In_304,In_993);
or U725 (N_725,In_696,In_419);
nand U726 (N_726,In_756,In_61);
nand U727 (N_727,In_146,In_678);
nor U728 (N_728,In_603,In_115);
nor U729 (N_729,In_567,In_706);
or U730 (N_730,In_157,In_550);
nor U731 (N_731,In_644,In_270);
nor U732 (N_732,In_987,In_118);
nand U733 (N_733,In_585,In_236);
nand U734 (N_734,In_204,In_370);
or U735 (N_735,In_818,In_324);
or U736 (N_736,In_546,In_996);
nand U737 (N_737,In_369,In_425);
or U738 (N_738,In_756,In_841);
or U739 (N_739,In_303,In_714);
or U740 (N_740,In_772,In_593);
xor U741 (N_741,In_686,In_126);
and U742 (N_742,In_218,In_18);
or U743 (N_743,In_582,In_437);
nand U744 (N_744,In_329,In_755);
nor U745 (N_745,In_231,In_472);
and U746 (N_746,In_717,In_183);
nand U747 (N_747,In_698,In_387);
or U748 (N_748,In_42,In_667);
or U749 (N_749,In_850,In_215);
or U750 (N_750,In_691,In_916);
or U751 (N_751,In_688,In_530);
xnor U752 (N_752,In_140,In_331);
nor U753 (N_753,In_791,In_355);
xor U754 (N_754,In_34,In_670);
nor U755 (N_755,In_480,In_209);
nor U756 (N_756,In_344,In_378);
nand U757 (N_757,In_673,In_742);
xor U758 (N_758,In_287,In_936);
xnor U759 (N_759,In_142,In_852);
or U760 (N_760,In_566,In_208);
and U761 (N_761,In_533,In_864);
or U762 (N_762,In_420,In_327);
or U763 (N_763,In_632,In_658);
nand U764 (N_764,In_944,In_772);
nand U765 (N_765,In_276,In_875);
or U766 (N_766,In_934,In_978);
nor U767 (N_767,In_402,In_823);
or U768 (N_768,In_39,In_980);
nand U769 (N_769,In_771,In_357);
or U770 (N_770,In_803,In_596);
or U771 (N_771,In_809,In_428);
xor U772 (N_772,In_428,In_27);
nand U773 (N_773,In_839,In_829);
xor U774 (N_774,In_706,In_373);
and U775 (N_775,In_955,In_283);
and U776 (N_776,In_859,In_297);
or U777 (N_777,In_472,In_794);
and U778 (N_778,In_132,In_58);
nor U779 (N_779,In_874,In_234);
or U780 (N_780,In_770,In_645);
and U781 (N_781,In_142,In_60);
and U782 (N_782,In_953,In_183);
and U783 (N_783,In_722,In_223);
and U784 (N_784,In_480,In_331);
nand U785 (N_785,In_565,In_640);
nand U786 (N_786,In_539,In_822);
or U787 (N_787,In_790,In_812);
nand U788 (N_788,In_298,In_16);
or U789 (N_789,In_57,In_72);
or U790 (N_790,In_653,In_935);
nor U791 (N_791,In_673,In_494);
or U792 (N_792,In_432,In_172);
nand U793 (N_793,In_97,In_382);
nand U794 (N_794,In_986,In_971);
nor U795 (N_795,In_609,In_269);
and U796 (N_796,In_850,In_736);
and U797 (N_797,In_22,In_667);
nor U798 (N_798,In_899,In_918);
nor U799 (N_799,In_531,In_623);
nand U800 (N_800,In_661,In_942);
nand U801 (N_801,In_836,In_241);
and U802 (N_802,In_308,In_641);
nor U803 (N_803,In_192,In_897);
or U804 (N_804,In_42,In_353);
and U805 (N_805,In_822,In_365);
and U806 (N_806,In_201,In_170);
xnor U807 (N_807,In_488,In_967);
nand U808 (N_808,In_917,In_957);
or U809 (N_809,In_139,In_307);
nand U810 (N_810,In_959,In_744);
nor U811 (N_811,In_30,In_417);
nor U812 (N_812,In_652,In_401);
or U813 (N_813,In_103,In_694);
nor U814 (N_814,In_608,In_406);
or U815 (N_815,In_99,In_384);
xor U816 (N_816,In_872,In_30);
or U817 (N_817,In_616,In_409);
and U818 (N_818,In_295,In_216);
or U819 (N_819,In_190,In_828);
nand U820 (N_820,In_302,In_603);
nand U821 (N_821,In_984,In_86);
nand U822 (N_822,In_17,In_800);
or U823 (N_823,In_337,In_643);
xnor U824 (N_824,In_266,In_726);
nor U825 (N_825,In_713,In_377);
nand U826 (N_826,In_853,In_322);
and U827 (N_827,In_209,In_310);
nand U828 (N_828,In_19,In_477);
or U829 (N_829,In_402,In_431);
nand U830 (N_830,In_154,In_725);
and U831 (N_831,In_504,In_179);
and U832 (N_832,In_772,In_472);
or U833 (N_833,In_154,In_519);
nor U834 (N_834,In_346,In_72);
nand U835 (N_835,In_712,In_802);
nand U836 (N_836,In_784,In_144);
xor U837 (N_837,In_775,In_737);
nand U838 (N_838,In_52,In_335);
nor U839 (N_839,In_812,In_196);
and U840 (N_840,In_890,In_27);
or U841 (N_841,In_223,In_414);
xnor U842 (N_842,In_120,In_268);
nor U843 (N_843,In_485,In_326);
nand U844 (N_844,In_528,In_827);
nor U845 (N_845,In_306,In_652);
xnor U846 (N_846,In_183,In_392);
xor U847 (N_847,In_25,In_944);
or U848 (N_848,In_204,In_342);
or U849 (N_849,In_503,In_368);
or U850 (N_850,In_485,In_199);
nor U851 (N_851,In_523,In_741);
nand U852 (N_852,In_190,In_398);
and U853 (N_853,In_508,In_531);
xor U854 (N_854,In_619,In_727);
and U855 (N_855,In_386,In_534);
nand U856 (N_856,In_601,In_279);
nand U857 (N_857,In_871,In_824);
and U858 (N_858,In_838,In_941);
nor U859 (N_859,In_477,In_454);
nor U860 (N_860,In_305,In_323);
and U861 (N_861,In_529,In_838);
and U862 (N_862,In_276,In_212);
nand U863 (N_863,In_735,In_698);
nor U864 (N_864,In_894,In_714);
nor U865 (N_865,In_517,In_105);
or U866 (N_866,In_869,In_944);
nor U867 (N_867,In_962,In_223);
and U868 (N_868,In_903,In_651);
nand U869 (N_869,In_42,In_805);
nand U870 (N_870,In_92,In_252);
nor U871 (N_871,In_87,In_237);
and U872 (N_872,In_24,In_700);
nor U873 (N_873,In_664,In_862);
xnor U874 (N_874,In_865,In_750);
nor U875 (N_875,In_821,In_407);
or U876 (N_876,In_143,In_253);
or U877 (N_877,In_285,In_168);
xnor U878 (N_878,In_878,In_271);
and U879 (N_879,In_555,In_421);
xor U880 (N_880,In_602,In_283);
or U881 (N_881,In_58,In_233);
or U882 (N_882,In_188,In_441);
nor U883 (N_883,In_446,In_821);
nand U884 (N_884,In_334,In_556);
xor U885 (N_885,In_819,In_799);
and U886 (N_886,In_285,In_485);
nor U887 (N_887,In_897,In_857);
or U888 (N_888,In_49,In_835);
nand U889 (N_889,In_60,In_521);
or U890 (N_890,In_920,In_180);
nand U891 (N_891,In_201,In_887);
and U892 (N_892,In_22,In_68);
and U893 (N_893,In_850,In_717);
nand U894 (N_894,In_585,In_848);
nor U895 (N_895,In_566,In_139);
nand U896 (N_896,In_762,In_592);
or U897 (N_897,In_43,In_241);
or U898 (N_898,In_4,In_391);
and U899 (N_899,In_191,In_376);
xor U900 (N_900,In_509,In_157);
nor U901 (N_901,In_236,In_827);
nor U902 (N_902,In_93,In_381);
nor U903 (N_903,In_73,In_99);
nor U904 (N_904,In_111,In_444);
nor U905 (N_905,In_417,In_62);
or U906 (N_906,In_773,In_893);
and U907 (N_907,In_91,In_353);
or U908 (N_908,In_239,In_774);
or U909 (N_909,In_895,In_957);
or U910 (N_910,In_397,In_34);
xor U911 (N_911,In_816,In_860);
and U912 (N_912,In_588,In_746);
nor U913 (N_913,In_544,In_271);
nor U914 (N_914,In_727,In_21);
nand U915 (N_915,In_178,In_270);
nand U916 (N_916,In_300,In_621);
nand U917 (N_917,In_771,In_70);
xnor U918 (N_918,In_155,In_255);
xnor U919 (N_919,In_175,In_880);
nand U920 (N_920,In_825,In_873);
or U921 (N_921,In_125,In_431);
or U922 (N_922,In_658,In_529);
xor U923 (N_923,In_203,In_348);
xnor U924 (N_924,In_972,In_533);
nand U925 (N_925,In_76,In_188);
nand U926 (N_926,In_491,In_455);
xnor U927 (N_927,In_472,In_375);
nand U928 (N_928,In_747,In_83);
nand U929 (N_929,In_592,In_250);
and U930 (N_930,In_531,In_319);
nand U931 (N_931,In_910,In_206);
and U932 (N_932,In_728,In_351);
and U933 (N_933,In_720,In_93);
or U934 (N_934,In_485,In_279);
nand U935 (N_935,In_755,In_312);
or U936 (N_936,In_827,In_521);
or U937 (N_937,In_143,In_205);
nand U938 (N_938,In_768,In_489);
nor U939 (N_939,In_8,In_786);
xor U940 (N_940,In_429,In_287);
and U941 (N_941,In_198,In_632);
or U942 (N_942,In_186,In_39);
xor U943 (N_943,In_242,In_15);
xnor U944 (N_944,In_49,In_357);
nor U945 (N_945,In_192,In_471);
and U946 (N_946,In_601,In_786);
or U947 (N_947,In_650,In_504);
or U948 (N_948,In_369,In_486);
nor U949 (N_949,In_668,In_110);
and U950 (N_950,In_83,In_177);
or U951 (N_951,In_188,In_845);
or U952 (N_952,In_985,In_954);
xor U953 (N_953,In_610,In_558);
or U954 (N_954,In_811,In_538);
nand U955 (N_955,In_101,In_904);
nand U956 (N_956,In_913,In_988);
and U957 (N_957,In_857,In_971);
nor U958 (N_958,In_28,In_535);
or U959 (N_959,In_691,In_230);
nand U960 (N_960,In_743,In_711);
nor U961 (N_961,In_37,In_158);
nand U962 (N_962,In_253,In_148);
nand U963 (N_963,In_969,In_794);
and U964 (N_964,In_293,In_801);
or U965 (N_965,In_285,In_892);
nor U966 (N_966,In_655,In_803);
and U967 (N_967,In_704,In_823);
nand U968 (N_968,In_6,In_475);
and U969 (N_969,In_530,In_907);
xnor U970 (N_970,In_232,In_959);
nand U971 (N_971,In_258,In_44);
xnor U972 (N_972,In_850,In_942);
and U973 (N_973,In_126,In_73);
or U974 (N_974,In_140,In_337);
nand U975 (N_975,In_475,In_416);
nor U976 (N_976,In_244,In_269);
nand U977 (N_977,In_927,In_591);
or U978 (N_978,In_222,In_931);
and U979 (N_979,In_878,In_675);
nor U980 (N_980,In_265,In_741);
or U981 (N_981,In_525,In_5);
and U982 (N_982,In_200,In_717);
and U983 (N_983,In_636,In_508);
nor U984 (N_984,In_161,In_396);
or U985 (N_985,In_980,In_495);
nor U986 (N_986,In_604,In_878);
or U987 (N_987,In_310,In_898);
or U988 (N_988,In_609,In_578);
nor U989 (N_989,In_53,In_392);
and U990 (N_990,In_133,In_549);
and U991 (N_991,In_664,In_268);
nand U992 (N_992,In_108,In_219);
xnor U993 (N_993,In_430,In_60);
or U994 (N_994,In_772,In_959);
or U995 (N_995,In_673,In_215);
nand U996 (N_996,In_292,In_221);
xor U997 (N_997,In_310,In_109);
xnor U998 (N_998,In_558,In_704);
nand U999 (N_999,In_726,In_99);
or U1000 (N_1000,In_163,In_164);
and U1001 (N_1001,In_630,In_487);
or U1002 (N_1002,In_1,In_343);
and U1003 (N_1003,In_719,In_449);
and U1004 (N_1004,In_169,In_723);
or U1005 (N_1005,In_5,In_162);
nand U1006 (N_1006,In_800,In_802);
nor U1007 (N_1007,In_879,In_576);
and U1008 (N_1008,In_733,In_171);
and U1009 (N_1009,In_224,In_148);
or U1010 (N_1010,In_534,In_347);
and U1011 (N_1011,In_825,In_239);
nor U1012 (N_1012,In_450,In_636);
nand U1013 (N_1013,In_60,In_328);
and U1014 (N_1014,In_520,In_386);
and U1015 (N_1015,In_796,In_3);
or U1016 (N_1016,In_636,In_506);
nand U1017 (N_1017,In_278,In_733);
or U1018 (N_1018,In_112,In_375);
or U1019 (N_1019,In_838,In_516);
nand U1020 (N_1020,In_79,In_881);
nand U1021 (N_1021,In_558,In_891);
nor U1022 (N_1022,In_955,In_222);
nand U1023 (N_1023,In_328,In_808);
nor U1024 (N_1024,In_551,In_765);
nor U1025 (N_1025,In_908,In_533);
nand U1026 (N_1026,In_372,In_226);
and U1027 (N_1027,In_299,In_676);
nand U1028 (N_1028,In_384,In_146);
nand U1029 (N_1029,In_255,In_504);
and U1030 (N_1030,In_377,In_712);
and U1031 (N_1031,In_523,In_379);
nor U1032 (N_1032,In_10,In_744);
and U1033 (N_1033,In_369,In_705);
nand U1034 (N_1034,In_189,In_686);
nor U1035 (N_1035,In_426,In_91);
and U1036 (N_1036,In_51,In_810);
or U1037 (N_1037,In_778,In_429);
nand U1038 (N_1038,In_277,In_453);
and U1039 (N_1039,In_630,In_666);
and U1040 (N_1040,In_290,In_837);
and U1041 (N_1041,In_815,In_914);
nor U1042 (N_1042,In_973,In_369);
nand U1043 (N_1043,In_223,In_371);
or U1044 (N_1044,In_153,In_401);
nor U1045 (N_1045,In_910,In_438);
and U1046 (N_1046,In_678,In_41);
or U1047 (N_1047,In_155,In_712);
or U1048 (N_1048,In_881,In_98);
and U1049 (N_1049,In_1,In_759);
or U1050 (N_1050,In_713,In_535);
or U1051 (N_1051,In_769,In_847);
or U1052 (N_1052,In_155,In_425);
xor U1053 (N_1053,In_395,In_696);
nand U1054 (N_1054,In_36,In_12);
nand U1055 (N_1055,In_499,In_978);
nand U1056 (N_1056,In_823,In_343);
xor U1057 (N_1057,In_295,In_662);
nand U1058 (N_1058,In_125,In_882);
and U1059 (N_1059,In_287,In_78);
nor U1060 (N_1060,In_514,In_538);
and U1061 (N_1061,In_983,In_684);
or U1062 (N_1062,In_606,In_517);
xnor U1063 (N_1063,In_7,In_891);
nand U1064 (N_1064,In_543,In_796);
nand U1065 (N_1065,In_31,In_800);
and U1066 (N_1066,In_760,In_463);
nand U1067 (N_1067,In_629,In_383);
xnor U1068 (N_1068,In_969,In_956);
and U1069 (N_1069,In_204,In_184);
or U1070 (N_1070,In_366,In_373);
nand U1071 (N_1071,In_533,In_861);
or U1072 (N_1072,In_587,In_783);
or U1073 (N_1073,In_51,In_111);
and U1074 (N_1074,In_757,In_347);
and U1075 (N_1075,In_939,In_25);
nand U1076 (N_1076,In_920,In_251);
or U1077 (N_1077,In_854,In_381);
and U1078 (N_1078,In_626,In_378);
and U1079 (N_1079,In_168,In_450);
nand U1080 (N_1080,In_174,In_794);
nor U1081 (N_1081,In_650,In_990);
and U1082 (N_1082,In_695,In_289);
nor U1083 (N_1083,In_149,In_707);
nor U1084 (N_1084,In_408,In_273);
and U1085 (N_1085,In_838,In_118);
nor U1086 (N_1086,In_413,In_921);
xnor U1087 (N_1087,In_748,In_931);
or U1088 (N_1088,In_910,In_909);
nor U1089 (N_1089,In_280,In_635);
and U1090 (N_1090,In_183,In_859);
nor U1091 (N_1091,In_747,In_487);
or U1092 (N_1092,In_133,In_391);
nand U1093 (N_1093,In_413,In_711);
nor U1094 (N_1094,In_283,In_806);
nor U1095 (N_1095,In_399,In_998);
nor U1096 (N_1096,In_26,In_601);
nor U1097 (N_1097,In_176,In_989);
nor U1098 (N_1098,In_779,In_85);
nand U1099 (N_1099,In_852,In_676);
nand U1100 (N_1100,In_190,In_128);
and U1101 (N_1101,In_932,In_972);
and U1102 (N_1102,In_469,In_92);
nand U1103 (N_1103,In_423,In_342);
and U1104 (N_1104,In_930,In_106);
or U1105 (N_1105,In_792,In_108);
nand U1106 (N_1106,In_225,In_521);
nand U1107 (N_1107,In_736,In_330);
and U1108 (N_1108,In_214,In_465);
nor U1109 (N_1109,In_214,In_419);
and U1110 (N_1110,In_222,In_83);
nand U1111 (N_1111,In_190,In_852);
nor U1112 (N_1112,In_536,In_549);
or U1113 (N_1113,In_124,In_489);
nor U1114 (N_1114,In_296,In_906);
or U1115 (N_1115,In_130,In_738);
nor U1116 (N_1116,In_368,In_238);
and U1117 (N_1117,In_141,In_943);
nand U1118 (N_1118,In_616,In_767);
xnor U1119 (N_1119,In_16,In_545);
and U1120 (N_1120,In_286,In_353);
and U1121 (N_1121,In_483,In_702);
nand U1122 (N_1122,In_554,In_444);
and U1123 (N_1123,In_859,In_379);
or U1124 (N_1124,In_661,In_330);
nor U1125 (N_1125,In_949,In_204);
or U1126 (N_1126,In_448,In_126);
xnor U1127 (N_1127,In_559,In_278);
nand U1128 (N_1128,In_679,In_974);
or U1129 (N_1129,In_270,In_172);
xor U1130 (N_1130,In_320,In_691);
xor U1131 (N_1131,In_360,In_372);
nor U1132 (N_1132,In_130,In_257);
and U1133 (N_1133,In_154,In_590);
nor U1134 (N_1134,In_557,In_138);
xnor U1135 (N_1135,In_241,In_254);
and U1136 (N_1136,In_57,In_829);
nor U1137 (N_1137,In_86,In_342);
xnor U1138 (N_1138,In_670,In_73);
and U1139 (N_1139,In_591,In_605);
nand U1140 (N_1140,In_212,In_27);
or U1141 (N_1141,In_544,In_420);
or U1142 (N_1142,In_781,In_25);
nor U1143 (N_1143,In_412,In_857);
or U1144 (N_1144,In_11,In_897);
and U1145 (N_1145,In_386,In_876);
nand U1146 (N_1146,In_814,In_872);
nand U1147 (N_1147,In_303,In_297);
nor U1148 (N_1148,In_251,In_478);
xor U1149 (N_1149,In_836,In_487);
nand U1150 (N_1150,In_939,In_595);
nand U1151 (N_1151,In_316,In_857);
nand U1152 (N_1152,In_484,In_190);
nor U1153 (N_1153,In_28,In_905);
nor U1154 (N_1154,In_553,In_422);
nand U1155 (N_1155,In_597,In_671);
and U1156 (N_1156,In_961,In_49);
nor U1157 (N_1157,In_650,In_823);
or U1158 (N_1158,In_697,In_708);
nor U1159 (N_1159,In_940,In_443);
nor U1160 (N_1160,In_183,In_799);
or U1161 (N_1161,In_272,In_149);
nand U1162 (N_1162,In_23,In_368);
or U1163 (N_1163,In_155,In_514);
and U1164 (N_1164,In_809,In_392);
or U1165 (N_1165,In_386,In_947);
and U1166 (N_1166,In_727,In_491);
nand U1167 (N_1167,In_934,In_32);
nor U1168 (N_1168,In_445,In_373);
nand U1169 (N_1169,In_927,In_317);
or U1170 (N_1170,In_445,In_613);
or U1171 (N_1171,In_121,In_147);
nor U1172 (N_1172,In_15,In_546);
or U1173 (N_1173,In_61,In_975);
nand U1174 (N_1174,In_876,In_236);
nand U1175 (N_1175,In_961,In_446);
xnor U1176 (N_1176,In_118,In_47);
and U1177 (N_1177,In_427,In_59);
and U1178 (N_1178,In_919,In_691);
xnor U1179 (N_1179,In_263,In_96);
or U1180 (N_1180,In_204,In_84);
nor U1181 (N_1181,In_711,In_151);
and U1182 (N_1182,In_86,In_572);
nor U1183 (N_1183,In_466,In_492);
nand U1184 (N_1184,In_175,In_64);
or U1185 (N_1185,In_74,In_159);
or U1186 (N_1186,In_313,In_987);
nor U1187 (N_1187,In_565,In_456);
nand U1188 (N_1188,In_785,In_802);
nand U1189 (N_1189,In_799,In_379);
and U1190 (N_1190,In_238,In_418);
nor U1191 (N_1191,In_597,In_91);
nor U1192 (N_1192,In_482,In_396);
nor U1193 (N_1193,In_826,In_975);
or U1194 (N_1194,In_693,In_933);
nor U1195 (N_1195,In_859,In_462);
or U1196 (N_1196,In_87,In_63);
nand U1197 (N_1197,In_91,In_705);
or U1198 (N_1198,In_905,In_750);
xnor U1199 (N_1199,In_474,In_60);
nand U1200 (N_1200,In_659,In_473);
or U1201 (N_1201,In_783,In_204);
or U1202 (N_1202,In_492,In_354);
nand U1203 (N_1203,In_644,In_481);
or U1204 (N_1204,In_758,In_38);
or U1205 (N_1205,In_438,In_511);
nand U1206 (N_1206,In_890,In_304);
nor U1207 (N_1207,In_441,In_306);
and U1208 (N_1208,In_24,In_336);
and U1209 (N_1209,In_723,In_728);
nor U1210 (N_1210,In_252,In_396);
nand U1211 (N_1211,In_24,In_399);
nor U1212 (N_1212,In_915,In_762);
nand U1213 (N_1213,In_485,In_980);
and U1214 (N_1214,In_890,In_862);
nand U1215 (N_1215,In_182,In_445);
nand U1216 (N_1216,In_401,In_967);
and U1217 (N_1217,In_201,In_935);
or U1218 (N_1218,In_362,In_486);
or U1219 (N_1219,In_235,In_441);
nand U1220 (N_1220,In_425,In_420);
nand U1221 (N_1221,In_955,In_508);
or U1222 (N_1222,In_473,In_894);
xor U1223 (N_1223,In_805,In_611);
or U1224 (N_1224,In_637,In_717);
or U1225 (N_1225,In_51,In_782);
nor U1226 (N_1226,In_124,In_909);
nand U1227 (N_1227,In_15,In_66);
xor U1228 (N_1228,In_52,In_458);
nor U1229 (N_1229,In_366,In_131);
xnor U1230 (N_1230,In_697,In_71);
nor U1231 (N_1231,In_442,In_246);
nand U1232 (N_1232,In_749,In_244);
nor U1233 (N_1233,In_89,In_253);
and U1234 (N_1234,In_152,In_603);
nand U1235 (N_1235,In_746,In_40);
nor U1236 (N_1236,In_136,In_518);
nand U1237 (N_1237,In_536,In_905);
nor U1238 (N_1238,In_260,In_202);
nor U1239 (N_1239,In_791,In_480);
nand U1240 (N_1240,In_578,In_629);
nor U1241 (N_1241,In_805,In_208);
nand U1242 (N_1242,In_69,In_781);
nand U1243 (N_1243,In_945,In_696);
nor U1244 (N_1244,In_569,In_843);
xnor U1245 (N_1245,In_126,In_854);
and U1246 (N_1246,In_685,In_721);
and U1247 (N_1247,In_516,In_228);
and U1248 (N_1248,In_585,In_260);
nor U1249 (N_1249,In_758,In_276);
nor U1250 (N_1250,In_752,In_264);
nand U1251 (N_1251,In_202,In_143);
xor U1252 (N_1252,In_838,In_211);
or U1253 (N_1253,In_28,In_214);
or U1254 (N_1254,In_104,In_335);
nand U1255 (N_1255,In_763,In_31);
and U1256 (N_1256,In_631,In_164);
nand U1257 (N_1257,In_435,In_876);
or U1258 (N_1258,In_434,In_315);
xor U1259 (N_1259,In_801,In_681);
nand U1260 (N_1260,In_563,In_656);
and U1261 (N_1261,In_399,In_818);
nor U1262 (N_1262,In_444,In_547);
or U1263 (N_1263,In_861,In_452);
and U1264 (N_1264,In_224,In_826);
nand U1265 (N_1265,In_490,In_94);
nor U1266 (N_1266,In_540,In_385);
nand U1267 (N_1267,In_79,In_901);
nand U1268 (N_1268,In_327,In_858);
nand U1269 (N_1269,In_737,In_143);
nand U1270 (N_1270,In_56,In_340);
nand U1271 (N_1271,In_889,In_693);
nor U1272 (N_1272,In_723,In_367);
or U1273 (N_1273,In_201,In_856);
or U1274 (N_1274,In_322,In_668);
and U1275 (N_1275,In_951,In_427);
xor U1276 (N_1276,In_328,In_561);
and U1277 (N_1277,In_990,In_974);
nand U1278 (N_1278,In_822,In_210);
xnor U1279 (N_1279,In_730,In_276);
nand U1280 (N_1280,In_811,In_379);
or U1281 (N_1281,In_426,In_400);
nor U1282 (N_1282,In_442,In_162);
nand U1283 (N_1283,In_169,In_73);
nand U1284 (N_1284,In_57,In_946);
or U1285 (N_1285,In_604,In_156);
and U1286 (N_1286,In_250,In_713);
nand U1287 (N_1287,In_144,In_186);
and U1288 (N_1288,In_636,In_149);
nor U1289 (N_1289,In_578,In_916);
and U1290 (N_1290,In_370,In_1);
nor U1291 (N_1291,In_660,In_729);
xnor U1292 (N_1292,In_398,In_968);
or U1293 (N_1293,In_373,In_213);
or U1294 (N_1294,In_432,In_852);
nand U1295 (N_1295,In_267,In_94);
or U1296 (N_1296,In_76,In_595);
nand U1297 (N_1297,In_240,In_798);
nand U1298 (N_1298,In_854,In_856);
xor U1299 (N_1299,In_790,In_161);
nor U1300 (N_1300,In_98,In_409);
nor U1301 (N_1301,In_634,In_882);
nand U1302 (N_1302,In_521,In_772);
or U1303 (N_1303,In_60,In_975);
xor U1304 (N_1304,In_348,In_383);
or U1305 (N_1305,In_646,In_133);
nor U1306 (N_1306,In_443,In_15);
xnor U1307 (N_1307,In_865,In_120);
nand U1308 (N_1308,In_331,In_956);
nand U1309 (N_1309,In_66,In_9);
and U1310 (N_1310,In_710,In_666);
nand U1311 (N_1311,In_523,In_629);
nand U1312 (N_1312,In_806,In_605);
nor U1313 (N_1313,In_429,In_993);
and U1314 (N_1314,In_337,In_191);
or U1315 (N_1315,In_148,In_585);
nand U1316 (N_1316,In_52,In_540);
or U1317 (N_1317,In_257,In_7);
nand U1318 (N_1318,In_547,In_658);
nand U1319 (N_1319,In_721,In_324);
nand U1320 (N_1320,In_113,In_222);
nor U1321 (N_1321,In_526,In_825);
nand U1322 (N_1322,In_403,In_800);
or U1323 (N_1323,In_491,In_229);
and U1324 (N_1324,In_613,In_865);
nand U1325 (N_1325,In_260,In_308);
and U1326 (N_1326,In_923,In_21);
and U1327 (N_1327,In_869,In_160);
nor U1328 (N_1328,In_238,In_889);
or U1329 (N_1329,In_90,In_841);
and U1330 (N_1330,In_494,In_540);
nor U1331 (N_1331,In_59,In_89);
and U1332 (N_1332,In_859,In_287);
nor U1333 (N_1333,In_8,In_776);
xnor U1334 (N_1334,In_616,In_756);
xor U1335 (N_1335,In_604,In_516);
nor U1336 (N_1336,In_75,In_440);
and U1337 (N_1337,In_868,In_75);
nand U1338 (N_1338,In_53,In_879);
nand U1339 (N_1339,In_968,In_360);
and U1340 (N_1340,In_625,In_877);
nor U1341 (N_1341,In_882,In_507);
and U1342 (N_1342,In_663,In_479);
nand U1343 (N_1343,In_5,In_393);
nand U1344 (N_1344,In_70,In_717);
nor U1345 (N_1345,In_130,In_868);
or U1346 (N_1346,In_337,In_325);
nor U1347 (N_1347,In_863,In_848);
or U1348 (N_1348,In_880,In_137);
nand U1349 (N_1349,In_106,In_680);
nor U1350 (N_1350,In_199,In_172);
nand U1351 (N_1351,In_535,In_184);
nand U1352 (N_1352,In_503,In_182);
xor U1353 (N_1353,In_149,In_542);
nor U1354 (N_1354,In_611,In_750);
nor U1355 (N_1355,In_342,In_349);
or U1356 (N_1356,In_30,In_696);
nor U1357 (N_1357,In_887,In_964);
and U1358 (N_1358,In_869,In_123);
nand U1359 (N_1359,In_785,In_106);
and U1360 (N_1360,In_302,In_158);
nor U1361 (N_1361,In_850,In_287);
nand U1362 (N_1362,In_567,In_515);
nand U1363 (N_1363,In_287,In_773);
and U1364 (N_1364,In_718,In_564);
nor U1365 (N_1365,In_261,In_987);
or U1366 (N_1366,In_211,In_708);
or U1367 (N_1367,In_309,In_374);
nor U1368 (N_1368,In_717,In_244);
nand U1369 (N_1369,In_686,In_423);
or U1370 (N_1370,In_672,In_181);
and U1371 (N_1371,In_665,In_104);
nand U1372 (N_1372,In_432,In_972);
and U1373 (N_1373,In_903,In_873);
nand U1374 (N_1374,In_279,In_258);
or U1375 (N_1375,In_207,In_901);
and U1376 (N_1376,In_15,In_862);
or U1377 (N_1377,In_819,In_716);
nand U1378 (N_1378,In_868,In_460);
nor U1379 (N_1379,In_675,In_646);
nand U1380 (N_1380,In_195,In_541);
xor U1381 (N_1381,In_884,In_763);
or U1382 (N_1382,In_968,In_314);
nand U1383 (N_1383,In_816,In_856);
nor U1384 (N_1384,In_814,In_64);
and U1385 (N_1385,In_125,In_428);
nand U1386 (N_1386,In_721,In_825);
and U1387 (N_1387,In_494,In_850);
nor U1388 (N_1388,In_671,In_967);
nor U1389 (N_1389,In_791,In_219);
nor U1390 (N_1390,In_676,In_256);
nand U1391 (N_1391,In_624,In_847);
or U1392 (N_1392,In_187,In_659);
nand U1393 (N_1393,In_28,In_861);
or U1394 (N_1394,In_143,In_265);
and U1395 (N_1395,In_662,In_402);
xor U1396 (N_1396,In_201,In_259);
and U1397 (N_1397,In_643,In_586);
nand U1398 (N_1398,In_323,In_62);
xnor U1399 (N_1399,In_302,In_851);
nand U1400 (N_1400,In_800,In_776);
or U1401 (N_1401,In_198,In_98);
and U1402 (N_1402,In_414,In_658);
nor U1403 (N_1403,In_519,In_118);
or U1404 (N_1404,In_553,In_544);
nor U1405 (N_1405,In_244,In_560);
xnor U1406 (N_1406,In_758,In_367);
or U1407 (N_1407,In_695,In_657);
nand U1408 (N_1408,In_523,In_828);
and U1409 (N_1409,In_529,In_409);
xnor U1410 (N_1410,In_122,In_795);
xor U1411 (N_1411,In_797,In_60);
or U1412 (N_1412,In_457,In_980);
nor U1413 (N_1413,In_670,In_846);
xor U1414 (N_1414,In_785,In_369);
nor U1415 (N_1415,In_80,In_646);
xnor U1416 (N_1416,In_123,In_496);
nand U1417 (N_1417,In_199,In_205);
nand U1418 (N_1418,In_765,In_812);
or U1419 (N_1419,In_212,In_607);
and U1420 (N_1420,In_362,In_882);
nand U1421 (N_1421,In_110,In_650);
nor U1422 (N_1422,In_174,In_534);
nand U1423 (N_1423,In_686,In_785);
nor U1424 (N_1424,In_476,In_806);
nand U1425 (N_1425,In_527,In_538);
or U1426 (N_1426,In_929,In_471);
or U1427 (N_1427,In_770,In_900);
or U1428 (N_1428,In_618,In_537);
and U1429 (N_1429,In_192,In_560);
and U1430 (N_1430,In_425,In_823);
or U1431 (N_1431,In_477,In_653);
and U1432 (N_1432,In_972,In_728);
nor U1433 (N_1433,In_869,In_725);
or U1434 (N_1434,In_945,In_239);
nor U1435 (N_1435,In_347,In_189);
or U1436 (N_1436,In_496,In_0);
or U1437 (N_1437,In_980,In_454);
nand U1438 (N_1438,In_582,In_111);
and U1439 (N_1439,In_301,In_90);
and U1440 (N_1440,In_573,In_68);
nor U1441 (N_1441,In_685,In_227);
xnor U1442 (N_1442,In_116,In_850);
nor U1443 (N_1443,In_329,In_999);
and U1444 (N_1444,In_481,In_389);
nor U1445 (N_1445,In_13,In_898);
nor U1446 (N_1446,In_766,In_888);
nand U1447 (N_1447,In_456,In_762);
nand U1448 (N_1448,In_254,In_142);
xor U1449 (N_1449,In_862,In_665);
or U1450 (N_1450,In_276,In_732);
nor U1451 (N_1451,In_300,In_72);
nand U1452 (N_1452,In_967,In_526);
or U1453 (N_1453,In_242,In_388);
or U1454 (N_1454,In_614,In_957);
or U1455 (N_1455,In_767,In_245);
or U1456 (N_1456,In_64,In_384);
and U1457 (N_1457,In_566,In_282);
nor U1458 (N_1458,In_743,In_474);
nand U1459 (N_1459,In_192,In_670);
nor U1460 (N_1460,In_258,In_817);
nor U1461 (N_1461,In_535,In_265);
and U1462 (N_1462,In_571,In_952);
nand U1463 (N_1463,In_639,In_357);
and U1464 (N_1464,In_469,In_697);
nand U1465 (N_1465,In_935,In_910);
nand U1466 (N_1466,In_766,In_388);
nand U1467 (N_1467,In_603,In_278);
nand U1468 (N_1468,In_718,In_581);
and U1469 (N_1469,In_561,In_57);
or U1470 (N_1470,In_619,In_458);
and U1471 (N_1471,In_649,In_433);
or U1472 (N_1472,In_103,In_766);
nor U1473 (N_1473,In_443,In_478);
or U1474 (N_1474,In_741,In_92);
or U1475 (N_1475,In_882,In_745);
xnor U1476 (N_1476,In_74,In_586);
nor U1477 (N_1477,In_376,In_403);
and U1478 (N_1478,In_760,In_845);
nor U1479 (N_1479,In_531,In_888);
or U1480 (N_1480,In_91,In_143);
nor U1481 (N_1481,In_651,In_536);
and U1482 (N_1482,In_97,In_145);
nor U1483 (N_1483,In_205,In_144);
nor U1484 (N_1484,In_595,In_412);
nand U1485 (N_1485,In_87,In_673);
and U1486 (N_1486,In_529,In_47);
nand U1487 (N_1487,In_164,In_706);
or U1488 (N_1488,In_42,In_124);
and U1489 (N_1489,In_201,In_737);
and U1490 (N_1490,In_432,In_684);
and U1491 (N_1491,In_416,In_338);
or U1492 (N_1492,In_899,In_310);
and U1493 (N_1493,In_484,In_870);
nor U1494 (N_1494,In_270,In_62);
nand U1495 (N_1495,In_868,In_254);
nand U1496 (N_1496,In_584,In_546);
and U1497 (N_1497,In_800,In_729);
nand U1498 (N_1498,In_863,In_876);
or U1499 (N_1499,In_293,In_523);
or U1500 (N_1500,In_276,In_941);
nor U1501 (N_1501,In_757,In_64);
nor U1502 (N_1502,In_507,In_156);
nand U1503 (N_1503,In_836,In_254);
or U1504 (N_1504,In_203,In_677);
and U1505 (N_1505,In_398,In_55);
or U1506 (N_1506,In_817,In_748);
nor U1507 (N_1507,In_351,In_746);
nand U1508 (N_1508,In_554,In_531);
xnor U1509 (N_1509,In_190,In_639);
xnor U1510 (N_1510,In_403,In_180);
xnor U1511 (N_1511,In_20,In_582);
xor U1512 (N_1512,In_925,In_56);
nor U1513 (N_1513,In_954,In_191);
nand U1514 (N_1514,In_341,In_820);
nor U1515 (N_1515,In_544,In_648);
or U1516 (N_1516,In_87,In_382);
and U1517 (N_1517,In_323,In_741);
and U1518 (N_1518,In_259,In_418);
nand U1519 (N_1519,In_501,In_571);
nor U1520 (N_1520,In_972,In_217);
or U1521 (N_1521,In_4,In_41);
and U1522 (N_1522,In_730,In_944);
nand U1523 (N_1523,In_211,In_542);
and U1524 (N_1524,In_615,In_774);
and U1525 (N_1525,In_614,In_203);
or U1526 (N_1526,In_575,In_927);
and U1527 (N_1527,In_242,In_18);
and U1528 (N_1528,In_929,In_904);
or U1529 (N_1529,In_602,In_529);
or U1530 (N_1530,In_130,In_344);
or U1531 (N_1531,In_929,In_355);
nand U1532 (N_1532,In_654,In_27);
nor U1533 (N_1533,In_573,In_346);
nor U1534 (N_1534,In_580,In_31);
xor U1535 (N_1535,In_39,In_919);
nor U1536 (N_1536,In_152,In_453);
and U1537 (N_1537,In_734,In_474);
nor U1538 (N_1538,In_505,In_122);
and U1539 (N_1539,In_150,In_606);
and U1540 (N_1540,In_18,In_283);
nand U1541 (N_1541,In_842,In_570);
or U1542 (N_1542,In_955,In_335);
and U1543 (N_1543,In_313,In_223);
and U1544 (N_1544,In_294,In_670);
and U1545 (N_1545,In_971,In_660);
or U1546 (N_1546,In_281,In_75);
nor U1547 (N_1547,In_255,In_542);
or U1548 (N_1548,In_274,In_763);
or U1549 (N_1549,In_818,In_63);
and U1550 (N_1550,In_352,In_122);
nor U1551 (N_1551,In_971,In_470);
and U1552 (N_1552,In_421,In_803);
nor U1553 (N_1553,In_107,In_253);
or U1554 (N_1554,In_311,In_154);
nand U1555 (N_1555,In_836,In_943);
xor U1556 (N_1556,In_810,In_3);
or U1557 (N_1557,In_132,In_272);
nor U1558 (N_1558,In_962,In_242);
xnor U1559 (N_1559,In_484,In_964);
or U1560 (N_1560,In_32,In_364);
or U1561 (N_1561,In_950,In_295);
nand U1562 (N_1562,In_524,In_271);
nor U1563 (N_1563,In_989,In_827);
nor U1564 (N_1564,In_798,In_709);
nor U1565 (N_1565,In_90,In_981);
or U1566 (N_1566,In_33,In_159);
or U1567 (N_1567,In_709,In_98);
nor U1568 (N_1568,In_524,In_283);
nand U1569 (N_1569,In_599,In_986);
nand U1570 (N_1570,In_532,In_993);
or U1571 (N_1571,In_582,In_633);
or U1572 (N_1572,In_143,In_123);
and U1573 (N_1573,In_295,In_278);
nand U1574 (N_1574,In_355,In_120);
nor U1575 (N_1575,In_323,In_272);
nor U1576 (N_1576,In_276,In_15);
or U1577 (N_1577,In_324,In_220);
and U1578 (N_1578,In_152,In_821);
xnor U1579 (N_1579,In_340,In_312);
and U1580 (N_1580,In_767,In_244);
or U1581 (N_1581,In_626,In_406);
nor U1582 (N_1582,In_620,In_832);
and U1583 (N_1583,In_104,In_823);
nand U1584 (N_1584,In_198,In_375);
nor U1585 (N_1585,In_125,In_716);
and U1586 (N_1586,In_750,In_267);
and U1587 (N_1587,In_256,In_219);
or U1588 (N_1588,In_435,In_4);
nor U1589 (N_1589,In_772,In_493);
nand U1590 (N_1590,In_200,In_494);
nand U1591 (N_1591,In_163,In_355);
nor U1592 (N_1592,In_706,In_354);
or U1593 (N_1593,In_429,In_385);
nor U1594 (N_1594,In_915,In_928);
nor U1595 (N_1595,In_939,In_394);
and U1596 (N_1596,In_794,In_402);
nand U1597 (N_1597,In_159,In_895);
or U1598 (N_1598,In_932,In_983);
or U1599 (N_1599,In_813,In_896);
nor U1600 (N_1600,In_48,In_781);
or U1601 (N_1601,In_48,In_855);
and U1602 (N_1602,In_574,In_378);
nor U1603 (N_1603,In_413,In_283);
nand U1604 (N_1604,In_344,In_282);
and U1605 (N_1605,In_804,In_971);
or U1606 (N_1606,In_399,In_822);
nand U1607 (N_1607,In_53,In_43);
nor U1608 (N_1608,In_640,In_152);
nand U1609 (N_1609,In_904,In_112);
or U1610 (N_1610,In_223,In_465);
nand U1611 (N_1611,In_715,In_589);
or U1612 (N_1612,In_780,In_228);
xor U1613 (N_1613,In_201,In_681);
xnor U1614 (N_1614,In_571,In_289);
nor U1615 (N_1615,In_349,In_99);
nand U1616 (N_1616,In_635,In_839);
nor U1617 (N_1617,In_264,In_565);
nand U1618 (N_1618,In_929,In_347);
and U1619 (N_1619,In_610,In_263);
or U1620 (N_1620,In_257,In_467);
and U1621 (N_1621,In_381,In_919);
or U1622 (N_1622,In_861,In_294);
nor U1623 (N_1623,In_292,In_736);
nor U1624 (N_1624,In_952,In_720);
and U1625 (N_1625,In_769,In_517);
and U1626 (N_1626,In_948,In_732);
nand U1627 (N_1627,In_256,In_370);
or U1628 (N_1628,In_956,In_29);
nand U1629 (N_1629,In_419,In_774);
nand U1630 (N_1630,In_81,In_360);
nor U1631 (N_1631,In_474,In_850);
and U1632 (N_1632,In_979,In_356);
xor U1633 (N_1633,In_575,In_694);
or U1634 (N_1634,In_296,In_84);
nor U1635 (N_1635,In_156,In_537);
nand U1636 (N_1636,In_610,In_27);
nor U1637 (N_1637,In_192,In_128);
or U1638 (N_1638,In_652,In_289);
and U1639 (N_1639,In_531,In_754);
or U1640 (N_1640,In_933,In_386);
nor U1641 (N_1641,In_583,In_810);
nor U1642 (N_1642,In_394,In_38);
nor U1643 (N_1643,In_141,In_874);
and U1644 (N_1644,In_246,In_992);
or U1645 (N_1645,In_264,In_581);
or U1646 (N_1646,In_865,In_844);
and U1647 (N_1647,In_740,In_567);
nor U1648 (N_1648,In_656,In_212);
or U1649 (N_1649,In_270,In_710);
nor U1650 (N_1650,In_833,In_699);
nand U1651 (N_1651,In_456,In_507);
xor U1652 (N_1652,In_125,In_861);
or U1653 (N_1653,In_866,In_285);
and U1654 (N_1654,In_548,In_731);
or U1655 (N_1655,In_160,In_333);
nor U1656 (N_1656,In_372,In_950);
xnor U1657 (N_1657,In_182,In_94);
nor U1658 (N_1658,In_620,In_314);
or U1659 (N_1659,In_590,In_65);
and U1660 (N_1660,In_58,In_342);
nor U1661 (N_1661,In_494,In_38);
nor U1662 (N_1662,In_114,In_300);
nor U1663 (N_1663,In_370,In_981);
xor U1664 (N_1664,In_431,In_633);
and U1665 (N_1665,In_8,In_622);
nand U1666 (N_1666,In_569,In_632);
nor U1667 (N_1667,In_353,In_381);
nand U1668 (N_1668,In_362,In_666);
nand U1669 (N_1669,In_982,In_320);
nand U1670 (N_1670,In_441,In_97);
nor U1671 (N_1671,In_940,In_104);
nor U1672 (N_1672,In_99,In_616);
nand U1673 (N_1673,In_732,In_222);
or U1674 (N_1674,In_208,In_894);
nand U1675 (N_1675,In_640,In_610);
and U1676 (N_1676,In_924,In_548);
and U1677 (N_1677,In_269,In_914);
and U1678 (N_1678,In_606,In_659);
or U1679 (N_1679,In_5,In_779);
or U1680 (N_1680,In_760,In_343);
nor U1681 (N_1681,In_863,In_933);
nand U1682 (N_1682,In_239,In_135);
nand U1683 (N_1683,In_341,In_527);
or U1684 (N_1684,In_623,In_694);
xor U1685 (N_1685,In_703,In_847);
and U1686 (N_1686,In_69,In_587);
xnor U1687 (N_1687,In_70,In_884);
nor U1688 (N_1688,In_225,In_783);
nor U1689 (N_1689,In_439,In_146);
or U1690 (N_1690,In_789,In_320);
and U1691 (N_1691,In_463,In_163);
or U1692 (N_1692,In_540,In_851);
or U1693 (N_1693,In_133,In_618);
nand U1694 (N_1694,In_862,In_437);
or U1695 (N_1695,In_76,In_856);
or U1696 (N_1696,In_772,In_195);
and U1697 (N_1697,In_34,In_342);
nand U1698 (N_1698,In_28,In_304);
or U1699 (N_1699,In_693,In_286);
or U1700 (N_1700,In_163,In_541);
xor U1701 (N_1701,In_312,In_897);
xor U1702 (N_1702,In_538,In_490);
nor U1703 (N_1703,In_30,In_344);
or U1704 (N_1704,In_553,In_313);
and U1705 (N_1705,In_909,In_497);
or U1706 (N_1706,In_503,In_303);
nand U1707 (N_1707,In_851,In_643);
and U1708 (N_1708,In_821,In_698);
or U1709 (N_1709,In_689,In_621);
and U1710 (N_1710,In_35,In_375);
and U1711 (N_1711,In_59,In_408);
xor U1712 (N_1712,In_900,In_328);
xor U1713 (N_1713,In_80,In_45);
nand U1714 (N_1714,In_461,In_57);
and U1715 (N_1715,In_681,In_651);
xor U1716 (N_1716,In_544,In_124);
or U1717 (N_1717,In_862,In_289);
nand U1718 (N_1718,In_943,In_494);
nand U1719 (N_1719,In_957,In_804);
nor U1720 (N_1720,In_462,In_460);
and U1721 (N_1721,In_932,In_947);
or U1722 (N_1722,In_511,In_585);
or U1723 (N_1723,In_253,In_568);
nor U1724 (N_1724,In_497,In_257);
nor U1725 (N_1725,In_756,In_284);
nand U1726 (N_1726,In_303,In_992);
nor U1727 (N_1727,In_361,In_322);
or U1728 (N_1728,In_893,In_70);
nor U1729 (N_1729,In_755,In_218);
xor U1730 (N_1730,In_232,In_211);
and U1731 (N_1731,In_224,In_664);
nor U1732 (N_1732,In_42,In_445);
nor U1733 (N_1733,In_237,In_915);
or U1734 (N_1734,In_423,In_753);
nand U1735 (N_1735,In_708,In_955);
nand U1736 (N_1736,In_190,In_722);
and U1737 (N_1737,In_710,In_751);
and U1738 (N_1738,In_542,In_119);
nor U1739 (N_1739,In_146,In_264);
nor U1740 (N_1740,In_99,In_149);
or U1741 (N_1741,In_378,In_859);
or U1742 (N_1742,In_788,In_951);
nor U1743 (N_1743,In_346,In_998);
nor U1744 (N_1744,In_802,In_801);
nand U1745 (N_1745,In_671,In_530);
xnor U1746 (N_1746,In_831,In_9);
xnor U1747 (N_1747,In_123,In_586);
nor U1748 (N_1748,In_87,In_531);
nand U1749 (N_1749,In_630,In_645);
and U1750 (N_1750,In_603,In_73);
or U1751 (N_1751,In_898,In_967);
nand U1752 (N_1752,In_347,In_366);
xor U1753 (N_1753,In_65,In_88);
or U1754 (N_1754,In_358,In_660);
or U1755 (N_1755,In_355,In_603);
or U1756 (N_1756,In_748,In_359);
and U1757 (N_1757,In_935,In_154);
nor U1758 (N_1758,In_173,In_921);
nand U1759 (N_1759,In_690,In_310);
nand U1760 (N_1760,In_429,In_447);
and U1761 (N_1761,In_793,In_43);
and U1762 (N_1762,In_53,In_55);
nor U1763 (N_1763,In_728,In_604);
or U1764 (N_1764,In_46,In_607);
and U1765 (N_1765,In_73,In_337);
or U1766 (N_1766,In_769,In_133);
nand U1767 (N_1767,In_720,In_165);
nor U1768 (N_1768,In_804,In_583);
and U1769 (N_1769,In_920,In_647);
nand U1770 (N_1770,In_902,In_68);
and U1771 (N_1771,In_289,In_672);
nand U1772 (N_1772,In_119,In_360);
or U1773 (N_1773,In_583,In_662);
nand U1774 (N_1774,In_11,In_807);
nand U1775 (N_1775,In_139,In_106);
nor U1776 (N_1776,In_137,In_879);
or U1777 (N_1777,In_201,In_197);
nor U1778 (N_1778,In_662,In_911);
and U1779 (N_1779,In_881,In_74);
and U1780 (N_1780,In_650,In_570);
or U1781 (N_1781,In_766,In_917);
or U1782 (N_1782,In_856,In_101);
nand U1783 (N_1783,In_893,In_955);
nand U1784 (N_1784,In_542,In_792);
and U1785 (N_1785,In_346,In_95);
xnor U1786 (N_1786,In_485,In_278);
or U1787 (N_1787,In_419,In_145);
nand U1788 (N_1788,In_955,In_700);
nand U1789 (N_1789,In_963,In_950);
nand U1790 (N_1790,In_393,In_842);
or U1791 (N_1791,In_269,In_633);
nor U1792 (N_1792,In_190,In_598);
nor U1793 (N_1793,In_126,In_460);
and U1794 (N_1794,In_146,In_205);
or U1795 (N_1795,In_138,In_605);
or U1796 (N_1796,In_71,In_535);
and U1797 (N_1797,In_212,In_44);
nand U1798 (N_1798,In_577,In_385);
nor U1799 (N_1799,In_592,In_434);
nand U1800 (N_1800,In_236,In_38);
nor U1801 (N_1801,In_103,In_308);
and U1802 (N_1802,In_911,In_400);
or U1803 (N_1803,In_554,In_433);
nor U1804 (N_1804,In_47,In_286);
and U1805 (N_1805,In_371,In_696);
nor U1806 (N_1806,In_183,In_72);
and U1807 (N_1807,In_123,In_865);
and U1808 (N_1808,In_839,In_130);
nor U1809 (N_1809,In_355,In_19);
nand U1810 (N_1810,In_244,In_499);
or U1811 (N_1811,In_591,In_742);
xor U1812 (N_1812,In_655,In_408);
xnor U1813 (N_1813,In_559,In_964);
nand U1814 (N_1814,In_319,In_853);
nor U1815 (N_1815,In_53,In_539);
and U1816 (N_1816,In_211,In_208);
or U1817 (N_1817,In_652,In_507);
or U1818 (N_1818,In_865,In_19);
xnor U1819 (N_1819,In_468,In_193);
xnor U1820 (N_1820,In_744,In_775);
xnor U1821 (N_1821,In_568,In_685);
nand U1822 (N_1822,In_395,In_821);
xor U1823 (N_1823,In_63,In_14);
xnor U1824 (N_1824,In_967,In_29);
nor U1825 (N_1825,In_292,In_973);
or U1826 (N_1826,In_475,In_154);
and U1827 (N_1827,In_850,In_685);
or U1828 (N_1828,In_117,In_854);
nand U1829 (N_1829,In_972,In_448);
or U1830 (N_1830,In_61,In_978);
or U1831 (N_1831,In_949,In_897);
nand U1832 (N_1832,In_982,In_523);
and U1833 (N_1833,In_907,In_984);
nand U1834 (N_1834,In_562,In_698);
xnor U1835 (N_1835,In_575,In_476);
or U1836 (N_1836,In_409,In_149);
and U1837 (N_1837,In_403,In_214);
and U1838 (N_1838,In_18,In_268);
nor U1839 (N_1839,In_731,In_728);
and U1840 (N_1840,In_173,In_706);
nand U1841 (N_1841,In_757,In_27);
or U1842 (N_1842,In_239,In_702);
or U1843 (N_1843,In_327,In_780);
xor U1844 (N_1844,In_688,In_800);
xnor U1845 (N_1845,In_282,In_541);
or U1846 (N_1846,In_282,In_688);
nand U1847 (N_1847,In_332,In_441);
or U1848 (N_1848,In_991,In_677);
nand U1849 (N_1849,In_118,In_27);
or U1850 (N_1850,In_591,In_201);
nor U1851 (N_1851,In_251,In_377);
nand U1852 (N_1852,In_599,In_628);
and U1853 (N_1853,In_201,In_389);
nand U1854 (N_1854,In_764,In_180);
nand U1855 (N_1855,In_503,In_560);
nand U1856 (N_1856,In_389,In_20);
nand U1857 (N_1857,In_609,In_635);
or U1858 (N_1858,In_621,In_54);
and U1859 (N_1859,In_574,In_374);
or U1860 (N_1860,In_790,In_70);
nor U1861 (N_1861,In_570,In_573);
nor U1862 (N_1862,In_192,In_97);
nor U1863 (N_1863,In_52,In_619);
nor U1864 (N_1864,In_810,In_783);
or U1865 (N_1865,In_862,In_224);
and U1866 (N_1866,In_688,In_312);
or U1867 (N_1867,In_317,In_3);
and U1868 (N_1868,In_234,In_383);
or U1869 (N_1869,In_309,In_953);
nor U1870 (N_1870,In_283,In_784);
nand U1871 (N_1871,In_976,In_750);
nor U1872 (N_1872,In_180,In_898);
or U1873 (N_1873,In_897,In_482);
nor U1874 (N_1874,In_211,In_787);
nor U1875 (N_1875,In_775,In_491);
xor U1876 (N_1876,In_345,In_523);
and U1877 (N_1877,In_604,In_285);
nand U1878 (N_1878,In_881,In_763);
nand U1879 (N_1879,In_118,In_158);
nand U1880 (N_1880,In_352,In_414);
or U1881 (N_1881,In_220,In_928);
nand U1882 (N_1882,In_538,In_608);
or U1883 (N_1883,In_204,In_387);
and U1884 (N_1884,In_428,In_643);
nor U1885 (N_1885,In_51,In_866);
or U1886 (N_1886,In_221,In_742);
and U1887 (N_1887,In_748,In_550);
or U1888 (N_1888,In_364,In_978);
nand U1889 (N_1889,In_129,In_36);
or U1890 (N_1890,In_965,In_325);
or U1891 (N_1891,In_588,In_702);
nor U1892 (N_1892,In_164,In_323);
or U1893 (N_1893,In_92,In_437);
or U1894 (N_1894,In_504,In_364);
nor U1895 (N_1895,In_809,In_301);
nand U1896 (N_1896,In_559,In_990);
nand U1897 (N_1897,In_116,In_483);
nor U1898 (N_1898,In_522,In_171);
nand U1899 (N_1899,In_793,In_271);
or U1900 (N_1900,In_771,In_117);
or U1901 (N_1901,In_637,In_650);
nor U1902 (N_1902,In_667,In_195);
nor U1903 (N_1903,In_678,In_667);
or U1904 (N_1904,In_280,In_484);
xor U1905 (N_1905,In_143,In_546);
nor U1906 (N_1906,In_24,In_49);
xor U1907 (N_1907,In_426,In_166);
or U1908 (N_1908,In_14,In_790);
nor U1909 (N_1909,In_453,In_590);
and U1910 (N_1910,In_175,In_448);
or U1911 (N_1911,In_582,In_807);
nor U1912 (N_1912,In_296,In_719);
and U1913 (N_1913,In_311,In_298);
nand U1914 (N_1914,In_954,In_632);
nor U1915 (N_1915,In_423,In_858);
nand U1916 (N_1916,In_785,In_114);
and U1917 (N_1917,In_259,In_728);
nand U1918 (N_1918,In_17,In_131);
or U1919 (N_1919,In_540,In_204);
nand U1920 (N_1920,In_255,In_213);
nand U1921 (N_1921,In_685,In_312);
nand U1922 (N_1922,In_521,In_29);
nand U1923 (N_1923,In_321,In_580);
xnor U1924 (N_1924,In_627,In_77);
and U1925 (N_1925,In_716,In_476);
and U1926 (N_1926,In_906,In_160);
nand U1927 (N_1927,In_494,In_74);
xor U1928 (N_1928,In_390,In_742);
nor U1929 (N_1929,In_937,In_472);
nand U1930 (N_1930,In_323,In_384);
and U1931 (N_1931,In_266,In_773);
or U1932 (N_1932,In_128,In_142);
nor U1933 (N_1933,In_171,In_787);
nand U1934 (N_1934,In_680,In_284);
or U1935 (N_1935,In_858,In_8);
nand U1936 (N_1936,In_295,In_124);
and U1937 (N_1937,In_765,In_762);
and U1938 (N_1938,In_862,In_534);
or U1939 (N_1939,In_528,In_2);
nand U1940 (N_1940,In_473,In_800);
nor U1941 (N_1941,In_491,In_782);
nor U1942 (N_1942,In_2,In_571);
and U1943 (N_1943,In_931,In_818);
nor U1944 (N_1944,In_119,In_309);
nand U1945 (N_1945,In_502,In_372);
or U1946 (N_1946,In_159,In_123);
or U1947 (N_1947,In_256,In_627);
and U1948 (N_1948,In_763,In_159);
or U1949 (N_1949,In_6,In_749);
and U1950 (N_1950,In_820,In_369);
or U1951 (N_1951,In_903,In_577);
nor U1952 (N_1952,In_566,In_459);
nor U1953 (N_1953,In_832,In_558);
nor U1954 (N_1954,In_907,In_84);
and U1955 (N_1955,In_888,In_426);
nand U1956 (N_1956,In_43,In_534);
or U1957 (N_1957,In_812,In_533);
and U1958 (N_1958,In_919,In_685);
nand U1959 (N_1959,In_872,In_17);
nor U1960 (N_1960,In_836,In_460);
or U1961 (N_1961,In_76,In_155);
nand U1962 (N_1962,In_519,In_159);
xor U1963 (N_1963,In_652,In_118);
nor U1964 (N_1964,In_680,In_749);
and U1965 (N_1965,In_14,In_546);
and U1966 (N_1966,In_575,In_407);
and U1967 (N_1967,In_424,In_681);
nor U1968 (N_1968,In_968,In_108);
nand U1969 (N_1969,In_602,In_422);
nor U1970 (N_1970,In_147,In_63);
and U1971 (N_1971,In_358,In_332);
xor U1972 (N_1972,In_107,In_551);
and U1973 (N_1973,In_406,In_840);
nor U1974 (N_1974,In_402,In_706);
or U1975 (N_1975,In_83,In_38);
nor U1976 (N_1976,In_192,In_713);
nor U1977 (N_1977,In_199,In_981);
nor U1978 (N_1978,In_340,In_466);
and U1979 (N_1979,In_36,In_196);
and U1980 (N_1980,In_945,In_647);
nand U1981 (N_1981,In_798,In_456);
nand U1982 (N_1982,In_601,In_103);
xnor U1983 (N_1983,In_49,In_39);
and U1984 (N_1984,In_89,In_454);
xor U1985 (N_1985,In_281,In_145);
and U1986 (N_1986,In_270,In_514);
and U1987 (N_1987,In_198,In_360);
xor U1988 (N_1988,In_403,In_961);
nand U1989 (N_1989,In_5,In_614);
nor U1990 (N_1990,In_915,In_611);
nand U1991 (N_1991,In_391,In_202);
and U1992 (N_1992,In_880,In_47);
and U1993 (N_1993,In_519,In_617);
nand U1994 (N_1994,In_767,In_187);
and U1995 (N_1995,In_624,In_53);
or U1996 (N_1996,In_262,In_144);
and U1997 (N_1997,In_373,In_856);
or U1998 (N_1998,In_25,In_437);
xor U1999 (N_1999,In_83,In_973);
and U2000 (N_2000,In_170,In_621);
nor U2001 (N_2001,In_238,In_788);
and U2002 (N_2002,In_831,In_490);
or U2003 (N_2003,In_963,In_253);
xor U2004 (N_2004,In_66,In_922);
or U2005 (N_2005,In_522,In_109);
or U2006 (N_2006,In_797,In_983);
or U2007 (N_2007,In_414,In_259);
nand U2008 (N_2008,In_320,In_230);
nor U2009 (N_2009,In_866,In_562);
xor U2010 (N_2010,In_252,In_241);
or U2011 (N_2011,In_798,In_830);
or U2012 (N_2012,In_618,In_152);
nor U2013 (N_2013,In_348,In_636);
and U2014 (N_2014,In_556,In_668);
and U2015 (N_2015,In_492,In_207);
or U2016 (N_2016,In_909,In_632);
nand U2017 (N_2017,In_417,In_216);
nor U2018 (N_2018,In_511,In_246);
or U2019 (N_2019,In_343,In_415);
xnor U2020 (N_2020,In_66,In_771);
and U2021 (N_2021,In_383,In_224);
or U2022 (N_2022,In_821,In_868);
nand U2023 (N_2023,In_857,In_106);
and U2024 (N_2024,In_166,In_580);
nor U2025 (N_2025,In_133,In_271);
or U2026 (N_2026,In_164,In_271);
or U2027 (N_2027,In_970,In_734);
or U2028 (N_2028,In_221,In_234);
or U2029 (N_2029,In_853,In_420);
nor U2030 (N_2030,In_22,In_264);
nor U2031 (N_2031,In_789,In_688);
or U2032 (N_2032,In_762,In_966);
nor U2033 (N_2033,In_364,In_100);
xnor U2034 (N_2034,In_679,In_800);
nor U2035 (N_2035,In_804,In_529);
or U2036 (N_2036,In_866,In_28);
nor U2037 (N_2037,In_943,In_112);
nand U2038 (N_2038,In_196,In_901);
or U2039 (N_2039,In_441,In_321);
or U2040 (N_2040,In_758,In_78);
nor U2041 (N_2041,In_512,In_290);
nand U2042 (N_2042,In_289,In_166);
nor U2043 (N_2043,In_34,In_992);
or U2044 (N_2044,In_764,In_352);
and U2045 (N_2045,In_316,In_328);
and U2046 (N_2046,In_589,In_240);
or U2047 (N_2047,In_324,In_986);
or U2048 (N_2048,In_217,In_449);
nor U2049 (N_2049,In_471,In_603);
or U2050 (N_2050,In_332,In_254);
nor U2051 (N_2051,In_903,In_289);
nor U2052 (N_2052,In_669,In_365);
nand U2053 (N_2053,In_76,In_242);
xnor U2054 (N_2054,In_690,In_925);
nor U2055 (N_2055,In_921,In_356);
nand U2056 (N_2056,In_556,In_76);
nand U2057 (N_2057,In_76,In_536);
nand U2058 (N_2058,In_972,In_880);
nand U2059 (N_2059,In_528,In_216);
nor U2060 (N_2060,In_888,In_620);
nand U2061 (N_2061,In_255,In_934);
and U2062 (N_2062,In_72,In_78);
nor U2063 (N_2063,In_362,In_832);
nand U2064 (N_2064,In_211,In_374);
nor U2065 (N_2065,In_149,In_8);
nor U2066 (N_2066,In_676,In_389);
xor U2067 (N_2067,In_633,In_198);
or U2068 (N_2068,In_524,In_911);
or U2069 (N_2069,In_523,In_198);
nor U2070 (N_2070,In_985,In_36);
or U2071 (N_2071,In_797,In_579);
or U2072 (N_2072,In_1,In_385);
nor U2073 (N_2073,In_428,In_529);
nor U2074 (N_2074,In_893,In_477);
nor U2075 (N_2075,In_504,In_452);
nand U2076 (N_2076,In_424,In_463);
xnor U2077 (N_2077,In_67,In_441);
nor U2078 (N_2078,In_527,In_882);
xor U2079 (N_2079,In_718,In_456);
nand U2080 (N_2080,In_53,In_762);
nor U2081 (N_2081,In_71,In_353);
and U2082 (N_2082,In_626,In_272);
or U2083 (N_2083,In_531,In_212);
and U2084 (N_2084,In_434,In_465);
or U2085 (N_2085,In_312,In_450);
nand U2086 (N_2086,In_962,In_530);
and U2087 (N_2087,In_887,In_969);
nand U2088 (N_2088,In_494,In_897);
nor U2089 (N_2089,In_450,In_299);
or U2090 (N_2090,In_295,In_992);
or U2091 (N_2091,In_98,In_833);
xor U2092 (N_2092,In_553,In_818);
or U2093 (N_2093,In_500,In_150);
nor U2094 (N_2094,In_627,In_267);
and U2095 (N_2095,In_521,In_443);
or U2096 (N_2096,In_889,In_224);
or U2097 (N_2097,In_701,In_340);
nand U2098 (N_2098,In_354,In_398);
and U2099 (N_2099,In_662,In_310);
or U2100 (N_2100,In_982,In_830);
and U2101 (N_2101,In_167,In_16);
and U2102 (N_2102,In_291,In_821);
and U2103 (N_2103,In_861,In_629);
xor U2104 (N_2104,In_933,In_983);
and U2105 (N_2105,In_378,In_2);
nand U2106 (N_2106,In_353,In_691);
xnor U2107 (N_2107,In_890,In_289);
nand U2108 (N_2108,In_246,In_510);
or U2109 (N_2109,In_221,In_356);
nor U2110 (N_2110,In_328,In_927);
nand U2111 (N_2111,In_486,In_829);
or U2112 (N_2112,In_451,In_59);
or U2113 (N_2113,In_429,In_235);
or U2114 (N_2114,In_739,In_563);
nand U2115 (N_2115,In_352,In_41);
nor U2116 (N_2116,In_695,In_681);
nand U2117 (N_2117,In_86,In_188);
nand U2118 (N_2118,In_855,In_305);
or U2119 (N_2119,In_541,In_389);
nor U2120 (N_2120,In_290,In_963);
nand U2121 (N_2121,In_680,In_289);
nand U2122 (N_2122,In_982,In_715);
nor U2123 (N_2123,In_309,In_655);
or U2124 (N_2124,In_921,In_150);
or U2125 (N_2125,In_107,In_460);
xnor U2126 (N_2126,In_646,In_345);
and U2127 (N_2127,In_53,In_332);
and U2128 (N_2128,In_715,In_463);
and U2129 (N_2129,In_848,In_578);
xor U2130 (N_2130,In_828,In_940);
nand U2131 (N_2131,In_847,In_944);
or U2132 (N_2132,In_725,In_239);
xor U2133 (N_2133,In_120,In_914);
or U2134 (N_2134,In_753,In_496);
or U2135 (N_2135,In_866,In_479);
xnor U2136 (N_2136,In_669,In_503);
nor U2137 (N_2137,In_382,In_914);
nor U2138 (N_2138,In_412,In_831);
nor U2139 (N_2139,In_682,In_773);
nand U2140 (N_2140,In_6,In_167);
nor U2141 (N_2141,In_621,In_820);
or U2142 (N_2142,In_584,In_641);
nor U2143 (N_2143,In_129,In_716);
or U2144 (N_2144,In_347,In_626);
nand U2145 (N_2145,In_544,In_300);
nand U2146 (N_2146,In_284,In_627);
or U2147 (N_2147,In_787,In_968);
or U2148 (N_2148,In_792,In_436);
nand U2149 (N_2149,In_908,In_114);
and U2150 (N_2150,In_319,In_612);
and U2151 (N_2151,In_474,In_482);
nor U2152 (N_2152,In_401,In_586);
nor U2153 (N_2153,In_911,In_14);
or U2154 (N_2154,In_900,In_204);
nand U2155 (N_2155,In_838,In_395);
nor U2156 (N_2156,In_478,In_299);
nor U2157 (N_2157,In_570,In_4);
and U2158 (N_2158,In_662,In_303);
or U2159 (N_2159,In_385,In_524);
xnor U2160 (N_2160,In_559,In_714);
or U2161 (N_2161,In_288,In_853);
or U2162 (N_2162,In_820,In_393);
nor U2163 (N_2163,In_619,In_421);
nand U2164 (N_2164,In_970,In_940);
or U2165 (N_2165,In_865,In_733);
nor U2166 (N_2166,In_638,In_640);
nor U2167 (N_2167,In_787,In_60);
nand U2168 (N_2168,In_615,In_174);
xor U2169 (N_2169,In_979,In_650);
or U2170 (N_2170,In_880,In_533);
and U2171 (N_2171,In_454,In_224);
or U2172 (N_2172,In_129,In_210);
or U2173 (N_2173,In_17,In_730);
nand U2174 (N_2174,In_677,In_279);
xor U2175 (N_2175,In_774,In_686);
nor U2176 (N_2176,In_594,In_490);
and U2177 (N_2177,In_540,In_47);
or U2178 (N_2178,In_136,In_137);
nand U2179 (N_2179,In_133,In_175);
and U2180 (N_2180,In_384,In_632);
or U2181 (N_2181,In_556,In_961);
nor U2182 (N_2182,In_430,In_213);
or U2183 (N_2183,In_73,In_512);
nand U2184 (N_2184,In_251,In_295);
nor U2185 (N_2185,In_19,In_59);
nor U2186 (N_2186,In_622,In_700);
or U2187 (N_2187,In_711,In_163);
xnor U2188 (N_2188,In_370,In_338);
and U2189 (N_2189,In_384,In_510);
or U2190 (N_2190,In_534,In_594);
or U2191 (N_2191,In_655,In_618);
and U2192 (N_2192,In_998,In_159);
or U2193 (N_2193,In_810,In_350);
nor U2194 (N_2194,In_549,In_220);
nand U2195 (N_2195,In_718,In_445);
or U2196 (N_2196,In_374,In_124);
nand U2197 (N_2197,In_512,In_179);
nor U2198 (N_2198,In_145,In_973);
nand U2199 (N_2199,In_274,In_927);
nand U2200 (N_2200,In_770,In_857);
nand U2201 (N_2201,In_824,In_577);
nor U2202 (N_2202,In_663,In_592);
nand U2203 (N_2203,In_15,In_445);
nand U2204 (N_2204,In_908,In_208);
xnor U2205 (N_2205,In_255,In_515);
nand U2206 (N_2206,In_618,In_905);
or U2207 (N_2207,In_9,In_575);
nor U2208 (N_2208,In_80,In_522);
or U2209 (N_2209,In_801,In_756);
nor U2210 (N_2210,In_714,In_625);
nand U2211 (N_2211,In_462,In_68);
nand U2212 (N_2212,In_757,In_607);
nand U2213 (N_2213,In_496,In_431);
nand U2214 (N_2214,In_263,In_276);
or U2215 (N_2215,In_379,In_594);
or U2216 (N_2216,In_900,In_220);
nand U2217 (N_2217,In_480,In_582);
nor U2218 (N_2218,In_177,In_77);
and U2219 (N_2219,In_541,In_805);
nand U2220 (N_2220,In_432,In_825);
nor U2221 (N_2221,In_795,In_95);
nor U2222 (N_2222,In_139,In_294);
and U2223 (N_2223,In_673,In_305);
nor U2224 (N_2224,In_688,In_826);
and U2225 (N_2225,In_197,In_727);
or U2226 (N_2226,In_770,In_333);
nand U2227 (N_2227,In_182,In_461);
or U2228 (N_2228,In_485,In_910);
or U2229 (N_2229,In_143,In_348);
nand U2230 (N_2230,In_575,In_744);
and U2231 (N_2231,In_900,In_155);
and U2232 (N_2232,In_743,In_817);
nand U2233 (N_2233,In_9,In_343);
xnor U2234 (N_2234,In_796,In_233);
nand U2235 (N_2235,In_567,In_19);
nand U2236 (N_2236,In_90,In_627);
or U2237 (N_2237,In_11,In_540);
xnor U2238 (N_2238,In_344,In_142);
nor U2239 (N_2239,In_269,In_334);
or U2240 (N_2240,In_104,In_749);
and U2241 (N_2241,In_956,In_84);
nor U2242 (N_2242,In_376,In_267);
nor U2243 (N_2243,In_876,In_791);
and U2244 (N_2244,In_48,In_630);
nor U2245 (N_2245,In_685,In_162);
and U2246 (N_2246,In_288,In_66);
nor U2247 (N_2247,In_721,In_658);
and U2248 (N_2248,In_39,In_666);
or U2249 (N_2249,In_673,In_246);
or U2250 (N_2250,In_515,In_396);
and U2251 (N_2251,In_247,In_287);
and U2252 (N_2252,In_420,In_751);
and U2253 (N_2253,In_168,In_511);
and U2254 (N_2254,In_986,In_431);
nand U2255 (N_2255,In_175,In_160);
nand U2256 (N_2256,In_901,In_157);
and U2257 (N_2257,In_479,In_861);
xor U2258 (N_2258,In_591,In_843);
or U2259 (N_2259,In_714,In_101);
xor U2260 (N_2260,In_462,In_364);
nand U2261 (N_2261,In_818,In_615);
or U2262 (N_2262,In_686,In_117);
and U2263 (N_2263,In_268,In_727);
and U2264 (N_2264,In_235,In_288);
nor U2265 (N_2265,In_194,In_709);
or U2266 (N_2266,In_48,In_817);
nand U2267 (N_2267,In_570,In_304);
nand U2268 (N_2268,In_850,In_243);
or U2269 (N_2269,In_537,In_826);
nor U2270 (N_2270,In_519,In_940);
nor U2271 (N_2271,In_923,In_874);
nor U2272 (N_2272,In_768,In_449);
or U2273 (N_2273,In_234,In_761);
or U2274 (N_2274,In_416,In_895);
and U2275 (N_2275,In_534,In_484);
nand U2276 (N_2276,In_450,In_154);
nor U2277 (N_2277,In_705,In_397);
nor U2278 (N_2278,In_330,In_875);
and U2279 (N_2279,In_482,In_803);
xor U2280 (N_2280,In_875,In_542);
and U2281 (N_2281,In_223,In_806);
nor U2282 (N_2282,In_457,In_935);
and U2283 (N_2283,In_981,In_71);
nor U2284 (N_2284,In_902,In_549);
and U2285 (N_2285,In_907,In_851);
nand U2286 (N_2286,In_590,In_384);
nor U2287 (N_2287,In_972,In_914);
nand U2288 (N_2288,In_16,In_382);
nor U2289 (N_2289,In_822,In_828);
nand U2290 (N_2290,In_693,In_105);
or U2291 (N_2291,In_89,In_136);
nand U2292 (N_2292,In_32,In_108);
and U2293 (N_2293,In_180,In_777);
nand U2294 (N_2294,In_992,In_810);
or U2295 (N_2295,In_481,In_561);
nand U2296 (N_2296,In_352,In_692);
nor U2297 (N_2297,In_143,In_858);
or U2298 (N_2298,In_852,In_361);
and U2299 (N_2299,In_206,In_251);
and U2300 (N_2300,In_806,In_427);
nor U2301 (N_2301,In_684,In_559);
and U2302 (N_2302,In_721,In_907);
nor U2303 (N_2303,In_591,In_707);
nand U2304 (N_2304,In_185,In_904);
nor U2305 (N_2305,In_372,In_251);
nand U2306 (N_2306,In_525,In_851);
nand U2307 (N_2307,In_27,In_46);
nand U2308 (N_2308,In_617,In_460);
nor U2309 (N_2309,In_719,In_503);
nand U2310 (N_2310,In_919,In_692);
nor U2311 (N_2311,In_289,In_859);
xnor U2312 (N_2312,In_868,In_700);
nand U2313 (N_2313,In_684,In_528);
nor U2314 (N_2314,In_911,In_741);
or U2315 (N_2315,In_357,In_780);
nand U2316 (N_2316,In_18,In_890);
and U2317 (N_2317,In_776,In_829);
nand U2318 (N_2318,In_876,In_750);
nand U2319 (N_2319,In_772,In_304);
nor U2320 (N_2320,In_252,In_194);
and U2321 (N_2321,In_486,In_656);
nand U2322 (N_2322,In_210,In_606);
nor U2323 (N_2323,In_110,In_444);
nand U2324 (N_2324,In_236,In_996);
nor U2325 (N_2325,In_415,In_935);
and U2326 (N_2326,In_160,In_930);
nand U2327 (N_2327,In_576,In_772);
and U2328 (N_2328,In_353,In_396);
nor U2329 (N_2329,In_307,In_246);
and U2330 (N_2330,In_663,In_564);
nor U2331 (N_2331,In_76,In_855);
nor U2332 (N_2332,In_969,In_122);
nand U2333 (N_2333,In_180,In_154);
nand U2334 (N_2334,In_550,In_313);
nor U2335 (N_2335,In_785,In_465);
and U2336 (N_2336,In_186,In_978);
or U2337 (N_2337,In_939,In_117);
nand U2338 (N_2338,In_117,In_97);
nor U2339 (N_2339,In_83,In_697);
nand U2340 (N_2340,In_343,In_625);
or U2341 (N_2341,In_263,In_444);
nor U2342 (N_2342,In_157,In_636);
and U2343 (N_2343,In_644,In_115);
and U2344 (N_2344,In_216,In_987);
nor U2345 (N_2345,In_923,In_54);
and U2346 (N_2346,In_73,In_522);
nand U2347 (N_2347,In_108,In_472);
nor U2348 (N_2348,In_318,In_562);
or U2349 (N_2349,In_27,In_21);
nand U2350 (N_2350,In_591,In_595);
or U2351 (N_2351,In_724,In_932);
or U2352 (N_2352,In_690,In_240);
nand U2353 (N_2353,In_339,In_564);
nor U2354 (N_2354,In_679,In_214);
nor U2355 (N_2355,In_70,In_846);
or U2356 (N_2356,In_785,In_603);
nand U2357 (N_2357,In_510,In_193);
and U2358 (N_2358,In_712,In_787);
nor U2359 (N_2359,In_299,In_812);
xnor U2360 (N_2360,In_782,In_565);
xor U2361 (N_2361,In_480,In_45);
xor U2362 (N_2362,In_393,In_521);
xor U2363 (N_2363,In_781,In_854);
or U2364 (N_2364,In_68,In_262);
nor U2365 (N_2365,In_275,In_452);
nor U2366 (N_2366,In_536,In_384);
nand U2367 (N_2367,In_958,In_39);
or U2368 (N_2368,In_499,In_938);
nor U2369 (N_2369,In_320,In_624);
or U2370 (N_2370,In_898,In_190);
and U2371 (N_2371,In_118,In_715);
nand U2372 (N_2372,In_395,In_929);
or U2373 (N_2373,In_570,In_909);
xor U2374 (N_2374,In_861,In_631);
or U2375 (N_2375,In_964,In_140);
or U2376 (N_2376,In_598,In_824);
or U2377 (N_2377,In_164,In_611);
nor U2378 (N_2378,In_649,In_923);
and U2379 (N_2379,In_239,In_52);
nor U2380 (N_2380,In_968,In_776);
nand U2381 (N_2381,In_513,In_701);
nor U2382 (N_2382,In_852,In_218);
nand U2383 (N_2383,In_792,In_977);
or U2384 (N_2384,In_192,In_521);
nor U2385 (N_2385,In_111,In_643);
and U2386 (N_2386,In_244,In_975);
nand U2387 (N_2387,In_278,In_6);
and U2388 (N_2388,In_415,In_152);
or U2389 (N_2389,In_781,In_484);
nand U2390 (N_2390,In_180,In_699);
nor U2391 (N_2391,In_850,In_820);
nand U2392 (N_2392,In_110,In_174);
and U2393 (N_2393,In_987,In_266);
and U2394 (N_2394,In_467,In_389);
nor U2395 (N_2395,In_803,In_689);
xor U2396 (N_2396,In_897,In_191);
or U2397 (N_2397,In_493,In_93);
nand U2398 (N_2398,In_465,In_382);
and U2399 (N_2399,In_514,In_777);
or U2400 (N_2400,In_587,In_522);
and U2401 (N_2401,In_79,In_258);
nor U2402 (N_2402,In_731,In_416);
nand U2403 (N_2403,In_8,In_94);
nor U2404 (N_2404,In_562,In_857);
or U2405 (N_2405,In_21,In_59);
nor U2406 (N_2406,In_843,In_547);
or U2407 (N_2407,In_901,In_426);
nand U2408 (N_2408,In_175,In_371);
nor U2409 (N_2409,In_883,In_496);
nor U2410 (N_2410,In_297,In_227);
or U2411 (N_2411,In_712,In_913);
xor U2412 (N_2412,In_334,In_910);
and U2413 (N_2413,In_250,In_635);
nor U2414 (N_2414,In_951,In_647);
nand U2415 (N_2415,In_546,In_708);
and U2416 (N_2416,In_152,In_914);
nor U2417 (N_2417,In_245,In_16);
or U2418 (N_2418,In_10,In_513);
nor U2419 (N_2419,In_582,In_386);
xnor U2420 (N_2420,In_427,In_197);
and U2421 (N_2421,In_433,In_387);
and U2422 (N_2422,In_452,In_926);
or U2423 (N_2423,In_84,In_51);
xor U2424 (N_2424,In_300,In_709);
nor U2425 (N_2425,In_933,In_329);
nand U2426 (N_2426,In_669,In_516);
nand U2427 (N_2427,In_679,In_776);
and U2428 (N_2428,In_224,In_680);
nand U2429 (N_2429,In_327,In_699);
nor U2430 (N_2430,In_337,In_648);
or U2431 (N_2431,In_860,In_453);
and U2432 (N_2432,In_17,In_27);
or U2433 (N_2433,In_507,In_431);
and U2434 (N_2434,In_187,In_991);
nand U2435 (N_2435,In_36,In_466);
or U2436 (N_2436,In_935,In_920);
and U2437 (N_2437,In_679,In_273);
nor U2438 (N_2438,In_186,In_747);
nand U2439 (N_2439,In_486,In_573);
or U2440 (N_2440,In_963,In_85);
xnor U2441 (N_2441,In_347,In_736);
or U2442 (N_2442,In_766,In_149);
xor U2443 (N_2443,In_916,In_123);
or U2444 (N_2444,In_601,In_630);
or U2445 (N_2445,In_581,In_257);
nor U2446 (N_2446,In_957,In_962);
nand U2447 (N_2447,In_648,In_692);
and U2448 (N_2448,In_347,In_906);
and U2449 (N_2449,In_178,In_458);
and U2450 (N_2450,In_548,In_484);
nand U2451 (N_2451,In_16,In_236);
or U2452 (N_2452,In_805,In_745);
xor U2453 (N_2453,In_760,In_790);
and U2454 (N_2454,In_230,In_667);
nor U2455 (N_2455,In_772,In_482);
xnor U2456 (N_2456,In_894,In_831);
or U2457 (N_2457,In_854,In_772);
nor U2458 (N_2458,In_267,In_406);
and U2459 (N_2459,In_912,In_984);
nand U2460 (N_2460,In_154,In_177);
and U2461 (N_2461,In_33,In_331);
and U2462 (N_2462,In_236,In_436);
nor U2463 (N_2463,In_279,In_585);
and U2464 (N_2464,In_789,In_704);
nand U2465 (N_2465,In_226,In_969);
and U2466 (N_2466,In_404,In_285);
nor U2467 (N_2467,In_292,In_402);
nand U2468 (N_2468,In_676,In_565);
xnor U2469 (N_2469,In_89,In_581);
or U2470 (N_2470,In_315,In_1);
or U2471 (N_2471,In_520,In_86);
and U2472 (N_2472,In_705,In_435);
or U2473 (N_2473,In_898,In_750);
or U2474 (N_2474,In_979,In_897);
nor U2475 (N_2475,In_984,In_575);
nor U2476 (N_2476,In_932,In_268);
nand U2477 (N_2477,In_739,In_368);
nand U2478 (N_2478,In_483,In_479);
nand U2479 (N_2479,In_266,In_36);
and U2480 (N_2480,In_13,In_93);
and U2481 (N_2481,In_859,In_529);
nor U2482 (N_2482,In_244,In_108);
nor U2483 (N_2483,In_751,In_472);
nor U2484 (N_2484,In_812,In_981);
and U2485 (N_2485,In_100,In_928);
and U2486 (N_2486,In_127,In_163);
and U2487 (N_2487,In_100,In_235);
xor U2488 (N_2488,In_403,In_583);
or U2489 (N_2489,In_764,In_530);
nand U2490 (N_2490,In_779,In_358);
nor U2491 (N_2491,In_532,In_110);
nor U2492 (N_2492,In_491,In_893);
or U2493 (N_2493,In_837,In_645);
nand U2494 (N_2494,In_287,In_24);
and U2495 (N_2495,In_138,In_711);
and U2496 (N_2496,In_832,In_745);
nand U2497 (N_2497,In_252,In_366);
or U2498 (N_2498,In_625,In_766);
nor U2499 (N_2499,In_703,In_199);
nor U2500 (N_2500,In_374,In_830);
and U2501 (N_2501,In_343,In_879);
xor U2502 (N_2502,In_101,In_536);
or U2503 (N_2503,In_621,In_55);
or U2504 (N_2504,In_497,In_340);
and U2505 (N_2505,In_617,In_693);
nand U2506 (N_2506,In_276,In_675);
or U2507 (N_2507,In_396,In_3);
or U2508 (N_2508,In_876,In_289);
xnor U2509 (N_2509,In_18,In_953);
and U2510 (N_2510,In_422,In_145);
nand U2511 (N_2511,In_270,In_572);
and U2512 (N_2512,In_97,In_599);
or U2513 (N_2513,In_927,In_809);
nand U2514 (N_2514,In_45,In_414);
or U2515 (N_2515,In_70,In_403);
or U2516 (N_2516,In_922,In_531);
nand U2517 (N_2517,In_33,In_547);
or U2518 (N_2518,In_501,In_489);
or U2519 (N_2519,In_88,In_609);
nand U2520 (N_2520,In_999,In_765);
nor U2521 (N_2521,In_131,In_105);
nor U2522 (N_2522,In_113,In_572);
nand U2523 (N_2523,In_382,In_231);
nand U2524 (N_2524,In_489,In_760);
nor U2525 (N_2525,In_747,In_392);
and U2526 (N_2526,In_47,In_763);
or U2527 (N_2527,In_888,In_546);
nor U2528 (N_2528,In_428,In_383);
nand U2529 (N_2529,In_826,In_338);
nor U2530 (N_2530,In_437,In_301);
nand U2531 (N_2531,In_528,In_370);
or U2532 (N_2532,In_428,In_280);
and U2533 (N_2533,In_707,In_42);
or U2534 (N_2534,In_757,In_886);
or U2535 (N_2535,In_355,In_716);
nor U2536 (N_2536,In_270,In_529);
or U2537 (N_2537,In_808,In_389);
and U2538 (N_2538,In_831,In_891);
and U2539 (N_2539,In_817,In_647);
and U2540 (N_2540,In_984,In_957);
or U2541 (N_2541,In_841,In_877);
or U2542 (N_2542,In_804,In_336);
nor U2543 (N_2543,In_591,In_563);
nor U2544 (N_2544,In_113,In_465);
nand U2545 (N_2545,In_566,In_992);
and U2546 (N_2546,In_750,In_440);
and U2547 (N_2547,In_245,In_190);
nor U2548 (N_2548,In_710,In_472);
and U2549 (N_2549,In_147,In_127);
and U2550 (N_2550,In_954,In_333);
or U2551 (N_2551,In_963,In_943);
nand U2552 (N_2552,In_552,In_404);
nand U2553 (N_2553,In_858,In_172);
and U2554 (N_2554,In_499,In_101);
nor U2555 (N_2555,In_778,In_645);
nor U2556 (N_2556,In_605,In_831);
nor U2557 (N_2557,In_34,In_17);
nand U2558 (N_2558,In_251,In_916);
and U2559 (N_2559,In_601,In_808);
or U2560 (N_2560,In_994,In_417);
or U2561 (N_2561,In_249,In_488);
nand U2562 (N_2562,In_492,In_664);
nor U2563 (N_2563,In_991,In_929);
nand U2564 (N_2564,In_56,In_463);
and U2565 (N_2565,In_215,In_419);
nor U2566 (N_2566,In_166,In_946);
or U2567 (N_2567,In_738,In_131);
or U2568 (N_2568,In_11,In_904);
or U2569 (N_2569,In_5,In_249);
and U2570 (N_2570,In_143,In_465);
nor U2571 (N_2571,In_799,In_412);
nand U2572 (N_2572,In_762,In_299);
nand U2573 (N_2573,In_733,In_957);
nand U2574 (N_2574,In_921,In_76);
nor U2575 (N_2575,In_192,In_524);
or U2576 (N_2576,In_482,In_989);
or U2577 (N_2577,In_1,In_413);
nand U2578 (N_2578,In_62,In_106);
nor U2579 (N_2579,In_624,In_470);
nand U2580 (N_2580,In_289,In_95);
nor U2581 (N_2581,In_526,In_856);
nor U2582 (N_2582,In_917,In_805);
and U2583 (N_2583,In_534,In_955);
and U2584 (N_2584,In_126,In_597);
nand U2585 (N_2585,In_188,In_512);
nor U2586 (N_2586,In_328,In_229);
or U2587 (N_2587,In_951,In_507);
nand U2588 (N_2588,In_524,In_882);
and U2589 (N_2589,In_187,In_567);
nor U2590 (N_2590,In_847,In_845);
and U2591 (N_2591,In_424,In_263);
nor U2592 (N_2592,In_812,In_452);
and U2593 (N_2593,In_987,In_48);
nand U2594 (N_2594,In_40,In_925);
nand U2595 (N_2595,In_387,In_839);
nand U2596 (N_2596,In_89,In_204);
and U2597 (N_2597,In_887,In_902);
nand U2598 (N_2598,In_689,In_275);
or U2599 (N_2599,In_214,In_280);
xor U2600 (N_2600,In_683,In_627);
nand U2601 (N_2601,In_702,In_738);
xor U2602 (N_2602,In_112,In_265);
nand U2603 (N_2603,In_70,In_238);
nand U2604 (N_2604,In_136,In_645);
xor U2605 (N_2605,In_414,In_665);
nand U2606 (N_2606,In_238,In_307);
and U2607 (N_2607,In_163,In_619);
and U2608 (N_2608,In_820,In_473);
and U2609 (N_2609,In_910,In_994);
nand U2610 (N_2610,In_803,In_871);
xnor U2611 (N_2611,In_23,In_833);
nand U2612 (N_2612,In_718,In_100);
nor U2613 (N_2613,In_264,In_760);
nand U2614 (N_2614,In_638,In_268);
nand U2615 (N_2615,In_792,In_734);
and U2616 (N_2616,In_772,In_328);
nor U2617 (N_2617,In_949,In_87);
or U2618 (N_2618,In_893,In_76);
and U2619 (N_2619,In_240,In_631);
xnor U2620 (N_2620,In_868,In_559);
and U2621 (N_2621,In_325,In_423);
nor U2622 (N_2622,In_80,In_567);
nand U2623 (N_2623,In_477,In_543);
and U2624 (N_2624,In_905,In_230);
and U2625 (N_2625,In_58,In_281);
and U2626 (N_2626,In_522,In_674);
xor U2627 (N_2627,In_125,In_611);
and U2628 (N_2628,In_430,In_613);
and U2629 (N_2629,In_584,In_4);
nand U2630 (N_2630,In_628,In_65);
and U2631 (N_2631,In_284,In_396);
or U2632 (N_2632,In_478,In_165);
and U2633 (N_2633,In_971,In_394);
and U2634 (N_2634,In_486,In_719);
xor U2635 (N_2635,In_580,In_907);
xor U2636 (N_2636,In_138,In_679);
nor U2637 (N_2637,In_888,In_383);
nor U2638 (N_2638,In_945,In_731);
nor U2639 (N_2639,In_754,In_894);
nor U2640 (N_2640,In_261,In_705);
or U2641 (N_2641,In_167,In_103);
nor U2642 (N_2642,In_726,In_466);
nor U2643 (N_2643,In_68,In_790);
or U2644 (N_2644,In_608,In_267);
nand U2645 (N_2645,In_660,In_550);
xnor U2646 (N_2646,In_818,In_269);
or U2647 (N_2647,In_527,In_471);
or U2648 (N_2648,In_25,In_933);
or U2649 (N_2649,In_843,In_759);
xor U2650 (N_2650,In_583,In_683);
nand U2651 (N_2651,In_562,In_85);
and U2652 (N_2652,In_956,In_445);
and U2653 (N_2653,In_98,In_866);
nor U2654 (N_2654,In_121,In_804);
and U2655 (N_2655,In_490,In_589);
and U2656 (N_2656,In_864,In_486);
or U2657 (N_2657,In_304,In_388);
or U2658 (N_2658,In_929,In_496);
and U2659 (N_2659,In_257,In_326);
and U2660 (N_2660,In_542,In_677);
nand U2661 (N_2661,In_120,In_29);
and U2662 (N_2662,In_546,In_140);
xnor U2663 (N_2663,In_692,In_213);
xnor U2664 (N_2664,In_212,In_476);
or U2665 (N_2665,In_340,In_399);
and U2666 (N_2666,In_707,In_200);
nand U2667 (N_2667,In_54,In_979);
nand U2668 (N_2668,In_294,In_365);
and U2669 (N_2669,In_87,In_585);
and U2670 (N_2670,In_27,In_145);
nand U2671 (N_2671,In_865,In_41);
nand U2672 (N_2672,In_376,In_52);
xnor U2673 (N_2673,In_334,In_847);
and U2674 (N_2674,In_452,In_454);
and U2675 (N_2675,In_258,In_555);
nor U2676 (N_2676,In_160,In_51);
nor U2677 (N_2677,In_231,In_987);
and U2678 (N_2678,In_208,In_405);
and U2679 (N_2679,In_794,In_497);
and U2680 (N_2680,In_905,In_604);
nor U2681 (N_2681,In_257,In_453);
or U2682 (N_2682,In_478,In_235);
nand U2683 (N_2683,In_945,In_244);
and U2684 (N_2684,In_72,In_994);
or U2685 (N_2685,In_663,In_452);
nor U2686 (N_2686,In_266,In_391);
nand U2687 (N_2687,In_161,In_301);
or U2688 (N_2688,In_71,In_171);
nand U2689 (N_2689,In_88,In_518);
nor U2690 (N_2690,In_63,In_487);
nand U2691 (N_2691,In_368,In_41);
nand U2692 (N_2692,In_16,In_856);
nand U2693 (N_2693,In_797,In_235);
nand U2694 (N_2694,In_595,In_647);
xnor U2695 (N_2695,In_848,In_766);
and U2696 (N_2696,In_521,In_870);
or U2697 (N_2697,In_587,In_819);
and U2698 (N_2698,In_531,In_140);
nand U2699 (N_2699,In_805,In_107);
nor U2700 (N_2700,In_483,In_33);
nand U2701 (N_2701,In_478,In_906);
nor U2702 (N_2702,In_863,In_469);
or U2703 (N_2703,In_144,In_131);
and U2704 (N_2704,In_811,In_136);
nor U2705 (N_2705,In_998,In_747);
or U2706 (N_2706,In_443,In_115);
or U2707 (N_2707,In_852,In_302);
and U2708 (N_2708,In_528,In_284);
nand U2709 (N_2709,In_988,In_481);
xnor U2710 (N_2710,In_150,In_164);
nor U2711 (N_2711,In_856,In_862);
or U2712 (N_2712,In_930,In_563);
nand U2713 (N_2713,In_750,In_260);
and U2714 (N_2714,In_972,In_368);
nand U2715 (N_2715,In_54,In_238);
or U2716 (N_2716,In_590,In_679);
nor U2717 (N_2717,In_151,In_115);
nor U2718 (N_2718,In_46,In_833);
and U2719 (N_2719,In_539,In_425);
nand U2720 (N_2720,In_923,In_238);
and U2721 (N_2721,In_463,In_68);
nand U2722 (N_2722,In_964,In_314);
nor U2723 (N_2723,In_923,In_125);
nor U2724 (N_2724,In_410,In_512);
nand U2725 (N_2725,In_478,In_714);
nand U2726 (N_2726,In_208,In_256);
and U2727 (N_2727,In_32,In_501);
nor U2728 (N_2728,In_892,In_910);
and U2729 (N_2729,In_338,In_69);
nor U2730 (N_2730,In_161,In_106);
and U2731 (N_2731,In_11,In_441);
nor U2732 (N_2732,In_281,In_946);
and U2733 (N_2733,In_177,In_320);
nand U2734 (N_2734,In_351,In_695);
or U2735 (N_2735,In_822,In_329);
and U2736 (N_2736,In_863,In_923);
and U2737 (N_2737,In_602,In_68);
and U2738 (N_2738,In_333,In_231);
nand U2739 (N_2739,In_733,In_168);
nor U2740 (N_2740,In_472,In_479);
nand U2741 (N_2741,In_975,In_596);
xnor U2742 (N_2742,In_120,In_842);
or U2743 (N_2743,In_108,In_48);
or U2744 (N_2744,In_874,In_832);
nor U2745 (N_2745,In_892,In_369);
nor U2746 (N_2746,In_888,In_492);
nand U2747 (N_2747,In_801,In_862);
and U2748 (N_2748,In_784,In_41);
nand U2749 (N_2749,In_540,In_469);
or U2750 (N_2750,In_877,In_514);
or U2751 (N_2751,In_79,In_393);
nor U2752 (N_2752,In_89,In_981);
and U2753 (N_2753,In_262,In_273);
nand U2754 (N_2754,In_253,In_474);
nor U2755 (N_2755,In_417,In_248);
nand U2756 (N_2756,In_812,In_412);
or U2757 (N_2757,In_287,In_203);
nand U2758 (N_2758,In_623,In_658);
xnor U2759 (N_2759,In_140,In_781);
or U2760 (N_2760,In_414,In_553);
or U2761 (N_2761,In_252,In_352);
xnor U2762 (N_2762,In_300,In_144);
nor U2763 (N_2763,In_268,In_412);
or U2764 (N_2764,In_447,In_743);
nor U2765 (N_2765,In_974,In_8);
nand U2766 (N_2766,In_625,In_525);
and U2767 (N_2767,In_576,In_5);
xor U2768 (N_2768,In_647,In_352);
nor U2769 (N_2769,In_297,In_652);
or U2770 (N_2770,In_735,In_369);
nor U2771 (N_2771,In_320,In_534);
nand U2772 (N_2772,In_23,In_60);
nor U2773 (N_2773,In_176,In_280);
xor U2774 (N_2774,In_960,In_342);
nor U2775 (N_2775,In_816,In_875);
nor U2776 (N_2776,In_479,In_934);
and U2777 (N_2777,In_356,In_845);
nand U2778 (N_2778,In_421,In_486);
nand U2779 (N_2779,In_226,In_268);
nand U2780 (N_2780,In_32,In_905);
xnor U2781 (N_2781,In_968,In_67);
nand U2782 (N_2782,In_200,In_346);
xor U2783 (N_2783,In_811,In_191);
or U2784 (N_2784,In_385,In_933);
nor U2785 (N_2785,In_424,In_371);
nand U2786 (N_2786,In_485,In_825);
nand U2787 (N_2787,In_971,In_431);
or U2788 (N_2788,In_542,In_653);
or U2789 (N_2789,In_437,In_781);
and U2790 (N_2790,In_38,In_601);
nand U2791 (N_2791,In_756,In_347);
xnor U2792 (N_2792,In_15,In_927);
nor U2793 (N_2793,In_337,In_977);
or U2794 (N_2794,In_601,In_330);
xor U2795 (N_2795,In_394,In_554);
xor U2796 (N_2796,In_122,In_623);
or U2797 (N_2797,In_217,In_29);
nor U2798 (N_2798,In_746,In_587);
nor U2799 (N_2799,In_85,In_463);
nand U2800 (N_2800,In_835,In_615);
nor U2801 (N_2801,In_140,In_911);
nand U2802 (N_2802,In_981,In_495);
and U2803 (N_2803,In_940,In_431);
nand U2804 (N_2804,In_594,In_756);
or U2805 (N_2805,In_699,In_557);
nor U2806 (N_2806,In_325,In_18);
nor U2807 (N_2807,In_767,In_892);
nor U2808 (N_2808,In_912,In_398);
and U2809 (N_2809,In_124,In_308);
xor U2810 (N_2810,In_93,In_516);
nand U2811 (N_2811,In_309,In_3);
and U2812 (N_2812,In_744,In_292);
and U2813 (N_2813,In_796,In_487);
nand U2814 (N_2814,In_223,In_743);
and U2815 (N_2815,In_104,In_743);
nor U2816 (N_2816,In_458,In_455);
nor U2817 (N_2817,In_671,In_770);
and U2818 (N_2818,In_24,In_141);
or U2819 (N_2819,In_858,In_742);
nand U2820 (N_2820,In_370,In_476);
or U2821 (N_2821,In_802,In_336);
nand U2822 (N_2822,In_710,In_775);
and U2823 (N_2823,In_796,In_535);
nor U2824 (N_2824,In_999,In_909);
nor U2825 (N_2825,In_25,In_883);
or U2826 (N_2826,In_903,In_735);
nor U2827 (N_2827,In_498,In_189);
or U2828 (N_2828,In_119,In_930);
or U2829 (N_2829,In_852,In_317);
xor U2830 (N_2830,In_68,In_272);
or U2831 (N_2831,In_862,In_436);
or U2832 (N_2832,In_532,In_217);
nand U2833 (N_2833,In_929,In_192);
nand U2834 (N_2834,In_610,In_131);
and U2835 (N_2835,In_755,In_270);
xnor U2836 (N_2836,In_403,In_593);
or U2837 (N_2837,In_148,In_368);
xor U2838 (N_2838,In_165,In_857);
or U2839 (N_2839,In_357,In_875);
or U2840 (N_2840,In_32,In_636);
nand U2841 (N_2841,In_89,In_621);
nand U2842 (N_2842,In_392,In_465);
or U2843 (N_2843,In_21,In_391);
or U2844 (N_2844,In_661,In_26);
or U2845 (N_2845,In_192,In_790);
or U2846 (N_2846,In_208,In_226);
or U2847 (N_2847,In_484,In_480);
nand U2848 (N_2848,In_29,In_795);
and U2849 (N_2849,In_192,In_438);
nand U2850 (N_2850,In_363,In_958);
xor U2851 (N_2851,In_471,In_65);
or U2852 (N_2852,In_506,In_663);
nor U2853 (N_2853,In_512,In_34);
and U2854 (N_2854,In_246,In_213);
or U2855 (N_2855,In_347,In_684);
or U2856 (N_2856,In_640,In_559);
or U2857 (N_2857,In_80,In_9);
or U2858 (N_2858,In_887,In_213);
nand U2859 (N_2859,In_876,In_486);
nor U2860 (N_2860,In_526,In_337);
nor U2861 (N_2861,In_221,In_487);
or U2862 (N_2862,In_97,In_331);
nand U2863 (N_2863,In_398,In_387);
nor U2864 (N_2864,In_297,In_57);
and U2865 (N_2865,In_82,In_738);
or U2866 (N_2866,In_265,In_200);
xnor U2867 (N_2867,In_509,In_230);
nand U2868 (N_2868,In_429,In_189);
and U2869 (N_2869,In_362,In_556);
and U2870 (N_2870,In_847,In_460);
or U2871 (N_2871,In_838,In_653);
xnor U2872 (N_2872,In_37,In_845);
xor U2873 (N_2873,In_97,In_467);
nand U2874 (N_2874,In_256,In_982);
nand U2875 (N_2875,In_874,In_486);
or U2876 (N_2876,In_475,In_936);
or U2877 (N_2877,In_384,In_628);
or U2878 (N_2878,In_951,In_441);
xor U2879 (N_2879,In_939,In_827);
nor U2880 (N_2880,In_561,In_194);
nand U2881 (N_2881,In_840,In_474);
nand U2882 (N_2882,In_968,In_844);
xnor U2883 (N_2883,In_188,In_836);
nand U2884 (N_2884,In_313,In_732);
or U2885 (N_2885,In_167,In_172);
and U2886 (N_2886,In_628,In_924);
and U2887 (N_2887,In_460,In_615);
nor U2888 (N_2888,In_171,In_546);
and U2889 (N_2889,In_742,In_321);
xor U2890 (N_2890,In_170,In_220);
nand U2891 (N_2891,In_604,In_710);
nor U2892 (N_2892,In_395,In_542);
or U2893 (N_2893,In_703,In_94);
nor U2894 (N_2894,In_198,In_796);
nor U2895 (N_2895,In_463,In_957);
or U2896 (N_2896,In_423,In_507);
xor U2897 (N_2897,In_466,In_821);
nand U2898 (N_2898,In_503,In_909);
and U2899 (N_2899,In_521,In_314);
nand U2900 (N_2900,In_248,In_587);
and U2901 (N_2901,In_940,In_407);
nor U2902 (N_2902,In_634,In_926);
nand U2903 (N_2903,In_958,In_488);
or U2904 (N_2904,In_444,In_525);
xnor U2905 (N_2905,In_530,In_936);
nand U2906 (N_2906,In_610,In_57);
nand U2907 (N_2907,In_412,In_177);
nand U2908 (N_2908,In_465,In_358);
and U2909 (N_2909,In_962,In_251);
or U2910 (N_2910,In_278,In_986);
xnor U2911 (N_2911,In_855,In_360);
or U2912 (N_2912,In_412,In_427);
nor U2913 (N_2913,In_205,In_604);
nor U2914 (N_2914,In_933,In_45);
and U2915 (N_2915,In_403,In_466);
or U2916 (N_2916,In_496,In_72);
nand U2917 (N_2917,In_865,In_915);
or U2918 (N_2918,In_521,In_539);
and U2919 (N_2919,In_739,In_651);
xnor U2920 (N_2920,In_984,In_169);
nor U2921 (N_2921,In_630,In_542);
or U2922 (N_2922,In_71,In_773);
xor U2923 (N_2923,In_24,In_458);
xor U2924 (N_2924,In_355,In_583);
xnor U2925 (N_2925,In_289,In_584);
or U2926 (N_2926,In_684,In_735);
or U2927 (N_2927,In_430,In_276);
and U2928 (N_2928,In_861,In_49);
and U2929 (N_2929,In_455,In_999);
nor U2930 (N_2930,In_41,In_693);
nand U2931 (N_2931,In_477,In_547);
nor U2932 (N_2932,In_737,In_363);
or U2933 (N_2933,In_120,In_257);
nand U2934 (N_2934,In_481,In_857);
xor U2935 (N_2935,In_715,In_531);
nand U2936 (N_2936,In_497,In_145);
nand U2937 (N_2937,In_698,In_697);
nand U2938 (N_2938,In_488,In_675);
and U2939 (N_2939,In_255,In_872);
nand U2940 (N_2940,In_752,In_354);
nand U2941 (N_2941,In_623,In_997);
and U2942 (N_2942,In_436,In_79);
nand U2943 (N_2943,In_839,In_492);
and U2944 (N_2944,In_126,In_673);
nor U2945 (N_2945,In_188,In_102);
nor U2946 (N_2946,In_56,In_464);
or U2947 (N_2947,In_912,In_276);
or U2948 (N_2948,In_549,In_501);
and U2949 (N_2949,In_316,In_147);
nand U2950 (N_2950,In_28,In_229);
nand U2951 (N_2951,In_544,In_260);
nor U2952 (N_2952,In_538,In_250);
xor U2953 (N_2953,In_811,In_296);
xnor U2954 (N_2954,In_318,In_459);
or U2955 (N_2955,In_32,In_930);
and U2956 (N_2956,In_981,In_677);
or U2957 (N_2957,In_960,In_630);
nor U2958 (N_2958,In_297,In_786);
nor U2959 (N_2959,In_611,In_606);
nand U2960 (N_2960,In_331,In_732);
nor U2961 (N_2961,In_125,In_146);
nor U2962 (N_2962,In_917,In_980);
nand U2963 (N_2963,In_954,In_282);
or U2964 (N_2964,In_741,In_597);
and U2965 (N_2965,In_364,In_782);
nor U2966 (N_2966,In_227,In_114);
nor U2967 (N_2967,In_722,In_916);
or U2968 (N_2968,In_607,In_585);
nor U2969 (N_2969,In_22,In_608);
or U2970 (N_2970,In_393,In_486);
xor U2971 (N_2971,In_341,In_52);
or U2972 (N_2972,In_532,In_612);
nand U2973 (N_2973,In_390,In_426);
nor U2974 (N_2974,In_145,In_184);
nand U2975 (N_2975,In_674,In_681);
nor U2976 (N_2976,In_685,In_18);
or U2977 (N_2977,In_434,In_162);
nor U2978 (N_2978,In_777,In_45);
nand U2979 (N_2979,In_59,In_30);
nor U2980 (N_2980,In_636,In_51);
or U2981 (N_2981,In_557,In_143);
or U2982 (N_2982,In_687,In_830);
nand U2983 (N_2983,In_238,In_503);
nor U2984 (N_2984,In_431,In_500);
nor U2985 (N_2985,In_767,In_954);
nor U2986 (N_2986,In_656,In_187);
or U2987 (N_2987,In_671,In_306);
xnor U2988 (N_2988,In_356,In_542);
and U2989 (N_2989,In_927,In_251);
or U2990 (N_2990,In_779,In_573);
nor U2991 (N_2991,In_105,In_950);
nand U2992 (N_2992,In_413,In_646);
and U2993 (N_2993,In_247,In_965);
or U2994 (N_2994,In_941,In_678);
nand U2995 (N_2995,In_108,In_654);
and U2996 (N_2996,In_592,In_845);
and U2997 (N_2997,In_553,In_837);
nand U2998 (N_2998,In_245,In_111);
and U2999 (N_2999,In_824,In_115);
nand U3000 (N_3000,In_806,In_384);
nor U3001 (N_3001,In_713,In_516);
nor U3002 (N_3002,In_431,In_307);
nor U3003 (N_3003,In_58,In_226);
nand U3004 (N_3004,In_525,In_360);
nand U3005 (N_3005,In_187,In_735);
xor U3006 (N_3006,In_954,In_494);
and U3007 (N_3007,In_5,In_250);
nor U3008 (N_3008,In_583,In_632);
xor U3009 (N_3009,In_766,In_515);
nor U3010 (N_3010,In_602,In_43);
xor U3011 (N_3011,In_864,In_431);
nor U3012 (N_3012,In_109,In_927);
xor U3013 (N_3013,In_323,In_642);
and U3014 (N_3014,In_742,In_11);
and U3015 (N_3015,In_40,In_356);
nor U3016 (N_3016,In_992,In_951);
or U3017 (N_3017,In_841,In_811);
nand U3018 (N_3018,In_562,In_435);
and U3019 (N_3019,In_243,In_659);
nor U3020 (N_3020,In_341,In_817);
xnor U3021 (N_3021,In_297,In_941);
and U3022 (N_3022,In_361,In_295);
nor U3023 (N_3023,In_714,In_914);
or U3024 (N_3024,In_197,In_544);
nor U3025 (N_3025,In_14,In_450);
or U3026 (N_3026,In_986,In_873);
and U3027 (N_3027,In_142,In_977);
nor U3028 (N_3028,In_671,In_891);
and U3029 (N_3029,In_852,In_972);
or U3030 (N_3030,In_939,In_383);
nor U3031 (N_3031,In_781,In_807);
nand U3032 (N_3032,In_406,In_924);
or U3033 (N_3033,In_67,In_645);
and U3034 (N_3034,In_756,In_246);
nor U3035 (N_3035,In_238,In_254);
nand U3036 (N_3036,In_793,In_77);
nand U3037 (N_3037,In_900,In_990);
nand U3038 (N_3038,In_261,In_643);
or U3039 (N_3039,In_880,In_999);
and U3040 (N_3040,In_517,In_155);
and U3041 (N_3041,In_476,In_999);
and U3042 (N_3042,In_518,In_755);
nor U3043 (N_3043,In_210,In_839);
or U3044 (N_3044,In_959,In_145);
nor U3045 (N_3045,In_585,In_309);
and U3046 (N_3046,In_434,In_73);
xor U3047 (N_3047,In_792,In_252);
or U3048 (N_3048,In_866,In_860);
nand U3049 (N_3049,In_440,In_935);
xnor U3050 (N_3050,In_568,In_440);
xnor U3051 (N_3051,In_114,In_580);
and U3052 (N_3052,In_47,In_76);
and U3053 (N_3053,In_183,In_150);
or U3054 (N_3054,In_351,In_720);
nand U3055 (N_3055,In_460,In_796);
or U3056 (N_3056,In_638,In_560);
nand U3057 (N_3057,In_881,In_777);
or U3058 (N_3058,In_84,In_911);
xnor U3059 (N_3059,In_519,In_997);
nand U3060 (N_3060,In_448,In_1);
or U3061 (N_3061,In_263,In_619);
nand U3062 (N_3062,In_476,In_389);
and U3063 (N_3063,In_672,In_932);
or U3064 (N_3064,In_918,In_758);
or U3065 (N_3065,In_925,In_136);
nor U3066 (N_3066,In_118,In_262);
or U3067 (N_3067,In_756,In_55);
xnor U3068 (N_3068,In_261,In_363);
nand U3069 (N_3069,In_463,In_15);
and U3070 (N_3070,In_47,In_370);
nor U3071 (N_3071,In_936,In_988);
and U3072 (N_3072,In_963,In_6);
and U3073 (N_3073,In_870,In_413);
or U3074 (N_3074,In_841,In_996);
nor U3075 (N_3075,In_351,In_911);
nand U3076 (N_3076,In_532,In_663);
nand U3077 (N_3077,In_462,In_801);
and U3078 (N_3078,In_140,In_328);
and U3079 (N_3079,In_822,In_592);
and U3080 (N_3080,In_356,In_140);
nand U3081 (N_3081,In_82,In_243);
or U3082 (N_3082,In_721,In_154);
nand U3083 (N_3083,In_347,In_165);
or U3084 (N_3084,In_292,In_601);
nor U3085 (N_3085,In_313,In_135);
nor U3086 (N_3086,In_523,In_354);
and U3087 (N_3087,In_919,In_206);
or U3088 (N_3088,In_343,In_764);
nor U3089 (N_3089,In_169,In_50);
nor U3090 (N_3090,In_504,In_506);
nor U3091 (N_3091,In_667,In_994);
nor U3092 (N_3092,In_332,In_998);
or U3093 (N_3093,In_376,In_61);
nand U3094 (N_3094,In_452,In_855);
or U3095 (N_3095,In_169,In_509);
or U3096 (N_3096,In_763,In_650);
or U3097 (N_3097,In_445,In_458);
nor U3098 (N_3098,In_936,In_558);
nor U3099 (N_3099,In_834,In_227);
and U3100 (N_3100,In_524,In_233);
nand U3101 (N_3101,In_620,In_428);
nand U3102 (N_3102,In_274,In_730);
and U3103 (N_3103,In_862,In_434);
and U3104 (N_3104,In_539,In_181);
or U3105 (N_3105,In_755,In_852);
or U3106 (N_3106,In_528,In_795);
nand U3107 (N_3107,In_503,In_99);
nor U3108 (N_3108,In_229,In_185);
nand U3109 (N_3109,In_614,In_61);
and U3110 (N_3110,In_682,In_150);
xor U3111 (N_3111,In_550,In_209);
or U3112 (N_3112,In_647,In_296);
or U3113 (N_3113,In_287,In_478);
or U3114 (N_3114,In_28,In_918);
nand U3115 (N_3115,In_220,In_862);
or U3116 (N_3116,In_258,In_998);
or U3117 (N_3117,In_911,In_606);
nand U3118 (N_3118,In_50,In_82);
or U3119 (N_3119,In_974,In_528);
xnor U3120 (N_3120,In_531,In_69);
or U3121 (N_3121,In_700,In_990);
xnor U3122 (N_3122,In_494,In_145);
or U3123 (N_3123,In_152,In_211);
nand U3124 (N_3124,In_561,In_351);
or U3125 (N_3125,In_214,In_253);
or U3126 (N_3126,In_103,In_936);
nand U3127 (N_3127,In_639,In_547);
nand U3128 (N_3128,In_84,In_372);
and U3129 (N_3129,In_204,In_940);
xnor U3130 (N_3130,In_672,In_884);
nand U3131 (N_3131,In_543,In_703);
and U3132 (N_3132,In_737,In_895);
nand U3133 (N_3133,In_403,In_220);
or U3134 (N_3134,In_276,In_408);
or U3135 (N_3135,In_709,In_977);
or U3136 (N_3136,In_18,In_497);
nor U3137 (N_3137,In_631,In_296);
nor U3138 (N_3138,In_594,In_266);
and U3139 (N_3139,In_594,In_865);
nand U3140 (N_3140,In_171,In_955);
nor U3141 (N_3141,In_754,In_344);
nor U3142 (N_3142,In_62,In_467);
or U3143 (N_3143,In_889,In_309);
nand U3144 (N_3144,In_964,In_457);
or U3145 (N_3145,In_487,In_853);
nand U3146 (N_3146,In_953,In_611);
and U3147 (N_3147,In_360,In_914);
or U3148 (N_3148,In_285,In_619);
xnor U3149 (N_3149,In_633,In_869);
nand U3150 (N_3150,In_781,In_597);
and U3151 (N_3151,In_974,In_764);
and U3152 (N_3152,In_849,In_632);
xor U3153 (N_3153,In_824,In_174);
and U3154 (N_3154,In_390,In_690);
xor U3155 (N_3155,In_403,In_532);
nand U3156 (N_3156,In_911,In_567);
and U3157 (N_3157,In_964,In_385);
or U3158 (N_3158,In_592,In_178);
and U3159 (N_3159,In_609,In_348);
or U3160 (N_3160,In_78,In_312);
nor U3161 (N_3161,In_114,In_158);
nor U3162 (N_3162,In_181,In_841);
nor U3163 (N_3163,In_620,In_493);
nor U3164 (N_3164,In_984,In_429);
and U3165 (N_3165,In_379,In_938);
nor U3166 (N_3166,In_586,In_574);
nor U3167 (N_3167,In_216,In_498);
and U3168 (N_3168,In_189,In_126);
nor U3169 (N_3169,In_725,In_189);
or U3170 (N_3170,In_666,In_658);
nor U3171 (N_3171,In_335,In_484);
and U3172 (N_3172,In_963,In_108);
nand U3173 (N_3173,In_777,In_285);
and U3174 (N_3174,In_570,In_225);
nor U3175 (N_3175,In_476,In_936);
and U3176 (N_3176,In_430,In_913);
or U3177 (N_3177,In_894,In_623);
nor U3178 (N_3178,In_818,In_813);
nand U3179 (N_3179,In_638,In_563);
nand U3180 (N_3180,In_918,In_113);
nand U3181 (N_3181,In_957,In_592);
xnor U3182 (N_3182,In_947,In_591);
and U3183 (N_3183,In_92,In_284);
nand U3184 (N_3184,In_285,In_983);
and U3185 (N_3185,In_670,In_668);
nor U3186 (N_3186,In_960,In_451);
and U3187 (N_3187,In_889,In_618);
xor U3188 (N_3188,In_571,In_92);
or U3189 (N_3189,In_199,In_86);
nand U3190 (N_3190,In_227,In_578);
or U3191 (N_3191,In_510,In_771);
nor U3192 (N_3192,In_492,In_493);
or U3193 (N_3193,In_654,In_825);
nand U3194 (N_3194,In_872,In_394);
nor U3195 (N_3195,In_242,In_841);
or U3196 (N_3196,In_490,In_140);
and U3197 (N_3197,In_815,In_213);
xnor U3198 (N_3198,In_561,In_485);
xor U3199 (N_3199,In_456,In_196);
or U3200 (N_3200,In_755,In_169);
nor U3201 (N_3201,In_578,In_952);
nand U3202 (N_3202,In_230,In_551);
nor U3203 (N_3203,In_266,In_264);
nor U3204 (N_3204,In_539,In_96);
and U3205 (N_3205,In_596,In_807);
nand U3206 (N_3206,In_599,In_352);
nor U3207 (N_3207,In_371,In_726);
or U3208 (N_3208,In_179,In_812);
or U3209 (N_3209,In_503,In_3);
xnor U3210 (N_3210,In_20,In_428);
nor U3211 (N_3211,In_198,In_278);
or U3212 (N_3212,In_37,In_281);
and U3213 (N_3213,In_710,In_930);
xor U3214 (N_3214,In_49,In_883);
nand U3215 (N_3215,In_528,In_636);
nand U3216 (N_3216,In_822,In_696);
and U3217 (N_3217,In_552,In_25);
and U3218 (N_3218,In_629,In_595);
or U3219 (N_3219,In_478,In_911);
nand U3220 (N_3220,In_392,In_381);
nor U3221 (N_3221,In_867,In_90);
nor U3222 (N_3222,In_802,In_236);
xnor U3223 (N_3223,In_185,In_583);
and U3224 (N_3224,In_496,In_712);
nor U3225 (N_3225,In_890,In_481);
nand U3226 (N_3226,In_130,In_537);
or U3227 (N_3227,In_682,In_242);
nor U3228 (N_3228,In_856,In_296);
and U3229 (N_3229,In_306,In_317);
xor U3230 (N_3230,In_774,In_267);
nor U3231 (N_3231,In_942,In_129);
nand U3232 (N_3232,In_579,In_335);
and U3233 (N_3233,In_544,In_941);
nor U3234 (N_3234,In_235,In_156);
nor U3235 (N_3235,In_495,In_96);
and U3236 (N_3236,In_751,In_218);
and U3237 (N_3237,In_672,In_729);
and U3238 (N_3238,In_585,In_966);
nand U3239 (N_3239,In_162,In_536);
and U3240 (N_3240,In_686,In_823);
and U3241 (N_3241,In_883,In_320);
and U3242 (N_3242,In_46,In_551);
or U3243 (N_3243,In_543,In_322);
nor U3244 (N_3244,In_860,In_574);
nor U3245 (N_3245,In_282,In_685);
nand U3246 (N_3246,In_683,In_324);
and U3247 (N_3247,In_251,In_603);
nand U3248 (N_3248,In_615,In_968);
nand U3249 (N_3249,In_429,In_616);
nand U3250 (N_3250,In_730,In_445);
xor U3251 (N_3251,In_685,In_226);
xor U3252 (N_3252,In_110,In_121);
nor U3253 (N_3253,In_761,In_839);
nand U3254 (N_3254,In_992,In_945);
or U3255 (N_3255,In_638,In_878);
xnor U3256 (N_3256,In_329,In_597);
nor U3257 (N_3257,In_440,In_195);
and U3258 (N_3258,In_608,In_440);
or U3259 (N_3259,In_141,In_416);
nor U3260 (N_3260,In_329,In_896);
xor U3261 (N_3261,In_722,In_995);
and U3262 (N_3262,In_846,In_265);
or U3263 (N_3263,In_878,In_170);
nor U3264 (N_3264,In_586,In_230);
or U3265 (N_3265,In_620,In_677);
nor U3266 (N_3266,In_219,In_553);
nor U3267 (N_3267,In_126,In_304);
nand U3268 (N_3268,In_960,In_554);
or U3269 (N_3269,In_406,In_462);
nand U3270 (N_3270,In_766,In_956);
and U3271 (N_3271,In_624,In_891);
nand U3272 (N_3272,In_990,In_604);
or U3273 (N_3273,In_804,In_337);
and U3274 (N_3274,In_666,In_413);
nor U3275 (N_3275,In_702,In_345);
nor U3276 (N_3276,In_131,In_854);
nand U3277 (N_3277,In_955,In_184);
and U3278 (N_3278,In_648,In_764);
xnor U3279 (N_3279,In_119,In_386);
nand U3280 (N_3280,In_647,In_765);
nand U3281 (N_3281,In_439,In_36);
or U3282 (N_3282,In_446,In_194);
or U3283 (N_3283,In_800,In_268);
or U3284 (N_3284,In_858,In_121);
nor U3285 (N_3285,In_820,In_38);
nor U3286 (N_3286,In_91,In_179);
xor U3287 (N_3287,In_599,In_810);
nand U3288 (N_3288,In_778,In_920);
nand U3289 (N_3289,In_529,In_360);
and U3290 (N_3290,In_543,In_968);
nor U3291 (N_3291,In_600,In_607);
xnor U3292 (N_3292,In_153,In_196);
nor U3293 (N_3293,In_793,In_877);
and U3294 (N_3294,In_555,In_924);
nor U3295 (N_3295,In_581,In_724);
and U3296 (N_3296,In_428,In_34);
nand U3297 (N_3297,In_182,In_478);
and U3298 (N_3298,In_608,In_16);
nand U3299 (N_3299,In_726,In_876);
and U3300 (N_3300,In_775,In_326);
xnor U3301 (N_3301,In_653,In_800);
or U3302 (N_3302,In_394,In_580);
and U3303 (N_3303,In_492,In_301);
and U3304 (N_3304,In_22,In_238);
or U3305 (N_3305,In_982,In_494);
or U3306 (N_3306,In_240,In_196);
nand U3307 (N_3307,In_471,In_578);
nor U3308 (N_3308,In_573,In_145);
nand U3309 (N_3309,In_230,In_403);
or U3310 (N_3310,In_675,In_942);
nand U3311 (N_3311,In_495,In_502);
nor U3312 (N_3312,In_308,In_242);
nand U3313 (N_3313,In_315,In_419);
xnor U3314 (N_3314,In_718,In_603);
and U3315 (N_3315,In_754,In_378);
nand U3316 (N_3316,In_157,In_872);
nand U3317 (N_3317,In_733,In_80);
xor U3318 (N_3318,In_927,In_605);
nand U3319 (N_3319,In_355,In_502);
xnor U3320 (N_3320,In_111,In_571);
or U3321 (N_3321,In_489,In_225);
and U3322 (N_3322,In_625,In_535);
nand U3323 (N_3323,In_302,In_530);
and U3324 (N_3324,In_796,In_749);
or U3325 (N_3325,In_653,In_526);
nor U3326 (N_3326,In_318,In_583);
nand U3327 (N_3327,In_703,In_173);
nand U3328 (N_3328,In_502,In_309);
nor U3329 (N_3329,In_711,In_569);
nand U3330 (N_3330,In_492,In_162);
or U3331 (N_3331,In_572,In_124);
and U3332 (N_3332,In_896,In_710);
nand U3333 (N_3333,In_528,In_28);
and U3334 (N_3334,In_446,In_792);
and U3335 (N_3335,In_835,In_269);
and U3336 (N_3336,In_89,In_517);
or U3337 (N_3337,In_858,In_494);
and U3338 (N_3338,In_464,In_823);
and U3339 (N_3339,In_236,In_296);
nor U3340 (N_3340,In_998,In_899);
or U3341 (N_3341,In_873,In_717);
xor U3342 (N_3342,In_546,In_557);
xnor U3343 (N_3343,In_784,In_63);
or U3344 (N_3344,In_831,In_240);
xnor U3345 (N_3345,In_499,In_474);
and U3346 (N_3346,In_768,In_848);
or U3347 (N_3347,In_707,In_739);
and U3348 (N_3348,In_849,In_718);
xor U3349 (N_3349,In_318,In_854);
and U3350 (N_3350,In_302,In_935);
nor U3351 (N_3351,In_535,In_396);
nor U3352 (N_3352,In_307,In_971);
nor U3353 (N_3353,In_335,In_629);
nor U3354 (N_3354,In_949,In_577);
nor U3355 (N_3355,In_792,In_129);
nand U3356 (N_3356,In_231,In_76);
nor U3357 (N_3357,In_128,In_164);
or U3358 (N_3358,In_350,In_550);
nand U3359 (N_3359,In_193,In_67);
nor U3360 (N_3360,In_1,In_522);
and U3361 (N_3361,In_35,In_740);
nor U3362 (N_3362,In_533,In_337);
nor U3363 (N_3363,In_773,In_990);
or U3364 (N_3364,In_894,In_443);
nand U3365 (N_3365,In_556,In_510);
and U3366 (N_3366,In_570,In_315);
nor U3367 (N_3367,In_500,In_958);
or U3368 (N_3368,In_281,In_190);
nor U3369 (N_3369,In_353,In_136);
or U3370 (N_3370,In_838,In_890);
nor U3371 (N_3371,In_946,In_720);
nand U3372 (N_3372,In_117,In_983);
and U3373 (N_3373,In_640,In_631);
nand U3374 (N_3374,In_25,In_787);
nor U3375 (N_3375,In_300,In_754);
and U3376 (N_3376,In_296,In_71);
or U3377 (N_3377,In_706,In_690);
xor U3378 (N_3378,In_106,In_798);
or U3379 (N_3379,In_808,In_92);
nor U3380 (N_3380,In_556,In_377);
or U3381 (N_3381,In_189,In_3);
nor U3382 (N_3382,In_460,In_219);
and U3383 (N_3383,In_973,In_982);
or U3384 (N_3384,In_798,In_504);
and U3385 (N_3385,In_697,In_270);
or U3386 (N_3386,In_605,In_945);
nand U3387 (N_3387,In_785,In_387);
and U3388 (N_3388,In_537,In_799);
and U3389 (N_3389,In_496,In_948);
nor U3390 (N_3390,In_372,In_115);
nand U3391 (N_3391,In_602,In_709);
xor U3392 (N_3392,In_309,In_135);
nand U3393 (N_3393,In_569,In_221);
or U3394 (N_3394,In_306,In_279);
nand U3395 (N_3395,In_937,In_194);
nand U3396 (N_3396,In_424,In_891);
and U3397 (N_3397,In_657,In_533);
or U3398 (N_3398,In_589,In_621);
nor U3399 (N_3399,In_31,In_77);
or U3400 (N_3400,In_27,In_209);
nor U3401 (N_3401,In_116,In_315);
or U3402 (N_3402,In_98,In_758);
xor U3403 (N_3403,In_293,In_601);
or U3404 (N_3404,In_704,In_753);
nand U3405 (N_3405,In_628,In_819);
and U3406 (N_3406,In_739,In_770);
nor U3407 (N_3407,In_209,In_983);
nand U3408 (N_3408,In_236,In_763);
or U3409 (N_3409,In_659,In_685);
and U3410 (N_3410,In_993,In_896);
xor U3411 (N_3411,In_568,In_886);
xnor U3412 (N_3412,In_788,In_337);
nor U3413 (N_3413,In_678,In_18);
and U3414 (N_3414,In_153,In_479);
nand U3415 (N_3415,In_628,In_43);
nor U3416 (N_3416,In_282,In_258);
or U3417 (N_3417,In_974,In_600);
or U3418 (N_3418,In_739,In_130);
and U3419 (N_3419,In_431,In_848);
xnor U3420 (N_3420,In_152,In_871);
nand U3421 (N_3421,In_429,In_361);
and U3422 (N_3422,In_294,In_901);
or U3423 (N_3423,In_417,In_380);
or U3424 (N_3424,In_876,In_241);
nand U3425 (N_3425,In_946,In_880);
or U3426 (N_3426,In_570,In_805);
or U3427 (N_3427,In_777,In_843);
nor U3428 (N_3428,In_432,In_344);
xnor U3429 (N_3429,In_78,In_922);
nor U3430 (N_3430,In_114,In_539);
nor U3431 (N_3431,In_663,In_30);
xor U3432 (N_3432,In_691,In_145);
and U3433 (N_3433,In_681,In_199);
xnor U3434 (N_3434,In_142,In_992);
or U3435 (N_3435,In_588,In_961);
nor U3436 (N_3436,In_569,In_374);
nor U3437 (N_3437,In_713,In_131);
or U3438 (N_3438,In_278,In_919);
xnor U3439 (N_3439,In_6,In_672);
or U3440 (N_3440,In_704,In_308);
and U3441 (N_3441,In_567,In_378);
and U3442 (N_3442,In_657,In_658);
nor U3443 (N_3443,In_553,In_472);
and U3444 (N_3444,In_592,In_524);
nand U3445 (N_3445,In_930,In_323);
nor U3446 (N_3446,In_752,In_526);
and U3447 (N_3447,In_508,In_75);
xnor U3448 (N_3448,In_909,In_434);
or U3449 (N_3449,In_84,In_817);
and U3450 (N_3450,In_794,In_506);
nand U3451 (N_3451,In_396,In_968);
nor U3452 (N_3452,In_950,In_478);
nand U3453 (N_3453,In_267,In_625);
nor U3454 (N_3454,In_930,In_272);
nand U3455 (N_3455,In_982,In_955);
nor U3456 (N_3456,In_598,In_64);
or U3457 (N_3457,In_839,In_830);
nor U3458 (N_3458,In_622,In_516);
or U3459 (N_3459,In_125,In_394);
xnor U3460 (N_3460,In_666,In_558);
and U3461 (N_3461,In_705,In_507);
nor U3462 (N_3462,In_277,In_777);
xor U3463 (N_3463,In_405,In_744);
nor U3464 (N_3464,In_207,In_255);
and U3465 (N_3465,In_414,In_920);
nand U3466 (N_3466,In_981,In_767);
or U3467 (N_3467,In_578,In_27);
and U3468 (N_3468,In_843,In_649);
or U3469 (N_3469,In_422,In_601);
nor U3470 (N_3470,In_872,In_13);
nand U3471 (N_3471,In_292,In_121);
nor U3472 (N_3472,In_214,In_170);
xor U3473 (N_3473,In_680,In_129);
nor U3474 (N_3474,In_230,In_728);
and U3475 (N_3475,In_278,In_141);
nand U3476 (N_3476,In_933,In_764);
and U3477 (N_3477,In_135,In_958);
nor U3478 (N_3478,In_211,In_862);
nand U3479 (N_3479,In_538,In_962);
or U3480 (N_3480,In_962,In_763);
nand U3481 (N_3481,In_295,In_379);
xor U3482 (N_3482,In_119,In_518);
nor U3483 (N_3483,In_349,In_593);
or U3484 (N_3484,In_325,In_436);
nor U3485 (N_3485,In_249,In_291);
or U3486 (N_3486,In_912,In_214);
nor U3487 (N_3487,In_90,In_187);
and U3488 (N_3488,In_881,In_316);
and U3489 (N_3489,In_553,In_308);
nor U3490 (N_3490,In_783,In_158);
xnor U3491 (N_3491,In_68,In_781);
nand U3492 (N_3492,In_595,In_386);
nor U3493 (N_3493,In_586,In_981);
or U3494 (N_3494,In_770,In_117);
or U3495 (N_3495,In_875,In_3);
and U3496 (N_3496,In_49,In_275);
nor U3497 (N_3497,In_95,In_421);
xnor U3498 (N_3498,In_54,In_996);
and U3499 (N_3499,In_168,In_337);
nor U3500 (N_3500,In_517,In_219);
and U3501 (N_3501,In_625,In_186);
and U3502 (N_3502,In_379,In_848);
nand U3503 (N_3503,In_599,In_379);
nor U3504 (N_3504,In_463,In_956);
nor U3505 (N_3505,In_593,In_179);
or U3506 (N_3506,In_168,In_213);
or U3507 (N_3507,In_808,In_600);
nand U3508 (N_3508,In_355,In_922);
nand U3509 (N_3509,In_158,In_597);
and U3510 (N_3510,In_711,In_36);
or U3511 (N_3511,In_190,In_918);
nand U3512 (N_3512,In_358,In_173);
xor U3513 (N_3513,In_437,In_64);
nand U3514 (N_3514,In_683,In_291);
or U3515 (N_3515,In_556,In_787);
or U3516 (N_3516,In_824,In_540);
or U3517 (N_3517,In_969,In_979);
and U3518 (N_3518,In_562,In_671);
or U3519 (N_3519,In_491,In_137);
or U3520 (N_3520,In_564,In_180);
and U3521 (N_3521,In_490,In_155);
and U3522 (N_3522,In_306,In_870);
nand U3523 (N_3523,In_49,In_120);
and U3524 (N_3524,In_901,In_966);
nor U3525 (N_3525,In_318,In_385);
or U3526 (N_3526,In_135,In_937);
and U3527 (N_3527,In_805,In_664);
or U3528 (N_3528,In_39,In_569);
and U3529 (N_3529,In_119,In_864);
nor U3530 (N_3530,In_948,In_388);
or U3531 (N_3531,In_48,In_808);
xor U3532 (N_3532,In_139,In_175);
xor U3533 (N_3533,In_400,In_588);
or U3534 (N_3534,In_599,In_774);
nand U3535 (N_3535,In_168,In_271);
or U3536 (N_3536,In_873,In_397);
nor U3537 (N_3537,In_876,In_284);
or U3538 (N_3538,In_139,In_81);
and U3539 (N_3539,In_972,In_960);
or U3540 (N_3540,In_996,In_9);
xor U3541 (N_3541,In_871,In_318);
and U3542 (N_3542,In_228,In_953);
or U3543 (N_3543,In_606,In_835);
nand U3544 (N_3544,In_375,In_804);
or U3545 (N_3545,In_127,In_637);
nor U3546 (N_3546,In_330,In_562);
or U3547 (N_3547,In_483,In_994);
nand U3548 (N_3548,In_460,In_247);
and U3549 (N_3549,In_855,In_293);
or U3550 (N_3550,In_322,In_380);
nand U3551 (N_3551,In_175,In_372);
nand U3552 (N_3552,In_936,In_919);
xor U3553 (N_3553,In_205,In_80);
or U3554 (N_3554,In_138,In_184);
nand U3555 (N_3555,In_613,In_567);
nor U3556 (N_3556,In_472,In_13);
or U3557 (N_3557,In_481,In_780);
nand U3558 (N_3558,In_977,In_531);
nor U3559 (N_3559,In_471,In_659);
or U3560 (N_3560,In_790,In_82);
xor U3561 (N_3561,In_971,In_131);
nor U3562 (N_3562,In_694,In_230);
nor U3563 (N_3563,In_778,In_158);
nor U3564 (N_3564,In_3,In_170);
nand U3565 (N_3565,In_437,In_579);
nor U3566 (N_3566,In_202,In_512);
and U3567 (N_3567,In_716,In_194);
or U3568 (N_3568,In_160,In_962);
nor U3569 (N_3569,In_918,In_346);
and U3570 (N_3570,In_202,In_999);
nand U3571 (N_3571,In_822,In_937);
nor U3572 (N_3572,In_91,In_711);
or U3573 (N_3573,In_808,In_852);
nor U3574 (N_3574,In_90,In_23);
or U3575 (N_3575,In_601,In_672);
or U3576 (N_3576,In_575,In_28);
and U3577 (N_3577,In_305,In_866);
and U3578 (N_3578,In_557,In_142);
and U3579 (N_3579,In_720,In_999);
nor U3580 (N_3580,In_356,In_738);
nor U3581 (N_3581,In_821,In_753);
or U3582 (N_3582,In_491,In_700);
nand U3583 (N_3583,In_643,In_386);
nand U3584 (N_3584,In_991,In_242);
and U3585 (N_3585,In_300,In_652);
nand U3586 (N_3586,In_700,In_714);
and U3587 (N_3587,In_618,In_226);
and U3588 (N_3588,In_566,In_870);
or U3589 (N_3589,In_457,In_473);
nand U3590 (N_3590,In_306,In_574);
or U3591 (N_3591,In_189,In_176);
nand U3592 (N_3592,In_164,In_181);
and U3593 (N_3593,In_127,In_526);
nand U3594 (N_3594,In_786,In_464);
or U3595 (N_3595,In_885,In_52);
and U3596 (N_3596,In_367,In_768);
xor U3597 (N_3597,In_596,In_713);
nor U3598 (N_3598,In_759,In_45);
or U3599 (N_3599,In_208,In_377);
and U3600 (N_3600,In_791,In_379);
nand U3601 (N_3601,In_117,In_369);
and U3602 (N_3602,In_886,In_781);
nand U3603 (N_3603,In_98,In_440);
xnor U3604 (N_3604,In_343,In_650);
or U3605 (N_3605,In_608,In_890);
nor U3606 (N_3606,In_254,In_89);
nor U3607 (N_3607,In_885,In_447);
nor U3608 (N_3608,In_234,In_904);
nand U3609 (N_3609,In_753,In_56);
xor U3610 (N_3610,In_19,In_873);
xor U3611 (N_3611,In_738,In_871);
nor U3612 (N_3612,In_528,In_560);
nand U3613 (N_3613,In_995,In_655);
and U3614 (N_3614,In_424,In_787);
and U3615 (N_3615,In_570,In_258);
nand U3616 (N_3616,In_824,In_667);
nor U3617 (N_3617,In_436,In_800);
nand U3618 (N_3618,In_607,In_245);
xnor U3619 (N_3619,In_749,In_624);
and U3620 (N_3620,In_55,In_463);
or U3621 (N_3621,In_765,In_525);
and U3622 (N_3622,In_954,In_24);
nand U3623 (N_3623,In_941,In_245);
nand U3624 (N_3624,In_284,In_339);
and U3625 (N_3625,In_183,In_958);
xnor U3626 (N_3626,In_647,In_35);
or U3627 (N_3627,In_978,In_445);
xnor U3628 (N_3628,In_313,In_522);
or U3629 (N_3629,In_9,In_429);
or U3630 (N_3630,In_135,In_71);
xor U3631 (N_3631,In_551,In_120);
nor U3632 (N_3632,In_721,In_714);
or U3633 (N_3633,In_627,In_492);
or U3634 (N_3634,In_381,In_283);
nor U3635 (N_3635,In_567,In_699);
nand U3636 (N_3636,In_769,In_868);
nand U3637 (N_3637,In_217,In_338);
nor U3638 (N_3638,In_663,In_317);
nor U3639 (N_3639,In_356,In_91);
xnor U3640 (N_3640,In_644,In_582);
nor U3641 (N_3641,In_825,In_455);
and U3642 (N_3642,In_100,In_792);
or U3643 (N_3643,In_62,In_68);
nor U3644 (N_3644,In_333,In_917);
nor U3645 (N_3645,In_508,In_650);
or U3646 (N_3646,In_384,In_612);
nor U3647 (N_3647,In_580,In_24);
and U3648 (N_3648,In_170,In_62);
nand U3649 (N_3649,In_290,In_438);
nand U3650 (N_3650,In_613,In_950);
nor U3651 (N_3651,In_36,In_391);
nor U3652 (N_3652,In_90,In_283);
or U3653 (N_3653,In_488,In_822);
and U3654 (N_3654,In_354,In_477);
nor U3655 (N_3655,In_686,In_671);
or U3656 (N_3656,In_334,In_855);
nor U3657 (N_3657,In_618,In_294);
xor U3658 (N_3658,In_77,In_803);
and U3659 (N_3659,In_193,In_121);
nor U3660 (N_3660,In_526,In_61);
nor U3661 (N_3661,In_147,In_400);
or U3662 (N_3662,In_6,In_391);
or U3663 (N_3663,In_975,In_833);
nand U3664 (N_3664,In_688,In_101);
and U3665 (N_3665,In_797,In_761);
or U3666 (N_3666,In_621,In_599);
xor U3667 (N_3667,In_397,In_114);
nand U3668 (N_3668,In_702,In_208);
or U3669 (N_3669,In_48,In_690);
nor U3670 (N_3670,In_139,In_675);
and U3671 (N_3671,In_173,In_374);
xor U3672 (N_3672,In_802,In_694);
or U3673 (N_3673,In_885,In_830);
nand U3674 (N_3674,In_415,In_576);
nor U3675 (N_3675,In_295,In_202);
and U3676 (N_3676,In_822,In_474);
and U3677 (N_3677,In_732,In_667);
nand U3678 (N_3678,In_979,In_32);
nor U3679 (N_3679,In_140,In_902);
nand U3680 (N_3680,In_513,In_49);
nor U3681 (N_3681,In_75,In_501);
and U3682 (N_3682,In_563,In_191);
nor U3683 (N_3683,In_131,In_248);
and U3684 (N_3684,In_374,In_393);
nor U3685 (N_3685,In_400,In_526);
nand U3686 (N_3686,In_834,In_320);
nand U3687 (N_3687,In_805,In_44);
or U3688 (N_3688,In_462,In_279);
and U3689 (N_3689,In_375,In_808);
nor U3690 (N_3690,In_970,In_456);
or U3691 (N_3691,In_804,In_372);
and U3692 (N_3692,In_344,In_755);
nor U3693 (N_3693,In_633,In_270);
or U3694 (N_3694,In_811,In_3);
nand U3695 (N_3695,In_241,In_58);
nand U3696 (N_3696,In_422,In_735);
and U3697 (N_3697,In_542,In_648);
nor U3698 (N_3698,In_970,In_774);
nand U3699 (N_3699,In_461,In_984);
and U3700 (N_3700,In_556,In_894);
nand U3701 (N_3701,In_224,In_851);
nor U3702 (N_3702,In_134,In_206);
or U3703 (N_3703,In_867,In_964);
nor U3704 (N_3704,In_769,In_824);
and U3705 (N_3705,In_629,In_160);
nand U3706 (N_3706,In_159,In_547);
xnor U3707 (N_3707,In_319,In_585);
nor U3708 (N_3708,In_364,In_60);
and U3709 (N_3709,In_64,In_484);
nand U3710 (N_3710,In_964,In_801);
and U3711 (N_3711,In_254,In_735);
nand U3712 (N_3712,In_282,In_532);
and U3713 (N_3713,In_18,In_575);
nand U3714 (N_3714,In_419,In_201);
nor U3715 (N_3715,In_386,In_361);
nand U3716 (N_3716,In_106,In_325);
nor U3717 (N_3717,In_134,In_471);
nand U3718 (N_3718,In_154,In_573);
nand U3719 (N_3719,In_368,In_651);
nor U3720 (N_3720,In_9,In_182);
nand U3721 (N_3721,In_850,In_432);
or U3722 (N_3722,In_743,In_782);
nor U3723 (N_3723,In_575,In_251);
and U3724 (N_3724,In_672,In_753);
and U3725 (N_3725,In_152,In_411);
and U3726 (N_3726,In_484,In_273);
nand U3727 (N_3727,In_154,In_24);
or U3728 (N_3728,In_468,In_660);
and U3729 (N_3729,In_240,In_146);
nand U3730 (N_3730,In_935,In_526);
nor U3731 (N_3731,In_841,In_700);
nor U3732 (N_3732,In_682,In_840);
xnor U3733 (N_3733,In_424,In_434);
or U3734 (N_3734,In_699,In_678);
and U3735 (N_3735,In_428,In_703);
nor U3736 (N_3736,In_94,In_324);
and U3737 (N_3737,In_152,In_117);
and U3738 (N_3738,In_785,In_226);
or U3739 (N_3739,In_611,In_348);
and U3740 (N_3740,In_273,In_680);
nand U3741 (N_3741,In_224,In_313);
or U3742 (N_3742,In_687,In_990);
nor U3743 (N_3743,In_719,In_701);
xor U3744 (N_3744,In_281,In_882);
or U3745 (N_3745,In_707,In_53);
xor U3746 (N_3746,In_247,In_649);
and U3747 (N_3747,In_110,In_635);
xor U3748 (N_3748,In_184,In_50);
nor U3749 (N_3749,In_527,In_518);
nor U3750 (N_3750,In_259,In_33);
nand U3751 (N_3751,In_739,In_15);
or U3752 (N_3752,In_697,In_175);
and U3753 (N_3753,In_103,In_772);
nor U3754 (N_3754,In_282,In_367);
nand U3755 (N_3755,In_937,In_405);
and U3756 (N_3756,In_985,In_613);
nor U3757 (N_3757,In_801,In_685);
or U3758 (N_3758,In_652,In_337);
or U3759 (N_3759,In_925,In_728);
nand U3760 (N_3760,In_427,In_610);
or U3761 (N_3761,In_995,In_143);
and U3762 (N_3762,In_421,In_112);
nand U3763 (N_3763,In_292,In_904);
nor U3764 (N_3764,In_771,In_298);
nand U3765 (N_3765,In_654,In_312);
and U3766 (N_3766,In_775,In_821);
or U3767 (N_3767,In_85,In_99);
and U3768 (N_3768,In_996,In_819);
nand U3769 (N_3769,In_729,In_824);
or U3770 (N_3770,In_831,In_703);
nor U3771 (N_3771,In_9,In_104);
nor U3772 (N_3772,In_547,In_27);
and U3773 (N_3773,In_866,In_802);
nand U3774 (N_3774,In_697,In_91);
nand U3775 (N_3775,In_407,In_154);
nor U3776 (N_3776,In_928,In_855);
and U3777 (N_3777,In_77,In_918);
and U3778 (N_3778,In_948,In_694);
or U3779 (N_3779,In_204,In_174);
xor U3780 (N_3780,In_45,In_795);
xnor U3781 (N_3781,In_264,In_866);
or U3782 (N_3782,In_975,In_136);
or U3783 (N_3783,In_600,In_763);
and U3784 (N_3784,In_939,In_593);
nand U3785 (N_3785,In_982,In_52);
nand U3786 (N_3786,In_845,In_145);
nor U3787 (N_3787,In_742,In_664);
and U3788 (N_3788,In_961,In_376);
xor U3789 (N_3789,In_427,In_360);
nand U3790 (N_3790,In_190,In_595);
and U3791 (N_3791,In_399,In_880);
nor U3792 (N_3792,In_43,In_507);
xnor U3793 (N_3793,In_373,In_493);
nor U3794 (N_3794,In_344,In_75);
or U3795 (N_3795,In_581,In_797);
nand U3796 (N_3796,In_17,In_295);
or U3797 (N_3797,In_264,In_296);
or U3798 (N_3798,In_992,In_207);
nand U3799 (N_3799,In_309,In_457);
and U3800 (N_3800,In_682,In_118);
xnor U3801 (N_3801,In_176,In_411);
and U3802 (N_3802,In_541,In_702);
or U3803 (N_3803,In_737,In_92);
or U3804 (N_3804,In_45,In_585);
nor U3805 (N_3805,In_621,In_198);
or U3806 (N_3806,In_848,In_812);
nor U3807 (N_3807,In_333,In_606);
xor U3808 (N_3808,In_975,In_396);
and U3809 (N_3809,In_707,In_954);
nand U3810 (N_3810,In_808,In_43);
and U3811 (N_3811,In_222,In_470);
nor U3812 (N_3812,In_92,In_503);
nor U3813 (N_3813,In_27,In_316);
nor U3814 (N_3814,In_440,In_520);
nor U3815 (N_3815,In_554,In_538);
nand U3816 (N_3816,In_502,In_741);
or U3817 (N_3817,In_641,In_993);
nand U3818 (N_3818,In_613,In_201);
and U3819 (N_3819,In_629,In_989);
and U3820 (N_3820,In_550,In_525);
nand U3821 (N_3821,In_397,In_256);
nor U3822 (N_3822,In_405,In_438);
and U3823 (N_3823,In_851,In_149);
nand U3824 (N_3824,In_822,In_600);
nor U3825 (N_3825,In_194,In_361);
xor U3826 (N_3826,In_65,In_559);
and U3827 (N_3827,In_240,In_552);
and U3828 (N_3828,In_632,In_115);
nand U3829 (N_3829,In_478,In_948);
nand U3830 (N_3830,In_273,In_621);
nand U3831 (N_3831,In_530,In_485);
or U3832 (N_3832,In_575,In_979);
or U3833 (N_3833,In_304,In_717);
xnor U3834 (N_3834,In_326,In_43);
nor U3835 (N_3835,In_194,In_304);
or U3836 (N_3836,In_176,In_373);
or U3837 (N_3837,In_928,In_844);
nand U3838 (N_3838,In_811,In_734);
and U3839 (N_3839,In_633,In_598);
nor U3840 (N_3840,In_668,In_874);
or U3841 (N_3841,In_777,In_201);
nor U3842 (N_3842,In_524,In_412);
nand U3843 (N_3843,In_864,In_644);
or U3844 (N_3844,In_154,In_936);
or U3845 (N_3845,In_571,In_785);
and U3846 (N_3846,In_230,In_363);
nor U3847 (N_3847,In_145,In_890);
or U3848 (N_3848,In_973,In_867);
nor U3849 (N_3849,In_470,In_999);
nand U3850 (N_3850,In_685,In_534);
and U3851 (N_3851,In_899,In_339);
nor U3852 (N_3852,In_858,In_116);
nand U3853 (N_3853,In_92,In_506);
nor U3854 (N_3854,In_756,In_515);
or U3855 (N_3855,In_197,In_366);
nand U3856 (N_3856,In_917,In_565);
xor U3857 (N_3857,In_965,In_958);
nor U3858 (N_3858,In_263,In_119);
or U3859 (N_3859,In_106,In_454);
and U3860 (N_3860,In_400,In_252);
or U3861 (N_3861,In_259,In_318);
xor U3862 (N_3862,In_570,In_796);
or U3863 (N_3863,In_893,In_81);
nand U3864 (N_3864,In_831,In_757);
or U3865 (N_3865,In_852,In_368);
and U3866 (N_3866,In_443,In_630);
nor U3867 (N_3867,In_708,In_608);
nand U3868 (N_3868,In_840,In_948);
nand U3869 (N_3869,In_400,In_537);
nand U3870 (N_3870,In_78,In_769);
and U3871 (N_3871,In_249,In_336);
nand U3872 (N_3872,In_401,In_393);
or U3873 (N_3873,In_429,In_752);
or U3874 (N_3874,In_865,In_693);
nor U3875 (N_3875,In_467,In_877);
or U3876 (N_3876,In_37,In_465);
nor U3877 (N_3877,In_726,In_592);
nor U3878 (N_3878,In_884,In_887);
nor U3879 (N_3879,In_400,In_163);
and U3880 (N_3880,In_804,In_639);
nor U3881 (N_3881,In_625,In_413);
nor U3882 (N_3882,In_67,In_975);
or U3883 (N_3883,In_194,In_831);
and U3884 (N_3884,In_555,In_466);
nor U3885 (N_3885,In_470,In_317);
and U3886 (N_3886,In_549,In_827);
or U3887 (N_3887,In_238,In_625);
and U3888 (N_3888,In_84,In_467);
nand U3889 (N_3889,In_344,In_25);
nand U3890 (N_3890,In_14,In_511);
or U3891 (N_3891,In_832,In_46);
and U3892 (N_3892,In_490,In_293);
and U3893 (N_3893,In_742,In_15);
xor U3894 (N_3894,In_282,In_970);
or U3895 (N_3895,In_583,In_610);
nand U3896 (N_3896,In_944,In_28);
xnor U3897 (N_3897,In_538,In_19);
nand U3898 (N_3898,In_311,In_494);
or U3899 (N_3899,In_408,In_831);
or U3900 (N_3900,In_870,In_915);
nand U3901 (N_3901,In_228,In_766);
nand U3902 (N_3902,In_838,In_812);
nand U3903 (N_3903,In_876,In_105);
nand U3904 (N_3904,In_504,In_198);
nor U3905 (N_3905,In_481,In_606);
nand U3906 (N_3906,In_719,In_644);
and U3907 (N_3907,In_998,In_597);
and U3908 (N_3908,In_112,In_739);
nand U3909 (N_3909,In_38,In_555);
xor U3910 (N_3910,In_114,In_890);
xor U3911 (N_3911,In_281,In_187);
and U3912 (N_3912,In_843,In_279);
xor U3913 (N_3913,In_679,In_113);
xnor U3914 (N_3914,In_55,In_196);
xor U3915 (N_3915,In_525,In_530);
nor U3916 (N_3916,In_177,In_693);
nor U3917 (N_3917,In_732,In_871);
nor U3918 (N_3918,In_437,In_367);
nor U3919 (N_3919,In_437,In_344);
or U3920 (N_3920,In_879,In_316);
nor U3921 (N_3921,In_886,In_130);
nand U3922 (N_3922,In_635,In_304);
xor U3923 (N_3923,In_662,In_829);
nor U3924 (N_3924,In_131,In_312);
or U3925 (N_3925,In_406,In_160);
nor U3926 (N_3926,In_36,In_442);
or U3927 (N_3927,In_312,In_713);
or U3928 (N_3928,In_386,In_870);
and U3929 (N_3929,In_636,In_166);
nand U3930 (N_3930,In_815,In_3);
or U3931 (N_3931,In_452,In_763);
nor U3932 (N_3932,In_69,In_49);
nor U3933 (N_3933,In_838,In_848);
and U3934 (N_3934,In_247,In_459);
nor U3935 (N_3935,In_792,In_689);
and U3936 (N_3936,In_406,In_552);
or U3937 (N_3937,In_179,In_638);
nand U3938 (N_3938,In_294,In_845);
or U3939 (N_3939,In_378,In_416);
xor U3940 (N_3940,In_324,In_542);
nand U3941 (N_3941,In_173,In_64);
or U3942 (N_3942,In_760,In_57);
nand U3943 (N_3943,In_145,In_151);
nor U3944 (N_3944,In_942,In_790);
nand U3945 (N_3945,In_83,In_165);
and U3946 (N_3946,In_391,In_884);
xnor U3947 (N_3947,In_615,In_244);
and U3948 (N_3948,In_314,In_439);
or U3949 (N_3949,In_58,In_101);
nand U3950 (N_3950,In_196,In_883);
nor U3951 (N_3951,In_996,In_292);
nor U3952 (N_3952,In_423,In_384);
or U3953 (N_3953,In_43,In_833);
or U3954 (N_3954,In_539,In_15);
nand U3955 (N_3955,In_576,In_932);
or U3956 (N_3956,In_986,In_157);
or U3957 (N_3957,In_4,In_660);
and U3958 (N_3958,In_625,In_292);
and U3959 (N_3959,In_197,In_265);
or U3960 (N_3960,In_522,In_100);
or U3961 (N_3961,In_987,In_362);
and U3962 (N_3962,In_104,In_708);
nor U3963 (N_3963,In_42,In_608);
xor U3964 (N_3964,In_690,In_721);
nand U3965 (N_3965,In_244,In_982);
nand U3966 (N_3966,In_926,In_742);
xor U3967 (N_3967,In_891,In_454);
or U3968 (N_3968,In_595,In_23);
nand U3969 (N_3969,In_574,In_715);
xor U3970 (N_3970,In_628,In_295);
nor U3971 (N_3971,In_866,In_876);
or U3972 (N_3972,In_272,In_158);
nor U3973 (N_3973,In_325,In_589);
or U3974 (N_3974,In_807,In_535);
or U3975 (N_3975,In_699,In_119);
nand U3976 (N_3976,In_842,In_832);
and U3977 (N_3977,In_11,In_34);
xor U3978 (N_3978,In_307,In_128);
nor U3979 (N_3979,In_624,In_836);
or U3980 (N_3980,In_709,In_42);
nor U3981 (N_3981,In_341,In_216);
nand U3982 (N_3982,In_539,In_799);
or U3983 (N_3983,In_725,In_24);
and U3984 (N_3984,In_380,In_607);
nand U3985 (N_3985,In_311,In_968);
nor U3986 (N_3986,In_410,In_308);
nor U3987 (N_3987,In_744,In_35);
and U3988 (N_3988,In_0,In_339);
or U3989 (N_3989,In_43,In_421);
nand U3990 (N_3990,In_369,In_462);
and U3991 (N_3991,In_705,In_297);
xnor U3992 (N_3992,In_959,In_318);
and U3993 (N_3993,In_289,In_868);
nor U3994 (N_3994,In_902,In_84);
xnor U3995 (N_3995,In_603,In_275);
nand U3996 (N_3996,In_822,In_615);
nor U3997 (N_3997,In_613,In_6);
nor U3998 (N_3998,In_899,In_262);
nand U3999 (N_3999,In_133,In_38);
nand U4000 (N_4000,In_874,In_639);
nand U4001 (N_4001,In_146,In_424);
nor U4002 (N_4002,In_217,In_118);
nand U4003 (N_4003,In_552,In_635);
or U4004 (N_4004,In_936,In_47);
nand U4005 (N_4005,In_730,In_910);
nand U4006 (N_4006,In_37,In_444);
xnor U4007 (N_4007,In_802,In_24);
and U4008 (N_4008,In_305,In_642);
nor U4009 (N_4009,In_306,In_293);
nor U4010 (N_4010,In_912,In_142);
and U4011 (N_4011,In_625,In_165);
or U4012 (N_4012,In_480,In_718);
or U4013 (N_4013,In_181,In_325);
and U4014 (N_4014,In_614,In_696);
nor U4015 (N_4015,In_868,In_907);
or U4016 (N_4016,In_686,In_755);
and U4017 (N_4017,In_298,In_53);
nor U4018 (N_4018,In_973,In_345);
nand U4019 (N_4019,In_664,In_180);
and U4020 (N_4020,In_713,In_650);
nand U4021 (N_4021,In_751,In_402);
nand U4022 (N_4022,In_554,In_992);
xnor U4023 (N_4023,In_308,In_583);
and U4024 (N_4024,In_93,In_410);
and U4025 (N_4025,In_588,In_545);
nand U4026 (N_4026,In_717,In_918);
or U4027 (N_4027,In_422,In_483);
or U4028 (N_4028,In_651,In_835);
and U4029 (N_4029,In_592,In_440);
xor U4030 (N_4030,In_743,In_115);
or U4031 (N_4031,In_380,In_33);
or U4032 (N_4032,In_463,In_543);
or U4033 (N_4033,In_143,In_932);
and U4034 (N_4034,In_482,In_544);
and U4035 (N_4035,In_751,In_469);
nor U4036 (N_4036,In_502,In_814);
or U4037 (N_4037,In_481,In_954);
nand U4038 (N_4038,In_53,In_760);
nand U4039 (N_4039,In_114,In_167);
nand U4040 (N_4040,In_119,In_701);
or U4041 (N_4041,In_365,In_488);
nor U4042 (N_4042,In_428,In_745);
nand U4043 (N_4043,In_187,In_538);
and U4044 (N_4044,In_430,In_185);
nand U4045 (N_4045,In_191,In_800);
nor U4046 (N_4046,In_173,In_517);
nand U4047 (N_4047,In_788,In_732);
or U4048 (N_4048,In_330,In_663);
nand U4049 (N_4049,In_172,In_409);
nor U4050 (N_4050,In_628,In_282);
nor U4051 (N_4051,In_851,In_799);
or U4052 (N_4052,In_910,In_391);
nand U4053 (N_4053,In_146,In_535);
nor U4054 (N_4054,In_182,In_570);
and U4055 (N_4055,In_586,In_565);
nand U4056 (N_4056,In_970,In_491);
or U4057 (N_4057,In_334,In_209);
or U4058 (N_4058,In_8,In_119);
nand U4059 (N_4059,In_248,In_809);
nor U4060 (N_4060,In_644,In_931);
xnor U4061 (N_4061,In_288,In_276);
and U4062 (N_4062,In_336,In_302);
nor U4063 (N_4063,In_297,In_589);
nand U4064 (N_4064,In_73,In_412);
nor U4065 (N_4065,In_699,In_306);
nand U4066 (N_4066,In_641,In_658);
and U4067 (N_4067,In_530,In_235);
nor U4068 (N_4068,In_788,In_334);
and U4069 (N_4069,In_217,In_810);
nand U4070 (N_4070,In_654,In_553);
nand U4071 (N_4071,In_685,In_969);
and U4072 (N_4072,In_751,In_868);
and U4073 (N_4073,In_358,In_407);
xor U4074 (N_4074,In_769,In_515);
nand U4075 (N_4075,In_269,In_109);
nor U4076 (N_4076,In_943,In_86);
or U4077 (N_4077,In_559,In_764);
nor U4078 (N_4078,In_198,In_271);
or U4079 (N_4079,In_813,In_486);
xnor U4080 (N_4080,In_293,In_554);
xnor U4081 (N_4081,In_308,In_910);
or U4082 (N_4082,In_874,In_80);
nand U4083 (N_4083,In_674,In_434);
and U4084 (N_4084,In_806,In_180);
nor U4085 (N_4085,In_924,In_330);
or U4086 (N_4086,In_689,In_665);
nor U4087 (N_4087,In_419,In_294);
nand U4088 (N_4088,In_462,In_815);
and U4089 (N_4089,In_601,In_206);
and U4090 (N_4090,In_252,In_187);
or U4091 (N_4091,In_779,In_650);
nand U4092 (N_4092,In_378,In_855);
xor U4093 (N_4093,In_130,In_901);
nand U4094 (N_4094,In_249,In_738);
nor U4095 (N_4095,In_284,In_298);
nor U4096 (N_4096,In_856,In_210);
nor U4097 (N_4097,In_645,In_866);
nor U4098 (N_4098,In_830,In_458);
or U4099 (N_4099,In_648,In_771);
nor U4100 (N_4100,In_73,In_612);
nor U4101 (N_4101,In_571,In_37);
or U4102 (N_4102,In_619,In_260);
and U4103 (N_4103,In_722,In_808);
or U4104 (N_4104,In_402,In_719);
and U4105 (N_4105,In_875,In_74);
or U4106 (N_4106,In_243,In_602);
nor U4107 (N_4107,In_151,In_381);
xnor U4108 (N_4108,In_322,In_790);
xnor U4109 (N_4109,In_654,In_959);
nand U4110 (N_4110,In_725,In_97);
or U4111 (N_4111,In_110,In_170);
nand U4112 (N_4112,In_85,In_383);
nand U4113 (N_4113,In_336,In_475);
and U4114 (N_4114,In_960,In_257);
and U4115 (N_4115,In_31,In_417);
nor U4116 (N_4116,In_957,In_445);
or U4117 (N_4117,In_473,In_924);
or U4118 (N_4118,In_286,In_391);
or U4119 (N_4119,In_31,In_205);
nor U4120 (N_4120,In_741,In_296);
and U4121 (N_4121,In_869,In_124);
and U4122 (N_4122,In_495,In_799);
and U4123 (N_4123,In_226,In_241);
or U4124 (N_4124,In_659,In_498);
nand U4125 (N_4125,In_277,In_312);
xnor U4126 (N_4126,In_516,In_943);
and U4127 (N_4127,In_750,In_217);
nor U4128 (N_4128,In_849,In_8);
nor U4129 (N_4129,In_890,In_185);
or U4130 (N_4130,In_307,In_477);
nor U4131 (N_4131,In_589,In_41);
or U4132 (N_4132,In_33,In_175);
nand U4133 (N_4133,In_807,In_54);
nand U4134 (N_4134,In_692,In_212);
xnor U4135 (N_4135,In_989,In_441);
and U4136 (N_4136,In_727,In_740);
and U4137 (N_4137,In_443,In_120);
xor U4138 (N_4138,In_380,In_305);
or U4139 (N_4139,In_873,In_99);
and U4140 (N_4140,In_446,In_815);
nand U4141 (N_4141,In_209,In_496);
and U4142 (N_4142,In_803,In_641);
or U4143 (N_4143,In_925,In_127);
nand U4144 (N_4144,In_929,In_505);
nand U4145 (N_4145,In_230,In_937);
nor U4146 (N_4146,In_877,In_124);
and U4147 (N_4147,In_442,In_883);
nor U4148 (N_4148,In_216,In_761);
and U4149 (N_4149,In_455,In_898);
and U4150 (N_4150,In_873,In_255);
or U4151 (N_4151,In_969,In_806);
nor U4152 (N_4152,In_475,In_905);
nor U4153 (N_4153,In_720,In_110);
xnor U4154 (N_4154,In_613,In_320);
nor U4155 (N_4155,In_86,In_576);
nor U4156 (N_4156,In_555,In_942);
and U4157 (N_4157,In_423,In_199);
nor U4158 (N_4158,In_513,In_98);
or U4159 (N_4159,In_983,In_136);
nor U4160 (N_4160,In_203,In_149);
or U4161 (N_4161,In_606,In_641);
nor U4162 (N_4162,In_86,In_795);
xnor U4163 (N_4163,In_376,In_407);
nand U4164 (N_4164,In_686,In_761);
nand U4165 (N_4165,In_819,In_499);
nor U4166 (N_4166,In_962,In_64);
xor U4167 (N_4167,In_31,In_749);
nor U4168 (N_4168,In_407,In_30);
nor U4169 (N_4169,In_524,In_33);
nand U4170 (N_4170,In_898,In_841);
or U4171 (N_4171,In_673,In_489);
and U4172 (N_4172,In_957,In_597);
nand U4173 (N_4173,In_186,In_590);
or U4174 (N_4174,In_77,In_566);
nand U4175 (N_4175,In_333,In_547);
or U4176 (N_4176,In_438,In_630);
and U4177 (N_4177,In_56,In_487);
nor U4178 (N_4178,In_39,In_779);
or U4179 (N_4179,In_846,In_826);
and U4180 (N_4180,In_367,In_867);
and U4181 (N_4181,In_546,In_437);
or U4182 (N_4182,In_948,In_965);
or U4183 (N_4183,In_586,In_923);
or U4184 (N_4184,In_632,In_168);
or U4185 (N_4185,In_979,In_20);
xnor U4186 (N_4186,In_395,In_109);
nand U4187 (N_4187,In_696,In_340);
nand U4188 (N_4188,In_565,In_828);
nor U4189 (N_4189,In_335,In_912);
or U4190 (N_4190,In_144,In_61);
nor U4191 (N_4191,In_776,In_663);
nor U4192 (N_4192,In_622,In_323);
and U4193 (N_4193,In_729,In_968);
or U4194 (N_4194,In_401,In_885);
xor U4195 (N_4195,In_681,In_280);
or U4196 (N_4196,In_867,In_300);
or U4197 (N_4197,In_424,In_691);
nand U4198 (N_4198,In_879,In_658);
nor U4199 (N_4199,In_881,In_439);
or U4200 (N_4200,In_290,In_101);
xnor U4201 (N_4201,In_996,In_828);
or U4202 (N_4202,In_855,In_319);
or U4203 (N_4203,In_239,In_925);
and U4204 (N_4204,In_172,In_833);
and U4205 (N_4205,In_467,In_585);
or U4206 (N_4206,In_563,In_594);
and U4207 (N_4207,In_149,In_159);
and U4208 (N_4208,In_979,In_114);
or U4209 (N_4209,In_790,In_345);
xor U4210 (N_4210,In_414,In_68);
or U4211 (N_4211,In_528,In_245);
and U4212 (N_4212,In_323,In_90);
nand U4213 (N_4213,In_440,In_698);
and U4214 (N_4214,In_576,In_768);
or U4215 (N_4215,In_387,In_97);
nor U4216 (N_4216,In_901,In_74);
xor U4217 (N_4217,In_787,In_165);
nand U4218 (N_4218,In_139,In_729);
xor U4219 (N_4219,In_616,In_304);
nand U4220 (N_4220,In_413,In_713);
nor U4221 (N_4221,In_842,In_652);
nand U4222 (N_4222,In_980,In_847);
nor U4223 (N_4223,In_943,In_496);
and U4224 (N_4224,In_334,In_876);
xnor U4225 (N_4225,In_8,In_250);
nand U4226 (N_4226,In_84,In_307);
and U4227 (N_4227,In_933,In_380);
nor U4228 (N_4228,In_3,In_217);
nor U4229 (N_4229,In_764,In_725);
nand U4230 (N_4230,In_13,In_950);
nor U4231 (N_4231,In_260,In_519);
nand U4232 (N_4232,In_523,In_704);
nor U4233 (N_4233,In_87,In_215);
xor U4234 (N_4234,In_821,In_747);
nor U4235 (N_4235,In_877,In_131);
nor U4236 (N_4236,In_804,In_558);
or U4237 (N_4237,In_375,In_712);
or U4238 (N_4238,In_286,In_850);
nand U4239 (N_4239,In_135,In_632);
and U4240 (N_4240,In_176,In_283);
nor U4241 (N_4241,In_206,In_459);
nand U4242 (N_4242,In_392,In_938);
or U4243 (N_4243,In_798,In_485);
and U4244 (N_4244,In_230,In_588);
and U4245 (N_4245,In_254,In_658);
nand U4246 (N_4246,In_233,In_405);
nand U4247 (N_4247,In_209,In_383);
or U4248 (N_4248,In_357,In_878);
or U4249 (N_4249,In_329,In_811);
or U4250 (N_4250,In_427,In_589);
nand U4251 (N_4251,In_92,In_598);
xor U4252 (N_4252,In_873,In_170);
xnor U4253 (N_4253,In_267,In_166);
or U4254 (N_4254,In_531,In_772);
and U4255 (N_4255,In_416,In_134);
or U4256 (N_4256,In_67,In_54);
nor U4257 (N_4257,In_723,In_179);
or U4258 (N_4258,In_701,In_728);
or U4259 (N_4259,In_630,In_232);
and U4260 (N_4260,In_295,In_833);
nand U4261 (N_4261,In_433,In_471);
nand U4262 (N_4262,In_5,In_750);
nand U4263 (N_4263,In_509,In_626);
nand U4264 (N_4264,In_70,In_879);
nand U4265 (N_4265,In_36,In_20);
nand U4266 (N_4266,In_630,In_858);
or U4267 (N_4267,In_564,In_973);
nor U4268 (N_4268,In_820,In_835);
and U4269 (N_4269,In_708,In_932);
or U4270 (N_4270,In_672,In_225);
nor U4271 (N_4271,In_74,In_351);
or U4272 (N_4272,In_816,In_769);
nor U4273 (N_4273,In_267,In_450);
or U4274 (N_4274,In_217,In_89);
nor U4275 (N_4275,In_640,In_624);
nor U4276 (N_4276,In_836,In_985);
xor U4277 (N_4277,In_413,In_242);
nor U4278 (N_4278,In_547,In_499);
nor U4279 (N_4279,In_196,In_79);
nand U4280 (N_4280,In_142,In_414);
or U4281 (N_4281,In_449,In_724);
and U4282 (N_4282,In_713,In_325);
nand U4283 (N_4283,In_207,In_815);
or U4284 (N_4284,In_73,In_458);
nand U4285 (N_4285,In_453,In_662);
and U4286 (N_4286,In_739,In_517);
and U4287 (N_4287,In_848,In_525);
or U4288 (N_4288,In_16,In_203);
or U4289 (N_4289,In_46,In_897);
nand U4290 (N_4290,In_459,In_894);
and U4291 (N_4291,In_844,In_363);
xnor U4292 (N_4292,In_820,In_36);
nand U4293 (N_4293,In_746,In_540);
nand U4294 (N_4294,In_402,In_604);
xor U4295 (N_4295,In_522,In_769);
nand U4296 (N_4296,In_95,In_743);
nand U4297 (N_4297,In_646,In_258);
nor U4298 (N_4298,In_753,In_969);
nor U4299 (N_4299,In_636,In_116);
or U4300 (N_4300,In_782,In_266);
and U4301 (N_4301,In_988,In_119);
nor U4302 (N_4302,In_4,In_932);
nor U4303 (N_4303,In_104,In_275);
nor U4304 (N_4304,In_759,In_282);
nand U4305 (N_4305,In_38,In_247);
nor U4306 (N_4306,In_988,In_361);
nor U4307 (N_4307,In_91,In_519);
and U4308 (N_4308,In_226,In_781);
nor U4309 (N_4309,In_189,In_387);
xnor U4310 (N_4310,In_191,In_478);
nand U4311 (N_4311,In_657,In_113);
nor U4312 (N_4312,In_882,In_557);
nor U4313 (N_4313,In_849,In_567);
nor U4314 (N_4314,In_53,In_97);
or U4315 (N_4315,In_635,In_168);
xor U4316 (N_4316,In_573,In_45);
or U4317 (N_4317,In_535,In_750);
and U4318 (N_4318,In_767,In_991);
or U4319 (N_4319,In_211,In_148);
and U4320 (N_4320,In_783,In_397);
nand U4321 (N_4321,In_875,In_621);
nand U4322 (N_4322,In_574,In_412);
nor U4323 (N_4323,In_476,In_789);
and U4324 (N_4324,In_745,In_727);
nand U4325 (N_4325,In_569,In_624);
and U4326 (N_4326,In_77,In_868);
and U4327 (N_4327,In_140,In_696);
or U4328 (N_4328,In_719,In_169);
xnor U4329 (N_4329,In_601,In_998);
nand U4330 (N_4330,In_359,In_300);
nor U4331 (N_4331,In_143,In_756);
or U4332 (N_4332,In_374,In_354);
nand U4333 (N_4333,In_818,In_390);
and U4334 (N_4334,In_952,In_681);
or U4335 (N_4335,In_568,In_385);
nand U4336 (N_4336,In_375,In_178);
and U4337 (N_4337,In_297,In_365);
nor U4338 (N_4338,In_276,In_175);
nand U4339 (N_4339,In_775,In_602);
nor U4340 (N_4340,In_428,In_15);
xnor U4341 (N_4341,In_704,In_605);
nand U4342 (N_4342,In_424,In_166);
nand U4343 (N_4343,In_422,In_64);
nor U4344 (N_4344,In_200,In_500);
or U4345 (N_4345,In_503,In_533);
nor U4346 (N_4346,In_383,In_357);
nand U4347 (N_4347,In_816,In_474);
or U4348 (N_4348,In_579,In_639);
or U4349 (N_4349,In_464,In_213);
nand U4350 (N_4350,In_489,In_801);
and U4351 (N_4351,In_289,In_918);
or U4352 (N_4352,In_490,In_444);
or U4353 (N_4353,In_205,In_414);
or U4354 (N_4354,In_992,In_212);
and U4355 (N_4355,In_441,In_277);
nand U4356 (N_4356,In_770,In_539);
or U4357 (N_4357,In_643,In_701);
nand U4358 (N_4358,In_936,In_612);
xnor U4359 (N_4359,In_638,In_345);
or U4360 (N_4360,In_923,In_513);
and U4361 (N_4361,In_596,In_722);
or U4362 (N_4362,In_465,In_3);
and U4363 (N_4363,In_595,In_443);
nor U4364 (N_4364,In_804,In_213);
nand U4365 (N_4365,In_230,In_392);
nand U4366 (N_4366,In_842,In_418);
and U4367 (N_4367,In_45,In_823);
nor U4368 (N_4368,In_304,In_853);
or U4369 (N_4369,In_143,In_814);
and U4370 (N_4370,In_488,In_844);
or U4371 (N_4371,In_263,In_878);
nor U4372 (N_4372,In_869,In_463);
nand U4373 (N_4373,In_15,In_875);
xor U4374 (N_4374,In_130,In_25);
nor U4375 (N_4375,In_962,In_129);
nor U4376 (N_4376,In_650,In_422);
xor U4377 (N_4377,In_56,In_687);
or U4378 (N_4378,In_648,In_893);
nand U4379 (N_4379,In_83,In_426);
nor U4380 (N_4380,In_386,In_142);
nor U4381 (N_4381,In_732,In_332);
and U4382 (N_4382,In_836,In_599);
xor U4383 (N_4383,In_522,In_180);
or U4384 (N_4384,In_727,In_863);
or U4385 (N_4385,In_51,In_534);
nand U4386 (N_4386,In_92,In_236);
or U4387 (N_4387,In_829,In_875);
and U4388 (N_4388,In_40,In_15);
and U4389 (N_4389,In_390,In_203);
or U4390 (N_4390,In_116,In_795);
or U4391 (N_4391,In_566,In_112);
nor U4392 (N_4392,In_457,In_695);
or U4393 (N_4393,In_550,In_202);
nor U4394 (N_4394,In_434,In_749);
nand U4395 (N_4395,In_230,In_618);
nand U4396 (N_4396,In_361,In_469);
nand U4397 (N_4397,In_3,In_876);
nor U4398 (N_4398,In_540,In_993);
or U4399 (N_4399,In_487,In_691);
nor U4400 (N_4400,In_751,In_328);
or U4401 (N_4401,In_64,In_519);
nor U4402 (N_4402,In_839,In_686);
and U4403 (N_4403,In_858,In_836);
nand U4404 (N_4404,In_76,In_463);
nand U4405 (N_4405,In_264,In_130);
nor U4406 (N_4406,In_784,In_683);
nor U4407 (N_4407,In_438,In_463);
nand U4408 (N_4408,In_737,In_505);
xnor U4409 (N_4409,In_884,In_826);
nand U4410 (N_4410,In_704,In_744);
or U4411 (N_4411,In_272,In_517);
or U4412 (N_4412,In_783,In_227);
or U4413 (N_4413,In_846,In_709);
or U4414 (N_4414,In_685,In_473);
and U4415 (N_4415,In_545,In_387);
nor U4416 (N_4416,In_418,In_63);
and U4417 (N_4417,In_637,In_762);
or U4418 (N_4418,In_873,In_158);
and U4419 (N_4419,In_516,In_823);
or U4420 (N_4420,In_714,In_934);
and U4421 (N_4421,In_153,In_801);
nor U4422 (N_4422,In_30,In_968);
and U4423 (N_4423,In_602,In_219);
nand U4424 (N_4424,In_269,In_455);
nand U4425 (N_4425,In_149,In_679);
xnor U4426 (N_4426,In_312,In_370);
nand U4427 (N_4427,In_241,In_275);
nand U4428 (N_4428,In_302,In_646);
nand U4429 (N_4429,In_125,In_150);
and U4430 (N_4430,In_168,In_571);
or U4431 (N_4431,In_927,In_319);
and U4432 (N_4432,In_269,In_372);
or U4433 (N_4433,In_338,In_858);
and U4434 (N_4434,In_175,In_167);
and U4435 (N_4435,In_681,In_422);
nand U4436 (N_4436,In_899,In_412);
nor U4437 (N_4437,In_158,In_538);
and U4438 (N_4438,In_34,In_642);
or U4439 (N_4439,In_201,In_385);
nor U4440 (N_4440,In_358,In_768);
and U4441 (N_4441,In_170,In_596);
and U4442 (N_4442,In_312,In_964);
or U4443 (N_4443,In_311,In_97);
and U4444 (N_4444,In_568,In_891);
nand U4445 (N_4445,In_950,In_292);
xnor U4446 (N_4446,In_508,In_67);
nor U4447 (N_4447,In_259,In_711);
or U4448 (N_4448,In_755,In_150);
and U4449 (N_4449,In_858,In_801);
or U4450 (N_4450,In_76,In_470);
or U4451 (N_4451,In_130,In_461);
nor U4452 (N_4452,In_875,In_277);
nand U4453 (N_4453,In_377,In_384);
or U4454 (N_4454,In_230,In_336);
xnor U4455 (N_4455,In_286,In_537);
nand U4456 (N_4456,In_190,In_662);
or U4457 (N_4457,In_84,In_393);
and U4458 (N_4458,In_209,In_656);
nand U4459 (N_4459,In_42,In_933);
xor U4460 (N_4460,In_394,In_274);
or U4461 (N_4461,In_834,In_560);
nor U4462 (N_4462,In_207,In_916);
nor U4463 (N_4463,In_24,In_609);
nand U4464 (N_4464,In_41,In_182);
or U4465 (N_4465,In_423,In_571);
nand U4466 (N_4466,In_686,In_375);
xor U4467 (N_4467,In_648,In_978);
xnor U4468 (N_4468,In_874,In_614);
nor U4469 (N_4469,In_640,In_977);
xor U4470 (N_4470,In_627,In_201);
nand U4471 (N_4471,In_709,In_647);
nor U4472 (N_4472,In_557,In_778);
or U4473 (N_4473,In_86,In_656);
or U4474 (N_4474,In_374,In_334);
or U4475 (N_4475,In_574,In_970);
nand U4476 (N_4476,In_884,In_813);
nor U4477 (N_4477,In_105,In_550);
nor U4478 (N_4478,In_841,In_856);
nor U4479 (N_4479,In_997,In_550);
and U4480 (N_4480,In_252,In_739);
and U4481 (N_4481,In_579,In_596);
and U4482 (N_4482,In_212,In_724);
and U4483 (N_4483,In_678,In_446);
nor U4484 (N_4484,In_902,In_937);
or U4485 (N_4485,In_575,In_557);
nand U4486 (N_4486,In_813,In_36);
nand U4487 (N_4487,In_568,In_0);
or U4488 (N_4488,In_840,In_521);
and U4489 (N_4489,In_941,In_359);
xnor U4490 (N_4490,In_298,In_562);
nand U4491 (N_4491,In_729,In_324);
or U4492 (N_4492,In_343,In_371);
and U4493 (N_4493,In_456,In_149);
or U4494 (N_4494,In_58,In_164);
nor U4495 (N_4495,In_934,In_756);
and U4496 (N_4496,In_439,In_132);
or U4497 (N_4497,In_108,In_936);
nor U4498 (N_4498,In_907,In_265);
nand U4499 (N_4499,In_722,In_298);
nand U4500 (N_4500,In_709,In_276);
nor U4501 (N_4501,In_82,In_151);
nor U4502 (N_4502,In_952,In_754);
or U4503 (N_4503,In_339,In_799);
and U4504 (N_4504,In_124,In_272);
nor U4505 (N_4505,In_21,In_602);
nor U4506 (N_4506,In_154,In_139);
and U4507 (N_4507,In_178,In_109);
xnor U4508 (N_4508,In_86,In_594);
or U4509 (N_4509,In_23,In_188);
and U4510 (N_4510,In_434,In_677);
nand U4511 (N_4511,In_279,In_449);
and U4512 (N_4512,In_561,In_706);
nor U4513 (N_4513,In_148,In_549);
nor U4514 (N_4514,In_179,In_70);
or U4515 (N_4515,In_359,In_229);
nor U4516 (N_4516,In_520,In_938);
or U4517 (N_4517,In_256,In_297);
nor U4518 (N_4518,In_380,In_952);
or U4519 (N_4519,In_203,In_490);
nor U4520 (N_4520,In_183,In_161);
nor U4521 (N_4521,In_997,In_814);
or U4522 (N_4522,In_177,In_81);
and U4523 (N_4523,In_450,In_674);
and U4524 (N_4524,In_925,In_72);
nor U4525 (N_4525,In_98,In_284);
and U4526 (N_4526,In_504,In_690);
and U4527 (N_4527,In_394,In_375);
nor U4528 (N_4528,In_817,In_619);
and U4529 (N_4529,In_599,In_732);
nand U4530 (N_4530,In_787,In_799);
nor U4531 (N_4531,In_434,In_98);
nand U4532 (N_4532,In_637,In_820);
nand U4533 (N_4533,In_938,In_538);
nor U4534 (N_4534,In_186,In_384);
nand U4535 (N_4535,In_503,In_207);
xnor U4536 (N_4536,In_303,In_398);
and U4537 (N_4537,In_531,In_780);
and U4538 (N_4538,In_584,In_71);
xor U4539 (N_4539,In_222,In_687);
and U4540 (N_4540,In_836,In_260);
nor U4541 (N_4541,In_358,In_476);
nor U4542 (N_4542,In_155,In_534);
nor U4543 (N_4543,In_653,In_819);
or U4544 (N_4544,In_508,In_725);
or U4545 (N_4545,In_503,In_650);
and U4546 (N_4546,In_153,In_418);
or U4547 (N_4547,In_881,In_183);
nor U4548 (N_4548,In_212,In_442);
and U4549 (N_4549,In_487,In_163);
or U4550 (N_4550,In_992,In_493);
xor U4551 (N_4551,In_342,In_325);
nor U4552 (N_4552,In_289,In_200);
xnor U4553 (N_4553,In_904,In_813);
or U4554 (N_4554,In_948,In_11);
xnor U4555 (N_4555,In_301,In_25);
or U4556 (N_4556,In_425,In_621);
nand U4557 (N_4557,In_719,In_245);
xnor U4558 (N_4558,In_986,In_42);
nand U4559 (N_4559,In_122,In_284);
and U4560 (N_4560,In_665,In_89);
nor U4561 (N_4561,In_622,In_122);
and U4562 (N_4562,In_878,In_43);
nand U4563 (N_4563,In_366,In_502);
nand U4564 (N_4564,In_750,In_76);
nand U4565 (N_4565,In_938,In_760);
or U4566 (N_4566,In_549,In_380);
and U4567 (N_4567,In_266,In_130);
xnor U4568 (N_4568,In_839,In_598);
xor U4569 (N_4569,In_593,In_758);
nand U4570 (N_4570,In_412,In_323);
nor U4571 (N_4571,In_990,In_464);
and U4572 (N_4572,In_600,In_486);
nor U4573 (N_4573,In_142,In_57);
nor U4574 (N_4574,In_151,In_218);
or U4575 (N_4575,In_185,In_930);
xor U4576 (N_4576,In_592,In_443);
xnor U4577 (N_4577,In_297,In_970);
nand U4578 (N_4578,In_525,In_169);
nand U4579 (N_4579,In_388,In_273);
or U4580 (N_4580,In_789,In_450);
or U4581 (N_4581,In_259,In_142);
nor U4582 (N_4582,In_644,In_485);
and U4583 (N_4583,In_191,In_453);
nand U4584 (N_4584,In_639,In_366);
or U4585 (N_4585,In_708,In_376);
xnor U4586 (N_4586,In_75,In_190);
and U4587 (N_4587,In_89,In_289);
or U4588 (N_4588,In_71,In_378);
nand U4589 (N_4589,In_266,In_3);
nor U4590 (N_4590,In_396,In_686);
or U4591 (N_4591,In_332,In_942);
and U4592 (N_4592,In_611,In_186);
nand U4593 (N_4593,In_194,In_701);
nand U4594 (N_4594,In_275,In_139);
and U4595 (N_4595,In_555,In_644);
and U4596 (N_4596,In_236,In_704);
nor U4597 (N_4597,In_294,In_33);
xnor U4598 (N_4598,In_339,In_744);
nor U4599 (N_4599,In_118,In_823);
nand U4600 (N_4600,In_327,In_717);
and U4601 (N_4601,In_315,In_944);
or U4602 (N_4602,In_746,In_803);
nor U4603 (N_4603,In_997,In_237);
nand U4604 (N_4604,In_526,In_542);
or U4605 (N_4605,In_859,In_774);
and U4606 (N_4606,In_38,In_869);
xor U4607 (N_4607,In_549,In_302);
and U4608 (N_4608,In_31,In_504);
nand U4609 (N_4609,In_154,In_679);
and U4610 (N_4610,In_979,In_139);
or U4611 (N_4611,In_118,In_967);
or U4612 (N_4612,In_674,In_989);
nand U4613 (N_4613,In_441,In_160);
nor U4614 (N_4614,In_763,In_287);
or U4615 (N_4615,In_306,In_9);
nand U4616 (N_4616,In_803,In_804);
xor U4617 (N_4617,In_230,In_527);
xor U4618 (N_4618,In_122,In_34);
and U4619 (N_4619,In_320,In_948);
nand U4620 (N_4620,In_21,In_858);
nand U4621 (N_4621,In_401,In_237);
nor U4622 (N_4622,In_724,In_772);
or U4623 (N_4623,In_466,In_215);
and U4624 (N_4624,In_900,In_261);
and U4625 (N_4625,In_248,In_382);
and U4626 (N_4626,In_311,In_198);
or U4627 (N_4627,In_704,In_79);
or U4628 (N_4628,In_700,In_148);
and U4629 (N_4629,In_489,In_240);
nand U4630 (N_4630,In_194,In_15);
nand U4631 (N_4631,In_839,In_150);
nor U4632 (N_4632,In_313,In_451);
nor U4633 (N_4633,In_965,In_733);
nor U4634 (N_4634,In_823,In_865);
nand U4635 (N_4635,In_813,In_119);
and U4636 (N_4636,In_583,In_449);
nor U4637 (N_4637,In_603,In_926);
nor U4638 (N_4638,In_93,In_531);
nand U4639 (N_4639,In_441,In_438);
and U4640 (N_4640,In_594,In_29);
xnor U4641 (N_4641,In_131,In_318);
nor U4642 (N_4642,In_504,In_971);
or U4643 (N_4643,In_644,In_336);
xnor U4644 (N_4644,In_758,In_148);
or U4645 (N_4645,In_771,In_635);
and U4646 (N_4646,In_483,In_348);
nand U4647 (N_4647,In_760,In_980);
nand U4648 (N_4648,In_782,In_624);
and U4649 (N_4649,In_356,In_164);
and U4650 (N_4650,In_404,In_916);
nand U4651 (N_4651,In_844,In_809);
and U4652 (N_4652,In_228,In_197);
or U4653 (N_4653,In_155,In_207);
xnor U4654 (N_4654,In_31,In_41);
nand U4655 (N_4655,In_810,In_804);
nor U4656 (N_4656,In_113,In_225);
nand U4657 (N_4657,In_249,In_794);
xor U4658 (N_4658,In_853,In_872);
and U4659 (N_4659,In_464,In_656);
nor U4660 (N_4660,In_656,In_313);
nor U4661 (N_4661,In_861,In_839);
and U4662 (N_4662,In_653,In_831);
nor U4663 (N_4663,In_305,In_400);
nor U4664 (N_4664,In_819,In_845);
or U4665 (N_4665,In_260,In_682);
nor U4666 (N_4666,In_893,In_456);
or U4667 (N_4667,In_446,In_10);
and U4668 (N_4668,In_686,In_419);
nand U4669 (N_4669,In_31,In_505);
nand U4670 (N_4670,In_329,In_339);
and U4671 (N_4671,In_784,In_487);
xnor U4672 (N_4672,In_971,In_83);
or U4673 (N_4673,In_636,In_243);
and U4674 (N_4674,In_672,In_525);
or U4675 (N_4675,In_693,In_605);
nand U4676 (N_4676,In_541,In_254);
and U4677 (N_4677,In_796,In_807);
or U4678 (N_4678,In_153,In_863);
xor U4679 (N_4679,In_560,In_852);
nor U4680 (N_4680,In_652,In_249);
and U4681 (N_4681,In_414,In_720);
nand U4682 (N_4682,In_960,In_983);
nor U4683 (N_4683,In_187,In_50);
nor U4684 (N_4684,In_344,In_583);
nand U4685 (N_4685,In_689,In_226);
and U4686 (N_4686,In_650,In_912);
and U4687 (N_4687,In_733,In_425);
nand U4688 (N_4688,In_234,In_22);
xnor U4689 (N_4689,In_918,In_515);
nor U4690 (N_4690,In_662,In_442);
or U4691 (N_4691,In_824,In_795);
xor U4692 (N_4692,In_827,In_514);
or U4693 (N_4693,In_842,In_866);
or U4694 (N_4694,In_975,In_670);
nor U4695 (N_4695,In_277,In_598);
nor U4696 (N_4696,In_184,In_464);
nor U4697 (N_4697,In_834,In_245);
or U4698 (N_4698,In_829,In_795);
or U4699 (N_4699,In_445,In_178);
nand U4700 (N_4700,In_8,In_983);
xor U4701 (N_4701,In_447,In_168);
and U4702 (N_4702,In_649,In_581);
xnor U4703 (N_4703,In_485,In_453);
nand U4704 (N_4704,In_132,In_295);
and U4705 (N_4705,In_434,In_264);
nand U4706 (N_4706,In_361,In_961);
nand U4707 (N_4707,In_507,In_475);
and U4708 (N_4708,In_869,In_876);
nor U4709 (N_4709,In_380,In_908);
and U4710 (N_4710,In_829,In_729);
nor U4711 (N_4711,In_144,In_605);
or U4712 (N_4712,In_575,In_383);
nor U4713 (N_4713,In_748,In_627);
and U4714 (N_4714,In_680,In_308);
and U4715 (N_4715,In_0,In_747);
xnor U4716 (N_4716,In_810,In_485);
nor U4717 (N_4717,In_895,In_571);
xor U4718 (N_4718,In_374,In_827);
nand U4719 (N_4719,In_308,In_428);
and U4720 (N_4720,In_578,In_684);
or U4721 (N_4721,In_546,In_736);
nor U4722 (N_4722,In_747,In_864);
and U4723 (N_4723,In_100,In_618);
or U4724 (N_4724,In_705,In_593);
nor U4725 (N_4725,In_646,In_693);
and U4726 (N_4726,In_271,In_672);
xnor U4727 (N_4727,In_330,In_468);
xnor U4728 (N_4728,In_707,In_539);
xor U4729 (N_4729,In_217,In_953);
or U4730 (N_4730,In_435,In_152);
nand U4731 (N_4731,In_44,In_688);
nand U4732 (N_4732,In_901,In_197);
xor U4733 (N_4733,In_715,In_665);
and U4734 (N_4734,In_706,In_998);
or U4735 (N_4735,In_649,In_665);
xnor U4736 (N_4736,In_512,In_822);
nor U4737 (N_4737,In_565,In_303);
xor U4738 (N_4738,In_108,In_184);
or U4739 (N_4739,In_880,In_895);
and U4740 (N_4740,In_909,In_794);
and U4741 (N_4741,In_623,In_571);
nor U4742 (N_4742,In_347,In_424);
xor U4743 (N_4743,In_767,In_679);
or U4744 (N_4744,In_367,In_77);
or U4745 (N_4745,In_536,In_398);
and U4746 (N_4746,In_190,In_515);
or U4747 (N_4747,In_563,In_151);
nor U4748 (N_4748,In_900,In_662);
or U4749 (N_4749,In_10,In_179);
nor U4750 (N_4750,In_385,In_38);
nor U4751 (N_4751,In_154,In_38);
nand U4752 (N_4752,In_858,In_812);
or U4753 (N_4753,In_879,In_597);
nor U4754 (N_4754,In_24,In_261);
and U4755 (N_4755,In_735,In_437);
or U4756 (N_4756,In_4,In_160);
xnor U4757 (N_4757,In_199,In_58);
nand U4758 (N_4758,In_484,In_321);
nor U4759 (N_4759,In_813,In_497);
and U4760 (N_4760,In_659,In_270);
and U4761 (N_4761,In_999,In_359);
nand U4762 (N_4762,In_448,In_848);
nand U4763 (N_4763,In_836,In_395);
nor U4764 (N_4764,In_276,In_414);
nor U4765 (N_4765,In_263,In_132);
nor U4766 (N_4766,In_151,In_45);
nand U4767 (N_4767,In_234,In_76);
xor U4768 (N_4768,In_618,In_763);
nand U4769 (N_4769,In_816,In_960);
and U4770 (N_4770,In_201,In_694);
nand U4771 (N_4771,In_254,In_100);
or U4772 (N_4772,In_540,In_404);
or U4773 (N_4773,In_374,In_177);
and U4774 (N_4774,In_637,In_785);
and U4775 (N_4775,In_931,In_233);
and U4776 (N_4776,In_198,In_361);
and U4777 (N_4777,In_802,In_777);
xnor U4778 (N_4778,In_952,In_12);
nor U4779 (N_4779,In_322,In_222);
or U4780 (N_4780,In_194,In_227);
nor U4781 (N_4781,In_487,In_535);
nand U4782 (N_4782,In_278,In_69);
nand U4783 (N_4783,In_14,In_337);
nor U4784 (N_4784,In_337,In_247);
xnor U4785 (N_4785,In_232,In_556);
nand U4786 (N_4786,In_326,In_559);
nor U4787 (N_4787,In_620,In_917);
nor U4788 (N_4788,In_112,In_665);
nand U4789 (N_4789,In_238,In_719);
xnor U4790 (N_4790,In_684,In_718);
nor U4791 (N_4791,In_337,In_180);
xnor U4792 (N_4792,In_730,In_474);
nor U4793 (N_4793,In_257,In_332);
xor U4794 (N_4794,In_614,In_859);
or U4795 (N_4795,In_767,In_285);
and U4796 (N_4796,In_920,In_204);
nand U4797 (N_4797,In_232,In_521);
nor U4798 (N_4798,In_225,In_383);
nor U4799 (N_4799,In_0,In_212);
or U4800 (N_4800,In_64,In_853);
nand U4801 (N_4801,In_177,In_159);
nor U4802 (N_4802,In_400,In_216);
or U4803 (N_4803,In_557,In_32);
and U4804 (N_4804,In_502,In_324);
nand U4805 (N_4805,In_713,In_842);
and U4806 (N_4806,In_927,In_454);
and U4807 (N_4807,In_818,In_539);
and U4808 (N_4808,In_449,In_340);
nand U4809 (N_4809,In_785,In_330);
nand U4810 (N_4810,In_124,In_655);
and U4811 (N_4811,In_643,In_395);
nor U4812 (N_4812,In_89,In_473);
or U4813 (N_4813,In_845,In_431);
nand U4814 (N_4814,In_132,In_95);
nand U4815 (N_4815,In_391,In_380);
and U4816 (N_4816,In_638,In_351);
and U4817 (N_4817,In_704,In_581);
or U4818 (N_4818,In_821,In_31);
nor U4819 (N_4819,In_47,In_843);
or U4820 (N_4820,In_312,In_84);
xor U4821 (N_4821,In_598,In_278);
nor U4822 (N_4822,In_317,In_713);
and U4823 (N_4823,In_419,In_307);
nor U4824 (N_4824,In_145,In_854);
or U4825 (N_4825,In_767,In_216);
nand U4826 (N_4826,In_396,In_911);
and U4827 (N_4827,In_967,In_178);
or U4828 (N_4828,In_984,In_651);
nand U4829 (N_4829,In_283,In_655);
nor U4830 (N_4830,In_623,In_938);
or U4831 (N_4831,In_31,In_67);
nand U4832 (N_4832,In_694,In_964);
xor U4833 (N_4833,In_332,In_669);
nor U4834 (N_4834,In_468,In_6);
nand U4835 (N_4835,In_919,In_501);
nand U4836 (N_4836,In_798,In_482);
nor U4837 (N_4837,In_501,In_667);
nand U4838 (N_4838,In_138,In_378);
nand U4839 (N_4839,In_193,In_230);
and U4840 (N_4840,In_445,In_783);
or U4841 (N_4841,In_838,In_901);
nand U4842 (N_4842,In_192,In_817);
nor U4843 (N_4843,In_753,In_81);
or U4844 (N_4844,In_686,In_431);
nor U4845 (N_4845,In_744,In_840);
or U4846 (N_4846,In_202,In_712);
nor U4847 (N_4847,In_125,In_547);
or U4848 (N_4848,In_42,In_74);
and U4849 (N_4849,In_967,In_353);
and U4850 (N_4850,In_490,In_763);
nand U4851 (N_4851,In_468,In_798);
xnor U4852 (N_4852,In_952,In_476);
nand U4853 (N_4853,In_712,In_180);
nor U4854 (N_4854,In_767,In_151);
or U4855 (N_4855,In_582,In_212);
and U4856 (N_4856,In_701,In_62);
nand U4857 (N_4857,In_481,In_388);
nor U4858 (N_4858,In_894,In_484);
nor U4859 (N_4859,In_732,In_410);
or U4860 (N_4860,In_229,In_674);
and U4861 (N_4861,In_319,In_667);
and U4862 (N_4862,In_860,In_960);
nand U4863 (N_4863,In_499,In_962);
nand U4864 (N_4864,In_272,In_342);
and U4865 (N_4865,In_628,In_259);
nand U4866 (N_4866,In_901,In_93);
or U4867 (N_4867,In_861,In_445);
nor U4868 (N_4868,In_620,In_592);
nand U4869 (N_4869,In_513,In_982);
nand U4870 (N_4870,In_155,In_469);
nand U4871 (N_4871,In_711,In_268);
xnor U4872 (N_4872,In_124,In_830);
or U4873 (N_4873,In_625,In_593);
nor U4874 (N_4874,In_252,In_335);
nor U4875 (N_4875,In_396,In_409);
nand U4876 (N_4876,In_346,In_479);
and U4877 (N_4877,In_445,In_569);
nand U4878 (N_4878,In_120,In_857);
xnor U4879 (N_4879,In_593,In_110);
nor U4880 (N_4880,In_237,In_980);
nor U4881 (N_4881,In_169,In_8);
nand U4882 (N_4882,In_619,In_108);
or U4883 (N_4883,In_210,In_983);
and U4884 (N_4884,In_78,In_184);
and U4885 (N_4885,In_913,In_230);
nor U4886 (N_4886,In_541,In_141);
or U4887 (N_4887,In_347,In_78);
nor U4888 (N_4888,In_575,In_668);
nor U4889 (N_4889,In_147,In_215);
nand U4890 (N_4890,In_474,In_404);
and U4891 (N_4891,In_192,In_284);
nand U4892 (N_4892,In_627,In_160);
nand U4893 (N_4893,In_789,In_439);
or U4894 (N_4894,In_820,In_243);
or U4895 (N_4895,In_947,In_653);
or U4896 (N_4896,In_186,In_171);
and U4897 (N_4897,In_553,In_817);
or U4898 (N_4898,In_908,In_486);
nor U4899 (N_4899,In_339,In_397);
or U4900 (N_4900,In_828,In_609);
nand U4901 (N_4901,In_933,In_384);
xor U4902 (N_4902,In_87,In_788);
nor U4903 (N_4903,In_974,In_50);
or U4904 (N_4904,In_849,In_605);
or U4905 (N_4905,In_701,In_366);
nor U4906 (N_4906,In_361,In_731);
nor U4907 (N_4907,In_570,In_894);
nand U4908 (N_4908,In_293,In_915);
nor U4909 (N_4909,In_578,In_682);
xnor U4910 (N_4910,In_495,In_394);
xor U4911 (N_4911,In_374,In_956);
nand U4912 (N_4912,In_615,In_603);
and U4913 (N_4913,In_835,In_96);
or U4914 (N_4914,In_491,In_865);
nor U4915 (N_4915,In_24,In_779);
nor U4916 (N_4916,In_38,In_574);
and U4917 (N_4917,In_199,In_948);
xnor U4918 (N_4918,In_278,In_981);
nand U4919 (N_4919,In_476,In_6);
nand U4920 (N_4920,In_92,In_303);
nand U4921 (N_4921,In_902,In_494);
nand U4922 (N_4922,In_837,In_106);
or U4923 (N_4923,In_226,In_116);
nor U4924 (N_4924,In_67,In_557);
or U4925 (N_4925,In_996,In_483);
or U4926 (N_4926,In_67,In_447);
xnor U4927 (N_4927,In_579,In_746);
and U4928 (N_4928,In_593,In_341);
nand U4929 (N_4929,In_145,In_177);
and U4930 (N_4930,In_223,In_774);
or U4931 (N_4931,In_865,In_99);
nor U4932 (N_4932,In_515,In_615);
xnor U4933 (N_4933,In_88,In_103);
and U4934 (N_4934,In_658,In_452);
and U4935 (N_4935,In_967,In_791);
or U4936 (N_4936,In_981,In_632);
or U4937 (N_4937,In_512,In_507);
and U4938 (N_4938,In_16,In_738);
or U4939 (N_4939,In_618,In_118);
and U4940 (N_4940,In_154,In_872);
nor U4941 (N_4941,In_592,In_540);
and U4942 (N_4942,In_496,In_354);
nor U4943 (N_4943,In_140,In_510);
or U4944 (N_4944,In_841,In_803);
nand U4945 (N_4945,In_934,In_615);
or U4946 (N_4946,In_947,In_676);
and U4947 (N_4947,In_121,In_483);
nand U4948 (N_4948,In_661,In_881);
nand U4949 (N_4949,In_189,In_689);
nand U4950 (N_4950,In_319,In_552);
and U4951 (N_4951,In_997,In_310);
nand U4952 (N_4952,In_904,In_702);
or U4953 (N_4953,In_987,In_588);
nor U4954 (N_4954,In_492,In_215);
nand U4955 (N_4955,In_742,In_230);
xor U4956 (N_4956,In_116,In_378);
and U4957 (N_4957,In_833,In_415);
and U4958 (N_4958,In_279,In_584);
nor U4959 (N_4959,In_356,In_332);
and U4960 (N_4960,In_188,In_907);
nor U4961 (N_4961,In_279,In_318);
and U4962 (N_4962,In_514,In_197);
or U4963 (N_4963,In_225,In_723);
xor U4964 (N_4964,In_851,In_0);
and U4965 (N_4965,In_717,In_281);
and U4966 (N_4966,In_360,In_237);
xor U4967 (N_4967,In_903,In_921);
nand U4968 (N_4968,In_457,In_290);
or U4969 (N_4969,In_627,In_792);
nand U4970 (N_4970,In_653,In_730);
and U4971 (N_4971,In_693,In_853);
and U4972 (N_4972,In_684,In_456);
and U4973 (N_4973,In_176,In_825);
xnor U4974 (N_4974,In_732,In_74);
nor U4975 (N_4975,In_212,In_281);
nand U4976 (N_4976,In_667,In_951);
xnor U4977 (N_4977,In_46,In_143);
nand U4978 (N_4978,In_485,In_66);
or U4979 (N_4979,In_801,In_675);
nor U4980 (N_4980,In_719,In_217);
or U4981 (N_4981,In_5,In_232);
xnor U4982 (N_4982,In_204,In_682);
and U4983 (N_4983,In_283,In_810);
xnor U4984 (N_4984,In_343,In_412);
nor U4985 (N_4985,In_179,In_992);
or U4986 (N_4986,In_740,In_538);
or U4987 (N_4987,In_650,In_760);
nor U4988 (N_4988,In_82,In_988);
nor U4989 (N_4989,In_286,In_878);
and U4990 (N_4990,In_829,In_359);
and U4991 (N_4991,In_469,In_581);
xnor U4992 (N_4992,In_200,In_642);
nor U4993 (N_4993,In_105,In_957);
or U4994 (N_4994,In_183,In_866);
or U4995 (N_4995,In_601,In_264);
and U4996 (N_4996,In_908,In_595);
or U4997 (N_4997,In_215,In_924);
or U4998 (N_4998,In_510,In_168);
nand U4999 (N_4999,In_598,In_975);
and U5000 (N_5000,N_2993,N_2797);
nor U5001 (N_5001,N_40,N_472);
nand U5002 (N_5002,N_4777,N_3493);
nor U5003 (N_5003,N_1716,N_1807);
nand U5004 (N_5004,N_1269,N_4296);
and U5005 (N_5005,N_3826,N_4426);
nor U5006 (N_5006,N_3412,N_4001);
and U5007 (N_5007,N_3623,N_4559);
nand U5008 (N_5008,N_4486,N_4344);
nand U5009 (N_5009,N_189,N_3257);
or U5010 (N_5010,N_3761,N_3479);
or U5011 (N_5011,N_417,N_166);
and U5012 (N_5012,N_2855,N_4314);
or U5013 (N_5013,N_904,N_4568);
or U5014 (N_5014,N_3009,N_424);
or U5015 (N_5015,N_1880,N_3325);
and U5016 (N_5016,N_2388,N_2214);
or U5017 (N_5017,N_1945,N_4576);
nor U5018 (N_5018,N_82,N_1219);
xnor U5019 (N_5019,N_996,N_1380);
and U5020 (N_5020,N_1841,N_829);
xor U5021 (N_5021,N_1637,N_1317);
or U5022 (N_5022,N_2881,N_3357);
xnor U5023 (N_5023,N_3705,N_2460);
xor U5024 (N_5024,N_489,N_3990);
nand U5025 (N_5025,N_4165,N_104);
nor U5026 (N_5026,N_4375,N_1700);
nand U5027 (N_5027,N_3063,N_4928);
and U5028 (N_5028,N_2077,N_3622);
xnor U5029 (N_5029,N_67,N_3133);
and U5030 (N_5030,N_4851,N_636);
or U5031 (N_5031,N_1672,N_3634);
nand U5032 (N_5032,N_3744,N_3079);
xor U5033 (N_5033,N_2637,N_3502);
nand U5034 (N_5034,N_4520,N_1001);
nor U5035 (N_5035,N_1053,N_3686);
or U5036 (N_5036,N_2358,N_4206);
and U5037 (N_5037,N_1514,N_1830);
or U5038 (N_5038,N_860,N_3427);
xor U5039 (N_5039,N_3684,N_4893);
nor U5040 (N_5040,N_3287,N_3296);
or U5041 (N_5041,N_603,N_4709);
nor U5042 (N_5042,N_1545,N_1937);
nor U5043 (N_5043,N_1467,N_1277);
xor U5044 (N_5044,N_3958,N_3323);
nor U5045 (N_5045,N_3532,N_4830);
and U5046 (N_5046,N_4698,N_626);
and U5047 (N_5047,N_461,N_4751);
and U5048 (N_5048,N_2449,N_3712);
and U5049 (N_5049,N_1926,N_2249);
or U5050 (N_5050,N_1237,N_4388);
xnor U5051 (N_5051,N_4909,N_4731);
and U5052 (N_5052,N_4645,N_1615);
nand U5053 (N_5053,N_4405,N_3980);
nor U5054 (N_5054,N_3887,N_2693);
or U5055 (N_5055,N_585,N_555);
and U5056 (N_5056,N_3458,N_1373);
nand U5057 (N_5057,N_3028,N_510);
or U5058 (N_5058,N_2166,N_2288);
or U5059 (N_5059,N_4607,N_4360);
nor U5060 (N_5060,N_2819,N_4288);
and U5061 (N_5061,N_2255,N_1749);
or U5062 (N_5062,N_2152,N_760);
and U5063 (N_5063,N_3938,N_1168);
or U5064 (N_5064,N_4594,N_2731);
nor U5065 (N_5065,N_2754,N_4438);
or U5066 (N_5066,N_1871,N_4646);
nor U5067 (N_5067,N_4113,N_1155);
or U5068 (N_5068,N_1264,N_3434);
nand U5069 (N_5069,N_3619,N_4549);
nand U5070 (N_5070,N_3656,N_3270);
nand U5071 (N_5071,N_4184,N_2656);
nor U5072 (N_5072,N_4975,N_4);
nor U5073 (N_5073,N_2704,N_4944);
nand U5074 (N_5074,N_3056,N_2368);
nand U5075 (N_5075,N_1726,N_2064);
nor U5076 (N_5076,N_854,N_3967);
and U5077 (N_5077,N_1013,N_3222);
or U5078 (N_5078,N_2114,N_275);
nand U5079 (N_5079,N_2371,N_1803);
and U5080 (N_5080,N_2685,N_3848);
or U5081 (N_5081,N_530,N_3783);
nor U5082 (N_5082,N_3536,N_776);
and U5083 (N_5083,N_4724,N_4318);
or U5084 (N_5084,N_477,N_4803);
or U5085 (N_5085,N_3422,N_4726);
and U5086 (N_5086,N_474,N_2765);
or U5087 (N_5087,N_511,N_2403);
or U5088 (N_5088,N_3209,N_222);
and U5089 (N_5089,N_2321,N_504);
nor U5090 (N_5090,N_2319,N_568);
or U5091 (N_5091,N_4605,N_1061);
nand U5092 (N_5092,N_3707,N_3109);
and U5093 (N_5093,N_3695,N_2200);
nor U5094 (N_5094,N_4179,N_1699);
and U5095 (N_5095,N_2921,N_1437);
nor U5096 (N_5096,N_2737,N_660);
and U5097 (N_5097,N_4653,N_3919);
xor U5098 (N_5098,N_4373,N_3577);
nor U5099 (N_5099,N_1338,N_3457);
and U5100 (N_5100,N_1466,N_3261);
nor U5101 (N_5101,N_2123,N_1202);
nor U5102 (N_5102,N_3450,N_2581);
nor U5103 (N_5103,N_264,N_1064);
nor U5104 (N_5104,N_4699,N_4313);
and U5105 (N_5105,N_3284,N_3642);
xor U5106 (N_5106,N_4337,N_4558);
nor U5107 (N_5107,N_3282,N_367);
nand U5108 (N_5108,N_1691,N_1402);
and U5109 (N_5109,N_3065,N_3503);
nand U5110 (N_5110,N_2472,N_2065);
nand U5111 (N_5111,N_2341,N_3500);
or U5112 (N_5112,N_2903,N_4585);
or U5113 (N_5113,N_1606,N_1439);
or U5114 (N_5114,N_4215,N_3982);
xor U5115 (N_5115,N_356,N_2565);
nor U5116 (N_5116,N_4850,N_3424);
nor U5117 (N_5117,N_4070,N_2506);
and U5118 (N_5118,N_2751,N_2886);
nor U5119 (N_5119,N_3926,N_1050);
nand U5120 (N_5120,N_1367,N_4458);
or U5121 (N_5121,N_2790,N_999);
nor U5122 (N_5122,N_3105,N_4095);
and U5123 (N_5123,N_617,N_3867);
and U5124 (N_5124,N_4162,N_1149);
nand U5125 (N_5125,N_3561,N_1023);
and U5126 (N_5126,N_3459,N_581);
nor U5127 (N_5127,N_2100,N_4094);
or U5128 (N_5128,N_3117,N_926);
and U5129 (N_5129,N_2399,N_249);
and U5130 (N_5130,N_1921,N_681);
and U5131 (N_5131,N_100,N_4315);
or U5132 (N_5132,N_4092,N_1640);
nand U5133 (N_5133,N_2401,N_955);
or U5134 (N_5134,N_2992,N_2503);
or U5135 (N_5135,N_1190,N_3135);
and U5136 (N_5136,N_4488,N_302);
nand U5137 (N_5137,N_1114,N_230);
and U5138 (N_5138,N_837,N_2684);
or U5139 (N_5139,N_3833,N_4744);
nand U5140 (N_5140,N_452,N_3831);
nand U5141 (N_5141,N_1528,N_741);
nand U5142 (N_5142,N_2818,N_3445);
nor U5143 (N_5143,N_3281,N_1136);
or U5144 (N_5144,N_4783,N_2753);
nor U5145 (N_5145,N_4679,N_3448);
or U5146 (N_5146,N_3004,N_1325);
xor U5147 (N_5147,N_1729,N_932);
nand U5148 (N_5148,N_3751,N_327);
xnor U5149 (N_5149,N_3240,N_3091);
and U5150 (N_5150,N_1026,N_3141);
nor U5151 (N_5151,N_3498,N_1907);
and U5152 (N_5152,N_3675,N_4140);
nand U5153 (N_5153,N_2889,N_1738);
nand U5154 (N_5154,N_2988,N_4236);
and U5155 (N_5155,N_3482,N_4204);
nor U5156 (N_5156,N_2720,N_4167);
nand U5157 (N_5157,N_2702,N_4856);
xor U5158 (N_5158,N_3734,N_4245);
nor U5159 (N_5159,N_1407,N_2750);
nor U5160 (N_5160,N_2582,N_1224);
xnor U5161 (N_5161,N_1475,N_4780);
nor U5162 (N_5162,N_1852,N_4505);
and U5163 (N_5163,N_2430,N_3771);
nor U5164 (N_5164,N_4734,N_4090);
nor U5165 (N_5165,N_4342,N_600);
xor U5166 (N_5166,N_1103,N_4616);
nand U5167 (N_5167,N_4685,N_4989);
nor U5168 (N_5168,N_4966,N_4498);
or U5169 (N_5169,N_1786,N_4742);
nand U5170 (N_5170,N_4769,N_404);
xor U5171 (N_5171,N_3256,N_2643);
or U5172 (N_5172,N_4496,N_3851);
and U5173 (N_5173,N_2650,N_1556);
or U5174 (N_5174,N_4183,N_4190);
and U5175 (N_5175,N_2208,N_3565);
and U5176 (N_5176,N_2682,N_3076);
nand U5177 (N_5177,N_1132,N_4810);
nand U5178 (N_5178,N_2300,N_3368);
nor U5179 (N_5179,N_1319,N_1774);
nor U5180 (N_5180,N_4358,N_1628);
and U5181 (N_5181,N_1660,N_4045);
nor U5182 (N_5182,N_4983,N_3013);
nor U5183 (N_5183,N_1034,N_4740);
nand U5184 (N_5184,N_954,N_3874);
or U5185 (N_5185,N_2777,N_2040);
nand U5186 (N_5186,N_871,N_758);
nand U5187 (N_5187,N_2946,N_4839);
nor U5188 (N_5188,N_528,N_3440);
xnor U5189 (N_5189,N_1707,N_2981);
or U5190 (N_5190,N_4534,N_4763);
nand U5191 (N_5191,N_4720,N_4471);
nand U5192 (N_5192,N_686,N_1265);
nor U5193 (N_5193,N_924,N_1505);
or U5194 (N_5194,N_1567,N_1713);
nor U5195 (N_5195,N_2044,N_1298);
or U5196 (N_5196,N_1827,N_4037);
and U5197 (N_5197,N_4655,N_4553);
nand U5198 (N_5198,N_1553,N_3101);
nand U5199 (N_5199,N_3904,N_1314);
or U5200 (N_5200,N_4050,N_967);
nor U5201 (N_5201,N_2768,N_2175);
xnor U5202 (N_5202,N_2824,N_1175);
or U5203 (N_5203,N_324,N_2461);
nor U5204 (N_5204,N_2260,N_1746);
nand U5205 (N_5205,N_3463,N_1472);
and U5206 (N_5206,N_2969,N_405);
nor U5207 (N_5207,N_4675,N_473);
xnor U5208 (N_5208,N_2714,N_144);
or U5209 (N_5209,N_1164,N_3676);
or U5210 (N_5210,N_418,N_1919);
nor U5211 (N_5211,N_929,N_2961);
or U5212 (N_5212,N_4287,N_593);
or U5213 (N_5213,N_194,N_4382);
nand U5214 (N_5214,N_3989,N_3704);
nand U5215 (N_5215,N_2063,N_3824);
nor U5216 (N_5216,N_4158,N_374);
nor U5217 (N_5217,N_2554,N_723);
xnor U5218 (N_5218,N_1722,N_3379);
or U5219 (N_5219,N_4087,N_4790);
nor U5220 (N_5220,N_1228,N_3782);
or U5221 (N_5221,N_2709,N_279);
or U5222 (N_5222,N_4543,N_1073);
and U5223 (N_5223,N_3398,N_3781);
nand U5224 (N_5224,N_649,N_3177);
nand U5225 (N_5225,N_2222,N_2967);
or U5226 (N_5226,N_2532,N_995);
or U5227 (N_5227,N_1413,N_369);
or U5228 (N_5228,N_3593,N_3384);
nor U5229 (N_5229,N_2631,N_4651);
or U5230 (N_5230,N_634,N_4570);
nor U5231 (N_5231,N_2484,N_4472);
nor U5232 (N_5232,N_2056,N_4331);
nand U5233 (N_5233,N_347,N_4916);
and U5234 (N_5234,N_3114,N_3311);
or U5235 (N_5235,N_4111,N_2259);
nand U5236 (N_5236,N_3346,N_3172);
nand U5237 (N_5237,N_4901,N_1750);
or U5238 (N_5238,N_1708,N_549);
or U5239 (N_5239,N_160,N_1872);
or U5240 (N_5240,N_485,N_688);
nor U5241 (N_5241,N_891,N_3762);
or U5242 (N_5242,N_1205,N_2130);
or U5243 (N_5243,N_4781,N_1352);
xnor U5244 (N_5244,N_65,N_3078);
nor U5245 (N_5245,N_3383,N_450);
nor U5246 (N_5246,N_59,N_4932);
nand U5247 (N_5247,N_670,N_4328);
or U5248 (N_5248,N_3529,N_4362);
and U5249 (N_5249,N_1186,N_2551);
nor U5250 (N_5250,N_4225,N_5);
and U5251 (N_5251,N_200,N_1516);
nand U5252 (N_5252,N_1560,N_2660);
nand U5253 (N_5253,N_4627,N_3594);
nand U5254 (N_5254,N_4809,N_518);
nor U5255 (N_5255,N_3799,N_2926);
or U5256 (N_5256,N_3030,N_917);
nand U5257 (N_5257,N_4067,N_52);
xor U5258 (N_5258,N_810,N_1171);
nor U5259 (N_5259,N_375,N_1574);
or U5260 (N_5260,N_1936,N_3343);
and U5261 (N_5261,N_1383,N_3171);
nand U5262 (N_5262,N_1564,N_4199);
or U5263 (N_5263,N_3018,N_4663);
xor U5264 (N_5264,N_4141,N_3241);
and U5265 (N_5265,N_2995,N_1123);
nand U5266 (N_5266,N_4500,N_3407);
or U5267 (N_5267,N_1953,N_2272);
and U5268 (N_5268,N_58,N_1977);
and U5269 (N_5269,N_2635,N_23);
and U5270 (N_5270,N_2671,N_4016);
and U5271 (N_5271,N_3406,N_2812);
nor U5272 (N_5272,N_3579,N_4899);
or U5273 (N_5273,N_4317,N_1820);
and U5274 (N_5274,N_1506,N_3258);
or U5275 (N_5275,N_1347,N_1826);
or U5276 (N_5276,N_812,N_139);
or U5277 (N_5277,N_3580,N_1635);
and U5278 (N_5278,N_396,N_1605);
nand U5279 (N_5279,N_2354,N_1748);
nor U5280 (N_5280,N_1282,N_3564);
or U5281 (N_5281,N_3721,N_976);
or U5282 (N_5282,N_4181,N_3745);
or U5283 (N_5283,N_586,N_3737);
or U5284 (N_5284,N_2396,N_4421);
and U5285 (N_5285,N_3150,N_1914);
and U5286 (N_5286,N_3962,N_2692);
or U5287 (N_5287,N_3116,N_1670);
and U5288 (N_5288,N_902,N_2746);
and U5289 (N_5289,N_614,N_1823);
nand U5290 (N_5290,N_346,N_3906);
or U5291 (N_5291,N_4692,N_1844);
xor U5292 (N_5292,N_3756,N_3167);
and U5293 (N_5293,N_4175,N_3560);
nor U5294 (N_5294,N_1372,N_3942);
nand U5295 (N_5295,N_3211,N_1249);
and U5296 (N_5296,N_1012,N_1244);
and U5297 (N_5297,N_1736,N_1889);
nand U5298 (N_5298,N_1197,N_1692);
nor U5299 (N_5299,N_2963,N_1459);
and U5300 (N_5300,N_3128,N_3333);
or U5301 (N_5301,N_219,N_3148);
or U5302 (N_5302,N_803,N_2030);
and U5303 (N_5303,N_3058,N_3681);
nor U5304 (N_5304,N_4670,N_608);
nand U5305 (N_5305,N_2075,N_3739);
nand U5306 (N_5306,N_4620,N_4606);
nor U5307 (N_5307,N_4355,N_717);
nand U5308 (N_5308,N_1084,N_2181);
and U5309 (N_5309,N_2320,N_4752);
or U5310 (N_5310,N_2990,N_1795);
nand U5311 (N_5311,N_4511,N_2932);
nand U5312 (N_5312,N_3677,N_4483);
or U5313 (N_5313,N_1327,N_2872);
nor U5314 (N_5314,N_2770,N_1311);
nor U5315 (N_5315,N_4213,N_1559);
or U5316 (N_5316,N_711,N_3191);
xor U5317 (N_5317,N_1394,N_1502);
or U5318 (N_5318,N_2322,N_1715);
nand U5319 (N_5319,N_1873,N_3868);
xnor U5320 (N_5320,N_355,N_363);
nand U5321 (N_5321,N_2562,N_4243);
or U5322 (N_5322,N_2176,N_1411);
nand U5323 (N_5323,N_3159,N_4361);
and U5324 (N_5324,N_3516,N_3129);
nand U5325 (N_5325,N_4435,N_68);
nor U5326 (N_5326,N_1705,N_77);
and U5327 (N_5327,N_1293,N_685);
nand U5328 (N_5328,N_1712,N_4530);
and U5329 (N_5329,N_4794,N_2463);
or U5330 (N_5330,N_3937,N_4682);
nor U5331 (N_5331,N_1482,N_2201);
nand U5332 (N_5332,N_1866,N_1141);
nor U5333 (N_5333,N_4256,N_3189);
nand U5334 (N_5334,N_2079,N_628);
nand U5335 (N_5335,N_246,N_1343);
or U5336 (N_5336,N_903,N_4604);
nand U5337 (N_5337,N_1610,N_1818);
or U5338 (N_5338,N_3059,N_1834);
xor U5339 (N_5339,N_3511,N_80);
or U5340 (N_5340,N_3016,N_2584);
nand U5341 (N_5341,N_2337,N_188);
xnor U5342 (N_5342,N_2864,N_3316);
or U5343 (N_5343,N_4918,N_4051);
nand U5344 (N_5344,N_3266,N_2060);
and U5345 (N_5345,N_894,N_4702);
nor U5346 (N_5346,N_1690,N_535);
and U5347 (N_5347,N_2909,N_3);
or U5348 (N_5348,N_4381,N_3236);
nand U5349 (N_5349,N_3208,N_2593);
xnor U5350 (N_5350,N_1143,N_1206);
nor U5351 (N_5351,N_2764,N_2221);
and U5352 (N_5352,N_3539,N_3596);
xor U5353 (N_5353,N_2977,N_9);
nor U5354 (N_5354,N_2140,N_2150);
xnor U5355 (N_5355,N_1231,N_2235);
and U5356 (N_5356,N_3408,N_1580);
nor U5357 (N_5357,N_2474,N_3069);
nor U5358 (N_5358,N_4883,N_3370);
xor U5359 (N_5359,N_3553,N_3404);
nor U5360 (N_5360,N_1461,N_4261);
and U5361 (N_5361,N_972,N_1965);
nand U5362 (N_5362,N_1315,N_247);
and U5363 (N_5363,N_2113,N_3274);
nor U5364 (N_5364,N_707,N_3181);
xnor U5365 (N_5365,N_2,N_4135);
nand U5366 (N_5366,N_3431,N_3390);
or U5367 (N_5367,N_1360,N_1170);
nor U5368 (N_5368,N_1732,N_3025);
nor U5369 (N_5369,N_3854,N_4914);
or U5370 (N_5370,N_2293,N_1201);
nand U5371 (N_5371,N_233,N_296);
and U5372 (N_5372,N_2223,N_4062);
nand U5373 (N_5373,N_881,N_1225);
nand U5374 (N_5374,N_4541,N_4833);
nand U5375 (N_5375,N_495,N_3504);
nand U5376 (N_5376,N_3402,N_1445);
nor U5377 (N_5377,N_3984,N_4160);
and U5378 (N_5378,N_151,N_2942);
nand U5379 (N_5379,N_1337,N_1718);
and U5380 (N_5380,N_3715,N_177);
and U5381 (N_5381,N_4995,N_574);
xnor U5382 (N_5382,N_2241,N_1377);
nand U5383 (N_5383,N_3415,N_2048);
nand U5384 (N_5384,N_1025,N_3462);
nor U5385 (N_5385,N_2149,N_3772);
nor U5386 (N_5386,N_2132,N_4867);
nand U5387 (N_5387,N_1891,N_468);
nand U5388 (N_5388,N_3071,N_1552);
or U5389 (N_5389,N_2829,N_1744);
and U5390 (N_5390,N_3336,N_2196);
xor U5391 (N_5391,N_4996,N_4115);
and U5392 (N_5392,N_3889,N_4696);
xor U5393 (N_5393,N_1994,N_2879);
or U5394 (N_5394,N_2105,N_744);
or U5395 (N_5395,N_2273,N_520);
nand U5396 (N_5396,N_4578,N_4778);
nor U5397 (N_5397,N_3007,N_4715);
nor U5398 (N_5398,N_2447,N_2772);
and U5399 (N_5399,N_4253,N_2070);
or U5400 (N_5400,N_4068,N_4272);
xor U5401 (N_5401,N_3625,N_656);
or U5402 (N_5402,N_4172,N_2359);
or U5403 (N_5403,N_1809,N_3574);
nor U5404 (N_5404,N_2561,N_3331);
and U5405 (N_5405,N_3041,N_1306);
nand U5406 (N_5406,N_2949,N_2187);
or U5407 (N_5407,N_1883,N_839);
nor U5408 (N_5408,N_4852,N_826);
or U5409 (N_5409,N_4054,N_2604);
nor U5410 (N_5410,N_1522,N_1757);
and U5411 (N_5411,N_951,N_3245);
nor U5412 (N_5412,N_74,N_2155);
xnor U5413 (N_5413,N_4625,N_865);
nor U5414 (N_5414,N_3365,N_1476);
nor U5415 (N_5415,N_4567,N_352);
and U5416 (N_5416,N_4286,N_2545);
or U5417 (N_5417,N_4716,N_4028);
and U5418 (N_5418,N_4465,N_3917);
or U5419 (N_5419,N_782,N_3521);
nand U5420 (N_5420,N_1385,N_2712);
and U5421 (N_5421,N_721,N_403);
xnor U5422 (N_5422,N_20,N_3275);
and U5423 (N_5423,N_272,N_4409);
nand U5424 (N_5424,N_414,N_2876);
nand U5425 (N_5425,N_2638,N_3183);
xnor U5426 (N_5426,N_728,N_1790);
nand U5427 (N_5427,N_98,N_3798);
and U5428 (N_5428,N_1200,N_4522);
nand U5429 (N_5429,N_2315,N_3871);
or U5430 (N_5430,N_3858,N_3436);
or U5431 (N_5431,N_2115,N_1646);
nand U5432 (N_5432,N_978,N_4484);
or U5433 (N_5433,N_2464,N_4687);
and U5434 (N_5434,N_4209,N_3785);
nand U5435 (N_5435,N_17,N_3347);
nand U5436 (N_5436,N_704,N_4592);
and U5437 (N_5437,N_455,N_2179);
nand U5438 (N_5438,N_1008,N_2453);
and U5439 (N_5439,N_3053,N_4499);
nand U5440 (N_5440,N_2045,N_2156);
or U5441 (N_5441,N_507,N_4007);
nand U5442 (N_5442,N_1000,N_2807);
xor U5443 (N_5443,N_3100,N_604);
nor U5444 (N_5444,N_1920,N_1330);
xor U5445 (N_5445,N_3216,N_3678);
nor U5446 (N_5446,N_1077,N_4903);
and U5447 (N_5447,N_3770,N_2280);
nor U5448 (N_5448,N_1817,N_2698);
nor U5449 (N_5449,N_1022,N_3235);
nand U5450 (N_5450,N_4582,N_2345);
nor U5451 (N_5451,N_2552,N_4517);
xor U5452 (N_5452,N_483,N_1800);
nand U5453 (N_5453,N_3127,N_26);
xnor U5454 (N_5454,N_251,N_4890);
xor U5455 (N_5455,N_3738,N_1566);
and U5456 (N_5456,N_43,N_4325);
or U5457 (N_5457,N_3724,N_934);
nand U5458 (N_5458,N_2933,N_538);
and U5459 (N_5459,N_4566,N_1032);
nor U5460 (N_5460,N_237,N_1877);
or U5461 (N_5461,N_3891,N_2182);
or U5462 (N_5462,N_3376,N_1855);
nand U5463 (N_5463,N_381,N_1821);
nand U5464 (N_5464,N_979,N_4531);
and U5465 (N_5465,N_178,N_3757);
and U5466 (N_5466,N_1323,N_4299);
nor U5467 (N_5467,N_1704,N_1333);
xnor U5468 (N_5468,N_3020,N_3363);
and U5469 (N_5469,N_2402,N_3915);
nor U5470 (N_5470,N_3923,N_428);
xnor U5471 (N_5471,N_393,N_3375);
and U5472 (N_5472,N_170,N_390);
xnor U5473 (N_5473,N_4502,N_605);
nor U5474 (N_5474,N_3327,N_2468);
nor U5475 (N_5475,N_6,N_759);
nor U5476 (N_5476,N_4469,N_3567);
nand U5477 (N_5477,N_328,N_2456);
or U5478 (N_5478,N_2325,N_2137);
nand U5479 (N_5479,N_2499,N_2571);
or U5480 (N_5480,N_1932,N_11);
or U5481 (N_5481,N_1875,N_813);
nor U5482 (N_5482,N_4665,N_654);
or U5483 (N_5483,N_4863,N_3293);
and U5484 (N_5484,N_544,N_3163);
and U5485 (N_5485,N_2502,N_2122);
or U5486 (N_5486,N_740,N_1091);
nand U5487 (N_5487,N_46,N_4601);
nor U5488 (N_5488,N_2015,N_1931);
nor U5489 (N_5489,N_1524,N_2494);
nor U5490 (N_5490,N_1204,N_3410);
and U5491 (N_5491,N_158,N_1568);
nor U5492 (N_5492,N_206,N_1667);
and U5493 (N_5493,N_130,N_126);
or U5494 (N_5494,N_2420,N_3339);
or U5495 (N_5495,N_157,N_597);
xor U5496 (N_5496,N_3048,N_3735);
nor U5497 (N_5497,N_3371,N_1794);
and U5498 (N_5498,N_3291,N_3870);
or U5499 (N_5499,N_4922,N_907);
and U5500 (N_5500,N_578,N_3358);
or U5501 (N_5501,N_1978,N_451);
and U5502 (N_5502,N_3229,N_1048);
or U5503 (N_5503,N_3470,N_2462);
nor U5504 (N_5504,N_4136,N_890);
or U5505 (N_5505,N_1003,N_15);
or U5506 (N_5506,N_3916,N_3843);
nor U5507 (N_5507,N_2603,N_2574);
and U5508 (N_5508,N_770,N_273);
nor U5509 (N_5509,N_4906,N_97);
and U5510 (N_5510,N_947,N_2939);
or U5511 (N_5511,N_3689,N_1428);
xnor U5512 (N_5512,N_1539,N_1430);
nor U5513 (N_5513,N_609,N_3232);
nand U5514 (N_5514,N_4324,N_62);
or U5515 (N_5515,N_3694,N_156);
xnor U5516 (N_5516,N_2711,N_2342);
or U5517 (N_5517,N_877,N_2034);
and U5518 (N_5518,N_496,N_4871);
and U5519 (N_5519,N_2883,N_1666);
or U5520 (N_5520,N_2073,N_2636);
nand U5521 (N_5521,N_3305,N_4595);
nand U5522 (N_5522,N_4292,N_1416);
and U5523 (N_5523,N_1874,N_4532);
or U5524 (N_5524,N_3491,N_1894);
or U5525 (N_5525,N_3153,N_4659);
xor U5526 (N_5526,N_3146,N_1530);
nor U5527 (N_5527,N_3790,N_4117);
nand U5528 (N_5528,N_1040,N_3354);
xnor U5529 (N_5529,N_2466,N_2126);
and U5530 (N_5530,N_2076,N_1088);
nor U5531 (N_5531,N_2590,N_480);
nand U5532 (N_5532,N_2815,N_1942);
nor U5533 (N_5533,N_3846,N_4987);
and U5534 (N_5534,N_4684,N_2487);
and U5535 (N_5535,N_774,N_3892);
xor U5536 (N_5536,N_962,N_1518);
nor U5537 (N_5537,N_1375,N_2111);
nor U5538 (N_5538,N_3556,N_1845);
nand U5539 (N_5539,N_1166,N_1102);
nor U5540 (N_5540,N_1954,N_3743);
and U5541 (N_5541,N_4211,N_1090);
nand U5542 (N_5542,N_2691,N_1253);
and U5543 (N_5543,N_2544,N_1620);
nand U5544 (N_5544,N_2124,N_1625);
nor U5545 (N_5545,N_1928,N_3476);
nor U5546 (N_5546,N_862,N_3897);
nor U5547 (N_5547,N_2483,N_1263);
and U5548 (N_5548,N_1527,N_86);
xor U5549 (N_5549,N_3960,N_3506);
nand U5550 (N_5550,N_900,N_847);
or U5551 (N_5551,N_1859,N_1976);
or U5552 (N_5552,N_3086,N_4341);
nand U5553 (N_5553,N_434,N_580);
nand U5554 (N_5554,N_4947,N_1836);
and U5555 (N_5555,N_2177,N_3158);
xnor U5556 (N_5556,N_3535,N_3344);
xnor U5557 (N_5557,N_2411,N_2163);
or U5558 (N_5558,N_2231,N_2431);
nand U5559 (N_5559,N_790,N_1621);
or U5560 (N_5560,N_1822,N_4902);
or U5561 (N_5561,N_992,N_3941);
nor U5562 (N_5562,N_554,N_2384);
nor U5563 (N_5563,N_259,N_4377);
or U5564 (N_5564,N_4806,N_4424);
xnor U5565 (N_5565,N_385,N_4557);
and U5566 (N_5566,N_1501,N_4835);
or U5567 (N_5567,N_4628,N_49);
xnor U5568 (N_5568,N_2350,N_1848);
or U5569 (N_5569,N_2563,N_792);
and U5570 (N_5570,N_3481,N_2882);
nand U5571 (N_5571,N_1256,N_1905);
nor U5572 (N_5572,N_4357,N_2266);
nand U5573 (N_5573,N_1612,N_3524);
or U5574 (N_5574,N_3309,N_261);
nor U5575 (N_5575,N_2726,N_2110);
nand U5576 (N_5576,N_3075,N_4473);
or U5577 (N_5577,N_3471,N_3433);
and U5578 (N_5578,N_1110,N_3921);
and U5579 (N_5579,N_630,N_290);
or U5580 (N_5580,N_3223,N_809);
nor U5581 (N_5581,N_3196,N_863);
nand U5582 (N_5582,N_4587,N_2190);
xor U5583 (N_5583,N_3050,N_4476);
nand U5584 (N_5584,N_1387,N_3237);
and U5585 (N_5585,N_4926,N_570);
or U5586 (N_5586,N_69,N_1128);
nor U5587 (N_5587,N_2007,N_4180);
or U5588 (N_5588,N_2811,N_205);
or U5589 (N_5589,N_2539,N_1238);
nand U5590 (N_5590,N_1677,N_506);
nand U5591 (N_5591,N_2490,N_2608);
nor U5592 (N_5592,N_3378,N_2756);
nor U5593 (N_5593,N_2805,N_1710);
nand U5594 (N_5594,N_4550,N_1235);
xor U5595 (N_5595,N_1882,N_3545);
nand U5596 (N_5596,N_4188,N_2804);
nor U5597 (N_5597,N_3000,N_2840);
or U5598 (N_5598,N_4937,N_3137);
or U5599 (N_5599,N_4750,N_2305);
or U5600 (N_5600,N_4800,N_362);
nand U5601 (N_5601,N_4992,N_2471);
nand U5602 (N_5602,N_2372,N_2413);
nor U5603 (N_5603,N_3497,N_1473);
nand U5604 (N_5604,N_204,N_1036);
and U5605 (N_5605,N_4609,N_3525);
or U5606 (N_5606,N_2640,N_3213);
xnor U5607 (N_5607,N_4254,N_3204);
and U5608 (N_5608,N_969,N_2159);
nor U5609 (N_5609,N_3943,N_2258);
or U5610 (N_5610,N_1104,N_778);
and U5611 (N_5611,N_905,N_2779);
and U5612 (N_5612,N_3420,N_2923);
or U5613 (N_5613,N_2511,N_1629);
and U5614 (N_5614,N_1869,N_2950);
and U5615 (N_5615,N_224,N_211);
or U5616 (N_5616,N_4635,N_4432);
and U5617 (N_5617,N_933,N_3277);
and U5618 (N_5618,N_3933,N_3038);
xor U5619 (N_5619,N_1184,N_3184);
nand U5620 (N_5620,N_4564,N_3125);
nand U5621 (N_5621,N_2173,N_3388);
nand U5622 (N_5622,N_4817,N_588);
xor U5623 (N_5623,N_1101,N_1199);
nor U5624 (N_5624,N_2517,N_1838);
and U5625 (N_5625,N_426,N_2618);
xnor U5626 (N_5626,N_382,N_4029);
nor U5627 (N_5627,N_2894,N_4281);
nor U5628 (N_5628,N_1938,N_3015);
or U5629 (N_5629,N_10,N_923);
nand U5630 (N_5630,N_3659,N_3262);
or U5631 (N_5631,N_4487,N_4949);
or U5632 (N_5632,N_4088,N_3042);
xnor U5633 (N_5633,N_4668,N_3823);
nor U5634 (N_5634,N_4142,N_874);
and U5635 (N_5635,N_906,N_225);
nand U5636 (N_5636,N_3667,N_4295);
and U5637 (N_5637,N_1085,N_4516);
and U5638 (N_5638,N_930,N_1831);
or U5639 (N_5639,N_1902,N_769);
nand U5640 (N_5640,N_4394,N_1582);
nor U5641 (N_5641,N_447,N_3162);
and U5642 (N_5642,N_2615,N_532);
nor U5643 (N_5643,N_1353,N_3691);
and U5644 (N_5644,N_3526,N_2701);
and U5645 (N_5645,N_3112,N_4759);
nand U5646 (N_5646,N_4304,N_2721);
xor U5647 (N_5647,N_203,N_2005);
nand U5648 (N_5648,N_3607,N_3718);
or U5649 (N_5649,N_1366,N_3246);
nand U5650 (N_5650,N_1543,N_4227);
or U5651 (N_5651,N_4451,N_2659);
nor U5652 (N_5652,N_590,N_4434);
nor U5653 (N_5653,N_4194,N_4754);
nand U5654 (N_5654,N_3731,N_4411);
nor U5655 (N_5655,N_3193,N_34);
nor U5656 (N_5656,N_1015,N_2717);
or U5657 (N_5657,N_3850,N_2778);
nand U5658 (N_5658,N_3813,N_500);
or U5659 (N_5659,N_4084,N_3072);
or U5660 (N_5660,N_270,N_351);
xor U5661 (N_5661,N_2645,N_4422);
or U5662 (N_5662,N_1607,N_1187);
nand U5663 (N_5663,N_2664,N_4077);
or U5664 (N_5664,N_2390,N_2766);
xor U5665 (N_5665,N_3883,N_3317);
nand U5666 (N_5666,N_99,N_4642);
or U5667 (N_5667,N_3366,N_2347);
or U5668 (N_5668,N_4010,N_3312);
nor U5669 (N_5669,N_3602,N_171);
nor U5670 (N_5670,N_1335,N_3838);
or U5671 (N_5671,N_1151,N_2039);
nor U5672 (N_5672,N_3138,N_4814);
nand U5673 (N_5673,N_2619,N_4746);
and U5674 (N_5674,N_729,N_4953);
nor U5675 (N_5675,N_4346,N_2180);
nand U5676 (N_5676,N_3429,N_2242);
nor U5677 (N_5677,N_3849,N_2728);
xor U5678 (N_5678,N_1232,N_2433);
nor U5679 (N_5679,N_2687,N_3061);
or U5680 (N_5680,N_2979,N_724);
nand U5681 (N_5681,N_950,N_1059);
xnor U5682 (N_5682,N_260,N_4491);
nand U5683 (N_5683,N_50,N_4957);
xnor U5684 (N_5684,N_3590,N_4598);
nor U5685 (N_5685,N_1631,N_332);
nor U5686 (N_5686,N_4834,N_2407);
nand U5687 (N_5687,N_4563,N_4440);
or U5688 (N_5688,N_2316,N_1198);
nand U5689 (N_5689,N_3049,N_516);
nand U5690 (N_5690,N_4691,N_4704);
nand U5691 (N_5691,N_12,N_3108);
or U5692 (N_5692,N_3180,N_181);
nand U5693 (N_5693,N_3628,N_4848);
nand U5694 (N_5694,N_113,N_4047);
and U5695 (N_5695,N_800,N_1);
nor U5696 (N_5696,N_1410,N_742);
and U5697 (N_5697,N_2445,N_2252);
or U5698 (N_5698,N_2880,N_3541);
and U5699 (N_5699,N_2160,N_557);
nor U5700 (N_5700,N_3991,N_75);
nor U5701 (N_5701,N_1140,N_3592);
or U5702 (N_5702,N_1510,N_1266);
nand U5703 (N_5703,N_3608,N_1989);
and U5704 (N_5704,N_30,N_3255);
nor U5705 (N_5705,N_2740,N_129);
and U5706 (N_5706,N_117,N_4707);
nand U5707 (N_5707,N_1208,N_2980);
nor U5708 (N_5708,N_3537,N_4186);
nand U5709 (N_5709,N_2108,N_3029);
nor U5710 (N_5710,N_2592,N_1734);
nand U5711 (N_5711,N_2412,N_4109);
and U5712 (N_5712,N_1010,N_1259);
nand U5713 (N_5713,N_625,N_527);
or U5714 (N_5714,N_1192,N_3454);
and U5715 (N_5715,N_364,N_4981);
nand U5716 (N_5716,N_1918,N_3488);
nor U5717 (N_5717,N_357,N_421);
and U5718 (N_5718,N_644,N_4976);
or U5719 (N_5719,N_1496,N_968);
nand U5720 (N_5720,N_2080,N_3759);
nand U5721 (N_5721,N_3494,N_1065);
and U5722 (N_5722,N_3505,N_4683);
nand U5723 (N_5723,N_2871,N_3332);
xnor U5724 (N_5724,N_2446,N_4705);
nand U5725 (N_5725,N_780,N_1728);
or U5726 (N_5726,N_3290,N_2304);
xnor U5727 (N_5727,N_591,N_2860);
nand U5728 (N_5728,N_1854,N_3742);
and U5729 (N_5729,N_2188,N_3732);
xor U5730 (N_5730,N_884,N_882);
nand U5731 (N_5731,N_1671,N_3095);
or U5732 (N_5732,N_4396,N_2526);
and U5733 (N_5733,N_4121,N_437);
nor U5734 (N_5734,N_2697,N_2218);
nor U5735 (N_5735,N_4756,N_4182);
nand U5736 (N_5736,N_4154,N_2212);
nand U5737 (N_5737,N_1188,N_2246);
or U5738 (N_5738,N_1074,N_3238);
and U5739 (N_5739,N_3834,N_146);
nor U5740 (N_5740,N_3242,N_2793);
and U5741 (N_5741,N_4634,N_4743);
or U5742 (N_5742,N_3700,N_4539);
nand U5743 (N_5743,N_3839,N_2579);
or U5744 (N_5744,N_2004,N_3377);
nand U5745 (N_5745,N_4501,N_1887);
xor U5746 (N_5746,N_2870,N_4573);
and U5747 (N_5747,N_2674,N_4100);
and U5748 (N_5748,N_3685,N_4450);
and U5749 (N_5749,N_3568,N_2822);
xnor U5750 (N_5750,N_795,N_4443);
or U5751 (N_5751,N_1630,N_4372);
nand U5752 (N_5752,N_4379,N_3558);
and U5753 (N_5753,N_913,N_4640);
and U5754 (N_5754,N_1477,N_548);
nand U5755 (N_5755,N_658,N_1763);
nor U5756 (N_5756,N_1986,N_3528);
and U5757 (N_5757,N_2008,N_2029);
nand U5758 (N_5758,N_2213,N_3083);
nand U5759 (N_5759,N_138,N_3819);
and U5760 (N_5760,N_2285,N_1997);
nand U5761 (N_5761,N_1068,N_2540);
nor U5762 (N_5762,N_935,N_2813);
nor U5763 (N_5763,N_1569,N_1575);
nor U5764 (N_5764,N_1047,N_2944);
and U5765 (N_5765,N_4226,N_4921);
nor U5766 (N_5766,N_3810,N_602);
nand U5767 (N_5767,N_3268,N_2943);
and U5768 (N_5768,N_659,N_4590);
or U5769 (N_5769,N_192,N_1424);
nand U5770 (N_5770,N_3627,N_14);
nand U5771 (N_5771,N_1292,N_2014);
nand U5772 (N_5772,N_4069,N_1131);
xnor U5773 (N_5773,N_2706,N_3549);
nand U5774 (N_5774,N_946,N_1272);
or U5775 (N_5775,N_1868,N_2862);
or U5776 (N_5776,N_749,N_2578);
nand U5777 (N_5777,N_3187,N_2957);
nand U5778 (N_5778,N_3643,N_1492);
nor U5779 (N_5779,N_3396,N_4721);
nand U5780 (N_5780,N_1180,N_2877);
nand U5781 (N_5781,N_2081,N_2143);
and U5782 (N_5782,N_3859,N_3950);
xor U5783 (N_5783,N_3423,N_612);
xnor U5784 (N_5784,N_2363,N_1913);
nor U5785 (N_5785,N_1546,N_4555);
xnor U5786 (N_5786,N_1028,N_3555);
nand U5787 (N_5787,N_1395,N_2836);
or U5788 (N_5788,N_2375,N_3609);
nor U5789 (N_5789,N_1161,N_4657);
and U5790 (N_5790,N_692,N_2243);
and U5791 (N_5791,N_4747,N_2101);
nor U5792 (N_5792,N_321,N_4026);
and U5793 (N_5793,N_1899,N_3725);
xnor U5794 (N_5794,N_2856,N_2795);
xor U5795 (N_5795,N_4453,N_1586);
nand U5796 (N_5796,N_2700,N_3690);
or U5797 (N_5797,N_2331,N_4250);
nor U5798 (N_5798,N_2282,N_3760);
xnor U5799 (N_5799,N_4770,N_462);
nand U5800 (N_5800,N_753,N_1756);
xor U5801 (N_5801,N_2896,N_3401);
nand U5802 (N_5802,N_2865,N_2928);
nor U5803 (N_5803,N_1351,N_3164);
nor U5804 (N_5804,N_1464,N_2542);
or U5805 (N_5805,N_1438,N_3382);
nand U5806 (N_5806,N_1011,N_1862);
and U5807 (N_5807,N_2703,N_4266);
nand U5808 (N_5808,N_1489,N_4329);
nand U5809 (N_5809,N_3961,N_4711);
or U5810 (N_5810,N_1488,N_1747);
nand U5811 (N_5811,N_4005,N_1896);
nand U5812 (N_5812,N_4941,N_4060);
nand U5813 (N_5813,N_4255,N_3748);
xnor U5814 (N_5814,N_1979,N_184);
and U5815 (N_5815,N_1099,N_1046);
or U5816 (N_5816,N_4464,N_4228);
and U5817 (N_5817,N_928,N_4290);
nand U5818 (N_5818,N_345,N_2941);
nor U5819 (N_5819,N_1376,N_4401);
or U5820 (N_5820,N_623,N_615);
nand U5821 (N_5821,N_4764,N_4086);
and U5822 (N_5822,N_4792,N_213);
or U5823 (N_5823,N_1515,N_4017);
or U5824 (N_5824,N_4729,N_1557);
and U5825 (N_5825,N_341,N_61);
nor U5826 (N_5826,N_1137,N_2234);
or U5827 (N_5827,N_821,N_1262);
nand U5828 (N_5828,N_4961,N_3952);
nor U5829 (N_5829,N_4391,N_4873);
and U5830 (N_5830,N_2639,N_1215);
and U5831 (N_5831,N_1719,N_3160);
nor U5832 (N_5832,N_1598,N_3501);
nor U5833 (N_5833,N_1446,N_1731);
and U5834 (N_5834,N_1572,N_1362);
or U5835 (N_5835,N_2019,N_4260);
and U5836 (N_5836,N_4030,N_3289);
nand U5837 (N_5837,N_571,N_402);
or U5838 (N_5838,N_766,N_1398);
or U5839 (N_5839,N_828,N_1092);
nand U5840 (N_5840,N_4536,N_1858);
nand U5841 (N_5841,N_4125,N_444);
nor U5842 (N_5842,N_2356,N_616);
and U5843 (N_5843,N_4343,N_1695);
nor U5844 (N_5844,N_1683,N_867);
or U5845 (N_5845,N_3977,N_4615);
xnor U5846 (N_5846,N_712,N_1801);
nor U5847 (N_5847,N_2560,N_3976);
nand U5848 (N_5848,N_377,N_4782);
nor U5849 (N_5849,N_343,N_2528);
or U5850 (N_5850,N_622,N_2586);
nor U5851 (N_5851,N_652,N_4629);
nor U5852 (N_5852,N_3768,N_1299);
and U5853 (N_5853,N_3863,N_386);
nand U5854 (N_5854,N_2215,N_174);
nor U5855 (N_5855,N_2607,N_3918);
or U5856 (N_5856,N_449,N_3932);
or U5857 (N_5857,N_2301,N_274);
nor U5858 (N_5858,N_2976,N_2343);
or U5859 (N_5859,N_3995,N_2847);
and U5860 (N_5860,N_4170,N_4268);
or U5861 (N_5861,N_4819,N_1770);
nand U5862 (N_5862,N_3066,N_3620);
nor U5863 (N_5863,N_4275,N_3008);
nor U5864 (N_5864,N_4579,N_825);
nor U5865 (N_5865,N_4812,N_4222);
nand U5866 (N_5866,N_2442,N_1191);
or U5867 (N_5867,N_2068,N_4677);
nand U5868 (N_5868,N_4506,N_2970);
nor U5869 (N_5869,N_713,N_3250);
or U5870 (N_5870,N_1178,N_3201);
or U5871 (N_5871,N_3827,N_2022);
nand U5872 (N_5872,N_1230,N_1142);
or U5873 (N_5873,N_3119,N_1908);
and U5874 (N_5874,N_4912,N_1214);
or U5875 (N_5875,N_2314,N_1541);
nand U5876 (N_5876,N_2251,N_2912);
nor U5877 (N_5877,N_4177,N_1449);
and U5878 (N_5878,N_4110,N_1361);
nand U5879 (N_5879,N_2290,N_2082);
nand U5880 (N_5880,N_2051,N_4978);
xnor U5881 (N_5881,N_2119,N_2585);
nor U5882 (N_5882,N_4521,N_1513);
nand U5883 (N_5883,N_2397,N_1243);
nor U5884 (N_5884,N_3249,N_310);
nand U5885 (N_5885,N_1662,N_2307);
and U5886 (N_5886,N_1536,N_3523);
nand U5887 (N_5887,N_1975,N_787);
or U5888 (N_5888,N_4942,N_4680);
and U5889 (N_5889,N_2935,N_752);
nor U5890 (N_5890,N_1456,N_553);
nor U5891 (N_5891,N_1203,N_1009);
nand U5892 (N_5892,N_1562,N_401);
nor U5893 (N_5893,N_2796,N_1441);
or U5894 (N_5894,N_2723,N_3954);
nor U5895 (N_5895,N_4080,N_540);
nor U5896 (N_5896,N_3922,N_4618);
nand U5897 (N_5897,N_2814,N_4366);
nor U5898 (N_5898,N_2973,N_3169);
nand U5899 (N_5899,N_4249,N_4815);
or U5900 (N_5900,N_3372,N_4697);
or U5901 (N_5901,N_3774,N_4876);
and U5902 (N_5902,N_952,N_2376);
or U5903 (N_5903,N_479,N_3645);
nor U5904 (N_5904,N_337,N_3067);
and U5905 (N_5905,N_1740,N_1331);
nand U5906 (N_5906,N_111,N_408);
or U5907 (N_5907,N_185,N_2760);
nand U5908 (N_5908,N_4258,N_3648);
and U5909 (N_5909,N_380,N_2666);
and U5910 (N_5910,N_3753,N_4482);
and U5911 (N_5911,N_1226,N_919);
and U5912 (N_5912,N_3419,N_716);
xor U5913 (N_5913,N_3983,N_3626);
nand U5914 (N_5914,N_372,N_1627);
or U5915 (N_5915,N_4112,N_1970);
and U5916 (N_5916,N_1533,N_1599);
or U5917 (N_5917,N_4445,N_3139);
and U5918 (N_5918,N_1252,N_3805);
or U5919 (N_5919,N_2194,N_4138);
or U5920 (N_5920,N_720,N_567);
nand U5921 (N_5921,N_2594,N_4303);
xor U5922 (N_5922,N_223,N_1217);
and U5923 (N_5923,N_703,N_4212);
and U5924 (N_5924,N_642,N_2543);
nand U5925 (N_5925,N_1895,N_957);
nor U5926 (N_5926,N_2694,N_3946);
nor U5927 (N_5927,N_4166,N_2135);
or U5928 (N_5928,N_1922,N_1165);
xnor U5929 (N_5929,N_221,N_1406);
nor U5930 (N_5930,N_3894,N_4178);
and U5931 (N_5931,N_4148,N_4297);
nor U5932 (N_5932,N_1324,N_4447);
nand U5933 (N_5933,N_2116,N_4565);
nor U5934 (N_5934,N_1982,N_4818);
and U5935 (N_5935,N_244,N_2053);
xor U5936 (N_5936,N_582,N_697);
and U5937 (N_5937,N_1643,N_2507);
xor U5938 (N_5938,N_3321,N_1499);
or U5939 (N_5939,N_4977,N_13);
nor U5940 (N_5940,N_2893,N_1390);
or U5941 (N_5941,N_763,N_2758);
nand U5942 (N_5942,N_458,N_624);
and U5943 (N_5943,N_4402,N_1884);
nor U5944 (N_5944,N_2432,N_3632);
nand U5945 (N_5945,N_767,N_3051);
xor U5946 (N_5946,N_3092,N_2352);
or U5947 (N_5947,N_879,N_2191);
nor U5948 (N_5948,N_4433,N_114);
nor U5949 (N_5949,N_702,N_738);
or U5950 (N_5950,N_3657,N_3439);
and U5951 (N_5951,N_4168,N_2839);
or U5952 (N_5952,N_2624,N_2178);
and U5953 (N_5953,N_3597,N_4802);
nor U5954 (N_5954,N_4972,N_4119);
nor U5955 (N_5955,N_2378,N_4836);
or U5956 (N_5956,N_765,N_3341);
or U5957 (N_5957,N_2168,N_4714);
nor U5958 (N_5958,N_859,N_4089);
and U5959 (N_5959,N_2172,N_4171);
and U5960 (N_5960,N_4241,N_376);
or U5961 (N_5961,N_3830,N_133);
or U5962 (N_5962,N_1959,N_980);
nor U5963 (N_5963,N_2676,N_4189);
and U5964 (N_5964,N_921,N_4647);
and U5965 (N_5965,N_734,N_2161);
nand U5966 (N_5966,N_4439,N_545);
or U5967 (N_5967,N_440,N_4319);
xnor U5968 (N_5968,N_2773,N_3780);
and U5969 (N_5969,N_3948,N_645);
nor U5970 (N_5970,N_4952,N_1534);
nor U5971 (N_5971,N_4351,N_1967);
and U5972 (N_5972,N_762,N_3149);
nand U5973 (N_5973,N_2400,N_2408);
xor U5974 (N_5974,N_229,N_3215);
nor U5975 (N_5975,N_748,N_484);
nand U5976 (N_5976,N_1903,N_79);
or U5977 (N_5977,N_1930,N_2127);
xor U5978 (N_5978,N_145,N_3896);
nand U5979 (N_5979,N_1531,N_1653);
or U5980 (N_5980,N_4561,N_3654);
and U5981 (N_5981,N_3472,N_3140);
nor U5982 (N_5982,N_3881,N_2605);
nand U5983 (N_5983,N_3492,N_2843);
nand U5984 (N_5984,N_1904,N_4326);
or U5985 (N_5985,N_4738,N_773);
and U5986 (N_5986,N_4693,N_3337);
and U5987 (N_5987,N_2470,N_2026);
xnor U5988 (N_5988,N_1641,N_2745);
nand U5989 (N_5989,N_4617,N_801);
xnor U5990 (N_5990,N_2616,N_2198);
and U5991 (N_5991,N_4147,N_499);
nor U5992 (N_5992,N_3453,N_4309);
and U5993 (N_5993,N_3658,N_1485);
nor U5994 (N_5994,N_4907,N_1041);
nor U5995 (N_5995,N_3951,N_1436);
nor U5996 (N_5996,N_4612,N_4455);
and U5997 (N_5997,N_312,N_1304);
xor U5998 (N_5998,N_354,N_3081);
and U5999 (N_5999,N_4233,N_2654);
nand U6000 (N_6000,N_2844,N_2644);
nand U6001 (N_6001,N_3857,N_359);
nor U6002 (N_6002,N_836,N_1596);
nand U6003 (N_6003,N_4927,N_3364);
and U6004 (N_6004,N_1468,N_164);
nor U6005 (N_6005,N_785,N_4237);
or U6006 (N_6006,N_1949,N_3687);
or U6007 (N_6007,N_3279,N_3713);
nand U6008 (N_6008,N_1307,N_2138);
nand U6009 (N_6009,N_2690,N_2783);
nand U6010 (N_6010,N_2689,N_986);
and U6011 (N_6011,N_2291,N_4347);
xor U6012 (N_6012,N_1429,N_1422);
and U6013 (N_6013,N_4507,N_3807);
or U6014 (N_6014,N_1342,N_4294);
or U6015 (N_6015,N_3741,N_1480);
nor U6016 (N_6016,N_1297,N_3652);
or U6017 (N_6017,N_1730,N_429);
or U6018 (N_6018,N_2473,N_1798);
and U6019 (N_6019,N_110,N_124);
nor U6020 (N_6020,N_1549,N_2416);
xor U6021 (N_6021,N_2052,N_3477);
nand U6022 (N_6022,N_2906,N_3430);
nand U6023 (N_6023,N_592,N_1082);
nand U6024 (N_6024,N_3836,N_269);
xor U6025 (N_6025,N_2404,N_848);
nor U6026 (N_6026,N_399,N_4123);
or U6027 (N_6027,N_1433,N_2380);
or U6028 (N_6028,N_4475,N_777);
or U6029 (N_6029,N_1529,N_994);
nor U6030 (N_6030,N_2769,N_2958);
nand U6031 (N_6031,N_2842,N_3668);
nand U6032 (N_6032,N_4775,N_2118);
or U6033 (N_6033,N_1503,N_1005);
nor U6034 (N_6034,N_1870,N_4333);
nor U6035 (N_6035,N_1301,N_1370);
nand U6036 (N_6036,N_3546,N_1765);
and U6037 (N_6037,N_2583,N_4837);
or U6038 (N_6038,N_2010,N_256);
and U6039 (N_6039,N_4205,N_550);
xor U6040 (N_6040,N_3252,N_55);
and U6041 (N_6041,N_814,N_4719);
nand U6042 (N_6042,N_3489,N_2833);
nand U6043 (N_6043,N_4575,N_36);
or U6044 (N_6044,N_1384,N_3582);
nand U6045 (N_6045,N_292,N_2033);
nand U6046 (N_6046,N_3355,N_2513);
nor U6047 (N_6047,N_2683,N_1910);
nor U6048 (N_6048,N_1956,N_197);
and U6049 (N_6049,N_2185,N_3860);
nor U6050 (N_6050,N_4230,N_278);
nand U6051 (N_6051,N_799,N_3040);
or U6052 (N_6052,N_521,N_1393);
nor U6053 (N_6053,N_407,N_664);
or U6054 (N_6054,N_1576,N_250);
nor U6055 (N_6055,N_2158,N_2930);
nor U6056 (N_6056,N_3403,N_2857);
or U6057 (N_6057,N_2042,N_820);
or U6058 (N_6058,N_209,N_678);
and U6059 (N_6059,N_3032,N_33);
or U6060 (N_6060,N_1281,N_1764);
nand U6061 (N_6061,N_1329,N_2938);
nand U6062 (N_6062,N_2296,N_3499);
nand U6063 (N_6063,N_1717,N_125);
and U6064 (N_6064,N_3683,N_3784);
and U6065 (N_6065,N_4631,N_3837);
nor U6066 (N_6066,N_1002,N_4984);
nand U6067 (N_6067,N_2146,N_1138);
nand U6068 (N_6068,N_727,N_559);
nand U6069 (N_6069,N_4428,N_4289);
nor U6070 (N_6070,N_3893,N_2575);
or U6071 (N_6071,N_827,N_4259);
or U6072 (N_6072,N_2066,N_3084);
nor U6073 (N_6073,N_4041,N_1985);
or U6074 (N_6074,N_239,N_1860);
nor U6075 (N_6075,N_283,N_2197);
xor U6076 (N_6076,N_2186,N_2955);
nand U6077 (N_6077,N_4198,N_4526);
nand U6078 (N_6078,N_2262,N_1863);
and U6079 (N_6079,N_4569,N_3123);
and U6080 (N_6080,N_459,N_3460);
xnor U6081 (N_6081,N_4503,N_4945);
or U6082 (N_6082,N_4881,N_4393);
xnor U6083 (N_6083,N_1698,N_4847);
or U6084 (N_6084,N_1355,N_2087);
and U6085 (N_6085,N_2261,N_1833);
nand U6086 (N_6086,N_3905,N_371);
or U6087 (N_6087,N_1955,N_970);
nand U6088 (N_6088,N_0,N_1639);
xnor U6089 (N_6089,N_3198,N_1520);
nor U6090 (N_6090,N_1703,N_4674);
nand U6091 (N_6091,N_4485,N_3763);
nand U6092 (N_6092,N_2142,N_2207);
and U6093 (N_6093,N_2405,N_1912);
or U6094 (N_6094,N_3769,N_122);
and U6095 (N_6095,N_1737,N_4277);
nor U6096 (N_6096,N_772,N_3306);
nand U6097 (N_6097,N_1209,N_2336);
nor U6098 (N_6098,N_4886,N_2667);
nor U6099 (N_6099,N_1221,N_3475);
or U6100 (N_6100,N_1124,N_841);
nor U6101 (N_6101,N_4669,N_4091);
nor U6102 (N_6102,N_3515,N_4270);
nand U6103 (N_6103,N_3217,N_433);
nand U6104 (N_6104,N_1935,N_2947);
and U6105 (N_6105,N_2580,N_2237);
or U6106 (N_6106,N_4397,N_4528);
nor U6107 (N_6107,N_2827,N_3544);
nor U6108 (N_6108,N_3711,N_1495);
nor U6109 (N_6109,N_832,N_2277);
nand U6110 (N_6110,N_1056,N_1350);
and U6111 (N_6111,N_3207,N_478);
nand U6112 (N_6112,N_3340,N_868);
and U6113 (N_6113,N_2611,N_2498);
nand U6114 (N_6114,N_1454,N_3787);
nor U6115 (N_6115,N_2508,N_525);
nand U6116 (N_6116,N_2657,N_2747);
nand U6117 (N_6117,N_2120,N_153);
or U6118 (N_6118,N_1081,N_3791);
or U6119 (N_6119,N_128,N_3754);
nand U6120 (N_6120,N_1060,N_4238);
or U6121 (N_6121,N_2617,N_971);
nand U6122 (N_6122,N_2046,N_737);
nor U6123 (N_6123,N_811,N_4776);
xnor U6124 (N_6124,N_3267,N_3027);
and U6125 (N_6125,N_3468,N_4958);
xnor U6126 (N_6126,N_276,N_4192);
or U6127 (N_6127,N_3190,N_4767);
xnor U6128 (N_6128,N_4096,N_3199);
and U6129 (N_6129,N_4700,N_4874);
nand U6130 (N_6130,N_3104,N_2128);
nand U6131 (N_6131,N_2279,N_262);
or U6132 (N_6132,N_2549,N_90);
xor U6133 (N_6133,N_2409,N_4114);
nand U6134 (N_6134,N_3212,N_3947);
nor U6135 (N_6135,N_2569,N_1655);
nand U6136 (N_6136,N_4694,N_2504);
or U6137 (N_6137,N_1451,N_2904);
xnor U6138 (N_6138,N_2264,N_4279);
nor U6139 (N_6139,N_263,N_1049);
and U6140 (N_6140,N_191,N_38);
nor U6141 (N_6141,N_1642,N_76);
nand U6142 (N_6142,N_1626,N_4269);
nor U6143 (N_6143,N_3033,N_2495);
or U6144 (N_6144,N_2238,N_18);
nand U6145 (N_6145,N_252,N_4998);
or U6146 (N_6146,N_430,N_2455);
or U6147 (N_6147,N_2808,N_4034);
nand U6148 (N_6148,N_4546,N_1320);
nor U6149 (N_6149,N_2351,N_4395);
or U6150 (N_6150,N_3972,N_4145);
xor U6151 (N_6151,N_2284,N_3243);
or U6152 (N_6152,N_875,N_4596);
xor U6153 (N_6153,N_2848,N_2340);
nand U6154 (N_6154,N_1697,N_4441);
and U6155 (N_6155,N_3278,N_1426);
nand U6156 (N_6156,N_4924,N_4202);
or U6157 (N_6157,N_4768,N_2609);
and U6158 (N_6158,N_4739,N_1080);
nand U6159 (N_6159,N_551,N_2098);
xnor U6160 (N_6160,N_2878,N_4855);
nor U6161 (N_6161,N_3173,N_983);
xor U6162 (N_6162,N_4994,N_3821);
and U6163 (N_6163,N_706,N_3912);
nor U6164 (N_6164,N_2910,N_3998);
nand U6165 (N_6165,N_2303,N_3945);
nor U6166 (N_6166,N_2379,N_4527);
and U6167 (N_6167,N_849,N_195);
nor U6168 (N_6168,N_412,N_1020);
nand U6169 (N_6169,N_3113,N_4150);
nand U6170 (N_6170,N_1267,N_4807);
and U6171 (N_6171,N_406,N_154);
nand U6172 (N_6172,N_2028,N_465);
or U6173 (N_6173,N_2035,N_3329);
or U6174 (N_6174,N_4345,N_8);
and U6175 (N_6175,N_3451,N_2085);
and U6176 (N_6176,N_2192,N_3485);
and U6177 (N_6177,N_3733,N_613);
nor U6178 (N_6178,N_48,N_3121);
nor U6179 (N_6179,N_1408,N_1760);
nand U6180 (N_6180,N_3520,N_2169);
xnor U6181 (N_6181,N_304,N_805);
and U6182 (N_6182,N_2803,N_2576);
nand U6183 (N_6183,N_2899,N_4878);
nor U6184 (N_6184,N_232,N_2673);
nor U6185 (N_6185,N_4788,N_4380);
and U6186 (N_6186,N_1766,N_2206);
nor U6187 (N_6187,N_4349,N_89);
nor U6188 (N_6188,N_326,N_3039);
nor U6189 (N_6189,N_1278,N_2663);
or U6190 (N_6190,N_3214,N_4173);
or U6191 (N_6191,N_4427,N_3898);
nand U6192 (N_6192,N_3188,N_3017);
nor U6193 (N_6193,N_1052,N_1302);
nor U6194 (N_6194,N_1992,N_3087);
and U6195 (N_6195,N_4784,N_689);
nand U6196 (N_6196,N_640,N_3519);
and U6197 (N_6197,N_4518,N_3474);
nor U6198 (N_6198,N_781,N_1851);
nand U6199 (N_6199,N_1067,N_4322);
nand U6200 (N_6200,N_3486,N_3861);
and U6201 (N_6201,N_3397,N_4265);
xnor U6202 (N_6202,N_3099,N_3507);
nand U6203 (N_6203,N_1815,N_4392);
and U6204 (N_6204,N_3464,N_2991);
and U6205 (N_6205,N_1427,N_4897);
and U6206 (N_6206,N_3437,N_1901);
nor U6207 (N_6207,N_45,N_3939);
nand U6208 (N_6208,N_1348,N_228);
nor U6209 (N_6209,N_3035,N_1876);
and U6210 (N_6210,N_1162,N_2629);
xor U6211 (N_6211,N_1106,N_4274);
and U6212 (N_6212,N_4436,N_1947);
nand U6213 (N_6213,N_3514,N_3914);
nor U6214 (N_6214,N_2134,N_1273);
and U6215 (N_6215,N_3969,N_4661);
and U6216 (N_6216,N_3688,N_446);
or U6217 (N_6217,N_2254,N_331);
and U6218 (N_6218,N_594,N_4191);
nand U6219 (N_6219,N_3132,N_2211);
or U6220 (N_6220,N_2846,N_3913);
nand U6221 (N_6221,N_596,N_1785);
and U6222 (N_6222,N_4544,N_199);
and U6223 (N_6223,N_1391,N_675);
xnor U6224 (N_6224,N_4547,N_141);
or U6225 (N_6225,N_217,N_699);
nor U6226 (N_6226,N_4474,N_3088);
nand U6227 (N_6227,N_4043,N_162);
nand U6228 (N_6228,N_2289,N_4301);
and U6229 (N_6229,N_843,N_3570);
nor U6230 (N_6230,N_3812,N_887);
or U6231 (N_6231,N_3749,N_1916);
or U6232 (N_6232,N_736,N_683);
nand U6233 (N_6233,N_784,N_143);
or U6234 (N_6234,N_4757,N_267);
and U6235 (N_6235,N_2210,N_83);
and U6236 (N_6236,N_648,N_1182);
or U6237 (N_6237,N_2787,N_383);
xor U6238 (N_6238,N_1042,N_2479);
or U6239 (N_6239,N_2344,N_3219);
nor U6240 (N_6240,N_1810,N_838);
and U6241 (N_6241,N_3931,N_1588);
and U6242 (N_6242,N_1941,N_3845);
or U6243 (N_6243,N_422,N_235);
or U6244 (N_6244,N_3272,N_991);
or U6245 (N_6245,N_4773,N_1962);
nand U6246 (N_6246,N_2089,N_680);
and U6247 (N_6247,N_1816,N_1972);
or U6248 (N_6248,N_4174,N_674);
xor U6249 (N_6249,N_163,N_3614);
and U6250 (N_6250,N_526,N_505);
or U6251 (N_6251,N_2348,N_3644);
nand U6252 (N_6252,N_3680,N_2013);
nor U6253 (N_6253,N_668,N_4811);
and U6254 (N_6254,N_1018,N_2821);
nor U6255 (N_6255,N_3467,N_2002);
nor U6256 (N_6256,N_1793,N_4826);
and U6257 (N_6257,N_722,N_3572);
and U6258 (N_6258,N_1120,N_910);
nor U6259 (N_6259,N_3111,N_3569);
or U6260 (N_6260,N_944,N_677);
or U6261 (N_6261,N_2699,N_1409);
or U6262 (N_6262,N_1295,N_3890);
and U6263 (N_6263,N_2103,N_4139);
nand U6264 (N_6264,N_4583,N_4905);
nor U6265 (N_6265,N_1542,N_1220);
or U6266 (N_6266,N_4887,N_4650);
nor U6267 (N_6267,N_2922,N_2588);
nor U6268 (N_6268,N_4430,N_3389);
nand U6269 (N_6269,N_2630,N_4658);
xnor U6270 (N_6270,N_611,N_519);
or U6271 (N_6271,N_1656,N_942);
nor U6272 (N_6272,N_1806,N_576);
nor U6273 (N_6273,N_207,N_3034);
or U6274 (N_6274,N_3046,N_1153);
xnor U6275 (N_6275,N_4036,N_1474);
nor U6276 (N_6276,N_2427,N_4735);
and U6277 (N_6277,N_1029,N_2898);
nand U6278 (N_6278,N_4031,N_3986);
nor U6279 (N_6279,N_2230,N_73);
nand U6280 (N_6280,N_4386,N_2677);
nand U6281 (N_6281,N_301,N_4383);
nand U6282 (N_6282,N_4127,N_2398);
or U6283 (N_6283,N_4155,N_4008);
nor U6284 (N_6284,N_1497,N_379);
nand U6285 (N_6285,N_3283,N_4470);
or U6286 (N_6286,N_750,N_4417);
and U6287 (N_6287,N_1973,N_3817);
nand U6288 (N_6288,N_1457,N_3400);
nor U6289 (N_6289,N_4321,N_4710);
nor U6290 (N_6290,N_2298,N_3443);
and U6291 (N_6291,N_155,N_2247);
or U6292 (N_6292,N_3900,N_1664);
nand U6293 (N_6293,N_4509,N_4872);
and U6294 (N_6294,N_1634,N_4666);
nand U6295 (N_6295,N_4580,N_1245);
and U6296 (N_6296,N_2602,N_2283);
xnor U6297 (N_6297,N_1943,N_4257);
or U6298 (N_6298,N_3953,N_1286);
or U6299 (N_6299,N_2422,N_4494);
or U6300 (N_6300,N_4385,N_202);
nor U6301 (N_6301,N_2951,N_3495);
and U6302 (N_6302,N_2897,N_4610);
nor U6303 (N_6303,N_241,N_4637);
xnor U6304 (N_6304,N_3227,N_3247);
nor U6305 (N_6305,N_4285,N_4262);
or U6306 (N_6306,N_2520,N_2547);
nor U6307 (N_6307,N_2193,N_2096);
or U6308 (N_6308,N_948,N_3697);
or U6309 (N_6309,N_4713,N_2802);
or U6310 (N_6310,N_2465,N_1274);
and U6311 (N_6311,N_4371,N_2968);
nand U6312 (N_6312,N_4760,N_1651);
nor U6313 (N_6313,N_4418,N_1172);
and U6314 (N_6314,N_1400,N_1727);
or U6315 (N_6315,N_4460,N_3324);
nand U6316 (N_6316,N_1702,N_365);
or U6317 (N_6317,N_2050,N_534);
and U6318 (N_6318,N_2792,N_1321);
nand U6319 (N_6319,N_3425,N_1819);
nand U6320 (N_6320,N_254,N_115);
nand U6321 (N_6321,N_1853,N_2716);
or U6322 (N_6322,N_1300,N_4997);
nor U6323 (N_6323,N_1752,N_3233);
or U6324 (N_6324,N_4200,N_1538);
nand U6325 (N_6325,N_4880,N_1946);
nor U6326 (N_6326,N_3796,N_3964);
and U6327 (N_6327,N_4974,N_119);
nand U6328 (N_6328,N_3304,N_1368);
and U6329 (N_6329,N_3975,N_899);
or U6330 (N_6330,N_4706,N_3822);
nor U6331 (N_6331,N_2998,N_4312);
nand U6332 (N_6332,N_3901,N_3651);
and U6333 (N_6333,N_1613,N_1799);
and U6334 (N_6334,N_587,N_1814);
nand U6335 (N_6335,N_4765,N_1886);
nor U6336 (N_6336,N_4083,N_370);
nand U6337 (N_6337,N_4467,N_293);
nand U6338 (N_6338,N_2370,N_309);
or U6339 (N_6339,N_1309,N_1289);
nor U6340 (N_6340,N_1280,N_3170);
or U6341 (N_6341,N_959,N_3985);
xnor U6342 (N_6342,N_2441,N_1517);
and U6343 (N_6343,N_2061,N_3758);
nand U6344 (N_6344,N_2820,N_682);
and U6345 (N_6345,N_2083,N_3024);
and U6346 (N_6346,N_2828,N_1213);
nand U6347 (N_6347,N_543,N_1688);
and U6348 (N_6348,N_2023,N_1647);
nand U6349 (N_6349,N_3145,N_2125);
and U6350 (N_6350,N_3010,N_1741);
nor U6351 (N_6351,N_1229,N_4232);
or U6352 (N_6352,N_714,N_2830);
or U6353 (N_6353,N_134,N_4689);
nor U6354 (N_6354,N_3205,N_4728);
xor U6355 (N_6355,N_180,N_4888);
nor U6356 (N_6356,N_3351,N_939);
nand U6357 (N_6357,N_2145,N_152);
nor U6358 (N_6358,N_4943,N_3872);
nor U6359 (N_6359,N_2020,N_4278);
or U6360 (N_6360,N_467,N_1775);
nand U6361 (N_6361,N_1813,N_4306);
and U6362 (N_6362,N_3663,N_3909);
or U6363 (N_6363,N_958,N_665);
or U6364 (N_6364,N_3775,N_666);
or U6365 (N_6365,N_1233,N_4452);
or U6366 (N_6366,N_4753,N_2043);
xor U6367 (N_6367,N_1284,N_3186);
xor U6368 (N_6368,N_4248,N_561);
nor U6369 (N_6369,N_165,N_1988);
nand U6370 (N_6370,N_497,N_1768);
xnor U6371 (N_6371,N_307,N_4367);
nor U6372 (N_6372,N_2931,N_731);
and U6373 (N_6373,N_844,N_4152);
xor U6374 (N_6374,N_101,N_1892);
and U6375 (N_6375,N_135,N_4986);
nand U6376 (N_6376,N_2867,N_39);
xnor U6377 (N_6377,N_1443,N_1758);
nand U6378 (N_6378,N_641,N_4894);
and U6379 (N_6379,N_1044,N_846);
nand U6380 (N_6380,N_306,N_2718);
nand U6381 (N_6381,N_537,N_3322);
and U6382 (N_6382,N_3548,N_1587);
nand U6383 (N_6383,N_3610,N_3461);
nand U6384 (N_6384,N_4950,N_3736);
or U6385 (N_6385,N_2199,N_3023);
xnor U6386 (N_6386,N_3533,N_4104);
or U6387 (N_6387,N_920,N_3518);
nor U6388 (N_6388,N_4869,N_2311);
or U6389 (N_6389,N_3706,N_4895);
or U6390 (N_6390,N_1974,N_3080);
nor U6391 (N_6391,N_852,N_2338);
nor U6392 (N_6392,N_1500,N_2868);
nor U6393 (N_6393,N_319,N_2559);
nor U6394 (N_6394,N_1900,N_1432);
and U6395 (N_6395,N_4664,N_1604);
and U6396 (N_6396,N_491,N_3650);
or U6397 (N_6397,N_3392,N_4384);
and U6398 (N_6398,N_4044,N_1885);
nor U6399 (N_6399,N_2573,N_966);
and U6400 (N_6400,N_1791,N_4196);
nand U6401 (N_6401,N_4551,N_855);
and U6402 (N_6402,N_1658,N_1125);
and U6403 (N_6403,N_3649,N_918);
nor U6404 (N_6404,N_1535,N_22);
nand U6405 (N_6405,N_2055,N_54);
nor U6406 (N_6406,N_739,N_2850);
and U6407 (N_6407,N_671,N_987);
nor U6408 (N_6408,N_4644,N_2032);
nand U6409 (N_6409,N_2866,N_1453);
or U6410 (N_6410,N_2710,N_4414);
and U6411 (N_6411,N_3465,N_3449);
or U6412 (N_6412,N_4915,N_1995);
nor U6413 (N_6413,N_4805,N_985);
or U6414 (N_6414,N_1753,N_2817);
nor U6415 (N_6415,N_1981,N_3618);
nor U6416 (N_6416,N_3696,N_300);
or U6417 (N_6417,N_2003,N_3852);
nand U6418 (N_6418,N_3653,N_1486);
or U6419 (N_6419,N_3174,N_66);
or U6420 (N_6420,N_1341,N_16);
and U6421 (N_6421,N_3944,N_1784);
and U6422 (N_6422,N_2481,N_3248);
or U6423 (N_6423,N_35,N_432);
nand U6424 (N_6424,N_2036,N_2274);
or U6425 (N_6425,N_4621,N_47);
and U6426 (N_6426,N_914,N_1004);
nor U6427 (N_6427,N_873,N_2406);
nor U6428 (N_6428,N_1379,N_1561);
nor U6429 (N_6429,N_3416,N_3730);
and U6430 (N_6430,N_4722,N_633);
or U6431 (N_6431,N_1917,N_1867);
nor U6432 (N_6432,N_2661,N_3936);
or U6433 (N_6433,N_3253,N_573);
and U6434 (N_6434,N_4828,N_2292);
or U6435 (N_6435,N_2287,N_853);
xnor U6436 (N_6436,N_998,N_552);
nand U6437 (N_6437,N_1070,N_1119);
xnor U6438 (N_6438,N_2377,N_305);
or U6439 (N_6439,N_1595,N_4000);
xnor U6440 (N_6440,N_397,N_3301);
nand U6441 (N_6441,N_531,N_2730);
or U6442 (N_6442,N_4857,N_4971);
or U6443 (N_6443,N_4796,N_940);
xnor U6444 (N_6444,N_4908,N_4608);
nor U6445 (N_6445,N_1223,N_243);
nor U6446 (N_6446,N_1017,N_2851);
nor U6447 (N_6447,N_1696,N_4925);
and U6448 (N_6448,N_2480,N_2387);
and U6449 (N_6449,N_3655,N_2501);
or U6450 (N_6450,N_2392,N_471);
nand U6451 (N_6451,N_127,N_672);
and U6452 (N_6452,N_466,N_3231);
and U6453 (N_6453,N_963,N_3806);
nor U6454 (N_6454,N_4201,N_4311);
or U6455 (N_6455,N_2286,N_2349);
nand U6456 (N_6456,N_2485,N_896);
and U6457 (N_6457,N_1276,N_4480);
and U6458 (N_6458,N_4350,N_4235);
or U6459 (N_6459,N_3924,N_4163);
nor U6460 (N_6460,N_529,N_2601);
or U6461 (N_6461,N_725,N_3970);
nand U6462 (N_6462,N_1923,N_2367);
nor U6463 (N_6463,N_3793,N_425);
nand U6464 (N_6464,N_861,N_2294);
nand U6465 (N_6465,N_2887,N_501);
and U6466 (N_6466,N_3068,N_3679);
nor U6467 (N_6467,N_1636,N_3043);
and U6468 (N_6468,N_1679,N_3795);
xnor U6469 (N_6469,N_3547,N_1216);
nand U6470 (N_6470,N_2477,N_2890);
nand U6471 (N_6471,N_2885,N_3288);
nand U6472 (N_6472,N_4143,N_4554);
or U6473 (N_6473,N_368,N_1864);
nor U6474 (N_6474,N_3968,N_94);
nor U6475 (N_6475,N_4730,N_662);
and U6476 (N_6476,N_4896,N_3230);
xnor U6477 (N_6477,N_1236,N_41);
or U6478 (N_6478,N_4840,N_4717);
nand U6479 (N_6479,N_4600,N_1033);
nor U6480 (N_6480,N_637,N_490);
and U6481 (N_6481,N_1071,N_182);
and U6482 (N_6482,N_142,N_4772);
nand U6483 (N_6483,N_3767,N_3090);
nand U6484 (N_6484,N_1007,N_4861);
nor U6485 (N_6485,N_3583,N_4239);
and U6486 (N_6486,N_1043,N_3907);
nor U6487 (N_6487,N_635,N_1909);
and U6488 (N_6488,N_1431,N_3517);
nor U6489 (N_6489,N_4504,N_1055);
xnor U6490 (N_6490,N_4853,N_779);
xor U6491 (N_6491,N_4866,N_4524);
nor U6492 (N_6492,N_4223,N_137);
nand U6493 (N_6493,N_3538,N_3152);
nor U6494 (N_6494,N_690,N_4293);
xnor U6495 (N_6495,N_1577,N_2153);
nand U6496 (N_6496,N_3239,N_318);
nor U6497 (N_6497,N_2900,N_512);
and U6498 (N_6498,N_3260,N_565);
nor U6499 (N_6499,N_3369,N_1150);
and U6500 (N_6500,N_579,N_2854);
nor U6501 (N_6501,N_78,N_1990);
and U6502 (N_6502,N_2424,N_4588);
or U6503 (N_6503,N_4523,N_1676);
nor U6504 (N_6504,N_895,N_2524);
or U6505 (N_6505,N_974,N_3055);
xnor U6506 (N_6506,N_3182,N_1460);
nand U6507 (N_6507,N_120,N_183);
and U6508 (N_6508,N_4512,N_311);
and U6509 (N_6509,N_1285,N_793);
and U6510 (N_6510,N_927,N_4708);
nand U6511 (N_6511,N_964,N_3194);
nand U6512 (N_6512,N_1837,N_1255);
or U6513 (N_6513,N_106,N_1346);
and U6514 (N_6514,N_1349,N_25);
or U6515 (N_6515,N_646,N_3166);
and U6516 (N_6516,N_3330,N_242);
and U6517 (N_6517,N_291,N_3314);
nor U6518 (N_6518,N_2109,N_1148);
nor U6519 (N_6519,N_2999,N_1602);
nand U6520 (N_6520,N_4654,N_2966);
and U6521 (N_6521,N_366,N_2916);
or U6522 (N_6522,N_2895,N_3380);
and U6523 (N_6523,N_4525,N_956);
and U6524 (N_6524,N_4951,N_4244);
xor U6525 (N_6525,N_4195,N_4132);
and U6526 (N_6526,N_284,N_3895);
nand U6527 (N_6527,N_32,N_2832);
nand U6528 (N_6528,N_3509,N_4688);
nand U6529 (N_6529,N_2600,N_2330);
nand U6530 (N_6530,N_2725,N_1847);
nand U6531 (N_6531,N_4146,N_1063);
and U6532 (N_6532,N_2675,N_4011);
nor U6533 (N_6533,N_1550,N_1195);
and U6534 (N_6534,N_4340,N_1850);
xor U6535 (N_6535,N_457,N_1771);
or U6536 (N_6536,N_4946,N_1571);
nor U6537 (N_6537,N_2965,N_925);
nor U6538 (N_6538,N_4048,N_909);
nand U6539 (N_6539,N_2510,N_1759);
or U6540 (N_6540,N_1835,N_3126);
nor U6541 (N_6541,N_298,N_257);
or U6542 (N_6542,N_1684,N_3853);
nor U6543 (N_6543,N_560,N_3963);
and U6544 (N_6544,N_2059,N_4673);
and U6545 (N_6545,N_2985,N_1211);
and U6546 (N_6546,N_416,N_650);
nand U6547 (N_6547,N_3551,N_3155);
or U6548 (N_6548,N_2536,N_2838);
nand U6549 (N_6549,N_3832,N_1754);
nor U6550 (N_6550,N_1419,N_1290);
xnor U6551 (N_6551,N_4962,N_2245);
nand U6552 (N_6552,N_4320,N_1675);
and U6553 (N_6553,N_3665,N_517);
nand U6554 (N_6554,N_2263,N_1723);
nand U6555 (N_6555,N_3888,N_679);
and U6556 (N_6556,N_4849,N_4798);
nor U6557 (N_6557,N_4082,N_3444);
nor U6558 (N_6558,N_1254,N_2776);
nor U6559 (N_6559,N_4108,N_2001);
xnor U6560 (N_6560,N_4038,N_4015);
nor U6561 (N_6561,N_1950,N_198);
or U6562 (N_6562,N_212,N_1452);
nor U6563 (N_6563,N_2360,N_1458);
and U6564 (N_6564,N_2577,N_487);
nand U6565 (N_6565,N_320,N_4370);
or U6566 (N_6566,N_29,N_2269);
xor U6567 (N_6567,N_4959,N_4352);
and U6568 (N_6568,N_280,N_4920);
nand U6569 (N_6569,N_2655,N_4560);
xnor U6570 (N_6570,N_757,N_4316);
nor U6571 (N_6571,N_1112,N_116);
nand U6572 (N_6572,N_3185,N_4364);
nand U6573 (N_6573,N_2228,N_2170);
nor U6574 (N_6574,N_3094,N_797);
nor U6575 (N_6575,N_3702,N_1396);
nor U6576 (N_6576,N_4508,N_1098);
xor U6577 (N_6577,N_1133,N_2672);
nor U6578 (N_6578,N_3530,N_1258);
nor U6579 (N_6579,N_2428,N_3527);
nor U6580 (N_6580,N_4099,N_1471);
nor U6581 (N_6581,N_409,N_1504);
nand U6582 (N_6582,N_3136,N_1927);
or U6583 (N_6583,N_696,N_2570);
xnor U6584 (N_6584,N_1334,N_1849);
or U6585 (N_6585,N_4390,N_4514);
xnor U6586 (N_6586,N_3280,N_589);
or U6587 (N_6587,N_4354,N_3348);
or U6588 (N_6588,N_2224,N_3362);
nor U6589 (N_6589,N_3107,N_3719);
nand U6590 (N_6590,N_176,N_2567);
nand U6591 (N_6591,N_378,N_2984);
nor U6592 (N_6592,N_1951,N_96);
nand U6593 (N_6593,N_542,N_2806);
xor U6594 (N_6594,N_1127,N_4779);
and U6595 (N_6595,N_411,N_3670);
nor U6596 (N_6596,N_2302,N_1762);
nor U6597 (N_6597,N_3661,N_3426);
nor U6598 (N_6598,N_541,N_4489);
or U6599 (N_6599,N_1157,N_2959);
or U6600 (N_6600,N_2798,N_2067);
nand U6601 (N_6601,N_1169,N_2994);
or U6602 (N_6602,N_4073,N_621);
nor U6603 (N_6603,N_1160,N_2164);
xor U6604 (N_6604,N_2708,N_584);
nand U6605 (N_6605,N_2275,N_3598);
nand U6606 (N_6606,N_2651,N_3825);
and U6607 (N_6607,N_4012,N_4013);
and U6608 (N_6608,N_1498,N_3765);
nand U6609 (N_6609,N_1193,N_3345);
or U6610 (N_6610,N_4298,N_3142);
nand U6611 (N_6611,N_1843,N_4749);
and U6612 (N_6612,N_4917,N_1879);
xor U6613 (N_6613,N_3130,N_3601);
nand U6614 (N_6614,N_2454,N_2521);
or U6615 (N_6615,N_4415,N_1525);
or U6616 (N_6616,N_1135,N_3522);
xnor U6617 (N_6617,N_234,N_107);
and U6618 (N_6618,N_502,N_1386);
or U6619 (N_6619,N_1579,N_4889);
nand U6620 (N_6620,N_1608,N_4919);
or U6621 (N_6621,N_3865,N_220);
nor U6622 (N_6622,N_3206,N_4302);
and U6623 (N_6623,N_3490,N_3106);
or U6624 (N_6624,N_1805,N_1532);
xor U6625 (N_6625,N_1600,N_2633);
nand U6626 (N_6626,N_2662,N_488);
nor U6627 (N_6627,N_2171,N_556);
and U6628 (N_6628,N_2309,N_3994);
and U6629 (N_6629,N_285,N_1404);
nand U6630 (N_6630,N_373,N_2104);
and U6631 (N_6631,N_4420,N_1693);
xnor U6632 (N_6632,N_3335,N_3701);
and U6633 (N_6633,N_4701,N_2232);
xor U6634 (N_6634,N_281,N_840);
or U6635 (N_6635,N_4808,N_1745);
and U6636 (N_6636,N_2049,N_4813);
nor U6637 (N_6637,N_4064,N_599);
and U6638 (N_6638,N_4078,N_2925);
or U6639 (N_6639,N_1663,N_1116);
xnor U6640 (N_6640,N_1305,N_1268);
nor U6641 (N_6641,N_4741,N_2884);
or U6642 (N_6642,N_2205,N_172);
and U6643 (N_6643,N_3302,N_2642);
nand U6644 (N_6644,N_3584,N_1414);
or U6645 (N_6645,N_2112,N_4841);
and U6646 (N_6646,N_4829,N_3993);
nand U6647 (N_6647,N_3606,N_168);
or U6648 (N_6648,N_2299,N_3098);
or U6649 (N_6649,N_638,N_4055);
nand U6650 (N_6650,N_2434,N_3005);
nor U6651 (N_6651,N_3624,N_2467);
nand U6652 (N_6652,N_3635,N_150);
nand U6653 (N_6653,N_558,N_1623);
and U6654 (N_6654,N_1357,N_857);
and U6655 (N_6655,N_4913,N_3037);
and U6656 (N_6656,N_3928,N_1294);
or U6657 (N_6657,N_3750,N_4468);
or U6658 (N_6658,N_4218,N_1483);
or U6659 (N_6659,N_3925,N_1971);
or U6660 (N_6660,N_2997,N_118);
and U6661 (N_6661,N_4956,N_4359);
or U6662 (N_6662,N_31,N_1644);
and U6663 (N_6663,N_4273,N_2011);
and U6664 (N_6664,N_4118,N_3636);
nand U6665 (N_6665,N_1313,N_4002);
nor U6666 (N_6666,N_2869,N_2278);
or U6667 (N_6667,N_4548,N_4242);
xnor U6668 (N_6668,N_2761,N_2591);
or U6669 (N_6669,N_3877,N_4247);
nor U6670 (N_6670,N_4785,N_3338);
and U6671 (N_6671,N_112,N_3022);
nand U6672 (N_6672,N_121,N_4774);
nor U6673 (N_6673,N_3483,N_1840);
nor U6674 (N_6674,N_2154,N_3956);
xnor U6675 (N_6675,N_655,N_4056);
nor U6676 (N_6676,N_2078,N_4407);
xnor U6677 (N_6677,N_695,N_4219);
or U6678 (N_6678,N_673,N_3074);
or U6679 (N_6679,N_2748,N_4151);
and U6680 (N_6680,N_92,N_4865);
nand U6681 (N_6681,N_2021,N_1364);
and U6682 (N_6682,N_872,N_3480);
and U6683 (N_6683,N_1083,N_726);
xor U6684 (N_6684,N_1558,N_2395);
xor U6685 (N_6685,N_4799,N_3973);
nor U6686 (N_6686,N_3531,N_2678);
nand U6687 (N_6687,N_1721,N_1096);
nor U6688 (N_6688,N_3326,N_1751);
nand U6689 (N_6689,N_456,N_3421);
nand U6690 (N_6690,N_700,N_4931);
nor U6691 (N_6691,N_931,N_4106);
nor U6692 (N_6692,N_3405,N_1177);
nand U6693 (N_6693,N_3797,N_1105);
and U6694 (N_6694,N_3637,N_3381);
or U6695 (N_6695,N_2558,N_938);
nor U6696 (N_6696,N_2324,N_2529);
xnor U6697 (N_6697,N_4059,N_4955);
and U6698 (N_6698,N_3276,N_3709);
xor U6699 (N_6699,N_791,N_3143);
nand U6700 (N_6700,N_4824,N_2845);
xor U6701 (N_6701,N_2415,N_824);
nor U6702 (N_6702,N_3286,N_1861);
nor U6703 (N_6703,N_2174,N_4571);
nor U6704 (N_6704,N_949,N_746);
and U6705 (N_6705,N_330,N_3641);
nor U6706 (N_6706,N_1487,N_2512);
nand U6707 (N_6707,N_1030,N_4885);
nand U6708 (N_6708,N_698,N_93);
nand U6709 (N_6709,N_266,N_4310);
or U6710 (N_6710,N_1957,N_3815);
nand U6711 (N_6711,N_2915,N_360);
nor U6712 (N_6712,N_2598,N_4858);
and U6713 (N_6713,N_431,N_2226);
and U6714 (N_6714,N_3226,N_4681);
or U6715 (N_6715,N_1126,N_3710);
and U6716 (N_6716,N_2357,N_851);
or U6717 (N_6717,N_1878,N_3571);
xor U6718 (N_6718,N_4980,N_1777);
nor U6719 (N_6719,N_912,N_56);
or U6720 (N_6720,N_719,N_1283);
nor U6721 (N_6721,N_282,N_4454);
nand U6722 (N_6722,N_607,N_3882);
or U6723 (N_6723,N_4334,N_2936);
and U6724 (N_6724,N_2681,N_4305);
or U6725 (N_6725,N_4497,N_1121);
nand U6726 (N_6726,N_691,N_2421);
nand U6727 (N_6727,N_508,N_427);
and U6728 (N_6728,N_3254,N_3210);
or U6729 (N_6729,N_1113,N_1181);
nor U6730 (N_6730,N_169,N_1308);
nor U6731 (N_6731,N_4789,N_3012);
nand U6732 (N_6732,N_1118,N_3203);
xnor U6733 (N_6733,N_1780,N_1681);
nor U6734 (N_6734,N_4662,N_876);
nor U6735 (N_6735,N_4461,N_989);
nor U6736 (N_6736,N_2141,N_4027);
and U6737 (N_6737,N_3835,N_1619);
nand U6738 (N_6738,N_1999,N_3674);
nand U6739 (N_6739,N_1189,N_2219);
and U6740 (N_6740,N_2312,N_2250);
or U6741 (N_6741,N_1270,N_610);
nor U6742 (N_6742,N_2491,N_1167);
nor U6743 (N_6743,N_1711,N_1772);
nor U6744 (N_6744,N_2204,N_3573);
and U6745 (N_6745,N_833,N_4493);
or U6746 (N_6746,N_1097,N_3811);
or U6747 (N_6747,N_4216,N_4862);
nor U6748 (N_6748,N_2705,N_3118);
nor U6749 (N_6749,N_4403,N_2362);
nor U6750 (N_6750,N_3057,N_4723);
or U6751 (N_6751,N_2696,N_1617);
nand U6752 (N_6752,N_1183,N_2093);
and U6753 (N_6753,N_667,N_227);
nor U6754 (N_6754,N_2133,N_4758);
nand U6755 (N_6755,N_1108,N_4586);
nor U6756 (N_6756,N_1094,N_831);
and U6757 (N_6757,N_1906,N_1767);
nand U6758 (N_6758,N_2436,N_436);
nand U6759 (N_6759,N_2695,N_413);
or U6760 (N_6760,N_2057,N_3534);
nor U6761 (N_6761,N_1421,N_4954);
nor U6762 (N_6762,N_4348,N_1714);
and U6763 (N_6763,N_4649,N_1260);
nand U6764 (N_6764,N_2927,N_3959);
or U6765 (N_6765,N_4973,N_4164);
and U6766 (N_6766,N_850,N_2444);
nand U6767 (N_6767,N_2971,N_4967);
and U6768 (N_6768,N_1563,N_2982);
nand U6769 (N_6769,N_226,N_1948);
nor U6770 (N_6770,N_4845,N_822);
xnor U6771 (N_6771,N_3600,N_186);
and U6772 (N_6772,N_2353,N_1991);
nand U6773 (N_6773,N_960,N_2566);
and U6774 (N_6774,N_3011,N_288);
and U6775 (N_6775,N_193,N_317);
or U6776 (N_6776,N_1797,N_1589);
and U6777 (N_6777,N_1019,N_3359);
nor U6778 (N_6778,N_1594,N_1540);
or U6779 (N_6779,N_2514,N_1743);
nand U6780 (N_6780,N_2486,N_3097);
and U6781 (N_6781,N_3115,N_419);
xnor U6782 (N_6782,N_503,N_1163);
or U6783 (N_6783,N_4671,N_4072);
nand U6784 (N_6784,N_4449,N_1444);
and U6785 (N_6785,N_3792,N_3391);
nand U6786 (N_6786,N_3469,N_823);
nor U6787 (N_6787,N_2334,N_3716);
nor U6788 (N_6788,N_922,N_3629);
or U6789 (N_6789,N_2531,N_3981);
nand U6790 (N_6790,N_1925,N_2131);
or U6791 (N_6791,N_2364,N_2875);
or U6792 (N_6792,N_533,N_2749);
or U6793 (N_6793,N_1678,N_3542);
and U6794 (N_6794,N_2874,N_4804);
or U6795 (N_6795,N_3134,N_693);
or U6796 (N_6796,N_494,N_864);
nand U6797 (N_6797,N_3292,N_4267);
nand U6798 (N_6798,N_1993,N_3353);
nor U6799 (N_6799,N_2732,N_2934);
nor U6800 (N_6800,N_4934,N_1363);
and U6801 (N_6801,N_4584,N_4032);
nand U6802 (N_6802,N_870,N_1897);
or U6803 (N_6803,N_277,N_1839);
and U6804 (N_6804,N_2355,N_175);
and U6805 (N_6805,N_1611,N_2913);
nor U6806 (N_6806,N_2784,N_2339);
or U6807 (N_6807,N_2074,N_1401);
xor U6808 (N_6808,N_1523,N_1511);
nand U6809 (N_6809,N_2535,N_1888);
nand U6810 (N_6810,N_2268,N_353);
or U6811 (N_6811,N_2686,N_60);
or U6812 (N_6812,N_2891,N_3566);
nand U6813 (N_6813,N_2439,N_3303);
and U6814 (N_6814,N_3992,N_3726);
nand U6815 (N_6815,N_2775,N_453);
or U6816 (N_6816,N_2069,N_2522);
or U6817 (N_6817,N_1463,N_1100);
nand U6818 (N_6818,N_2658,N_1673);
nand U6819 (N_6819,N_2475,N_2072);
nor U6820 (N_6820,N_1583,N_1782);
nor U6821 (N_6821,N_4457,N_2589);
or U6822 (N_6822,N_3432,N_4911);
and U6823 (N_6823,N_3878,N_3263);
nor U6824 (N_6824,N_4791,N_4842);
nand U6825 (N_6825,N_1680,N_1397);
nand U6826 (N_6826,N_2741,N_1491);
nand U6827 (N_6827,N_1733,N_3717);
nor U6828 (N_6828,N_4006,N_4599);
xor U6829 (N_6829,N_2739,N_4965);
nand U6830 (N_6830,N_3124,N_3021);
nand U6831 (N_6831,N_4825,N_4999);
nor U6832 (N_6832,N_2789,N_4376);
xnor U6833 (N_6833,N_2613,N_3840);
nand U6834 (N_6834,N_1983,N_2587);
or U6835 (N_6835,N_3144,N_732);
nand U6836 (N_6836,N_1789,N_3996);
nor U6837 (N_6837,N_1303,N_1739);
or U6838 (N_6838,N_4712,N_2018);
nor U6839 (N_6839,N_3006,N_1435);
or U6840 (N_6840,N_2329,N_410);
or U6841 (N_6841,N_2548,N_569);
or U6842 (N_6842,N_4879,N_3788);
nor U6843 (N_6843,N_2757,N_583);
nor U6844 (N_6844,N_577,N_3285);
nor U6845 (N_6845,N_1685,N_1006);
nor U6846 (N_6846,N_2665,N_2799);
and U6847 (N_6847,N_2823,N_4988);
or U6848 (N_6848,N_3350,N_420);
nand U6849 (N_6849,N_3664,N_3615);
and U6850 (N_6850,N_4076,N_3352);
nor U6851 (N_6851,N_1591,N_936);
nand U6852 (N_6852,N_1724,N_1829);
nand U6853 (N_6853,N_1519,N_3014);
nand U6854 (N_6854,N_2849,N_1735);
xnor U6855 (N_6855,N_4910,N_3019);
and U6856 (N_6856,N_3979,N_2062);
nor U6857 (N_6857,N_161,N_901);
nand U6858 (N_6858,N_2627,N_513);
or U6859 (N_6859,N_2914,N_2774);
nor U6860 (N_6860,N_4964,N_2438);
nand U6861 (N_6861,N_3708,N_2516);
and U6862 (N_6862,N_2217,N_463);
or U6863 (N_6863,N_3640,N_19);
nand U6864 (N_6864,N_4538,N_941);
nand U6865 (N_6865,N_2530,N_619);
and U6866 (N_6866,N_4933,N_1156);
nor U6867 (N_6867,N_4042,N_2071);
and U6868 (N_6868,N_2385,N_2435);
nand U6869 (N_6869,N_1369,N_3342);
nand U6870 (N_6870,N_349,N_4098);
and U6871 (N_6871,N_3587,N_745);
nand U6872 (N_6872,N_663,N_245);
and U6873 (N_6873,N_2918,N_4797);
and U6874 (N_6874,N_4408,N_2006);
or U6875 (N_6875,N_4611,N_3297);
nand U6876 (N_6876,N_1494,N_2121);
nand U6877 (N_6877,N_915,N_2670);
xor U6878 (N_6878,N_2620,N_179);
nor U6879 (N_6879,N_2129,N_3361);
or U6880 (N_6880,N_3093,N_2478);
nor U6881 (N_6881,N_1322,N_3478);
and U6882 (N_6882,N_64,N_344);
nor U6883 (N_6883,N_2107,N_2310);
nand U6884 (N_6884,N_808,N_3179);
nor U6885 (N_6885,N_522,N_509);
nor U6886 (N_6886,N_2386,N_973);
or U6887 (N_6887,N_1420,N_4378);
nand U6888 (N_6888,N_2090,N_2450);
or U6889 (N_6889,N_2785,N_4217);
nor U6890 (N_6890,N_4624,N_159);
or U6891 (N_6891,N_764,N_687);
nand U6892 (N_6892,N_4144,N_1144);
nand U6893 (N_6893,N_2715,N_3829);
nor U6894 (N_6894,N_1890,N_2518);
nand U6895 (N_6895,N_3496,N_1075);
nor U6896 (N_6896,N_4827,N_4389);
nor U6897 (N_6897,N_2326,N_4816);
or U6898 (N_6898,N_1996,N_4021);
or U6899 (N_6899,N_1469,N_1146);
nor U6900 (N_6900,N_3054,N_4291);
nand U6901 (N_6901,N_339,N_438);
or U6902 (N_6902,N_4843,N_514);
nor U6903 (N_6903,N_1980,N_3886);
nor U6904 (N_6904,N_2908,N_806);
or U6905 (N_6905,N_2907,N_4737);
and U6906 (N_6906,N_1952,N_1403);
xnor U6907 (N_6907,N_4821,N_2458);
nand U6908 (N_6908,N_1940,N_547);
nand U6909 (N_6909,N_3802,N_761);
nand U6910 (N_6910,N_4363,N_469);
or U6911 (N_6911,N_1933,N_44);
or U6912 (N_6912,N_4875,N_2572);
nand U6913 (N_6913,N_4229,N_4982);
nor U6914 (N_6914,N_3927,N_4891);
and U6915 (N_6915,N_3764,N_2835);
nand U6916 (N_6916,N_4748,N_4820);
and U6917 (N_6917,N_2500,N_563);
and U6918 (N_6918,N_3244,N_3554);
or U6919 (N_6919,N_1016,N_2233);
and U6920 (N_6920,N_755,N_2646);
nor U6921 (N_6921,N_57,N_705);
and U6922 (N_6922,N_2165,N_2983);
and U6923 (N_6923,N_2306,N_448);
nand U6924 (N_6924,N_908,N_3755);
and U6925 (N_6925,N_627,N_4014);
nor U6926 (N_6926,N_3631,N_2948);
and U6927 (N_6927,N_4283,N_1312);
nor U6928 (N_6928,N_1054,N_2295);
nand U6929 (N_6929,N_3864,N_4214);
and U6930 (N_6930,N_2451,N_4365);
nor U6931 (N_6931,N_3752,N_1442);
or U6932 (N_6932,N_27,N_4446);
or U6933 (N_6933,N_1374,N_1434);
nand U6934 (N_6934,N_4844,N_2443);
nand U6935 (N_6935,N_3395,N_3671);
nor U6936 (N_6936,N_2920,N_1570);
and U6937 (N_6937,N_3698,N_4593);
and U6938 (N_6938,N_2729,N_3920);
and U6939 (N_6939,N_1565,N_2482);
and U6940 (N_6940,N_1968,N_880);
nor U6941 (N_6941,N_3265,N_3096);
xor U6942 (N_6942,N_2009,N_1316);
or U6943 (N_6943,N_1381,N_3856);
nand U6944 (N_6944,N_708,N_3666);
or U6945 (N_6945,N_620,N_1669);
nand U6946 (N_6946,N_4513,N_2027);
or U6947 (N_6947,N_2393,N_3603);
nand U6948 (N_6948,N_818,N_2738);
or U6949 (N_6949,N_3747,N_361);
nor U6950 (N_6950,N_4122,N_1584);
nor U6951 (N_6951,N_2425,N_1031);
or U6952 (N_6952,N_3077,N_3411);
and U6953 (N_6953,N_3512,N_2653);
or U6954 (N_6954,N_4936,N_1893);
nand U6955 (N_6955,N_4632,N_2905);
or U6956 (N_6956,N_2978,N_4103);
nor U6957 (N_6957,N_3908,N_4656);
or U6958 (N_6958,N_916,N_24);
nand U6959 (N_6959,N_2556,N_4336);
nand U6960 (N_6960,N_4786,N_796);
xor U6961 (N_6961,N_2374,N_4046);
nor U6962 (N_6962,N_3586,N_1694);
and U6963 (N_6963,N_1291,N_1241);
xnor U6964 (N_6964,N_2555,N_3466);
xnor U6965 (N_6965,N_3612,N_2058);
and U6966 (N_6966,N_2954,N_3875);
nor U6967 (N_6967,N_253,N_3801);
and U6968 (N_6968,N_3999,N_3880);
and U6969 (N_6969,N_482,N_1493);
nand U6970 (N_6970,N_886,N_2634);
nand U6971 (N_6971,N_1686,N_3955);
or U6972 (N_6972,N_2335,N_2538);
and U6973 (N_6973,N_4795,N_735);
nand U6974 (N_6974,N_3576,N_4134);
nand U6975 (N_6975,N_4510,N_3513);
nand U6976 (N_6976,N_3334,N_2244);
nor U6977 (N_6977,N_4429,N_3585);
or U6978 (N_6978,N_2791,N_2323);
nor U6979 (N_6979,N_1609,N_4633);
and U6980 (N_6980,N_2313,N_4495);
nor U6981 (N_6981,N_1079,N_4019);
or U6982 (N_6982,N_2986,N_3319);
or U6983 (N_6983,N_1687,N_2550);
and U6984 (N_6984,N_2183,N_1210);
or U6985 (N_6985,N_3729,N_1246);
or U6986 (N_6986,N_2136,N_1218);
nor U6987 (N_6987,N_335,N_3360);
or U6988 (N_6988,N_4058,N_336);
or U6989 (N_6989,N_3828,N_4490);
and U6990 (N_6990,N_108,N_3638);
nand U6991 (N_6991,N_4308,N_878);
or U6992 (N_6992,N_2265,N_4766);
nand U6993 (N_6993,N_1652,N_4330);
nand U6994 (N_6994,N_391,N_167);
or U6995 (N_6995,N_2391,N_2091);
nor U6996 (N_6996,N_2236,N_2888);
nor U6997 (N_6997,N_786,N_91);
xnor U6998 (N_6998,N_990,N_1107);
xnor U6999 (N_6999,N_4149,N_1573);
nand U7000 (N_7000,N_3766,N_982);
xnor U7001 (N_7001,N_1659,N_3669);
nor U7002 (N_7002,N_4284,N_4246);
and U7003 (N_7003,N_4280,N_3387);
xor U7004 (N_7004,N_1062,N_2996);
nor U7005 (N_7005,N_2733,N_4868);
or U7006 (N_7006,N_2744,N_231);
nand U7007 (N_7007,N_289,N_747);
and U7008 (N_7008,N_804,N_4398);
and U7009 (N_7009,N_684,N_3313);
xor U7010 (N_7010,N_3195,N_4846);
or U7011 (N_7011,N_2755,N_4993);
nand U7012 (N_7012,N_4678,N_1296);
nand U7013 (N_7013,N_1111,N_4572);
nor U7014 (N_7014,N_2092,N_4300);
nand U7015 (N_7015,N_4832,N_1846);
xor U7016 (N_7016,N_3779,N_4033);
and U7017 (N_7017,N_733,N_3809);
or U7018 (N_7018,N_4276,N_4630);
nor U7019 (N_7019,N_1130,N_334);
or U7020 (N_7020,N_1340,N_308);
and U7021 (N_7021,N_3418,N_470);
nor U7022 (N_7022,N_3605,N_3259);
xnor U7023 (N_7023,N_3949,N_768);
nor U7024 (N_7024,N_4234,N_1185);
or U7025 (N_7025,N_2861,N_1674);
nand U7026 (N_7026,N_2497,N_1248);
nand U7027 (N_7027,N_3156,N_3808);
nand U7028 (N_7028,N_4870,N_524);
nand U7029 (N_7029,N_4400,N_2975);
or U7030 (N_7030,N_3386,N_3385);
and U7031 (N_7031,N_4745,N_893);
nand U7032 (N_7032,N_4282,N_1769);
and U7033 (N_7033,N_783,N_2621);
and U7034 (N_7034,N_1388,N_1792);
nor U7035 (N_7035,N_3786,N_1021);
nor U7036 (N_7036,N_1881,N_3456);
xnor U7037 (N_7037,N_3855,N_1371);
and U7038 (N_7038,N_1345,N_4970);
or U7039 (N_7039,N_1551,N_4128);
nor U7040 (N_7040,N_651,N_4552);
or U7041 (N_7041,N_1648,N_3935);
and U7042 (N_7042,N_3589,N_2713);
nand U7043 (N_7043,N_4703,N_4672);
or U7044 (N_7044,N_4626,N_2469);
or U7045 (N_7045,N_3723,N_394);
or U7046 (N_7046,N_4801,N_3308);
nor U7047 (N_7047,N_1761,N_1037);
nor U7048 (N_7048,N_1939,N_1787);
nand U7049 (N_7049,N_2945,N_4622);
and U7050 (N_7050,N_492,N_1638);
and U7051 (N_7051,N_2606,N_2102);
and U7052 (N_7052,N_4537,N_1275);
nor U7053 (N_7053,N_4623,N_1808);
or U7054 (N_7054,N_70,N_1045);
and U7055 (N_7055,N_2649,N_816);
nor U7056 (N_7056,N_2267,N_3803);
nor U7057 (N_7057,N_2834,N_268);
nor U7058 (N_7058,N_945,N_2297);
or U7059 (N_7059,N_2037,N_3264);
or U7060 (N_7060,N_1227,N_1624);
nor U7061 (N_7061,N_1856,N_1481);
xnor U7062 (N_7062,N_1318,N_3800);
or U7063 (N_7063,N_3438,N_975);
and U7064 (N_7064,N_294,N_4187);
nand U7065 (N_7065,N_3722,N_2227);
or U7066 (N_7066,N_3298,N_4574);
or U7067 (N_7067,N_2382,N_1271);
nor U7068 (N_7068,N_1087,N_314);
or U7069 (N_7069,N_2623,N_4220);
and U7070 (N_7070,N_2229,N_657);
or U7071 (N_7071,N_1359,N_4968);
nand U7072 (N_7072,N_2940,N_1706);
and U7073 (N_7073,N_3026,N_2781);
xor U7074 (N_7074,N_3814,N_2270);
or U7075 (N_7075,N_2722,N_3374);
nand U7076 (N_7076,N_3789,N_4353);
or U7077 (N_7077,N_2151,N_2256);
and U7078 (N_7078,N_4963,N_618);
nor U7079 (N_7079,N_988,N_4718);
or U7080 (N_7080,N_1554,N_4207);
and U7081 (N_7081,N_1593,N_3616);
nor U7082 (N_7082,N_1776,N_3693);
or U7083 (N_7083,N_389,N_715);
nand U7084 (N_7084,N_325,N_1078);
or U7085 (N_7085,N_2626,N_3873);
nand U7086 (N_7086,N_2892,N_2383);
nor U7087 (N_7087,N_400,N_4185);
nor U7088 (N_7088,N_2628,N_443);
and U7089 (N_7089,N_4466,N_1179);
nor U7090 (N_7090,N_3647,N_3175);
and U7091 (N_7091,N_3866,N_63);
nand U7092 (N_7092,N_1122,N_2117);
and U7093 (N_7093,N_4252,N_1423);
and U7094 (N_7094,N_4898,N_3446);
and U7095 (N_7095,N_4332,N_350);
nand U7096 (N_7096,N_3673,N_4271);
nor U7097 (N_7097,N_2184,N_4193);
nor U7098 (N_7098,N_1812,N_2366);
nor U7099 (N_7099,N_754,N_1963);
xor U7100 (N_7100,N_961,N_295);
or U7101 (N_7101,N_1581,N_4053);
and U7102 (N_7102,N_2533,N_4831);
nor U7103 (N_7103,N_2144,N_1247);
or U7104 (N_7104,N_4904,N_4203);
or U7105 (N_7105,N_2937,N_2964);
nand U7106 (N_7106,N_1250,N_4462);
nand U7107 (N_7107,N_4437,N_1093);
or U7108 (N_7108,N_4787,N_3971);
or U7109 (N_7109,N_2534,N_4210);
xnor U7110 (N_7110,N_216,N_271);
nand U7111 (N_7111,N_1147,N_4732);
nor U7112 (N_7112,N_3060,N_3911);
xor U7113 (N_7113,N_1392,N_3168);
or U7114 (N_7114,N_709,N_536);
nand U7115 (N_7115,N_102,N_632);
or U7116 (N_7116,N_4416,N_2953);
or U7117 (N_7117,N_3089,N_3307);
or U7118 (N_7118,N_392,N_4130);
and U7119 (N_7119,N_2167,N_4156);
or U7120 (N_7120,N_842,N_2956);
and U7121 (N_7121,N_4413,N_4107);
or U7122 (N_7122,N_3510,N_2962);
or U7123 (N_7123,N_2094,N_3957);
and U7124 (N_7124,N_1134,N_1645);
nor U7125 (N_7125,N_4169,N_3617);
nor U7126 (N_7126,N_4613,N_4463);
nand U7127 (N_7127,N_1779,N_1509);
nand U7128 (N_7128,N_2782,N_2189);
nand U7129 (N_7129,N_4938,N_4884);
and U7130 (N_7130,N_3176,N_2742);
nor U7131 (N_7131,N_4251,N_387);
nor U7132 (N_7132,N_2719,N_3294);
nand U7133 (N_7133,N_3563,N_1632);
and U7134 (N_7134,N_2762,N_2459);
or U7135 (N_7135,N_435,N_1633);
or U7136 (N_7136,N_3910,N_4556);
xnor U7137 (N_7137,N_2088,N_2041);
nand U7138 (N_7138,N_4882,N_835);
or U7139 (N_7139,N_3987,N_2763);
nor U7140 (N_7140,N_3660,N_2752);
xor U7141 (N_7141,N_313,N_4838);
and U7142 (N_7142,N_2084,N_4040);
and U7143 (N_7143,N_1832,N_384);
or U7144 (N_7144,N_4061,N_2972);
nor U7145 (N_7145,N_3441,N_4991);
xnor U7146 (N_7146,N_493,N_3251);
and U7147 (N_7147,N_2911,N_85);
and U7148 (N_7148,N_3978,N_2568);
nand U7149 (N_7149,N_4519,N_1310);
nor U7150 (N_7150,N_4695,N_3884);
nor U7151 (N_7151,N_866,N_1929);
nand U7152 (N_7152,N_3070,N_1773);
nor U7153 (N_7153,N_2505,N_3613);
nor U7154 (N_7154,N_4101,N_981);
nand U7155 (N_7155,N_3393,N_3842);
nand U7156 (N_7156,N_3727,N_2253);
nand U7157 (N_7157,N_4264,N_4074);
and U7158 (N_7158,N_476,N_149);
nor U7159 (N_7159,N_2724,N_1960);
nand U7160 (N_7160,N_4431,N_3611);
nand U7161 (N_7161,N_4410,N_2557);
xnor U7162 (N_7162,N_1592,N_3562);
nand U7163 (N_7163,N_1176,N_1661);
nor U7164 (N_7164,N_2381,N_1682);
and U7165 (N_7165,N_2426,N_2317);
nand U7166 (N_7166,N_2493,N_3934);
xnor U7167 (N_7167,N_3002,N_1944);
xor U7168 (N_7168,N_937,N_1115);
nand U7169 (N_7169,N_81,N_3940);
and U7170 (N_7170,N_214,N_255);
nor U7171 (N_7171,N_515,N_3997);
nor U7172 (N_7172,N_1399,N_1601);
and U7173 (N_7173,N_2429,N_3588);
nor U7174 (N_7174,N_187,N_2622);
xnor U7175 (N_7175,N_3550,N_1998);
and U7176 (N_7176,N_1066,N_338);
nor U7177 (N_7177,N_442,N_2012);
nand U7178 (N_7178,N_4157,N_1058);
or U7179 (N_7179,N_1287,N_718);
nor U7180 (N_7180,N_539,N_1415);
xor U7181 (N_7181,N_103,N_2328);
xnor U7182 (N_7182,N_1450,N_1194);
nor U7183 (N_7183,N_1382,N_4969);
nand U7184 (N_7184,N_4399,N_4097);
xnor U7185 (N_7185,N_2225,N_322);
and U7186 (N_7186,N_3876,N_2974);
or U7187 (N_7187,N_53,N_3328);
and U7188 (N_7188,N_136,N_286);
or U7189 (N_7189,N_3202,N_572);
nand U7190 (N_7190,N_2410,N_441);
and U7191 (N_7191,N_2515,N_4515);
nor U7192 (N_7192,N_3367,N_3228);
or U7193 (N_7193,N_1222,N_3703);
nand U7194 (N_7194,N_42,N_4529);
or U7195 (N_7195,N_2652,N_4456);
or U7196 (N_7196,N_1802,N_51);
or U7197 (N_7197,N_1616,N_4690);
and U7198 (N_7198,N_4339,N_4929);
nor U7199 (N_7199,N_240,N_1207);
and U7200 (N_7200,N_464,N_888);
nand U7201 (N_7201,N_1478,N_3844);
or U7202 (N_7202,N_2457,N_2148);
or U7203 (N_7203,N_2476,N_1649);
and U7204 (N_7204,N_566,N_1069);
or U7205 (N_7205,N_303,N_1668);
nor U7206 (N_7206,N_562,N_4930);
or U7207 (N_7207,N_3776,N_3604);
or U7208 (N_7208,N_4356,N_775);
or U7209 (N_7209,N_4369,N_3200);
nor U7210 (N_7210,N_653,N_4733);
nor U7211 (N_7211,N_395,N_2271);
nor U7212 (N_7212,N_595,N_1288);
nand U7213 (N_7213,N_2318,N_3122);
nand U7214 (N_7214,N_2801,N_4423);
or U7215 (N_7215,N_911,N_2599);
nand U7216 (N_7216,N_4323,N_4643);
nand U7217 (N_7217,N_2489,N_2767);
nor U7218 (N_7218,N_2239,N_883);
nor U7219 (N_7219,N_1857,N_215);
nor U7220 (N_7220,N_897,N_2452);
and U7221 (N_7221,N_3599,N_1618);
or U7222 (N_7222,N_1578,N_3373);
and U7223 (N_7223,N_4822,N_2025);
xnor U7224 (N_7224,N_3044,N_3052);
nor U7225 (N_7225,N_2734,N_4057);
and U7226 (N_7226,N_2873,N_287);
and U7227 (N_7227,N_3699,N_2054);
or U7228 (N_7228,N_4124,N_1755);
nand U7229 (N_7229,N_4614,N_4577);
nand U7230 (N_7230,N_1261,N_1865);
nor U7231 (N_7231,N_3455,N_1742);
nand U7232 (N_7232,N_2553,N_3862);
nor U7233 (N_7233,N_807,N_4075);
nand U7234 (N_7234,N_4533,N_123);
or U7235 (N_7235,N_1811,N_4641);
and U7236 (N_7236,N_4020,N_131);
nor U7237 (N_7237,N_4406,N_2440);
and U7238 (N_7238,N_4049,N_1783);
or U7239 (N_7239,N_1038,N_3409);
nand U7240 (N_7240,N_4660,N_4478);
nor U7241 (N_7241,N_2220,N_4161);
and U7242 (N_7242,N_997,N_1701);
and U7243 (N_7243,N_1824,N_3930);
nand U7244 (N_7244,N_1484,N_4591);
and U7245 (N_7245,N_892,N_3552);
nor U7246 (N_7246,N_4176,N_2853);
or U7247 (N_7247,N_4892,N_3728);
and U7248 (N_7248,N_481,N_4442);
nor U7249 (N_7249,N_2418,N_953);
or U7250 (N_7250,N_3320,N_4063);
nand U7251 (N_7251,N_4603,N_4923);
nand U7252 (N_7252,N_2610,N_388);
xnor U7253 (N_7253,N_95,N_3639);
or U7254 (N_7254,N_3575,N_2735);
nor U7255 (N_7255,N_2800,N_3082);
and U7256 (N_7256,N_2423,N_2162);
nor U7257 (N_7257,N_1035,N_669);
nand U7258 (N_7258,N_643,N_1657);
and U7259 (N_7259,N_4648,N_4562);
nor U7260 (N_7260,N_3484,N_1129);
xor U7261 (N_7261,N_1915,N_3929);
xor U7262 (N_7262,N_4116,N_3047);
nand U7263 (N_7263,N_1508,N_4003);
nand U7264 (N_7264,N_4859,N_3591);
nor U7265 (N_7265,N_1257,N_3165);
xnor U7266 (N_7266,N_4153,N_4137);
nor U7267 (N_7267,N_1154,N_3045);
nor U7268 (N_7268,N_1490,N_1328);
nand U7269 (N_7269,N_4022,N_4900);
or U7270 (N_7270,N_88,N_889);
and U7271 (N_7271,N_37,N_661);
and U7272 (N_7272,N_2595,N_1479);
or U7273 (N_7273,N_1251,N_4727);
and U7274 (N_7274,N_3902,N_1465);
or U7275 (N_7275,N_21,N_3414);
or U7276 (N_7276,N_3269,N_2276);
or U7277 (N_7277,N_2448,N_3001);
and U7278 (N_7278,N_3224,N_2047);
or U7279 (N_7279,N_3841,N_4535);
and U7280 (N_7280,N_2523,N_109);
and U7281 (N_7281,N_4619,N_1969);
nor U7282 (N_7282,N_4133,N_3595);
nor U7283 (N_7283,N_1139,N_1781);
nor U7284 (N_7284,N_2816,N_2917);
and U7285 (N_7285,N_28,N_4102);
and U7286 (N_7286,N_3197,N_4327);
nor U7287 (N_7287,N_2794,N_3487);
nor U7288 (N_7288,N_2327,N_423);
and U7289 (N_7289,N_710,N_1548);
nor U7290 (N_7290,N_1412,N_4652);
nor U7291 (N_7291,N_316,N_4066);
nand U7292 (N_7292,N_4636,N_3273);
or U7293 (N_7293,N_1057,N_3318);
nor U7294 (N_7294,N_265,N_4823);
and U7295 (N_7295,N_834,N_3349);
or U7296 (N_7296,N_4686,N_2202);
or U7297 (N_7297,N_2248,N_1089);
and U7298 (N_7298,N_1603,N_1455);
nand U7299 (N_7299,N_3399,N_2437);
nand U7300 (N_7300,N_3062,N_2858);
nand U7301 (N_7301,N_2825,N_2333);
xor U7302 (N_7302,N_2902,N_1117);
and U7303 (N_7303,N_2417,N_2612);
and U7304 (N_7304,N_3452,N_1804);
nand U7305 (N_7305,N_2901,N_2419);
nand U7306 (N_7306,N_4208,N_3234);
nand U7307 (N_7307,N_3816,N_1332);
and U7308 (N_7308,N_1796,N_3633);
nor U7309 (N_7309,N_977,N_523);
nor U7310 (N_7310,N_4736,N_2361);
nand U7311 (N_7311,N_1614,N_132);
and U7312 (N_7312,N_4221,N_3621);
nand U7313 (N_7313,N_3662,N_3120);
or U7314 (N_7314,N_258,N_3746);
xnor U7315 (N_7315,N_4105,N_4990);
and U7316 (N_7316,N_1076,N_856);
or U7317 (N_7317,N_4412,N_2668);
nand U7318 (N_7318,N_71,N_3031);
and U7319 (N_7319,N_4263,N_4985);
nor U7320 (N_7320,N_858,N_358);
and U7321 (N_7321,N_694,N_2863);
and U7322 (N_7322,N_3740,N_2960);
and U7323 (N_7323,N_208,N_348);
or U7324 (N_7324,N_2837,N_2492);
nand U7325 (N_7325,N_3300,N_218);
xor U7326 (N_7326,N_2147,N_2679);
and U7327 (N_7327,N_2216,N_1358);
or U7328 (N_7328,N_3447,N_299);
nor U7329 (N_7329,N_3869,N_1825);
xnor U7330 (N_7330,N_2759,N_210);
and U7331 (N_7331,N_869,N_575);
nand U7332 (N_7332,N_3773,N_4126);
xnor U7333 (N_7333,N_1507,N_1086);
and U7334 (N_7334,N_4542,N_3646);
or U7335 (N_7335,N_342,N_2780);
and U7336 (N_7336,N_631,N_4065);
nand U7337 (N_7337,N_1958,N_1212);
xor U7338 (N_7338,N_798,N_4004);
nand U7339 (N_7339,N_1665,N_3394);
and U7340 (N_7340,N_1109,N_4159);
or U7341 (N_7341,N_3879,N_2106);
or U7342 (N_7342,N_1964,N_1356);
and U7343 (N_7343,N_1788,N_4338);
or U7344 (N_7344,N_398,N_4419);
or U7345 (N_7345,N_2826,N_1378);
nand U7346 (N_7346,N_4052,N_3003);
and U7347 (N_7347,N_105,N_3581);
nand U7348 (N_7348,N_1240,N_2496);
or U7349 (N_7349,N_2680,N_4639);
nand U7350 (N_7350,N_4240,N_3073);
nand U7351 (N_7351,N_2389,N_817);
or U7352 (N_7352,N_201,N_2240);
nor U7353 (N_7353,N_1622,N_4071);
nor U7354 (N_7354,N_4425,N_3557);
and U7355 (N_7355,N_3225,N_3085);
or U7356 (N_7356,N_333,N_3147);
nand U7357 (N_7357,N_4860,N_2771);
nor U7358 (N_7358,N_1336,N_87);
or U7359 (N_7359,N_2810,N_4755);
nand U7360 (N_7360,N_2688,N_943);
nor U7361 (N_7361,N_329,N_3413);
and U7362 (N_7362,N_439,N_4035);
nand U7363 (N_7363,N_1027,N_4762);
nor U7364 (N_7364,N_2632,N_3714);
or U7365 (N_7365,N_2597,N_190);
nor U7366 (N_7366,N_1709,N_3794);
or U7367 (N_7367,N_1440,N_1095);
nor U7368 (N_7368,N_1425,N_819);
or U7369 (N_7369,N_4081,N_2809);
or U7370 (N_7370,N_2281,N_297);
or U7371 (N_7371,N_1924,N_3064);
nand U7372 (N_7372,N_1152,N_1966);
nor U7373 (N_7373,N_2209,N_2831);
and U7374 (N_7374,N_4581,N_2541);
and U7375 (N_7375,N_2203,N_845);
and U7376 (N_7376,N_4131,N_2086);
nand U7377 (N_7377,N_2788,N_3161);
or U7378 (N_7378,N_629,N_1470);
and U7379 (N_7379,N_830,N_1778);
and U7380 (N_7380,N_4793,N_3192);
xnor U7381 (N_7381,N_730,N_3299);
and U7382 (N_7382,N_3966,N_4444);
or U7383 (N_7383,N_4481,N_1158);
or U7384 (N_7384,N_4854,N_2859);
nand U7385 (N_7385,N_1521,N_3804);
nor U7386 (N_7386,N_4079,N_2038);
xnor U7387 (N_7387,N_4725,N_3271);
and U7388 (N_7388,N_173,N_1961);
and U7389 (N_7389,N_4948,N_475);
and U7390 (N_7390,N_3988,N_2841);
nand U7391 (N_7391,N_4085,N_2394);
or U7392 (N_7392,N_2139,N_4540);
or U7393 (N_7393,N_1279,N_564);
xnor U7394 (N_7394,N_3899,N_4667);
nor U7395 (N_7395,N_1828,N_647);
or U7396 (N_7396,N_2614,N_4939);
nor U7397 (N_7397,N_3777,N_498);
and U7398 (N_7398,N_4864,N_771);
or U7399 (N_7399,N_4448,N_3178);
xor U7400 (N_7400,N_3540,N_1239);
nor U7401 (N_7401,N_1526,N_1417);
nand U7402 (N_7402,N_3847,N_2016);
nand U7403 (N_7403,N_1234,N_4877);
nand U7404 (N_7404,N_2987,N_788);
and U7405 (N_7405,N_1447,N_2257);
or U7406 (N_7406,N_1911,N_751);
or U7407 (N_7407,N_140,N_3435);
nor U7408 (N_7408,N_2157,N_1842);
xor U7409 (N_7409,N_1339,N_601);
or U7410 (N_7410,N_3157,N_885);
or U7411 (N_7411,N_1418,N_1898);
nor U7412 (N_7412,N_1174,N_3720);
nor U7413 (N_7413,N_196,N_1654);
and U7414 (N_7414,N_1934,N_1984);
nand U7415 (N_7415,N_4979,N_4231);
nor U7416 (N_7416,N_1326,N_445);
nor U7417 (N_7417,N_3131,N_3036);
or U7418 (N_7418,N_2564,N_2537);
xnor U7419 (N_7419,N_3428,N_3559);
or U7420 (N_7420,N_4404,N_3442);
nor U7421 (N_7421,N_4009,N_315);
nor U7422 (N_7422,N_3315,N_2743);
and U7423 (N_7423,N_1024,N_1145);
nor U7424 (N_7424,N_3295,N_4479);
nor U7425 (N_7425,N_3974,N_84);
or U7426 (N_7426,N_3682,N_1597);
nor U7427 (N_7427,N_4093,N_4307);
and U7428 (N_7428,N_2924,N_4023);
and U7429 (N_7429,N_639,N_1405);
and U7430 (N_7430,N_1344,N_2641);
or U7431 (N_7431,N_2786,N_238);
nand U7432 (N_7432,N_3154,N_4589);
nand U7433 (N_7433,N_4761,N_2369);
and U7434 (N_7434,N_4387,N_3310);
nor U7435 (N_7435,N_3672,N_4638);
and U7436 (N_7436,N_248,N_3356);
xnor U7437 (N_7437,N_2017,N_3885);
nor U7438 (N_7438,N_1650,N_1159);
nand U7439 (N_7439,N_3218,N_743);
or U7440 (N_7440,N_3417,N_1555);
nand U7441 (N_7441,N_1547,N_756);
and U7442 (N_7442,N_2952,N_2332);
or U7443 (N_7443,N_3220,N_789);
nor U7444 (N_7444,N_2365,N_4025);
and U7445 (N_7445,N_3820,N_3110);
nand U7446 (N_7446,N_898,N_2373);
nand U7447 (N_7447,N_1987,N_2596);
or U7448 (N_7448,N_4024,N_1039);
or U7449 (N_7449,N_2736,N_2195);
nand U7450 (N_7450,N_1590,N_148);
and U7451 (N_7451,N_546,N_3103);
and U7452 (N_7452,N_2852,N_2414);
and U7453 (N_7453,N_2527,N_2989);
nor U7454 (N_7454,N_4935,N_2647);
nand U7455 (N_7455,N_4492,N_340);
and U7456 (N_7456,N_2000,N_1014);
and U7457 (N_7457,N_2095,N_701);
and U7458 (N_7458,N_2488,N_3903);
nor U7459 (N_7459,N_3818,N_1389);
and U7460 (N_7460,N_1585,N_3221);
nand U7461 (N_7461,N_984,N_1720);
xor U7462 (N_7462,N_147,N_2024);
and U7463 (N_7463,N_7,N_3151);
or U7464 (N_7464,N_4224,N_4676);
nor U7465 (N_7465,N_606,N_2919);
nor U7466 (N_7466,N_2669,N_4368);
nand U7467 (N_7467,N_3543,N_794);
or U7468 (N_7468,N_323,N_676);
xor U7469 (N_7469,N_3473,N_2519);
nand U7470 (N_7470,N_1051,N_3102);
nand U7471 (N_7471,N_486,N_2929);
and U7472 (N_7472,N_965,N_2346);
or U7473 (N_7473,N_4960,N_1354);
or U7474 (N_7474,N_815,N_4374);
nand U7475 (N_7475,N_415,N_4545);
nand U7476 (N_7476,N_4477,N_4940);
nand U7477 (N_7477,N_2648,N_993);
nand U7478 (N_7478,N_2546,N_3508);
or U7479 (N_7479,N_2707,N_2625);
nand U7480 (N_7480,N_4771,N_3965);
xnor U7481 (N_7481,N_3692,N_4602);
and U7482 (N_7482,N_1365,N_1725);
or U7483 (N_7483,N_4459,N_2031);
nand U7484 (N_7484,N_1196,N_4335);
and U7485 (N_7485,N_4039,N_1462);
nor U7486 (N_7486,N_4120,N_4597);
nand U7487 (N_7487,N_2097,N_802);
nor U7488 (N_7488,N_460,N_1537);
nor U7489 (N_7489,N_2727,N_1173);
or U7490 (N_7490,N_3630,N_1544);
or U7491 (N_7491,N_4018,N_3778);
nand U7492 (N_7492,N_72,N_2308);
and U7493 (N_7493,N_2509,N_3578);
xor U7494 (N_7494,N_236,N_1448);
or U7495 (N_7495,N_4129,N_2525);
and U7496 (N_7496,N_4197,N_1512);
nand U7497 (N_7497,N_2099,N_1072);
xor U7498 (N_7498,N_1242,N_454);
nand U7499 (N_7499,N_1689,N_598);
nand U7500 (N_7500,N_4954,N_508);
and U7501 (N_7501,N_4673,N_4211);
nand U7502 (N_7502,N_3527,N_65);
and U7503 (N_7503,N_4603,N_3730);
or U7504 (N_7504,N_516,N_1771);
nand U7505 (N_7505,N_47,N_2379);
or U7506 (N_7506,N_1185,N_2078);
xnor U7507 (N_7507,N_1547,N_496);
nand U7508 (N_7508,N_4252,N_71);
and U7509 (N_7509,N_2484,N_2660);
or U7510 (N_7510,N_176,N_4302);
nor U7511 (N_7511,N_1297,N_3364);
nor U7512 (N_7512,N_4450,N_2442);
nor U7513 (N_7513,N_1461,N_2033);
and U7514 (N_7514,N_1400,N_4863);
nor U7515 (N_7515,N_498,N_1212);
nor U7516 (N_7516,N_2592,N_2185);
or U7517 (N_7517,N_2348,N_3565);
nand U7518 (N_7518,N_2225,N_1585);
or U7519 (N_7519,N_1772,N_1501);
or U7520 (N_7520,N_3982,N_2781);
nor U7521 (N_7521,N_1492,N_1493);
nor U7522 (N_7522,N_60,N_168);
nor U7523 (N_7523,N_127,N_1293);
or U7524 (N_7524,N_4741,N_4406);
or U7525 (N_7525,N_3579,N_1530);
nor U7526 (N_7526,N_1358,N_2200);
and U7527 (N_7527,N_4256,N_1636);
and U7528 (N_7528,N_4218,N_1888);
xnor U7529 (N_7529,N_1771,N_2658);
nand U7530 (N_7530,N_4615,N_357);
and U7531 (N_7531,N_4894,N_4328);
nand U7532 (N_7532,N_221,N_2571);
or U7533 (N_7533,N_4060,N_3235);
nor U7534 (N_7534,N_1923,N_4732);
or U7535 (N_7535,N_4725,N_65);
or U7536 (N_7536,N_2458,N_4219);
xnor U7537 (N_7537,N_491,N_3434);
and U7538 (N_7538,N_2615,N_1043);
xnor U7539 (N_7539,N_4078,N_1799);
or U7540 (N_7540,N_799,N_1164);
or U7541 (N_7541,N_530,N_3966);
nand U7542 (N_7542,N_2118,N_4748);
or U7543 (N_7543,N_433,N_2598);
nor U7544 (N_7544,N_1428,N_417);
or U7545 (N_7545,N_1293,N_2130);
and U7546 (N_7546,N_1756,N_2508);
nor U7547 (N_7547,N_1226,N_1956);
nor U7548 (N_7548,N_2259,N_2820);
and U7549 (N_7549,N_1601,N_3781);
or U7550 (N_7550,N_1434,N_3135);
or U7551 (N_7551,N_3730,N_4634);
nor U7552 (N_7552,N_2652,N_1652);
or U7553 (N_7553,N_447,N_1434);
and U7554 (N_7554,N_436,N_4541);
nand U7555 (N_7555,N_1264,N_3400);
nor U7556 (N_7556,N_4331,N_1369);
xnor U7557 (N_7557,N_4888,N_4966);
nor U7558 (N_7558,N_4436,N_2273);
nor U7559 (N_7559,N_4655,N_854);
nor U7560 (N_7560,N_3933,N_629);
and U7561 (N_7561,N_1820,N_2242);
xnor U7562 (N_7562,N_1051,N_4494);
xnor U7563 (N_7563,N_3127,N_2966);
nor U7564 (N_7564,N_3210,N_97);
nand U7565 (N_7565,N_1909,N_702);
or U7566 (N_7566,N_1701,N_3071);
and U7567 (N_7567,N_1747,N_1007);
nand U7568 (N_7568,N_2684,N_1315);
nand U7569 (N_7569,N_3948,N_361);
nor U7570 (N_7570,N_3771,N_2938);
or U7571 (N_7571,N_4458,N_3616);
xor U7572 (N_7572,N_2692,N_1463);
nor U7573 (N_7573,N_1848,N_2827);
nor U7574 (N_7574,N_240,N_4635);
nand U7575 (N_7575,N_85,N_2016);
nand U7576 (N_7576,N_1805,N_3604);
nand U7577 (N_7577,N_2541,N_4151);
nand U7578 (N_7578,N_237,N_2192);
nand U7579 (N_7579,N_575,N_430);
or U7580 (N_7580,N_3470,N_1465);
nand U7581 (N_7581,N_4239,N_2176);
and U7582 (N_7582,N_4275,N_4458);
nor U7583 (N_7583,N_2909,N_3369);
nor U7584 (N_7584,N_1682,N_4544);
or U7585 (N_7585,N_1394,N_194);
nand U7586 (N_7586,N_1140,N_982);
and U7587 (N_7587,N_4240,N_4200);
nor U7588 (N_7588,N_2314,N_437);
nor U7589 (N_7589,N_1767,N_2450);
or U7590 (N_7590,N_4647,N_4839);
nand U7591 (N_7591,N_3155,N_4951);
nand U7592 (N_7592,N_402,N_4038);
xnor U7593 (N_7593,N_4442,N_592);
and U7594 (N_7594,N_3689,N_2179);
nor U7595 (N_7595,N_4992,N_616);
xor U7596 (N_7596,N_1046,N_4006);
and U7597 (N_7597,N_3667,N_1670);
and U7598 (N_7598,N_1757,N_1914);
and U7599 (N_7599,N_3296,N_2915);
nor U7600 (N_7600,N_2803,N_3710);
or U7601 (N_7601,N_1928,N_4277);
and U7602 (N_7602,N_3863,N_414);
or U7603 (N_7603,N_4098,N_3525);
or U7604 (N_7604,N_4063,N_1743);
nor U7605 (N_7605,N_2889,N_4236);
or U7606 (N_7606,N_4474,N_2226);
nor U7607 (N_7607,N_3628,N_2085);
and U7608 (N_7608,N_3092,N_4116);
nand U7609 (N_7609,N_1281,N_2682);
nand U7610 (N_7610,N_3617,N_4744);
nand U7611 (N_7611,N_3826,N_1235);
nor U7612 (N_7612,N_1791,N_3853);
and U7613 (N_7613,N_846,N_1685);
or U7614 (N_7614,N_4997,N_2873);
nand U7615 (N_7615,N_536,N_3222);
nor U7616 (N_7616,N_1891,N_2842);
xor U7617 (N_7617,N_2095,N_4022);
nor U7618 (N_7618,N_3303,N_235);
nand U7619 (N_7619,N_4766,N_4187);
or U7620 (N_7620,N_1731,N_1356);
nor U7621 (N_7621,N_739,N_4206);
and U7622 (N_7622,N_900,N_65);
xnor U7623 (N_7623,N_2261,N_60);
nand U7624 (N_7624,N_4689,N_1194);
and U7625 (N_7625,N_378,N_4207);
nand U7626 (N_7626,N_4621,N_4717);
nand U7627 (N_7627,N_847,N_1544);
and U7628 (N_7628,N_1383,N_870);
or U7629 (N_7629,N_285,N_342);
xor U7630 (N_7630,N_684,N_322);
nand U7631 (N_7631,N_1690,N_900);
or U7632 (N_7632,N_3363,N_1084);
nor U7633 (N_7633,N_4962,N_3517);
or U7634 (N_7634,N_4972,N_2123);
or U7635 (N_7635,N_2345,N_884);
nand U7636 (N_7636,N_3851,N_990);
or U7637 (N_7637,N_2359,N_4239);
nor U7638 (N_7638,N_1176,N_3705);
nor U7639 (N_7639,N_3283,N_3622);
or U7640 (N_7640,N_4507,N_4425);
nor U7641 (N_7641,N_3339,N_3008);
and U7642 (N_7642,N_1789,N_2473);
nand U7643 (N_7643,N_2842,N_220);
nand U7644 (N_7644,N_1709,N_1582);
and U7645 (N_7645,N_2207,N_1402);
or U7646 (N_7646,N_4751,N_2782);
or U7647 (N_7647,N_3546,N_1675);
nor U7648 (N_7648,N_2007,N_1901);
nor U7649 (N_7649,N_889,N_3413);
nand U7650 (N_7650,N_4680,N_996);
nand U7651 (N_7651,N_4528,N_2760);
nand U7652 (N_7652,N_2631,N_4102);
or U7653 (N_7653,N_2498,N_730);
and U7654 (N_7654,N_4094,N_2468);
nand U7655 (N_7655,N_1499,N_1234);
nor U7656 (N_7656,N_3591,N_2094);
nand U7657 (N_7657,N_882,N_1597);
and U7658 (N_7658,N_251,N_2706);
or U7659 (N_7659,N_2953,N_2993);
nor U7660 (N_7660,N_943,N_4026);
nor U7661 (N_7661,N_3958,N_2843);
and U7662 (N_7662,N_2285,N_3568);
or U7663 (N_7663,N_3314,N_4511);
xor U7664 (N_7664,N_1239,N_2751);
or U7665 (N_7665,N_2524,N_3627);
nand U7666 (N_7666,N_2220,N_342);
and U7667 (N_7667,N_2944,N_1586);
or U7668 (N_7668,N_3371,N_1055);
nand U7669 (N_7669,N_2675,N_4690);
and U7670 (N_7670,N_2436,N_4243);
nand U7671 (N_7671,N_1156,N_518);
and U7672 (N_7672,N_2950,N_1447);
nand U7673 (N_7673,N_3181,N_2559);
nor U7674 (N_7674,N_367,N_4188);
nor U7675 (N_7675,N_4191,N_4013);
and U7676 (N_7676,N_271,N_2908);
nand U7677 (N_7677,N_1764,N_4007);
nor U7678 (N_7678,N_540,N_1002);
nor U7679 (N_7679,N_2503,N_3993);
nor U7680 (N_7680,N_531,N_3220);
and U7681 (N_7681,N_1957,N_2249);
xnor U7682 (N_7682,N_1408,N_3857);
nor U7683 (N_7683,N_2437,N_4139);
or U7684 (N_7684,N_2160,N_535);
nand U7685 (N_7685,N_3583,N_4404);
nor U7686 (N_7686,N_2435,N_2701);
nand U7687 (N_7687,N_367,N_4388);
xor U7688 (N_7688,N_2041,N_3373);
and U7689 (N_7689,N_2132,N_2612);
xnor U7690 (N_7690,N_4105,N_210);
and U7691 (N_7691,N_4624,N_4728);
or U7692 (N_7692,N_2836,N_4279);
and U7693 (N_7693,N_4958,N_251);
nand U7694 (N_7694,N_4081,N_271);
nor U7695 (N_7695,N_4074,N_4787);
nand U7696 (N_7696,N_4972,N_2994);
nor U7697 (N_7697,N_408,N_3432);
and U7698 (N_7698,N_1074,N_4280);
nor U7699 (N_7699,N_3540,N_4262);
and U7700 (N_7700,N_3028,N_4104);
nor U7701 (N_7701,N_1111,N_1768);
nand U7702 (N_7702,N_3340,N_1291);
nand U7703 (N_7703,N_4241,N_4273);
xor U7704 (N_7704,N_68,N_4244);
or U7705 (N_7705,N_1583,N_2730);
nand U7706 (N_7706,N_2950,N_306);
nor U7707 (N_7707,N_4036,N_1962);
and U7708 (N_7708,N_3392,N_3562);
and U7709 (N_7709,N_1070,N_3830);
nand U7710 (N_7710,N_3447,N_889);
nor U7711 (N_7711,N_365,N_4207);
or U7712 (N_7712,N_3664,N_4999);
nand U7713 (N_7713,N_1745,N_2213);
and U7714 (N_7714,N_2246,N_27);
and U7715 (N_7715,N_1526,N_1541);
nor U7716 (N_7716,N_867,N_1937);
or U7717 (N_7717,N_4179,N_3307);
nor U7718 (N_7718,N_458,N_4249);
or U7719 (N_7719,N_2315,N_1902);
or U7720 (N_7720,N_1166,N_2500);
nand U7721 (N_7721,N_4462,N_272);
or U7722 (N_7722,N_1519,N_2696);
or U7723 (N_7723,N_2328,N_4767);
nor U7724 (N_7724,N_4840,N_2861);
nor U7725 (N_7725,N_3522,N_2541);
and U7726 (N_7726,N_3018,N_4953);
or U7727 (N_7727,N_1310,N_851);
or U7728 (N_7728,N_2891,N_1319);
and U7729 (N_7729,N_366,N_4347);
or U7730 (N_7730,N_1366,N_3476);
nor U7731 (N_7731,N_4208,N_2945);
and U7732 (N_7732,N_3250,N_4169);
nand U7733 (N_7733,N_229,N_428);
or U7734 (N_7734,N_3007,N_4094);
nor U7735 (N_7735,N_4253,N_4432);
nor U7736 (N_7736,N_1376,N_4340);
nand U7737 (N_7737,N_58,N_696);
nor U7738 (N_7738,N_1861,N_2847);
nor U7739 (N_7739,N_4834,N_1209);
or U7740 (N_7740,N_748,N_3360);
nor U7741 (N_7741,N_4756,N_1983);
or U7742 (N_7742,N_2836,N_2329);
xnor U7743 (N_7743,N_3352,N_471);
and U7744 (N_7744,N_464,N_4773);
and U7745 (N_7745,N_4946,N_2496);
and U7746 (N_7746,N_4428,N_2663);
nand U7747 (N_7747,N_563,N_3816);
or U7748 (N_7748,N_2400,N_896);
or U7749 (N_7749,N_4321,N_286);
nor U7750 (N_7750,N_1634,N_1798);
nor U7751 (N_7751,N_3969,N_3463);
and U7752 (N_7752,N_3196,N_2156);
or U7753 (N_7753,N_3513,N_4856);
nor U7754 (N_7754,N_1154,N_4150);
nand U7755 (N_7755,N_1532,N_3312);
or U7756 (N_7756,N_1478,N_1741);
and U7757 (N_7757,N_2866,N_4931);
xor U7758 (N_7758,N_4607,N_2444);
and U7759 (N_7759,N_276,N_2761);
nor U7760 (N_7760,N_783,N_4311);
and U7761 (N_7761,N_4658,N_3309);
nor U7762 (N_7762,N_1454,N_4643);
or U7763 (N_7763,N_1558,N_3211);
or U7764 (N_7764,N_2194,N_1197);
or U7765 (N_7765,N_4309,N_3583);
xor U7766 (N_7766,N_3432,N_3466);
and U7767 (N_7767,N_1379,N_4920);
or U7768 (N_7768,N_2484,N_3815);
nor U7769 (N_7769,N_793,N_1409);
or U7770 (N_7770,N_2091,N_2650);
and U7771 (N_7771,N_1470,N_4433);
and U7772 (N_7772,N_4842,N_2715);
nand U7773 (N_7773,N_4953,N_2705);
xnor U7774 (N_7774,N_4053,N_2914);
or U7775 (N_7775,N_1558,N_2716);
or U7776 (N_7776,N_1829,N_4320);
and U7777 (N_7777,N_1898,N_3438);
nor U7778 (N_7778,N_2993,N_4134);
xor U7779 (N_7779,N_1921,N_3283);
and U7780 (N_7780,N_3250,N_2215);
and U7781 (N_7781,N_1082,N_3358);
xnor U7782 (N_7782,N_1975,N_3487);
xnor U7783 (N_7783,N_4496,N_236);
nand U7784 (N_7784,N_748,N_4036);
and U7785 (N_7785,N_1972,N_268);
and U7786 (N_7786,N_1812,N_1547);
xnor U7787 (N_7787,N_129,N_646);
nor U7788 (N_7788,N_2803,N_2126);
nand U7789 (N_7789,N_1706,N_4253);
and U7790 (N_7790,N_30,N_2347);
or U7791 (N_7791,N_3217,N_3976);
xnor U7792 (N_7792,N_2442,N_4621);
or U7793 (N_7793,N_1251,N_3261);
and U7794 (N_7794,N_1797,N_4083);
or U7795 (N_7795,N_228,N_3208);
xor U7796 (N_7796,N_4186,N_244);
nor U7797 (N_7797,N_2380,N_4201);
nand U7798 (N_7798,N_22,N_4312);
nand U7799 (N_7799,N_1418,N_3454);
nor U7800 (N_7800,N_2220,N_3796);
xnor U7801 (N_7801,N_4957,N_4216);
xor U7802 (N_7802,N_4599,N_563);
and U7803 (N_7803,N_4676,N_3426);
xor U7804 (N_7804,N_2222,N_1702);
and U7805 (N_7805,N_4621,N_559);
nand U7806 (N_7806,N_2928,N_3638);
nor U7807 (N_7807,N_656,N_2947);
or U7808 (N_7808,N_2284,N_2804);
nand U7809 (N_7809,N_209,N_9);
nand U7810 (N_7810,N_2422,N_3171);
nand U7811 (N_7811,N_3423,N_1223);
or U7812 (N_7812,N_1853,N_4482);
or U7813 (N_7813,N_504,N_1133);
and U7814 (N_7814,N_3717,N_361);
nor U7815 (N_7815,N_1079,N_128);
nor U7816 (N_7816,N_3820,N_3807);
nand U7817 (N_7817,N_2622,N_1974);
nor U7818 (N_7818,N_3775,N_1504);
or U7819 (N_7819,N_1064,N_3682);
nand U7820 (N_7820,N_3680,N_4667);
nor U7821 (N_7821,N_1689,N_4124);
and U7822 (N_7822,N_1183,N_333);
and U7823 (N_7823,N_1470,N_1260);
nor U7824 (N_7824,N_1631,N_2676);
and U7825 (N_7825,N_2087,N_4753);
and U7826 (N_7826,N_4417,N_266);
or U7827 (N_7827,N_3521,N_4151);
nor U7828 (N_7828,N_4379,N_4527);
nand U7829 (N_7829,N_3858,N_2122);
and U7830 (N_7830,N_2592,N_3483);
and U7831 (N_7831,N_4291,N_3241);
nor U7832 (N_7832,N_2510,N_2958);
xor U7833 (N_7833,N_4228,N_2842);
nand U7834 (N_7834,N_3869,N_340);
nand U7835 (N_7835,N_830,N_931);
nor U7836 (N_7836,N_4339,N_2980);
or U7837 (N_7837,N_220,N_266);
or U7838 (N_7838,N_4410,N_2718);
xor U7839 (N_7839,N_4209,N_4099);
nand U7840 (N_7840,N_2186,N_789);
nand U7841 (N_7841,N_3722,N_82);
nor U7842 (N_7842,N_1889,N_1666);
nor U7843 (N_7843,N_2691,N_2454);
nand U7844 (N_7844,N_145,N_1046);
nand U7845 (N_7845,N_2451,N_3340);
and U7846 (N_7846,N_848,N_3959);
xor U7847 (N_7847,N_3281,N_4229);
nand U7848 (N_7848,N_1188,N_1576);
or U7849 (N_7849,N_4571,N_159);
and U7850 (N_7850,N_2108,N_4314);
xor U7851 (N_7851,N_385,N_1656);
and U7852 (N_7852,N_384,N_3749);
nand U7853 (N_7853,N_1149,N_4677);
nand U7854 (N_7854,N_4226,N_2256);
nor U7855 (N_7855,N_20,N_4825);
xor U7856 (N_7856,N_3169,N_4590);
or U7857 (N_7857,N_4548,N_3845);
or U7858 (N_7858,N_4977,N_27);
or U7859 (N_7859,N_2151,N_3724);
or U7860 (N_7860,N_593,N_2499);
nand U7861 (N_7861,N_4384,N_4299);
and U7862 (N_7862,N_4875,N_4680);
or U7863 (N_7863,N_2607,N_3385);
nand U7864 (N_7864,N_4702,N_3067);
nand U7865 (N_7865,N_4073,N_3140);
or U7866 (N_7866,N_73,N_3161);
nand U7867 (N_7867,N_1774,N_3126);
or U7868 (N_7868,N_4372,N_4701);
nor U7869 (N_7869,N_500,N_2350);
nand U7870 (N_7870,N_3092,N_3991);
nor U7871 (N_7871,N_4288,N_2490);
nand U7872 (N_7872,N_1011,N_4469);
nand U7873 (N_7873,N_1054,N_1173);
nand U7874 (N_7874,N_3601,N_109);
or U7875 (N_7875,N_354,N_2641);
or U7876 (N_7876,N_1378,N_3526);
nand U7877 (N_7877,N_3030,N_3746);
nand U7878 (N_7878,N_3432,N_3348);
or U7879 (N_7879,N_175,N_4815);
nor U7880 (N_7880,N_4508,N_2210);
and U7881 (N_7881,N_1453,N_1648);
nand U7882 (N_7882,N_3815,N_4489);
and U7883 (N_7883,N_2692,N_4554);
nor U7884 (N_7884,N_1231,N_1696);
and U7885 (N_7885,N_3802,N_740);
or U7886 (N_7886,N_2162,N_1425);
nor U7887 (N_7887,N_1047,N_4937);
nor U7888 (N_7888,N_3244,N_2154);
and U7889 (N_7889,N_1321,N_4944);
nor U7890 (N_7890,N_3263,N_2338);
nand U7891 (N_7891,N_3028,N_2470);
nand U7892 (N_7892,N_353,N_2144);
and U7893 (N_7893,N_491,N_2005);
nand U7894 (N_7894,N_2535,N_4915);
or U7895 (N_7895,N_4439,N_671);
nor U7896 (N_7896,N_1223,N_3219);
and U7897 (N_7897,N_2327,N_4617);
and U7898 (N_7898,N_1924,N_4084);
and U7899 (N_7899,N_3943,N_2488);
and U7900 (N_7900,N_817,N_2157);
nand U7901 (N_7901,N_4275,N_162);
or U7902 (N_7902,N_2819,N_663);
nand U7903 (N_7903,N_3509,N_1324);
nand U7904 (N_7904,N_2584,N_130);
nor U7905 (N_7905,N_2207,N_3818);
or U7906 (N_7906,N_3811,N_1431);
nand U7907 (N_7907,N_3005,N_1518);
or U7908 (N_7908,N_1929,N_3899);
nor U7909 (N_7909,N_585,N_1324);
or U7910 (N_7910,N_4500,N_2233);
nor U7911 (N_7911,N_1060,N_56);
and U7912 (N_7912,N_2319,N_1844);
or U7913 (N_7913,N_1337,N_2770);
xor U7914 (N_7914,N_2313,N_4441);
and U7915 (N_7915,N_4401,N_56);
and U7916 (N_7916,N_1033,N_1073);
and U7917 (N_7917,N_1027,N_1642);
nand U7918 (N_7918,N_14,N_1042);
and U7919 (N_7919,N_2057,N_938);
nor U7920 (N_7920,N_1994,N_4474);
nand U7921 (N_7921,N_1114,N_3506);
and U7922 (N_7922,N_207,N_4687);
xnor U7923 (N_7923,N_1705,N_2550);
nand U7924 (N_7924,N_2139,N_1445);
and U7925 (N_7925,N_3003,N_737);
or U7926 (N_7926,N_4423,N_2448);
nor U7927 (N_7927,N_1404,N_2063);
nand U7928 (N_7928,N_4380,N_1560);
or U7929 (N_7929,N_1315,N_4788);
or U7930 (N_7930,N_1979,N_3930);
nand U7931 (N_7931,N_3377,N_3011);
or U7932 (N_7932,N_2856,N_1504);
or U7933 (N_7933,N_1586,N_3677);
and U7934 (N_7934,N_3598,N_2992);
xor U7935 (N_7935,N_2794,N_1078);
or U7936 (N_7936,N_3162,N_3413);
nor U7937 (N_7937,N_4371,N_666);
or U7938 (N_7938,N_1392,N_3311);
or U7939 (N_7939,N_1141,N_468);
or U7940 (N_7940,N_597,N_2588);
nor U7941 (N_7941,N_1984,N_2777);
and U7942 (N_7942,N_960,N_4798);
and U7943 (N_7943,N_495,N_4171);
or U7944 (N_7944,N_1117,N_4990);
nor U7945 (N_7945,N_3629,N_1037);
nor U7946 (N_7946,N_184,N_4500);
or U7947 (N_7947,N_4554,N_3501);
nand U7948 (N_7948,N_1161,N_661);
or U7949 (N_7949,N_3722,N_2613);
or U7950 (N_7950,N_1942,N_907);
nor U7951 (N_7951,N_1213,N_4879);
and U7952 (N_7952,N_4727,N_2051);
nor U7953 (N_7953,N_1652,N_2916);
nand U7954 (N_7954,N_4660,N_650);
nand U7955 (N_7955,N_3461,N_1286);
or U7956 (N_7956,N_1248,N_3983);
or U7957 (N_7957,N_1991,N_1498);
nor U7958 (N_7958,N_396,N_1572);
and U7959 (N_7959,N_1504,N_4215);
or U7960 (N_7960,N_2667,N_3228);
xor U7961 (N_7961,N_3,N_1221);
nor U7962 (N_7962,N_3670,N_4682);
or U7963 (N_7963,N_13,N_248);
nor U7964 (N_7964,N_653,N_2778);
nor U7965 (N_7965,N_3607,N_4830);
or U7966 (N_7966,N_798,N_64);
nand U7967 (N_7967,N_4905,N_903);
or U7968 (N_7968,N_778,N_926);
and U7969 (N_7969,N_2885,N_1321);
nor U7970 (N_7970,N_1423,N_1016);
nand U7971 (N_7971,N_1916,N_4150);
and U7972 (N_7972,N_274,N_2197);
nand U7973 (N_7973,N_868,N_2973);
or U7974 (N_7974,N_329,N_1771);
and U7975 (N_7975,N_3061,N_2887);
nand U7976 (N_7976,N_2873,N_769);
and U7977 (N_7977,N_3442,N_3880);
and U7978 (N_7978,N_3772,N_3370);
nor U7979 (N_7979,N_4965,N_606);
and U7980 (N_7980,N_643,N_3285);
nor U7981 (N_7981,N_1161,N_1765);
nor U7982 (N_7982,N_3248,N_1260);
nor U7983 (N_7983,N_4968,N_2285);
or U7984 (N_7984,N_4614,N_4256);
nor U7985 (N_7985,N_1664,N_2251);
xnor U7986 (N_7986,N_3232,N_3480);
or U7987 (N_7987,N_4669,N_4319);
nor U7988 (N_7988,N_2589,N_2796);
nand U7989 (N_7989,N_3305,N_92);
nor U7990 (N_7990,N_2735,N_2081);
nand U7991 (N_7991,N_2704,N_479);
or U7992 (N_7992,N_4476,N_2342);
or U7993 (N_7993,N_3788,N_2521);
nor U7994 (N_7994,N_1968,N_1685);
nand U7995 (N_7995,N_4577,N_2947);
xnor U7996 (N_7996,N_3785,N_1111);
and U7997 (N_7997,N_3793,N_3660);
nand U7998 (N_7998,N_576,N_4583);
or U7999 (N_7999,N_1635,N_634);
nand U8000 (N_8000,N_3331,N_3418);
or U8001 (N_8001,N_4227,N_4463);
xnor U8002 (N_8002,N_2852,N_3168);
nand U8003 (N_8003,N_2842,N_4655);
nor U8004 (N_8004,N_2085,N_3387);
xor U8005 (N_8005,N_545,N_4239);
or U8006 (N_8006,N_82,N_2215);
or U8007 (N_8007,N_2801,N_3781);
nand U8008 (N_8008,N_2967,N_756);
or U8009 (N_8009,N_3106,N_2007);
nand U8010 (N_8010,N_1271,N_815);
xnor U8011 (N_8011,N_1374,N_1547);
nor U8012 (N_8012,N_2587,N_2719);
or U8013 (N_8013,N_40,N_3796);
or U8014 (N_8014,N_853,N_2112);
or U8015 (N_8015,N_3050,N_4123);
and U8016 (N_8016,N_310,N_2908);
and U8017 (N_8017,N_1706,N_4683);
xor U8018 (N_8018,N_861,N_3920);
and U8019 (N_8019,N_3350,N_1203);
xor U8020 (N_8020,N_51,N_3638);
or U8021 (N_8021,N_1483,N_516);
and U8022 (N_8022,N_1967,N_454);
nor U8023 (N_8023,N_1182,N_4580);
nand U8024 (N_8024,N_489,N_4394);
and U8025 (N_8025,N_1971,N_2538);
or U8026 (N_8026,N_1444,N_2282);
or U8027 (N_8027,N_305,N_1221);
and U8028 (N_8028,N_4256,N_1582);
or U8029 (N_8029,N_4590,N_246);
and U8030 (N_8030,N_1768,N_4059);
nand U8031 (N_8031,N_1279,N_1478);
or U8032 (N_8032,N_1025,N_1642);
nand U8033 (N_8033,N_4371,N_254);
nor U8034 (N_8034,N_1046,N_4866);
nand U8035 (N_8035,N_2166,N_4759);
xor U8036 (N_8036,N_1164,N_4403);
xnor U8037 (N_8037,N_1039,N_443);
and U8038 (N_8038,N_564,N_463);
or U8039 (N_8039,N_1810,N_4133);
nand U8040 (N_8040,N_1912,N_834);
nand U8041 (N_8041,N_3490,N_4802);
and U8042 (N_8042,N_3651,N_4826);
and U8043 (N_8043,N_4947,N_3557);
or U8044 (N_8044,N_4174,N_3081);
or U8045 (N_8045,N_1960,N_2199);
and U8046 (N_8046,N_665,N_2919);
and U8047 (N_8047,N_725,N_4057);
and U8048 (N_8048,N_684,N_4509);
or U8049 (N_8049,N_1542,N_2026);
and U8050 (N_8050,N_4861,N_3849);
nor U8051 (N_8051,N_1655,N_1391);
nand U8052 (N_8052,N_1302,N_2296);
or U8053 (N_8053,N_630,N_3659);
nor U8054 (N_8054,N_594,N_1824);
nand U8055 (N_8055,N_2394,N_4660);
or U8056 (N_8056,N_1713,N_2503);
and U8057 (N_8057,N_850,N_2049);
or U8058 (N_8058,N_621,N_3036);
or U8059 (N_8059,N_2092,N_4272);
nand U8060 (N_8060,N_1575,N_1288);
and U8061 (N_8061,N_3642,N_95);
or U8062 (N_8062,N_2672,N_3371);
nor U8063 (N_8063,N_873,N_4705);
or U8064 (N_8064,N_1254,N_4459);
or U8065 (N_8065,N_2486,N_2582);
xnor U8066 (N_8066,N_4702,N_1966);
or U8067 (N_8067,N_2377,N_267);
nand U8068 (N_8068,N_4450,N_4351);
nand U8069 (N_8069,N_3397,N_2155);
xor U8070 (N_8070,N_2871,N_2110);
or U8071 (N_8071,N_2399,N_3295);
or U8072 (N_8072,N_1013,N_4112);
xor U8073 (N_8073,N_1560,N_1923);
nand U8074 (N_8074,N_3670,N_354);
nand U8075 (N_8075,N_2033,N_4760);
and U8076 (N_8076,N_4500,N_4287);
xor U8077 (N_8077,N_3933,N_2857);
and U8078 (N_8078,N_3791,N_3592);
and U8079 (N_8079,N_2465,N_750);
nor U8080 (N_8080,N_2425,N_4524);
nand U8081 (N_8081,N_694,N_888);
or U8082 (N_8082,N_1364,N_2456);
nor U8083 (N_8083,N_3685,N_1723);
and U8084 (N_8084,N_3637,N_3640);
nor U8085 (N_8085,N_1753,N_102);
xor U8086 (N_8086,N_3428,N_4274);
nor U8087 (N_8087,N_1542,N_2843);
nand U8088 (N_8088,N_3869,N_4548);
nor U8089 (N_8089,N_1597,N_3310);
or U8090 (N_8090,N_3085,N_350);
nor U8091 (N_8091,N_4758,N_3859);
and U8092 (N_8092,N_1982,N_4450);
nand U8093 (N_8093,N_149,N_1325);
or U8094 (N_8094,N_2075,N_1934);
nand U8095 (N_8095,N_3505,N_2830);
nand U8096 (N_8096,N_3715,N_2284);
and U8097 (N_8097,N_4682,N_4433);
xor U8098 (N_8098,N_1805,N_305);
nor U8099 (N_8099,N_2189,N_1388);
nor U8100 (N_8100,N_4709,N_698);
nor U8101 (N_8101,N_2848,N_2408);
xor U8102 (N_8102,N_1297,N_3619);
and U8103 (N_8103,N_276,N_1764);
and U8104 (N_8104,N_3267,N_2160);
or U8105 (N_8105,N_299,N_2520);
nand U8106 (N_8106,N_212,N_1712);
or U8107 (N_8107,N_2081,N_3949);
nor U8108 (N_8108,N_2903,N_4101);
nand U8109 (N_8109,N_1756,N_1767);
and U8110 (N_8110,N_1302,N_3309);
and U8111 (N_8111,N_2390,N_3338);
and U8112 (N_8112,N_4575,N_2522);
xor U8113 (N_8113,N_1700,N_217);
nor U8114 (N_8114,N_375,N_1232);
and U8115 (N_8115,N_284,N_2350);
or U8116 (N_8116,N_941,N_3948);
nor U8117 (N_8117,N_3539,N_3781);
nor U8118 (N_8118,N_4570,N_389);
nor U8119 (N_8119,N_2928,N_3381);
xor U8120 (N_8120,N_2946,N_3568);
nand U8121 (N_8121,N_2619,N_2367);
and U8122 (N_8122,N_3174,N_2358);
nand U8123 (N_8123,N_3674,N_4128);
or U8124 (N_8124,N_1307,N_2294);
nand U8125 (N_8125,N_2880,N_371);
and U8126 (N_8126,N_2066,N_3739);
and U8127 (N_8127,N_3614,N_1038);
and U8128 (N_8128,N_3360,N_4345);
nand U8129 (N_8129,N_4097,N_569);
nor U8130 (N_8130,N_2055,N_59);
xor U8131 (N_8131,N_1646,N_3720);
nor U8132 (N_8132,N_2158,N_3514);
or U8133 (N_8133,N_4088,N_710);
and U8134 (N_8134,N_1665,N_2567);
nand U8135 (N_8135,N_2647,N_412);
nand U8136 (N_8136,N_4817,N_4684);
nand U8137 (N_8137,N_261,N_2215);
xor U8138 (N_8138,N_4154,N_428);
and U8139 (N_8139,N_307,N_2165);
or U8140 (N_8140,N_1934,N_927);
and U8141 (N_8141,N_730,N_4782);
nor U8142 (N_8142,N_3069,N_3626);
or U8143 (N_8143,N_646,N_2077);
nor U8144 (N_8144,N_383,N_4674);
nand U8145 (N_8145,N_4107,N_4941);
xor U8146 (N_8146,N_4890,N_4066);
xnor U8147 (N_8147,N_2005,N_4481);
or U8148 (N_8148,N_4750,N_4873);
nand U8149 (N_8149,N_2109,N_4747);
and U8150 (N_8150,N_186,N_390);
nor U8151 (N_8151,N_4036,N_3904);
and U8152 (N_8152,N_745,N_4131);
nor U8153 (N_8153,N_3165,N_4550);
and U8154 (N_8154,N_1087,N_3323);
nor U8155 (N_8155,N_1223,N_4695);
nand U8156 (N_8156,N_670,N_2585);
and U8157 (N_8157,N_392,N_2895);
xor U8158 (N_8158,N_3283,N_14);
and U8159 (N_8159,N_2318,N_3644);
or U8160 (N_8160,N_3406,N_370);
nand U8161 (N_8161,N_2108,N_3323);
and U8162 (N_8162,N_4424,N_3988);
and U8163 (N_8163,N_3899,N_3787);
or U8164 (N_8164,N_3292,N_3665);
or U8165 (N_8165,N_310,N_2530);
and U8166 (N_8166,N_1983,N_699);
nand U8167 (N_8167,N_2061,N_632);
and U8168 (N_8168,N_3310,N_2616);
or U8169 (N_8169,N_4667,N_1631);
nand U8170 (N_8170,N_327,N_2496);
nand U8171 (N_8171,N_526,N_424);
nand U8172 (N_8172,N_943,N_622);
nand U8173 (N_8173,N_1403,N_4748);
nand U8174 (N_8174,N_344,N_3760);
nor U8175 (N_8175,N_1368,N_4600);
or U8176 (N_8176,N_2310,N_1825);
nor U8177 (N_8177,N_3381,N_857);
nor U8178 (N_8178,N_1079,N_933);
and U8179 (N_8179,N_4102,N_598);
nand U8180 (N_8180,N_2207,N_3651);
xor U8181 (N_8181,N_670,N_2881);
nand U8182 (N_8182,N_3350,N_804);
nand U8183 (N_8183,N_451,N_3505);
nand U8184 (N_8184,N_2096,N_2178);
or U8185 (N_8185,N_2276,N_1339);
or U8186 (N_8186,N_1955,N_3789);
and U8187 (N_8187,N_101,N_3796);
and U8188 (N_8188,N_2344,N_3545);
nor U8189 (N_8189,N_4893,N_256);
or U8190 (N_8190,N_4837,N_3345);
nor U8191 (N_8191,N_4139,N_3057);
and U8192 (N_8192,N_4846,N_3661);
nand U8193 (N_8193,N_201,N_2026);
or U8194 (N_8194,N_274,N_2623);
nand U8195 (N_8195,N_4589,N_3144);
nor U8196 (N_8196,N_4560,N_2840);
and U8197 (N_8197,N_1881,N_3042);
nand U8198 (N_8198,N_486,N_1352);
nand U8199 (N_8199,N_445,N_4650);
nor U8200 (N_8200,N_2913,N_4837);
nand U8201 (N_8201,N_607,N_1791);
nand U8202 (N_8202,N_1730,N_829);
and U8203 (N_8203,N_3983,N_262);
xnor U8204 (N_8204,N_465,N_3971);
nor U8205 (N_8205,N_2283,N_4517);
or U8206 (N_8206,N_3087,N_4457);
xnor U8207 (N_8207,N_1330,N_4825);
nor U8208 (N_8208,N_160,N_659);
or U8209 (N_8209,N_3201,N_2708);
nand U8210 (N_8210,N_3242,N_531);
and U8211 (N_8211,N_1789,N_176);
or U8212 (N_8212,N_2353,N_2323);
and U8213 (N_8213,N_4929,N_1880);
or U8214 (N_8214,N_1500,N_3729);
nand U8215 (N_8215,N_1923,N_3898);
nand U8216 (N_8216,N_199,N_3142);
nand U8217 (N_8217,N_4352,N_787);
xnor U8218 (N_8218,N_1186,N_3038);
and U8219 (N_8219,N_1277,N_989);
or U8220 (N_8220,N_3616,N_2479);
nor U8221 (N_8221,N_4621,N_4406);
or U8222 (N_8222,N_2716,N_4265);
and U8223 (N_8223,N_124,N_2885);
or U8224 (N_8224,N_792,N_2306);
and U8225 (N_8225,N_4676,N_4907);
nor U8226 (N_8226,N_3628,N_728);
nand U8227 (N_8227,N_24,N_4266);
nand U8228 (N_8228,N_2076,N_2315);
nor U8229 (N_8229,N_1343,N_4696);
nand U8230 (N_8230,N_1682,N_2818);
and U8231 (N_8231,N_2976,N_4588);
nand U8232 (N_8232,N_1788,N_3818);
or U8233 (N_8233,N_4232,N_1446);
or U8234 (N_8234,N_3892,N_514);
or U8235 (N_8235,N_1157,N_4462);
and U8236 (N_8236,N_1546,N_2904);
nor U8237 (N_8237,N_1649,N_1541);
nand U8238 (N_8238,N_2175,N_1460);
or U8239 (N_8239,N_1608,N_827);
nor U8240 (N_8240,N_2889,N_1226);
nor U8241 (N_8241,N_4936,N_4119);
and U8242 (N_8242,N_4739,N_1229);
nor U8243 (N_8243,N_584,N_624);
nor U8244 (N_8244,N_2103,N_1869);
nand U8245 (N_8245,N_1318,N_3607);
nand U8246 (N_8246,N_2536,N_2196);
or U8247 (N_8247,N_1227,N_1845);
and U8248 (N_8248,N_1903,N_1944);
or U8249 (N_8249,N_238,N_1319);
xor U8250 (N_8250,N_811,N_3902);
xor U8251 (N_8251,N_953,N_803);
nand U8252 (N_8252,N_1490,N_4155);
or U8253 (N_8253,N_3863,N_1716);
nand U8254 (N_8254,N_2620,N_3515);
and U8255 (N_8255,N_3766,N_3567);
nor U8256 (N_8256,N_4084,N_3550);
nor U8257 (N_8257,N_3592,N_2014);
nand U8258 (N_8258,N_1256,N_1065);
or U8259 (N_8259,N_413,N_2760);
nand U8260 (N_8260,N_4480,N_3338);
xor U8261 (N_8261,N_1669,N_4748);
nand U8262 (N_8262,N_2157,N_4932);
or U8263 (N_8263,N_1762,N_3858);
or U8264 (N_8264,N_1585,N_3500);
xnor U8265 (N_8265,N_2635,N_1445);
xor U8266 (N_8266,N_1120,N_3282);
nor U8267 (N_8267,N_4607,N_3953);
and U8268 (N_8268,N_4980,N_4392);
nand U8269 (N_8269,N_4262,N_3203);
nor U8270 (N_8270,N_1365,N_1145);
nor U8271 (N_8271,N_3636,N_4290);
nand U8272 (N_8272,N_1456,N_933);
nand U8273 (N_8273,N_2299,N_4824);
nor U8274 (N_8274,N_1714,N_509);
and U8275 (N_8275,N_4013,N_4206);
and U8276 (N_8276,N_4996,N_4573);
and U8277 (N_8277,N_2300,N_3313);
nand U8278 (N_8278,N_2624,N_2833);
or U8279 (N_8279,N_1239,N_1123);
nor U8280 (N_8280,N_1656,N_700);
or U8281 (N_8281,N_2600,N_2559);
or U8282 (N_8282,N_2699,N_1266);
and U8283 (N_8283,N_3494,N_3486);
xor U8284 (N_8284,N_1828,N_605);
and U8285 (N_8285,N_2936,N_4830);
or U8286 (N_8286,N_595,N_1915);
nor U8287 (N_8287,N_1979,N_4542);
nand U8288 (N_8288,N_3497,N_4065);
or U8289 (N_8289,N_3505,N_3811);
nand U8290 (N_8290,N_3156,N_4416);
nand U8291 (N_8291,N_3163,N_1836);
nor U8292 (N_8292,N_2038,N_3512);
and U8293 (N_8293,N_855,N_2597);
xnor U8294 (N_8294,N_4340,N_3607);
xnor U8295 (N_8295,N_2994,N_452);
xnor U8296 (N_8296,N_898,N_973);
and U8297 (N_8297,N_168,N_1566);
xor U8298 (N_8298,N_2772,N_1909);
nor U8299 (N_8299,N_2043,N_2797);
nand U8300 (N_8300,N_162,N_4676);
nor U8301 (N_8301,N_4425,N_784);
xnor U8302 (N_8302,N_2589,N_3395);
nor U8303 (N_8303,N_4565,N_864);
xnor U8304 (N_8304,N_3843,N_1545);
nor U8305 (N_8305,N_2661,N_824);
and U8306 (N_8306,N_4543,N_1356);
xnor U8307 (N_8307,N_3022,N_1931);
or U8308 (N_8308,N_4411,N_1531);
nand U8309 (N_8309,N_2678,N_3759);
nand U8310 (N_8310,N_4705,N_1615);
and U8311 (N_8311,N_4367,N_1296);
xor U8312 (N_8312,N_4088,N_3546);
and U8313 (N_8313,N_636,N_2950);
nor U8314 (N_8314,N_791,N_3397);
or U8315 (N_8315,N_3490,N_2555);
nor U8316 (N_8316,N_2237,N_1397);
nand U8317 (N_8317,N_3095,N_3884);
xnor U8318 (N_8318,N_1012,N_4581);
nor U8319 (N_8319,N_4872,N_1902);
nor U8320 (N_8320,N_991,N_4172);
or U8321 (N_8321,N_2676,N_3636);
and U8322 (N_8322,N_431,N_4776);
nand U8323 (N_8323,N_3197,N_2114);
and U8324 (N_8324,N_2127,N_4649);
or U8325 (N_8325,N_4868,N_2081);
or U8326 (N_8326,N_4583,N_2356);
nor U8327 (N_8327,N_640,N_2469);
and U8328 (N_8328,N_940,N_1733);
and U8329 (N_8329,N_2859,N_2523);
nand U8330 (N_8330,N_999,N_773);
nand U8331 (N_8331,N_4341,N_3811);
nand U8332 (N_8332,N_1650,N_3164);
nor U8333 (N_8333,N_4284,N_1744);
nand U8334 (N_8334,N_1544,N_1435);
and U8335 (N_8335,N_4429,N_4821);
and U8336 (N_8336,N_364,N_2886);
and U8337 (N_8337,N_4630,N_446);
xor U8338 (N_8338,N_4056,N_1481);
and U8339 (N_8339,N_2550,N_805);
nor U8340 (N_8340,N_669,N_1935);
nor U8341 (N_8341,N_4803,N_4055);
nand U8342 (N_8342,N_1141,N_644);
nor U8343 (N_8343,N_1194,N_864);
nor U8344 (N_8344,N_661,N_361);
nand U8345 (N_8345,N_1529,N_2504);
nor U8346 (N_8346,N_3184,N_3860);
and U8347 (N_8347,N_1064,N_1155);
and U8348 (N_8348,N_2981,N_4066);
and U8349 (N_8349,N_1317,N_3174);
nor U8350 (N_8350,N_2972,N_1042);
xor U8351 (N_8351,N_3613,N_1738);
nor U8352 (N_8352,N_3629,N_2566);
or U8353 (N_8353,N_2972,N_754);
nand U8354 (N_8354,N_3154,N_769);
nand U8355 (N_8355,N_1858,N_4552);
and U8356 (N_8356,N_3679,N_2157);
nor U8357 (N_8357,N_2252,N_3313);
and U8358 (N_8358,N_59,N_1223);
xnor U8359 (N_8359,N_802,N_774);
xor U8360 (N_8360,N_836,N_4155);
or U8361 (N_8361,N_2510,N_2830);
nand U8362 (N_8362,N_1501,N_804);
or U8363 (N_8363,N_335,N_2887);
nand U8364 (N_8364,N_2845,N_4298);
and U8365 (N_8365,N_4235,N_1682);
nor U8366 (N_8366,N_1561,N_3370);
or U8367 (N_8367,N_1446,N_3456);
or U8368 (N_8368,N_417,N_2575);
and U8369 (N_8369,N_41,N_2224);
nor U8370 (N_8370,N_3643,N_1010);
nand U8371 (N_8371,N_3784,N_4386);
nand U8372 (N_8372,N_3761,N_4563);
and U8373 (N_8373,N_3940,N_2457);
nand U8374 (N_8374,N_2477,N_4652);
or U8375 (N_8375,N_4818,N_4579);
or U8376 (N_8376,N_4996,N_4376);
nor U8377 (N_8377,N_2687,N_3723);
or U8378 (N_8378,N_4281,N_2995);
and U8379 (N_8379,N_3829,N_2318);
nor U8380 (N_8380,N_534,N_2256);
and U8381 (N_8381,N_3768,N_1802);
or U8382 (N_8382,N_2616,N_197);
nor U8383 (N_8383,N_1465,N_4921);
xor U8384 (N_8384,N_4844,N_2885);
and U8385 (N_8385,N_3627,N_2572);
and U8386 (N_8386,N_3520,N_937);
and U8387 (N_8387,N_3611,N_4278);
nor U8388 (N_8388,N_3777,N_1162);
nor U8389 (N_8389,N_1672,N_4643);
nand U8390 (N_8390,N_3457,N_3360);
xor U8391 (N_8391,N_4068,N_1667);
or U8392 (N_8392,N_1882,N_3461);
or U8393 (N_8393,N_3705,N_284);
nor U8394 (N_8394,N_3550,N_452);
and U8395 (N_8395,N_994,N_3905);
or U8396 (N_8396,N_4180,N_3315);
nor U8397 (N_8397,N_3503,N_4525);
and U8398 (N_8398,N_3982,N_569);
or U8399 (N_8399,N_155,N_650);
or U8400 (N_8400,N_1065,N_828);
nand U8401 (N_8401,N_4326,N_4658);
nor U8402 (N_8402,N_2081,N_3734);
nor U8403 (N_8403,N_1120,N_2299);
and U8404 (N_8404,N_1787,N_3110);
xor U8405 (N_8405,N_620,N_2240);
xor U8406 (N_8406,N_2532,N_354);
xnor U8407 (N_8407,N_2124,N_3613);
nor U8408 (N_8408,N_1915,N_4490);
and U8409 (N_8409,N_1170,N_2647);
or U8410 (N_8410,N_1676,N_2289);
nor U8411 (N_8411,N_1735,N_3480);
nand U8412 (N_8412,N_1878,N_3352);
nor U8413 (N_8413,N_293,N_950);
nand U8414 (N_8414,N_407,N_1487);
nor U8415 (N_8415,N_1460,N_1638);
or U8416 (N_8416,N_69,N_1643);
or U8417 (N_8417,N_1197,N_356);
nor U8418 (N_8418,N_1421,N_250);
nor U8419 (N_8419,N_4991,N_3078);
or U8420 (N_8420,N_3778,N_1045);
and U8421 (N_8421,N_702,N_3517);
and U8422 (N_8422,N_3438,N_4836);
and U8423 (N_8423,N_3097,N_4176);
nand U8424 (N_8424,N_3534,N_383);
and U8425 (N_8425,N_3026,N_2025);
nor U8426 (N_8426,N_1864,N_2168);
nor U8427 (N_8427,N_4172,N_4040);
and U8428 (N_8428,N_2260,N_3022);
and U8429 (N_8429,N_589,N_3235);
and U8430 (N_8430,N_2773,N_265);
xnor U8431 (N_8431,N_4192,N_3948);
nand U8432 (N_8432,N_4966,N_4311);
nor U8433 (N_8433,N_2562,N_2176);
and U8434 (N_8434,N_95,N_1616);
nand U8435 (N_8435,N_3882,N_2963);
and U8436 (N_8436,N_1362,N_1794);
xnor U8437 (N_8437,N_1635,N_3686);
nand U8438 (N_8438,N_751,N_1126);
and U8439 (N_8439,N_1205,N_491);
nand U8440 (N_8440,N_4718,N_3814);
xnor U8441 (N_8441,N_2125,N_3753);
xnor U8442 (N_8442,N_4665,N_1859);
or U8443 (N_8443,N_4554,N_4);
nor U8444 (N_8444,N_1461,N_3923);
nand U8445 (N_8445,N_126,N_4379);
nand U8446 (N_8446,N_4535,N_2190);
or U8447 (N_8447,N_4479,N_1378);
nor U8448 (N_8448,N_330,N_3053);
or U8449 (N_8449,N_3421,N_3894);
nor U8450 (N_8450,N_1397,N_4620);
or U8451 (N_8451,N_2364,N_264);
nand U8452 (N_8452,N_4486,N_2950);
and U8453 (N_8453,N_3786,N_4063);
xor U8454 (N_8454,N_3799,N_738);
xor U8455 (N_8455,N_2331,N_3518);
xnor U8456 (N_8456,N_908,N_3216);
nor U8457 (N_8457,N_974,N_4073);
and U8458 (N_8458,N_1897,N_843);
or U8459 (N_8459,N_4670,N_2125);
nand U8460 (N_8460,N_572,N_4139);
nor U8461 (N_8461,N_524,N_2185);
xnor U8462 (N_8462,N_1539,N_1073);
or U8463 (N_8463,N_2278,N_3466);
nor U8464 (N_8464,N_4189,N_3472);
nor U8465 (N_8465,N_2797,N_87);
xnor U8466 (N_8466,N_2536,N_732);
nand U8467 (N_8467,N_4106,N_1615);
nor U8468 (N_8468,N_4719,N_1456);
nand U8469 (N_8469,N_2335,N_1152);
nor U8470 (N_8470,N_4911,N_3686);
nor U8471 (N_8471,N_2042,N_2358);
or U8472 (N_8472,N_2041,N_2114);
nor U8473 (N_8473,N_3696,N_3721);
or U8474 (N_8474,N_4657,N_3124);
nand U8475 (N_8475,N_2924,N_1178);
nor U8476 (N_8476,N_3083,N_799);
or U8477 (N_8477,N_2621,N_4064);
and U8478 (N_8478,N_1935,N_4479);
nor U8479 (N_8479,N_157,N_4905);
nor U8480 (N_8480,N_2780,N_2393);
nor U8481 (N_8481,N_4006,N_2534);
or U8482 (N_8482,N_1886,N_2531);
nor U8483 (N_8483,N_3177,N_1022);
or U8484 (N_8484,N_4609,N_1311);
nor U8485 (N_8485,N_3289,N_3871);
nor U8486 (N_8486,N_2356,N_1842);
and U8487 (N_8487,N_3118,N_1204);
and U8488 (N_8488,N_1145,N_3076);
nand U8489 (N_8489,N_231,N_4458);
nand U8490 (N_8490,N_1768,N_3200);
nor U8491 (N_8491,N_4234,N_2724);
or U8492 (N_8492,N_4405,N_715);
nand U8493 (N_8493,N_1348,N_1011);
and U8494 (N_8494,N_2607,N_2957);
and U8495 (N_8495,N_758,N_192);
nand U8496 (N_8496,N_4518,N_1171);
or U8497 (N_8497,N_776,N_3986);
xor U8498 (N_8498,N_2700,N_2761);
nand U8499 (N_8499,N_6,N_1297);
or U8500 (N_8500,N_4100,N_4198);
nor U8501 (N_8501,N_3499,N_2720);
nor U8502 (N_8502,N_47,N_3575);
and U8503 (N_8503,N_967,N_4482);
xor U8504 (N_8504,N_3982,N_1927);
nor U8505 (N_8505,N_3783,N_9);
and U8506 (N_8506,N_809,N_3879);
nand U8507 (N_8507,N_4031,N_2538);
nor U8508 (N_8508,N_434,N_4613);
nor U8509 (N_8509,N_3535,N_1636);
nand U8510 (N_8510,N_1017,N_813);
or U8511 (N_8511,N_4596,N_317);
or U8512 (N_8512,N_2822,N_1778);
nand U8513 (N_8513,N_2992,N_3207);
nand U8514 (N_8514,N_3512,N_1774);
or U8515 (N_8515,N_2930,N_1898);
nor U8516 (N_8516,N_4360,N_4437);
and U8517 (N_8517,N_3397,N_564);
xnor U8518 (N_8518,N_1621,N_2755);
nor U8519 (N_8519,N_1053,N_4443);
nand U8520 (N_8520,N_2124,N_3436);
or U8521 (N_8521,N_1646,N_2023);
nand U8522 (N_8522,N_4070,N_4756);
and U8523 (N_8523,N_194,N_1081);
or U8524 (N_8524,N_1783,N_2955);
and U8525 (N_8525,N_2613,N_4959);
or U8526 (N_8526,N_2658,N_4953);
nand U8527 (N_8527,N_2435,N_4413);
nand U8528 (N_8528,N_239,N_2261);
nor U8529 (N_8529,N_3736,N_3311);
and U8530 (N_8530,N_4479,N_1270);
and U8531 (N_8531,N_2476,N_3613);
nand U8532 (N_8532,N_82,N_4759);
nand U8533 (N_8533,N_260,N_921);
nor U8534 (N_8534,N_4705,N_3369);
nand U8535 (N_8535,N_193,N_1258);
or U8536 (N_8536,N_2369,N_3408);
nand U8537 (N_8537,N_3898,N_2489);
and U8538 (N_8538,N_1511,N_1256);
xor U8539 (N_8539,N_1963,N_1498);
or U8540 (N_8540,N_1821,N_4131);
or U8541 (N_8541,N_2824,N_3681);
or U8542 (N_8542,N_1325,N_1692);
and U8543 (N_8543,N_4394,N_4121);
nor U8544 (N_8544,N_2978,N_3098);
nand U8545 (N_8545,N_1811,N_1365);
nor U8546 (N_8546,N_4433,N_4335);
xor U8547 (N_8547,N_3223,N_1874);
or U8548 (N_8548,N_1223,N_4678);
nor U8549 (N_8549,N_746,N_842);
xnor U8550 (N_8550,N_2588,N_2221);
nor U8551 (N_8551,N_3237,N_2054);
nor U8552 (N_8552,N_3074,N_0);
or U8553 (N_8553,N_908,N_522);
and U8554 (N_8554,N_3379,N_3552);
or U8555 (N_8555,N_2670,N_2862);
nor U8556 (N_8556,N_3838,N_4717);
nor U8557 (N_8557,N_1375,N_4805);
nand U8558 (N_8558,N_3820,N_294);
nor U8559 (N_8559,N_733,N_572);
or U8560 (N_8560,N_3611,N_1507);
and U8561 (N_8561,N_2673,N_306);
nand U8562 (N_8562,N_4154,N_4877);
xnor U8563 (N_8563,N_445,N_4831);
and U8564 (N_8564,N_953,N_4815);
and U8565 (N_8565,N_3151,N_4763);
nor U8566 (N_8566,N_2843,N_512);
nand U8567 (N_8567,N_3144,N_2481);
nor U8568 (N_8568,N_1979,N_768);
and U8569 (N_8569,N_2706,N_2985);
nor U8570 (N_8570,N_1457,N_186);
nand U8571 (N_8571,N_314,N_3067);
or U8572 (N_8572,N_544,N_1854);
or U8573 (N_8573,N_1677,N_1375);
nor U8574 (N_8574,N_2894,N_1658);
xnor U8575 (N_8575,N_282,N_2702);
nand U8576 (N_8576,N_1200,N_3902);
or U8577 (N_8577,N_1601,N_1448);
nor U8578 (N_8578,N_1436,N_3875);
and U8579 (N_8579,N_466,N_307);
and U8580 (N_8580,N_3351,N_2745);
and U8581 (N_8581,N_56,N_181);
nor U8582 (N_8582,N_2472,N_4035);
nand U8583 (N_8583,N_1942,N_345);
nor U8584 (N_8584,N_1539,N_2226);
nand U8585 (N_8585,N_2036,N_1610);
nor U8586 (N_8586,N_2685,N_894);
and U8587 (N_8587,N_4975,N_2215);
nand U8588 (N_8588,N_1414,N_1137);
or U8589 (N_8589,N_2704,N_3191);
nand U8590 (N_8590,N_3144,N_2075);
nand U8591 (N_8591,N_1893,N_4093);
or U8592 (N_8592,N_2594,N_42);
and U8593 (N_8593,N_401,N_3962);
or U8594 (N_8594,N_4671,N_4772);
nor U8595 (N_8595,N_1300,N_3612);
or U8596 (N_8596,N_814,N_941);
and U8597 (N_8597,N_4738,N_3585);
nand U8598 (N_8598,N_3300,N_4010);
or U8599 (N_8599,N_4323,N_3257);
and U8600 (N_8600,N_1731,N_4026);
xor U8601 (N_8601,N_3689,N_3802);
nand U8602 (N_8602,N_4482,N_4395);
or U8603 (N_8603,N_4371,N_3843);
xnor U8604 (N_8604,N_1923,N_4074);
nor U8605 (N_8605,N_1755,N_3968);
nand U8606 (N_8606,N_416,N_1028);
nand U8607 (N_8607,N_857,N_1427);
nand U8608 (N_8608,N_1777,N_1612);
or U8609 (N_8609,N_1797,N_295);
and U8610 (N_8610,N_4768,N_3627);
and U8611 (N_8611,N_4963,N_1873);
xor U8612 (N_8612,N_4140,N_3663);
and U8613 (N_8613,N_2441,N_4027);
or U8614 (N_8614,N_1183,N_2580);
or U8615 (N_8615,N_1221,N_2569);
and U8616 (N_8616,N_4567,N_3837);
nand U8617 (N_8617,N_1515,N_2114);
and U8618 (N_8618,N_2846,N_1244);
nor U8619 (N_8619,N_665,N_2920);
and U8620 (N_8620,N_55,N_4320);
nor U8621 (N_8621,N_3268,N_990);
nor U8622 (N_8622,N_2978,N_2651);
and U8623 (N_8623,N_2880,N_189);
nor U8624 (N_8624,N_1683,N_3195);
and U8625 (N_8625,N_1604,N_1576);
or U8626 (N_8626,N_645,N_2461);
and U8627 (N_8627,N_1795,N_623);
and U8628 (N_8628,N_1851,N_3251);
nand U8629 (N_8629,N_2932,N_3365);
or U8630 (N_8630,N_1735,N_3832);
nand U8631 (N_8631,N_3679,N_3651);
nor U8632 (N_8632,N_4066,N_1748);
xnor U8633 (N_8633,N_2703,N_750);
nand U8634 (N_8634,N_3536,N_2565);
nor U8635 (N_8635,N_4776,N_3599);
nand U8636 (N_8636,N_1918,N_1627);
nor U8637 (N_8637,N_3926,N_1291);
or U8638 (N_8638,N_2898,N_1664);
or U8639 (N_8639,N_1244,N_1665);
or U8640 (N_8640,N_2088,N_510);
nor U8641 (N_8641,N_1916,N_2323);
nor U8642 (N_8642,N_2428,N_2074);
and U8643 (N_8643,N_76,N_4137);
nand U8644 (N_8644,N_4815,N_1788);
and U8645 (N_8645,N_1957,N_3794);
or U8646 (N_8646,N_4596,N_1656);
or U8647 (N_8647,N_2286,N_2150);
nor U8648 (N_8648,N_4420,N_517);
nor U8649 (N_8649,N_2580,N_4168);
nand U8650 (N_8650,N_3197,N_3455);
xor U8651 (N_8651,N_3364,N_3230);
or U8652 (N_8652,N_2340,N_997);
nor U8653 (N_8653,N_1608,N_2147);
nor U8654 (N_8654,N_4646,N_2392);
nor U8655 (N_8655,N_1363,N_2420);
nand U8656 (N_8656,N_2092,N_257);
nand U8657 (N_8657,N_1640,N_1326);
nand U8658 (N_8658,N_4092,N_4729);
xnor U8659 (N_8659,N_4155,N_4972);
nand U8660 (N_8660,N_2902,N_3734);
or U8661 (N_8661,N_1967,N_866);
and U8662 (N_8662,N_2497,N_2532);
nand U8663 (N_8663,N_4421,N_4109);
xor U8664 (N_8664,N_2672,N_580);
xnor U8665 (N_8665,N_2537,N_4988);
nor U8666 (N_8666,N_82,N_2869);
and U8667 (N_8667,N_4654,N_4561);
xnor U8668 (N_8668,N_4159,N_4327);
and U8669 (N_8669,N_4026,N_4644);
nand U8670 (N_8670,N_3641,N_4275);
or U8671 (N_8671,N_59,N_2983);
nor U8672 (N_8672,N_186,N_3798);
xnor U8673 (N_8673,N_1741,N_1411);
nand U8674 (N_8674,N_104,N_3969);
or U8675 (N_8675,N_4620,N_511);
or U8676 (N_8676,N_2854,N_1823);
or U8677 (N_8677,N_483,N_1989);
nor U8678 (N_8678,N_2177,N_1329);
nand U8679 (N_8679,N_3659,N_2351);
and U8680 (N_8680,N_2068,N_877);
nor U8681 (N_8681,N_3875,N_1954);
nand U8682 (N_8682,N_2002,N_3088);
and U8683 (N_8683,N_4745,N_2191);
nand U8684 (N_8684,N_1727,N_3218);
and U8685 (N_8685,N_377,N_3639);
nor U8686 (N_8686,N_4715,N_3848);
nor U8687 (N_8687,N_876,N_4804);
xnor U8688 (N_8688,N_2809,N_3729);
and U8689 (N_8689,N_106,N_3372);
and U8690 (N_8690,N_1970,N_4590);
or U8691 (N_8691,N_2224,N_852);
nor U8692 (N_8692,N_36,N_263);
nand U8693 (N_8693,N_1882,N_3041);
or U8694 (N_8694,N_3674,N_1426);
and U8695 (N_8695,N_648,N_634);
nand U8696 (N_8696,N_4050,N_3887);
nand U8697 (N_8697,N_2947,N_2144);
or U8698 (N_8698,N_3623,N_111);
nor U8699 (N_8699,N_821,N_1952);
nor U8700 (N_8700,N_3127,N_142);
nand U8701 (N_8701,N_3339,N_1976);
or U8702 (N_8702,N_4077,N_2579);
and U8703 (N_8703,N_4362,N_1165);
and U8704 (N_8704,N_2651,N_2948);
nor U8705 (N_8705,N_1739,N_4965);
or U8706 (N_8706,N_3942,N_1807);
nand U8707 (N_8707,N_2994,N_2353);
xnor U8708 (N_8708,N_3816,N_2836);
or U8709 (N_8709,N_2512,N_1355);
or U8710 (N_8710,N_4390,N_359);
nor U8711 (N_8711,N_2002,N_1103);
nand U8712 (N_8712,N_1325,N_1853);
and U8713 (N_8713,N_2528,N_647);
nor U8714 (N_8714,N_1700,N_4947);
and U8715 (N_8715,N_1064,N_1989);
or U8716 (N_8716,N_4424,N_3542);
nor U8717 (N_8717,N_4010,N_4615);
nor U8718 (N_8718,N_2902,N_4133);
nor U8719 (N_8719,N_2297,N_2615);
nor U8720 (N_8720,N_3382,N_786);
or U8721 (N_8721,N_2688,N_3647);
or U8722 (N_8722,N_3652,N_369);
or U8723 (N_8723,N_3510,N_1048);
nor U8724 (N_8724,N_3980,N_193);
xor U8725 (N_8725,N_3951,N_2657);
nor U8726 (N_8726,N_1961,N_852);
and U8727 (N_8727,N_10,N_4302);
nand U8728 (N_8728,N_1249,N_1637);
nor U8729 (N_8729,N_15,N_2582);
nand U8730 (N_8730,N_2356,N_3462);
or U8731 (N_8731,N_4512,N_2448);
nand U8732 (N_8732,N_3374,N_2270);
xor U8733 (N_8733,N_947,N_968);
nand U8734 (N_8734,N_1109,N_1878);
or U8735 (N_8735,N_4184,N_4642);
nor U8736 (N_8736,N_4491,N_1240);
nand U8737 (N_8737,N_4730,N_3714);
xor U8738 (N_8738,N_1632,N_278);
nand U8739 (N_8739,N_96,N_3109);
and U8740 (N_8740,N_1533,N_1169);
nor U8741 (N_8741,N_4622,N_2057);
nand U8742 (N_8742,N_1551,N_1216);
nor U8743 (N_8743,N_2143,N_1119);
and U8744 (N_8744,N_3897,N_2860);
and U8745 (N_8745,N_4572,N_1428);
xor U8746 (N_8746,N_2429,N_2621);
xor U8747 (N_8747,N_3412,N_4750);
nand U8748 (N_8748,N_3797,N_1290);
nand U8749 (N_8749,N_1808,N_2641);
or U8750 (N_8750,N_4447,N_2161);
or U8751 (N_8751,N_2708,N_439);
xnor U8752 (N_8752,N_4236,N_1460);
and U8753 (N_8753,N_3487,N_2002);
nor U8754 (N_8754,N_4912,N_4180);
or U8755 (N_8755,N_4976,N_2022);
and U8756 (N_8756,N_2490,N_3980);
nand U8757 (N_8757,N_1759,N_683);
and U8758 (N_8758,N_1362,N_4265);
nand U8759 (N_8759,N_4345,N_1917);
nor U8760 (N_8760,N_3937,N_4840);
and U8761 (N_8761,N_656,N_3966);
or U8762 (N_8762,N_4941,N_2916);
nor U8763 (N_8763,N_1208,N_1342);
nand U8764 (N_8764,N_3523,N_2008);
and U8765 (N_8765,N_2963,N_4756);
and U8766 (N_8766,N_3402,N_614);
or U8767 (N_8767,N_4394,N_3218);
nand U8768 (N_8768,N_3256,N_2719);
and U8769 (N_8769,N_105,N_859);
and U8770 (N_8770,N_1260,N_2024);
and U8771 (N_8771,N_1893,N_4645);
xnor U8772 (N_8772,N_1177,N_256);
nor U8773 (N_8773,N_77,N_3262);
and U8774 (N_8774,N_800,N_3781);
nand U8775 (N_8775,N_2320,N_1414);
nand U8776 (N_8776,N_4478,N_2158);
nor U8777 (N_8777,N_778,N_1444);
or U8778 (N_8778,N_4185,N_729);
nand U8779 (N_8779,N_1647,N_1878);
or U8780 (N_8780,N_4966,N_3306);
nand U8781 (N_8781,N_1487,N_505);
nand U8782 (N_8782,N_1962,N_2517);
or U8783 (N_8783,N_2782,N_92);
and U8784 (N_8784,N_3836,N_1473);
nor U8785 (N_8785,N_1620,N_91);
nor U8786 (N_8786,N_337,N_2780);
xor U8787 (N_8787,N_471,N_1766);
nand U8788 (N_8788,N_1782,N_1826);
nor U8789 (N_8789,N_3198,N_4722);
or U8790 (N_8790,N_4576,N_3699);
nand U8791 (N_8791,N_1761,N_4805);
xor U8792 (N_8792,N_4004,N_3106);
and U8793 (N_8793,N_196,N_2690);
nand U8794 (N_8794,N_2879,N_1438);
xnor U8795 (N_8795,N_2535,N_4086);
and U8796 (N_8796,N_2314,N_207);
or U8797 (N_8797,N_1022,N_3727);
nor U8798 (N_8798,N_3947,N_806);
and U8799 (N_8799,N_2209,N_15);
nand U8800 (N_8800,N_4201,N_1061);
nand U8801 (N_8801,N_4455,N_4065);
and U8802 (N_8802,N_610,N_3804);
nor U8803 (N_8803,N_1226,N_3238);
nor U8804 (N_8804,N_206,N_4489);
xnor U8805 (N_8805,N_1367,N_907);
xor U8806 (N_8806,N_817,N_1871);
or U8807 (N_8807,N_313,N_2327);
and U8808 (N_8808,N_4665,N_2660);
or U8809 (N_8809,N_3699,N_105);
nand U8810 (N_8810,N_1033,N_4950);
nand U8811 (N_8811,N_1027,N_4058);
and U8812 (N_8812,N_4668,N_3029);
xnor U8813 (N_8813,N_1930,N_2033);
nand U8814 (N_8814,N_2759,N_203);
nor U8815 (N_8815,N_2,N_2342);
nand U8816 (N_8816,N_3874,N_997);
nand U8817 (N_8817,N_3985,N_4830);
and U8818 (N_8818,N_3396,N_3810);
or U8819 (N_8819,N_2795,N_83);
or U8820 (N_8820,N_3316,N_2044);
xnor U8821 (N_8821,N_539,N_2100);
xnor U8822 (N_8822,N_560,N_4208);
nand U8823 (N_8823,N_4948,N_4860);
and U8824 (N_8824,N_3125,N_3346);
and U8825 (N_8825,N_4212,N_2785);
nor U8826 (N_8826,N_823,N_2434);
nor U8827 (N_8827,N_4398,N_3324);
nand U8828 (N_8828,N_1314,N_2051);
nand U8829 (N_8829,N_2802,N_4315);
and U8830 (N_8830,N_1519,N_3616);
xor U8831 (N_8831,N_1669,N_2866);
or U8832 (N_8832,N_4585,N_4683);
or U8833 (N_8833,N_91,N_2111);
xor U8834 (N_8834,N_678,N_2235);
nand U8835 (N_8835,N_2806,N_4285);
nand U8836 (N_8836,N_1700,N_286);
nor U8837 (N_8837,N_1020,N_1216);
nand U8838 (N_8838,N_3934,N_3921);
xnor U8839 (N_8839,N_3427,N_2381);
nor U8840 (N_8840,N_4814,N_1710);
nand U8841 (N_8841,N_866,N_2240);
and U8842 (N_8842,N_4455,N_2611);
and U8843 (N_8843,N_1842,N_2270);
and U8844 (N_8844,N_3819,N_507);
and U8845 (N_8845,N_4307,N_2154);
nor U8846 (N_8846,N_3813,N_2294);
or U8847 (N_8847,N_3159,N_2625);
xnor U8848 (N_8848,N_3106,N_1676);
nor U8849 (N_8849,N_4360,N_4275);
and U8850 (N_8850,N_2442,N_2556);
or U8851 (N_8851,N_1920,N_1686);
nor U8852 (N_8852,N_4566,N_4730);
nor U8853 (N_8853,N_4365,N_2157);
xnor U8854 (N_8854,N_1538,N_2542);
nor U8855 (N_8855,N_4400,N_1160);
nand U8856 (N_8856,N_4866,N_1735);
nand U8857 (N_8857,N_2851,N_242);
or U8858 (N_8858,N_4134,N_644);
or U8859 (N_8859,N_3037,N_3714);
xor U8860 (N_8860,N_4571,N_941);
or U8861 (N_8861,N_1992,N_4332);
and U8862 (N_8862,N_4220,N_4200);
nand U8863 (N_8863,N_4452,N_4851);
nand U8864 (N_8864,N_390,N_2126);
or U8865 (N_8865,N_1271,N_2517);
xor U8866 (N_8866,N_212,N_3727);
nor U8867 (N_8867,N_1478,N_3439);
or U8868 (N_8868,N_1484,N_1381);
xor U8869 (N_8869,N_1247,N_87);
or U8870 (N_8870,N_3679,N_4681);
nor U8871 (N_8871,N_1016,N_3518);
nor U8872 (N_8872,N_569,N_1530);
nand U8873 (N_8873,N_4080,N_2815);
and U8874 (N_8874,N_3654,N_14);
xor U8875 (N_8875,N_4226,N_3911);
nand U8876 (N_8876,N_4489,N_64);
and U8877 (N_8877,N_3663,N_4426);
nand U8878 (N_8878,N_3798,N_4914);
nor U8879 (N_8879,N_545,N_1388);
nand U8880 (N_8880,N_864,N_826);
and U8881 (N_8881,N_4514,N_4627);
nor U8882 (N_8882,N_3755,N_4151);
nor U8883 (N_8883,N_3736,N_22);
and U8884 (N_8884,N_2091,N_4638);
or U8885 (N_8885,N_686,N_1204);
and U8886 (N_8886,N_2610,N_3646);
nor U8887 (N_8887,N_1917,N_1077);
or U8888 (N_8888,N_4680,N_2486);
and U8889 (N_8889,N_3820,N_1827);
and U8890 (N_8890,N_4830,N_3194);
or U8891 (N_8891,N_2684,N_4879);
nand U8892 (N_8892,N_888,N_547);
nand U8893 (N_8893,N_4180,N_3799);
nor U8894 (N_8894,N_4775,N_3009);
or U8895 (N_8895,N_3358,N_4827);
or U8896 (N_8896,N_2395,N_2481);
xor U8897 (N_8897,N_1864,N_68);
or U8898 (N_8898,N_3339,N_1945);
or U8899 (N_8899,N_357,N_4414);
or U8900 (N_8900,N_3431,N_4072);
nand U8901 (N_8901,N_713,N_4622);
or U8902 (N_8902,N_340,N_4272);
or U8903 (N_8903,N_435,N_2487);
nand U8904 (N_8904,N_3795,N_1936);
nand U8905 (N_8905,N_2770,N_635);
nand U8906 (N_8906,N_2637,N_4258);
xnor U8907 (N_8907,N_2746,N_38);
nand U8908 (N_8908,N_4078,N_1613);
or U8909 (N_8909,N_1085,N_1261);
nor U8910 (N_8910,N_4394,N_4636);
nand U8911 (N_8911,N_1462,N_119);
or U8912 (N_8912,N_4176,N_2679);
and U8913 (N_8913,N_2404,N_472);
nor U8914 (N_8914,N_2430,N_2061);
or U8915 (N_8915,N_1260,N_1377);
nand U8916 (N_8916,N_2537,N_4684);
and U8917 (N_8917,N_4644,N_1650);
nor U8918 (N_8918,N_1519,N_3581);
nor U8919 (N_8919,N_2975,N_1875);
nor U8920 (N_8920,N_2243,N_1040);
xnor U8921 (N_8921,N_2938,N_244);
xnor U8922 (N_8922,N_591,N_4264);
nand U8923 (N_8923,N_2677,N_1786);
and U8924 (N_8924,N_1606,N_738);
or U8925 (N_8925,N_4604,N_1847);
nand U8926 (N_8926,N_3741,N_4650);
nand U8927 (N_8927,N_4254,N_883);
and U8928 (N_8928,N_1984,N_2197);
xor U8929 (N_8929,N_4366,N_3342);
nand U8930 (N_8930,N_1570,N_602);
xor U8931 (N_8931,N_1844,N_3771);
nor U8932 (N_8932,N_2265,N_1668);
xnor U8933 (N_8933,N_2171,N_1892);
nand U8934 (N_8934,N_1115,N_1648);
and U8935 (N_8935,N_2342,N_4837);
nand U8936 (N_8936,N_2547,N_1655);
nor U8937 (N_8937,N_2394,N_3611);
nand U8938 (N_8938,N_3451,N_2039);
and U8939 (N_8939,N_3554,N_2180);
nor U8940 (N_8940,N_3769,N_4814);
nand U8941 (N_8941,N_2390,N_4798);
or U8942 (N_8942,N_214,N_243);
nor U8943 (N_8943,N_3449,N_1928);
and U8944 (N_8944,N_1972,N_2487);
or U8945 (N_8945,N_990,N_2605);
or U8946 (N_8946,N_854,N_1875);
nor U8947 (N_8947,N_2587,N_3532);
and U8948 (N_8948,N_2589,N_603);
nor U8949 (N_8949,N_2779,N_4930);
or U8950 (N_8950,N_3060,N_2132);
xor U8951 (N_8951,N_4486,N_569);
nor U8952 (N_8952,N_2750,N_4614);
nor U8953 (N_8953,N_2889,N_2164);
xor U8954 (N_8954,N_3696,N_1481);
nor U8955 (N_8955,N_4379,N_3154);
xnor U8956 (N_8956,N_4796,N_295);
nand U8957 (N_8957,N_1445,N_3112);
nand U8958 (N_8958,N_3537,N_4216);
xnor U8959 (N_8959,N_2173,N_2379);
nand U8960 (N_8960,N_4341,N_367);
or U8961 (N_8961,N_610,N_3147);
nand U8962 (N_8962,N_464,N_2200);
xnor U8963 (N_8963,N_792,N_769);
nand U8964 (N_8964,N_2518,N_3323);
and U8965 (N_8965,N_1933,N_3152);
and U8966 (N_8966,N_3109,N_156);
nor U8967 (N_8967,N_328,N_3235);
and U8968 (N_8968,N_4778,N_785);
and U8969 (N_8969,N_2407,N_1385);
nand U8970 (N_8970,N_2543,N_1738);
nand U8971 (N_8971,N_160,N_3642);
or U8972 (N_8972,N_3826,N_4414);
xnor U8973 (N_8973,N_3885,N_953);
nor U8974 (N_8974,N_3069,N_2340);
nand U8975 (N_8975,N_117,N_4148);
xnor U8976 (N_8976,N_1576,N_302);
and U8977 (N_8977,N_512,N_3491);
xnor U8978 (N_8978,N_650,N_364);
nor U8979 (N_8979,N_1844,N_2567);
nor U8980 (N_8980,N_3265,N_2777);
and U8981 (N_8981,N_2544,N_4065);
or U8982 (N_8982,N_1269,N_2612);
xor U8983 (N_8983,N_466,N_714);
nor U8984 (N_8984,N_3146,N_2413);
and U8985 (N_8985,N_4979,N_4658);
nor U8986 (N_8986,N_272,N_1025);
or U8987 (N_8987,N_1902,N_720);
nand U8988 (N_8988,N_2601,N_586);
nand U8989 (N_8989,N_1736,N_1745);
xor U8990 (N_8990,N_1406,N_2659);
and U8991 (N_8991,N_1274,N_1084);
nand U8992 (N_8992,N_3037,N_4851);
nand U8993 (N_8993,N_2712,N_1946);
nor U8994 (N_8994,N_3249,N_866);
nor U8995 (N_8995,N_3019,N_4239);
xor U8996 (N_8996,N_2555,N_2589);
or U8997 (N_8997,N_1477,N_375);
nand U8998 (N_8998,N_4072,N_2524);
or U8999 (N_8999,N_822,N_4824);
and U9000 (N_9000,N_2203,N_788);
or U9001 (N_9001,N_4016,N_117);
nor U9002 (N_9002,N_4804,N_277);
and U9003 (N_9003,N_1376,N_4762);
or U9004 (N_9004,N_1843,N_3421);
and U9005 (N_9005,N_2705,N_2100);
xnor U9006 (N_9006,N_2292,N_2089);
or U9007 (N_9007,N_1693,N_4450);
and U9008 (N_9008,N_1084,N_2605);
nand U9009 (N_9009,N_2208,N_1414);
nor U9010 (N_9010,N_491,N_4615);
nand U9011 (N_9011,N_433,N_651);
nand U9012 (N_9012,N_1429,N_1844);
nor U9013 (N_9013,N_1761,N_2305);
or U9014 (N_9014,N_1816,N_123);
or U9015 (N_9015,N_180,N_236);
nor U9016 (N_9016,N_4107,N_4340);
nand U9017 (N_9017,N_71,N_2735);
xnor U9018 (N_9018,N_3184,N_555);
nor U9019 (N_9019,N_4319,N_4375);
nor U9020 (N_9020,N_339,N_180);
nand U9021 (N_9021,N_3364,N_4964);
nand U9022 (N_9022,N_4444,N_4799);
nand U9023 (N_9023,N_4426,N_4190);
and U9024 (N_9024,N_1514,N_1615);
or U9025 (N_9025,N_633,N_2388);
nand U9026 (N_9026,N_461,N_1610);
xor U9027 (N_9027,N_4824,N_714);
and U9028 (N_9028,N_4806,N_1215);
nor U9029 (N_9029,N_618,N_2099);
nor U9030 (N_9030,N_78,N_0);
nor U9031 (N_9031,N_364,N_1955);
and U9032 (N_9032,N_4070,N_2497);
xor U9033 (N_9033,N_1090,N_3351);
xnor U9034 (N_9034,N_1811,N_1121);
nand U9035 (N_9035,N_911,N_4539);
or U9036 (N_9036,N_1840,N_1622);
or U9037 (N_9037,N_3179,N_3671);
nand U9038 (N_9038,N_3876,N_3441);
nand U9039 (N_9039,N_4495,N_1732);
or U9040 (N_9040,N_578,N_790);
or U9041 (N_9041,N_3821,N_3833);
nand U9042 (N_9042,N_4246,N_4881);
or U9043 (N_9043,N_4811,N_1797);
nor U9044 (N_9044,N_1438,N_3003);
and U9045 (N_9045,N_3821,N_4485);
xnor U9046 (N_9046,N_2475,N_823);
or U9047 (N_9047,N_3802,N_1087);
nand U9048 (N_9048,N_3158,N_2150);
or U9049 (N_9049,N_2969,N_105);
nand U9050 (N_9050,N_988,N_674);
nor U9051 (N_9051,N_1778,N_395);
nor U9052 (N_9052,N_2695,N_896);
and U9053 (N_9053,N_1262,N_2552);
and U9054 (N_9054,N_878,N_105);
nand U9055 (N_9055,N_2250,N_4181);
and U9056 (N_9056,N_4001,N_212);
or U9057 (N_9057,N_254,N_411);
and U9058 (N_9058,N_1860,N_4242);
nor U9059 (N_9059,N_1748,N_722);
and U9060 (N_9060,N_4582,N_1611);
and U9061 (N_9061,N_3503,N_3956);
nor U9062 (N_9062,N_4385,N_1994);
nand U9063 (N_9063,N_4053,N_3217);
nand U9064 (N_9064,N_1498,N_614);
and U9065 (N_9065,N_1779,N_4615);
nor U9066 (N_9066,N_3301,N_2823);
nor U9067 (N_9067,N_2485,N_3243);
and U9068 (N_9068,N_2849,N_2056);
or U9069 (N_9069,N_1918,N_3028);
nand U9070 (N_9070,N_4108,N_3578);
and U9071 (N_9071,N_753,N_4502);
or U9072 (N_9072,N_4895,N_154);
nand U9073 (N_9073,N_2475,N_1236);
and U9074 (N_9074,N_867,N_4923);
xor U9075 (N_9075,N_3481,N_235);
nor U9076 (N_9076,N_564,N_4955);
nand U9077 (N_9077,N_4340,N_2285);
nand U9078 (N_9078,N_871,N_1224);
or U9079 (N_9079,N_4782,N_2144);
nor U9080 (N_9080,N_4304,N_2196);
or U9081 (N_9081,N_2211,N_1404);
nor U9082 (N_9082,N_384,N_848);
xnor U9083 (N_9083,N_890,N_4722);
xnor U9084 (N_9084,N_4315,N_4584);
nor U9085 (N_9085,N_1936,N_2078);
or U9086 (N_9086,N_2770,N_1645);
or U9087 (N_9087,N_1223,N_4017);
nor U9088 (N_9088,N_3670,N_4334);
nor U9089 (N_9089,N_258,N_4026);
or U9090 (N_9090,N_3349,N_4690);
xor U9091 (N_9091,N_3263,N_3360);
and U9092 (N_9092,N_3961,N_3093);
and U9093 (N_9093,N_1518,N_1736);
nor U9094 (N_9094,N_1018,N_1422);
nand U9095 (N_9095,N_4475,N_3563);
nand U9096 (N_9096,N_4629,N_1192);
nor U9097 (N_9097,N_2,N_695);
or U9098 (N_9098,N_2999,N_2871);
or U9099 (N_9099,N_2645,N_4112);
nand U9100 (N_9100,N_922,N_1029);
or U9101 (N_9101,N_1483,N_3448);
nand U9102 (N_9102,N_177,N_3025);
xnor U9103 (N_9103,N_2497,N_4897);
or U9104 (N_9104,N_2867,N_3105);
nand U9105 (N_9105,N_4037,N_4526);
and U9106 (N_9106,N_2858,N_1340);
nor U9107 (N_9107,N_1788,N_2716);
xor U9108 (N_9108,N_973,N_4588);
and U9109 (N_9109,N_1172,N_4412);
nand U9110 (N_9110,N_3836,N_4555);
or U9111 (N_9111,N_1989,N_89);
nor U9112 (N_9112,N_132,N_295);
and U9113 (N_9113,N_4979,N_4178);
and U9114 (N_9114,N_4487,N_2126);
or U9115 (N_9115,N_4694,N_4466);
or U9116 (N_9116,N_4258,N_1858);
nor U9117 (N_9117,N_216,N_2077);
xor U9118 (N_9118,N_3300,N_251);
and U9119 (N_9119,N_1346,N_2467);
or U9120 (N_9120,N_2943,N_231);
or U9121 (N_9121,N_3906,N_3475);
or U9122 (N_9122,N_3113,N_4494);
or U9123 (N_9123,N_1442,N_1943);
or U9124 (N_9124,N_3428,N_2620);
nor U9125 (N_9125,N_1359,N_4505);
or U9126 (N_9126,N_2988,N_1421);
nor U9127 (N_9127,N_1865,N_2450);
nor U9128 (N_9128,N_21,N_267);
nand U9129 (N_9129,N_3409,N_151);
and U9130 (N_9130,N_1993,N_1544);
and U9131 (N_9131,N_4558,N_2223);
or U9132 (N_9132,N_2385,N_2236);
nor U9133 (N_9133,N_4454,N_1354);
nor U9134 (N_9134,N_2845,N_490);
nand U9135 (N_9135,N_4072,N_1923);
nand U9136 (N_9136,N_81,N_3979);
nand U9137 (N_9137,N_1136,N_2851);
nor U9138 (N_9138,N_1055,N_3278);
nor U9139 (N_9139,N_647,N_4892);
nor U9140 (N_9140,N_2913,N_4399);
xor U9141 (N_9141,N_3088,N_3950);
nor U9142 (N_9142,N_1135,N_190);
nand U9143 (N_9143,N_1016,N_2565);
and U9144 (N_9144,N_4072,N_105);
nand U9145 (N_9145,N_1078,N_1337);
and U9146 (N_9146,N_2361,N_1775);
or U9147 (N_9147,N_88,N_917);
nor U9148 (N_9148,N_4137,N_167);
nor U9149 (N_9149,N_4279,N_2258);
nand U9150 (N_9150,N_4446,N_1991);
nor U9151 (N_9151,N_2659,N_1616);
nor U9152 (N_9152,N_2724,N_2102);
and U9153 (N_9153,N_53,N_1708);
nor U9154 (N_9154,N_1457,N_3271);
nand U9155 (N_9155,N_651,N_2645);
and U9156 (N_9156,N_2528,N_461);
nand U9157 (N_9157,N_1653,N_1777);
and U9158 (N_9158,N_470,N_709);
nand U9159 (N_9159,N_4422,N_373);
nor U9160 (N_9160,N_2151,N_1620);
or U9161 (N_9161,N_1546,N_346);
nor U9162 (N_9162,N_187,N_144);
xor U9163 (N_9163,N_4024,N_4520);
nand U9164 (N_9164,N_3480,N_1983);
nand U9165 (N_9165,N_3257,N_3053);
and U9166 (N_9166,N_1322,N_1368);
or U9167 (N_9167,N_2671,N_2281);
nor U9168 (N_9168,N_3683,N_1839);
or U9169 (N_9169,N_2913,N_2474);
and U9170 (N_9170,N_259,N_2398);
nand U9171 (N_9171,N_2798,N_769);
and U9172 (N_9172,N_4709,N_4788);
nor U9173 (N_9173,N_1596,N_2622);
nand U9174 (N_9174,N_240,N_1351);
nor U9175 (N_9175,N_4137,N_2495);
or U9176 (N_9176,N_3778,N_2603);
or U9177 (N_9177,N_719,N_3253);
or U9178 (N_9178,N_2230,N_1084);
or U9179 (N_9179,N_4644,N_1364);
xnor U9180 (N_9180,N_4014,N_2838);
nor U9181 (N_9181,N_2572,N_1092);
nor U9182 (N_9182,N_3919,N_2209);
and U9183 (N_9183,N_3099,N_1384);
nand U9184 (N_9184,N_1051,N_3025);
xor U9185 (N_9185,N_4077,N_4158);
nand U9186 (N_9186,N_1616,N_3365);
and U9187 (N_9187,N_4870,N_1415);
or U9188 (N_9188,N_2721,N_173);
nor U9189 (N_9189,N_255,N_1918);
nand U9190 (N_9190,N_79,N_3576);
nand U9191 (N_9191,N_4488,N_105);
nor U9192 (N_9192,N_3125,N_533);
nand U9193 (N_9193,N_740,N_2281);
nand U9194 (N_9194,N_2974,N_2319);
or U9195 (N_9195,N_1490,N_1769);
nand U9196 (N_9196,N_1654,N_2885);
nor U9197 (N_9197,N_1103,N_1394);
xnor U9198 (N_9198,N_838,N_4886);
nand U9199 (N_9199,N_8,N_2414);
nand U9200 (N_9200,N_854,N_3083);
xor U9201 (N_9201,N_566,N_2700);
nand U9202 (N_9202,N_4025,N_1100);
or U9203 (N_9203,N_858,N_908);
nand U9204 (N_9204,N_3092,N_3165);
nand U9205 (N_9205,N_148,N_550);
or U9206 (N_9206,N_4457,N_2178);
and U9207 (N_9207,N_1815,N_4516);
or U9208 (N_9208,N_2688,N_3380);
nand U9209 (N_9209,N_2516,N_299);
and U9210 (N_9210,N_2632,N_362);
xnor U9211 (N_9211,N_959,N_4262);
and U9212 (N_9212,N_3055,N_1709);
xnor U9213 (N_9213,N_3844,N_1919);
nand U9214 (N_9214,N_3822,N_4248);
nor U9215 (N_9215,N_3933,N_1591);
nor U9216 (N_9216,N_3112,N_3470);
nand U9217 (N_9217,N_3,N_2580);
nand U9218 (N_9218,N_2530,N_4074);
nor U9219 (N_9219,N_616,N_692);
and U9220 (N_9220,N_1688,N_1503);
or U9221 (N_9221,N_3114,N_4369);
or U9222 (N_9222,N_4330,N_2542);
and U9223 (N_9223,N_593,N_181);
and U9224 (N_9224,N_1319,N_115);
nor U9225 (N_9225,N_3024,N_2340);
xnor U9226 (N_9226,N_3961,N_1999);
and U9227 (N_9227,N_3662,N_1267);
xor U9228 (N_9228,N_4525,N_346);
nand U9229 (N_9229,N_910,N_1778);
and U9230 (N_9230,N_1932,N_182);
and U9231 (N_9231,N_3712,N_1343);
nor U9232 (N_9232,N_718,N_3358);
and U9233 (N_9233,N_861,N_2604);
xnor U9234 (N_9234,N_2514,N_1841);
and U9235 (N_9235,N_1960,N_2706);
or U9236 (N_9236,N_4702,N_3731);
nor U9237 (N_9237,N_2464,N_1488);
nand U9238 (N_9238,N_4697,N_3506);
and U9239 (N_9239,N_104,N_4067);
and U9240 (N_9240,N_4138,N_1521);
and U9241 (N_9241,N_3979,N_3714);
nand U9242 (N_9242,N_2313,N_2540);
or U9243 (N_9243,N_1422,N_3310);
and U9244 (N_9244,N_4946,N_1166);
or U9245 (N_9245,N_505,N_1884);
nor U9246 (N_9246,N_215,N_4909);
or U9247 (N_9247,N_3448,N_1081);
and U9248 (N_9248,N_1852,N_25);
nor U9249 (N_9249,N_2278,N_4058);
xnor U9250 (N_9250,N_2950,N_986);
and U9251 (N_9251,N_3468,N_4572);
or U9252 (N_9252,N_3937,N_4890);
nor U9253 (N_9253,N_1000,N_3651);
and U9254 (N_9254,N_1586,N_3908);
and U9255 (N_9255,N_3149,N_4239);
and U9256 (N_9256,N_3075,N_3357);
and U9257 (N_9257,N_253,N_4645);
nor U9258 (N_9258,N_4129,N_3906);
or U9259 (N_9259,N_1250,N_656);
nand U9260 (N_9260,N_2979,N_2069);
nand U9261 (N_9261,N_3677,N_183);
nor U9262 (N_9262,N_2108,N_353);
and U9263 (N_9263,N_3154,N_2410);
or U9264 (N_9264,N_4099,N_426);
nand U9265 (N_9265,N_903,N_1880);
nand U9266 (N_9266,N_3276,N_2232);
or U9267 (N_9267,N_3504,N_3294);
nand U9268 (N_9268,N_1239,N_3234);
nor U9269 (N_9269,N_3933,N_3315);
and U9270 (N_9270,N_1470,N_3054);
or U9271 (N_9271,N_3331,N_4003);
xor U9272 (N_9272,N_2116,N_2957);
nand U9273 (N_9273,N_388,N_2710);
nand U9274 (N_9274,N_2195,N_3471);
nor U9275 (N_9275,N_876,N_2074);
nor U9276 (N_9276,N_1296,N_2948);
nand U9277 (N_9277,N_4202,N_3568);
and U9278 (N_9278,N_2412,N_3474);
nand U9279 (N_9279,N_4636,N_4262);
nor U9280 (N_9280,N_887,N_2712);
nor U9281 (N_9281,N_3940,N_553);
nor U9282 (N_9282,N_2557,N_2788);
xor U9283 (N_9283,N_4767,N_3487);
and U9284 (N_9284,N_2539,N_284);
nor U9285 (N_9285,N_2971,N_1090);
xnor U9286 (N_9286,N_992,N_2823);
nor U9287 (N_9287,N_2010,N_4166);
nor U9288 (N_9288,N_150,N_3173);
or U9289 (N_9289,N_3328,N_1586);
nand U9290 (N_9290,N_3511,N_4293);
and U9291 (N_9291,N_1793,N_2808);
xnor U9292 (N_9292,N_1473,N_2378);
nand U9293 (N_9293,N_2870,N_3488);
or U9294 (N_9294,N_4483,N_3849);
or U9295 (N_9295,N_1279,N_2661);
xor U9296 (N_9296,N_1216,N_2853);
nor U9297 (N_9297,N_2500,N_3854);
and U9298 (N_9298,N_3193,N_939);
nor U9299 (N_9299,N_3158,N_1943);
nor U9300 (N_9300,N_2248,N_2465);
and U9301 (N_9301,N_1077,N_4698);
and U9302 (N_9302,N_38,N_3331);
nor U9303 (N_9303,N_3465,N_4661);
xnor U9304 (N_9304,N_3624,N_125);
and U9305 (N_9305,N_3872,N_141);
nor U9306 (N_9306,N_3008,N_2237);
nor U9307 (N_9307,N_4425,N_1165);
nor U9308 (N_9308,N_4970,N_4852);
nor U9309 (N_9309,N_4094,N_2235);
or U9310 (N_9310,N_3017,N_1365);
nand U9311 (N_9311,N_3916,N_1333);
and U9312 (N_9312,N_4837,N_275);
nor U9313 (N_9313,N_4888,N_144);
or U9314 (N_9314,N_74,N_2828);
or U9315 (N_9315,N_2480,N_4165);
nand U9316 (N_9316,N_1209,N_3910);
and U9317 (N_9317,N_2002,N_3876);
nor U9318 (N_9318,N_982,N_3654);
nor U9319 (N_9319,N_3737,N_3548);
xor U9320 (N_9320,N_1022,N_581);
and U9321 (N_9321,N_4499,N_595);
nor U9322 (N_9322,N_2124,N_3386);
xor U9323 (N_9323,N_4573,N_2196);
nand U9324 (N_9324,N_1627,N_1341);
nor U9325 (N_9325,N_1654,N_4581);
or U9326 (N_9326,N_347,N_3527);
or U9327 (N_9327,N_3617,N_30);
nand U9328 (N_9328,N_1162,N_4622);
and U9329 (N_9329,N_3664,N_1751);
or U9330 (N_9330,N_4853,N_3036);
nand U9331 (N_9331,N_555,N_3409);
xnor U9332 (N_9332,N_2216,N_132);
xnor U9333 (N_9333,N_2040,N_3847);
nand U9334 (N_9334,N_790,N_663);
or U9335 (N_9335,N_2539,N_3172);
and U9336 (N_9336,N_2481,N_2763);
and U9337 (N_9337,N_3592,N_2886);
nand U9338 (N_9338,N_1931,N_3953);
nor U9339 (N_9339,N_1570,N_1304);
nor U9340 (N_9340,N_1090,N_1587);
and U9341 (N_9341,N_4287,N_4125);
or U9342 (N_9342,N_1854,N_396);
and U9343 (N_9343,N_1185,N_2431);
and U9344 (N_9344,N_2031,N_2900);
nor U9345 (N_9345,N_2088,N_79);
and U9346 (N_9346,N_4930,N_267);
and U9347 (N_9347,N_4056,N_2204);
or U9348 (N_9348,N_4319,N_2574);
nor U9349 (N_9349,N_3577,N_2587);
xnor U9350 (N_9350,N_4182,N_1780);
or U9351 (N_9351,N_2341,N_4317);
and U9352 (N_9352,N_4351,N_4543);
nor U9353 (N_9353,N_3600,N_85);
xnor U9354 (N_9354,N_3719,N_2782);
or U9355 (N_9355,N_3420,N_1897);
nor U9356 (N_9356,N_4523,N_1331);
nand U9357 (N_9357,N_4395,N_1787);
or U9358 (N_9358,N_3135,N_800);
nor U9359 (N_9359,N_2734,N_4022);
xor U9360 (N_9360,N_4646,N_2246);
nor U9361 (N_9361,N_4016,N_4575);
and U9362 (N_9362,N_3295,N_2886);
xor U9363 (N_9363,N_3449,N_1148);
nor U9364 (N_9364,N_2600,N_2117);
nor U9365 (N_9365,N_1674,N_2357);
or U9366 (N_9366,N_3110,N_3305);
nor U9367 (N_9367,N_1161,N_1511);
or U9368 (N_9368,N_2930,N_4603);
and U9369 (N_9369,N_2468,N_4652);
nand U9370 (N_9370,N_990,N_314);
xor U9371 (N_9371,N_560,N_3840);
nor U9372 (N_9372,N_2960,N_159);
nand U9373 (N_9373,N_4738,N_2268);
nand U9374 (N_9374,N_520,N_4395);
or U9375 (N_9375,N_4814,N_2334);
xor U9376 (N_9376,N_857,N_4047);
and U9377 (N_9377,N_2304,N_591);
nand U9378 (N_9378,N_1418,N_3265);
nor U9379 (N_9379,N_3945,N_2585);
or U9380 (N_9380,N_2262,N_1468);
or U9381 (N_9381,N_3672,N_3739);
or U9382 (N_9382,N_2099,N_4788);
nand U9383 (N_9383,N_805,N_255);
or U9384 (N_9384,N_2381,N_500);
nand U9385 (N_9385,N_77,N_1609);
and U9386 (N_9386,N_3120,N_2120);
nand U9387 (N_9387,N_3948,N_258);
nor U9388 (N_9388,N_3730,N_4233);
xnor U9389 (N_9389,N_4757,N_2785);
nand U9390 (N_9390,N_1602,N_4327);
nand U9391 (N_9391,N_2832,N_4597);
or U9392 (N_9392,N_2405,N_1307);
nand U9393 (N_9393,N_1513,N_4555);
and U9394 (N_9394,N_3039,N_3991);
nand U9395 (N_9395,N_1776,N_3261);
nor U9396 (N_9396,N_1542,N_4446);
nor U9397 (N_9397,N_3661,N_1893);
and U9398 (N_9398,N_2823,N_1030);
nor U9399 (N_9399,N_86,N_3910);
or U9400 (N_9400,N_424,N_2412);
xnor U9401 (N_9401,N_1487,N_3703);
nand U9402 (N_9402,N_4237,N_3724);
or U9403 (N_9403,N_4897,N_3092);
xor U9404 (N_9404,N_537,N_3292);
nand U9405 (N_9405,N_1888,N_1464);
and U9406 (N_9406,N_3670,N_398);
xor U9407 (N_9407,N_807,N_275);
or U9408 (N_9408,N_494,N_509);
xnor U9409 (N_9409,N_3044,N_2260);
nor U9410 (N_9410,N_1615,N_464);
and U9411 (N_9411,N_3979,N_4612);
or U9412 (N_9412,N_4424,N_4079);
and U9413 (N_9413,N_534,N_4719);
nor U9414 (N_9414,N_437,N_3723);
nor U9415 (N_9415,N_3866,N_3679);
nor U9416 (N_9416,N_3122,N_3442);
and U9417 (N_9417,N_1798,N_1144);
nor U9418 (N_9418,N_3816,N_3923);
and U9419 (N_9419,N_2422,N_2665);
xnor U9420 (N_9420,N_450,N_2630);
and U9421 (N_9421,N_2803,N_1678);
and U9422 (N_9422,N_1879,N_2803);
and U9423 (N_9423,N_1906,N_2653);
xnor U9424 (N_9424,N_3399,N_2642);
or U9425 (N_9425,N_4402,N_4118);
xnor U9426 (N_9426,N_598,N_512);
xnor U9427 (N_9427,N_788,N_2194);
nor U9428 (N_9428,N_1672,N_3717);
and U9429 (N_9429,N_1034,N_2384);
xnor U9430 (N_9430,N_3343,N_134);
nand U9431 (N_9431,N_3712,N_4204);
nor U9432 (N_9432,N_1978,N_685);
and U9433 (N_9433,N_796,N_4833);
xnor U9434 (N_9434,N_4815,N_4993);
nor U9435 (N_9435,N_1786,N_2069);
or U9436 (N_9436,N_300,N_1644);
or U9437 (N_9437,N_504,N_2958);
nand U9438 (N_9438,N_304,N_3010);
nor U9439 (N_9439,N_2400,N_3751);
nor U9440 (N_9440,N_1579,N_2405);
and U9441 (N_9441,N_2451,N_0);
or U9442 (N_9442,N_3885,N_3345);
or U9443 (N_9443,N_492,N_3830);
nor U9444 (N_9444,N_2867,N_2176);
xor U9445 (N_9445,N_3940,N_4684);
or U9446 (N_9446,N_127,N_1357);
nor U9447 (N_9447,N_509,N_3276);
nor U9448 (N_9448,N_567,N_1431);
nor U9449 (N_9449,N_2832,N_2199);
nand U9450 (N_9450,N_3199,N_3910);
nor U9451 (N_9451,N_1022,N_162);
xor U9452 (N_9452,N_3969,N_1661);
or U9453 (N_9453,N_55,N_4227);
nor U9454 (N_9454,N_4006,N_4979);
or U9455 (N_9455,N_156,N_464);
or U9456 (N_9456,N_897,N_4752);
or U9457 (N_9457,N_2281,N_2662);
nor U9458 (N_9458,N_2261,N_2833);
or U9459 (N_9459,N_2752,N_953);
or U9460 (N_9460,N_3248,N_2999);
nor U9461 (N_9461,N_4445,N_1308);
and U9462 (N_9462,N_1957,N_1161);
nand U9463 (N_9463,N_3184,N_3188);
nand U9464 (N_9464,N_512,N_590);
nor U9465 (N_9465,N_2216,N_4219);
nand U9466 (N_9466,N_2330,N_2337);
and U9467 (N_9467,N_2631,N_1269);
nand U9468 (N_9468,N_340,N_2196);
or U9469 (N_9469,N_2283,N_392);
nand U9470 (N_9470,N_794,N_1659);
nor U9471 (N_9471,N_3175,N_8);
xnor U9472 (N_9472,N_2152,N_3455);
nor U9473 (N_9473,N_940,N_2018);
or U9474 (N_9474,N_888,N_1395);
and U9475 (N_9475,N_3801,N_4181);
nand U9476 (N_9476,N_3037,N_762);
nor U9477 (N_9477,N_2441,N_30);
and U9478 (N_9478,N_946,N_2662);
and U9479 (N_9479,N_2869,N_3673);
nand U9480 (N_9480,N_3302,N_3882);
nand U9481 (N_9481,N_381,N_3031);
nor U9482 (N_9482,N_4718,N_154);
xor U9483 (N_9483,N_4090,N_2377);
and U9484 (N_9484,N_3043,N_4190);
or U9485 (N_9485,N_551,N_4292);
nand U9486 (N_9486,N_4714,N_965);
nand U9487 (N_9487,N_3614,N_1945);
nor U9488 (N_9488,N_1665,N_281);
nor U9489 (N_9489,N_4455,N_3601);
nor U9490 (N_9490,N_4675,N_602);
and U9491 (N_9491,N_2946,N_2506);
nor U9492 (N_9492,N_831,N_4971);
nor U9493 (N_9493,N_2595,N_1113);
xor U9494 (N_9494,N_2576,N_372);
nand U9495 (N_9495,N_4502,N_4878);
or U9496 (N_9496,N_4972,N_1673);
and U9497 (N_9497,N_1806,N_288);
or U9498 (N_9498,N_3886,N_4097);
nor U9499 (N_9499,N_89,N_4004);
and U9500 (N_9500,N_3145,N_3619);
and U9501 (N_9501,N_3123,N_2247);
or U9502 (N_9502,N_287,N_3419);
xor U9503 (N_9503,N_965,N_4324);
or U9504 (N_9504,N_2653,N_1615);
or U9505 (N_9505,N_2822,N_2110);
and U9506 (N_9506,N_833,N_3137);
or U9507 (N_9507,N_522,N_4358);
or U9508 (N_9508,N_2596,N_3477);
and U9509 (N_9509,N_3490,N_2402);
nor U9510 (N_9510,N_361,N_3867);
nand U9511 (N_9511,N_1252,N_263);
nand U9512 (N_9512,N_473,N_4289);
nor U9513 (N_9513,N_4313,N_3716);
nor U9514 (N_9514,N_307,N_2499);
nor U9515 (N_9515,N_4775,N_2707);
and U9516 (N_9516,N_1726,N_1851);
xor U9517 (N_9517,N_3966,N_209);
nand U9518 (N_9518,N_1580,N_3636);
nand U9519 (N_9519,N_2256,N_4561);
and U9520 (N_9520,N_2112,N_816);
nand U9521 (N_9521,N_4761,N_704);
nor U9522 (N_9522,N_309,N_4903);
and U9523 (N_9523,N_4459,N_2178);
nor U9524 (N_9524,N_1367,N_655);
nor U9525 (N_9525,N_2215,N_1382);
nor U9526 (N_9526,N_2326,N_4580);
and U9527 (N_9527,N_263,N_1793);
nand U9528 (N_9528,N_2549,N_2366);
xnor U9529 (N_9529,N_3895,N_4005);
nand U9530 (N_9530,N_4788,N_317);
and U9531 (N_9531,N_3743,N_221);
nor U9532 (N_9532,N_3578,N_103);
nand U9533 (N_9533,N_2697,N_4449);
xor U9534 (N_9534,N_2804,N_895);
nor U9535 (N_9535,N_3245,N_1233);
or U9536 (N_9536,N_3384,N_3532);
and U9537 (N_9537,N_4284,N_105);
nor U9538 (N_9538,N_3969,N_2284);
or U9539 (N_9539,N_4931,N_2125);
nor U9540 (N_9540,N_2181,N_2915);
nor U9541 (N_9541,N_4820,N_3460);
and U9542 (N_9542,N_3668,N_977);
and U9543 (N_9543,N_4913,N_1673);
nand U9544 (N_9544,N_2611,N_2718);
or U9545 (N_9545,N_3631,N_1871);
xnor U9546 (N_9546,N_3667,N_379);
xnor U9547 (N_9547,N_4567,N_2446);
nor U9548 (N_9548,N_3287,N_2989);
nor U9549 (N_9549,N_2169,N_3235);
or U9550 (N_9550,N_3279,N_2691);
and U9551 (N_9551,N_605,N_2534);
or U9552 (N_9552,N_77,N_574);
or U9553 (N_9553,N_3973,N_2045);
nor U9554 (N_9554,N_2919,N_4549);
nor U9555 (N_9555,N_2053,N_4300);
nand U9556 (N_9556,N_147,N_4775);
and U9557 (N_9557,N_1814,N_4041);
xor U9558 (N_9558,N_2927,N_1114);
nor U9559 (N_9559,N_2813,N_1067);
and U9560 (N_9560,N_3925,N_3745);
nand U9561 (N_9561,N_2608,N_4604);
nor U9562 (N_9562,N_2420,N_2862);
and U9563 (N_9563,N_18,N_3384);
xor U9564 (N_9564,N_1959,N_2809);
or U9565 (N_9565,N_138,N_1777);
nand U9566 (N_9566,N_1323,N_4180);
or U9567 (N_9567,N_4584,N_1018);
or U9568 (N_9568,N_1405,N_2879);
nand U9569 (N_9569,N_699,N_1787);
and U9570 (N_9570,N_1795,N_2103);
and U9571 (N_9571,N_3126,N_3542);
nor U9572 (N_9572,N_595,N_389);
or U9573 (N_9573,N_4931,N_4918);
or U9574 (N_9574,N_4559,N_437);
or U9575 (N_9575,N_1770,N_3032);
xnor U9576 (N_9576,N_1639,N_2834);
nor U9577 (N_9577,N_63,N_2800);
nand U9578 (N_9578,N_2100,N_2750);
nand U9579 (N_9579,N_4318,N_389);
or U9580 (N_9580,N_2415,N_4507);
nand U9581 (N_9581,N_4494,N_1183);
xnor U9582 (N_9582,N_1819,N_3946);
nand U9583 (N_9583,N_2746,N_4955);
nor U9584 (N_9584,N_1126,N_880);
or U9585 (N_9585,N_917,N_1470);
nor U9586 (N_9586,N_4079,N_3499);
nand U9587 (N_9587,N_4395,N_792);
nand U9588 (N_9588,N_4553,N_1646);
and U9589 (N_9589,N_4122,N_2162);
nand U9590 (N_9590,N_1556,N_2198);
xnor U9591 (N_9591,N_1001,N_2317);
or U9592 (N_9592,N_425,N_3609);
and U9593 (N_9593,N_175,N_2069);
xnor U9594 (N_9594,N_4397,N_2289);
xor U9595 (N_9595,N_4217,N_3337);
xnor U9596 (N_9596,N_4204,N_680);
or U9597 (N_9597,N_1927,N_2061);
and U9598 (N_9598,N_3800,N_932);
or U9599 (N_9599,N_844,N_894);
nor U9600 (N_9600,N_2915,N_945);
nand U9601 (N_9601,N_847,N_4729);
and U9602 (N_9602,N_1465,N_4792);
and U9603 (N_9603,N_2064,N_857);
nor U9604 (N_9604,N_2737,N_4592);
and U9605 (N_9605,N_2553,N_661);
or U9606 (N_9606,N_646,N_4407);
nand U9607 (N_9607,N_1137,N_2301);
or U9608 (N_9608,N_2017,N_362);
and U9609 (N_9609,N_1411,N_4900);
or U9610 (N_9610,N_2369,N_1083);
xnor U9611 (N_9611,N_2922,N_2866);
xor U9612 (N_9612,N_1921,N_4846);
and U9613 (N_9613,N_4468,N_4687);
or U9614 (N_9614,N_184,N_2374);
nor U9615 (N_9615,N_1777,N_4949);
nand U9616 (N_9616,N_432,N_1009);
nor U9617 (N_9617,N_2823,N_1861);
or U9618 (N_9618,N_790,N_1863);
nor U9619 (N_9619,N_4601,N_3755);
or U9620 (N_9620,N_3144,N_3088);
or U9621 (N_9621,N_2411,N_4819);
xnor U9622 (N_9622,N_2048,N_2473);
or U9623 (N_9623,N_2178,N_3395);
nand U9624 (N_9624,N_2424,N_1722);
or U9625 (N_9625,N_49,N_4289);
or U9626 (N_9626,N_3588,N_3672);
and U9627 (N_9627,N_4727,N_408);
nand U9628 (N_9628,N_1678,N_598);
or U9629 (N_9629,N_3565,N_2205);
nand U9630 (N_9630,N_85,N_1753);
or U9631 (N_9631,N_3343,N_1394);
or U9632 (N_9632,N_296,N_319);
and U9633 (N_9633,N_4941,N_1999);
nor U9634 (N_9634,N_4595,N_869);
or U9635 (N_9635,N_3132,N_1549);
nor U9636 (N_9636,N_4696,N_1080);
nand U9637 (N_9637,N_2450,N_2310);
and U9638 (N_9638,N_725,N_3261);
nor U9639 (N_9639,N_4739,N_518);
nand U9640 (N_9640,N_3639,N_1775);
and U9641 (N_9641,N_4038,N_2802);
and U9642 (N_9642,N_1545,N_1523);
nor U9643 (N_9643,N_325,N_2744);
nand U9644 (N_9644,N_568,N_4722);
or U9645 (N_9645,N_4029,N_2047);
nand U9646 (N_9646,N_4399,N_62);
or U9647 (N_9647,N_1277,N_3025);
nor U9648 (N_9648,N_4538,N_608);
nand U9649 (N_9649,N_665,N_4099);
nor U9650 (N_9650,N_99,N_3405);
or U9651 (N_9651,N_9,N_3341);
or U9652 (N_9652,N_3321,N_1870);
nor U9653 (N_9653,N_417,N_475);
nor U9654 (N_9654,N_3377,N_3767);
nor U9655 (N_9655,N_1092,N_2768);
nor U9656 (N_9656,N_4567,N_1773);
or U9657 (N_9657,N_4309,N_1885);
nor U9658 (N_9658,N_1664,N_4128);
nor U9659 (N_9659,N_2886,N_407);
or U9660 (N_9660,N_3474,N_2071);
xnor U9661 (N_9661,N_2151,N_3311);
or U9662 (N_9662,N_3672,N_877);
nand U9663 (N_9663,N_3981,N_3855);
nand U9664 (N_9664,N_2559,N_2432);
nand U9665 (N_9665,N_2379,N_57);
nand U9666 (N_9666,N_1204,N_4266);
or U9667 (N_9667,N_3212,N_4921);
and U9668 (N_9668,N_4413,N_1246);
and U9669 (N_9669,N_4160,N_281);
and U9670 (N_9670,N_4694,N_2368);
nand U9671 (N_9671,N_2003,N_2740);
nand U9672 (N_9672,N_3652,N_864);
nand U9673 (N_9673,N_1426,N_3890);
nand U9674 (N_9674,N_94,N_4066);
nor U9675 (N_9675,N_1156,N_1842);
nand U9676 (N_9676,N_4888,N_3861);
and U9677 (N_9677,N_4831,N_401);
nor U9678 (N_9678,N_3892,N_1467);
or U9679 (N_9679,N_48,N_3230);
and U9680 (N_9680,N_4261,N_2786);
or U9681 (N_9681,N_4353,N_1255);
nand U9682 (N_9682,N_4396,N_3519);
nor U9683 (N_9683,N_3327,N_980);
nand U9684 (N_9684,N_3419,N_1592);
nor U9685 (N_9685,N_2311,N_3695);
nand U9686 (N_9686,N_601,N_4905);
xor U9687 (N_9687,N_1956,N_3465);
nand U9688 (N_9688,N_742,N_1539);
nor U9689 (N_9689,N_1947,N_4644);
nor U9690 (N_9690,N_1716,N_1509);
nor U9691 (N_9691,N_2783,N_4653);
or U9692 (N_9692,N_2055,N_3699);
nor U9693 (N_9693,N_2390,N_3643);
nor U9694 (N_9694,N_1940,N_2867);
and U9695 (N_9695,N_1725,N_2382);
nand U9696 (N_9696,N_2277,N_3284);
and U9697 (N_9697,N_3516,N_2858);
or U9698 (N_9698,N_4282,N_587);
nand U9699 (N_9699,N_4583,N_4885);
and U9700 (N_9700,N_4146,N_1131);
nand U9701 (N_9701,N_3532,N_2741);
xor U9702 (N_9702,N_1552,N_3742);
xnor U9703 (N_9703,N_3714,N_1727);
nor U9704 (N_9704,N_3870,N_594);
nor U9705 (N_9705,N_3266,N_3531);
or U9706 (N_9706,N_4676,N_3212);
nand U9707 (N_9707,N_1724,N_4421);
and U9708 (N_9708,N_1030,N_4);
nor U9709 (N_9709,N_2503,N_71);
xnor U9710 (N_9710,N_1756,N_2281);
nand U9711 (N_9711,N_1254,N_732);
nor U9712 (N_9712,N_1335,N_911);
xnor U9713 (N_9713,N_2709,N_2930);
nand U9714 (N_9714,N_2303,N_3700);
and U9715 (N_9715,N_3673,N_2493);
nor U9716 (N_9716,N_2067,N_2293);
nor U9717 (N_9717,N_4548,N_3314);
nand U9718 (N_9718,N_1366,N_3129);
xor U9719 (N_9719,N_1008,N_3151);
xor U9720 (N_9720,N_2365,N_257);
nand U9721 (N_9721,N_4468,N_4760);
and U9722 (N_9722,N_3942,N_1285);
and U9723 (N_9723,N_437,N_2225);
nor U9724 (N_9724,N_1314,N_4877);
or U9725 (N_9725,N_172,N_641);
or U9726 (N_9726,N_1092,N_2630);
nand U9727 (N_9727,N_2480,N_3002);
or U9728 (N_9728,N_1414,N_3681);
and U9729 (N_9729,N_2558,N_1529);
nor U9730 (N_9730,N_3223,N_4901);
nand U9731 (N_9731,N_557,N_2939);
and U9732 (N_9732,N_241,N_1892);
nor U9733 (N_9733,N_22,N_3912);
and U9734 (N_9734,N_4005,N_712);
and U9735 (N_9735,N_178,N_1771);
or U9736 (N_9736,N_543,N_1788);
nand U9737 (N_9737,N_1746,N_4414);
nand U9738 (N_9738,N_1232,N_2454);
nor U9739 (N_9739,N_4646,N_3950);
nand U9740 (N_9740,N_800,N_868);
xor U9741 (N_9741,N_16,N_1809);
nor U9742 (N_9742,N_4218,N_3623);
nand U9743 (N_9743,N_4323,N_3235);
nand U9744 (N_9744,N_3147,N_2992);
or U9745 (N_9745,N_3583,N_709);
or U9746 (N_9746,N_4482,N_60);
or U9747 (N_9747,N_3723,N_84);
xor U9748 (N_9748,N_1909,N_1598);
or U9749 (N_9749,N_870,N_772);
nor U9750 (N_9750,N_2410,N_1197);
and U9751 (N_9751,N_4158,N_3648);
or U9752 (N_9752,N_3989,N_2613);
or U9753 (N_9753,N_1938,N_3722);
nand U9754 (N_9754,N_2322,N_1779);
nor U9755 (N_9755,N_2277,N_1152);
nor U9756 (N_9756,N_4682,N_4705);
nand U9757 (N_9757,N_2932,N_2835);
or U9758 (N_9758,N_2881,N_2886);
or U9759 (N_9759,N_1125,N_4356);
or U9760 (N_9760,N_2925,N_4344);
nor U9761 (N_9761,N_2724,N_1371);
and U9762 (N_9762,N_1590,N_4476);
and U9763 (N_9763,N_4287,N_4565);
xor U9764 (N_9764,N_3673,N_471);
nand U9765 (N_9765,N_4802,N_3817);
nor U9766 (N_9766,N_4608,N_553);
or U9767 (N_9767,N_1544,N_2558);
nor U9768 (N_9768,N_4233,N_2465);
nand U9769 (N_9769,N_1973,N_796);
or U9770 (N_9770,N_680,N_983);
or U9771 (N_9771,N_2473,N_1585);
nor U9772 (N_9772,N_315,N_2880);
nand U9773 (N_9773,N_3038,N_976);
or U9774 (N_9774,N_2872,N_2649);
nand U9775 (N_9775,N_1128,N_1078);
nor U9776 (N_9776,N_3602,N_3153);
nor U9777 (N_9777,N_4566,N_1814);
nand U9778 (N_9778,N_2987,N_1815);
nand U9779 (N_9779,N_3372,N_3652);
and U9780 (N_9780,N_2427,N_3260);
nor U9781 (N_9781,N_2702,N_3877);
or U9782 (N_9782,N_2419,N_348);
xnor U9783 (N_9783,N_1378,N_3855);
and U9784 (N_9784,N_2590,N_2610);
or U9785 (N_9785,N_2394,N_994);
nor U9786 (N_9786,N_2153,N_1011);
or U9787 (N_9787,N_1688,N_2844);
nand U9788 (N_9788,N_967,N_991);
and U9789 (N_9789,N_972,N_1979);
xor U9790 (N_9790,N_4922,N_311);
or U9791 (N_9791,N_3056,N_312);
or U9792 (N_9792,N_1380,N_1845);
and U9793 (N_9793,N_2317,N_1714);
xor U9794 (N_9794,N_2838,N_2107);
xnor U9795 (N_9795,N_4013,N_2734);
nor U9796 (N_9796,N_1826,N_2375);
nand U9797 (N_9797,N_4196,N_3143);
nor U9798 (N_9798,N_2292,N_1624);
and U9799 (N_9799,N_2404,N_3303);
nand U9800 (N_9800,N_4518,N_4807);
xnor U9801 (N_9801,N_4933,N_341);
nor U9802 (N_9802,N_3693,N_404);
nand U9803 (N_9803,N_2200,N_4949);
nor U9804 (N_9804,N_3736,N_4234);
nand U9805 (N_9805,N_4474,N_2232);
nand U9806 (N_9806,N_3856,N_1590);
nor U9807 (N_9807,N_3164,N_3271);
or U9808 (N_9808,N_175,N_1456);
or U9809 (N_9809,N_2474,N_4549);
nand U9810 (N_9810,N_2944,N_4655);
nor U9811 (N_9811,N_1548,N_859);
xnor U9812 (N_9812,N_3081,N_4267);
and U9813 (N_9813,N_3836,N_3786);
nand U9814 (N_9814,N_4404,N_3425);
nand U9815 (N_9815,N_4387,N_3700);
xnor U9816 (N_9816,N_4970,N_429);
nor U9817 (N_9817,N_653,N_3708);
and U9818 (N_9818,N_3807,N_882);
and U9819 (N_9819,N_2812,N_1198);
and U9820 (N_9820,N_1766,N_4313);
xor U9821 (N_9821,N_3889,N_783);
and U9822 (N_9822,N_2997,N_199);
nand U9823 (N_9823,N_600,N_1048);
nor U9824 (N_9824,N_1962,N_1612);
nor U9825 (N_9825,N_2190,N_2020);
and U9826 (N_9826,N_3949,N_2838);
nand U9827 (N_9827,N_2208,N_854);
or U9828 (N_9828,N_683,N_4834);
nand U9829 (N_9829,N_45,N_3847);
and U9830 (N_9830,N_4214,N_2496);
xnor U9831 (N_9831,N_3618,N_1023);
nor U9832 (N_9832,N_4439,N_2851);
nor U9833 (N_9833,N_443,N_3189);
nand U9834 (N_9834,N_2167,N_666);
nor U9835 (N_9835,N_4576,N_2610);
and U9836 (N_9836,N_4565,N_1972);
or U9837 (N_9837,N_1625,N_1827);
and U9838 (N_9838,N_2761,N_2876);
nor U9839 (N_9839,N_2746,N_3189);
or U9840 (N_9840,N_641,N_4151);
and U9841 (N_9841,N_2546,N_1384);
and U9842 (N_9842,N_2928,N_4565);
nor U9843 (N_9843,N_3135,N_4694);
nand U9844 (N_9844,N_2768,N_2204);
nor U9845 (N_9845,N_3885,N_2778);
nor U9846 (N_9846,N_4299,N_921);
and U9847 (N_9847,N_2506,N_1899);
xor U9848 (N_9848,N_418,N_647);
and U9849 (N_9849,N_3958,N_472);
or U9850 (N_9850,N_1590,N_1385);
nor U9851 (N_9851,N_4713,N_2063);
or U9852 (N_9852,N_4004,N_3114);
xnor U9853 (N_9853,N_1755,N_1607);
or U9854 (N_9854,N_338,N_1478);
and U9855 (N_9855,N_1078,N_3679);
nand U9856 (N_9856,N_4290,N_3575);
nand U9857 (N_9857,N_2074,N_4226);
and U9858 (N_9858,N_1269,N_204);
xnor U9859 (N_9859,N_907,N_997);
and U9860 (N_9860,N_1642,N_52);
or U9861 (N_9861,N_3252,N_3632);
or U9862 (N_9862,N_1019,N_4938);
or U9863 (N_9863,N_2432,N_2834);
nand U9864 (N_9864,N_2488,N_1473);
and U9865 (N_9865,N_953,N_998);
or U9866 (N_9866,N_2096,N_307);
and U9867 (N_9867,N_4947,N_2401);
nor U9868 (N_9868,N_782,N_4749);
and U9869 (N_9869,N_2107,N_2512);
and U9870 (N_9870,N_4933,N_3107);
or U9871 (N_9871,N_2426,N_4734);
or U9872 (N_9872,N_2349,N_1465);
nand U9873 (N_9873,N_4189,N_3308);
and U9874 (N_9874,N_4342,N_2670);
nand U9875 (N_9875,N_649,N_2987);
and U9876 (N_9876,N_2790,N_1771);
or U9877 (N_9877,N_4024,N_2396);
nand U9878 (N_9878,N_4710,N_3153);
or U9879 (N_9879,N_3426,N_2554);
nand U9880 (N_9880,N_2297,N_3328);
and U9881 (N_9881,N_4853,N_3561);
and U9882 (N_9882,N_3518,N_4269);
xnor U9883 (N_9883,N_1459,N_4491);
or U9884 (N_9884,N_1424,N_1599);
and U9885 (N_9885,N_3906,N_888);
xor U9886 (N_9886,N_1608,N_2826);
or U9887 (N_9887,N_2166,N_4447);
nand U9888 (N_9888,N_817,N_2894);
or U9889 (N_9889,N_2289,N_325);
nor U9890 (N_9890,N_2609,N_972);
or U9891 (N_9891,N_1666,N_2313);
nor U9892 (N_9892,N_2105,N_3551);
nor U9893 (N_9893,N_170,N_2794);
and U9894 (N_9894,N_3620,N_3312);
nand U9895 (N_9895,N_1281,N_4336);
nand U9896 (N_9896,N_2989,N_3574);
nand U9897 (N_9897,N_3649,N_3976);
and U9898 (N_9898,N_1378,N_1812);
and U9899 (N_9899,N_4769,N_1675);
and U9900 (N_9900,N_30,N_2936);
nor U9901 (N_9901,N_169,N_3368);
and U9902 (N_9902,N_4792,N_2580);
xnor U9903 (N_9903,N_2896,N_2109);
and U9904 (N_9904,N_2865,N_3983);
or U9905 (N_9905,N_1848,N_4218);
xor U9906 (N_9906,N_4358,N_4567);
xnor U9907 (N_9907,N_4234,N_3283);
nand U9908 (N_9908,N_497,N_1488);
and U9909 (N_9909,N_2940,N_191);
nand U9910 (N_9910,N_486,N_2840);
or U9911 (N_9911,N_2901,N_2021);
nand U9912 (N_9912,N_3630,N_4453);
and U9913 (N_9913,N_1700,N_1918);
and U9914 (N_9914,N_4973,N_2509);
or U9915 (N_9915,N_1250,N_377);
nor U9916 (N_9916,N_4901,N_1798);
nand U9917 (N_9917,N_3799,N_921);
and U9918 (N_9918,N_701,N_723);
nand U9919 (N_9919,N_821,N_3791);
or U9920 (N_9920,N_2889,N_3169);
nor U9921 (N_9921,N_4503,N_3088);
or U9922 (N_9922,N_1248,N_2866);
nand U9923 (N_9923,N_4583,N_2086);
nor U9924 (N_9924,N_3578,N_494);
nor U9925 (N_9925,N_3525,N_2528);
nand U9926 (N_9926,N_1626,N_2558);
nand U9927 (N_9927,N_674,N_1235);
nand U9928 (N_9928,N_3422,N_1094);
nor U9929 (N_9929,N_2419,N_4760);
xor U9930 (N_9930,N_1320,N_2355);
nand U9931 (N_9931,N_988,N_4190);
nor U9932 (N_9932,N_4048,N_2989);
and U9933 (N_9933,N_4479,N_200);
nand U9934 (N_9934,N_1271,N_2028);
nor U9935 (N_9935,N_2025,N_1967);
or U9936 (N_9936,N_3929,N_560);
and U9937 (N_9937,N_3127,N_3814);
and U9938 (N_9938,N_850,N_1411);
and U9939 (N_9939,N_819,N_3617);
nand U9940 (N_9940,N_1101,N_1179);
and U9941 (N_9941,N_1313,N_955);
and U9942 (N_9942,N_3265,N_4116);
or U9943 (N_9943,N_34,N_4562);
nand U9944 (N_9944,N_732,N_4845);
nor U9945 (N_9945,N_4846,N_4515);
and U9946 (N_9946,N_2289,N_1588);
and U9947 (N_9947,N_722,N_3275);
and U9948 (N_9948,N_3811,N_1047);
xnor U9949 (N_9949,N_4004,N_2700);
nor U9950 (N_9950,N_2209,N_3135);
and U9951 (N_9951,N_929,N_304);
and U9952 (N_9952,N_25,N_468);
nor U9953 (N_9953,N_979,N_348);
and U9954 (N_9954,N_4488,N_1670);
nor U9955 (N_9955,N_295,N_3482);
xor U9956 (N_9956,N_3186,N_3685);
or U9957 (N_9957,N_2494,N_4493);
and U9958 (N_9958,N_598,N_4537);
nand U9959 (N_9959,N_1722,N_4020);
and U9960 (N_9960,N_1805,N_3755);
nor U9961 (N_9961,N_4260,N_659);
nand U9962 (N_9962,N_884,N_3547);
or U9963 (N_9963,N_1862,N_827);
nor U9964 (N_9964,N_1049,N_1397);
or U9965 (N_9965,N_3072,N_3259);
xor U9966 (N_9966,N_4449,N_3039);
or U9967 (N_9967,N_2865,N_640);
and U9968 (N_9968,N_2452,N_3388);
xnor U9969 (N_9969,N_2256,N_2986);
and U9970 (N_9970,N_25,N_982);
nand U9971 (N_9971,N_1667,N_4769);
nand U9972 (N_9972,N_235,N_3607);
nor U9973 (N_9973,N_745,N_1561);
nand U9974 (N_9974,N_4428,N_3968);
nand U9975 (N_9975,N_3124,N_615);
xor U9976 (N_9976,N_4484,N_1203);
and U9977 (N_9977,N_4035,N_3459);
nand U9978 (N_9978,N_4834,N_3138);
nor U9979 (N_9979,N_2584,N_1923);
nor U9980 (N_9980,N_972,N_2532);
or U9981 (N_9981,N_2852,N_2438);
nand U9982 (N_9982,N_383,N_4684);
or U9983 (N_9983,N_842,N_3253);
nor U9984 (N_9984,N_4946,N_2619);
nor U9985 (N_9985,N_2310,N_556);
nor U9986 (N_9986,N_268,N_3110);
nor U9987 (N_9987,N_1787,N_1957);
and U9988 (N_9988,N_4502,N_1610);
and U9989 (N_9989,N_814,N_4216);
xnor U9990 (N_9990,N_1604,N_361);
and U9991 (N_9991,N_72,N_154);
and U9992 (N_9992,N_2078,N_2964);
nand U9993 (N_9993,N_4375,N_4009);
or U9994 (N_9994,N_2312,N_4271);
xnor U9995 (N_9995,N_248,N_958);
and U9996 (N_9996,N_4007,N_367);
nor U9997 (N_9997,N_3631,N_2587);
and U9998 (N_9998,N_4389,N_2545);
nand U9999 (N_9999,N_4916,N_514);
xor UO_0 (O_0,N_6770,N_5270);
or UO_1 (O_1,N_5175,N_7689);
or UO_2 (O_2,N_8686,N_7529);
or UO_3 (O_3,N_6040,N_5228);
and UO_4 (O_4,N_8062,N_6187);
and UO_5 (O_5,N_5208,N_5235);
and UO_6 (O_6,N_5979,N_7862);
xor UO_7 (O_7,N_8180,N_6823);
nor UO_8 (O_8,N_6490,N_7586);
xnor UO_9 (O_9,N_7148,N_8512);
or UO_10 (O_10,N_5904,N_9851);
nand UO_11 (O_11,N_7280,N_5065);
or UO_12 (O_12,N_9692,N_8432);
nor UO_13 (O_13,N_5252,N_9997);
and UO_14 (O_14,N_5715,N_6748);
or UO_15 (O_15,N_9878,N_6357);
or UO_16 (O_16,N_6976,N_7986);
nor UO_17 (O_17,N_8519,N_9864);
or UO_18 (O_18,N_7056,N_5107);
xor UO_19 (O_19,N_7776,N_5874);
nand UO_20 (O_20,N_8918,N_8074);
xor UO_21 (O_21,N_6798,N_5358);
or UO_22 (O_22,N_7196,N_9955);
and UO_23 (O_23,N_6465,N_8007);
xor UO_24 (O_24,N_7916,N_8258);
and UO_25 (O_25,N_5736,N_8466);
or UO_26 (O_26,N_8371,N_7758);
nor UO_27 (O_27,N_8951,N_6230);
nor UO_28 (O_28,N_8095,N_8043);
nor UO_29 (O_29,N_9369,N_9417);
nand UO_30 (O_30,N_8099,N_5286);
and UO_31 (O_31,N_8214,N_6827);
or UO_32 (O_32,N_7402,N_6227);
and UO_33 (O_33,N_6917,N_6668);
nor UO_34 (O_34,N_7768,N_8010);
and UO_35 (O_35,N_7628,N_9235);
or UO_36 (O_36,N_7960,N_7054);
nor UO_37 (O_37,N_8633,N_6160);
and UO_38 (O_38,N_6458,N_6611);
nand UO_39 (O_39,N_8736,N_6268);
and UO_40 (O_40,N_5763,N_8564);
nand UO_41 (O_41,N_5556,N_6244);
nor UO_42 (O_42,N_5000,N_6751);
or UO_43 (O_43,N_8740,N_5101);
nand UO_44 (O_44,N_7572,N_9629);
nor UO_45 (O_45,N_8810,N_5610);
nand UO_46 (O_46,N_6636,N_8735);
and UO_47 (O_47,N_7759,N_7958);
nor UO_48 (O_48,N_5439,N_8813);
xor UO_49 (O_49,N_7642,N_8334);
nand UO_50 (O_50,N_9133,N_8756);
nand UO_51 (O_51,N_6715,N_8039);
or UO_52 (O_52,N_7130,N_9113);
and UO_53 (O_53,N_9734,N_9298);
and UO_54 (O_54,N_9948,N_8719);
nand UO_55 (O_55,N_5120,N_7560);
nand UO_56 (O_56,N_7446,N_7975);
nor UO_57 (O_57,N_7151,N_7968);
or UO_58 (O_58,N_9167,N_9403);
nand UO_59 (O_59,N_6546,N_5577);
and UO_60 (O_60,N_8666,N_7172);
and UO_61 (O_61,N_8793,N_7220);
or UO_62 (O_62,N_5207,N_9392);
nor UO_63 (O_63,N_6764,N_9199);
xor UO_64 (O_64,N_6693,N_7704);
nor UO_65 (O_65,N_8833,N_7005);
or UO_66 (O_66,N_5550,N_6997);
and UO_67 (O_67,N_6552,N_9993);
nand UO_68 (O_68,N_7578,N_9285);
nand UO_69 (O_69,N_6441,N_5435);
nand UO_70 (O_70,N_8779,N_5970);
and UO_71 (O_71,N_9248,N_9796);
nand UO_72 (O_72,N_6815,N_5012);
or UO_73 (O_73,N_9447,N_9558);
or UO_74 (O_74,N_7688,N_7580);
and UO_75 (O_75,N_8430,N_9435);
and UO_76 (O_76,N_9548,N_6947);
and UO_77 (O_77,N_6648,N_5745);
or UO_78 (O_78,N_8473,N_5968);
or UO_79 (O_79,N_9555,N_6398);
nand UO_80 (O_80,N_6891,N_8961);
xnor UO_81 (O_81,N_6713,N_6363);
and UO_82 (O_82,N_7488,N_8695);
nand UO_83 (O_83,N_9452,N_8706);
nand UO_84 (O_84,N_7679,N_7551);
nor UO_85 (O_85,N_9426,N_8534);
or UO_86 (O_86,N_6568,N_9825);
nor UO_87 (O_87,N_9320,N_9895);
or UO_88 (O_88,N_9516,N_8861);
xor UO_89 (O_89,N_9779,N_7493);
or UO_90 (O_90,N_5196,N_9632);
or UO_91 (O_91,N_6451,N_6733);
and UO_92 (O_92,N_8264,N_7246);
and UO_93 (O_93,N_5250,N_5394);
nand UO_94 (O_94,N_7015,N_9464);
and UO_95 (O_95,N_8130,N_8622);
nor UO_96 (O_96,N_9179,N_8767);
or UO_97 (O_97,N_9277,N_8004);
xor UO_98 (O_98,N_8591,N_6328);
or UO_99 (O_99,N_6353,N_5748);
or UO_100 (O_100,N_5637,N_5386);
or UO_101 (O_101,N_8167,N_7019);
or UO_102 (O_102,N_6466,N_6232);
nand UO_103 (O_103,N_7569,N_7420);
and UO_104 (O_104,N_7814,N_5621);
nor UO_105 (O_105,N_9151,N_6418);
and UO_106 (O_106,N_7545,N_8694);
nand UO_107 (O_107,N_8376,N_8186);
xor UO_108 (O_108,N_7946,N_8805);
or UO_109 (O_109,N_6861,N_7271);
or UO_110 (O_110,N_8569,N_9837);
and UO_111 (O_111,N_5367,N_9745);
nand UO_112 (O_112,N_6728,N_9960);
nor UO_113 (O_113,N_7046,N_9703);
nand UO_114 (O_114,N_9434,N_6410);
nor UO_115 (O_115,N_9917,N_7310);
xor UO_116 (O_116,N_8903,N_6304);
nor UO_117 (O_117,N_8057,N_9255);
nand UO_118 (O_118,N_9511,N_9666);
nand UO_119 (O_119,N_6974,N_6639);
nor UO_120 (O_120,N_6523,N_6395);
and UO_121 (O_121,N_9784,N_6542);
or UO_122 (O_122,N_5393,N_7588);
nand UO_123 (O_123,N_8696,N_5587);
nor UO_124 (O_124,N_5074,N_9067);
nand UO_125 (O_125,N_5727,N_6958);
or UO_126 (O_126,N_8143,N_6107);
nand UO_127 (O_127,N_5562,N_7353);
and UO_128 (O_128,N_6281,N_6133);
nor UO_129 (O_129,N_6135,N_8021);
or UO_130 (O_130,N_7816,N_7226);
or UO_131 (O_131,N_5329,N_6803);
nand UO_132 (O_132,N_6746,N_6509);
or UO_133 (O_133,N_9247,N_7608);
nor UO_134 (O_134,N_6525,N_6696);
nand UO_135 (O_135,N_7256,N_5628);
and UO_136 (O_136,N_5268,N_8920);
and UO_137 (O_137,N_5044,N_9090);
xnor UO_138 (O_138,N_6050,N_5530);
nor UO_139 (O_139,N_9495,N_9265);
and UO_140 (O_140,N_5411,N_9420);
xnor UO_141 (O_141,N_5023,N_6838);
nand UO_142 (O_142,N_7548,N_7191);
xnor UO_143 (O_143,N_7648,N_6768);
nor UO_144 (O_144,N_9181,N_7247);
and UO_145 (O_145,N_7400,N_5838);
or UO_146 (O_146,N_9946,N_6140);
nor UO_147 (O_147,N_7825,N_5547);
nor UO_148 (O_148,N_6347,N_8855);
nand UO_149 (O_149,N_6309,N_5723);
or UO_150 (O_150,N_6178,N_7504);
nand UO_151 (O_151,N_7435,N_7932);
nor UO_152 (O_152,N_5740,N_7736);
xnor UO_153 (O_153,N_7443,N_6291);
nand UO_154 (O_154,N_5842,N_7926);
nand UO_155 (O_155,N_5718,N_9036);
and UO_156 (O_156,N_7371,N_9873);
nor UO_157 (O_157,N_5466,N_5659);
nand UO_158 (O_158,N_5097,N_7654);
and UO_159 (O_159,N_9184,N_8864);
nor UO_160 (O_160,N_8956,N_9968);
and UO_161 (O_161,N_9858,N_9951);
nor UO_162 (O_162,N_7300,N_6651);
xnor UO_163 (O_163,N_9297,N_7397);
and UO_164 (O_164,N_5333,N_7842);
and UO_165 (O_165,N_5630,N_6323);
or UO_166 (O_166,N_6753,N_8191);
and UO_167 (O_167,N_7751,N_5456);
or UO_168 (O_168,N_7020,N_6782);
nand UO_169 (O_169,N_8478,N_7718);
nor UO_170 (O_170,N_8710,N_9210);
nand UO_171 (O_171,N_7407,N_5670);
or UO_172 (O_172,N_6780,N_6174);
and UO_173 (O_173,N_5942,N_6483);
nor UO_174 (O_174,N_9686,N_9479);
or UO_175 (O_175,N_5040,N_5130);
nand UO_176 (O_176,N_7132,N_6002);
nor UO_177 (O_177,N_5241,N_9517);
nor UO_178 (O_178,N_5519,N_6358);
nor UO_179 (O_179,N_7441,N_6329);
and UO_180 (O_180,N_7624,N_6723);
nand UO_181 (O_181,N_9860,N_9468);
or UO_182 (O_182,N_9428,N_6065);
and UO_183 (O_183,N_8230,N_9135);
xnor UO_184 (O_184,N_5622,N_5331);
or UO_185 (O_185,N_5450,N_6888);
nor UO_186 (O_186,N_9861,N_9419);
nand UO_187 (O_187,N_5284,N_9412);
and UO_188 (O_188,N_5339,N_7991);
and UO_189 (O_189,N_7531,N_9207);
and UO_190 (O_190,N_9079,N_5691);
xnor UO_191 (O_191,N_9883,N_7659);
or UO_192 (O_192,N_7045,N_6908);
nor UO_193 (O_193,N_5453,N_8117);
nor UO_194 (O_194,N_7253,N_6667);
nor UO_195 (O_195,N_7634,N_7442);
nor UO_196 (O_196,N_8356,N_8602);
and UO_197 (O_197,N_6327,N_9009);
and UO_198 (O_198,N_7161,N_8012);
nand UO_199 (O_199,N_6967,N_8225);
nand UO_200 (O_200,N_5377,N_7176);
xor UO_201 (O_201,N_5275,N_5912);
nand UO_202 (O_202,N_5242,N_8731);
nor UO_203 (O_203,N_6405,N_7336);
xor UO_204 (O_204,N_8570,N_6868);
nor UO_205 (O_205,N_7022,N_6734);
xnor UO_206 (O_206,N_7099,N_9990);
and UO_207 (O_207,N_7168,N_5364);
nor UO_208 (O_208,N_8407,N_7765);
xor UO_209 (O_209,N_6622,N_9357);
nand UO_210 (O_210,N_7516,N_9896);
nand UO_211 (O_211,N_5714,N_7413);
xor UO_212 (O_212,N_9083,N_7092);
and UO_213 (O_213,N_5271,N_9981);
nor UO_214 (O_214,N_6897,N_9114);
and UO_215 (O_215,N_7575,N_8557);
nor UO_216 (O_216,N_7109,N_7849);
nand UO_217 (O_217,N_6303,N_5548);
or UO_218 (O_218,N_8307,N_9925);
and UO_219 (O_219,N_8965,N_6158);
nand UO_220 (O_220,N_7309,N_7143);
and UO_221 (O_221,N_5708,N_7083);
nand UO_222 (O_222,N_7331,N_9939);
nor UO_223 (O_223,N_8263,N_5030);
nand UO_224 (O_224,N_6654,N_8635);
nor UO_225 (O_225,N_7500,N_7913);
and UO_226 (O_226,N_8597,N_6008);
nand UO_227 (O_227,N_6023,N_7055);
and UO_228 (O_228,N_5848,N_6545);
and UO_229 (O_229,N_5226,N_5455);
and UO_230 (O_230,N_6125,N_7165);
or UO_231 (O_231,N_6207,N_7093);
and UO_232 (O_232,N_9892,N_5588);
or UO_233 (O_233,N_8626,N_5581);
nor UO_234 (O_234,N_5945,N_8273);
and UO_235 (O_235,N_7379,N_8325);
nor UO_236 (O_236,N_8081,N_5353);
xnor UO_237 (O_237,N_7599,N_7291);
nor UO_238 (O_238,N_7567,N_5494);
and UO_239 (O_239,N_6324,N_5863);
or UO_240 (O_240,N_7279,N_8808);
nand UO_241 (O_241,N_5491,N_7517);
and UO_242 (O_242,N_8136,N_7684);
and UO_243 (O_243,N_9502,N_5502);
nor UO_244 (O_244,N_8536,N_8406);
nand UO_245 (O_245,N_5167,N_7095);
nor UO_246 (O_246,N_9268,N_8111);
nand UO_247 (O_247,N_6840,N_9042);
nor UO_248 (O_248,N_5933,N_8579);
nand UO_249 (O_249,N_9049,N_5820);
and UO_250 (O_250,N_8025,N_9243);
or UO_251 (O_251,N_5325,N_5645);
and UO_252 (O_252,N_6881,N_6496);
and UO_253 (O_253,N_5583,N_6689);
and UO_254 (O_254,N_9584,N_5761);
and UO_255 (O_255,N_5255,N_8960);
nor UO_256 (O_256,N_9767,N_7542);
nor UO_257 (O_257,N_7273,N_7002);
nand UO_258 (O_258,N_9828,N_9752);
nand UO_259 (O_259,N_6811,N_5159);
and UO_260 (O_260,N_9590,N_5619);
or UO_261 (O_261,N_6677,N_6257);
or UO_262 (O_262,N_6727,N_9020);
nand UO_263 (O_263,N_6522,N_5582);
xor UO_264 (O_264,N_7506,N_6557);
nand UO_265 (O_265,N_8262,N_5403);
nand UO_266 (O_266,N_5123,N_9589);
or UO_267 (O_267,N_7409,N_7249);
or UO_268 (O_268,N_7252,N_7389);
nand UO_269 (O_269,N_8384,N_5202);
and UO_270 (O_270,N_7620,N_5513);
or UO_271 (O_271,N_6092,N_8194);
nand UO_272 (O_272,N_7676,N_9797);
and UO_273 (O_273,N_8505,N_8929);
nor UO_274 (O_274,N_8601,N_6448);
nor UO_275 (O_275,N_6348,N_8341);
and UO_276 (O_276,N_8218,N_9719);
nand UO_277 (O_277,N_7138,N_7934);
nand UO_278 (O_278,N_8902,N_6331);
nand UO_279 (O_279,N_6384,N_6122);
and UO_280 (O_280,N_6415,N_7909);
or UO_281 (O_281,N_5446,N_9252);
nand UO_282 (O_282,N_9700,N_5893);
nand UO_283 (O_283,N_6952,N_6832);
or UO_284 (O_284,N_8868,N_9263);
and UO_285 (O_285,N_7163,N_8798);
nand UO_286 (O_286,N_7826,N_7125);
or UO_287 (O_287,N_7555,N_7683);
nand UO_288 (O_288,N_7292,N_8107);
nand UO_289 (O_289,N_7865,N_5110);
or UO_290 (O_290,N_7464,N_9577);
nand UO_291 (O_291,N_8983,N_5010);
nand UO_292 (O_292,N_7422,N_5374);
nand UO_293 (O_293,N_8209,N_6657);
or UO_294 (O_294,N_8817,N_6368);
or UO_295 (O_295,N_5853,N_5140);
and UO_296 (O_296,N_8690,N_8742);
or UO_297 (O_297,N_5066,N_6758);
and UO_298 (O_298,N_5758,N_6836);
nor UO_299 (O_299,N_7111,N_8231);
or UO_300 (O_300,N_6456,N_7269);
or UO_301 (O_301,N_8576,N_8522);
or UO_302 (O_302,N_9319,N_8465);
or UO_303 (O_303,N_5317,N_6873);
nor UO_304 (O_304,N_6739,N_8562);
nor UO_305 (O_305,N_6156,N_9764);
nand UO_306 (O_306,N_5535,N_6822);
nor UO_307 (O_307,N_6921,N_8245);
nor UO_308 (O_308,N_9775,N_9986);
nand UO_309 (O_309,N_9585,N_7466);
nor UO_310 (O_310,N_9786,N_6695);
and UO_311 (O_311,N_5383,N_6396);
and UO_312 (O_312,N_9085,N_6137);
nand UO_313 (O_313,N_8667,N_7147);
nor UO_314 (O_314,N_9910,N_5495);
nand UO_315 (O_315,N_5815,N_7031);
or UO_316 (O_316,N_7963,N_6287);
nand UO_317 (O_317,N_5388,N_6126);
or UO_318 (O_318,N_6749,N_5919);
nand UO_319 (O_319,N_6280,N_6212);
or UO_320 (O_320,N_5033,N_9660);
nand UO_321 (O_321,N_7121,N_5350);
nand UO_322 (O_322,N_9003,N_9901);
nor UO_323 (O_323,N_6108,N_9900);
or UO_324 (O_324,N_9762,N_7739);
xnor UO_325 (O_325,N_9073,N_8379);
nor UO_326 (O_326,N_9544,N_9250);
nor UO_327 (O_327,N_6901,N_7011);
xnor UO_328 (O_328,N_7017,N_7576);
nand UO_329 (O_329,N_8832,N_9066);
and UO_330 (O_330,N_6196,N_7326);
nand UO_331 (O_331,N_8521,N_9724);
nand UO_332 (O_332,N_7972,N_7737);
or UO_333 (O_333,N_7368,N_9217);
xor UO_334 (O_334,N_8016,N_9429);
nand UO_335 (O_335,N_8450,N_7396);
and UO_336 (O_336,N_5057,N_9538);
nor UO_337 (O_337,N_5644,N_6019);
nand UO_338 (O_338,N_8061,N_5128);
and UO_339 (O_339,N_6500,N_8027);
nand UO_340 (O_340,N_5669,N_7728);
nor UO_341 (O_341,N_9021,N_5267);
and UO_342 (O_342,N_7004,N_7501);
or UO_343 (O_343,N_5134,N_5785);
or UO_344 (O_344,N_5024,N_5307);
and UO_345 (O_345,N_6350,N_8036);
nor UO_346 (O_346,N_6067,N_6217);
xnor UO_347 (O_347,N_6834,N_7479);
nand UO_348 (O_348,N_7480,N_9756);
and UO_349 (O_349,N_7533,N_6539);
or UO_350 (O_350,N_8722,N_6605);
xnor UO_351 (O_351,N_9606,N_5218);
xnor UO_352 (O_352,N_5117,N_7394);
or UO_353 (O_353,N_5139,N_8673);
and UO_354 (O_354,N_9927,N_7964);
nor UO_355 (O_355,N_9404,N_9230);
nor UO_356 (O_356,N_8045,N_5096);
and UO_357 (O_357,N_7470,N_7519);
and UO_358 (O_358,N_7999,N_6098);
nand UO_359 (O_359,N_6761,N_9176);
or UO_360 (O_360,N_6419,N_7050);
and UO_361 (O_361,N_6162,N_9826);
nand UO_362 (O_362,N_7698,N_6297);
and UO_363 (O_363,N_9096,N_6634);
or UO_364 (O_364,N_7622,N_8758);
or UO_365 (O_365,N_9792,N_6799);
and UO_366 (O_366,N_8051,N_9368);
nand UO_367 (O_367,N_5730,N_5080);
nand UO_368 (O_368,N_7665,N_5198);
and UO_369 (O_369,N_9611,N_8571);
nor UO_370 (O_370,N_9805,N_7742);
nand UO_371 (O_371,N_9455,N_5867);
xnor UO_372 (O_372,N_5082,N_5844);
nand UO_373 (O_373,N_5314,N_8708);
nand UO_374 (O_374,N_6860,N_7908);
and UO_375 (O_375,N_6383,N_5533);
nand UO_376 (O_376,N_6660,N_9137);
or UO_377 (O_377,N_5655,N_7229);
nand UO_378 (O_378,N_8946,N_6111);
nor UO_379 (O_379,N_6276,N_8838);
nor UO_380 (O_380,N_7115,N_7360);
nor UO_381 (O_381,N_7085,N_9057);
nor UO_382 (O_382,N_6431,N_7503);
or UO_383 (O_383,N_5459,N_5506);
and UO_384 (O_384,N_8524,N_8018);
and UO_385 (O_385,N_8504,N_8125);
nand UO_386 (O_386,N_5295,N_7887);
nand UO_387 (O_387,N_5552,N_7127);
or UO_388 (O_388,N_7613,N_7839);
nor UO_389 (O_389,N_5183,N_8358);
nand UO_390 (O_390,N_9982,N_7320);
nor UO_391 (O_391,N_8594,N_6903);
xor UO_392 (O_392,N_5611,N_8786);
and UO_393 (O_393,N_9458,N_9162);
nand UO_394 (O_394,N_6988,N_7073);
nor UO_395 (O_395,N_6537,N_6474);
or UO_396 (O_396,N_5857,N_5319);
and UO_397 (O_397,N_8785,N_6950);
and UO_398 (O_398,N_6105,N_8424);
and UO_399 (O_399,N_6965,N_5825);
nor UO_400 (O_400,N_6745,N_8795);
nand UO_401 (O_401,N_5993,N_5342);
nand UO_402 (O_402,N_8005,N_6747);
or UO_403 (O_403,N_7602,N_7415);
or UO_404 (O_404,N_7417,N_9559);
xor UO_405 (O_405,N_5373,N_6293);
or UO_406 (O_406,N_5733,N_5877);
nor UO_407 (O_407,N_9448,N_8691);
nand UO_408 (O_408,N_8458,N_8219);
or UO_409 (O_409,N_8857,N_5344);
and UO_410 (O_410,N_7583,N_6837);
nor UO_411 (O_411,N_8459,N_6186);
nand UO_412 (O_412,N_7706,N_5716);
and UO_413 (O_413,N_8925,N_5629);
nand UO_414 (O_414,N_5505,N_5118);
nand UO_415 (O_415,N_8816,N_6189);
xnor UO_416 (O_416,N_9233,N_9682);
and UO_417 (O_417,N_9527,N_7527);
xnor UO_418 (O_418,N_8869,N_5467);
nand UO_419 (O_419,N_7880,N_6077);
xor UO_420 (O_420,N_9336,N_7301);
xnor UO_421 (O_421,N_7770,N_5472);
and UO_422 (O_422,N_9523,N_5937);
and UO_423 (O_423,N_8076,N_9496);
and UO_424 (O_424,N_6058,N_5633);
nor UO_425 (O_425,N_9650,N_7465);
and UO_426 (O_426,N_9803,N_7129);
nand UO_427 (O_427,N_7060,N_6031);
nor UO_428 (O_428,N_7871,N_9424);
nand UO_429 (O_429,N_5759,N_6045);
nand UO_430 (O_430,N_5019,N_5396);
or UO_431 (O_431,N_5966,N_8975);
nand UO_432 (O_432,N_7875,N_7203);
or UO_433 (O_433,N_5778,N_7752);
or UO_434 (O_434,N_7745,N_9220);
nand UO_435 (O_435,N_5070,N_6390);
and UO_436 (O_436,N_9329,N_9237);
or UO_437 (O_437,N_8939,N_8105);
xor UO_438 (O_438,N_8775,N_9765);
nand UO_439 (O_439,N_5754,N_8393);
or UO_440 (O_440,N_5807,N_8663);
nor UO_441 (O_441,N_9224,N_9875);
and UO_442 (O_442,N_9308,N_5961);
nor UO_443 (O_443,N_8717,N_6754);
and UO_444 (O_444,N_7423,N_8531);
and UO_445 (O_445,N_6147,N_9662);
nand UO_446 (O_446,N_8907,N_8019);
and UO_447 (O_447,N_9531,N_7190);
nor UO_448 (O_448,N_9552,N_7117);
or UO_449 (O_449,N_5692,N_8778);
nand UO_450 (O_450,N_5965,N_9716);
nor UO_451 (O_451,N_7873,N_8616);
and UO_452 (O_452,N_9942,N_6020);
nor UO_453 (O_453,N_6346,N_6878);
xor UO_454 (O_454,N_7359,N_6843);
nand UO_455 (O_455,N_9713,N_6269);
nor UO_456 (O_456,N_5773,N_8984);
nor UO_457 (O_457,N_8181,N_7355);
nor UO_458 (O_458,N_6612,N_9105);
nor UO_459 (O_459,N_7180,N_5083);
nor UO_460 (O_460,N_8471,N_7463);
xnor UO_461 (O_461,N_8528,N_5184);
and UO_462 (O_462,N_7925,N_9833);
nand UO_463 (O_463,N_5928,N_8347);
and UO_464 (O_464,N_5667,N_8968);
xor UO_465 (O_465,N_9087,N_5543);
nor UO_466 (O_466,N_9778,N_6237);
xnor UO_467 (O_467,N_8041,N_8713);
and UO_468 (O_468,N_5632,N_7255);
and UO_469 (O_469,N_6344,N_5626);
nor UO_470 (O_470,N_9674,N_7486);
and UO_471 (O_471,N_9602,N_6618);
xor UO_472 (O_472,N_7156,N_6641);
nor UO_473 (O_473,N_7189,N_9299);
nand UO_474 (O_474,N_6286,N_7796);
nor UO_475 (O_475,N_8260,N_9306);
or UO_476 (O_476,N_7462,N_5043);
xor UO_477 (O_477,N_8103,N_8653);
or UO_478 (O_478,N_7308,N_7072);
nand UO_479 (O_479,N_6769,N_5157);
or UO_480 (O_480,N_9835,N_8862);
nor UO_481 (O_481,N_6084,N_9394);
xor UO_482 (O_482,N_7079,N_9922);
nand UO_483 (O_483,N_8692,N_6176);
xnor UO_484 (O_484,N_5496,N_8281);
nand UO_485 (O_485,N_9112,N_9882);
nor UO_486 (O_486,N_9385,N_8535);
xnor UO_487 (O_487,N_6561,N_7267);
and UO_488 (O_488,N_6517,N_7753);
nor UO_489 (O_489,N_5521,N_6424);
and UO_490 (O_490,N_8912,N_5846);
or UO_491 (O_491,N_8584,N_8502);
or UO_492 (O_492,N_6587,N_9549);
or UO_493 (O_493,N_8174,N_9342);
and UO_494 (O_494,N_6809,N_7982);
nand UO_495 (O_495,N_8177,N_8060);
or UO_496 (O_496,N_8561,N_9958);
or UO_497 (O_497,N_6529,N_6777);
nand UO_498 (O_498,N_8998,N_8000);
nor UO_499 (O_499,N_7918,N_7799);
nand UO_500 (O_500,N_5302,N_6364);
nor UO_501 (O_501,N_5263,N_6828);
and UO_502 (O_502,N_9165,N_7579);
nand UO_503 (O_503,N_6371,N_6676);
or UO_504 (O_504,N_7087,N_9507);
and UO_505 (O_505,N_8993,N_9023);
or UO_506 (O_506,N_7597,N_5999);
xnor UO_507 (O_507,N_9290,N_9363);
or UO_508 (O_508,N_8215,N_7007);
and UO_509 (O_509,N_8905,N_6128);
and UO_510 (O_510,N_9171,N_6316);
or UO_511 (O_511,N_7811,N_8792);
nand UO_512 (O_512,N_6263,N_6659);
nand UO_513 (O_513,N_8441,N_7043);
or UO_514 (O_514,N_5076,N_8400);
nor UO_515 (O_515,N_6972,N_8515);
xnor UO_516 (O_516,N_7106,N_5826);
nand UO_517 (O_517,N_5693,N_7123);
nor UO_518 (O_518,N_9920,N_8370);
nor UO_519 (O_519,N_9229,N_8088);
or UO_520 (O_520,N_5894,N_9869);
nand UO_521 (O_521,N_5953,N_6533);
or UO_522 (O_522,N_5606,N_9402);
nand UO_523 (O_523,N_5664,N_8295);
or UO_524 (O_524,N_5917,N_7094);
nor UO_525 (O_525,N_7534,N_5300);
nand UO_526 (O_526,N_9249,N_6295);
nor UO_527 (O_527,N_8444,N_6294);
nor UO_528 (O_528,N_5855,N_9366);
nor UO_529 (O_529,N_5498,N_7090);
nor UO_530 (O_530,N_5812,N_9831);
nor UO_531 (O_531,N_9493,N_7860);
nand UO_532 (O_532,N_7289,N_8001);
or UO_533 (O_533,N_6985,N_9142);
or UO_534 (O_534,N_8359,N_9031);
xor UO_535 (O_535,N_6859,N_8852);
nand UO_536 (O_536,N_5954,N_9156);
or UO_537 (O_537,N_5501,N_9132);
and UO_538 (O_538,N_5077,N_8484);
and UO_539 (O_539,N_8734,N_6895);
nand UO_540 (O_540,N_6172,N_8607);
xnor UO_541 (O_541,N_9065,N_5634);
or UO_542 (O_542,N_5658,N_7003);
and UO_543 (O_543,N_8070,N_6277);
nor UO_544 (O_544,N_6200,N_6422);
and UO_545 (O_545,N_8460,N_9407);
nand UO_546 (O_546,N_5280,N_5346);
or UO_547 (O_547,N_8727,N_8870);
nand UO_548 (O_548,N_5660,N_6446);
nor UO_549 (O_549,N_5803,N_6219);
or UO_550 (O_550,N_8682,N_5234);
or UO_551 (O_551,N_8101,N_8585);
or UO_552 (O_552,N_8092,N_9726);
nand UO_553 (O_553,N_6998,N_6617);
and UO_554 (O_554,N_6204,N_8685);
nor UO_555 (O_555,N_6018,N_9194);
nand UO_556 (O_556,N_7395,N_5760);
nand UO_557 (O_557,N_6491,N_5404);
and UO_558 (O_558,N_9581,N_6786);
or UO_559 (O_559,N_5108,N_7921);
and UO_560 (O_560,N_8169,N_9760);
and UO_561 (O_561,N_8765,N_6551);
nor UO_562 (O_562,N_6194,N_7059);
nand UO_563 (O_563,N_8461,N_9274);
nor UO_564 (O_564,N_5567,N_6678);
or UO_565 (O_565,N_7969,N_5162);
nor UO_566 (O_566,N_7794,N_9406);
nor UO_567 (O_567,N_6646,N_5964);
or UO_568 (O_568,N_8129,N_9935);
nor UO_569 (O_569,N_5440,N_6510);
nand UO_570 (O_570,N_9999,N_8298);
nand UO_571 (O_571,N_6149,N_9919);
xnor UO_572 (O_572,N_6885,N_9187);
and UO_573 (O_573,N_8831,N_5007);
nand UO_574 (O_574,N_8316,N_7941);
and UO_575 (O_575,N_7281,N_5725);
xnor UO_576 (O_576,N_6349,N_5131);
or UO_577 (O_577,N_8135,N_8418);
or UO_578 (O_578,N_9654,N_8590);
or UO_579 (O_579,N_7455,N_8159);
nor UO_580 (O_580,N_8698,N_6097);
nor UO_581 (O_581,N_5151,N_7530);
nand UO_582 (O_582,N_7234,N_8513);
or UO_583 (O_583,N_7663,N_5203);
or UO_584 (O_584,N_9633,N_5086);
nor UO_585 (O_585,N_9382,N_8412);
nor UO_586 (O_586,N_8991,N_5525);
and UO_587 (O_587,N_5251,N_7146);
xor UO_588 (O_588,N_8324,N_6145);
nand UO_589 (O_589,N_6870,N_7110);
nor UO_590 (O_590,N_9197,N_8054);
nor UO_591 (O_591,N_9761,N_6497);
nand UO_592 (O_592,N_8291,N_6402);
or UO_593 (O_593,N_7984,N_8807);
or UO_594 (O_594,N_9275,N_9123);
nor UO_595 (O_595,N_5819,N_5324);
nor UO_596 (O_596,N_6710,N_8503);
nand UO_597 (O_597,N_9373,N_8718);
xor UO_598 (O_598,N_8006,N_8739);
and UO_599 (O_599,N_9758,N_5794);
nor UO_600 (O_600,N_6342,N_6375);
nand UO_601 (O_601,N_7223,N_8380);
nor UO_602 (O_602,N_6812,N_9741);
nand UO_603 (O_603,N_9739,N_7366);
nor UO_604 (O_604,N_5986,N_9293);
nor UO_605 (O_605,N_6225,N_6979);
nor UO_606 (O_606,N_5639,N_8620);
and UO_607 (O_607,N_8532,N_8318);
and UO_608 (O_608,N_7134,N_7844);
and UO_609 (O_609,N_6004,N_7403);
and UO_610 (O_610,N_6919,N_7725);
nor UO_611 (O_611,N_8055,N_9117);
nand UO_612 (O_612,N_9387,N_8335);
or UO_613 (O_613,N_8020,N_8958);
and UO_614 (O_614,N_6896,N_9084);
and UO_615 (O_615,N_6948,N_9222);
nor UO_616 (O_616,N_9198,N_8467);
nor UO_617 (O_617,N_6935,N_9723);
nand UO_618 (O_618,N_8419,N_7013);
xnor UO_619 (O_619,N_5821,N_8788);
or UO_620 (O_620,N_5164,N_7122);
nand UO_621 (O_621,N_8189,N_6794);
and UO_622 (O_622,N_9152,N_5220);
nand UO_623 (O_623,N_5069,N_7427);
or UO_624 (O_624,N_7606,N_5902);
xnor UO_625 (O_625,N_5950,N_5854);
and UO_626 (O_626,N_8163,N_8963);
or UO_627 (O_627,N_9928,N_7448);
and UO_628 (O_628,N_8455,N_9494);
xnor UO_629 (O_629,N_6355,N_6425);
nand UO_630 (O_630,N_8362,N_8543);
or UO_631 (O_631,N_5109,N_9678);
nand UO_632 (O_632,N_5746,N_8097);
nand UO_633 (O_633,N_8676,N_6080);
nand UO_634 (O_634,N_6642,N_7756);
nand UO_635 (O_635,N_9370,N_8434);
or UO_636 (O_636,N_7869,N_5310);
nand UO_637 (O_637,N_7762,N_6265);
nor UO_638 (O_638,N_9963,N_9620);
or UO_639 (O_639,N_5484,N_6797);
or UO_640 (O_640,N_7169,N_7956);
or UO_641 (O_641,N_9473,N_5071);
nor UO_642 (O_642,N_7640,N_8650);
xor UO_643 (O_643,N_9477,N_5136);
nand UO_644 (O_644,N_5004,N_8477);
nand UO_645 (O_645,N_9449,N_8178);
nor UO_646 (O_646,N_8642,N_7966);
or UO_647 (O_647,N_9995,N_5915);
nand UO_648 (O_648,N_9720,N_5817);
nor UO_649 (O_649,N_9027,N_9912);
and UO_650 (O_650,N_8402,N_9149);
and UO_651 (O_651,N_8403,N_5783);
nand UO_652 (O_652,N_6892,N_7509);
nor UO_653 (O_653,N_5997,N_9649);
or UO_654 (O_654,N_7297,N_5982);
nand UO_655 (O_655,N_5355,N_7820);
and UO_656 (O_656,N_6957,N_7483);
or UO_657 (O_657,N_6742,N_9499);
and UO_658 (O_658,N_7910,N_6995);
or UO_659 (O_659,N_6254,N_8881);
and UO_660 (O_660,N_5523,N_5764);
and UO_661 (O_661,N_9415,N_5884);
or UO_662 (O_662,N_9467,N_7096);
or UO_663 (O_663,N_7717,N_9753);
and UO_664 (O_664,N_6684,N_7644);
nor UO_665 (O_665,N_7347,N_5540);
xor UO_666 (O_666,N_8850,N_9601);
and UO_667 (O_667,N_9604,N_6598);
and UO_668 (O_668,N_8102,N_8538);
or UO_669 (O_669,N_8542,N_9457);
nor UO_670 (O_670,N_6201,N_9699);
and UO_671 (O_671,N_9124,N_8374);
nor UO_672 (O_672,N_8104,N_6071);
or UO_673 (O_673,N_5542,N_6132);
or UO_674 (O_674,N_5642,N_5259);
nor UO_675 (O_675,N_9380,N_6905);
and UO_676 (O_676,N_7631,N_9725);
nand UO_677 (O_677,N_9603,N_5775);
nand UO_678 (O_678,N_7781,N_9809);
xor UO_679 (O_679,N_8274,N_9343);
nand UO_680 (O_680,N_5221,N_8408);
nand UO_681 (O_681,N_7216,N_7254);
nand UO_682 (O_682,N_5122,N_7905);
xor UO_683 (O_683,N_9742,N_9550);
xor UO_684 (O_684,N_6171,N_9906);
or UO_685 (O_685,N_5514,N_6984);
and UO_686 (O_686,N_9030,N_7681);
xnor UO_687 (O_687,N_6279,N_6464);
xor UO_688 (O_688,N_9498,N_9594);
or UO_689 (O_689,N_9232,N_9868);
nor UO_690 (O_690,N_7929,N_6003);
xor UO_691 (O_691,N_6824,N_8259);
and UO_692 (O_692,N_5338,N_8669);
nor UO_693 (O_693,N_8530,N_8581);
nand UO_694 (O_694,N_6153,N_5870);
or UO_695 (O_695,N_7459,N_8085);
nand UO_696 (O_696,N_8820,N_7870);
and UO_697 (O_697,N_5721,N_6702);
and UO_698 (O_698,N_8275,N_7513);
and UO_699 (O_699,N_6658,N_5766);
nand UO_700 (O_700,N_6063,N_5625);
and UO_701 (O_701,N_6221,N_9506);
nand UO_702 (O_702,N_7537,N_7965);
and UO_703 (O_703,N_6216,N_6721);
and UO_704 (O_704,N_5356,N_6030);
and UO_705 (O_705,N_5470,N_7696);
nor UO_706 (O_706,N_9623,N_8957);
nand UO_707 (O_707,N_9565,N_6032);
nor UO_708 (O_708,N_9240,N_6662);
and UO_709 (O_709,N_9657,N_6544);
and UO_710 (O_710,N_9106,N_8243);
nor UO_711 (O_711,N_7307,N_6101);
or UO_712 (O_712,N_9119,N_9150);
and UO_713 (O_713,N_5719,N_7646);
nor UO_714 (O_714,N_8548,N_6179);
or UO_715 (O_715,N_9988,N_8517);
or UO_716 (O_716,N_5990,N_8702);
nand UO_717 (O_717,N_9192,N_8728);
nand UO_718 (O_718,N_6681,N_5429);
and UO_719 (O_719,N_7701,N_6652);
or UO_720 (O_720,N_9183,N_8002);
nand UO_721 (O_721,N_7290,N_6492);
nor UO_722 (O_722,N_7853,N_6027);
nor UO_723 (O_723,N_6688,N_6220);
nor UO_724 (O_724,N_8026,N_6123);
nor UO_725 (O_725,N_8014,N_6601);
or UO_726 (O_726,N_9505,N_6009);
nand UO_727 (O_727,N_5451,N_9337);
or UO_728 (O_728,N_8979,N_5801);
and UO_729 (O_729,N_6454,N_8416);
and UO_730 (O_730,N_9488,N_5049);
nand UO_731 (O_731,N_6487,N_8636);
and UO_732 (O_732,N_7014,N_6089);
nand UO_733 (O_733,N_6938,N_7288);
nor UO_734 (O_734,N_5378,N_8414);
nand UO_735 (O_735,N_6115,N_5090);
and UO_736 (O_736,N_8574,N_6796);
and UO_737 (O_737,N_5017,N_7993);
nor UO_738 (O_738,N_5054,N_7823);
nor UO_739 (O_739,N_6914,N_8445);
nor UO_740 (O_740,N_5189,N_9593);
nand UO_741 (O_741,N_9358,N_9812);
and UO_742 (O_742,N_5294,N_9874);
nand UO_743 (O_743,N_6356,N_6307);
xor UO_744 (O_744,N_8413,N_8614);
and UO_745 (O_745,N_6131,N_6447);
xor UO_746 (O_746,N_6503,N_5651);
nor UO_747 (O_747,N_5390,N_5962);
and UO_748 (O_748,N_5767,N_8761);
or UO_749 (O_749,N_7703,N_8138);
and UO_750 (O_750,N_9754,N_8799);
nor UO_751 (O_751,N_9076,N_8748);
nor UO_752 (O_752,N_5059,N_9781);
xnor UO_753 (O_753,N_5354,N_9396);
or UO_754 (O_754,N_5504,N_5266);
and UO_755 (O_755,N_7846,N_6707);
nand UO_756 (O_756,N_7980,N_9879);
or UO_757 (O_757,N_7617,N_5555);
and UO_758 (O_758,N_8580,N_5975);
xnor UO_759 (O_759,N_7894,N_7318);
or UO_760 (O_760,N_9024,N_8658);
and UO_761 (O_761,N_9526,N_6576);
or UO_762 (O_762,N_9007,N_8415);
xnor UO_763 (O_763,N_9116,N_9731);
nor UO_764 (O_764,N_5316,N_8496);
nor UO_765 (O_765,N_9190,N_8329);
nand UO_766 (O_766,N_7390,N_6912);
nor UO_767 (O_767,N_7218,N_5636);
or UO_768 (O_768,N_7239,N_7433);
or UO_769 (O_769,N_5687,N_9612);
xor UO_770 (O_770,N_8032,N_7494);
xor UO_771 (O_771,N_9006,N_8405);
and UO_772 (O_772,N_7323,N_8646);
xor UO_773 (O_773,N_8192,N_7328);
nand UO_774 (O_774,N_5438,N_8206);
nand UO_775 (O_775,N_9454,N_8743);
or UO_776 (O_776,N_9980,N_8959);
or UO_777 (O_777,N_7573,N_9362);
nor UO_778 (O_778,N_7748,N_9656);
nand UO_779 (O_779,N_9281,N_8127);
or UO_780 (O_780,N_9715,N_7804);
nor UO_781 (O_781,N_5677,N_9153);
or UO_782 (O_782,N_9389,N_6213);
nor UO_783 (O_783,N_5230,N_5039);
nand UO_784 (O_784,N_5868,N_9820);
or UO_785 (O_785,N_7299,N_8132);
nand UO_786 (O_786,N_8472,N_6528);
nor UO_787 (O_787,N_9055,N_6978);
nor UO_788 (O_788,N_7035,N_5798);
and UO_789 (O_789,N_9391,N_6462);
and UO_790 (O_790,N_8897,N_9344);
or UO_791 (O_791,N_8464,N_9547);
or UO_792 (O_792,N_8269,N_9641);
xor UO_793 (O_793,N_8688,N_5124);
and UO_794 (O_794,N_9553,N_5865);
and UO_795 (O_795,N_8649,N_7051);
nand UO_796 (O_796,N_6626,N_9818);
nand UO_797 (O_797,N_6690,N_8320);
nand UO_798 (O_798,N_6296,N_9186);
nor UO_799 (O_799,N_8630,N_9608);
nand UO_800 (O_800,N_5322,N_8520);
or UO_801 (O_801,N_7981,N_9286);
nor UO_802 (O_802,N_7920,N_6595);
nand UO_803 (O_803,N_9576,N_8293);
nor UO_804 (O_804,N_7655,N_5214);
nor UO_805 (O_805,N_8108,N_8977);
and UO_806 (O_806,N_7375,N_8851);
nor UO_807 (O_807,N_9052,N_8615);
or UO_808 (O_808,N_8997,N_6619);
nand UO_809 (O_809,N_7449,N_8760);
nor UO_810 (O_810,N_8257,N_5022);
and UO_811 (O_811,N_5088,N_6638);
nor UO_812 (O_812,N_6531,N_8453);
nand UO_813 (O_813,N_9214,N_7915);
nor UO_814 (O_814,N_5907,N_6206);
and UO_815 (O_815,N_9711,N_9634);
or UO_816 (O_816,N_8940,N_8701);
or UO_817 (O_817,N_6061,N_5113);
and UO_818 (O_818,N_8428,N_8797);
and UO_819 (O_819,N_6233,N_7726);
nand UO_820 (O_820,N_8063,N_8865);
nor UO_821 (O_821,N_5638,N_8843);
nor UO_822 (O_822,N_8729,N_8352);
or UO_823 (O_823,N_5303,N_5922);
and UO_824 (O_824,N_6981,N_8008);
and UO_825 (O_825,N_8368,N_5601);
and UO_826 (O_826,N_7711,N_8715);
and UO_827 (O_827,N_5998,N_9289);
nor UO_828 (O_828,N_7953,N_7278);
and UO_829 (O_829,N_9216,N_8198);
and UO_830 (O_830,N_7061,N_6238);
nor UO_831 (O_831,N_9242,N_8628);
and UO_832 (O_832,N_9880,N_5534);
or UO_833 (O_833,N_6603,N_8351);
and UO_834 (O_834,N_9376,N_6910);
nor UO_835 (O_835,N_9738,N_6472);
and UO_836 (O_836,N_6203,N_6954);
nor UO_837 (O_837,N_5111,N_7142);
and UO_838 (O_838,N_5656,N_6006);
and UO_839 (O_839,N_5987,N_7619);
nor UO_840 (O_840,N_9077,N_7044);
nor UO_841 (O_841,N_5372,N_8689);
nor UO_842 (O_842,N_7208,N_7937);
nand UO_843 (O_843,N_8300,N_6564);
nor UO_844 (O_844,N_9834,N_5710);
xor UO_845 (O_845,N_9510,N_8139);
nand UO_846 (O_846,N_6182,N_6426);
or UO_847 (O_847,N_5809,N_8592);
and UO_848 (O_848,N_8398,N_5304);
or UO_849 (O_849,N_8849,N_9866);
nor UO_850 (O_850,N_6936,N_9645);
nand UO_851 (O_851,N_9721,N_6876);
nand UO_852 (O_852,N_7743,N_7401);
nand UO_853 (O_853,N_8475,N_8087);
or UO_854 (O_854,N_8879,N_6442);
and UO_855 (O_855,N_9921,N_6756);
or UO_856 (O_856,N_9575,N_6513);
nand UO_857 (O_857,N_5094,N_6055);
and UO_858 (O_858,N_6113,N_8899);
nand UO_859 (O_859,N_7514,N_5881);
nor UO_860 (O_860,N_8773,N_9850);
nand UO_861 (O_861,N_7227,N_7593);
nand UO_862 (O_862,N_6035,N_9798);
nor UO_863 (O_863,N_7577,N_8995);
nor UO_864 (O_864,N_5604,N_5948);
or UO_865 (O_865,N_5464,N_7955);
and UO_866 (O_866,N_9206,N_9282);
or UO_867 (O_867,N_9004,N_6675);
nor UO_868 (O_868,N_7668,N_9722);
nand UO_869 (O_869,N_7732,N_8853);
nand UO_870 (O_870,N_8035,N_6880);
nand UO_871 (O_871,N_5011,N_6795);
and UO_872 (O_872,N_7261,N_8674);
and UO_873 (O_873,N_8506,N_6818);
or UO_874 (O_874,N_7774,N_8880);
and UO_875 (O_875,N_7891,N_7052);
nor UO_876 (O_876,N_6508,N_8469);
or UO_877 (O_877,N_8553,N_6923);
nand UO_878 (O_878,N_7878,N_6977);
nand UO_879 (O_879,N_9118,N_5477);
nand UO_880 (O_880,N_8160,N_5887);
nand UO_881 (O_881,N_9044,N_8552);
nand UO_882 (O_882,N_7543,N_5570);
nand UO_883 (O_883,N_8967,N_8559);
and UO_884 (O_884,N_5443,N_9859);
nand UO_885 (O_885,N_9876,N_6574);
and UO_886 (O_886,N_6590,N_6223);
and UO_887 (O_887,N_7345,N_8118);
and UO_888 (O_888,N_9940,N_5285);
nor UO_889 (O_889,N_6940,N_6514);
or UO_890 (O_890,N_5614,N_8643);
nor UO_891 (O_891,N_8009,N_8497);
nand UO_892 (O_892,N_7036,N_9838);
nor UO_893 (O_893,N_9648,N_7312);
and UO_894 (O_894,N_7852,N_9377);
and UO_895 (O_895,N_9321,N_7919);
nor UO_896 (O_896,N_6195,N_5231);
nor UO_897 (O_897,N_7460,N_7033);
nand UO_898 (O_898,N_8151,N_6581);
nor UO_899 (O_899,N_8752,N_7611);
and UO_900 (O_900,N_6929,N_9459);
nand UO_901 (O_901,N_5509,N_8640);
nand UO_902 (O_902,N_9975,N_9219);
xnor UO_903 (O_903,N_9551,N_7450);
nand UO_904 (O_904,N_7957,N_5858);
or UO_905 (O_905,N_7369,N_5436);
xnor UO_906 (O_906,N_8612,N_5402);
nor UO_907 (O_907,N_7840,N_8480);
or UO_908 (O_908,N_5379,N_7935);
xor UO_909 (O_909,N_8144,N_6072);
nand UO_910 (O_910,N_8279,N_5592);
and UO_911 (O_911,N_8284,N_8927);
and UO_912 (O_912,N_9887,N_5566);
nor UO_913 (O_913,N_7245,N_5493);
or UO_914 (O_914,N_9346,N_9461);
nor UO_915 (O_915,N_9058,N_8369);
nand UO_916 (O_916,N_8487,N_9037);
xor UO_917 (O_917,N_6906,N_6007);
and UO_918 (O_918,N_7818,N_6501);
nor UO_919 (O_919,N_7171,N_5298);
or UO_920 (O_920,N_7848,N_8050);
nor UO_921 (O_921,N_8457,N_5729);
nor UO_922 (O_922,N_9463,N_8211);
nand UO_923 (O_923,N_9080,N_5434);
or UO_924 (O_924,N_8110,N_5428);
and UO_925 (O_925,N_6175,N_5261);
xnor UO_926 (O_926,N_7373,N_5205);
and UO_927 (O_927,N_6712,N_8901);
nor UO_928 (O_928,N_7761,N_7612);
and UO_929 (O_929,N_8750,N_6991);
nand UO_930 (O_930,N_5934,N_9774);
xnor UO_931 (O_931,N_8323,N_7805);
and UO_932 (O_932,N_8312,N_7221);
nand UO_933 (O_933,N_9973,N_9422);
nor UO_934 (O_934,N_7518,N_9173);
or UO_935 (O_935,N_8395,N_6409);
or UO_936 (O_936,N_8829,N_8510);
nand UO_937 (O_937,N_5784,N_8937);
nand UO_938 (O_938,N_6502,N_8826);
xor UO_939 (O_939,N_7675,N_7747);
nor UO_940 (O_940,N_5002,N_7831);
nand UO_941 (O_941,N_7062,N_9451);
nand UO_942 (O_942,N_5974,N_6168);
xor UO_943 (O_943,N_7207,N_7179);
nor UO_944 (O_944,N_5685,N_5576);
nand UO_945 (O_945,N_9439,N_9795);
nor UO_946 (O_946,N_7694,N_8309);
and UO_947 (O_947,N_8410,N_5891);
and UO_948 (O_948,N_5376,N_8800);
and UO_949 (O_949,N_8634,N_9166);
nor UO_950 (O_950,N_5194,N_6022);
nor UO_951 (O_951,N_6714,N_7760);
and UO_952 (O_952,N_5770,N_5847);
nand UO_953 (O_953,N_6530,N_6983);
nand UO_954 (O_954,N_8839,N_6317);
and UO_955 (O_955,N_5910,N_7550);
and UO_956 (O_956,N_7876,N_6130);
nor UO_957 (O_957,N_6644,N_8096);
or UO_958 (O_958,N_5983,N_6173);
or UO_959 (O_959,N_8704,N_5177);
nand UO_960 (O_960,N_8603,N_9899);
or UO_961 (O_961,N_7610,N_5616);
and UO_962 (O_962,N_8411,N_6208);
xor UO_963 (O_963,N_9894,N_8197);
and UO_964 (O_964,N_7173,N_7510);
or UO_965 (O_965,N_6680,N_5900);
nand UO_966 (O_966,N_5834,N_8896);
nand UO_967 (O_967,N_5006,N_7357);
or UO_968 (O_968,N_8866,N_6498);
or UO_969 (O_969,N_6504,N_9082);
nor UO_970 (O_970,N_8239,N_8587);
and UO_971 (O_971,N_9513,N_9907);
or UO_972 (O_972,N_8809,N_5182);
or UO_973 (O_973,N_8846,N_6924);
xor UO_974 (O_974,N_6479,N_6591);
nand UO_975 (O_975,N_5119,N_8610);
and UO_976 (O_976,N_5739,N_6499);
and UO_977 (O_977,N_6907,N_5262);
nor UO_978 (O_978,N_7485,N_5288);
or UO_979 (O_979,N_6527,N_6157);
nor UO_980 (O_980,N_5700,N_6665);
or UO_981 (O_981,N_5750,N_5232);
xor UO_982 (O_982,N_5914,N_8426);
or UO_983 (O_983,N_6083,N_6093);
or UO_984 (O_984,N_7211,N_6586);
and UO_985 (O_985,N_8875,N_7240);
or UO_986 (O_986,N_6185,N_7734);
and UO_987 (O_987,N_5561,N_6776);
nand UO_988 (O_988,N_9514,N_8053);
or UO_989 (O_989,N_8109,N_8910);
nor UO_990 (O_990,N_6024,N_6743);
nor UO_991 (O_991,N_9312,N_6151);
nand UO_992 (O_992,N_7750,N_6752);
xnor UO_993 (O_993,N_9016,N_7650);
nand UO_994 (O_994,N_8121,N_9992);
and UO_995 (O_995,N_6036,N_7641);
and UO_996 (O_996,N_6251,N_8086);
nor UO_997 (O_997,N_7898,N_6750);
and UO_998 (O_998,N_5876,N_8340);
and UO_999 (O_999,N_7192,N_6589);
or UO_1000 (O_1000,N_7847,N_9534);
nand UO_1001 (O_1001,N_5776,N_9182);
or UO_1002 (O_1002,N_5737,N_7445);
nand UO_1003 (O_1003,N_7376,N_6231);
and UO_1004 (O_1004,N_7626,N_6310);
nand UO_1005 (O_1005,N_9053,N_8935);
nand UO_1006 (O_1006,N_8123,N_5816);
nand UO_1007 (O_1007,N_9102,N_8237);
xor UO_1008 (O_1008,N_8712,N_8812);
nor UO_1009 (O_1009,N_6515,N_6521);
and UO_1010 (O_1010,N_8280,N_8776);
nor UO_1011 (O_1011,N_6953,N_9015);
nor UO_1012 (O_1012,N_5522,N_7568);
nand UO_1013 (O_1013,N_5481,N_7474);
nand UO_1014 (O_1014,N_5507,N_8306);
nor UO_1015 (O_1015,N_8917,N_8661);
and UO_1016 (O_1016,N_9733,N_7962);
nand UO_1017 (O_1017,N_7119,N_9705);
xor UO_1018 (O_1018,N_8754,N_5959);
nor UO_1019 (O_1019,N_8985,N_9349);
and UO_1020 (O_1020,N_6235,N_8094);
or UO_1021 (O_1021,N_6429,N_6394);
nor UO_1022 (O_1022,N_7066,N_5363);
nand UO_1023 (O_1023,N_6305,N_8119);
nand UO_1024 (O_1024,N_7992,N_8578);
nor UO_1025 (O_1025,N_7528,N_9827);
xnor UO_1026 (O_1026,N_6420,N_6671);
and UO_1027 (O_1027,N_5041,N_9431);
and UO_1028 (O_1028,N_8976,N_5654);
and UO_1029 (O_1029,N_7081,N_8987);
nor UO_1030 (O_1030,N_7763,N_5048);
nand UO_1031 (O_1031,N_7574,N_9413);
or UO_1032 (O_1032,N_7340,N_8251);
nor UO_1033 (O_1033,N_9035,N_8923);
xnor UO_1034 (O_1034,N_7744,N_8244);
and UO_1035 (O_1035,N_6583,N_6592);
nand UO_1036 (O_1036,N_6144,N_5544);
xor UO_1037 (O_1037,N_8962,N_8745);
nor UO_1038 (O_1038,N_8781,N_8488);
nand UO_1039 (O_1039,N_8648,N_6289);
xor UO_1040 (O_1040,N_6106,N_8252);
nand UO_1041 (O_1041,N_6155,N_8945);
xor UO_1042 (O_1042,N_8794,N_9423);
nand UO_1043 (O_1043,N_9897,N_8483);
and UO_1044 (O_1044,N_8527,N_5768);
nor UO_1045 (O_1045,N_7635,N_7859);
nand UO_1046 (O_1046,N_8265,N_7931);
xor UO_1047 (O_1047,N_6438,N_7419);
xnor UO_1048 (O_1048,N_8595,N_8877);
nor UO_1049 (O_1049,N_9688,N_5253);
or UO_1050 (O_1050,N_7077,N_5988);
nor UO_1051 (O_1051,N_5967,N_5273);
or UO_1052 (O_1052,N_7382,N_5901);
or UO_1053 (O_1053,N_6961,N_5095);
nand UO_1054 (O_1054,N_5811,N_5518);
or UO_1055 (O_1055,N_7023,N_5594);
nor UO_1056 (O_1056,N_6033,N_6148);
or UO_1057 (O_1057,N_8147,N_8098);
nand UO_1058 (O_1058,N_8749,N_6461);
and UO_1059 (O_1059,N_5055,N_9311);
nor UO_1060 (O_1060,N_5777,N_5078);
xnor UO_1061 (O_1061,N_7193,N_8438);
nor UO_1062 (O_1062,N_5397,N_5448);
and UO_1063 (O_1063,N_7828,N_7499);
nor UO_1064 (O_1064,N_5445,N_6159);
nor UO_1065 (O_1065,N_6647,N_7434);
xnor UO_1066 (O_1066,N_7888,N_5541);
nand UO_1067 (O_1067,N_5617,N_7538);
or UO_1068 (O_1068,N_5292,N_7636);
nor UO_1069 (O_1069,N_6489,N_6452);
nor UO_1070 (O_1070,N_5384,N_7936);
and UO_1071 (O_1071,N_7817,N_8716);
and UO_1072 (O_1072,N_7362,N_9545);
nand UO_1073 (O_1073,N_5906,N_7815);
nand UO_1074 (O_1074,N_8289,N_6849);
nor UO_1075 (O_1075,N_5392,N_8860);
and UO_1076 (O_1076,N_7942,N_5960);
nor UO_1077 (O_1077,N_8777,N_9408);
xor UO_1078 (O_1078,N_5574,N_9962);
and UO_1079 (O_1079,N_6493,N_5222);
or UO_1080 (O_1080,N_9918,N_5084);
nor UO_1081 (O_1081,N_9625,N_9470);
and UO_1082 (O_1082,N_9260,N_7144);
and UO_1083 (O_1083,N_8372,N_5103);
and UO_1084 (O_1084,N_7771,N_5873);
or UO_1085 (O_1085,N_7549,N_6444);
or UO_1086 (O_1086,N_7028,N_8498);
nand UO_1087 (O_1087,N_7590,N_7778);
and UO_1088 (O_1088,N_9653,N_9375);
nor UO_1089 (O_1089,N_7589,N_7235);
and UO_1090 (O_1090,N_5698,N_9790);
nand UO_1091 (O_1091,N_5753,N_6211);
and UO_1092 (O_1092,N_5612,N_8737);
or UO_1093 (O_1093,N_8836,N_7733);
and UO_1094 (O_1094,N_9639,N_5282);
xor UO_1095 (O_1095,N_9804,N_9257);
nor UO_1096 (O_1096,N_6202,N_7363);
nand UO_1097 (O_1097,N_8942,N_9668);
nor UO_1098 (O_1098,N_7496,N_6535);
nand UO_1099 (O_1099,N_9141,N_6703);
and UO_1100 (O_1100,N_5254,N_5417);
nand UO_1101 (O_1101,N_6726,N_5586);
nor UO_1102 (O_1102,N_9709,N_6550);
nor UO_1103 (O_1103,N_5839,N_6579);
and UO_1104 (O_1104,N_9310,N_8394);
nor UO_1105 (O_1105,N_8898,N_8637);
or UO_1106 (O_1106,N_5034,N_9278);
nand UO_1107 (O_1107,N_9223,N_9676);
nor UO_1108 (O_1108,N_5323,N_6143);
xnor UO_1109 (O_1109,N_6679,N_6562);
and UO_1110 (O_1110,N_9772,N_8278);
xnor UO_1111 (O_1111,N_6801,N_9444);
nor UO_1112 (O_1112,N_5869,N_6694);
and UO_1113 (O_1113,N_5488,N_6266);
xor UO_1114 (O_1114,N_6850,N_7983);
or UO_1115 (O_1115,N_9195,N_6596);
xor UO_1116 (O_1116,N_6765,N_8321);
or UO_1117 (O_1117,N_6793,N_5240);
nor UO_1118 (O_1118,N_8433,N_6166);
xnor UO_1119 (O_1119,N_7749,N_5029);
nor UO_1120 (O_1120,N_5166,N_9582);
and UO_1121 (O_1121,N_7316,N_7344);
nand UO_1122 (O_1122,N_9635,N_6495);
and UO_1123 (O_1123,N_5133,N_7071);
nor UO_1124 (O_1124,N_5064,N_9627);
nor UO_1125 (O_1125,N_7911,N_6673);
xnor UO_1126 (O_1126,N_6469,N_5500);
nand UO_1127 (O_1127,N_8364,N_9228);
and UO_1128 (O_1128,N_7766,N_9414);
nand UO_1129 (O_1129,N_8678,N_9793);
xnor UO_1130 (O_1130,N_5357,N_9208);
and UO_1131 (O_1131,N_8242,N_9669);
nor UO_1132 (O_1132,N_6047,N_9092);
nand UO_1133 (O_1133,N_8254,N_9372);
nor UO_1134 (O_1134,N_6112,N_5699);
nand UO_1135 (O_1135,N_5480,N_9333);
nand UO_1136 (O_1136,N_5600,N_8886);
and UO_1137 (O_1137,N_9144,N_9120);
and UO_1138 (O_1138,N_7670,N_7552);
nor UO_1139 (O_1139,N_7645,N_5941);
nor UO_1140 (O_1140,N_7959,N_6767);
nand UO_1141 (O_1141,N_8971,N_9714);
or UO_1142 (O_1142,N_6524,N_6477);
and UO_1143 (O_1143,N_5465,N_8854);
or UO_1144 (O_1144,N_6049,N_5106);
or UO_1145 (O_1145,N_9134,N_9147);
and UO_1146 (O_1146,N_6379,N_9442);
and UO_1147 (O_1147,N_8083,N_8670);
and UO_1148 (O_1148,N_6825,N_9355);
or UO_1149 (O_1149,N_7961,N_5474);
and UO_1150 (O_1150,N_5102,N_7884);
xor UO_1151 (O_1151,N_5421,N_9307);
nor UO_1152 (O_1152,N_5441,N_6494);
or UO_1153 (O_1153,N_6340,N_7472);
nor UO_1154 (O_1154,N_8892,N_9390);
or UO_1155 (O_1155,N_7741,N_6021);
nand UO_1156 (O_1156,N_7775,N_5156);
nor UO_1157 (O_1157,N_7251,N_8246);
or UO_1158 (O_1158,N_5327,N_6081);
xor UO_1159 (O_1159,N_5473,N_6898);
nor UO_1160 (O_1160,N_9996,N_9747);
nor UO_1161 (O_1161,N_7000,N_5318);
and UO_1162 (O_1162,N_9115,N_6518);
and UO_1163 (O_1163,N_7440,N_7903);
and UO_1164 (O_1164,N_6435,N_8913);
nand UO_1165 (O_1165,N_9884,N_8271);
nor UO_1166 (O_1166,N_6110,N_5994);
and UO_1167 (O_1167,N_9287,N_9288);
or UO_1168 (O_1168,N_6785,N_5199);
or UO_1169 (O_1169,N_9322,N_9227);
nor UO_1170 (O_1170,N_7988,N_6139);
nor UO_1171 (O_1171,N_6872,N_7049);
or UO_1172 (O_1172,N_9283,N_5399);
and UO_1173 (O_1173,N_6109,N_5536);
or UO_1174 (O_1174,N_8508,N_5557);
nand UO_1175 (O_1175,N_6884,N_6079);
and UO_1176 (O_1176,N_7603,N_5368);
and UO_1177 (O_1177,N_9949,N_7215);
nor UO_1178 (O_1178,N_9291,N_8417);
or UO_1179 (O_1179,N_8801,N_8873);
nand UO_1180 (O_1180,N_8367,N_8931);
nand UO_1181 (O_1181,N_7660,N_9976);
nand UO_1182 (O_1182,N_8071,N_6312);
nor UO_1183 (O_1183,N_6321,N_5143);
and UO_1184 (O_1184,N_7558,N_5458);
and UO_1185 (O_1185,N_5274,N_6190);
and UO_1186 (O_1186,N_5946,N_5163);
or UO_1187 (O_1187,N_8828,N_7174);
nor UO_1188 (O_1188,N_5546,N_5814);
nand UO_1189 (O_1189,N_5188,N_6334);
nor UO_1190 (O_1190,N_6248,N_5415);
xor UO_1191 (O_1191,N_8613,N_6858);
nor UO_1192 (O_1192,N_8030,N_9456);
or UO_1193 (O_1193,N_5153,N_8825);
nand UO_1194 (O_1194,N_7943,N_8915);
or UO_1195 (O_1195,N_8529,N_5864);
or UO_1196 (O_1196,N_6674,N_7108);
nand UO_1197 (O_1197,N_7365,N_9395);
and UO_1198 (O_1198,N_6116,N_8100);
or UO_1199 (O_1199,N_7907,N_8811);
and UO_1200 (O_1200,N_8114,N_6637);
nor UO_1201 (O_1201,N_9091,N_9628);
and UO_1202 (O_1202,N_7715,N_9854);
and UO_1203 (O_1203,N_6046,N_8988);
and UO_1204 (O_1204,N_7114,N_9196);
nor UO_1205 (O_1205,N_6198,N_5969);
nand UO_1206 (O_1206,N_7638,N_8906);
nand UO_1207 (O_1207,N_7720,N_8681);
nor UO_1208 (O_1208,N_6655,N_6760);
nand UO_1209 (O_1209,N_9770,N_7789);
and UO_1210 (O_1210,N_7901,N_8768);
nand UO_1211 (O_1211,N_5916,N_9212);
nand UO_1212 (O_1212,N_8150,N_8516);
nand UO_1213 (O_1213,N_5210,N_5137);
xor UO_1214 (O_1214,N_8397,N_9131);
nor UO_1215 (O_1215,N_9626,N_7571);
or UO_1216 (O_1216,N_5042,N_8523);
and UO_1217 (O_1217,N_5671,N_6306);
xor UO_1218 (O_1218,N_6082,N_6345);
and UO_1219 (O_1219,N_6725,N_7133);
xnor UO_1220 (O_1220,N_9646,N_6580);
nand UO_1221 (O_1221,N_8383,N_6778);
or UO_1222 (O_1222,N_5414,N_7813);
xnor UO_1223 (O_1223,N_7615,N_7194);
nor UO_1224 (O_1224,N_9110,N_7649);
nand UO_1225 (O_1225,N_7100,N_7438);
and UO_1226 (O_1226,N_6275,N_7709);
nand UO_1227 (O_1227,N_9746,N_8660);
or UO_1228 (O_1228,N_6913,N_7864);
xnor UO_1229 (O_1229,N_9520,N_7468);
nand UO_1230 (O_1230,N_7139,N_7024);
or UO_1231 (O_1231,N_9979,N_5705);
nand UO_1232 (O_1232,N_9480,N_5905);
and UO_1233 (O_1233,N_6904,N_5047);
nor UO_1234 (O_1234,N_5115,N_5972);
nand UO_1235 (O_1235,N_6086,N_8762);
xor UO_1236 (O_1236,N_7639,N_7735);
nand UO_1237 (O_1237,N_8217,N_8604);
nor UO_1238 (O_1238,N_6845,N_8210);
or UO_1239 (O_1239,N_5100,N_7167);
or UO_1240 (O_1240,N_6060,N_8588);
nand UO_1241 (O_1241,N_5053,N_6430);
and UO_1242 (O_1242,N_6103,N_5808);
and UO_1243 (O_1243,N_7797,N_8556);
nand UO_1244 (O_1244,N_7260,N_5330);
and UO_1245 (O_1245,N_7896,N_6548);
and UO_1246 (O_1246,N_6573,N_7041);
nand UO_1247 (O_1247,N_6519,N_9614);
or UO_1248 (O_1248,N_7313,N_8126);
and UO_1249 (O_1249,N_9556,N_8267);
nor UO_1250 (O_1250,N_8182,N_5224);
or UO_1251 (O_1251,N_5885,N_6433);
xor UO_1252 (O_1252,N_8774,N_5749);
nand UO_1253 (O_1253,N_8544,N_8495);
or UO_1254 (O_1254,N_8605,N_8994);
xnor UO_1255 (O_1255,N_7270,N_5683);
or UO_1256 (O_1256,N_6585,N_5291);
or UO_1257 (O_1257,N_7091,N_6352);
or UO_1258 (O_1258,N_6854,N_9740);
and UO_1259 (O_1259,N_9701,N_5038);
nand UO_1260 (O_1260,N_5056,N_5932);
nand UO_1261 (O_1261,N_6547,N_7783);
or UO_1262 (O_1262,N_6989,N_8304);
nor UO_1263 (O_1263,N_6980,N_9913);
or UO_1264 (O_1264,N_7784,N_7845);
nor UO_1265 (O_1265,N_9453,N_6210);
and UO_1266 (O_1266,N_6706,N_9484);
xnor UO_1267 (O_1267,N_6301,N_7372);
xnor UO_1268 (O_1268,N_8617,N_7063);
and UO_1269 (O_1269,N_7600,N_6445);
nor UO_1270 (O_1270,N_5956,N_8079);
and UO_1271 (O_1271,N_5026,N_8133);
and UO_1272 (O_1272,N_9170,N_5244);
and UO_1273 (O_1273,N_5454,N_7653);
nor UO_1274 (O_1274,N_9367,N_5145);
nand UO_1275 (O_1275,N_6255,N_5528);
nand UO_1276 (O_1276,N_9836,N_8707);
nor UO_1277 (O_1277,N_5485,N_9847);
nand UO_1278 (O_1278,N_8720,N_8375);
or UO_1279 (O_1279,N_6893,N_9580);
or UO_1280 (O_1280,N_5589,N_7604);
xnor UO_1281 (O_1281,N_7047,N_5813);
xnor UO_1282 (O_1282,N_8149,N_7327);
nand UO_1283 (O_1283,N_7520,N_6607);
or UO_1284 (O_1284,N_8044,N_6724);
and UO_1285 (O_1285,N_6538,N_6273);
or UO_1286 (O_1286,N_9093,N_7940);
nand UO_1287 (O_1287,N_9497,N_7755);
nor UO_1288 (O_1288,N_5947,N_7886);
nand UO_1289 (O_1289,N_7669,N_7324);
and UO_1290 (O_1290,N_8693,N_9384);
or UO_1291 (O_1291,N_5173,N_6387);
or UO_1292 (O_1292,N_8859,N_5938);
or UO_1293 (O_1293,N_8355,N_5471);
or UO_1294 (O_1294,N_9075,N_6010);
nor UO_1295 (O_1295,N_5335,N_7697);
nand UO_1296 (O_1296,N_8338,N_9998);
nor UO_1297 (O_1297,N_7667,N_8029);
xor UO_1298 (O_1298,N_9088,N_7708);
xnor UO_1299 (O_1299,N_7078,N_9279);
xnor UO_1300 (O_1300,N_8479,N_8385);
and UO_1301 (O_1301,N_5223,N_5370);
xor UO_1302 (O_1302,N_9350,N_5829);
nor UO_1303 (O_1303,N_9618,N_7008);
xnor UO_1304 (O_1304,N_6330,N_5219);
xnor UO_1305 (O_1305,N_5127,N_9103);
and UO_1306 (O_1306,N_7467,N_7954);
and UO_1307 (O_1307,N_9068,N_5883);
nor UO_1308 (O_1308,N_5831,N_9681);
or UO_1309 (O_1309,N_9122,N_7458);
or UO_1310 (O_1310,N_7228,N_6191);
and UO_1311 (O_1311,N_8357,N_6653);
nand UO_1312 (O_1312,N_8566,N_9280);
nor UO_1313 (O_1313,N_5349,N_5981);
nor UO_1314 (O_1314,N_6971,N_5684);
nor UO_1315 (O_1315,N_6597,N_7625);
or UO_1316 (O_1316,N_7523,N_5762);
nand UO_1317 (O_1317,N_8228,N_7838);
nand UO_1318 (O_1318,N_6318,N_7136);
xor UO_1319 (O_1319,N_8802,N_9032);
nor UO_1320 (O_1320,N_5409,N_7356);
xnor UO_1321 (O_1321,N_6711,N_8554);
and UO_1322 (O_1322,N_7927,N_5886);
or UO_1323 (O_1323,N_9663,N_7367);
xor UO_1324 (O_1324,N_5179,N_7032);
nand UO_1325 (O_1325,N_7478,N_6987);
or UO_1326 (O_1326,N_6319,N_6781);
or UO_1327 (O_1327,N_5879,N_8272);
or UO_1328 (O_1328,N_9244,N_7951);
xor UO_1329 (O_1329,N_9766,N_9807);
or UO_1330 (O_1330,N_9155,N_8627);
nand UO_1331 (O_1331,N_8089,N_5924);
and UO_1332 (O_1332,N_7112,N_9658);
and UO_1333 (O_1333,N_6014,N_6366);
and UO_1334 (O_1334,N_5790,N_5401);
and UO_1335 (O_1335,N_6076,N_7009);
nand UO_1336 (O_1336,N_6338,N_8662);
or UO_1337 (O_1337,N_9236,N_9005);
nand UO_1338 (O_1338,N_9683,N_5696);
nand UO_1339 (O_1339,N_5195,N_8423);
or UO_1340 (O_1340,N_7195,N_9652);
or UO_1341 (O_1341,N_8422,N_5551);
or UO_1342 (O_1342,N_5247,N_5497);
nand UO_1343 (O_1343,N_7439,N_6934);
and UO_1344 (O_1344,N_8345,N_9040);
nand UO_1345 (O_1345,N_8609,N_5640);
or UO_1346 (O_1346,N_7374,N_6326);
nand UO_1347 (O_1347,N_5832,N_6095);
nor UO_1348 (O_1348,N_6242,N_5890);
or UO_1349 (O_1349,N_6184,N_7037);
nand UO_1350 (O_1350,N_8090,N_7507);
nor UO_1351 (O_1351,N_9022,N_5646);
nor UO_1352 (O_1352,N_8339,N_5320);
nor UO_1353 (O_1353,N_9399,N_7724);
nand UO_1354 (O_1354,N_9416,N_5793);
and UO_1355 (O_1355,N_5618,N_8589);
nand UO_1356 (O_1356,N_7822,N_8705);
nand UO_1357 (O_1357,N_7350,N_8619);
or UO_1358 (O_1358,N_8560,N_9610);
nand UO_1359 (O_1359,N_9318,N_6732);
xnor UO_1360 (O_1360,N_9773,N_7764);
and UO_1361 (O_1361,N_8337,N_6925);
nand UO_1362 (O_1362,N_8733,N_7384);
nor UO_1363 (O_1363,N_5105,N_8463);
xor UO_1364 (O_1364,N_8148,N_5125);
nand UO_1365 (O_1365,N_9339,N_6399);
xnor UO_1366 (O_1366,N_5146,N_8282);
or UO_1367 (O_1367,N_9270,N_9817);
or UO_1368 (O_1368,N_9871,N_5596);
nand UO_1369 (O_1369,N_9471,N_5661);
nor UO_1370 (O_1370,N_9211,N_7492);
nand UO_1371 (O_1371,N_9158,N_8080);
or UO_1372 (O_1372,N_7259,N_6028);
nand UO_1373 (O_1373,N_7025,N_9146);
and UO_1374 (O_1374,N_9991,N_9911);
nor UO_1375 (O_1375,N_6830,N_8396);
and UO_1376 (O_1376,N_6167,N_8624);
nand UO_1377 (O_1377,N_9326,N_5822);
xor UO_1378 (O_1378,N_9783,N_9238);
and UO_1379 (O_1379,N_7217,N_8069);
and UO_1380 (O_1380,N_7800,N_6959);
or UO_1381 (O_1381,N_6057,N_5849);
nor UO_1382 (O_1382,N_8950,N_7973);
or UO_1383 (O_1383,N_7782,N_8507);
nor UO_1384 (O_1384,N_8470,N_6807);
or UO_1385 (O_1385,N_6367,N_6025);
or UO_1386 (O_1386,N_5688,N_9491);
or UO_1387 (O_1387,N_7719,N_9543);
or UO_1388 (O_1388,N_9271,N_5169);
and UO_1389 (O_1389,N_6805,N_8113);
and UO_1390 (O_1390,N_8420,N_6005);
nand UO_1391 (O_1391,N_7821,N_6866);
nand UO_1392 (O_1392,N_6391,N_6918);
nor UO_1393 (O_1393,N_5246,N_8818);
xnor UO_1394 (O_1394,N_5233,N_5486);
and UO_1395 (O_1395,N_5888,N_9665);
or UO_1396 (O_1396,N_6669,N_5387);
nor UO_1397 (O_1397,N_7175,N_6729);
and UO_1398 (O_1398,N_7857,N_9425);
nand UO_1399 (O_1399,N_8806,N_6704);
nor UO_1400 (O_1400,N_5672,N_8311);
nand UO_1401 (O_1401,N_5452,N_6867);
nand UO_1402 (O_1402,N_9872,N_7695);
or UO_1403 (O_1403,N_7787,N_5571);
and UO_1404 (O_1404,N_8916,N_9748);
nand UO_1405 (O_1405,N_7664,N_6656);
nand UO_1406 (O_1406,N_6847,N_5774);
and UO_1407 (O_1407,N_8573,N_9750);
or UO_1408 (O_1408,N_8638,N_5008);
nand UO_1409 (O_1409,N_6274,N_7137);
nor UO_1410 (O_1410,N_6593,N_5925);
or UO_1411 (O_1411,N_5895,N_6205);
or UO_1412 (O_1412,N_6455,N_7377);
and UO_1413 (O_1413,N_9097,N_5201);
nor UO_1414 (O_1414,N_6240,N_6374);
nand UO_1415 (O_1415,N_5306,N_5675);
or UO_1416 (O_1416,N_9664,N_9327);
xor UO_1417 (O_1417,N_8330,N_8596);
and UO_1418 (O_1418,N_5385,N_5833);
nor UO_1419 (O_1419,N_5431,N_6048);
and UO_1420 (O_1420,N_7867,N_6283);
nor UO_1421 (O_1421,N_6359,N_7311);
nand UO_1422 (O_1422,N_6054,N_8288);
nor UO_1423 (O_1423,N_6624,N_7135);
or UO_1424 (O_1424,N_5697,N_9978);
or UO_1425 (O_1425,N_9672,N_7339);
or UO_1426 (O_1426,N_9010,N_7205);
xor UO_1427 (O_1427,N_7677,N_7505);
nand UO_1428 (O_1428,N_5178,N_5695);
nand UO_1429 (O_1429,N_9813,N_7412);
nor UO_1430 (O_1430,N_7030,N_5512);
nor UO_1431 (O_1431,N_5031,N_7788);
nor UO_1432 (O_1432,N_8684,N_9296);
nor UO_1433 (O_1433,N_6250,N_9671);
nand UO_1434 (O_1434,N_7354,N_6610);
nand UO_1435 (O_1435,N_8294,N_7661);
nand UO_1436 (O_1436,N_7672,N_6705);
nor UO_1437 (O_1437,N_8212,N_5782);
or UO_1438 (O_1438,N_7585,N_9047);
or UO_1439 (O_1439,N_9554,N_9855);
and UO_1440 (O_1440,N_8827,N_7065);
nand UO_1441 (O_1441,N_8425,N_6253);
nor UO_1442 (O_1442,N_7358,N_5861);
or UO_1443 (O_1443,N_9014,N_5992);
or UO_1444 (O_1444,N_6853,N_6336);
and UO_1445 (O_1445,N_7900,N_8170);
or UO_1446 (O_1446,N_8183,N_7088);
nand UO_1447 (O_1447,N_5072,N_9691);
nor UO_1448 (O_1448,N_7700,N_6315);
and UO_1449 (O_1449,N_6672,N_9712);
nor UO_1450 (O_1450,N_8365,N_6453);
nand UO_1451 (O_1451,N_9771,N_5236);
nor UO_1452 (O_1452,N_7557,N_8558);
nand UO_1453 (O_1453,N_9630,N_6628);
and UO_1454 (O_1454,N_9852,N_5418);
or UO_1455 (O_1455,N_7333,N_7564);
xor UO_1456 (O_1456,N_9401,N_9695);
xor UO_1457 (O_1457,N_9661,N_7950);
xor UO_1458 (O_1458,N_6209,N_9839);
nor UO_1459 (O_1459,N_6857,N_5927);
nor UO_1460 (O_1460,N_5882,N_7398);
or UO_1461 (O_1461,N_7785,N_8348);
nor UO_1462 (O_1462,N_5360,N_5001);
xor UO_1463 (O_1463,N_9361,N_9504);
nor UO_1464 (O_1464,N_9525,N_8196);
nand UO_1465 (O_1465,N_6540,N_9586);
nand UO_1466 (O_1466,N_8732,N_9863);
or UO_1467 (O_1467,N_8072,N_9069);
or UO_1468 (O_1468,N_9987,N_6763);
nand UO_1469 (O_1469,N_8711,N_5757);
and UO_1470 (O_1470,N_7330,N_5944);
nand UO_1471 (O_1471,N_6241,N_7702);
nand UO_1472 (O_1472,N_7502,N_9735);
nand UO_1473 (O_1473,N_7447,N_9157);
or UO_1474 (O_1474,N_5840,N_7224);
xnor UO_1475 (O_1475,N_7241,N_6874);
and UO_1476 (O_1476,N_5248,N_7157);
nor UO_1477 (O_1477,N_7456,N_6053);
and UO_1478 (O_1478,N_6731,N_9659);
nor UO_1479 (O_1479,N_8052,N_9421);
nand UO_1480 (O_1480,N_5442,N_7057);
nor UO_1481 (O_1481,N_6813,N_7924);
nand UO_1482 (O_1482,N_9254,N_9086);
nand UO_1483 (O_1483,N_8106,N_9690);
nand UO_1484 (O_1484,N_8645,N_7792);
nand UO_1485 (O_1485,N_7563,N_8499);
nand UO_1486 (O_1486,N_5174,N_6506);
xor UO_1487 (O_1487,N_8763,N_8780);
xnor UO_1488 (O_1488,N_8791,N_6920);
xnor UO_1489 (O_1489,N_6829,N_5641);
nor UO_1490 (O_1490,N_9418,N_5311);
and UO_1491 (O_1491,N_9541,N_7378);
nand UO_1492 (O_1492,N_8378,N_9379);
or UO_1493 (O_1493,N_8944,N_6569);
nand UO_1494 (O_1494,N_9600,N_6839);
or UO_1495 (O_1495,N_6392,N_8909);
nor UO_1496 (O_1496,N_7690,N_5539);
and UO_1497 (O_1497,N_5681,N_7995);
and UO_1498 (O_1498,N_7540,N_6852);
nor UO_1499 (O_1499,N_9026,N_7874);
endmodule