module basic_1500_15000_2000_20_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_886,In_246);
nand U1 (N_1,In_919,In_365);
nand U2 (N_2,In_1314,In_601);
xor U3 (N_3,In_1172,In_1098);
and U4 (N_4,In_540,In_1190);
nor U5 (N_5,In_294,In_362);
xnor U6 (N_6,In_762,In_1400);
nand U7 (N_7,In_605,In_580);
or U8 (N_8,In_532,In_1008);
and U9 (N_9,In_1263,In_41);
nor U10 (N_10,In_1403,In_198);
nand U11 (N_11,In_591,In_479);
and U12 (N_12,In_992,In_117);
or U13 (N_13,In_91,In_1175);
nor U14 (N_14,In_779,In_135);
nor U15 (N_15,In_1137,In_386);
and U16 (N_16,In_775,In_471);
xor U17 (N_17,In_1473,In_678);
nor U18 (N_18,In_217,In_255);
xor U19 (N_19,In_381,In_965);
xor U20 (N_20,In_895,In_936);
xor U21 (N_21,In_1277,In_885);
nand U22 (N_22,In_1496,In_1162);
xnor U23 (N_23,In_538,In_777);
nand U24 (N_24,In_1282,In_660);
or U25 (N_25,In_124,In_745);
and U26 (N_26,In_1124,In_1227);
and U27 (N_27,In_1458,In_707);
or U28 (N_28,In_69,In_1006);
or U29 (N_29,In_1122,In_1086);
nand U30 (N_30,In_59,In_593);
and U31 (N_31,In_407,In_1468);
and U32 (N_32,In_1389,In_93);
xnor U33 (N_33,In_1102,In_307);
nor U34 (N_34,In_419,In_872);
nor U35 (N_35,In_1344,In_331);
nand U36 (N_36,In_611,In_652);
nand U37 (N_37,In_349,In_1460);
nor U38 (N_38,In_1335,In_796);
xnor U39 (N_39,In_154,In_1211);
or U40 (N_40,In_68,In_1372);
xnor U41 (N_41,In_159,In_803);
xnor U42 (N_42,In_1443,In_1163);
nor U43 (N_43,In_1101,In_1244);
xor U44 (N_44,In_375,In_1093);
or U45 (N_45,In_145,In_764);
xnor U46 (N_46,In_379,In_941);
or U47 (N_47,In_1380,In_814);
or U48 (N_48,In_1415,In_85);
and U49 (N_49,In_212,In_1146);
and U50 (N_50,In_837,In_1136);
xor U51 (N_51,In_256,In_168);
and U52 (N_52,In_845,In_202);
or U53 (N_53,In_735,In_710);
xor U54 (N_54,In_647,In_1209);
or U55 (N_55,In_499,In_692);
xnor U56 (N_56,In_480,In_914);
nand U57 (N_57,In_295,In_865);
nand U58 (N_58,In_498,In_950);
nor U59 (N_59,In_1355,In_1265);
xnor U60 (N_60,In_976,In_98);
nor U61 (N_61,In_995,In_1082);
nand U62 (N_62,In_747,In_1268);
and U63 (N_63,In_638,In_902);
or U64 (N_64,In_1429,In_358);
nand U65 (N_65,In_208,In_94);
nor U66 (N_66,In_830,In_959);
or U67 (N_67,In_1378,In_999);
nor U68 (N_68,In_292,In_1187);
nand U69 (N_69,In_1181,In_937);
and U70 (N_70,In_700,In_1345);
nor U71 (N_71,In_33,In_1143);
nand U72 (N_72,In_756,In_1352);
or U73 (N_73,In_1305,In_1308);
or U74 (N_74,In_447,In_812);
xnor U75 (N_75,In_786,In_718);
xnor U76 (N_76,In_582,In_1410);
xnor U77 (N_77,In_1159,In_542);
or U78 (N_78,In_1363,In_674);
nand U79 (N_79,In_1270,In_1393);
nor U80 (N_80,In_685,In_146);
nand U81 (N_81,In_951,In_699);
xnor U82 (N_82,In_1408,In_221);
and U83 (N_83,In_541,In_403);
nand U84 (N_84,In_1022,In_1317);
or U85 (N_85,In_1100,In_196);
or U86 (N_86,In_1286,In_1201);
xnor U87 (N_87,In_1271,In_414);
or U88 (N_88,In_1302,In_1319);
and U89 (N_89,In_84,In_86);
nor U90 (N_90,In_251,In_826);
nor U91 (N_91,In_1450,In_383);
xnor U92 (N_92,In_957,In_904);
xnor U93 (N_93,In_485,In_1068);
nor U94 (N_94,In_555,In_483);
xnor U95 (N_95,In_486,In_352);
and U96 (N_96,In_460,In_335);
nand U97 (N_97,In_793,In_1440);
nor U98 (N_98,In_750,In_179);
and U99 (N_99,In_426,In_1366);
xnor U100 (N_100,In_56,In_846);
nor U101 (N_101,In_417,In_1276);
nand U102 (N_102,In_1016,In_1248);
and U103 (N_103,In_204,In_63);
and U104 (N_104,In_943,In_308);
or U105 (N_105,In_406,In_1413);
nor U106 (N_106,In_437,In_1471);
nor U107 (N_107,In_266,In_1260);
or U108 (N_108,In_157,In_971);
or U109 (N_109,In_1310,In_1139);
or U110 (N_110,In_393,In_1485);
or U111 (N_111,In_50,In_724);
and U112 (N_112,In_521,In_1338);
nand U113 (N_113,In_1430,In_1166);
nand U114 (N_114,In_224,In_115);
or U115 (N_115,In_1035,In_96);
xnor U116 (N_116,In_972,In_1199);
or U117 (N_117,In_1313,In_215);
xnor U118 (N_118,In_634,In_899);
and U119 (N_119,In_1032,In_684);
or U120 (N_120,In_702,In_596);
nor U121 (N_121,In_942,In_740);
and U122 (N_122,In_148,In_276);
nor U123 (N_123,In_1452,In_657);
nand U124 (N_124,In_495,In_164);
nand U125 (N_125,In_935,In_161);
and U126 (N_126,In_840,In_90);
nor U127 (N_127,In_1092,In_1229);
nand U128 (N_128,In_565,In_676);
nand U129 (N_129,In_366,In_852);
nor U130 (N_130,In_420,In_597);
nor U131 (N_131,In_245,In_488);
nand U132 (N_132,In_1288,In_1097);
nor U133 (N_133,In_968,In_277);
nand U134 (N_134,In_1048,In_1295);
xnor U135 (N_135,In_927,In_434);
nor U136 (N_136,In_780,In_169);
or U137 (N_137,In_66,In_1438);
nand U138 (N_138,In_1498,In_165);
or U139 (N_139,In_956,In_1034);
xor U140 (N_140,In_1499,In_810);
or U141 (N_141,In_1251,In_1356);
or U142 (N_142,In_126,In_454);
nor U143 (N_143,In_1367,In_633);
and U144 (N_144,In_642,In_1129);
nor U145 (N_145,In_549,In_932);
or U146 (N_146,In_921,In_288);
nand U147 (N_147,In_1434,In_961);
nor U148 (N_148,In_506,In_432);
nand U149 (N_149,In_416,In_566);
nand U150 (N_150,In_1484,In_1466);
xor U151 (N_151,In_109,In_1018);
nor U152 (N_152,In_1328,In_749);
xnor U153 (N_153,In_1495,In_1297);
nand U154 (N_154,In_1259,In_817);
nor U155 (N_155,In_1064,In_618);
and U156 (N_156,In_1174,In_278);
nor U157 (N_157,In_931,In_1170);
and U158 (N_158,In_274,In_818);
xor U159 (N_159,In_797,In_873);
xnor U160 (N_160,In_1158,In_834);
or U161 (N_161,In_329,In_1448);
nand U162 (N_162,In_934,In_828);
or U163 (N_163,In_1472,In_283);
nor U164 (N_164,In_82,In_909);
or U165 (N_165,In_782,In_1108);
xor U166 (N_166,In_1379,In_727);
nor U167 (N_167,In_127,In_472);
or U168 (N_168,In_1368,In_1349);
nor U169 (N_169,In_44,In_205);
xnor U170 (N_170,In_848,In_1353);
or U171 (N_171,In_1283,In_649);
nor U172 (N_172,In_16,In_241);
nor U173 (N_173,In_1059,In_24);
xnor U174 (N_174,In_1447,In_286);
and U175 (N_175,In_10,In_871);
and U176 (N_176,In_265,In_481);
or U177 (N_177,In_639,In_564);
or U178 (N_178,In_1463,In_658);
nor U179 (N_179,In_854,In_705);
nor U180 (N_180,In_1052,In_102);
or U181 (N_181,In_856,In_673);
or U182 (N_182,In_150,In_1090);
or U183 (N_183,In_51,In_1207);
and U184 (N_184,In_1320,In_1334);
or U185 (N_185,In_588,In_509);
nand U186 (N_186,In_1073,In_248);
nand U187 (N_187,In_262,In_1128);
xnor U188 (N_188,In_821,In_1331);
nand U189 (N_189,In_1192,In_79);
nor U190 (N_190,In_34,In_39);
nor U191 (N_191,In_1116,In_332);
xor U192 (N_192,In_516,In_133);
xnor U193 (N_193,In_617,In_436);
xnor U194 (N_194,In_1401,In_418);
or U195 (N_195,In_189,In_1074);
xnor U196 (N_196,In_963,In_1218);
nand U197 (N_197,In_1405,In_773);
xnor U198 (N_198,In_1036,In_178);
xnor U199 (N_199,In_1258,In_1444);
nand U200 (N_200,In_125,In_608);
xnor U201 (N_201,In_389,In_1112);
nor U202 (N_202,In_667,In_97);
nor U203 (N_203,In_484,In_551);
nand U204 (N_204,In_1493,In_1080);
nand U205 (N_205,In_546,In_670);
nand U206 (N_206,In_567,In_788);
nand U207 (N_207,In_827,In_759);
nand U208 (N_208,In_574,In_839);
and U209 (N_209,In_1113,In_1414);
and U210 (N_210,In_443,In_257);
xnor U211 (N_211,In_725,In_328);
nand U212 (N_212,In_1228,In_1252);
nand U213 (N_213,In_207,In_402);
nand U214 (N_214,In_1233,In_132);
nor U215 (N_215,In_1156,In_514);
xor U216 (N_216,In_815,In_1070);
and U217 (N_217,In_975,In_1195);
nand U218 (N_218,In_809,In_798);
nand U219 (N_219,In_1294,In_1041);
nand U220 (N_220,In_1083,In_232);
or U221 (N_221,In_1293,In_1107);
nand U222 (N_222,In_804,In_890);
xor U223 (N_223,In_138,In_1423);
xor U224 (N_224,In_147,In_691);
and U225 (N_225,In_905,In_1173);
and U226 (N_226,In_29,In_630);
and U227 (N_227,In_5,In_825);
xor U228 (N_228,In_625,In_847);
nand U229 (N_229,In_831,In_915);
nor U230 (N_230,In_330,In_833);
nor U231 (N_231,In_261,In_510);
or U232 (N_232,In_734,In_1391);
nor U233 (N_233,In_568,In_1455);
and U234 (N_234,In_421,In_1341);
xor U235 (N_235,In_1402,In_71);
or U236 (N_236,In_345,In_1135);
and U237 (N_237,In_1103,In_160);
and U238 (N_238,In_761,In_1386);
nand U239 (N_239,In_1232,In_758);
or U240 (N_240,In_722,In_322);
or U241 (N_241,In_1011,In_1240);
nor U242 (N_242,In_340,In_163);
nor U243 (N_243,In_615,In_43);
or U244 (N_244,In_237,In_518);
and U245 (N_245,In_622,In_1001);
nor U246 (N_246,In_808,In_477);
and U247 (N_247,In_993,In_412);
or U248 (N_248,In_629,In_739);
or U249 (N_249,In_1039,In_1104);
and U250 (N_250,In_428,In_190);
xor U251 (N_251,In_321,In_1406);
nand U252 (N_252,In_348,In_226);
nand U253 (N_253,In_171,In_153);
nor U254 (N_254,In_874,In_1065);
and U255 (N_255,In_341,In_800);
nor U256 (N_256,In_113,In_369);
nor U257 (N_257,In_1223,In_628);
nand U258 (N_258,In_1214,In_632);
nand U259 (N_259,In_285,In_859);
or U260 (N_260,In_1058,In_1189);
and U261 (N_261,In_181,In_698);
xor U262 (N_262,In_1024,In_1118);
xnor U263 (N_263,In_423,In_1084);
nor U264 (N_264,In_1177,In_1028);
or U265 (N_265,In_570,In_250);
or U266 (N_266,In_534,In_714);
xor U267 (N_267,In_731,In_1131);
nor U268 (N_268,In_881,In_1327);
and U269 (N_269,In_989,In_1225);
or U270 (N_270,In_879,In_1387);
or U271 (N_271,In_768,In_575);
nand U272 (N_272,In_716,In_1075);
nor U273 (N_273,In_167,In_1081);
nand U274 (N_274,In_1106,In_1040);
nor U275 (N_275,In_451,In_501);
nor U276 (N_276,In_519,In_377);
nor U277 (N_277,In_1152,In_966);
or U278 (N_278,In_1219,In_526);
and U279 (N_279,In_216,In_563);
nand U280 (N_280,In_336,In_1196);
xnor U281 (N_281,In_1224,In_515);
nor U282 (N_282,In_911,In_755);
and U283 (N_283,In_695,In_1442);
nand U284 (N_284,In_560,In_721);
xnor U285 (N_285,In_228,In_4);
nand U286 (N_286,In_67,In_141);
or U287 (N_287,In_372,In_924);
nand U288 (N_288,In_1148,In_304);
or U289 (N_289,In_58,In_864);
xor U290 (N_290,In_333,In_766);
xnor U291 (N_291,In_1306,In_589);
or U292 (N_292,In_405,In_547);
nor U293 (N_293,In_291,In_18);
nand U294 (N_294,In_343,In_1150);
nor U295 (N_295,In_267,In_457);
and U296 (N_296,In_603,In_1347);
and U297 (N_297,In_1004,In_119);
nor U298 (N_298,In_1066,In_1247);
and U299 (N_299,In_281,In_155);
or U300 (N_300,In_12,In_1115);
nand U301 (N_301,In_88,In_693);
or U302 (N_302,In_1357,In_548);
or U303 (N_303,In_537,In_1492);
or U304 (N_304,In_680,In_1254);
nand U305 (N_305,In_819,In_77);
and U306 (N_306,In_1337,In_577);
xnor U307 (N_307,In_1125,In_974);
and U308 (N_308,In_867,In_980);
xor U309 (N_309,In_361,In_1375);
or U310 (N_310,In_287,In_1340);
and U311 (N_311,In_1279,In_30);
xnor U312 (N_312,In_1291,In_607);
or U313 (N_313,In_1369,In_7);
or U314 (N_314,In_176,In_1117);
xor U315 (N_315,In_390,In_75);
and U316 (N_316,In_1256,In_813);
nor U317 (N_317,In_524,In_0);
nor U318 (N_318,In_991,In_1044);
or U319 (N_319,In_1309,In_1287);
nor U320 (N_320,In_600,In_1494);
and U321 (N_321,In_1222,In_1350);
xor U322 (N_322,In_1383,In_843);
and U323 (N_323,In_757,In_87);
nor U324 (N_324,In_891,In_23);
or U325 (N_325,In_60,In_954);
nor U326 (N_326,In_592,In_1395);
xor U327 (N_327,In_1020,In_763);
nand U328 (N_328,In_602,In_970);
nor U329 (N_329,In_1269,In_289);
or U330 (N_330,In_967,In_1290);
and U331 (N_331,In_121,In_1374);
xnor U332 (N_332,In_236,In_354);
or U333 (N_333,In_945,In_829);
xnor U334 (N_334,In_263,In_1210);
nor U335 (N_335,In_732,In_987);
nand U336 (N_336,In_496,In_1339);
or U337 (N_337,In_952,In_1437);
and U338 (N_338,In_318,In_370);
xor U339 (N_339,In_453,In_535);
and U340 (N_340,In_1456,In_284);
and U341 (N_341,In_184,In_270);
and U342 (N_342,In_877,In_475);
nor U343 (N_343,In_238,In_1243);
and U344 (N_344,In_408,In_1274);
or U345 (N_345,In_411,In_1280);
xor U346 (N_346,In_1149,In_449);
nand U347 (N_347,In_1482,In_1457);
nor U348 (N_348,In_222,In_641);
nor U349 (N_349,In_556,In_253);
or U350 (N_350,In_820,In_1109);
or U351 (N_351,In_173,In_1031);
and U352 (N_352,In_778,In_824);
xor U353 (N_353,In_492,In_1422);
nand U354 (N_354,In_861,In_1479);
and U355 (N_355,In_137,In_717);
or U356 (N_356,In_197,In_209);
xor U357 (N_357,In_394,In_712);
or U358 (N_358,In_371,In_1428);
nand U359 (N_359,In_823,In_720);
nand U360 (N_360,In_1216,In_1478);
xnor U361 (N_361,In_938,In_1105);
nand U362 (N_362,In_579,In_726);
nor U363 (N_363,In_1354,In_903);
or U364 (N_364,In_1300,In_889);
and U365 (N_365,In_646,In_269);
or U366 (N_366,In_80,In_162);
or U367 (N_367,In_2,In_464);
nand U368 (N_368,In_1246,In_953);
or U369 (N_369,In_1026,In_787);
nand U370 (N_370,In_690,In_1407);
nand U371 (N_371,In_1316,In_1132);
or U372 (N_372,In_22,In_404);
and U373 (N_373,In_1469,In_438);
nor U374 (N_374,In_1394,In_401);
or U375 (N_375,In_1062,In_998);
or U376 (N_376,In_1061,In_1332);
nor U377 (N_377,In_20,In_252);
nor U378 (N_378,In_1095,In_870);
and U379 (N_379,In_118,In_35);
or U380 (N_380,In_1373,In_737);
xor U381 (N_381,In_1441,In_853);
nor U382 (N_382,In_1009,In_884);
xor U383 (N_383,In_268,In_363);
xnor U384 (N_384,In_573,In_367);
xor U385 (N_385,In_397,In_784);
or U386 (N_386,In_857,In_595);
nor U387 (N_387,In_324,In_1182);
xor U388 (N_388,In_156,In_1346);
xor U389 (N_389,In_384,In_355);
nand U390 (N_390,In_1250,In_186);
or U391 (N_391,In_1436,In_765);
nand U392 (N_392,In_719,In_648);
or U393 (N_393,In_612,In_1432);
nor U394 (N_394,In_892,In_444);
or U395 (N_395,In_467,In_296);
and U396 (N_396,In_666,In_374);
nand U397 (N_397,In_940,In_1416);
or U398 (N_398,In_45,In_323);
nor U399 (N_399,In_604,In_503);
and U400 (N_400,In_247,In_424);
nand U401 (N_401,In_616,In_982);
and U402 (N_402,In_1141,In_400);
and U403 (N_403,In_1161,In_385);
nor U404 (N_404,In_1446,In_53);
nand U405 (N_405,In_131,In_623);
or U406 (N_406,In_668,In_1289);
nand U407 (N_407,In_581,In_1358);
nor U408 (N_408,In_104,In_1176);
nand U409 (N_409,In_1202,In_123);
and U410 (N_410,In_1043,In_836);
or U411 (N_411,In_599,In_225);
xor U412 (N_412,In_913,In_327);
nor U413 (N_413,In_711,In_880);
and U414 (N_414,In_832,In_1164);
nand U415 (N_415,In_175,In_1480);
or U416 (N_416,In_1003,In_1325);
nand U417 (N_417,In_11,In_427);
or U418 (N_418,In_410,In_1002);
nand U419 (N_419,In_511,In_949);
nand U420 (N_420,In_789,In_624);
xnor U421 (N_421,In_380,In_469);
nor U422 (N_422,In_1063,In_1120);
xor U423 (N_423,In_1488,In_440);
or U424 (N_424,In_578,In_230);
xor U425 (N_425,In_585,In_1239);
nand U426 (N_426,In_134,In_42);
xnor U427 (N_427,In_979,In_1160);
or U428 (N_428,In_1281,In_468);
xnor U429 (N_429,In_1390,In_741);
and U430 (N_430,In_746,In_1014);
nor U431 (N_431,In_898,In_754);
nor U432 (N_432,In_1023,In_130);
nor U433 (N_433,In_470,In_1411);
nand U434 (N_434,In_1015,In_1396);
and U435 (N_435,In_74,In_413);
xor U436 (N_436,In_116,In_507);
or U437 (N_437,In_785,In_76);
xnor U438 (N_438,In_1491,In_517);
xnor U439 (N_439,In_458,In_696);
and U440 (N_440,In_528,In_1094);
nor U441 (N_441,In_679,In_26);
nand U442 (N_442,In_728,In_1114);
or U443 (N_443,In_1205,In_910);
nor U444 (N_444,In_311,In_918);
nand U445 (N_445,In_305,In_1005);
nor U446 (N_446,In_1307,In_107);
xnor U447 (N_447,In_1235,In_213);
nand U448 (N_448,In_770,In_89);
nor U449 (N_449,In_1010,In_206);
nand U450 (N_450,In_1180,In_996);
nor U451 (N_451,In_522,In_504);
and U452 (N_452,In_558,In_536);
and U453 (N_453,In_1236,In_378);
nor U454 (N_454,In_733,In_1133);
xnor U455 (N_455,In_994,In_342);
and U456 (N_456,In_31,In_704);
xor U457 (N_457,In_1111,In_933);
nand U458 (N_458,In_1257,In_64);
and U459 (N_459,In_461,In_357);
xnor U460 (N_460,In_1025,In_1377);
nand U461 (N_461,In_1315,In_431);
nand U462 (N_462,In_923,In_1019);
and U463 (N_463,In_1056,In_571);
or U464 (N_464,In_822,In_106);
nand U465 (N_465,In_955,In_1203);
nor U466 (N_466,In_1330,In_1454);
nand U467 (N_467,In_100,In_806);
nand U468 (N_468,In_306,In_319);
nor U469 (N_469,In_663,In_944);
nand U470 (N_470,In_95,In_613);
nand U471 (N_471,In_52,In_1483);
and U472 (N_472,In_1194,In_751);
or U473 (N_473,In_36,In_1419);
xnor U474 (N_474,In_1096,In_191);
or U475 (N_475,In_631,In_356);
xor U476 (N_476,In_152,In_1237);
nor U477 (N_477,In_653,In_1130);
nand U478 (N_478,In_491,In_1050);
nor U479 (N_479,In_774,In_260);
nor U480 (N_480,In_1329,In_701);
nor U481 (N_481,In_120,In_767);
or U482 (N_482,In_300,In_863);
nand U483 (N_483,In_723,In_303);
xnor U484 (N_484,In_1140,In_1459);
nand U485 (N_485,In_1230,In_513);
xnor U486 (N_486,In_1200,In_455);
xnor U487 (N_487,In_738,In_878);
nand U488 (N_488,In_271,In_1445);
or U489 (N_489,In_841,In_561);
and U490 (N_490,In_1266,In_1012);
or U491 (N_491,In_533,In_272);
nand U492 (N_492,In_706,In_664);
and U493 (N_493,In_866,In_298);
or U494 (N_494,In_1435,In_344);
or U495 (N_495,In_450,In_1088);
xnor U496 (N_496,In_1360,In_211);
or U497 (N_497,In_1119,In_81);
nor U498 (N_498,In_1241,In_697);
xnor U499 (N_499,In_1217,In_531);
and U500 (N_500,In_1326,In_376);
and U501 (N_501,In_544,In_456);
nand U502 (N_502,In_1204,In_883);
nor U503 (N_503,In_838,In_49);
nand U504 (N_504,In_258,In_473);
nand U505 (N_505,In_487,In_550);
nor U506 (N_506,In_771,In_908);
nor U507 (N_507,In_1489,In_1299);
nand U508 (N_508,In_1198,In_855);
nand U509 (N_509,In_235,In_729);
and U510 (N_510,In_662,In_1231);
nand U511 (N_511,In_493,In_654);
and U512 (N_512,In_844,In_1371);
or U513 (N_513,In_129,In_614);
nor U514 (N_514,In_743,In_1151);
nor U515 (N_515,In_435,In_439);
nand U516 (N_516,In_143,In_1476);
and U517 (N_517,In_1186,In_1053);
nand U518 (N_518,In_83,In_1212);
and U519 (N_519,In_875,In_1486);
xnor U520 (N_520,In_985,In_1067);
nand U521 (N_521,In_792,In_665);
xor U522 (N_522,In_490,In_1385);
or U523 (N_523,In_17,In_234);
xor U524 (N_524,In_359,In_425);
nor U525 (N_525,In_1215,In_1462);
or U526 (N_526,In_1197,In_1123);
xnor U527 (N_527,In_112,In_474);
nand U528 (N_528,In_110,In_218);
nor U529 (N_529,In_219,In_229);
xor U530 (N_530,In_1049,In_930);
or U531 (N_531,In_1298,In_1311);
xnor U532 (N_532,In_1046,In_317);
nand U533 (N_533,In_947,In_199);
xor U534 (N_534,In_520,In_708);
xor U535 (N_535,In_543,In_187);
nand U536 (N_536,In_21,In_13);
or U537 (N_537,In_1168,In_48);
nor U538 (N_538,In_897,In_610);
and U539 (N_539,In_958,In_1421);
nor U540 (N_540,In_185,In_1348);
xor U541 (N_541,In_1333,In_791);
or U542 (N_542,In_587,In_1370);
or U543 (N_543,In_203,In_606);
nand U544 (N_544,In_494,In_776);
xor U545 (N_545,In_32,In_61);
and U546 (N_546,In_772,In_1398);
and U547 (N_547,In_273,In_635);
and U548 (N_548,In_790,In_1425);
xnor U549 (N_549,In_1155,In_802);
nand U550 (N_550,In_1312,In_105);
xor U551 (N_551,In_1321,In_1253);
xnor U552 (N_552,In_1076,In_27);
and U553 (N_553,In_1138,In_282);
nand U554 (N_554,In_65,In_1077);
nor U555 (N_555,In_876,In_835);
or U556 (N_556,In_244,In_46);
nor U557 (N_557,In_849,In_136);
or U558 (N_558,In_1206,In_525);
nand U559 (N_559,In_887,In_1284);
xor U560 (N_560,In_816,In_429);
or U561 (N_561,In_553,In_1275);
or U562 (N_562,In_860,In_960);
nor U563 (N_563,In_922,In_313);
and U564 (N_564,In_1126,In_687);
or U565 (N_565,In_851,In_382);
nor U566 (N_566,In_512,In_301);
xor U567 (N_567,In_681,In_103);
xor U568 (N_568,In_1365,In_325);
and U569 (N_569,In_1296,In_346);
or U570 (N_570,In_445,In_730);
and U571 (N_571,In_671,In_900);
nor U572 (N_572,In_783,In_360);
and U573 (N_573,In_715,In_290);
nor U574 (N_574,In_1071,In_586);
nor U575 (N_575,In_174,In_858);
or U576 (N_576,In_626,In_441);
xor U577 (N_577,In_1134,In_1060);
nor U578 (N_578,In_465,In_1343);
xor U579 (N_579,In_299,In_1021);
nor U580 (N_580,In_214,In_142);
nor U581 (N_581,In_1145,In_326);
or U582 (N_582,In_675,In_1409);
nand U583 (N_583,In_1245,In_552);
and U584 (N_584,In_1388,In_1467);
xor U585 (N_585,In_523,In_459);
xor U586 (N_586,In_170,In_108);
or U587 (N_587,In_1382,In_478);
nand U588 (N_588,In_280,In_279);
nand U589 (N_589,In_1418,In_907);
nor U590 (N_590,In_144,In_231);
nand U591 (N_591,In_920,In_57);
and U592 (N_592,In_1262,In_896);
xnor U593 (N_593,In_557,In_906);
and U594 (N_594,In_1007,In_1242);
and U595 (N_595,In_1381,In_54);
nand U596 (N_596,In_1042,In_1465);
xor U597 (N_597,In_929,In_677);
nor U598 (N_598,In_1420,In_339);
xor U599 (N_599,In_569,In_1361);
nor U600 (N_600,In_925,In_193);
and U601 (N_601,In_1078,In_901);
xnor U602 (N_602,In_1089,In_505);
nand U603 (N_603,In_1470,In_893);
or U604 (N_604,In_192,In_753);
xor U605 (N_605,In_1142,In_1157);
nand U606 (N_606,In_264,In_1153);
nand U607 (N_607,In_850,In_1185);
and U608 (N_608,In_243,In_1054);
nand U609 (N_609,In_1392,In_489);
and U610 (N_610,In_584,In_986);
xnor U611 (N_611,In_656,In_645);
or U612 (N_612,In_1261,In_47);
nor U613 (N_613,In_194,In_939);
and U614 (N_614,In_1234,In_977);
nand U615 (N_615,In_964,In_1069);
or U616 (N_616,In_1364,In_223);
xnor U617 (N_617,In_398,In_562);
nand U618 (N_618,In_482,In_769);
nor U619 (N_619,In_220,In_62);
nand U620 (N_620,In_683,In_409);
and U621 (N_621,In_430,In_1384);
xor U622 (N_622,In_166,In_807);
xor U623 (N_623,In_1301,In_446);
xor U624 (N_624,In_1091,In_1318);
and U625 (N_625,In_983,In_794);
or U626 (N_626,In_962,In_894);
and U627 (N_627,In_78,In_1249);
xnor U628 (N_628,In_111,In_1017);
or U629 (N_629,In_392,In_452);
xor U630 (N_630,In_805,In_1399);
and U631 (N_631,In_1426,In_1474);
nor U632 (N_632,In_655,In_703);
and U633 (N_633,In_1255,In_554);
and U634 (N_634,In_686,In_25);
nor U635 (N_635,In_15,In_912);
or U636 (N_636,In_9,In_28);
xor U637 (N_637,In_981,In_92);
nand U638 (N_638,In_182,In_928);
or U639 (N_639,In_1,In_1264);
or U640 (N_640,In_353,In_752);
xor U641 (N_641,In_347,In_316);
and U642 (N_642,In_1272,In_415);
and U643 (N_643,In_101,In_1449);
and U644 (N_644,In_1292,In_1453);
and U645 (N_645,In_1464,In_527);
or U646 (N_646,In_781,In_395);
and U647 (N_647,In_1000,In_609);
nand U648 (N_648,In_1051,In_640);
or U649 (N_649,In_1397,In_1497);
or U650 (N_650,In_1037,In_1087);
or U651 (N_651,In_1027,In_40);
and U652 (N_652,In_1342,In_1304);
xnor U653 (N_653,In_1324,In_1336);
nor U654 (N_654,In_799,In_19);
and U655 (N_655,In_709,In_1055);
nand U656 (N_656,In_650,In_988);
or U657 (N_657,In_842,In_1033);
and U658 (N_658,In_1178,In_969);
nor U659 (N_659,In_254,In_659);
xnor U660 (N_660,In_1273,In_1144);
xnor U661 (N_661,In_1285,In_448);
nor U662 (N_662,In_502,In_1433);
or U663 (N_663,In_1045,In_736);
and U664 (N_664,In_149,In_210);
nor U665 (N_665,In_1220,In_862);
nand U666 (N_666,In_368,In_651);
nand U667 (N_667,In_984,In_545);
and U668 (N_668,In_1013,In_1323);
or U669 (N_669,In_1322,In_882);
nor U670 (N_670,In_1461,In_530);
nor U671 (N_671,In_312,In_1072);
nor U672 (N_672,In_990,In_1427);
nand U673 (N_673,In_433,In_590);
or U674 (N_674,In_37,In_497);
or U675 (N_675,In_1303,In_233);
nand U676 (N_676,In_73,In_637);
or U677 (N_677,In_1191,In_6);
or U678 (N_678,In_309,In_636);
nand U679 (N_679,In_1431,In_1154);
nand U680 (N_680,In_916,In_1184);
and U681 (N_681,In_8,In_688);
and U682 (N_682,In_310,In_38);
xnor U683 (N_683,In_462,In_151);
or U684 (N_684,In_869,In_195);
nor U685 (N_685,In_795,In_917);
nand U686 (N_686,In_643,In_388);
and U687 (N_687,In_242,In_669);
nor U688 (N_688,In_240,In_334);
nor U689 (N_689,In_463,In_320);
nor U690 (N_690,In_1376,In_1213);
or U691 (N_691,In_3,In_275);
nand U692 (N_692,In_249,In_1171);
or U693 (N_693,In_1038,In_297);
and U694 (N_694,In_713,In_466);
and U695 (N_695,In_1029,In_293);
nand U696 (N_696,In_1267,In_387);
and U697 (N_697,In_1127,In_508);
nor U698 (N_698,In_14,In_619);
nand U699 (N_699,In_888,In_1424);
and U700 (N_700,In_997,In_978);
and U701 (N_701,In_1359,In_572);
nand U702 (N_702,In_373,In_1417);
or U703 (N_703,In_442,In_946);
and U704 (N_704,In_948,In_422);
nand U705 (N_705,In_1487,In_1238);
nor U706 (N_706,In_1183,In_259);
nor U707 (N_707,In_476,In_1477);
or U708 (N_708,In_598,In_1404);
nor U709 (N_709,In_239,In_1179);
nor U710 (N_710,In_529,In_742);
nor U711 (N_711,In_183,In_744);
or U712 (N_712,In_661,In_177);
nor U713 (N_713,In_55,In_644);
and U714 (N_714,In_1110,In_1351);
and U715 (N_715,In_99,In_627);
nand U716 (N_716,In_1099,In_364);
nand U717 (N_717,In_689,In_559);
and U718 (N_718,In_801,In_114);
and U719 (N_719,In_200,In_201);
nand U720 (N_720,In_391,In_72);
nor U721 (N_721,In_1362,In_1188);
and U722 (N_722,In_576,In_1208);
nand U723 (N_723,In_128,In_1475);
nand U724 (N_724,In_672,In_811);
xnor U725 (N_725,In_1451,In_868);
or U726 (N_726,In_1147,In_760);
xnor U727 (N_727,In_1167,In_399);
nor U728 (N_728,In_1490,In_314);
nand U729 (N_729,In_1278,In_158);
xor U730 (N_730,In_1221,In_139);
xor U731 (N_731,In_621,In_1085);
or U732 (N_732,In_1169,In_539);
and U733 (N_733,In_1439,In_1030);
nand U734 (N_734,In_1412,In_583);
xnor U735 (N_735,In_172,In_338);
nand U736 (N_736,In_926,In_188);
xnor U737 (N_737,In_1226,In_351);
or U738 (N_738,In_1481,In_1193);
xnor U739 (N_739,In_1165,In_500);
or U740 (N_740,In_973,In_620);
and U741 (N_741,In_1121,In_694);
and U742 (N_742,In_1047,In_302);
and U743 (N_743,In_180,In_122);
xnor U744 (N_744,In_682,In_1079);
nand U745 (N_745,In_227,In_70);
or U746 (N_746,In_350,In_337);
xor U747 (N_747,In_315,In_594);
nand U748 (N_748,In_748,In_396);
nor U749 (N_749,In_1057,In_140);
and U750 (N_750,N_30,N_552);
nand U751 (N_751,N_708,N_495);
nor U752 (N_752,N_301,N_542);
nand U753 (N_753,N_689,N_524);
and U754 (N_754,N_73,N_169);
xnor U755 (N_755,N_366,N_71);
and U756 (N_756,N_704,N_685);
nor U757 (N_757,N_715,N_386);
nor U758 (N_758,N_458,N_218);
nand U759 (N_759,N_637,N_151);
and U760 (N_760,N_467,N_729);
and U761 (N_761,N_713,N_201);
nor U762 (N_762,N_247,N_735);
or U763 (N_763,N_320,N_677);
xnor U764 (N_764,N_562,N_720);
or U765 (N_765,N_266,N_354);
nor U766 (N_766,N_272,N_402);
and U767 (N_767,N_457,N_550);
xor U768 (N_768,N_722,N_5);
nand U769 (N_769,N_268,N_614);
xor U770 (N_770,N_687,N_167);
nand U771 (N_771,N_84,N_516);
nor U772 (N_772,N_517,N_257);
nand U773 (N_773,N_630,N_97);
nor U774 (N_774,N_711,N_326);
nor U775 (N_775,N_592,N_2);
or U776 (N_776,N_621,N_283);
nor U777 (N_777,N_34,N_349);
nand U778 (N_778,N_565,N_277);
and U779 (N_779,N_246,N_703);
nor U780 (N_780,N_16,N_615);
or U781 (N_781,N_184,N_357);
nand U782 (N_782,N_649,N_398);
and U783 (N_783,N_665,N_700);
nor U784 (N_784,N_577,N_271);
or U785 (N_785,N_96,N_510);
or U786 (N_786,N_578,N_198);
nand U787 (N_787,N_11,N_165);
nor U788 (N_788,N_119,N_748);
nor U789 (N_789,N_551,N_26);
or U790 (N_790,N_709,N_323);
xor U791 (N_791,N_555,N_408);
and U792 (N_792,N_50,N_199);
and U793 (N_793,N_481,N_444);
and U794 (N_794,N_436,N_237);
and U795 (N_795,N_439,N_705);
nor U796 (N_796,N_308,N_233);
and U797 (N_797,N_528,N_75);
nor U798 (N_798,N_168,N_372);
nand U799 (N_799,N_632,N_92);
xnor U800 (N_800,N_429,N_23);
and U801 (N_801,N_314,N_527);
and U802 (N_802,N_497,N_362);
xor U803 (N_803,N_412,N_673);
nor U804 (N_804,N_728,N_482);
nand U805 (N_805,N_724,N_142);
or U806 (N_806,N_437,N_139);
xnor U807 (N_807,N_342,N_638);
nand U808 (N_808,N_440,N_202);
and U809 (N_809,N_148,N_253);
xnor U810 (N_810,N_57,N_19);
and U811 (N_811,N_701,N_537);
nand U812 (N_812,N_146,N_573);
nand U813 (N_813,N_593,N_411);
nand U814 (N_814,N_273,N_426);
or U815 (N_815,N_302,N_579);
or U816 (N_816,N_667,N_491);
or U817 (N_817,N_209,N_397);
nand U818 (N_818,N_441,N_417);
nand U819 (N_819,N_175,N_640);
xor U820 (N_820,N_616,N_446);
nand U821 (N_821,N_217,N_35);
nor U822 (N_822,N_191,N_331);
xnor U823 (N_823,N_594,N_694);
nand U824 (N_824,N_737,N_631);
and U825 (N_825,N_636,N_582);
nor U826 (N_826,N_298,N_24);
nor U827 (N_827,N_154,N_157);
xnor U828 (N_828,N_628,N_33);
xor U829 (N_829,N_43,N_313);
and U830 (N_830,N_507,N_619);
and U831 (N_831,N_477,N_341);
and U832 (N_832,N_605,N_546);
xnor U833 (N_833,N_414,N_221);
or U834 (N_834,N_89,N_442);
and U835 (N_835,N_663,N_473);
or U836 (N_836,N_378,N_275);
nor U837 (N_837,N_211,N_435);
and U838 (N_838,N_560,N_415);
nor U839 (N_839,N_425,N_145);
nand U840 (N_840,N_364,N_282);
or U841 (N_841,N_557,N_658);
and U842 (N_842,N_674,N_219);
nand U843 (N_843,N_493,N_574);
nand U844 (N_844,N_120,N_171);
or U845 (N_845,N_147,N_177);
nand U846 (N_846,N_186,N_393);
or U847 (N_847,N_624,N_395);
and U848 (N_848,N_488,N_185);
nor U849 (N_849,N_498,N_589);
nor U850 (N_850,N_133,N_305);
or U851 (N_851,N_403,N_152);
nand U852 (N_852,N_492,N_545);
or U853 (N_853,N_194,N_261);
nor U854 (N_854,N_170,N_262);
nand U855 (N_855,N_114,N_127);
nor U856 (N_856,N_315,N_113);
xnor U857 (N_857,N_483,N_93);
and U858 (N_858,N_377,N_264);
nand U859 (N_859,N_732,N_68);
xor U860 (N_860,N_633,N_613);
or U861 (N_861,N_438,N_249);
nor U862 (N_862,N_723,N_310);
nand U863 (N_863,N_197,N_454);
or U864 (N_864,N_486,N_714);
and U865 (N_865,N_459,N_462);
nand U866 (N_866,N_598,N_375);
xnor U867 (N_867,N_309,N_269);
nand U868 (N_868,N_245,N_99);
or U869 (N_869,N_427,N_83);
or U870 (N_870,N_501,N_285);
and U871 (N_871,N_278,N_222);
or U872 (N_872,N_718,N_404);
nand U873 (N_873,N_466,N_215);
xor U874 (N_874,N_596,N_340);
nor U875 (N_875,N_334,N_286);
nor U876 (N_876,N_746,N_153);
nor U877 (N_877,N_472,N_480);
or U878 (N_878,N_259,N_409);
or U879 (N_879,N_679,N_654);
nand U880 (N_880,N_164,N_39);
nor U881 (N_881,N_210,N_413);
xnor U882 (N_882,N_379,N_626);
nor U883 (N_883,N_248,N_112);
xor U884 (N_884,N_163,N_660);
nor U885 (N_885,N_287,N_59);
xnor U886 (N_886,N_242,N_150);
nor U887 (N_887,N_586,N_470);
nand U888 (N_888,N_355,N_489);
and U889 (N_889,N_647,N_428);
and U890 (N_890,N_474,N_290);
or U891 (N_891,N_680,N_612);
xor U892 (N_892,N_289,N_144);
nor U893 (N_893,N_235,N_200);
nor U894 (N_894,N_9,N_584);
and U895 (N_895,N_622,N_155);
or U896 (N_896,N_223,N_69);
nor U897 (N_897,N_333,N_338);
nor U898 (N_898,N_239,N_123);
and U899 (N_899,N_38,N_696);
nor U900 (N_900,N_125,N_182);
nor U901 (N_901,N_588,N_580);
nand U902 (N_902,N_388,N_747);
and U903 (N_903,N_618,N_452);
or U904 (N_904,N_360,N_190);
or U905 (N_905,N_321,N_585);
or U906 (N_906,N_361,N_387);
xnor U907 (N_907,N_293,N_743);
and U908 (N_908,N_686,N_672);
xor U909 (N_909,N_443,N_183);
xor U910 (N_910,N_553,N_207);
and U911 (N_911,N_424,N_79);
nand U912 (N_912,N_433,N_118);
nor U913 (N_913,N_47,N_692);
and U914 (N_914,N_234,N_396);
or U915 (N_915,N_319,N_14);
nor U916 (N_916,N_487,N_549);
or U917 (N_917,N_250,N_52);
or U918 (N_918,N_464,N_742);
nand U919 (N_919,N_284,N_351);
nor U920 (N_920,N_243,N_554);
or U921 (N_921,N_116,N_325);
and U922 (N_922,N_85,N_206);
xnor U923 (N_923,N_611,N_121);
nand U924 (N_924,N_258,N_350);
or U925 (N_925,N_451,N_385);
and U926 (N_926,N_140,N_571);
xnor U927 (N_927,N_311,N_670);
or U928 (N_928,N_664,N_279);
xnor U929 (N_929,N_421,N_359);
xnor U930 (N_930,N_179,N_77);
nand U931 (N_931,N_371,N_126);
nand U932 (N_932,N_41,N_352);
or U933 (N_933,N_365,N_539);
nand U934 (N_934,N_336,N_490);
nor U935 (N_935,N_6,N_270);
nor U936 (N_936,N_343,N_27);
nand U937 (N_937,N_12,N_499);
nand U938 (N_938,N_511,N_540);
nand U939 (N_939,N_115,N_382);
and U940 (N_940,N_274,N_690);
or U941 (N_941,N_641,N_203);
xor U942 (N_942,N_373,N_42);
and U943 (N_943,N_263,N_204);
nor U944 (N_944,N_58,N_716);
and U945 (N_945,N_731,N_111);
nor U946 (N_946,N_399,N_383);
and U947 (N_947,N_668,N_188);
nand U948 (N_948,N_90,N_122);
nor U949 (N_949,N_66,N_564);
or U950 (N_950,N_644,N_535);
nor U951 (N_951,N_538,N_740);
and U952 (N_952,N_353,N_478);
xor U953 (N_953,N_244,N_513);
xor U954 (N_954,N_617,N_518);
xnor U955 (N_955,N_189,N_337);
nand U956 (N_956,N_318,N_512);
nor U957 (N_957,N_707,N_335);
nor U958 (N_958,N_31,N_590);
nor U959 (N_959,N_381,N_607);
xor U960 (N_960,N_659,N_25);
and U961 (N_961,N_160,N_698);
nor U962 (N_962,N_136,N_392);
nor U963 (N_963,N_423,N_608);
or U964 (N_964,N_176,N_260);
nand U965 (N_965,N_505,N_520);
or U966 (N_966,N_655,N_306);
nor U967 (N_967,N_141,N_471);
xor U968 (N_968,N_529,N_62);
nand U969 (N_969,N_651,N_149);
nor U970 (N_970,N_48,N_702);
nand U971 (N_971,N_627,N_297);
or U972 (N_972,N_220,N_479);
or U973 (N_973,N_61,N_254);
nor U974 (N_974,N_216,N_156);
nor U975 (N_975,N_128,N_556);
nand U976 (N_976,N_132,N_347);
nand U977 (N_977,N_602,N_54);
or U978 (N_978,N_135,N_653);
or U979 (N_979,N_80,N_389);
nand U980 (N_980,N_238,N_374);
xor U981 (N_981,N_32,N_496);
nand U982 (N_982,N_662,N_706);
and U983 (N_983,N_671,N_604);
nor U984 (N_984,N_205,N_712);
and U985 (N_985,N_502,N_240);
or U986 (N_986,N_51,N_161);
and U987 (N_987,N_67,N_460);
nor U988 (N_988,N_46,N_195);
and U989 (N_989,N_583,N_212);
xor U990 (N_990,N_504,N_695);
nor U991 (N_991,N_70,N_358);
xor U992 (N_992,N_87,N_610);
and U993 (N_993,N_453,N_676);
nor U994 (N_994,N_106,N_107);
or U995 (N_995,N_400,N_60);
and U996 (N_996,N_569,N_316);
and U997 (N_997,N_434,N_265);
xor U998 (N_998,N_44,N_251);
nand U999 (N_999,N_575,N_213);
or U1000 (N_1000,N_652,N_566);
and U1001 (N_1001,N_241,N_523);
or U1002 (N_1002,N_697,N_558);
and U1003 (N_1003,N_563,N_448);
nor U1004 (N_1004,N_101,N_669);
xor U1005 (N_1005,N_288,N_304);
nor U1006 (N_1006,N_29,N_603);
or U1007 (N_1007,N_280,N_410);
and U1008 (N_1008,N_744,N_208);
xor U1009 (N_1009,N_406,N_226);
nor U1010 (N_1010,N_0,N_678);
nor U1011 (N_1011,N_532,N_100);
nand U1012 (N_1012,N_431,N_508);
xnor U1013 (N_1013,N_368,N_521);
nand U1014 (N_1014,N_228,N_173);
or U1015 (N_1015,N_291,N_739);
nand U1016 (N_1016,N_4,N_339);
nor U1017 (N_1017,N_683,N_587);
or U1018 (N_1018,N_475,N_256);
and U1019 (N_1019,N_432,N_420);
or U1020 (N_1020,N_623,N_648);
xor U1021 (N_1021,N_231,N_348);
xor U1022 (N_1022,N_595,N_634);
nand U1023 (N_1023,N_419,N_95);
or U1024 (N_1024,N_500,N_28);
xnor U1025 (N_1025,N_620,N_193);
xnor U1026 (N_1026,N_78,N_710);
xnor U1027 (N_1027,N_18,N_643);
and U1028 (N_1028,N_717,N_736);
nand U1029 (N_1029,N_65,N_172);
xnor U1030 (N_1030,N_738,N_721);
xor U1031 (N_1031,N_559,N_682);
nor U1032 (N_1032,N_447,N_324);
nor U1033 (N_1033,N_416,N_450);
xor U1034 (N_1034,N_503,N_22);
xnor U1035 (N_1035,N_646,N_327);
xnor U1036 (N_1036,N_294,N_267);
nand U1037 (N_1037,N_40,N_749);
nand U1038 (N_1038,N_21,N_53);
xnor U1039 (N_1039,N_681,N_576);
nand U1040 (N_1040,N_192,N_380);
and U1041 (N_1041,N_162,N_449);
nor U1042 (N_1042,N_86,N_329);
xnor U1043 (N_1043,N_129,N_376);
or U1044 (N_1044,N_137,N_300);
and U1045 (N_1045,N_105,N_699);
nor U1046 (N_1046,N_158,N_691);
and U1047 (N_1047,N_312,N_405);
xnor U1048 (N_1048,N_461,N_15);
nor U1049 (N_1049,N_606,N_572);
or U1050 (N_1050,N_130,N_322);
xor U1051 (N_1051,N_224,N_591);
xor U1052 (N_1052,N_629,N_548);
or U1053 (N_1053,N_561,N_346);
nor U1054 (N_1054,N_401,N_196);
or U1055 (N_1055,N_635,N_544);
and U1056 (N_1056,N_255,N_124);
xor U1057 (N_1057,N_7,N_64);
and U1058 (N_1058,N_91,N_36);
and U1059 (N_1059,N_656,N_317);
and U1060 (N_1060,N_407,N_102);
xor U1061 (N_1061,N_642,N_296);
nor U1062 (N_1062,N_650,N_688);
nor U1063 (N_1063,N_369,N_609);
nand U1064 (N_1064,N_63,N_236);
or U1065 (N_1065,N_675,N_476);
nor U1066 (N_1066,N_295,N_20);
and U1067 (N_1067,N_485,N_465);
or U1068 (N_1068,N_657,N_117);
nand U1069 (N_1069,N_494,N_456);
xnor U1070 (N_1070,N_567,N_82);
or U1071 (N_1071,N_8,N_187);
xor U1072 (N_1072,N_547,N_328);
or U1073 (N_1073,N_230,N_98);
xor U1074 (N_1074,N_639,N_109);
nor U1075 (N_1075,N_108,N_509);
or U1076 (N_1076,N_276,N_536);
and U1077 (N_1077,N_370,N_74);
or U1078 (N_1078,N_1,N_143);
and U1079 (N_1079,N_134,N_726);
nor U1080 (N_1080,N_344,N_225);
nand U1081 (N_1081,N_94,N_110);
or U1082 (N_1082,N_367,N_81);
nor U1083 (N_1083,N_430,N_445);
nand U1084 (N_1084,N_390,N_391);
and U1085 (N_1085,N_345,N_541);
or U1086 (N_1086,N_741,N_166);
nor U1087 (N_1087,N_684,N_17);
and U1088 (N_1088,N_468,N_356);
xnor U1089 (N_1089,N_104,N_76);
xor U1090 (N_1090,N_159,N_394);
xnor U1091 (N_1091,N_418,N_181);
xnor U1092 (N_1092,N_292,N_463);
and U1093 (N_1093,N_88,N_384);
nor U1094 (N_1094,N_227,N_745);
and U1095 (N_1095,N_37,N_3);
or U1096 (N_1096,N_730,N_229);
nor U1097 (N_1097,N_484,N_180);
or U1098 (N_1098,N_599,N_533);
xor U1099 (N_1099,N_56,N_55);
nor U1100 (N_1100,N_330,N_45);
or U1101 (N_1101,N_601,N_303);
or U1102 (N_1102,N_725,N_49);
nor U1103 (N_1103,N_666,N_597);
and U1104 (N_1104,N_469,N_525);
nor U1105 (N_1105,N_530,N_299);
xor U1106 (N_1106,N_568,N_733);
nor U1107 (N_1107,N_693,N_232);
or U1108 (N_1108,N_534,N_131);
nor U1109 (N_1109,N_514,N_734);
nor U1110 (N_1110,N_543,N_522);
and U1111 (N_1111,N_252,N_10);
nor U1112 (N_1112,N_214,N_727);
nor U1113 (N_1113,N_645,N_570);
xnor U1114 (N_1114,N_531,N_455);
or U1115 (N_1115,N_515,N_600);
xnor U1116 (N_1116,N_178,N_506);
nand U1117 (N_1117,N_519,N_174);
and U1118 (N_1118,N_13,N_581);
nand U1119 (N_1119,N_363,N_719);
and U1120 (N_1120,N_307,N_72);
nand U1121 (N_1121,N_526,N_661);
nor U1122 (N_1122,N_625,N_281);
nand U1123 (N_1123,N_138,N_103);
nand U1124 (N_1124,N_422,N_332);
or U1125 (N_1125,N_196,N_534);
xor U1126 (N_1126,N_227,N_660);
nor U1127 (N_1127,N_249,N_604);
nor U1128 (N_1128,N_557,N_429);
xnor U1129 (N_1129,N_550,N_559);
or U1130 (N_1130,N_408,N_115);
xnor U1131 (N_1131,N_48,N_197);
nor U1132 (N_1132,N_32,N_151);
or U1133 (N_1133,N_231,N_91);
and U1134 (N_1134,N_461,N_59);
and U1135 (N_1135,N_616,N_339);
nand U1136 (N_1136,N_156,N_83);
or U1137 (N_1137,N_535,N_263);
nand U1138 (N_1138,N_538,N_54);
xor U1139 (N_1139,N_699,N_612);
nor U1140 (N_1140,N_522,N_235);
nand U1141 (N_1141,N_623,N_184);
nand U1142 (N_1142,N_193,N_275);
xnor U1143 (N_1143,N_519,N_623);
nor U1144 (N_1144,N_223,N_594);
or U1145 (N_1145,N_513,N_78);
nand U1146 (N_1146,N_459,N_246);
nor U1147 (N_1147,N_218,N_148);
xor U1148 (N_1148,N_369,N_749);
nor U1149 (N_1149,N_383,N_262);
or U1150 (N_1150,N_427,N_512);
xor U1151 (N_1151,N_109,N_631);
or U1152 (N_1152,N_3,N_689);
xnor U1153 (N_1153,N_136,N_127);
or U1154 (N_1154,N_694,N_550);
nor U1155 (N_1155,N_145,N_103);
and U1156 (N_1156,N_692,N_700);
nor U1157 (N_1157,N_402,N_201);
nor U1158 (N_1158,N_73,N_447);
nor U1159 (N_1159,N_145,N_35);
xor U1160 (N_1160,N_63,N_411);
and U1161 (N_1161,N_120,N_584);
nand U1162 (N_1162,N_463,N_624);
or U1163 (N_1163,N_350,N_320);
nor U1164 (N_1164,N_72,N_57);
and U1165 (N_1165,N_65,N_595);
or U1166 (N_1166,N_258,N_364);
nor U1167 (N_1167,N_428,N_381);
nand U1168 (N_1168,N_468,N_324);
nor U1169 (N_1169,N_321,N_196);
nand U1170 (N_1170,N_162,N_199);
nand U1171 (N_1171,N_711,N_14);
and U1172 (N_1172,N_32,N_16);
and U1173 (N_1173,N_549,N_396);
nor U1174 (N_1174,N_194,N_419);
nand U1175 (N_1175,N_223,N_304);
nand U1176 (N_1176,N_152,N_609);
xor U1177 (N_1177,N_369,N_516);
nor U1178 (N_1178,N_654,N_668);
nor U1179 (N_1179,N_674,N_401);
nor U1180 (N_1180,N_73,N_511);
and U1181 (N_1181,N_500,N_603);
or U1182 (N_1182,N_278,N_101);
xnor U1183 (N_1183,N_284,N_559);
nor U1184 (N_1184,N_402,N_135);
xor U1185 (N_1185,N_340,N_47);
nand U1186 (N_1186,N_565,N_223);
and U1187 (N_1187,N_655,N_690);
nand U1188 (N_1188,N_208,N_502);
nand U1189 (N_1189,N_517,N_471);
nor U1190 (N_1190,N_605,N_450);
or U1191 (N_1191,N_37,N_29);
nor U1192 (N_1192,N_384,N_625);
nand U1193 (N_1193,N_236,N_160);
nor U1194 (N_1194,N_435,N_414);
xor U1195 (N_1195,N_496,N_104);
nand U1196 (N_1196,N_383,N_30);
and U1197 (N_1197,N_260,N_285);
or U1198 (N_1198,N_469,N_493);
nand U1199 (N_1199,N_573,N_36);
or U1200 (N_1200,N_584,N_215);
and U1201 (N_1201,N_610,N_51);
xor U1202 (N_1202,N_668,N_115);
xnor U1203 (N_1203,N_302,N_50);
nor U1204 (N_1204,N_192,N_220);
nor U1205 (N_1205,N_405,N_680);
nor U1206 (N_1206,N_83,N_380);
nor U1207 (N_1207,N_130,N_635);
nand U1208 (N_1208,N_423,N_506);
nor U1209 (N_1209,N_434,N_701);
nor U1210 (N_1210,N_695,N_485);
xnor U1211 (N_1211,N_553,N_562);
xnor U1212 (N_1212,N_607,N_302);
or U1213 (N_1213,N_625,N_284);
xnor U1214 (N_1214,N_746,N_516);
xnor U1215 (N_1215,N_293,N_127);
or U1216 (N_1216,N_379,N_466);
or U1217 (N_1217,N_95,N_512);
nand U1218 (N_1218,N_378,N_211);
nor U1219 (N_1219,N_407,N_489);
xor U1220 (N_1220,N_490,N_529);
or U1221 (N_1221,N_231,N_673);
nor U1222 (N_1222,N_168,N_353);
and U1223 (N_1223,N_448,N_514);
nor U1224 (N_1224,N_662,N_293);
or U1225 (N_1225,N_223,N_66);
xor U1226 (N_1226,N_487,N_520);
xnor U1227 (N_1227,N_724,N_737);
or U1228 (N_1228,N_355,N_213);
nor U1229 (N_1229,N_584,N_479);
xor U1230 (N_1230,N_537,N_164);
nand U1231 (N_1231,N_16,N_151);
and U1232 (N_1232,N_292,N_220);
nor U1233 (N_1233,N_194,N_491);
nand U1234 (N_1234,N_341,N_177);
or U1235 (N_1235,N_377,N_334);
or U1236 (N_1236,N_33,N_146);
nand U1237 (N_1237,N_184,N_353);
nand U1238 (N_1238,N_370,N_569);
nor U1239 (N_1239,N_223,N_588);
or U1240 (N_1240,N_201,N_327);
or U1241 (N_1241,N_683,N_136);
nand U1242 (N_1242,N_617,N_570);
nand U1243 (N_1243,N_408,N_92);
or U1244 (N_1244,N_645,N_670);
or U1245 (N_1245,N_435,N_550);
xnor U1246 (N_1246,N_638,N_201);
nor U1247 (N_1247,N_619,N_380);
nor U1248 (N_1248,N_269,N_276);
nor U1249 (N_1249,N_699,N_220);
and U1250 (N_1250,N_744,N_291);
nand U1251 (N_1251,N_325,N_310);
nor U1252 (N_1252,N_167,N_4);
nand U1253 (N_1253,N_456,N_695);
xnor U1254 (N_1254,N_204,N_305);
xor U1255 (N_1255,N_214,N_373);
or U1256 (N_1256,N_147,N_589);
nand U1257 (N_1257,N_328,N_530);
xnor U1258 (N_1258,N_33,N_89);
xnor U1259 (N_1259,N_34,N_355);
and U1260 (N_1260,N_744,N_564);
nand U1261 (N_1261,N_561,N_78);
or U1262 (N_1262,N_243,N_699);
or U1263 (N_1263,N_704,N_180);
nor U1264 (N_1264,N_542,N_167);
nor U1265 (N_1265,N_416,N_94);
and U1266 (N_1266,N_711,N_721);
or U1267 (N_1267,N_395,N_182);
xnor U1268 (N_1268,N_234,N_700);
nor U1269 (N_1269,N_551,N_94);
nand U1270 (N_1270,N_492,N_445);
nand U1271 (N_1271,N_279,N_620);
nor U1272 (N_1272,N_176,N_544);
nor U1273 (N_1273,N_554,N_735);
or U1274 (N_1274,N_129,N_563);
and U1275 (N_1275,N_58,N_457);
and U1276 (N_1276,N_672,N_725);
xnor U1277 (N_1277,N_191,N_501);
nor U1278 (N_1278,N_744,N_599);
nor U1279 (N_1279,N_719,N_340);
xor U1280 (N_1280,N_97,N_677);
or U1281 (N_1281,N_434,N_505);
and U1282 (N_1282,N_29,N_126);
and U1283 (N_1283,N_85,N_680);
and U1284 (N_1284,N_296,N_25);
nand U1285 (N_1285,N_352,N_287);
nand U1286 (N_1286,N_269,N_577);
nor U1287 (N_1287,N_102,N_716);
xor U1288 (N_1288,N_637,N_611);
xor U1289 (N_1289,N_690,N_106);
nor U1290 (N_1290,N_264,N_54);
nand U1291 (N_1291,N_131,N_454);
or U1292 (N_1292,N_62,N_579);
nor U1293 (N_1293,N_116,N_648);
xor U1294 (N_1294,N_45,N_568);
nor U1295 (N_1295,N_485,N_164);
and U1296 (N_1296,N_349,N_653);
nor U1297 (N_1297,N_659,N_353);
or U1298 (N_1298,N_97,N_590);
and U1299 (N_1299,N_221,N_539);
or U1300 (N_1300,N_11,N_99);
xor U1301 (N_1301,N_13,N_571);
and U1302 (N_1302,N_324,N_405);
xor U1303 (N_1303,N_143,N_275);
nor U1304 (N_1304,N_259,N_731);
nand U1305 (N_1305,N_642,N_186);
or U1306 (N_1306,N_213,N_318);
or U1307 (N_1307,N_468,N_722);
nand U1308 (N_1308,N_196,N_471);
or U1309 (N_1309,N_607,N_606);
nor U1310 (N_1310,N_56,N_583);
nand U1311 (N_1311,N_400,N_740);
nor U1312 (N_1312,N_412,N_450);
or U1313 (N_1313,N_241,N_151);
and U1314 (N_1314,N_143,N_548);
nand U1315 (N_1315,N_210,N_212);
nand U1316 (N_1316,N_679,N_211);
xor U1317 (N_1317,N_723,N_652);
or U1318 (N_1318,N_61,N_99);
or U1319 (N_1319,N_114,N_575);
and U1320 (N_1320,N_271,N_92);
and U1321 (N_1321,N_126,N_96);
nand U1322 (N_1322,N_501,N_207);
and U1323 (N_1323,N_103,N_379);
and U1324 (N_1324,N_688,N_385);
nand U1325 (N_1325,N_635,N_501);
nand U1326 (N_1326,N_413,N_236);
xnor U1327 (N_1327,N_422,N_198);
and U1328 (N_1328,N_214,N_131);
nor U1329 (N_1329,N_615,N_158);
or U1330 (N_1330,N_408,N_398);
xor U1331 (N_1331,N_703,N_411);
and U1332 (N_1332,N_663,N_591);
xor U1333 (N_1333,N_165,N_93);
xor U1334 (N_1334,N_53,N_594);
xnor U1335 (N_1335,N_600,N_384);
nor U1336 (N_1336,N_270,N_635);
nand U1337 (N_1337,N_545,N_377);
nor U1338 (N_1338,N_331,N_332);
or U1339 (N_1339,N_392,N_249);
or U1340 (N_1340,N_400,N_331);
and U1341 (N_1341,N_661,N_457);
xor U1342 (N_1342,N_57,N_15);
and U1343 (N_1343,N_452,N_578);
nor U1344 (N_1344,N_593,N_475);
nand U1345 (N_1345,N_320,N_249);
and U1346 (N_1346,N_134,N_343);
and U1347 (N_1347,N_394,N_438);
and U1348 (N_1348,N_247,N_293);
and U1349 (N_1349,N_621,N_402);
or U1350 (N_1350,N_393,N_471);
nand U1351 (N_1351,N_194,N_54);
or U1352 (N_1352,N_210,N_489);
and U1353 (N_1353,N_71,N_337);
xnor U1354 (N_1354,N_439,N_430);
nor U1355 (N_1355,N_46,N_643);
nand U1356 (N_1356,N_250,N_262);
xnor U1357 (N_1357,N_39,N_575);
or U1358 (N_1358,N_233,N_711);
and U1359 (N_1359,N_668,N_232);
nor U1360 (N_1360,N_253,N_574);
and U1361 (N_1361,N_142,N_6);
nor U1362 (N_1362,N_65,N_28);
nand U1363 (N_1363,N_558,N_265);
and U1364 (N_1364,N_587,N_518);
nand U1365 (N_1365,N_382,N_40);
nor U1366 (N_1366,N_65,N_563);
and U1367 (N_1367,N_630,N_483);
nand U1368 (N_1368,N_268,N_379);
or U1369 (N_1369,N_461,N_347);
or U1370 (N_1370,N_271,N_500);
nor U1371 (N_1371,N_599,N_315);
or U1372 (N_1372,N_245,N_451);
nor U1373 (N_1373,N_131,N_373);
and U1374 (N_1374,N_699,N_326);
xor U1375 (N_1375,N_360,N_662);
and U1376 (N_1376,N_223,N_158);
xor U1377 (N_1377,N_407,N_471);
nor U1378 (N_1378,N_530,N_457);
nor U1379 (N_1379,N_411,N_662);
and U1380 (N_1380,N_109,N_698);
and U1381 (N_1381,N_358,N_442);
nor U1382 (N_1382,N_592,N_702);
nand U1383 (N_1383,N_220,N_435);
nand U1384 (N_1384,N_537,N_670);
nand U1385 (N_1385,N_733,N_216);
nand U1386 (N_1386,N_604,N_740);
xor U1387 (N_1387,N_538,N_405);
xnor U1388 (N_1388,N_132,N_582);
nand U1389 (N_1389,N_743,N_676);
and U1390 (N_1390,N_557,N_128);
or U1391 (N_1391,N_176,N_500);
or U1392 (N_1392,N_56,N_64);
nor U1393 (N_1393,N_655,N_679);
xnor U1394 (N_1394,N_590,N_197);
nand U1395 (N_1395,N_635,N_489);
nor U1396 (N_1396,N_318,N_614);
nor U1397 (N_1397,N_21,N_257);
xor U1398 (N_1398,N_723,N_298);
nand U1399 (N_1399,N_517,N_488);
or U1400 (N_1400,N_261,N_431);
and U1401 (N_1401,N_312,N_161);
nand U1402 (N_1402,N_83,N_239);
nand U1403 (N_1403,N_475,N_356);
nor U1404 (N_1404,N_411,N_480);
and U1405 (N_1405,N_35,N_334);
and U1406 (N_1406,N_156,N_351);
xor U1407 (N_1407,N_446,N_141);
nand U1408 (N_1408,N_540,N_493);
nand U1409 (N_1409,N_250,N_240);
nand U1410 (N_1410,N_502,N_593);
xnor U1411 (N_1411,N_143,N_680);
xor U1412 (N_1412,N_655,N_383);
xnor U1413 (N_1413,N_222,N_81);
or U1414 (N_1414,N_670,N_388);
or U1415 (N_1415,N_557,N_347);
or U1416 (N_1416,N_175,N_676);
nor U1417 (N_1417,N_632,N_723);
and U1418 (N_1418,N_681,N_472);
nand U1419 (N_1419,N_428,N_203);
xor U1420 (N_1420,N_343,N_141);
and U1421 (N_1421,N_474,N_312);
nand U1422 (N_1422,N_425,N_691);
nor U1423 (N_1423,N_536,N_481);
or U1424 (N_1424,N_593,N_435);
nor U1425 (N_1425,N_428,N_220);
xnor U1426 (N_1426,N_446,N_554);
nand U1427 (N_1427,N_694,N_281);
and U1428 (N_1428,N_729,N_87);
nor U1429 (N_1429,N_653,N_332);
or U1430 (N_1430,N_562,N_431);
nand U1431 (N_1431,N_109,N_95);
or U1432 (N_1432,N_431,N_654);
and U1433 (N_1433,N_293,N_426);
and U1434 (N_1434,N_160,N_490);
or U1435 (N_1435,N_119,N_388);
nand U1436 (N_1436,N_407,N_173);
or U1437 (N_1437,N_38,N_608);
nand U1438 (N_1438,N_63,N_611);
or U1439 (N_1439,N_536,N_615);
and U1440 (N_1440,N_674,N_3);
and U1441 (N_1441,N_119,N_323);
xnor U1442 (N_1442,N_392,N_174);
xnor U1443 (N_1443,N_522,N_192);
xnor U1444 (N_1444,N_109,N_64);
or U1445 (N_1445,N_650,N_181);
xor U1446 (N_1446,N_261,N_94);
xnor U1447 (N_1447,N_34,N_559);
nand U1448 (N_1448,N_436,N_292);
nand U1449 (N_1449,N_685,N_473);
nand U1450 (N_1450,N_730,N_101);
nand U1451 (N_1451,N_201,N_527);
nor U1452 (N_1452,N_211,N_474);
nor U1453 (N_1453,N_542,N_29);
nand U1454 (N_1454,N_422,N_619);
nand U1455 (N_1455,N_114,N_124);
or U1456 (N_1456,N_591,N_329);
nor U1457 (N_1457,N_564,N_51);
nor U1458 (N_1458,N_199,N_264);
nor U1459 (N_1459,N_93,N_67);
nand U1460 (N_1460,N_206,N_264);
nand U1461 (N_1461,N_575,N_565);
nand U1462 (N_1462,N_629,N_500);
nor U1463 (N_1463,N_222,N_31);
or U1464 (N_1464,N_196,N_332);
xnor U1465 (N_1465,N_107,N_187);
nand U1466 (N_1466,N_287,N_516);
and U1467 (N_1467,N_482,N_207);
or U1468 (N_1468,N_652,N_473);
nand U1469 (N_1469,N_437,N_568);
and U1470 (N_1470,N_383,N_307);
or U1471 (N_1471,N_88,N_3);
nand U1472 (N_1472,N_320,N_393);
or U1473 (N_1473,N_197,N_433);
and U1474 (N_1474,N_647,N_181);
or U1475 (N_1475,N_204,N_659);
nand U1476 (N_1476,N_236,N_524);
xor U1477 (N_1477,N_462,N_348);
or U1478 (N_1478,N_64,N_276);
nor U1479 (N_1479,N_11,N_155);
and U1480 (N_1480,N_404,N_432);
and U1481 (N_1481,N_652,N_35);
nand U1482 (N_1482,N_133,N_411);
or U1483 (N_1483,N_189,N_27);
nor U1484 (N_1484,N_414,N_683);
xnor U1485 (N_1485,N_448,N_387);
and U1486 (N_1486,N_583,N_199);
or U1487 (N_1487,N_397,N_624);
nor U1488 (N_1488,N_112,N_414);
or U1489 (N_1489,N_495,N_605);
xor U1490 (N_1490,N_481,N_494);
and U1491 (N_1491,N_204,N_81);
xnor U1492 (N_1492,N_413,N_174);
nor U1493 (N_1493,N_130,N_640);
and U1494 (N_1494,N_530,N_20);
xor U1495 (N_1495,N_421,N_707);
and U1496 (N_1496,N_726,N_581);
xor U1497 (N_1497,N_451,N_570);
nor U1498 (N_1498,N_269,N_294);
nand U1499 (N_1499,N_327,N_662);
and U1500 (N_1500,N_958,N_845);
and U1501 (N_1501,N_984,N_1344);
nor U1502 (N_1502,N_1119,N_1436);
and U1503 (N_1503,N_1117,N_1282);
xor U1504 (N_1504,N_856,N_1074);
nand U1505 (N_1505,N_1192,N_1419);
or U1506 (N_1506,N_1176,N_753);
and U1507 (N_1507,N_1464,N_1247);
and U1508 (N_1508,N_1058,N_1337);
or U1509 (N_1509,N_794,N_898);
xnor U1510 (N_1510,N_760,N_1342);
or U1511 (N_1511,N_1311,N_1267);
and U1512 (N_1512,N_1110,N_1275);
xnor U1513 (N_1513,N_790,N_989);
xor U1514 (N_1514,N_1321,N_1017);
nor U1515 (N_1515,N_955,N_943);
nand U1516 (N_1516,N_1162,N_979);
xor U1517 (N_1517,N_1450,N_1491);
nand U1518 (N_1518,N_833,N_1047);
and U1519 (N_1519,N_1483,N_1052);
and U1520 (N_1520,N_1233,N_1087);
nand U1521 (N_1521,N_1187,N_776);
nand U1522 (N_1522,N_1349,N_942);
xnor U1523 (N_1523,N_859,N_1240);
nor U1524 (N_1524,N_1227,N_815);
nor U1525 (N_1525,N_1433,N_1265);
or U1526 (N_1526,N_1134,N_1099);
xnor U1527 (N_1527,N_1094,N_1408);
nand U1528 (N_1528,N_1010,N_1116);
or U1529 (N_1529,N_1118,N_1249);
nand U1530 (N_1530,N_1331,N_822);
xnor U1531 (N_1531,N_1487,N_824);
xor U1532 (N_1532,N_1077,N_851);
nor U1533 (N_1533,N_1068,N_812);
nor U1534 (N_1534,N_1031,N_1092);
or U1535 (N_1535,N_1071,N_892);
and U1536 (N_1536,N_1237,N_1406);
or U1537 (N_1537,N_1132,N_860);
nor U1538 (N_1538,N_768,N_1015);
and U1539 (N_1539,N_894,N_983);
and U1540 (N_1540,N_1289,N_1486);
nor U1541 (N_1541,N_1199,N_802);
nand U1542 (N_1542,N_820,N_1318);
nor U1543 (N_1543,N_974,N_1159);
and U1544 (N_1544,N_949,N_1059);
nand U1545 (N_1545,N_1498,N_1194);
nand U1546 (N_1546,N_1044,N_1332);
nand U1547 (N_1547,N_863,N_901);
or U1548 (N_1548,N_1231,N_987);
nand U1549 (N_1549,N_995,N_1365);
nor U1550 (N_1550,N_993,N_1163);
nand U1551 (N_1551,N_1209,N_1285);
nor U1552 (N_1552,N_1447,N_915);
nand U1553 (N_1553,N_778,N_1413);
nor U1554 (N_1554,N_1293,N_1355);
nand U1555 (N_1555,N_767,N_811);
nand U1556 (N_1556,N_880,N_1135);
xnor U1557 (N_1557,N_1012,N_950);
and U1558 (N_1558,N_1338,N_785);
xnor U1559 (N_1559,N_954,N_1198);
xor U1560 (N_1560,N_1426,N_1496);
and U1561 (N_1561,N_862,N_1095);
nor U1562 (N_1562,N_902,N_1383);
nand U1563 (N_1563,N_766,N_1394);
or U1564 (N_1564,N_826,N_1213);
or U1565 (N_1565,N_927,N_1003);
or U1566 (N_1566,N_816,N_1211);
or U1567 (N_1567,N_809,N_1361);
xor U1568 (N_1568,N_1229,N_928);
nor U1569 (N_1569,N_1066,N_1232);
and U1570 (N_1570,N_1272,N_1024);
xor U1571 (N_1571,N_962,N_827);
xor U1572 (N_1572,N_1401,N_1477);
xnor U1573 (N_1573,N_1151,N_1054);
nor U1574 (N_1574,N_946,N_1287);
and U1575 (N_1575,N_1370,N_1205);
and U1576 (N_1576,N_837,N_1298);
or U1577 (N_1577,N_1183,N_1167);
or U1578 (N_1578,N_1429,N_1043);
or U1579 (N_1579,N_934,N_960);
nor U1580 (N_1580,N_1421,N_1326);
xor U1581 (N_1581,N_900,N_913);
xnor U1582 (N_1582,N_1157,N_893);
nor U1583 (N_1583,N_1112,N_975);
xor U1584 (N_1584,N_821,N_825);
or U1585 (N_1585,N_1234,N_990);
nand U1586 (N_1586,N_770,N_1493);
nor U1587 (N_1587,N_1360,N_980);
xnor U1588 (N_1588,N_1263,N_930);
nand U1589 (N_1589,N_940,N_931);
or U1590 (N_1590,N_1432,N_945);
or U1591 (N_1591,N_1372,N_959);
nand U1592 (N_1592,N_1007,N_1105);
and U1593 (N_1593,N_1420,N_1171);
nor U1594 (N_1594,N_1316,N_764);
and U1595 (N_1595,N_921,N_999);
nor U1596 (N_1596,N_1352,N_1062);
and U1597 (N_1597,N_896,N_883);
and U1598 (N_1598,N_1441,N_1463);
xnor U1599 (N_1599,N_965,N_1301);
nor U1600 (N_1600,N_1107,N_1019);
and U1601 (N_1601,N_1423,N_976);
or U1602 (N_1602,N_1081,N_1091);
and U1603 (N_1603,N_1050,N_972);
nor U1604 (N_1604,N_904,N_1461);
nand U1605 (N_1605,N_879,N_850);
xnor U1606 (N_1606,N_1489,N_1359);
nor U1607 (N_1607,N_1482,N_1324);
nand U1608 (N_1608,N_1008,N_772);
or U1609 (N_1609,N_1350,N_1467);
or U1610 (N_1610,N_805,N_1197);
or U1611 (N_1611,N_1149,N_857);
nand U1612 (N_1612,N_933,N_1250);
xnor U1613 (N_1613,N_1085,N_813);
nor U1614 (N_1614,N_1177,N_1079);
and U1615 (N_1615,N_1204,N_874);
nor U1616 (N_1616,N_1458,N_819);
or U1617 (N_1617,N_1224,N_763);
nand U1618 (N_1618,N_1238,N_1174);
or U1619 (N_1619,N_951,N_1106);
nor U1620 (N_1620,N_1103,N_1312);
nand U1621 (N_1621,N_886,N_868);
nor U1622 (N_1622,N_761,N_1225);
or U1623 (N_1623,N_865,N_1184);
or U1624 (N_1624,N_1390,N_969);
xor U1625 (N_1625,N_1492,N_1290);
or U1626 (N_1626,N_1279,N_1442);
and U1627 (N_1627,N_973,N_1367);
nor U1628 (N_1628,N_1256,N_1283);
nor U1629 (N_1629,N_1303,N_905);
or U1630 (N_1630,N_1195,N_1378);
or U1631 (N_1631,N_1023,N_1366);
or U1632 (N_1632,N_1428,N_1154);
and U1633 (N_1633,N_1065,N_953);
or U1634 (N_1634,N_1111,N_1364);
xnor U1635 (N_1635,N_1398,N_1488);
and U1636 (N_1636,N_1029,N_1064);
nand U1637 (N_1637,N_1353,N_992);
and U1638 (N_1638,N_1152,N_1206);
or U1639 (N_1639,N_843,N_1327);
xor U1640 (N_1640,N_952,N_777);
nand U1641 (N_1641,N_996,N_1212);
and U1642 (N_1642,N_861,N_926);
xor U1643 (N_1643,N_1333,N_1030);
or U1644 (N_1644,N_1221,N_795);
xnor U1645 (N_1645,N_1158,N_1465);
or U1646 (N_1646,N_907,N_1278);
xor U1647 (N_1647,N_1258,N_1271);
nand U1648 (N_1648,N_783,N_1323);
or U1649 (N_1649,N_1389,N_1207);
nor U1650 (N_1650,N_1038,N_1244);
xnor U1651 (N_1651,N_957,N_1425);
and U1652 (N_1652,N_1392,N_1381);
xnor U1653 (N_1653,N_852,N_985);
and U1654 (N_1654,N_1228,N_1306);
nor U1655 (N_1655,N_1485,N_1322);
nand U1656 (N_1656,N_910,N_908);
xor U1657 (N_1657,N_831,N_1056);
xor U1658 (N_1658,N_1472,N_1276);
or U1659 (N_1659,N_938,N_1039);
and U1660 (N_1660,N_1295,N_869);
nor U1661 (N_1661,N_1016,N_1480);
xnor U1662 (N_1662,N_1264,N_1385);
and U1663 (N_1663,N_1438,N_1376);
or U1664 (N_1664,N_937,N_1411);
and U1665 (N_1665,N_1310,N_911);
nor U1666 (N_1666,N_1335,N_840);
nand U1667 (N_1667,N_887,N_836);
nand U1668 (N_1668,N_1393,N_889);
and U1669 (N_1669,N_855,N_1073);
and U1670 (N_1670,N_891,N_1454);
and U1671 (N_1671,N_1453,N_781);
nand U1672 (N_1672,N_1082,N_1302);
nor U1673 (N_1673,N_780,N_1001);
nand U1674 (N_1674,N_1127,N_1072);
and U1675 (N_1675,N_1443,N_1304);
or U1676 (N_1676,N_1236,N_978);
nand U1677 (N_1677,N_1113,N_839);
xor U1678 (N_1678,N_1076,N_846);
and U1679 (N_1679,N_1202,N_1128);
xor U1680 (N_1680,N_1096,N_1011);
and U1681 (N_1681,N_1277,N_924);
xor U1682 (N_1682,N_1169,N_1098);
nor U1683 (N_1683,N_1230,N_759);
xnor U1684 (N_1684,N_947,N_932);
nand U1685 (N_1685,N_754,N_1037);
nand U1686 (N_1686,N_1270,N_1291);
nor U1687 (N_1687,N_1185,N_798);
nor U1688 (N_1688,N_1122,N_1346);
nand U1689 (N_1689,N_1060,N_1343);
xor U1690 (N_1690,N_1242,N_882);
and U1691 (N_1691,N_828,N_864);
nand U1692 (N_1692,N_1178,N_1446);
or U1693 (N_1693,N_935,N_920);
and U1694 (N_1694,N_1495,N_1336);
nor U1695 (N_1695,N_1402,N_1469);
xor U1696 (N_1696,N_1269,N_838);
and U1697 (N_1697,N_866,N_1173);
or U1698 (N_1698,N_1048,N_787);
or U1699 (N_1699,N_1124,N_823);
and U1700 (N_1700,N_1033,N_1317);
nor U1701 (N_1701,N_1422,N_1186);
xor U1702 (N_1702,N_1188,N_1448);
nand U1703 (N_1703,N_1339,N_1191);
and U1704 (N_1704,N_1329,N_1175);
xor U1705 (N_1705,N_1210,N_1299);
xor U1706 (N_1706,N_873,N_1475);
xnor U1707 (N_1707,N_1086,N_1035);
and U1708 (N_1708,N_1430,N_1165);
xor U1709 (N_1709,N_1404,N_1179);
xnor U1710 (N_1710,N_1319,N_1036);
and U1711 (N_1711,N_1215,N_1140);
and U1712 (N_1712,N_1101,N_1196);
xnor U1713 (N_1713,N_1032,N_1403);
nand U1714 (N_1714,N_803,N_1220);
xor U1715 (N_1715,N_853,N_906);
nand U1716 (N_1716,N_1371,N_1396);
nor U1717 (N_1717,N_1320,N_1004);
nand U1718 (N_1718,N_1143,N_1459);
xnor U1719 (N_1719,N_1046,N_1253);
xor U1720 (N_1720,N_964,N_1142);
and U1721 (N_1721,N_1248,N_1348);
nand U1722 (N_1722,N_1104,N_751);
xnor U1723 (N_1723,N_792,N_1499);
nor U1724 (N_1724,N_1083,N_1241);
nand U1725 (N_1725,N_1377,N_1013);
or U1726 (N_1726,N_1400,N_1075);
or U1727 (N_1727,N_1497,N_1380);
nor U1728 (N_1728,N_1435,N_1476);
nand U1729 (N_1729,N_1150,N_771);
xnor U1730 (N_1730,N_1002,N_796);
xnor U1731 (N_1731,N_1455,N_1217);
and U1732 (N_1732,N_1180,N_895);
nand U1733 (N_1733,N_1161,N_1300);
xor U1734 (N_1734,N_841,N_1051);
xor U1735 (N_1735,N_1284,N_871);
and U1736 (N_1736,N_769,N_994);
and U1737 (N_1737,N_1144,N_800);
nand U1738 (N_1738,N_848,N_1470);
and U1739 (N_1739,N_888,N_1172);
nand U1740 (N_1740,N_799,N_936);
nand U1741 (N_1741,N_1181,N_1414);
or U1742 (N_1742,N_1042,N_1424);
xnor U1743 (N_1743,N_1292,N_854);
nor U1744 (N_1744,N_1452,N_1208);
or U1745 (N_1745,N_1356,N_877);
nor U1746 (N_1746,N_1468,N_1216);
xor U1747 (N_1747,N_1391,N_909);
nor U1748 (N_1748,N_1351,N_765);
nor U1749 (N_1749,N_1239,N_1246);
nor U1750 (N_1750,N_914,N_1368);
or U1751 (N_1751,N_1375,N_1369);
nor U1752 (N_1752,N_1025,N_788);
or U1753 (N_1753,N_844,N_1379);
nor U1754 (N_1754,N_1245,N_1412);
xnor U1755 (N_1755,N_1286,N_991);
nor U1756 (N_1756,N_786,N_757);
nor U1757 (N_1757,N_1397,N_1407);
nor U1758 (N_1758,N_1328,N_835);
nor U1759 (N_1759,N_775,N_961);
nor U1760 (N_1760,N_1462,N_1363);
and U1761 (N_1761,N_1314,N_1146);
nand U1762 (N_1762,N_1473,N_1069);
and U1763 (N_1763,N_791,N_1490);
nand U1764 (N_1764,N_1139,N_750);
xor U1765 (N_1765,N_1294,N_1022);
nand U1766 (N_1766,N_1166,N_1141);
xor U1767 (N_1767,N_944,N_1057);
nand U1768 (N_1768,N_782,N_1431);
or U1769 (N_1769,N_1108,N_1340);
xnor U1770 (N_1770,N_1266,N_756);
or U1771 (N_1771,N_1014,N_804);
and U1772 (N_1772,N_1131,N_1026);
nor U1773 (N_1773,N_1427,N_922);
nor U1774 (N_1774,N_982,N_1388);
or U1775 (N_1775,N_998,N_1214);
nor U1776 (N_1776,N_1251,N_1410);
nand U1777 (N_1777,N_1070,N_1354);
nand U1778 (N_1778,N_774,N_1138);
nand U1779 (N_1779,N_1474,N_1126);
xor U1780 (N_1780,N_1494,N_1034);
or U1781 (N_1781,N_872,N_1481);
nor U1782 (N_1782,N_1274,N_1005);
nor U1783 (N_1783,N_1384,N_956);
or U1784 (N_1784,N_1203,N_847);
nand U1785 (N_1785,N_1078,N_818);
xnor U1786 (N_1786,N_929,N_1386);
and U1787 (N_1787,N_1288,N_1164);
or U1788 (N_1788,N_1148,N_925);
and U1789 (N_1789,N_1451,N_1102);
nand U1790 (N_1790,N_793,N_1254);
xor U1791 (N_1791,N_806,N_1456);
or U1792 (N_1792,N_1219,N_1260);
nor U1793 (N_1793,N_1045,N_1315);
and U1794 (N_1794,N_1416,N_1281);
nand U1795 (N_1795,N_1021,N_1100);
nand U1796 (N_1796,N_1261,N_1020);
and U1797 (N_1797,N_1307,N_1330);
xor U1798 (N_1798,N_1109,N_1439);
nand U1799 (N_1799,N_878,N_758);
and U1800 (N_1800,N_1235,N_1374);
or U1801 (N_1801,N_1006,N_1189);
or U1802 (N_1802,N_797,N_1345);
and U1803 (N_1803,N_1418,N_1160);
or U1804 (N_1804,N_876,N_1089);
nand U1805 (N_1805,N_916,N_1357);
and U1806 (N_1806,N_1280,N_899);
nand U1807 (N_1807,N_1129,N_1305);
nor U1808 (N_1808,N_1478,N_801);
xnor U1809 (N_1809,N_1362,N_762);
xor U1810 (N_1810,N_1193,N_981);
and U1811 (N_1811,N_1313,N_1090);
or U1812 (N_1812,N_1009,N_1055);
nor U1813 (N_1813,N_1457,N_1471);
nor U1814 (N_1814,N_1137,N_1334);
or U1815 (N_1815,N_1308,N_1061);
nor U1816 (N_1816,N_1200,N_807);
xnor U1817 (N_1817,N_1252,N_1147);
nand U1818 (N_1818,N_1097,N_1460);
and U1819 (N_1819,N_967,N_808);
nand U1820 (N_1820,N_1347,N_1417);
xnor U1821 (N_1821,N_1395,N_919);
xor U1822 (N_1822,N_1434,N_1136);
nor U1823 (N_1823,N_1120,N_1123);
nor U1824 (N_1824,N_1382,N_1297);
and U1825 (N_1825,N_903,N_1156);
nor U1826 (N_1826,N_1226,N_1309);
and U1827 (N_1827,N_810,N_1201);
nor U1828 (N_1828,N_1440,N_966);
nor U1829 (N_1829,N_1268,N_923);
and U1830 (N_1830,N_1088,N_814);
nor U1831 (N_1831,N_870,N_1027);
xnor U1832 (N_1832,N_1296,N_1133);
or U1833 (N_1833,N_1000,N_1145);
nand U1834 (N_1834,N_1041,N_970);
and U1835 (N_1835,N_1373,N_789);
and U1836 (N_1836,N_1273,N_875);
nor U1837 (N_1837,N_1223,N_1484);
nand U1838 (N_1838,N_971,N_1437);
xnor U1839 (N_1839,N_1063,N_1121);
or U1840 (N_1840,N_1479,N_1182);
or U1841 (N_1841,N_1130,N_912);
and U1842 (N_1842,N_1444,N_988);
xor U1843 (N_1843,N_1259,N_1049);
nand U1844 (N_1844,N_1358,N_941);
nor U1845 (N_1845,N_1190,N_1153);
or U1846 (N_1846,N_939,N_897);
or U1847 (N_1847,N_1040,N_1053);
nand U1848 (N_1848,N_1125,N_1445);
xor U1849 (N_1849,N_1449,N_784);
nand U1850 (N_1850,N_1466,N_986);
and U1851 (N_1851,N_849,N_1255);
nor U1852 (N_1852,N_817,N_1409);
nand U1853 (N_1853,N_890,N_963);
or U1854 (N_1854,N_1115,N_830);
xor U1855 (N_1855,N_968,N_977);
xor U1856 (N_1856,N_858,N_842);
xor U1857 (N_1857,N_1028,N_1168);
nand U1858 (N_1858,N_1170,N_885);
nor U1859 (N_1859,N_997,N_832);
nand U1860 (N_1860,N_752,N_1114);
nand U1861 (N_1861,N_755,N_834);
and U1862 (N_1862,N_1084,N_1155);
or U1863 (N_1863,N_1399,N_881);
or U1864 (N_1864,N_829,N_1387);
xor U1865 (N_1865,N_1415,N_1067);
or U1866 (N_1866,N_918,N_884);
xor U1867 (N_1867,N_1257,N_948);
xor U1868 (N_1868,N_1405,N_867);
nor U1869 (N_1869,N_1093,N_1243);
nor U1870 (N_1870,N_917,N_1218);
and U1871 (N_1871,N_1080,N_1325);
xnor U1872 (N_1872,N_773,N_779);
and U1873 (N_1873,N_1341,N_1018);
and U1874 (N_1874,N_1262,N_1222);
and U1875 (N_1875,N_1005,N_885);
xor U1876 (N_1876,N_1308,N_776);
nor U1877 (N_1877,N_1172,N_793);
and U1878 (N_1878,N_1444,N_900);
or U1879 (N_1879,N_824,N_1309);
xor U1880 (N_1880,N_1308,N_792);
or U1881 (N_1881,N_883,N_1406);
nor U1882 (N_1882,N_1480,N_1021);
xnor U1883 (N_1883,N_775,N_930);
or U1884 (N_1884,N_791,N_1208);
xor U1885 (N_1885,N_1210,N_1418);
nor U1886 (N_1886,N_1230,N_1009);
or U1887 (N_1887,N_860,N_851);
and U1888 (N_1888,N_1033,N_764);
or U1889 (N_1889,N_1025,N_1330);
xnor U1890 (N_1890,N_1179,N_988);
xor U1891 (N_1891,N_1252,N_1286);
and U1892 (N_1892,N_1409,N_1255);
and U1893 (N_1893,N_1342,N_1221);
nand U1894 (N_1894,N_1426,N_1117);
xnor U1895 (N_1895,N_1340,N_1320);
xnor U1896 (N_1896,N_858,N_937);
nand U1897 (N_1897,N_926,N_1010);
or U1898 (N_1898,N_1315,N_1350);
nand U1899 (N_1899,N_888,N_1422);
nand U1900 (N_1900,N_1268,N_988);
and U1901 (N_1901,N_1443,N_923);
nor U1902 (N_1902,N_1459,N_934);
or U1903 (N_1903,N_1033,N_848);
xnor U1904 (N_1904,N_1385,N_1008);
nand U1905 (N_1905,N_1375,N_807);
and U1906 (N_1906,N_769,N_900);
or U1907 (N_1907,N_961,N_854);
or U1908 (N_1908,N_1141,N_920);
xor U1909 (N_1909,N_784,N_1155);
xnor U1910 (N_1910,N_1179,N_1086);
or U1911 (N_1911,N_988,N_1247);
and U1912 (N_1912,N_1483,N_1270);
nor U1913 (N_1913,N_1293,N_1447);
nor U1914 (N_1914,N_1455,N_1107);
nand U1915 (N_1915,N_924,N_755);
nand U1916 (N_1916,N_1365,N_1222);
nand U1917 (N_1917,N_847,N_1270);
and U1918 (N_1918,N_937,N_921);
xor U1919 (N_1919,N_1194,N_1089);
or U1920 (N_1920,N_890,N_1204);
nand U1921 (N_1921,N_1213,N_1448);
nand U1922 (N_1922,N_948,N_1091);
and U1923 (N_1923,N_1130,N_1325);
nor U1924 (N_1924,N_893,N_1073);
nor U1925 (N_1925,N_999,N_894);
nand U1926 (N_1926,N_1144,N_1297);
xor U1927 (N_1927,N_1059,N_1398);
nor U1928 (N_1928,N_927,N_1218);
xnor U1929 (N_1929,N_1364,N_1176);
and U1930 (N_1930,N_1358,N_979);
and U1931 (N_1931,N_755,N_1130);
xor U1932 (N_1932,N_1164,N_1456);
or U1933 (N_1933,N_1410,N_825);
nand U1934 (N_1934,N_1453,N_1301);
xor U1935 (N_1935,N_1272,N_1263);
and U1936 (N_1936,N_987,N_1259);
nor U1937 (N_1937,N_1373,N_760);
nand U1938 (N_1938,N_1349,N_1381);
nand U1939 (N_1939,N_1299,N_1445);
and U1940 (N_1940,N_900,N_1380);
or U1941 (N_1941,N_862,N_1230);
and U1942 (N_1942,N_1049,N_1412);
xnor U1943 (N_1943,N_1071,N_1089);
or U1944 (N_1944,N_1082,N_1266);
nand U1945 (N_1945,N_1184,N_852);
xor U1946 (N_1946,N_1056,N_756);
or U1947 (N_1947,N_1325,N_1219);
nor U1948 (N_1948,N_1445,N_1066);
and U1949 (N_1949,N_1317,N_1238);
or U1950 (N_1950,N_1307,N_1369);
xor U1951 (N_1951,N_754,N_1307);
nor U1952 (N_1952,N_1240,N_1196);
xor U1953 (N_1953,N_1487,N_1031);
and U1954 (N_1954,N_1345,N_995);
nand U1955 (N_1955,N_1026,N_782);
nand U1956 (N_1956,N_883,N_1458);
xnor U1957 (N_1957,N_807,N_979);
xnor U1958 (N_1958,N_1328,N_1364);
or U1959 (N_1959,N_833,N_1481);
and U1960 (N_1960,N_1358,N_789);
nor U1961 (N_1961,N_1302,N_999);
nand U1962 (N_1962,N_849,N_1260);
nand U1963 (N_1963,N_1026,N_1214);
nor U1964 (N_1964,N_1099,N_812);
and U1965 (N_1965,N_1214,N_810);
and U1966 (N_1966,N_1329,N_1100);
or U1967 (N_1967,N_1243,N_1233);
and U1968 (N_1968,N_933,N_975);
and U1969 (N_1969,N_1331,N_1269);
nand U1970 (N_1970,N_876,N_1100);
nor U1971 (N_1971,N_1137,N_1013);
or U1972 (N_1972,N_1494,N_1296);
and U1973 (N_1973,N_1082,N_795);
or U1974 (N_1974,N_1036,N_1252);
and U1975 (N_1975,N_1402,N_1235);
nor U1976 (N_1976,N_1481,N_936);
and U1977 (N_1977,N_883,N_868);
or U1978 (N_1978,N_1133,N_1222);
or U1979 (N_1979,N_1064,N_1347);
nand U1980 (N_1980,N_1169,N_754);
and U1981 (N_1981,N_1210,N_1457);
xor U1982 (N_1982,N_829,N_1112);
nor U1983 (N_1983,N_1021,N_799);
and U1984 (N_1984,N_888,N_1389);
xor U1985 (N_1985,N_1312,N_1060);
and U1986 (N_1986,N_991,N_1340);
or U1987 (N_1987,N_1249,N_1478);
nor U1988 (N_1988,N_974,N_944);
and U1989 (N_1989,N_925,N_1292);
xnor U1990 (N_1990,N_1304,N_980);
xor U1991 (N_1991,N_971,N_1315);
or U1992 (N_1992,N_911,N_1353);
nand U1993 (N_1993,N_1290,N_758);
or U1994 (N_1994,N_1382,N_834);
xnor U1995 (N_1995,N_1019,N_840);
or U1996 (N_1996,N_1059,N_861);
nor U1997 (N_1997,N_925,N_1320);
xor U1998 (N_1998,N_1483,N_834);
xor U1999 (N_1999,N_1048,N_1155);
nand U2000 (N_2000,N_1421,N_1113);
nand U2001 (N_2001,N_809,N_1290);
nor U2002 (N_2002,N_1032,N_1061);
or U2003 (N_2003,N_971,N_809);
nand U2004 (N_2004,N_1117,N_1083);
and U2005 (N_2005,N_925,N_1080);
and U2006 (N_2006,N_1083,N_933);
and U2007 (N_2007,N_951,N_1047);
xnor U2008 (N_2008,N_979,N_933);
or U2009 (N_2009,N_1098,N_1154);
or U2010 (N_2010,N_1228,N_1078);
xnor U2011 (N_2011,N_1078,N_770);
xnor U2012 (N_2012,N_1208,N_1354);
nor U2013 (N_2013,N_1480,N_822);
xor U2014 (N_2014,N_1294,N_950);
or U2015 (N_2015,N_1391,N_915);
or U2016 (N_2016,N_1056,N_1198);
xor U2017 (N_2017,N_866,N_1376);
nor U2018 (N_2018,N_1460,N_1017);
and U2019 (N_2019,N_863,N_1106);
or U2020 (N_2020,N_1005,N_1000);
nor U2021 (N_2021,N_1157,N_771);
or U2022 (N_2022,N_1098,N_1486);
nor U2023 (N_2023,N_1086,N_1287);
nand U2024 (N_2024,N_853,N_1488);
xor U2025 (N_2025,N_885,N_772);
and U2026 (N_2026,N_1451,N_1294);
and U2027 (N_2027,N_1015,N_834);
xor U2028 (N_2028,N_1316,N_857);
or U2029 (N_2029,N_1079,N_809);
nor U2030 (N_2030,N_799,N_1077);
or U2031 (N_2031,N_1400,N_1074);
or U2032 (N_2032,N_1035,N_924);
xnor U2033 (N_2033,N_911,N_1229);
nor U2034 (N_2034,N_1085,N_792);
nor U2035 (N_2035,N_1395,N_1275);
nand U2036 (N_2036,N_765,N_784);
or U2037 (N_2037,N_1225,N_754);
nand U2038 (N_2038,N_1487,N_1443);
nand U2039 (N_2039,N_1150,N_1284);
xnor U2040 (N_2040,N_958,N_995);
xor U2041 (N_2041,N_1019,N_937);
or U2042 (N_2042,N_1322,N_898);
nand U2043 (N_2043,N_842,N_1306);
nor U2044 (N_2044,N_1407,N_1336);
xnor U2045 (N_2045,N_779,N_968);
nor U2046 (N_2046,N_996,N_1121);
xor U2047 (N_2047,N_895,N_832);
and U2048 (N_2048,N_876,N_1073);
nor U2049 (N_2049,N_1414,N_992);
xor U2050 (N_2050,N_771,N_1086);
or U2051 (N_2051,N_987,N_1168);
or U2052 (N_2052,N_755,N_1006);
and U2053 (N_2053,N_1188,N_1202);
nor U2054 (N_2054,N_776,N_1037);
xnor U2055 (N_2055,N_1245,N_825);
xnor U2056 (N_2056,N_872,N_1091);
or U2057 (N_2057,N_1096,N_1230);
nor U2058 (N_2058,N_935,N_1469);
or U2059 (N_2059,N_1159,N_1397);
nand U2060 (N_2060,N_899,N_1335);
xor U2061 (N_2061,N_1284,N_976);
or U2062 (N_2062,N_929,N_1260);
or U2063 (N_2063,N_1048,N_1485);
xnor U2064 (N_2064,N_1423,N_915);
nor U2065 (N_2065,N_877,N_1184);
xor U2066 (N_2066,N_1129,N_1344);
or U2067 (N_2067,N_1090,N_1029);
nor U2068 (N_2068,N_962,N_1162);
xnor U2069 (N_2069,N_940,N_993);
nor U2070 (N_2070,N_1356,N_1324);
or U2071 (N_2071,N_903,N_1232);
nand U2072 (N_2072,N_879,N_807);
and U2073 (N_2073,N_1406,N_1313);
or U2074 (N_2074,N_1173,N_1408);
nor U2075 (N_2075,N_873,N_1427);
and U2076 (N_2076,N_1436,N_1451);
xnor U2077 (N_2077,N_1221,N_1334);
xnor U2078 (N_2078,N_1172,N_960);
xnor U2079 (N_2079,N_1400,N_831);
nor U2080 (N_2080,N_1217,N_1257);
nand U2081 (N_2081,N_890,N_1071);
nor U2082 (N_2082,N_827,N_781);
or U2083 (N_2083,N_911,N_968);
xor U2084 (N_2084,N_1275,N_1342);
nand U2085 (N_2085,N_1293,N_811);
or U2086 (N_2086,N_1326,N_1416);
nand U2087 (N_2087,N_984,N_1011);
and U2088 (N_2088,N_1148,N_789);
nor U2089 (N_2089,N_882,N_1017);
nand U2090 (N_2090,N_913,N_1223);
or U2091 (N_2091,N_806,N_891);
xnor U2092 (N_2092,N_765,N_934);
and U2093 (N_2093,N_799,N_1062);
xnor U2094 (N_2094,N_951,N_1010);
or U2095 (N_2095,N_1046,N_1346);
or U2096 (N_2096,N_1022,N_822);
or U2097 (N_2097,N_1144,N_1467);
nand U2098 (N_2098,N_972,N_759);
and U2099 (N_2099,N_829,N_1221);
or U2100 (N_2100,N_1044,N_1402);
nor U2101 (N_2101,N_1300,N_798);
or U2102 (N_2102,N_1333,N_1340);
and U2103 (N_2103,N_1089,N_1316);
nor U2104 (N_2104,N_931,N_1047);
nor U2105 (N_2105,N_1099,N_1469);
and U2106 (N_2106,N_1056,N_986);
xnor U2107 (N_2107,N_1043,N_1037);
nand U2108 (N_2108,N_1009,N_1395);
nand U2109 (N_2109,N_1173,N_927);
xnor U2110 (N_2110,N_1288,N_833);
nor U2111 (N_2111,N_1175,N_1299);
nand U2112 (N_2112,N_958,N_888);
nor U2113 (N_2113,N_1275,N_1252);
nand U2114 (N_2114,N_1104,N_1188);
and U2115 (N_2115,N_1130,N_1100);
xnor U2116 (N_2116,N_1092,N_1097);
and U2117 (N_2117,N_1413,N_1032);
xor U2118 (N_2118,N_961,N_787);
nor U2119 (N_2119,N_943,N_752);
nor U2120 (N_2120,N_1099,N_1059);
nor U2121 (N_2121,N_1171,N_991);
or U2122 (N_2122,N_1178,N_966);
xnor U2123 (N_2123,N_1167,N_1408);
nor U2124 (N_2124,N_1455,N_776);
nor U2125 (N_2125,N_1455,N_1085);
xnor U2126 (N_2126,N_1195,N_1221);
nand U2127 (N_2127,N_996,N_1097);
nand U2128 (N_2128,N_786,N_1417);
and U2129 (N_2129,N_1043,N_1166);
nor U2130 (N_2130,N_917,N_1458);
nand U2131 (N_2131,N_1403,N_1029);
nand U2132 (N_2132,N_1420,N_894);
nor U2133 (N_2133,N_1451,N_985);
or U2134 (N_2134,N_832,N_1215);
and U2135 (N_2135,N_1254,N_901);
nor U2136 (N_2136,N_1368,N_1361);
xnor U2137 (N_2137,N_808,N_1210);
xor U2138 (N_2138,N_858,N_1484);
or U2139 (N_2139,N_857,N_1440);
nand U2140 (N_2140,N_876,N_1026);
nor U2141 (N_2141,N_1234,N_888);
and U2142 (N_2142,N_1231,N_1201);
nand U2143 (N_2143,N_1386,N_1071);
xor U2144 (N_2144,N_792,N_1028);
or U2145 (N_2145,N_753,N_1058);
and U2146 (N_2146,N_1316,N_1253);
and U2147 (N_2147,N_1139,N_807);
xnor U2148 (N_2148,N_866,N_1252);
nor U2149 (N_2149,N_1368,N_1206);
nand U2150 (N_2150,N_1192,N_1352);
nand U2151 (N_2151,N_856,N_890);
and U2152 (N_2152,N_1316,N_1293);
or U2153 (N_2153,N_1176,N_836);
nor U2154 (N_2154,N_1247,N_861);
and U2155 (N_2155,N_1359,N_1165);
nor U2156 (N_2156,N_1377,N_1064);
and U2157 (N_2157,N_1289,N_893);
or U2158 (N_2158,N_1003,N_1147);
nor U2159 (N_2159,N_1301,N_880);
and U2160 (N_2160,N_1145,N_1379);
nand U2161 (N_2161,N_1183,N_1402);
and U2162 (N_2162,N_1485,N_1054);
or U2163 (N_2163,N_1345,N_1222);
nor U2164 (N_2164,N_1022,N_1187);
or U2165 (N_2165,N_1353,N_1392);
nor U2166 (N_2166,N_922,N_1355);
nand U2167 (N_2167,N_862,N_854);
and U2168 (N_2168,N_1375,N_1190);
or U2169 (N_2169,N_1055,N_1026);
xnor U2170 (N_2170,N_1152,N_1125);
xnor U2171 (N_2171,N_1275,N_957);
nand U2172 (N_2172,N_872,N_922);
xor U2173 (N_2173,N_896,N_1167);
nor U2174 (N_2174,N_989,N_1075);
or U2175 (N_2175,N_832,N_1189);
nor U2176 (N_2176,N_844,N_822);
xor U2177 (N_2177,N_1476,N_1120);
xor U2178 (N_2178,N_1344,N_1189);
nand U2179 (N_2179,N_1380,N_1018);
nand U2180 (N_2180,N_1044,N_782);
and U2181 (N_2181,N_1204,N_1297);
nor U2182 (N_2182,N_757,N_1427);
and U2183 (N_2183,N_1425,N_864);
or U2184 (N_2184,N_978,N_977);
and U2185 (N_2185,N_1365,N_1351);
or U2186 (N_2186,N_849,N_1126);
nand U2187 (N_2187,N_1063,N_1416);
nor U2188 (N_2188,N_1002,N_1237);
xor U2189 (N_2189,N_932,N_1234);
xor U2190 (N_2190,N_1001,N_1126);
and U2191 (N_2191,N_1217,N_932);
or U2192 (N_2192,N_868,N_1343);
and U2193 (N_2193,N_1473,N_998);
xor U2194 (N_2194,N_1398,N_994);
and U2195 (N_2195,N_1333,N_1200);
and U2196 (N_2196,N_1046,N_1488);
nand U2197 (N_2197,N_1493,N_1393);
xnor U2198 (N_2198,N_1440,N_870);
xnor U2199 (N_2199,N_1244,N_922);
nand U2200 (N_2200,N_1304,N_1250);
and U2201 (N_2201,N_1097,N_1457);
xor U2202 (N_2202,N_1326,N_1200);
or U2203 (N_2203,N_998,N_901);
nor U2204 (N_2204,N_897,N_1075);
nand U2205 (N_2205,N_819,N_1227);
and U2206 (N_2206,N_1073,N_812);
or U2207 (N_2207,N_1229,N_809);
nand U2208 (N_2208,N_862,N_963);
nand U2209 (N_2209,N_1237,N_1348);
or U2210 (N_2210,N_1095,N_1085);
and U2211 (N_2211,N_901,N_1338);
nand U2212 (N_2212,N_1317,N_1418);
nand U2213 (N_2213,N_841,N_843);
nand U2214 (N_2214,N_1428,N_1046);
or U2215 (N_2215,N_1087,N_1355);
or U2216 (N_2216,N_934,N_1068);
nor U2217 (N_2217,N_1249,N_1062);
xor U2218 (N_2218,N_1308,N_1259);
and U2219 (N_2219,N_1045,N_835);
nand U2220 (N_2220,N_795,N_890);
and U2221 (N_2221,N_1394,N_1292);
nand U2222 (N_2222,N_1493,N_800);
nor U2223 (N_2223,N_1466,N_1154);
or U2224 (N_2224,N_1033,N_928);
and U2225 (N_2225,N_976,N_1274);
xor U2226 (N_2226,N_841,N_791);
nor U2227 (N_2227,N_832,N_1091);
or U2228 (N_2228,N_1268,N_1076);
and U2229 (N_2229,N_1435,N_932);
and U2230 (N_2230,N_1064,N_1178);
and U2231 (N_2231,N_1197,N_1195);
xnor U2232 (N_2232,N_867,N_1426);
or U2233 (N_2233,N_1137,N_986);
or U2234 (N_2234,N_1353,N_1465);
nand U2235 (N_2235,N_1039,N_1411);
and U2236 (N_2236,N_1225,N_1487);
nand U2237 (N_2237,N_1338,N_1074);
and U2238 (N_2238,N_1240,N_1350);
or U2239 (N_2239,N_1257,N_1176);
xor U2240 (N_2240,N_1183,N_1140);
or U2241 (N_2241,N_1182,N_1460);
xor U2242 (N_2242,N_1239,N_1260);
nor U2243 (N_2243,N_1306,N_1230);
and U2244 (N_2244,N_768,N_1332);
nand U2245 (N_2245,N_1409,N_938);
nand U2246 (N_2246,N_933,N_1369);
xor U2247 (N_2247,N_1226,N_1233);
xnor U2248 (N_2248,N_1029,N_1431);
nor U2249 (N_2249,N_806,N_1340);
and U2250 (N_2250,N_2011,N_1834);
nor U2251 (N_2251,N_1809,N_1547);
or U2252 (N_2252,N_1561,N_1802);
or U2253 (N_2253,N_1540,N_1875);
and U2254 (N_2254,N_2203,N_1947);
and U2255 (N_2255,N_2165,N_2192);
nand U2256 (N_2256,N_2233,N_1510);
and U2257 (N_2257,N_1535,N_2062);
or U2258 (N_2258,N_2018,N_1543);
nand U2259 (N_2259,N_1603,N_1639);
and U2260 (N_2260,N_2071,N_1849);
nand U2261 (N_2261,N_1913,N_1766);
or U2262 (N_2262,N_1563,N_1537);
nor U2263 (N_2263,N_1974,N_1773);
or U2264 (N_2264,N_2221,N_1881);
nor U2265 (N_2265,N_1523,N_1858);
nor U2266 (N_2266,N_1565,N_1631);
xor U2267 (N_2267,N_1978,N_1894);
nor U2268 (N_2268,N_2040,N_2241);
or U2269 (N_2269,N_2019,N_1811);
nand U2270 (N_2270,N_1599,N_1711);
xnor U2271 (N_2271,N_1911,N_1666);
and U2272 (N_2272,N_1677,N_2180);
nor U2273 (N_2273,N_1892,N_1519);
nor U2274 (N_2274,N_1800,N_1676);
nand U2275 (N_2275,N_2125,N_1832);
xnor U2276 (N_2276,N_1693,N_1774);
and U2277 (N_2277,N_2219,N_2127);
xnor U2278 (N_2278,N_2081,N_1979);
xnor U2279 (N_2279,N_1816,N_2074);
nor U2280 (N_2280,N_1899,N_1943);
and U2281 (N_2281,N_1727,N_1756);
and U2282 (N_2282,N_2025,N_1648);
nor U2283 (N_2283,N_1514,N_1709);
nor U2284 (N_2284,N_1882,N_1734);
nand U2285 (N_2285,N_1532,N_1889);
xor U2286 (N_2286,N_1931,N_2089);
xnor U2287 (N_2287,N_1571,N_1655);
or U2288 (N_2288,N_2128,N_2001);
or U2289 (N_2289,N_1914,N_2190);
or U2290 (N_2290,N_1819,N_1524);
nand U2291 (N_2291,N_2187,N_2134);
nor U2292 (N_2292,N_1966,N_2045);
nor U2293 (N_2293,N_1794,N_2055);
xnor U2294 (N_2294,N_1907,N_2120);
or U2295 (N_2295,N_2207,N_2100);
nand U2296 (N_2296,N_1691,N_1526);
nand U2297 (N_2297,N_2141,N_1634);
nand U2298 (N_2298,N_1778,N_1873);
or U2299 (N_2299,N_1912,N_2114);
or U2300 (N_2300,N_1705,N_1527);
or U2301 (N_2301,N_1653,N_1877);
nor U2302 (N_2302,N_1857,N_1845);
and U2303 (N_2303,N_2247,N_1829);
or U2304 (N_2304,N_2131,N_1923);
xor U2305 (N_2305,N_1684,N_1716);
nor U2306 (N_2306,N_1635,N_1638);
or U2307 (N_2307,N_1598,N_2143);
nand U2308 (N_2308,N_2158,N_2068);
xnor U2309 (N_2309,N_1939,N_1852);
xnor U2310 (N_2310,N_1826,N_2046);
nor U2311 (N_2311,N_1654,N_2079);
or U2312 (N_2312,N_2249,N_1995);
nor U2313 (N_2313,N_2237,N_2231);
xor U2314 (N_2314,N_2196,N_1799);
xnor U2315 (N_2315,N_2216,N_1950);
xor U2316 (N_2316,N_2234,N_2013);
and U2317 (N_2317,N_1708,N_1812);
and U2318 (N_2318,N_1506,N_1577);
and U2319 (N_2319,N_2033,N_1515);
xor U2320 (N_2320,N_1872,N_1968);
nor U2321 (N_2321,N_1970,N_2174);
nor U2322 (N_2322,N_1539,N_2063);
or U2323 (N_2323,N_1567,N_1851);
nor U2324 (N_2324,N_1536,N_2113);
and U2325 (N_2325,N_2050,N_1868);
and U2326 (N_2326,N_1604,N_1895);
xnor U2327 (N_2327,N_1742,N_1793);
and U2328 (N_2328,N_2155,N_1859);
nor U2329 (N_2329,N_1694,N_1879);
nand U2330 (N_2330,N_1797,N_1745);
nand U2331 (N_2331,N_2172,N_1548);
or U2332 (N_2332,N_1623,N_1674);
and U2333 (N_2333,N_1695,N_2194);
xnor U2334 (N_2334,N_2225,N_2191);
nor U2335 (N_2335,N_2167,N_2154);
xor U2336 (N_2336,N_2137,N_2181);
nor U2337 (N_2337,N_2210,N_2092);
nand U2338 (N_2338,N_1673,N_2088);
or U2339 (N_2339,N_1600,N_1521);
or U2340 (N_2340,N_2006,N_1863);
nor U2341 (N_2341,N_2135,N_2130);
nand U2342 (N_2342,N_1976,N_1622);
or U2343 (N_2343,N_1870,N_1888);
and U2344 (N_2344,N_1739,N_1737);
nor U2345 (N_2345,N_2205,N_2099);
or U2346 (N_2346,N_2177,N_1568);
nand U2347 (N_2347,N_1721,N_1828);
and U2348 (N_2348,N_1796,N_2093);
nand U2349 (N_2349,N_1779,N_2198);
or U2350 (N_2350,N_1722,N_1746);
xor U2351 (N_2351,N_2182,N_2080);
nor U2352 (N_2352,N_1781,N_1838);
and U2353 (N_2353,N_1720,N_2124);
nand U2354 (N_2354,N_1592,N_2026);
nor U2355 (N_2355,N_2035,N_2168);
xnor U2356 (N_2356,N_2076,N_1841);
or U2357 (N_2357,N_1618,N_2206);
or U2358 (N_2358,N_1696,N_2094);
nand U2359 (N_2359,N_2160,N_1637);
xnor U2360 (N_2360,N_2054,N_1699);
or U2361 (N_2361,N_1730,N_1546);
xnor U2362 (N_2362,N_2103,N_2204);
and U2363 (N_2363,N_1560,N_1953);
xor U2364 (N_2364,N_2086,N_1701);
or U2365 (N_2365,N_1559,N_1712);
xnor U2366 (N_2366,N_1844,N_1996);
nor U2367 (N_2367,N_1955,N_1780);
or U2368 (N_2368,N_2214,N_1817);
xnor U2369 (N_2369,N_1919,N_1957);
xor U2370 (N_2370,N_1962,N_1807);
or U2371 (N_2371,N_1702,N_1723);
nand U2372 (N_2372,N_1507,N_1847);
xnor U2373 (N_2373,N_1810,N_2090);
xor U2374 (N_2374,N_1920,N_2148);
nor U2375 (N_2375,N_1752,N_1554);
nor U2376 (N_2376,N_2039,N_2075);
nor U2377 (N_2377,N_1516,N_1835);
or U2378 (N_2378,N_1650,N_1736);
xor U2379 (N_2379,N_1997,N_1596);
or U2380 (N_2380,N_1659,N_1893);
and U2381 (N_2381,N_1704,N_2162);
xor U2382 (N_2382,N_2049,N_2215);
xnor U2383 (N_2383,N_2059,N_1961);
nand U2384 (N_2384,N_1967,N_1531);
xor U2385 (N_2385,N_2029,N_1985);
nor U2386 (N_2386,N_2188,N_1934);
xnor U2387 (N_2387,N_1628,N_1775);
nor U2388 (N_2388,N_1710,N_1751);
xnor U2389 (N_2389,N_1612,N_1761);
xor U2390 (N_2390,N_1770,N_2101);
xnor U2391 (N_2391,N_2183,N_2157);
nand U2392 (N_2392,N_1517,N_1789);
xor U2393 (N_2393,N_1856,N_1665);
nand U2394 (N_2394,N_2023,N_2171);
and U2395 (N_2395,N_1508,N_1593);
and U2396 (N_2396,N_1777,N_1795);
nor U2397 (N_2397,N_2139,N_1725);
and U2398 (N_2398,N_1549,N_1602);
xor U2399 (N_2399,N_2052,N_1876);
xnor U2400 (N_2400,N_1700,N_1741);
or U2401 (N_2401,N_2122,N_1509);
or U2402 (N_2402,N_2057,N_1581);
nand U2403 (N_2403,N_1784,N_1715);
xor U2404 (N_2404,N_1830,N_2179);
and U2405 (N_2405,N_1994,N_1848);
nor U2406 (N_2406,N_2002,N_1839);
nor U2407 (N_2407,N_2084,N_2056);
nor U2408 (N_2408,N_2236,N_2043);
and U2409 (N_2409,N_1959,N_1647);
or U2410 (N_2410,N_1884,N_1971);
nand U2411 (N_2411,N_2217,N_1550);
nand U2412 (N_2412,N_1556,N_2149);
nor U2413 (N_2413,N_2146,N_2087);
xnor U2414 (N_2414,N_2243,N_1606);
nand U2415 (N_2415,N_1890,N_2041);
nor U2416 (N_2416,N_1946,N_1866);
nor U2417 (N_2417,N_2201,N_2166);
nor U2418 (N_2418,N_1505,N_1867);
and U2419 (N_2419,N_1552,N_1644);
or U2420 (N_2420,N_2132,N_2021);
nor U2421 (N_2421,N_1649,N_1625);
or U2422 (N_2422,N_1749,N_1754);
xor U2423 (N_2423,N_1590,N_1977);
nor U2424 (N_2424,N_1587,N_2119);
xnor U2425 (N_2425,N_1748,N_1679);
xor U2426 (N_2426,N_2105,N_1733);
nand U2427 (N_2427,N_1986,N_1818);
nand U2428 (N_2428,N_1886,N_1764);
and U2429 (N_2429,N_2108,N_2032);
or U2430 (N_2430,N_1763,N_2042);
or U2431 (N_2431,N_1806,N_2095);
xor U2432 (N_2432,N_2235,N_2170);
and U2433 (N_2433,N_2230,N_1878);
and U2434 (N_2434,N_1572,N_1518);
and U2435 (N_2435,N_2010,N_2005);
nor U2436 (N_2436,N_2051,N_1591);
or U2437 (N_2437,N_1898,N_2218);
xor U2438 (N_2438,N_1940,N_2212);
or U2439 (N_2439,N_2195,N_1573);
nand U2440 (N_2440,N_1740,N_1883);
and U2441 (N_2441,N_1902,N_1897);
nor U2442 (N_2442,N_1597,N_2111);
nand U2443 (N_2443,N_1688,N_2227);
nand U2444 (N_2444,N_1562,N_1891);
and U2445 (N_2445,N_2185,N_1703);
nor U2446 (N_2446,N_1904,N_2102);
and U2447 (N_2447,N_1626,N_1588);
xor U2448 (N_2448,N_2015,N_1951);
xnor U2449 (N_2449,N_1909,N_2176);
nor U2450 (N_2450,N_2121,N_1735);
and U2451 (N_2451,N_1831,N_1580);
nor U2452 (N_2452,N_1714,N_1726);
nand U2453 (N_2453,N_2069,N_1854);
or U2454 (N_2454,N_2159,N_1991);
or U2455 (N_2455,N_2030,N_2224);
nand U2456 (N_2456,N_1900,N_1956);
nor U2457 (N_2457,N_2016,N_1993);
and U2458 (N_2458,N_1935,N_2144);
xnor U2459 (N_2459,N_1570,N_2096);
nor U2460 (N_2460,N_1885,N_1713);
nor U2461 (N_2461,N_1594,N_1564);
or U2462 (N_2462,N_2014,N_2009);
nor U2463 (N_2463,N_1732,N_1855);
and U2464 (N_2464,N_1724,N_1840);
xor U2465 (N_2465,N_1617,N_1982);
or U2466 (N_2466,N_1689,N_2228);
nand U2467 (N_2467,N_1758,N_1698);
xor U2468 (N_2468,N_2061,N_1528);
and U2469 (N_2469,N_1706,N_1621);
nand U2470 (N_2470,N_1964,N_2020);
and U2471 (N_2471,N_2048,N_2008);
nand U2472 (N_2472,N_2150,N_1921);
nor U2473 (N_2473,N_1942,N_2085);
xor U2474 (N_2474,N_1553,N_2145);
or U2475 (N_2475,N_2110,N_1948);
xnor U2476 (N_2476,N_1928,N_2000);
nand U2477 (N_2477,N_1916,N_2138);
nand U2478 (N_2478,N_1944,N_2242);
nor U2479 (N_2479,N_2058,N_2133);
nor U2480 (N_2480,N_1960,N_2065);
nand U2481 (N_2481,N_1887,N_2106);
nor U2482 (N_2482,N_1798,N_2036);
nand U2483 (N_2483,N_2116,N_1813);
or U2484 (N_2484,N_1788,N_1999);
and U2485 (N_2485,N_1584,N_2213);
and U2486 (N_2486,N_2034,N_2064);
and U2487 (N_2487,N_1901,N_2175);
or U2488 (N_2488,N_1690,N_2173);
nor U2489 (N_2489,N_2047,N_1992);
nand U2490 (N_2490,N_1717,N_1915);
and U2491 (N_2491,N_1760,N_1757);
xor U2492 (N_2492,N_1922,N_2078);
xnor U2493 (N_2493,N_2017,N_1786);
and U2494 (N_2494,N_1566,N_1640);
or U2495 (N_2495,N_2117,N_1808);
or U2496 (N_2496,N_2199,N_2140);
and U2497 (N_2497,N_1759,N_1729);
xnor U2498 (N_2498,N_1504,N_1685);
xor U2499 (N_2499,N_1896,N_1719);
nand U2500 (N_2500,N_1989,N_1513);
nand U2501 (N_2501,N_1678,N_2072);
or U2502 (N_2502,N_2186,N_1917);
nor U2503 (N_2503,N_1769,N_1614);
or U2504 (N_2504,N_1657,N_1538);
xor U2505 (N_2505,N_2027,N_1557);
and U2506 (N_2506,N_2248,N_1541);
nand U2507 (N_2507,N_1718,N_2022);
and U2508 (N_2508,N_1670,N_2164);
xnor U2509 (N_2509,N_1743,N_1667);
xor U2510 (N_2510,N_1824,N_1608);
or U2511 (N_2511,N_1972,N_1501);
nand U2512 (N_2512,N_1833,N_2060);
and U2513 (N_2513,N_2142,N_1925);
and U2514 (N_2514,N_1975,N_2044);
and U2515 (N_2515,N_1980,N_1785);
or U2516 (N_2516,N_2244,N_2151);
xnor U2517 (N_2517,N_2129,N_1983);
xor U2518 (N_2518,N_1932,N_1776);
xnor U2519 (N_2519,N_1990,N_1579);
nand U2520 (N_2520,N_1620,N_1927);
nand U2521 (N_2521,N_1707,N_1952);
and U2522 (N_2522,N_1503,N_2037);
nor U2523 (N_2523,N_1762,N_1869);
or U2524 (N_2524,N_2097,N_2238);
or U2525 (N_2525,N_1998,N_2082);
nor U2526 (N_2526,N_1929,N_2126);
nand U2527 (N_2527,N_2123,N_1663);
or U2528 (N_2528,N_1664,N_1636);
xnor U2529 (N_2529,N_1697,N_2031);
or U2530 (N_2530,N_1534,N_1500);
and U2531 (N_2531,N_1656,N_2073);
nand U2532 (N_2532,N_1905,N_1755);
and U2533 (N_2533,N_1583,N_1820);
or U2534 (N_2534,N_1601,N_1672);
and U2535 (N_2535,N_1520,N_2067);
nor U2536 (N_2536,N_1569,N_1803);
nor U2537 (N_2537,N_1941,N_1753);
nand U2538 (N_2538,N_2197,N_1629);
nand U2539 (N_2539,N_1682,N_1981);
nand U2540 (N_2540,N_1973,N_1836);
nand U2541 (N_2541,N_2161,N_1822);
nor U2542 (N_2542,N_1768,N_1681);
xor U2543 (N_2543,N_1949,N_1850);
xnor U2544 (N_2544,N_1692,N_1683);
or U2545 (N_2545,N_1871,N_1984);
xnor U2546 (N_2546,N_2118,N_1965);
nand U2547 (N_2547,N_1512,N_1918);
and U2548 (N_2548,N_1529,N_2109);
nand U2549 (N_2549,N_1880,N_1846);
xnor U2550 (N_2550,N_1864,N_1687);
xor U2551 (N_2551,N_1611,N_1511);
nand U2552 (N_2552,N_1791,N_1660);
and U2553 (N_2553,N_1750,N_1937);
nor U2554 (N_2554,N_2107,N_1661);
and U2555 (N_2555,N_1906,N_1630);
or U2556 (N_2556,N_1963,N_1954);
nand U2557 (N_2557,N_1578,N_1910);
and U2558 (N_2558,N_2229,N_1645);
or U2559 (N_2559,N_1815,N_2209);
and U2560 (N_2560,N_1987,N_1651);
xor U2561 (N_2561,N_1675,N_1805);
nor U2562 (N_2562,N_1662,N_2163);
nor U2563 (N_2563,N_2136,N_1533);
xor U2564 (N_2564,N_1643,N_1619);
and U2565 (N_2565,N_1624,N_1585);
and U2566 (N_2566,N_1924,N_1823);
and U2567 (N_2567,N_2232,N_2223);
or U2568 (N_2568,N_1574,N_1744);
nand U2569 (N_2569,N_1843,N_2200);
nor U2570 (N_2570,N_1627,N_1969);
nand U2571 (N_2571,N_1936,N_2222);
and U2572 (N_2572,N_1926,N_1790);
xnor U2573 (N_2573,N_1642,N_2007);
nand U2574 (N_2574,N_1607,N_1738);
xor U2575 (N_2575,N_2178,N_2147);
nand U2576 (N_2576,N_2028,N_2239);
nor U2577 (N_2577,N_1575,N_2169);
xor U2578 (N_2578,N_2112,N_2189);
nor U2579 (N_2579,N_1609,N_1586);
nand U2580 (N_2580,N_2240,N_1680);
and U2581 (N_2581,N_2004,N_1747);
xor U2582 (N_2582,N_1903,N_2156);
or U2583 (N_2583,N_1842,N_1853);
xor U2584 (N_2584,N_1782,N_1731);
or U2585 (N_2585,N_1544,N_2091);
or U2586 (N_2586,N_1525,N_1641);
xnor U2587 (N_2587,N_1988,N_1765);
and U2588 (N_2588,N_1502,N_2193);
and U2589 (N_2589,N_1551,N_1555);
xor U2590 (N_2590,N_2115,N_1771);
nor U2591 (N_2591,N_2038,N_1522);
or U2592 (N_2592,N_1616,N_1938);
nand U2593 (N_2593,N_1933,N_2202);
nor U2594 (N_2594,N_1671,N_2012);
nand U2595 (N_2595,N_2083,N_2220);
nor U2596 (N_2596,N_2208,N_1633);
and U2597 (N_2597,N_1605,N_1804);
nand U2598 (N_2598,N_2098,N_1837);
nand U2599 (N_2599,N_2077,N_1772);
xnor U2600 (N_2600,N_2024,N_1558);
nor U2601 (N_2601,N_1787,N_1668);
and U2602 (N_2602,N_1646,N_1861);
or U2603 (N_2603,N_2053,N_1860);
or U2604 (N_2604,N_1610,N_1908);
and U2605 (N_2605,N_1589,N_1821);
nand U2606 (N_2606,N_1827,N_1783);
nor U2607 (N_2607,N_1945,N_1595);
nor U2608 (N_2608,N_2211,N_1632);
or U2609 (N_2609,N_2153,N_2226);
xnor U2610 (N_2610,N_1652,N_2246);
xor U2611 (N_2611,N_2003,N_1825);
nor U2612 (N_2612,N_1862,N_2070);
or U2613 (N_2613,N_1545,N_1613);
or U2614 (N_2614,N_1686,N_1582);
and U2615 (N_2615,N_2104,N_1801);
nand U2616 (N_2616,N_2245,N_1792);
xor U2617 (N_2617,N_1542,N_1615);
xnor U2618 (N_2618,N_2066,N_1530);
and U2619 (N_2619,N_1728,N_1865);
nor U2620 (N_2620,N_2184,N_1669);
and U2621 (N_2621,N_2152,N_1958);
nor U2622 (N_2622,N_1658,N_1767);
xor U2623 (N_2623,N_1576,N_1930);
nand U2624 (N_2624,N_1874,N_1814);
xor U2625 (N_2625,N_1601,N_1945);
or U2626 (N_2626,N_1780,N_1614);
or U2627 (N_2627,N_2188,N_1698);
nor U2628 (N_2628,N_2123,N_1867);
nand U2629 (N_2629,N_1659,N_2130);
or U2630 (N_2630,N_2208,N_2064);
or U2631 (N_2631,N_1910,N_1662);
nor U2632 (N_2632,N_1512,N_2005);
nand U2633 (N_2633,N_1893,N_1858);
or U2634 (N_2634,N_1577,N_1555);
and U2635 (N_2635,N_1992,N_1983);
nor U2636 (N_2636,N_2117,N_2156);
or U2637 (N_2637,N_1831,N_2029);
and U2638 (N_2638,N_1803,N_2173);
and U2639 (N_2639,N_1812,N_1644);
and U2640 (N_2640,N_1894,N_1829);
nand U2641 (N_2641,N_2200,N_2155);
nor U2642 (N_2642,N_1872,N_1922);
nand U2643 (N_2643,N_1539,N_1996);
xor U2644 (N_2644,N_2064,N_2027);
nor U2645 (N_2645,N_2131,N_2029);
nor U2646 (N_2646,N_1839,N_1974);
and U2647 (N_2647,N_1857,N_2101);
nand U2648 (N_2648,N_1785,N_1899);
nor U2649 (N_2649,N_1546,N_2045);
xor U2650 (N_2650,N_2164,N_1532);
xor U2651 (N_2651,N_2007,N_1944);
or U2652 (N_2652,N_1541,N_1946);
xnor U2653 (N_2653,N_1638,N_1683);
or U2654 (N_2654,N_2243,N_1760);
nand U2655 (N_2655,N_1684,N_1694);
nor U2656 (N_2656,N_2157,N_2211);
nor U2657 (N_2657,N_1973,N_1978);
nor U2658 (N_2658,N_1940,N_1990);
nand U2659 (N_2659,N_1857,N_2117);
or U2660 (N_2660,N_1987,N_1691);
nand U2661 (N_2661,N_1788,N_1716);
xor U2662 (N_2662,N_2018,N_1821);
nor U2663 (N_2663,N_1544,N_1856);
and U2664 (N_2664,N_1648,N_2095);
nand U2665 (N_2665,N_2127,N_1768);
and U2666 (N_2666,N_2224,N_2058);
and U2667 (N_2667,N_2174,N_2229);
nor U2668 (N_2668,N_1799,N_1879);
nor U2669 (N_2669,N_1985,N_1906);
and U2670 (N_2670,N_1511,N_2073);
xnor U2671 (N_2671,N_2041,N_1768);
nor U2672 (N_2672,N_2186,N_2190);
or U2673 (N_2673,N_1847,N_1720);
and U2674 (N_2674,N_1680,N_1586);
xor U2675 (N_2675,N_1635,N_1822);
and U2676 (N_2676,N_1925,N_1601);
nand U2677 (N_2677,N_2138,N_1766);
or U2678 (N_2678,N_2002,N_1668);
nor U2679 (N_2679,N_1794,N_1735);
and U2680 (N_2680,N_2126,N_1972);
and U2681 (N_2681,N_1973,N_1654);
nand U2682 (N_2682,N_2190,N_2125);
nor U2683 (N_2683,N_1922,N_1609);
xor U2684 (N_2684,N_2048,N_1804);
xnor U2685 (N_2685,N_1557,N_1795);
or U2686 (N_2686,N_2164,N_2154);
xor U2687 (N_2687,N_1704,N_1900);
and U2688 (N_2688,N_1660,N_1661);
nand U2689 (N_2689,N_1699,N_1559);
or U2690 (N_2690,N_1524,N_1513);
nor U2691 (N_2691,N_1592,N_2231);
and U2692 (N_2692,N_2136,N_1738);
or U2693 (N_2693,N_1990,N_1534);
and U2694 (N_2694,N_1583,N_2163);
nand U2695 (N_2695,N_1845,N_1651);
and U2696 (N_2696,N_1593,N_1558);
and U2697 (N_2697,N_1829,N_1978);
nand U2698 (N_2698,N_2069,N_2028);
nor U2699 (N_2699,N_1889,N_1824);
nand U2700 (N_2700,N_2191,N_2028);
xor U2701 (N_2701,N_2178,N_2219);
nand U2702 (N_2702,N_1655,N_2061);
or U2703 (N_2703,N_2224,N_1571);
xnor U2704 (N_2704,N_2086,N_1904);
nor U2705 (N_2705,N_1686,N_1991);
or U2706 (N_2706,N_2106,N_1535);
nor U2707 (N_2707,N_1905,N_1582);
or U2708 (N_2708,N_2165,N_2060);
nor U2709 (N_2709,N_1867,N_1555);
nor U2710 (N_2710,N_1609,N_2008);
xnor U2711 (N_2711,N_2169,N_1601);
or U2712 (N_2712,N_1645,N_2192);
nand U2713 (N_2713,N_1942,N_1871);
nand U2714 (N_2714,N_1925,N_2189);
or U2715 (N_2715,N_2072,N_1673);
and U2716 (N_2716,N_2214,N_2173);
or U2717 (N_2717,N_1857,N_2215);
and U2718 (N_2718,N_1892,N_2157);
and U2719 (N_2719,N_2116,N_1920);
nor U2720 (N_2720,N_1757,N_1989);
or U2721 (N_2721,N_1597,N_1743);
or U2722 (N_2722,N_1827,N_1504);
nand U2723 (N_2723,N_1581,N_1626);
and U2724 (N_2724,N_2113,N_1627);
or U2725 (N_2725,N_1687,N_1926);
or U2726 (N_2726,N_2228,N_1691);
nor U2727 (N_2727,N_1981,N_1581);
and U2728 (N_2728,N_1639,N_1884);
xnor U2729 (N_2729,N_2246,N_1508);
nor U2730 (N_2730,N_1788,N_1547);
nand U2731 (N_2731,N_2105,N_1830);
xnor U2732 (N_2732,N_1823,N_2204);
or U2733 (N_2733,N_1831,N_1662);
xnor U2734 (N_2734,N_1764,N_1650);
nand U2735 (N_2735,N_1749,N_2068);
and U2736 (N_2736,N_2132,N_2233);
nor U2737 (N_2737,N_2001,N_1715);
and U2738 (N_2738,N_1787,N_1684);
nand U2739 (N_2739,N_1550,N_1615);
and U2740 (N_2740,N_1635,N_2152);
nand U2741 (N_2741,N_1981,N_1883);
nor U2742 (N_2742,N_2055,N_1987);
and U2743 (N_2743,N_2124,N_1527);
nand U2744 (N_2744,N_2095,N_1926);
or U2745 (N_2745,N_2003,N_2218);
xor U2746 (N_2746,N_2150,N_2066);
or U2747 (N_2747,N_1915,N_1687);
xor U2748 (N_2748,N_2087,N_1830);
xnor U2749 (N_2749,N_1918,N_1982);
nor U2750 (N_2750,N_1798,N_2191);
and U2751 (N_2751,N_1689,N_2006);
and U2752 (N_2752,N_1614,N_1729);
nor U2753 (N_2753,N_1871,N_1713);
xor U2754 (N_2754,N_1591,N_1816);
and U2755 (N_2755,N_1618,N_1725);
nand U2756 (N_2756,N_2125,N_2243);
or U2757 (N_2757,N_2032,N_1556);
nand U2758 (N_2758,N_2106,N_2207);
xor U2759 (N_2759,N_1623,N_1566);
nand U2760 (N_2760,N_2162,N_1705);
or U2761 (N_2761,N_2049,N_1969);
and U2762 (N_2762,N_1598,N_2101);
or U2763 (N_2763,N_1736,N_2036);
and U2764 (N_2764,N_1614,N_1782);
or U2765 (N_2765,N_1580,N_2016);
xor U2766 (N_2766,N_2160,N_1787);
nand U2767 (N_2767,N_1517,N_1769);
nor U2768 (N_2768,N_2172,N_1640);
or U2769 (N_2769,N_1586,N_1569);
nor U2770 (N_2770,N_1833,N_1951);
xor U2771 (N_2771,N_1762,N_1956);
or U2772 (N_2772,N_1695,N_1902);
or U2773 (N_2773,N_2163,N_1538);
xor U2774 (N_2774,N_1983,N_1540);
or U2775 (N_2775,N_1717,N_1901);
and U2776 (N_2776,N_1739,N_1895);
nor U2777 (N_2777,N_2063,N_1956);
xor U2778 (N_2778,N_1739,N_1964);
xnor U2779 (N_2779,N_2007,N_2057);
or U2780 (N_2780,N_1658,N_1747);
xor U2781 (N_2781,N_1789,N_2044);
nor U2782 (N_2782,N_1594,N_1772);
and U2783 (N_2783,N_1838,N_1718);
nand U2784 (N_2784,N_1936,N_1568);
nand U2785 (N_2785,N_1741,N_1783);
xnor U2786 (N_2786,N_1977,N_1564);
nor U2787 (N_2787,N_1508,N_1891);
nand U2788 (N_2788,N_1959,N_1864);
nand U2789 (N_2789,N_1762,N_1562);
nand U2790 (N_2790,N_2122,N_2114);
or U2791 (N_2791,N_2177,N_1736);
or U2792 (N_2792,N_2069,N_1590);
or U2793 (N_2793,N_1698,N_2075);
and U2794 (N_2794,N_1801,N_2187);
and U2795 (N_2795,N_1858,N_1882);
nand U2796 (N_2796,N_1682,N_1660);
nand U2797 (N_2797,N_1719,N_2023);
nand U2798 (N_2798,N_1823,N_1830);
and U2799 (N_2799,N_1902,N_1981);
nand U2800 (N_2800,N_2064,N_2160);
nor U2801 (N_2801,N_1769,N_1765);
nand U2802 (N_2802,N_1598,N_1849);
or U2803 (N_2803,N_1648,N_1844);
and U2804 (N_2804,N_1763,N_1698);
xnor U2805 (N_2805,N_1866,N_2116);
nand U2806 (N_2806,N_1669,N_1894);
or U2807 (N_2807,N_2088,N_1950);
and U2808 (N_2808,N_1633,N_1948);
or U2809 (N_2809,N_1805,N_2158);
or U2810 (N_2810,N_2032,N_1600);
nor U2811 (N_2811,N_1692,N_2082);
or U2812 (N_2812,N_1814,N_1821);
nand U2813 (N_2813,N_2001,N_1794);
nor U2814 (N_2814,N_2166,N_1982);
and U2815 (N_2815,N_1845,N_1932);
nand U2816 (N_2816,N_1504,N_2244);
and U2817 (N_2817,N_1535,N_1945);
or U2818 (N_2818,N_1885,N_1562);
nand U2819 (N_2819,N_1829,N_1544);
and U2820 (N_2820,N_1869,N_2061);
nor U2821 (N_2821,N_1972,N_1648);
xor U2822 (N_2822,N_1966,N_1802);
nand U2823 (N_2823,N_2150,N_2045);
nand U2824 (N_2824,N_1998,N_1760);
or U2825 (N_2825,N_1923,N_1840);
nor U2826 (N_2826,N_2200,N_2142);
and U2827 (N_2827,N_1721,N_2012);
nor U2828 (N_2828,N_1632,N_2000);
nand U2829 (N_2829,N_2232,N_1580);
nor U2830 (N_2830,N_2109,N_2141);
or U2831 (N_2831,N_2079,N_1570);
xor U2832 (N_2832,N_2052,N_2032);
nor U2833 (N_2833,N_2230,N_2229);
or U2834 (N_2834,N_1578,N_1942);
nand U2835 (N_2835,N_1710,N_1917);
xnor U2836 (N_2836,N_1650,N_1586);
nor U2837 (N_2837,N_1647,N_2191);
nand U2838 (N_2838,N_2080,N_2113);
nand U2839 (N_2839,N_1505,N_1548);
or U2840 (N_2840,N_1780,N_1605);
and U2841 (N_2841,N_1705,N_2136);
nand U2842 (N_2842,N_1831,N_1563);
nor U2843 (N_2843,N_2052,N_1679);
or U2844 (N_2844,N_1576,N_1868);
and U2845 (N_2845,N_1632,N_1758);
nand U2846 (N_2846,N_1685,N_2104);
or U2847 (N_2847,N_1612,N_1605);
nor U2848 (N_2848,N_1914,N_2162);
nand U2849 (N_2849,N_1619,N_1906);
nor U2850 (N_2850,N_2012,N_1899);
nor U2851 (N_2851,N_1596,N_1748);
nor U2852 (N_2852,N_1880,N_1825);
and U2853 (N_2853,N_1523,N_1690);
nor U2854 (N_2854,N_1859,N_1962);
and U2855 (N_2855,N_1736,N_1868);
or U2856 (N_2856,N_2132,N_1734);
or U2857 (N_2857,N_1780,N_2116);
xnor U2858 (N_2858,N_1699,N_1674);
xnor U2859 (N_2859,N_1687,N_1592);
or U2860 (N_2860,N_2077,N_2062);
nor U2861 (N_2861,N_2169,N_2136);
xnor U2862 (N_2862,N_1776,N_1857);
xor U2863 (N_2863,N_1587,N_2040);
nand U2864 (N_2864,N_2009,N_1674);
nor U2865 (N_2865,N_1834,N_1805);
and U2866 (N_2866,N_2131,N_1805);
nand U2867 (N_2867,N_1743,N_1529);
nand U2868 (N_2868,N_1653,N_1672);
xor U2869 (N_2869,N_2178,N_1818);
xor U2870 (N_2870,N_2065,N_1711);
nand U2871 (N_2871,N_1501,N_1560);
nor U2872 (N_2872,N_1842,N_1902);
or U2873 (N_2873,N_2040,N_2028);
nand U2874 (N_2874,N_1610,N_2102);
and U2875 (N_2875,N_1745,N_2227);
and U2876 (N_2876,N_2227,N_1699);
xor U2877 (N_2877,N_1501,N_1764);
xnor U2878 (N_2878,N_1943,N_1772);
and U2879 (N_2879,N_1522,N_1689);
and U2880 (N_2880,N_1534,N_1711);
and U2881 (N_2881,N_1962,N_2015);
and U2882 (N_2882,N_1867,N_2195);
nand U2883 (N_2883,N_1755,N_1618);
and U2884 (N_2884,N_1933,N_1685);
xnor U2885 (N_2885,N_1657,N_2066);
and U2886 (N_2886,N_1780,N_2018);
or U2887 (N_2887,N_2249,N_1907);
nor U2888 (N_2888,N_1922,N_1968);
nor U2889 (N_2889,N_2208,N_1767);
or U2890 (N_2890,N_2243,N_2189);
and U2891 (N_2891,N_1794,N_1730);
or U2892 (N_2892,N_1966,N_1583);
or U2893 (N_2893,N_1552,N_2063);
and U2894 (N_2894,N_1626,N_1609);
nand U2895 (N_2895,N_1732,N_1524);
nand U2896 (N_2896,N_1905,N_1511);
and U2897 (N_2897,N_1742,N_1992);
xor U2898 (N_2898,N_1672,N_1880);
nor U2899 (N_2899,N_2044,N_1660);
nor U2900 (N_2900,N_1505,N_2075);
or U2901 (N_2901,N_1686,N_2246);
and U2902 (N_2902,N_1669,N_1844);
nor U2903 (N_2903,N_2178,N_1689);
nor U2904 (N_2904,N_1893,N_2160);
nand U2905 (N_2905,N_1757,N_1528);
nor U2906 (N_2906,N_2183,N_1855);
xnor U2907 (N_2907,N_2114,N_1893);
nor U2908 (N_2908,N_2018,N_2149);
xor U2909 (N_2909,N_2211,N_2117);
and U2910 (N_2910,N_1695,N_1977);
or U2911 (N_2911,N_1575,N_1634);
or U2912 (N_2912,N_1967,N_1684);
nand U2913 (N_2913,N_2168,N_1890);
xnor U2914 (N_2914,N_1992,N_2169);
nor U2915 (N_2915,N_2213,N_1712);
nand U2916 (N_2916,N_1559,N_1878);
nor U2917 (N_2917,N_1838,N_1895);
or U2918 (N_2918,N_1502,N_1656);
xnor U2919 (N_2919,N_1646,N_2211);
and U2920 (N_2920,N_1572,N_1562);
nand U2921 (N_2921,N_2185,N_2136);
and U2922 (N_2922,N_1978,N_1548);
and U2923 (N_2923,N_1515,N_1638);
nor U2924 (N_2924,N_2021,N_1751);
or U2925 (N_2925,N_2006,N_1866);
and U2926 (N_2926,N_1845,N_1650);
or U2927 (N_2927,N_2011,N_1700);
xor U2928 (N_2928,N_1599,N_1768);
xnor U2929 (N_2929,N_1659,N_1762);
nand U2930 (N_2930,N_1648,N_2067);
or U2931 (N_2931,N_2202,N_1851);
and U2932 (N_2932,N_1791,N_2224);
nand U2933 (N_2933,N_1738,N_1662);
nor U2934 (N_2934,N_2131,N_2018);
or U2935 (N_2935,N_2148,N_1619);
nor U2936 (N_2936,N_2092,N_1501);
or U2937 (N_2937,N_1952,N_1591);
or U2938 (N_2938,N_1594,N_1730);
or U2939 (N_2939,N_1515,N_1698);
nand U2940 (N_2940,N_1721,N_1716);
nor U2941 (N_2941,N_2108,N_1514);
nand U2942 (N_2942,N_1825,N_2076);
nand U2943 (N_2943,N_2020,N_1673);
and U2944 (N_2944,N_1845,N_1654);
xor U2945 (N_2945,N_1557,N_2054);
or U2946 (N_2946,N_1887,N_2065);
or U2947 (N_2947,N_1679,N_1869);
nand U2948 (N_2948,N_1955,N_2070);
xor U2949 (N_2949,N_2018,N_1622);
nand U2950 (N_2950,N_1626,N_1549);
nor U2951 (N_2951,N_1929,N_2143);
nor U2952 (N_2952,N_2203,N_1776);
nand U2953 (N_2953,N_1920,N_2140);
or U2954 (N_2954,N_1632,N_2073);
xor U2955 (N_2955,N_2168,N_1859);
nor U2956 (N_2956,N_1687,N_1933);
xnor U2957 (N_2957,N_1657,N_1557);
and U2958 (N_2958,N_1561,N_2223);
nor U2959 (N_2959,N_1959,N_2027);
and U2960 (N_2960,N_1720,N_2068);
xnor U2961 (N_2961,N_1795,N_1946);
and U2962 (N_2962,N_1892,N_1725);
xor U2963 (N_2963,N_1822,N_1664);
xnor U2964 (N_2964,N_2209,N_2152);
nor U2965 (N_2965,N_2242,N_2112);
and U2966 (N_2966,N_2090,N_2137);
and U2967 (N_2967,N_1771,N_1952);
and U2968 (N_2968,N_1638,N_2158);
or U2969 (N_2969,N_2169,N_1569);
nor U2970 (N_2970,N_2057,N_2130);
and U2971 (N_2971,N_2238,N_2012);
and U2972 (N_2972,N_1716,N_1791);
or U2973 (N_2973,N_2208,N_1613);
xor U2974 (N_2974,N_1829,N_1951);
nand U2975 (N_2975,N_1691,N_2027);
xnor U2976 (N_2976,N_2195,N_2097);
nand U2977 (N_2977,N_2031,N_2192);
or U2978 (N_2978,N_1846,N_2031);
nor U2979 (N_2979,N_2215,N_1570);
xor U2980 (N_2980,N_1723,N_1738);
and U2981 (N_2981,N_2127,N_1605);
xnor U2982 (N_2982,N_1808,N_2131);
or U2983 (N_2983,N_1655,N_1525);
nor U2984 (N_2984,N_2170,N_1810);
and U2985 (N_2985,N_1549,N_1935);
xor U2986 (N_2986,N_1626,N_1734);
xnor U2987 (N_2987,N_2132,N_1985);
nor U2988 (N_2988,N_1784,N_1671);
nor U2989 (N_2989,N_1500,N_2118);
xor U2990 (N_2990,N_1834,N_1730);
or U2991 (N_2991,N_1518,N_2064);
xor U2992 (N_2992,N_1790,N_1632);
and U2993 (N_2993,N_2016,N_1950);
nor U2994 (N_2994,N_2128,N_1608);
nor U2995 (N_2995,N_2185,N_1610);
xnor U2996 (N_2996,N_2103,N_1731);
nand U2997 (N_2997,N_1833,N_1893);
and U2998 (N_2998,N_1914,N_2115);
or U2999 (N_2999,N_1762,N_2184);
nor U3000 (N_3000,N_2918,N_2792);
and U3001 (N_3001,N_2430,N_2274);
nor U3002 (N_3002,N_2574,N_2538);
and U3003 (N_3003,N_2373,N_2816);
and U3004 (N_3004,N_2714,N_2415);
nand U3005 (N_3005,N_2524,N_2600);
or U3006 (N_3006,N_2523,N_2854);
or U3007 (N_3007,N_2475,N_2972);
nand U3008 (N_3008,N_2550,N_2681);
and U3009 (N_3009,N_2751,N_2670);
and U3010 (N_3010,N_2990,N_2323);
and U3011 (N_3011,N_2951,N_2336);
nand U3012 (N_3012,N_2709,N_2535);
and U3013 (N_3013,N_2431,N_2326);
and U3014 (N_3014,N_2954,N_2702);
and U3015 (N_3015,N_2590,N_2517);
nand U3016 (N_3016,N_2963,N_2891);
nand U3017 (N_3017,N_2484,N_2878);
or U3018 (N_3018,N_2465,N_2541);
or U3019 (N_3019,N_2664,N_2700);
xor U3020 (N_3020,N_2426,N_2438);
or U3021 (N_3021,N_2901,N_2254);
or U3022 (N_3022,N_2307,N_2689);
nor U3023 (N_3023,N_2761,N_2947);
and U3024 (N_3024,N_2937,N_2850);
xnor U3025 (N_3025,N_2722,N_2748);
or U3026 (N_3026,N_2643,N_2626);
nor U3027 (N_3027,N_2644,N_2340);
and U3028 (N_3028,N_2788,N_2707);
nor U3029 (N_3029,N_2335,N_2776);
nand U3030 (N_3030,N_2394,N_2741);
and U3031 (N_3031,N_2488,N_2468);
xor U3032 (N_3032,N_2455,N_2253);
nor U3033 (N_3033,N_2530,N_2531);
nand U3034 (N_3034,N_2623,N_2851);
nor U3035 (N_3035,N_2942,N_2258);
nand U3036 (N_3036,N_2889,N_2865);
nand U3037 (N_3037,N_2601,N_2656);
nand U3038 (N_3038,N_2858,N_2435);
nor U3039 (N_3039,N_2364,N_2270);
and U3040 (N_3040,N_2938,N_2405);
xnor U3041 (N_3041,N_2647,N_2553);
and U3042 (N_3042,N_2318,N_2305);
nand U3043 (N_3043,N_2312,N_2817);
xor U3044 (N_3044,N_2402,N_2559);
or U3045 (N_3045,N_2347,N_2434);
xor U3046 (N_3046,N_2683,N_2775);
and U3047 (N_3047,N_2471,N_2502);
nand U3048 (N_3048,N_2487,N_2380);
nor U3049 (N_3049,N_2387,N_2799);
xnor U3050 (N_3050,N_2446,N_2639);
nor U3051 (N_3051,N_2718,N_2806);
nor U3052 (N_3052,N_2259,N_2450);
nand U3053 (N_3053,N_2859,N_2328);
nand U3054 (N_3054,N_2795,N_2971);
xnor U3055 (N_3055,N_2786,N_2818);
or U3056 (N_3056,N_2866,N_2470);
nor U3057 (N_3057,N_2390,N_2310);
or U3058 (N_3058,N_2992,N_2606);
xnor U3059 (N_3059,N_2584,N_2991);
or U3060 (N_3060,N_2422,N_2619);
and U3061 (N_3061,N_2356,N_2561);
xor U3062 (N_3062,N_2263,N_2410);
xnor U3063 (N_3063,N_2466,N_2374);
and U3064 (N_3064,N_2663,N_2874);
or U3065 (N_3065,N_2887,N_2883);
nand U3066 (N_3066,N_2908,N_2445);
xor U3067 (N_3067,N_2986,N_2367);
nand U3068 (N_3068,N_2311,N_2962);
or U3069 (N_3069,N_2782,N_2618);
nor U3070 (N_3070,N_2463,N_2745);
xor U3071 (N_3071,N_2712,N_2399);
nand U3072 (N_3072,N_2697,N_2351);
nor U3073 (N_3073,N_2354,N_2691);
and U3074 (N_3074,N_2558,N_2357);
or U3075 (N_3075,N_2526,N_2638);
xnor U3076 (N_3076,N_2542,N_2375);
nand U3077 (N_3077,N_2406,N_2515);
nand U3078 (N_3078,N_2621,N_2327);
xnor U3079 (N_3079,N_2716,N_2605);
xor U3080 (N_3080,N_2358,N_2384);
nor U3081 (N_3081,N_2899,N_2540);
or U3082 (N_3082,N_2687,N_2770);
nand U3083 (N_3083,N_2674,N_2407);
xor U3084 (N_3084,N_2966,N_2864);
or U3085 (N_3085,N_2424,N_2950);
nor U3086 (N_3086,N_2876,N_2863);
and U3087 (N_3087,N_2759,N_2699);
nor U3088 (N_3088,N_2442,N_2796);
nor U3089 (N_3089,N_2955,N_2439);
nor U3090 (N_3090,N_2295,N_2765);
nor U3091 (N_3091,N_2843,N_2580);
xnor U3092 (N_3092,N_2694,N_2490);
nor U3093 (N_3093,N_2255,N_2652);
xnor U3094 (N_3094,N_2520,N_2428);
and U3095 (N_3095,N_2945,N_2627);
xnor U3096 (N_3096,N_2568,N_2291);
xnor U3097 (N_3097,N_2729,N_2754);
xor U3098 (N_3098,N_2585,N_2570);
nor U3099 (N_3099,N_2653,N_2688);
or U3100 (N_3100,N_2649,N_2974);
nor U3101 (N_3101,N_2365,N_2802);
nand U3102 (N_3102,N_2979,N_2416);
xnor U3103 (N_3103,N_2845,N_2432);
nand U3104 (N_3104,N_2642,N_2299);
nand U3105 (N_3105,N_2982,N_2824);
nand U3106 (N_3106,N_2698,N_2360);
xnor U3107 (N_3107,N_2717,N_2659);
xnor U3108 (N_3108,N_2926,N_2277);
nor U3109 (N_3109,N_2682,N_2680);
or U3110 (N_3110,N_2830,N_2667);
nand U3111 (N_3111,N_2267,N_2904);
nand U3112 (N_3112,N_2331,N_2884);
xnor U3113 (N_3113,N_2777,N_2496);
nor U3114 (N_3114,N_2345,N_2313);
or U3115 (N_3115,N_2798,N_2975);
and U3116 (N_3116,N_2289,N_2730);
and U3117 (N_3117,N_2497,N_2467);
and U3118 (N_3118,N_2793,N_2921);
or U3119 (N_3119,N_2368,N_2723);
nor U3120 (N_3120,N_2564,N_2720);
or U3121 (N_3121,N_2361,N_2257);
or U3122 (N_3122,N_2632,N_2493);
nand U3123 (N_3123,N_2482,N_2575);
and U3124 (N_3124,N_2448,N_2890);
and U3125 (N_3125,N_2393,N_2780);
or U3126 (N_3126,N_2505,N_2593);
xnor U3127 (N_3127,N_2984,N_2569);
xor U3128 (N_3128,N_2855,N_2602);
and U3129 (N_3129,N_2755,N_2592);
nand U3130 (N_3130,N_2703,N_2747);
xnor U3131 (N_3131,N_2304,N_2612);
nand U3132 (N_3132,N_2923,N_2783);
xor U3133 (N_3133,N_2516,N_2711);
nor U3134 (N_3134,N_2427,N_2298);
and U3135 (N_3135,N_2543,N_2847);
and U3136 (N_3136,N_2977,N_2348);
or U3137 (N_3137,N_2460,N_2774);
xnor U3138 (N_3138,N_2337,N_2338);
nor U3139 (N_3139,N_2481,N_2300);
xnor U3140 (N_3140,N_2737,N_2370);
xnor U3141 (N_3141,N_2614,N_2451);
nand U3142 (N_3142,N_2693,N_2763);
xor U3143 (N_3143,N_2309,N_2322);
nor U3144 (N_3144,N_2772,N_2732);
and U3145 (N_3145,N_2603,N_2419);
and U3146 (N_3146,N_2953,N_2476);
nor U3147 (N_3147,N_2743,N_2790);
and U3148 (N_3148,N_2549,N_2853);
nand U3149 (N_3149,N_2967,N_2939);
xnor U3150 (N_3150,N_2286,N_2452);
or U3151 (N_3151,N_2268,N_2636);
nand U3152 (N_3152,N_2925,N_2646);
and U3153 (N_3153,N_2981,N_2701);
and U3154 (N_3154,N_2705,N_2260);
xnor U3155 (N_3155,N_2607,N_2400);
nor U3156 (N_3156,N_2555,N_2290);
xor U3157 (N_3157,N_2521,N_2522);
xor U3158 (N_3158,N_2385,N_2457);
or U3159 (N_3159,N_2856,N_2495);
nor U3160 (N_3160,N_2650,N_2911);
and U3161 (N_3161,N_2486,N_2789);
nand U3162 (N_3162,N_2746,N_2803);
or U3163 (N_3163,N_2848,N_2534);
xnor U3164 (N_3164,N_2846,N_2713);
or U3165 (N_3165,N_2425,N_2871);
nor U3166 (N_3166,N_2492,N_2279);
nand U3167 (N_3167,N_2936,N_2423);
nor U3168 (N_3168,N_2464,N_2999);
and U3169 (N_3169,N_2869,N_2302);
and U3170 (N_3170,N_2897,N_2836);
xor U3171 (N_3171,N_2778,N_2868);
nand U3172 (N_3172,N_2912,N_2379);
xor U3173 (N_3173,N_2376,N_2959);
and U3174 (N_3174,N_2581,N_2742);
xnor U3175 (N_3175,N_2640,N_2414);
nand U3176 (N_3176,N_2898,N_2572);
nand U3177 (N_3177,N_2329,N_2319);
and U3178 (N_3178,N_2334,N_2609);
nand U3179 (N_3179,N_2766,N_2834);
and U3180 (N_3180,N_2444,N_2436);
nor U3181 (N_3181,N_2504,N_2749);
nand U3182 (N_3182,N_2395,N_2801);
nand U3183 (N_3183,N_2833,N_2661);
or U3184 (N_3184,N_2562,N_2842);
nor U3185 (N_3185,N_2731,N_2511);
nand U3186 (N_3186,N_2800,N_2815);
nand U3187 (N_3187,N_2736,N_2769);
nor U3188 (N_3188,N_2403,N_2757);
xor U3189 (N_3189,N_2401,N_2507);
xor U3190 (N_3190,N_2919,N_2610);
and U3191 (N_3191,N_2281,N_2762);
and U3192 (N_3192,N_2679,N_2383);
xnor U3193 (N_3193,N_2886,N_2797);
nand U3194 (N_3194,N_2785,N_2684);
nor U3195 (N_3195,N_2764,N_2784);
xnor U3196 (N_3196,N_2760,N_2449);
nand U3197 (N_3197,N_2733,N_2849);
xor U3198 (N_3198,N_2655,N_2840);
nor U3199 (N_3199,N_2728,N_2261);
nand U3200 (N_3200,N_2758,N_2862);
and U3201 (N_3201,N_2724,N_2350);
xor U3202 (N_3202,N_2624,N_2514);
nor U3203 (N_3203,N_2989,N_2819);
or U3204 (N_3204,N_2491,N_2506);
and U3205 (N_3205,N_2404,N_2461);
xor U3206 (N_3206,N_2630,N_2995);
nor U3207 (N_3207,N_2651,N_2927);
nor U3208 (N_3208,N_2994,N_2931);
or U3209 (N_3209,N_2325,N_2536);
nand U3210 (N_3210,N_2417,N_2576);
or U3211 (N_3211,N_2831,N_2894);
nand U3212 (N_3212,N_2509,N_2631);
nor U3213 (N_3213,N_2301,N_2969);
or U3214 (N_3214,N_2895,N_2316);
or U3215 (N_3215,N_2922,N_2993);
nor U3216 (N_3216,N_2529,N_2372);
xor U3217 (N_3217,N_2821,N_2551);
nor U3218 (N_3218,N_2537,N_2499);
and U3219 (N_3219,N_2589,N_2998);
xor U3220 (N_3220,N_2381,N_2478);
xor U3221 (N_3221,N_2933,N_2944);
nor U3222 (N_3222,N_2948,N_2317);
or U3223 (N_3223,N_2658,N_2418);
nor U3224 (N_3224,N_2976,N_2917);
nor U3225 (N_3225,N_2935,N_2265);
or U3226 (N_3226,N_2494,N_2706);
and U3227 (N_3227,N_2861,N_2508);
or U3228 (N_3228,N_2678,N_2293);
xnor U3229 (N_3229,N_2586,N_2719);
or U3230 (N_3230,N_2420,N_2896);
nor U3231 (N_3231,N_2413,N_2598);
or U3232 (N_3232,N_2665,N_2805);
xor U3233 (N_3233,N_2756,N_2512);
nand U3234 (N_3234,N_2675,N_2928);
or U3235 (N_3235,N_2366,N_2264);
xnor U3236 (N_3236,N_2885,N_2548);
or U3237 (N_3237,N_2750,N_2888);
or U3238 (N_3238,N_2662,N_2710);
and U3239 (N_3239,N_2285,N_2635);
xnor U3240 (N_3240,N_2625,N_2909);
nand U3241 (N_3241,N_2276,N_2980);
nand U3242 (N_3242,N_2565,N_2518);
nand U3243 (N_3243,N_2773,N_2941);
and U3244 (N_3244,N_2804,N_2458);
nand U3245 (N_3245,N_2296,N_2477);
nor U3246 (N_3246,N_2839,N_2837);
xor U3247 (N_3247,N_2734,N_2657);
and U3248 (N_3248,N_2794,N_2314);
nor U3249 (N_3249,N_2835,N_2900);
or U3250 (N_3250,N_2411,N_2272);
nand U3251 (N_3251,N_2280,N_2672);
nand U3252 (N_3252,N_2352,N_2582);
and U3253 (N_3253,N_2857,N_2519);
or U3254 (N_3254,N_2595,N_2771);
or U3255 (N_3255,N_2852,N_2692);
nand U3256 (N_3256,N_2303,N_2573);
or U3257 (N_3257,N_2251,N_2828);
and U3258 (N_3258,N_2708,N_2282);
and U3259 (N_3259,N_2563,N_2344);
xor U3260 (N_3260,N_2462,N_2382);
xor U3261 (N_3261,N_2739,N_2753);
xor U3262 (N_3262,N_2250,N_2278);
nand U3263 (N_3263,N_2292,N_2978);
and U3264 (N_3264,N_2829,N_2297);
nor U3265 (N_3265,N_2578,N_2472);
xor U3266 (N_3266,N_2532,N_2500);
xnor U3267 (N_3267,N_2641,N_2949);
nor U3268 (N_3268,N_2877,N_2875);
xor U3269 (N_3269,N_2525,N_2744);
xnor U3270 (N_3270,N_2544,N_2870);
nand U3271 (N_3271,N_2902,N_2892);
or U3272 (N_3272,N_2832,N_2355);
and U3273 (N_3273,N_2617,N_2447);
nand U3274 (N_3274,N_2867,N_2628);
xnor U3275 (N_3275,N_2970,N_2807);
and U3276 (N_3276,N_2704,N_2579);
xnor U3277 (N_3277,N_2860,N_2934);
or U3278 (N_3278,N_2905,N_2668);
or U3279 (N_3279,N_2913,N_2533);
nor U3280 (N_3280,N_2915,N_2841);
and U3281 (N_3281,N_2485,N_2676);
nor U3282 (N_3282,N_2583,N_2914);
and U3283 (N_3283,N_2988,N_2459);
and U3284 (N_3284,N_2392,N_2654);
xnor U3285 (N_3285,N_2513,N_2546);
nor U3286 (N_3286,N_2596,N_2363);
and U3287 (N_3287,N_2985,N_2554);
nand U3288 (N_3288,N_2273,N_2397);
or U3289 (N_3289,N_2408,N_2726);
and U3290 (N_3290,N_2725,N_2369);
nand U3291 (N_3291,N_2910,N_2552);
or U3292 (N_3292,N_2341,N_2827);
xor U3293 (N_3293,N_2440,N_2930);
nor U3294 (N_3294,N_2321,N_2346);
xnor U3295 (N_3295,N_2671,N_2547);
nor U3296 (N_3296,N_2881,N_2262);
and U3297 (N_3297,N_2443,N_2820);
nor U3298 (N_3298,N_2362,N_2940);
and U3299 (N_3299,N_2964,N_2811);
nand U3300 (N_3300,N_2660,N_2973);
or U3301 (N_3301,N_2727,N_2594);
nand U3302 (N_3302,N_2353,N_2308);
nor U3303 (N_3303,N_2412,N_2906);
nor U3304 (N_3304,N_2965,N_2620);
or U3305 (N_3305,N_2695,N_2768);
or U3306 (N_3306,N_2409,N_2677);
and U3307 (N_3307,N_2377,N_2907);
and U3308 (N_3308,N_2571,N_2645);
or U3309 (N_3309,N_2634,N_2738);
nor U3310 (N_3310,N_2320,N_2287);
xor U3311 (N_3311,N_2556,N_2893);
nor U3312 (N_3312,N_2479,N_2903);
or U3313 (N_3313,N_2378,N_2275);
or U3314 (N_3314,N_2838,N_2597);
and U3315 (N_3315,N_2557,N_2315);
nor U3316 (N_3316,N_2616,N_2528);
nor U3317 (N_3317,N_2956,N_2473);
nand U3318 (N_3318,N_2604,N_2599);
xnor U3319 (N_3319,N_2501,N_2987);
nand U3320 (N_3320,N_2721,N_2813);
or U3321 (N_3321,N_2740,N_2997);
nand U3322 (N_3322,N_2545,N_2330);
or U3323 (N_3323,N_2685,N_2715);
nor U3324 (N_3324,N_2983,N_2343);
nand U3325 (N_3325,N_2608,N_2648);
nand U3326 (N_3326,N_2283,N_2916);
nand U3327 (N_3327,N_2791,N_2880);
and U3328 (N_3328,N_2629,N_2591);
nand U3329 (N_3329,N_2735,N_2615);
nand U3330 (N_3330,N_2342,N_2808);
or U3331 (N_3331,N_2873,N_2433);
or U3332 (N_3332,N_2256,N_2996);
nor U3333 (N_3333,N_2396,N_2391);
or U3334 (N_3334,N_2527,N_2577);
nor U3335 (N_3335,N_2456,N_2666);
and U3336 (N_3336,N_2333,N_2294);
nor U3337 (N_3337,N_2371,N_2474);
or U3338 (N_3338,N_2844,N_2673);
xor U3339 (N_3339,N_2929,N_2686);
nand U3340 (N_3340,N_2284,N_2489);
or U3341 (N_3341,N_2588,N_2437);
xnor U3342 (N_3342,N_2946,N_2386);
nand U3343 (N_3343,N_2812,N_2339);
nor U3344 (N_3344,N_2510,N_2441);
and U3345 (N_3345,N_2567,N_2388);
xnor U3346 (N_3346,N_2924,N_2480);
and U3347 (N_3347,N_2810,N_2822);
nand U3348 (N_3348,N_2566,N_2252);
xor U3349 (N_3349,N_2779,N_2696);
xnor U3350 (N_3350,N_2349,N_2823);
and U3351 (N_3351,N_2271,N_2587);
nand U3352 (N_3352,N_2469,N_2952);
or U3353 (N_3353,N_2872,N_2814);
nor U3354 (N_3354,N_2690,N_2622);
xor U3355 (N_3355,N_2539,N_2882);
nand U3356 (N_3356,N_2389,N_2429);
nand U3357 (N_3357,N_2611,N_2398);
and U3358 (N_3358,N_2961,N_2920);
nor U3359 (N_3359,N_2809,N_2787);
and U3360 (N_3360,N_2943,N_2879);
nand U3361 (N_3361,N_2266,N_2288);
nor U3362 (N_3362,N_2958,N_2421);
nor U3363 (N_3363,N_2454,N_2324);
and U3364 (N_3364,N_2957,N_2483);
nand U3365 (N_3365,N_2826,N_2637);
xor U3366 (N_3366,N_2633,N_2669);
nand U3367 (N_3367,N_2503,N_2498);
nor U3368 (N_3368,N_2613,N_2752);
nor U3369 (N_3369,N_2560,N_2960);
and U3370 (N_3370,N_2781,N_2767);
xor U3371 (N_3371,N_2306,N_2269);
xor U3372 (N_3372,N_2332,N_2359);
and U3373 (N_3373,N_2932,N_2453);
xnor U3374 (N_3374,N_2825,N_2968);
nor U3375 (N_3375,N_2376,N_2497);
and U3376 (N_3376,N_2252,N_2945);
nand U3377 (N_3377,N_2592,N_2442);
and U3378 (N_3378,N_2469,N_2346);
nor U3379 (N_3379,N_2462,N_2594);
nand U3380 (N_3380,N_2819,N_2611);
nand U3381 (N_3381,N_2878,N_2987);
nand U3382 (N_3382,N_2981,N_2840);
and U3383 (N_3383,N_2298,N_2423);
or U3384 (N_3384,N_2850,N_2430);
or U3385 (N_3385,N_2450,N_2431);
nor U3386 (N_3386,N_2972,N_2818);
or U3387 (N_3387,N_2962,N_2439);
nand U3388 (N_3388,N_2922,N_2612);
xor U3389 (N_3389,N_2454,N_2567);
xor U3390 (N_3390,N_2342,N_2725);
and U3391 (N_3391,N_2607,N_2448);
nand U3392 (N_3392,N_2820,N_2675);
xnor U3393 (N_3393,N_2921,N_2726);
and U3394 (N_3394,N_2955,N_2713);
nand U3395 (N_3395,N_2770,N_2445);
nand U3396 (N_3396,N_2803,N_2756);
or U3397 (N_3397,N_2768,N_2712);
or U3398 (N_3398,N_2640,N_2716);
nand U3399 (N_3399,N_2590,N_2793);
or U3400 (N_3400,N_2631,N_2993);
xnor U3401 (N_3401,N_2344,N_2653);
nor U3402 (N_3402,N_2526,N_2411);
and U3403 (N_3403,N_2536,N_2652);
or U3404 (N_3404,N_2430,N_2648);
nand U3405 (N_3405,N_2904,N_2434);
and U3406 (N_3406,N_2930,N_2758);
and U3407 (N_3407,N_2830,N_2998);
and U3408 (N_3408,N_2462,N_2415);
xnor U3409 (N_3409,N_2970,N_2347);
xnor U3410 (N_3410,N_2341,N_2735);
xor U3411 (N_3411,N_2964,N_2637);
nand U3412 (N_3412,N_2830,N_2890);
and U3413 (N_3413,N_2348,N_2732);
nor U3414 (N_3414,N_2604,N_2590);
nor U3415 (N_3415,N_2998,N_2610);
and U3416 (N_3416,N_2942,N_2939);
nor U3417 (N_3417,N_2724,N_2710);
nand U3418 (N_3418,N_2899,N_2497);
or U3419 (N_3419,N_2563,N_2987);
nand U3420 (N_3420,N_2484,N_2756);
or U3421 (N_3421,N_2416,N_2970);
or U3422 (N_3422,N_2484,N_2313);
and U3423 (N_3423,N_2613,N_2480);
and U3424 (N_3424,N_2584,N_2722);
nand U3425 (N_3425,N_2551,N_2855);
or U3426 (N_3426,N_2931,N_2424);
xor U3427 (N_3427,N_2288,N_2818);
xor U3428 (N_3428,N_2637,N_2423);
or U3429 (N_3429,N_2840,N_2384);
or U3430 (N_3430,N_2532,N_2632);
nand U3431 (N_3431,N_2899,N_2538);
xnor U3432 (N_3432,N_2702,N_2354);
and U3433 (N_3433,N_2766,N_2979);
nand U3434 (N_3434,N_2836,N_2462);
and U3435 (N_3435,N_2709,N_2657);
or U3436 (N_3436,N_2414,N_2673);
nand U3437 (N_3437,N_2521,N_2318);
or U3438 (N_3438,N_2774,N_2859);
and U3439 (N_3439,N_2439,N_2566);
or U3440 (N_3440,N_2456,N_2278);
nor U3441 (N_3441,N_2272,N_2300);
or U3442 (N_3442,N_2250,N_2592);
xor U3443 (N_3443,N_2408,N_2306);
nand U3444 (N_3444,N_2279,N_2925);
xor U3445 (N_3445,N_2295,N_2470);
nand U3446 (N_3446,N_2737,N_2592);
or U3447 (N_3447,N_2968,N_2831);
nor U3448 (N_3448,N_2906,N_2717);
or U3449 (N_3449,N_2480,N_2683);
or U3450 (N_3450,N_2623,N_2654);
and U3451 (N_3451,N_2814,N_2543);
or U3452 (N_3452,N_2941,N_2474);
or U3453 (N_3453,N_2985,N_2717);
or U3454 (N_3454,N_2859,N_2909);
xor U3455 (N_3455,N_2611,N_2253);
xor U3456 (N_3456,N_2824,N_2860);
xnor U3457 (N_3457,N_2499,N_2285);
nand U3458 (N_3458,N_2591,N_2523);
and U3459 (N_3459,N_2961,N_2323);
nand U3460 (N_3460,N_2357,N_2712);
xnor U3461 (N_3461,N_2624,N_2763);
or U3462 (N_3462,N_2440,N_2443);
or U3463 (N_3463,N_2645,N_2406);
xnor U3464 (N_3464,N_2544,N_2269);
nand U3465 (N_3465,N_2869,N_2456);
xor U3466 (N_3466,N_2582,N_2599);
or U3467 (N_3467,N_2894,N_2298);
nand U3468 (N_3468,N_2436,N_2282);
and U3469 (N_3469,N_2793,N_2786);
nand U3470 (N_3470,N_2489,N_2430);
nor U3471 (N_3471,N_2371,N_2444);
and U3472 (N_3472,N_2777,N_2953);
and U3473 (N_3473,N_2258,N_2541);
and U3474 (N_3474,N_2833,N_2296);
nor U3475 (N_3475,N_2862,N_2737);
nand U3476 (N_3476,N_2916,N_2883);
nor U3477 (N_3477,N_2840,N_2255);
xor U3478 (N_3478,N_2620,N_2727);
or U3479 (N_3479,N_2278,N_2401);
or U3480 (N_3480,N_2326,N_2647);
nand U3481 (N_3481,N_2310,N_2618);
nand U3482 (N_3482,N_2473,N_2903);
or U3483 (N_3483,N_2441,N_2957);
or U3484 (N_3484,N_2604,N_2757);
and U3485 (N_3485,N_2962,N_2869);
and U3486 (N_3486,N_2628,N_2713);
and U3487 (N_3487,N_2469,N_2265);
nand U3488 (N_3488,N_2473,N_2260);
nor U3489 (N_3489,N_2329,N_2432);
nand U3490 (N_3490,N_2500,N_2650);
or U3491 (N_3491,N_2749,N_2386);
nor U3492 (N_3492,N_2767,N_2932);
xnor U3493 (N_3493,N_2296,N_2816);
or U3494 (N_3494,N_2259,N_2391);
nand U3495 (N_3495,N_2753,N_2530);
nand U3496 (N_3496,N_2467,N_2676);
and U3497 (N_3497,N_2696,N_2890);
and U3498 (N_3498,N_2362,N_2696);
nor U3499 (N_3499,N_2760,N_2979);
and U3500 (N_3500,N_2419,N_2855);
nand U3501 (N_3501,N_2777,N_2790);
nor U3502 (N_3502,N_2963,N_2515);
and U3503 (N_3503,N_2940,N_2751);
or U3504 (N_3504,N_2341,N_2730);
or U3505 (N_3505,N_2373,N_2253);
or U3506 (N_3506,N_2900,N_2309);
xor U3507 (N_3507,N_2971,N_2914);
or U3508 (N_3508,N_2565,N_2682);
xor U3509 (N_3509,N_2801,N_2948);
or U3510 (N_3510,N_2784,N_2931);
xor U3511 (N_3511,N_2979,N_2643);
nand U3512 (N_3512,N_2663,N_2526);
or U3513 (N_3513,N_2897,N_2465);
nand U3514 (N_3514,N_2741,N_2491);
and U3515 (N_3515,N_2537,N_2542);
nor U3516 (N_3516,N_2284,N_2298);
nor U3517 (N_3517,N_2307,N_2799);
or U3518 (N_3518,N_2250,N_2520);
nand U3519 (N_3519,N_2476,N_2963);
or U3520 (N_3520,N_2488,N_2943);
xor U3521 (N_3521,N_2669,N_2303);
nor U3522 (N_3522,N_2484,N_2476);
or U3523 (N_3523,N_2401,N_2893);
and U3524 (N_3524,N_2304,N_2895);
or U3525 (N_3525,N_2919,N_2446);
nand U3526 (N_3526,N_2962,N_2750);
and U3527 (N_3527,N_2367,N_2638);
nor U3528 (N_3528,N_2936,N_2584);
and U3529 (N_3529,N_2359,N_2762);
xor U3530 (N_3530,N_2762,N_2529);
or U3531 (N_3531,N_2628,N_2539);
xnor U3532 (N_3532,N_2754,N_2668);
xor U3533 (N_3533,N_2834,N_2274);
nand U3534 (N_3534,N_2351,N_2649);
or U3535 (N_3535,N_2814,N_2450);
xor U3536 (N_3536,N_2704,N_2976);
or U3537 (N_3537,N_2288,N_2640);
nor U3538 (N_3538,N_2353,N_2386);
nand U3539 (N_3539,N_2509,N_2457);
xnor U3540 (N_3540,N_2711,N_2917);
nor U3541 (N_3541,N_2408,N_2293);
xor U3542 (N_3542,N_2856,N_2962);
nor U3543 (N_3543,N_2726,N_2998);
xor U3544 (N_3544,N_2437,N_2822);
xnor U3545 (N_3545,N_2550,N_2644);
or U3546 (N_3546,N_2449,N_2932);
or U3547 (N_3547,N_2252,N_2775);
xor U3548 (N_3548,N_2596,N_2262);
nor U3549 (N_3549,N_2922,N_2568);
xor U3550 (N_3550,N_2979,N_2802);
xnor U3551 (N_3551,N_2977,N_2665);
nand U3552 (N_3552,N_2922,N_2456);
nand U3553 (N_3553,N_2941,N_2739);
nor U3554 (N_3554,N_2456,N_2775);
and U3555 (N_3555,N_2686,N_2462);
nand U3556 (N_3556,N_2761,N_2569);
nand U3557 (N_3557,N_2490,N_2515);
and U3558 (N_3558,N_2429,N_2278);
nand U3559 (N_3559,N_2880,N_2431);
xnor U3560 (N_3560,N_2696,N_2501);
or U3561 (N_3561,N_2796,N_2292);
or U3562 (N_3562,N_2818,N_2982);
nor U3563 (N_3563,N_2748,N_2578);
nand U3564 (N_3564,N_2344,N_2683);
nand U3565 (N_3565,N_2885,N_2765);
xor U3566 (N_3566,N_2844,N_2823);
nor U3567 (N_3567,N_2347,N_2949);
nand U3568 (N_3568,N_2459,N_2915);
xor U3569 (N_3569,N_2749,N_2994);
xnor U3570 (N_3570,N_2823,N_2554);
or U3571 (N_3571,N_2458,N_2540);
or U3572 (N_3572,N_2341,N_2402);
xnor U3573 (N_3573,N_2509,N_2627);
or U3574 (N_3574,N_2433,N_2973);
nor U3575 (N_3575,N_2507,N_2952);
nand U3576 (N_3576,N_2801,N_2976);
nor U3577 (N_3577,N_2720,N_2746);
and U3578 (N_3578,N_2412,N_2651);
nor U3579 (N_3579,N_2755,N_2937);
nor U3580 (N_3580,N_2387,N_2560);
and U3581 (N_3581,N_2948,N_2397);
or U3582 (N_3582,N_2604,N_2338);
nor U3583 (N_3583,N_2623,N_2618);
nor U3584 (N_3584,N_2799,N_2672);
nand U3585 (N_3585,N_2427,N_2571);
nor U3586 (N_3586,N_2647,N_2481);
nand U3587 (N_3587,N_2931,N_2772);
nor U3588 (N_3588,N_2574,N_2397);
or U3589 (N_3589,N_2493,N_2336);
nor U3590 (N_3590,N_2689,N_2514);
and U3591 (N_3591,N_2472,N_2628);
or U3592 (N_3592,N_2544,N_2712);
nor U3593 (N_3593,N_2911,N_2759);
or U3594 (N_3594,N_2439,N_2721);
and U3595 (N_3595,N_2554,N_2801);
xnor U3596 (N_3596,N_2800,N_2758);
nand U3597 (N_3597,N_2747,N_2301);
and U3598 (N_3598,N_2537,N_2475);
or U3599 (N_3599,N_2325,N_2915);
and U3600 (N_3600,N_2689,N_2279);
nand U3601 (N_3601,N_2383,N_2797);
nand U3602 (N_3602,N_2347,N_2412);
and U3603 (N_3603,N_2691,N_2477);
nand U3604 (N_3604,N_2502,N_2453);
and U3605 (N_3605,N_2849,N_2546);
or U3606 (N_3606,N_2387,N_2266);
nand U3607 (N_3607,N_2511,N_2610);
and U3608 (N_3608,N_2753,N_2427);
and U3609 (N_3609,N_2597,N_2431);
and U3610 (N_3610,N_2896,N_2828);
nor U3611 (N_3611,N_2311,N_2868);
xor U3612 (N_3612,N_2396,N_2486);
or U3613 (N_3613,N_2736,N_2778);
or U3614 (N_3614,N_2571,N_2893);
nand U3615 (N_3615,N_2692,N_2331);
xnor U3616 (N_3616,N_2456,N_2931);
xnor U3617 (N_3617,N_2856,N_2929);
or U3618 (N_3618,N_2475,N_2743);
xor U3619 (N_3619,N_2967,N_2605);
xor U3620 (N_3620,N_2802,N_2400);
nor U3621 (N_3621,N_2326,N_2651);
nand U3622 (N_3622,N_2667,N_2996);
nand U3623 (N_3623,N_2459,N_2683);
and U3624 (N_3624,N_2768,N_2507);
xnor U3625 (N_3625,N_2878,N_2554);
and U3626 (N_3626,N_2796,N_2830);
nand U3627 (N_3627,N_2530,N_2592);
nor U3628 (N_3628,N_2606,N_2591);
and U3629 (N_3629,N_2480,N_2388);
or U3630 (N_3630,N_2423,N_2520);
or U3631 (N_3631,N_2317,N_2611);
or U3632 (N_3632,N_2844,N_2607);
nand U3633 (N_3633,N_2687,N_2720);
and U3634 (N_3634,N_2892,N_2537);
nor U3635 (N_3635,N_2591,N_2830);
xor U3636 (N_3636,N_2997,N_2725);
xnor U3637 (N_3637,N_2559,N_2382);
xor U3638 (N_3638,N_2625,N_2402);
nor U3639 (N_3639,N_2369,N_2859);
nor U3640 (N_3640,N_2854,N_2616);
nand U3641 (N_3641,N_2377,N_2332);
xnor U3642 (N_3642,N_2772,N_2444);
nor U3643 (N_3643,N_2440,N_2809);
nand U3644 (N_3644,N_2937,N_2973);
xor U3645 (N_3645,N_2432,N_2740);
and U3646 (N_3646,N_2575,N_2994);
and U3647 (N_3647,N_2319,N_2317);
and U3648 (N_3648,N_2630,N_2528);
or U3649 (N_3649,N_2833,N_2355);
and U3650 (N_3650,N_2883,N_2387);
nor U3651 (N_3651,N_2623,N_2873);
nor U3652 (N_3652,N_2725,N_2499);
nor U3653 (N_3653,N_2735,N_2442);
nand U3654 (N_3654,N_2740,N_2482);
nand U3655 (N_3655,N_2508,N_2712);
nor U3656 (N_3656,N_2873,N_2348);
or U3657 (N_3657,N_2396,N_2977);
nand U3658 (N_3658,N_2999,N_2384);
nor U3659 (N_3659,N_2716,N_2281);
and U3660 (N_3660,N_2771,N_2926);
or U3661 (N_3661,N_2558,N_2509);
or U3662 (N_3662,N_2562,N_2952);
and U3663 (N_3663,N_2472,N_2749);
or U3664 (N_3664,N_2743,N_2377);
nand U3665 (N_3665,N_2856,N_2500);
xor U3666 (N_3666,N_2776,N_2663);
or U3667 (N_3667,N_2292,N_2919);
or U3668 (N_3668,N_2932,N_2409);
nor U3669 (N_3669,N_2624,N_2801);
nand U3670 (N_3670,N_2485,N_2322);
nand U3671 (N_3671,N_2811,N_2979);
nor U3672 (N_3672,N_2893,N_2485);
nand U3673 (N_3673,N_2638,N_2503);
and U3674 (N_3674,N_2257,N_2324);
xnor U3675 (N_3675,N_2499,N_2870);
nand U3676 (N_3676,N_2400,N_2479);
or U3677 (N_3677,N_2939,N_2924);
and U3678 (N_3678,N_2841,N_2342);
nand U3679 (N_3679,N_2812,N_2503);
and U3680 (N_3680,N_2821,N_2754);
and U3681 (N_3681,N_2469,N_2415);
xor U3682 (N_3682,N_2582,N_2486);
or U3683 (N_3683,N_2554,N_2345);
nand U3684 (N_3684,N_2774,N_2937);
xnor U3685 (N_3685,N_2386,N_2272);
and U3686 (N_3686,N_2559,N_2357);
nand U3687 (N_3687,N_2834,N_2399);
or U3688 (N_3688,N_2782,N_2792);
or U3689 (N_3689,N_2354,N_2864);
and U3690 (N_3690,N_2311,N_2329);
and U3691 (N_3691,N_2558,N_2267);
xnor U3692 (N_3692,N_2566,N_2770);
and U3693 (N_3693,N_2786,N_2859);
nand U3694 (N_3694,N_2596,N_2905);
and U3695 (N_3695,N_2972,N_2359);
or U3696 (N_3696,N_2524,N_2352);
nand U3697 (N_3697,N_2462,N_2327);
nand U3698 (N_3698,N_2985,N_2962);
xor U3699 (N_3699,N_2406,N_2781);
or U3700 (N_3700,N_2372,N_2622);
nand U3701 (N_3701,N_2557,N_2304);
xnor U3702 (N_3702,N_2985,N_2711);
xor U3703 (N_3703,N_2593,N_2819);
nand U3704 (N_3704,N_2888,N_2955);
xor U3705 (N_3705,N_2753,N_2907);
nor U3706 (N_3706,N_2936,N_2969);
and U3707 (N_3707,N_2922,N_2372);
nor U3708 (N_3708,N_2735,N_2280);
xor U3709 (N_3709,N_2610,N_2748);
or U3710 (N_3710,N_2569,N_2453);
nand U3711 (N_3711,N_2297,N_2784);
or U3712 (N_3712,N_2404,N_2658);
nor U3713 (N_3713,N_2254,N_2935);
nor U3714 (N_3714,N_2691,N_2819);
nand U3715 (N_3715,N_2352,N_2411);
xnor U3716 (N_3716,N_2285,N_2325);
nand U3717 (N_3717,N_2872,N_2409);
nor U3718 (N_3718,N_2867,N_2882);
or U3719 (N_3719,N_2333,N_2691);
and U3720 (N_3720,N_2632,N_2514);
and U3721 (N_3721,N_2455,N_2591);
xor U3722 (N_3722,N_2562,N_2417);
nor U3723 (N_3723,N_2363,N_2863);
xnor U3724 (N_3724,N_2996,N_2332);
or U3725 (N_3725,N_2469,N_2773);
nand U3726 (N_3726,N_2317,N_2979);
nand U3727 (N_3727,N_2527,N_2928);
nand U3728 (N_3728,N_2477,N_2498);
nand U3729 (N_3729,N_2890,N_2889);
and U3730 (N_3730,N_2480,N_2839);
nand U3731 (N_3731,N_2704,N_2907);
nand U3732 (N_3732,N_2357,N_2773);
nor U3733 (N_3733,N_2711,N_2281);
or U3734 (N_3734,N_2773,N_2463);
or U3735 (N_3735,N_2670,N_2866);
nor U3736 (N_3736,N_2486,N_2805);
and U3737 (N_3737,N_2351,N_2643);
or U3738 (N_3738,N_2614,N_2279);
or U3739 (N_3739,N_2712,N_2581);
and U3740 (N_3740,N_2919,N_2434);
xnor U3741 (N_3741,N_2634,N_2283);
nor U3742 (N_3742,N_2875,N_2772);
nand U3743 (N_3743,N_2397,N_2519);
nand U3744 (N_3744,N_2652,N_2670);
or U3745 (N_3745,N_2761,N_2902);
nor U3746 (N_3746,N_2560,N_2313);
nand U3747 (N_3747,N_2757,N_2818);
nor U3748 (N_3748,N_2628,N_2886);
xor U3749 (N_3749,N_2255,N_2693);
xor U3750 (N_3750,N_3474,N_3186);
and U3751 (N_3751,N_3091,N_3512);
xnor U3752 (N_3752,N_3323,N_3661);
and U3753 (N_3753,N_3353,N_3424);
and U3754 (N_3754,N_3171,N_3730);
xnor U3755 (N_3755,N_3033,N_3552);
or U3756 (N_3756,N_3471,N_3703);
xor U3757 (N_3757,N_3333,N_3510);
xnor U3758 (N_3758,N_3725,N_3056);
nor U3759 (N_3759,N_3090,N_3148);
nand U3760 (N_3760,N_3364,N_3008);
and U3761 (N_3761,N_3619,N_3487);
xnor U3762 (N_3762,N_3551,N_3629);
or U3763 (N_3763,N_3669,N_3178);
nor U3764 (N_3764,N_3531,N_3037);
xor U3765 (N_3765,N_3234,N_3155);
or U3766 (N_3766,N_3328,N_3034);
or U3767 (N_3767,N_3267,N_3406);
or U3768 (N_3768,N_3057,N_3276);
nor U3769 (N_3769,N_3292,N_3457);
or U3770 (N_3770,N_3615,N_3383);
nor U3771 (N_3771,N_3451,N_3075);
nor U3772 (N_3772,N_3385,N_3047);
xor U3773 (N_3773,N_3243,N_3278);
xor U3774 (N_3774,N_3442,N_3588);
or U3775 (N_3775,N_3724,N_3696);
nand U3776 (N_3776,N_3470,N_3183);
nand U3777 (N_3777,N_3310,N_3388);
xnor U3778 (N_3778,N_3735,N_3184);
and U3779 (N_3779,N_3676,N_3632);
or U3780 (N_3780,N_3108,N_3158);
and U3781 (N_3781,N_3702,N_3706);
xnor U3782 (N_3782,N_3347,N_3521);
xnor U3783 (N_3783,N_3045,N_3204);
nand U3784 (N_3784,N_3738,N_3105);
nand U3785 (N_3785,N_3192,N_3281);
or U3786 (N_3786,N_3550,N_3187);
or U3787 (N_3787,N_3340,N_3527);
nand U3788 (N_3788,N_3175,N_3371);
nand U3789 (N_3789,N_3579,N_3377);
xor U3790 (N_3790,N_3603,N_3680);
nor U3791 (N_3791,N_3199,N_3188);
nand U3792 (N_3792,N_3745,N_3461);
xor U3793 (N_3793,N_3672,N_3205);
nor U3794 (N_3794,N_3011,N_3475);
nor U3795 (N_3795,N_3386,N_3196);
and U3796 (N_3796,N_3226,N_3722);
nor U3797 (N_3797,N_3248,N_3421);
and U3798 (N_3798,N_3397,N_3093);
nand U3799 (N_3799,N_3502,N_3219);
nand U3800 (N_3800,N_3143,N_3013);
or U3801 (N_3801,N_3391,N_3410);
xnor U3802 (N_3802,N_3414,N_3417);
xnor U3803 (N_3803,N_3520,N_3060);
and U3804 (N_3804,N_3295,N_3287);
nor U3805 (N_3805,N_3541,N_3251);
nor U3806 (N_3806,N_3335,N_3288);
or U3807 (N_3807,N_3157,N_3538);
or U3808 (N_3808,N_3246,N_3712);
and U3809 (N_3809,N_3181,N_3220);
nor U3810 (N_3810,N_3587,N_3555);
nor U3811 (N_3811,N_3425,N_3433);
xor U3812 (N_3812,N_3170,N_3086);
nand U3813 (N_3813,N_3727,N_3304);
or U3814 (N_3814,N_3539,N_3350);
nor U3815 (N_3815,N_3100,N_3339);
and U3816 (N_3816,N_3000,N_3194);
nor U3817 (N_3817,N_3134,N_3465);
or U3818 (N_3818,N_3296,N_3098);
xor U3819 (N_3819,N_3411,N_3051);
or U3820 (N_3820,N_3644,N_3687);
nand U3821 (N_3821,N_3382,N_3711);
or U3822 (N_3822,N_3453,N_3628);
nor U3823 (N_3823,N_3577,N_3623);
and U3824 (N_3824,N_3341,N_3558);
nand U3825 (N_3825,N_3656,N_3543);
nand U3826 (N_3826,N_3467,N_3561);
nand U3827 (N_3827,N_3027,N_3375);
and U3828 (N_3828,N_3643,N_3572);
and U3829 (N_3829,N_3376,N_3069);
xor U3830 (N_3830,N_3492,N_3046);
xnor U3831 (N_3831,N_3351,N_3532);
xnor U3832 (N_3832,N_3673,N_3638);
xnor U3833 (N_3833,N_3431,N_3168);
nand U3834 (N_3834,N_3320,N_3537);
xnor U3835 (N_3835,N_3529,N_3720);
or U3836 (N_3836,N_3614,N_3023);
and U3837 (N_3837,N_3124,N_3079);
nand U3838 (N_3838,N_3307,N_3118);
nand U3839 (N_3839,N_3260,N_3159);
nor U3840 (N_3840,N_3454,N_3648);
nor U3841 (N_3841,N_3218,N_3518);
xnor U3842 (N_3842,N_3272,N_3161);
and U3843 (N_3843,N_3334,N_3262);
nand U3844 (N_3844,N_3122,N_3139);
nor U3845 (N_3845,N_3390,N_3526);
or U3846 (N_3846,N_3244,N_3275);
nand U3847 (N_3847,N_3191,N_3257);
nand U3848 (N_3848,N_3040,N_3324);
or U3849 (N_3849,N_3713,N_3140);
nor U3850 (N_3850,N_3096,N_3416);
nor U3851 (N_3851,N_3338,N_3035);
xnor U3852 (N_3852,N_3400,N_3723);
or U3853 (N_3853,N_3654,N_3142);
or U3854 (N_3854,N_3372,N_3115);
and U3855 (N_3855,N_3022,N_3675);
nand U3856 (N_3856,N_3437,N_3315);
xor U3857 (N_3857,N_3209,N_3015);
nor U3858 (N_3858,N_3409,N_3686);
or U3859 (N_3859,N_3683,N_3326);
and U3860 (N_3860,N_3349,N_3432);
nor U3861 (N_3861,N_3360,N_3065);
and U3862 (N_3862,N_3695,N_3700);
xnor U3863 (N_3863,N_3007,N_3710);
or U3864 (N_3864,N_3741,N_3238);
nand U3865 (N_3865,N_3516,N_3571);
and U3866 (N_3866,N_3059,N_3601);
nor U3867 (N_3867,N_3355,N_3228);
nand U3868 (N_3868,N_3121,N_3744);
or U3869 (N_3869,N_3380,N_3670);
and U3870 (N_3870,N_3151,N_3441);
nor U3871 (N_3871,N_3450,N_3742);
nand U3872 (N_3872,N_3627,N_3305);
nand U3873 (N_3873,N_3210,N_3112);
nor U3874 (N_3874,N_3519,N_3428);
nor U3875 (N_3875,N_3036,N_3484);
and U3876 (N_3876,N_3041,N_3277);
xor U3877 (N_3877,N_3594,N_3581);
and U3878 (N_3878,N_3708,N_3524);
or U3879 (N_3879,N_3265,N_3255);
or U3880 (N_3880,N_3429,N_3678);
or U3881 (N_3881,N_3651,N_3068);
nand U3882 (N_3882,N_3229,N_3482);
xnor U3883 (N_3883,N_3689,N_3256);
nor U3884 (N_3884,N_3418,N_3449);
nor U3885 (N_3885,N_3299,N_3652);
xor U3886 (N_3886,N_3133,N_3247);
and U3887 (N_3887,N_3331,N_3662);
and U3888 (N_3888,N_3358,N_3200);
nor U3889 (N_3889,N_3591,N_3213);
or U3890 (N_3890,N_3602,N_3279);
and U3891 (N_3891,N_3554,N_3640);
xnor U3892 (N_3892,N_3719,N_3458);
nand U3893 (N_3893,N_3620,N_3354);
or U3894 (N_3894,N_3309,N_3317);
nand U3895 (N_3895,N_3674,N_3180);
and U3896 (N_3896,N_3154,N_3740);
nor U3897 (N_3897,N_3547,N_3490);
xnor U3898 (N_3898,N_3626,N_3663);
nand U3899 (N_3899,N_3359,N_3387);
xor U3900 (N_3900,N_3621,N_3690);
and U3901 (N_3901,N_3254,N_3314);
xnor U3902 (N_3902,N_3009,N_3422);
or U3903 (N_3903,N_3636,N_3312);
and U3904 (N_3904,N_3381,N_3645);
nand U3905 (N_3905,N_3066,N_3479);
and U3906 (N_3906,N_3513,N_3500);
or U3907 (N_3907,N_3608,N_3448);
nand U3908 (N_3908,N_3052,N_3348);
or U3909 (N_3909,N_3293,N_3396);
or U3910 (N_3910,N_3363,N_3478);
nor U3911 (N_3911,N_3352,N_3123);
nor U3912 (N_3912,N_3156,N_3217);
nor U3913 (N_3913,N_3596,N_3094);
or U3914 (N_3914,N_3172,N_3061);
xor U3915 (N_3915,N_3286,N_3102);
xor U3916 (N_3916,N_3024,N_3495);
or U3917 (N_3917,N_3503,N_3370);
nor U3918 (N_3918,N_3497,N_3523);
nor U3919 (N_3919,N_3600,N_3111);
nand U3920 (N_3920,N_3245,N_3426);
or U3921 (N_3921,N_3447,N_3699);
or U3922 (N_3922,N_3622,N_3707);
nand U3923 (N_3923,N_3044,N_3542);
nor U3924 (N_3924,N_3634,N_3684);
or U3925 (N_3925,N_3736,N_3266);
or U3926 (N_3926,N_3250,N_3419);
nand U3927 (N_3927,N_3625,N_3473);
and U3928 (N_3928,N_3544,N_3164);
xnor U3929 (N_3929,N_3010,N_3055);
nor U3930 (N_3930,N_3198,N_3104);
or U3931 (N_3931,N_3249,N_3223);
nand U3932 (N_3932,N_3452,N_3412);
xnor U3933 (N_3933,N_3427,N_3235);
or U3934 (N_3934,N_3574,N_3677);
nand U3935 (N_3935,N_3368,N_3085);
nand U3936 (N_3936,N_3095,N_3322);
nor U3937 (N_3937,N_3336,N_3241);
nand U3938 (N_3938,N_3746,N_3087);
xor U3939 (N_3939,N_3264,N_3076);
or U3940 (N_3940,N_3081,N_3545);
and U3941 (N_3941,N_3717,N_3477);
nor U3942 (N_3942,N_3599,N_3062);
xnor U3943 (N_3943,N_3166,N_3119);
nor U3944 (N_3944,N_3273,N_3446);
and U3945 (N_3945,N_3197,N_3070);
or U3946 (N_3946,N_3728,N_3053);
xor U3947 (N_3947,N_3019,N_3297);
nand U3948 (N_3948,N_3697,N_3659);
or U3949 (N_3949,N_3704,N_3568);
or U3950 (N_3950,N_3378,N_3570);
nor U3951 (N_3951,N_3459,N_3405);
nand U3952 (N_3952,N_3236,N_3514);
nor U3953 (N_3953,N_3083,N_3444);
xnor U3954 (N_3954,N_3089,N_3306);
or U3955 (N_3955,N_3384,N_3329);
and U3956 (N_3956,N_3120,N_3612);
xnor U3957 (N_3957,N_3014,N_3284);
or U3958 (N_3958,N_3576,N_3285);
nor U3959 (N_3959,N_3435,N_3099);
and U3960 (N_3960,N_3026,N_3101);
nor U3961 (N_3961,N_3274,N_3580);
and U3962 (N_3962,N_3110,N_3508);
xnor U3963 (N_3963,N_3694,N_3145);
nand U3964 (N_3964,N_3438,N_3589);
nand U3965 (N_3965,N_3038,N_3506);
and U3966 (N_3966,N_3637,N_3107);
and U3967 (N_3967,N_3650,N_3436);
nand U3968 (N_3968,N_3567,N_3361);
or U3969 (N_3969,N_3595,N_3660);
or U3970 (N_3970,N_3682,N_3729);
xnor U3971 (N_3971,N_3413,N_3227);
or U3972 (N_3972,N_3714,N_3592);
nand U3973 (N_3973,N_3001,N_3379);
and U3974 (N_3974,N_3434,N_3671);
nor U3975 (N_3975,N_3127,N_3501);
xor U3976 (N_3976,N_3269,N_3135);
and U3977 (N_3977,N_3106,N_3582);
nand U3978 (N_3978,N_3511,N_3504);
or U3979 (N_3979,N_3731,N_3395);
or U3980 (N_3980,N_3282,N_3049);
or U3981 (N_3981,N_3709,N_3207);
nand U3982 (N_3982,N_3017,N_3613);
nand U3983 (N_3983,N_3646,N_3463);
or U3984 (N_3984,N_3734,N_3182);
xor U3985 (N_3985,N_3679,N_3562);
xor U3986 (N_3986,N_3617,N_3404);
or U3987 (N_3987,N_3721,N_3546);
or U3988 (N_3988,N_3583,N_3462);
and U3989 (N_3989,N_3138,N_3030);
nor U3990 (N_3990,N_3584,N_3018);
nand U3991 (N_3991,N_3560,N_3607);
or U3992 (N_3992,N_3499,N_3743);
nor U3993 (N_3993,N_3125,N_3058);
nand U3994 (N_3994,N_3715,N_3165);
or U3995 (N_3995,N_3189,N_3630);
nand U3996 (N_3996,N_3193,N_3153);
or U3997 (N_3997,N_3491,N_3149);
nand U3998 (N_3998,N_3162,N_3590);
and U3999 (N_3999,N_3002,N_3103);
and U4000 (N_4000,N_3618,N_3169);
or U4001 (N_4001,N_3078,N_3203);
or U4002 (N_4002,N_3394,N_3150);
nor U4003 (N_4003,N_3642,N_3319);
nand U4004 (N_4004,N_3144,N_3748);
and U4005 (N_4005,N_3214,N_3283);
or U4006 (N_4006,N_3559,N_3747);
nand U4007 (N_4007,N_3088,N_3318);
xnor U4008 (N_4008,N_3224,N_3530);
nor U4009 (N_4009,N_3252,N_3667);
and U4010 (N_4010,N_3496,N_3476);
xnor U4011 (N_4011,N_3303,N_3016);
or U4012 (N_4012,N_3598,N_3050);
and U4013 (N_4013,N_3401,N_3606);
nor U4014 (N_4014,N_3367,N_3649);
or U4015 (N_4015,N_3536,N_3486);
and U4016 (N_4016,N_3298,N_3566);
xnor U4017 (N_4017,N_3136,N_3215);
nand U4018 (N_4018,N_3407,N_3097);
xor U4019 (N_4019,N_3393,N_3494);
nor U4020 (N_4020,N_3485,N_3517);
nand U4021 (N_4021,N_3633,N_3698);
and U4022 (N_4022,N_3525,N_3029);
nor U4023 (N_4023,N_3374,N_3006);
nand U4024 (N_4024,N_3109,N_3167);
xor U4025 (N_4025,N_3681,N_3268);
nand U4026 (N_4026,N_3263,N_3420);
and U4027 (N_4027,N_3032,N_3445);
nand U4028 (N_4028,N_3232,N_3553);
nand U4029 (N_4029,N_3160,N_3259);
and U4030 (N_4030,N_3597,N_3732);
nor U4031 (N_4031,N_3239,N_3020);
xor U4032 (N_4032,N_3460,N_3399);
or U4033 (N_4033,N_3222,N_3739);
nor U4034 (N_4034,N_3366,N_3240);
and U4035 (N_4035,N_3258,N_3356);
nand U4036 (N_4036,N_3332,N_3179);
nor U4037 (N_4037,N_3655,N_3357);
xor U4038 (N_4038,N_3593,N_3337);
xnor U4039 (N_4039,N_3201,N_3126);
nand U4040 (N_4040,N_3321,N_3130);
or U4041 (N_4041,N_3208,N_3177);
nor U4042 (N_4042,N_3141,N_3084);
nor U4043 (N_4043,N_3290,N_3311);
and U4044 (N_4044,N_3392,N_3345);
xor U4045 (N_4045,N_3609,N_3330);
xor U4046 (N_4046,N_3564,N_3389);
or U4047 (N_4047,N_3147,N_3117);
xor U4048 (N_4048,N_3131,N_3472);
or U4049 (N_4049,N_3624,N_3693);
nor U4050 (N_4050,N_3430,N_3469);
and U4051 (N_4051,N_3611,N_3585);
nand U4052 (N_4052,N_3221,N_3152);
nor U4053 (N_4053,N_3507,N_3185);
and U4054 (N_4054,N_3190,N_3586);
and U4055 (N_4055,N_3505,N_3344);
xnor U4056 (N_4056,N_3569,N_3291);
nand U4057 (N_4057,N_3128,N_3408);
xor U4058 (N_4058,N_3028,N_3233);
and U4059 (N_4059,N_3173,N_3231);
or U4060 (N_4060,N_3074,N_3515);
or U4061 (N_4061,N_3664,N_3327);
or U4062 (N_4062,N_3666,N_3261);
nor U4063 (N_4063,N_3692,N_3080);
nand U4064 (N_4064,N_3528,N_3365);
and U4065 (N_4065,N_3316,N_3423);
and U4066 (N_4066,N_3493,N_3003);
or U4067 (N_4067,N_3202,N_3216);
nand U4068 (N_4068,N_3362,N_3575);
xnor U4069 (N_4069,N_3132,N_3701);
nor U4070 (N_4070,N_3685,N_3373);
xor U4071 (N_4071,N_3073,N_3114);
xor U4072 (N_4072,N_3439,N_3289);
nor U4073 (N_4073,N_3534,N_3737);
nand U4074 (N_4074,N_3346,N_3610);
and U4075 (N_4075,N_3212,N_3705);
xor U4076 (N_4076,N_3031,N_3653);
xnor U4077 (N_4077,N_3540,N_3398);
xnor U4078 (N_4078,N_3113,N_3402);
nand U4079 (N_4079,N_3733,N_3325);
nand U4080 (N_4080,N_3498,N_3242);
nor U4081 (N_4081,N_3043,N_3129);
nand U4082 (N_4082,N_3464,N_3647);
or U4083 (N_4083,N_3468,N_3206);
nor U4084 (N_4084,N_3294,N_3369);
xnor U4085 (N_4085,N_3726,N_3021);
and U4086 (N_4086,N_3176,N_3071);
and U4087 (N_4087,N_3616,N_3082);
nand U4088 (N_4088,N_3556,N_3509);
nor U4089 (N_4089,N_3481,N_3456);
and U4090 (N_4090,N_3004,N_3749);
and U4091 (N_4091,N_3549,N_3688);
xnor U4092 (N_4092,N_3573,N_3565);
nand U4093 (N_4093,N_3535,N_3691);
nor U4094 (N_4094,N_3657,N_3483);
and U4095 (N_4095,N_3489,N_3280);
and U4096 (N_4096,N_3308,N_3237);
or U4097 (N_4097,N_3480,N_3146);
xor U4098 (N_4098,N_3658,N_3533);
nor U4099 (N_4099,N_3342,N_3072);
or U4100 (N_4100,N_3302,N_3137);
and U4101 (N_4101,N_3270,N_3578);
xor U4102 (N_4102,N_3665,N_3163);
nor U4103 (N_4103,N_3605,N_3300);
nor U4104 (N_4104,N_3313,N_3639);
xnor U4105 (N_4105,N_3271,N_3005);
and U4106 (N_4106,N_3455,N_3563);
or U4107 (N_4107,N_3548,N_3225);
xor U4108 (N_4108,N_3064,N_3716);
xnor U4109 (N_4109,N_3063,N_3012);
nand U4110 (N_4110,N_3067,N_3025);
or U4111 (N_4111,N_3466,N_3635);
xnor U4112 (N_4112,N_3230,N_3557);
nor U4113 (N_4113,N_3092,N_3174);
or U4114 (N_4114,N_3211,N_3042);
and U4115 (N_4115,N_3301,N_3443);
xnor U4116 (N_4116,N_3718,N_3048);
nor U4117 (N_4117,N_3641,N_3403);
or U4118 (N_4118,N_3440,N_3195);
or U4119 (N_4119,N_3522,N_3343);
nand U4120 (N_4120,N_3604,N_3253);
nand U4121 (N_4121,N_3488,N_3631);
xnor U4122 (N_4122,N_3077,N_3054);
nand U4123 (N_4123,N_3039,N_3668);
nor U4124 (N_4124,N_3116,N_3415);
or U4125 (N_4125,N_3597,N_3113);
nand U4126 (N_4126,N_3078,N_3721);
nand U4127 (N_4127,N_3205,N_3142);
nor U4128 (N_4128,N_3445,N_3331);
nand U4129 (N_4129,N_3013,N_3058);
nand U4130 (N_4130,N_3562,N_3036);
xor U4131 (N_4131,N_3344,N_3625);
nand U4132 (N_4132,N_3181,N_3547);
xor U4133 (N_4133,N_3164,N_3227);
xor U4134 (N_4134,N_3026,N_3188);
nor U4135 (N_4135,N_3248,N_3163);
nor U4136 (N_4136,N_3559,N_3537);
nand U4137 (N_4137,N_3385,N_3153);
or U4138 (N_4138,N_3344,N_3175);
and U4139 (N_4139,N_3362,N_3171);
nor U4140 (N_4140,N_3519,N_3550);
and U4141 (N_4141,N_3345,N_3328);
or U4142 (N_4142,N_3226,N_3509);
nor U4143 (N_4143,N_3658,N_3209);
nand U4144 (N_4144,N_3112,N_3104);
xnor U4145 (N_4145,N_3693,N_3402);
or U4146 (N_4146,N_3553,N_3396);
nor U4147 (N_4147,N_3203,N_3742);
nor U4148 (N_4148,N_3038,N_3543);
nor U4149 (N_4149,N_3516,N_3414);
and U4150 (N_4150,N_3485,N_3701);
xnor U4151 (N_4151,N_3440,N_3450);
nor U4152 (N_4152,N_3334,N_3688);
xor U4153 (N_4153,N_3683,N_3697);
and U4154 (N_4154,N_3294,N_3132);
and U4155 (N_4155,N_3490,N_3380);
and U4156 (N_4156,N_3450,N_3346);
or U4157 (N_4157,N_3218,N_3459);
nor U4158 (N_4158,N_3624,N_3181);
xnor U4159 (N_4159,N_3065,N_3397);
nand U4160 (N_4160,N_3043,N_3180);
and U4161 (N_4161,N_3246,N_3349);
nor U4162 (N_4162,N_3157,N_3019);
nor U4163 (N_4163,N_3070,N_3615);
nand U4164 (N_4164,N_3295,N_3461);
or U4165 (N_4165,N_3374,N_3041);
nand U4166 (N_4166,N_3122,N_3663);
nor U4167 (N_4167,N_3553,N_3341);
nand U4168 (N_4168,N_3488,N_3124);
xnor U4169 (N_4169,N_3531,N_3404);
or U4170 (N_4170,N_3228,N_3322);
and U4171 (N_4171,N_3176,N_3646);
nor U4172 (N_4172,N_3347,N_3531);
and U4173 (N_4173,N_3144,N_3603);
xnor U4174 (N_4174,N_3496,N_3497);
nor U4175 (N_4175,N_3127,N_3590);
or U4176 (N_4176,N_3381,N_3330);
or U4177 (N_4177,N_3603,N_3256);
or U4178 (N_4178,N_3002,N_3596);
nand U4179 (N_4179,N_3589,N_3437);
or U4180 (N_4180,N_3440,N_3358);
xnor U4181 (N_4181,N_3484,N_3219);
and U4182 (N_4182,N_3359,N_3144);
nand U4183 (N_4183,N_3641,N_3369);
or U4184 (N_4184,N_3645,N_3345);
nor U4185 (N_4185,N_3032,N_3449);
xnor U4186 (N_4186,N_3693,N_3022);
nand U4187 (N_4187,N_3561,N_3608);
and U4188 (N_4188,N_3499,N_3150);
or U4189 (N_4189,N_3081,N_3051);
nand U4190 (N_4190,N_3526,N_3506);
and U4191 (N_4191,N_3683,N_3428);
and U4192 (N_4192,N_3413,N_3577);
and U4193 (N_4193,N_3201,N_3466);
xnor U4194 (N_4194,N_3137,N_3065);
xor U4195 (N_4195,N_3448,N_3074);
and U4196 (N_4196,N_3221,N_3096);
nor U4197 (N_4197,N_3406,N_3747);
nand U4198 (N_4198,N_3494,N_3244);
nand U4199 (N_4199,N_3631,N_3546);
xnor U4200 (N_4200,N_3164,N_3238);
and U4201 (N_4201,N_3015,N_3692);
xnor U4202 (N_4202,N_3445,N_3748);
and U4203 (N_4203,N_3737,N_3194);
xor U4204 (N_4204,N_3290,N_3397);
nand U4205 (N_4205,N_3618,N_3677);
xor U4206 (N_4206,N_3347,N_3032);
or U4207 (N_4207,N_3712,N_3506);
xnor U4208 (N_4208,N_3654,N_3065);
and U4209 (N_4209,N_3166,N_3322);
or U4210 (N_4210,N_3625,N_3454);
nor U4211 (N_4211,N_3024,N_3574);
nand U4212 (N_4212,N_3391,N_3208);
nand U4213 (N_4213,N_3512,N_3109);
and U4214 (N_4214,N_3171,N_3053);
and U4215 (N_4215,N_3379,N_3022);
or U4216 (N_4216,N_3363,N_3583);
nand U4217 (N_4217,N_3104,N_3396);
xor U4218 (N_4218,N_3101,N_3176);
nand U4219 (N_4219,N_3595,N_3653);
and U4220 (N_4220,N_3117,N_3105);
nor U4221 (N_4221,N_3079,N_3496);
xor U4222 (N_4222,N_3498,N_3723);
or U4223 (N_4223,N_3748,N_3086);
xor U4224 (N_4224,N_3616,N_3246);
nand U4225 (N_4225,N_3396,N_3559);
or U4226 (N_4226,N_3211,N_3582);
and U4227 (N_4227,N_3035,N_3268);
xnor U4228 (N_4228,N_3556,N_3397);
or U4229 (N_4229,N_3400,N_3743);
or U4230 (N_4230,N_3685,N_3233);
or U4231 (N_4231,N_3614,N_3106);
nor U4232 (N_4232,N_3402,N_3332);
and U4233 (N_4233,N_3685,N_3599);
xnor U4234 (N_4234,N_3444,N_3071);
or U4235 (N_4235,N_3311,N_3375);
nor U4236 (N_4236,N_3612,N_3403);
xnor U4237 (N_4237,N_3596,N_3485);
xor U4238 (N_4238,N_3091,N_3034);
nor U4239 (N_4239,N_3345,N_3332);
and U4240 (N_4240,N_3379,N_3279);
xnor U4241 (N_4241,N_3278,N_3469);
and U4242 (N_4242,N_3335,N_3590);
or U4243 (N_4243,N_3157,N_3625);
nor U4244 (N_4244,N_3190,N_3020);
nand U4245 (N_4245,N_3474,N_3728);
nand U4246 (N_4246,N_3022,N_3747);
or U4247 (N_4247,N_3575,N_3193);
nor U4248 (N_4248,N_3256,N_3061);
or U4249 (N_4249,N_3357,N_3358);
and U4250 (N_4250,N_3529,N_3659);
xor U4251 (N_4251,N_3330,N_3075);
xor U4252 (N_4252,N_3077,N_3727);
or U4253 (N_4253,N_3059,N_3389);
or U4254 (N_4254,N_3090,N_3717);
xor U4255 (N_4255,N_3074,N_3196);
nand U4256 (N_4256,N_3543,N_3740);
nor U4257 (N_4257,N_3263,N_3160);
xor U4258 (N_4258,N_3668,N_3310);
xor U4259 (N_4259,N_3411,N_3476);
or U4260 (N_4260,N_3624,N_3557);
and U4261 (N_4261,N_3068,N_3553);
or U4262 (N_4262,N_3299,N_3401);
nand U4263 (N_4263,N_3304,N_3104);
and U4264 (N_4264,N_3311,N_3085);
xnor U4265 (N_4265,N_3244,N_3682);
nand U4266 (N_4266,N_3073,N_3227);
nor U4267 (N_4267,N_3737,N_3575);
and U4268 (N_4268,N_3660,N_3484);
xnor U4269 (N_4269,N_3282,N_3713);
nand U4270 (N_4270,N_3309,N_3570);
nor U4271 (N_4271,N_3372,N_3196);
nor U4272 (N_4272,N_3095,N_3033);
xor U4273 (N_4273,N_3745,N_3418);
and U4274 (N_4274,N_3562,N_3268);
and U4275 (N_4275,N_3174,N_3309);
xnor U4276 (N_4276,N_3441,N_3034);
xnor U4277 (N_4277,N_3431,N_3639);
and U4278 (N_4278,N_3503,N_3736);
or U4279 (N_4279,N_3404,N_3130);
or U4280 (N_4280,N_3044,N_3408);
nor U4281 (N_4281,N_3157,N_3026);
xnor U4282 (N_4282,N_3118,N_3238);
and U4283 (N_4283,N_3148,N_3466);
and U4284 (N_4284,N_3634,N_3203);
xor U4285 (N_4285,N_3512,N_3275);
and U4286 (N_4286,N_3495,N_3235);
and U4287 (N_4287,N_3051,N_3035);
or U4288 (N_4288,N_3546,N_3589);
and U4289 (N_4289,N_3580,N_3475);
nand U4290 (N_4290,N_3404,N_3708);
or U4291 (N_4291,N_3365,N_3081);
xor U4292 (N_4292,N_3546,N_3616);
or U4293 (N_4293,N_3037,N_3636);
nand U4294 (N_4294,N_3569,N_3242);
nor U4295 (N_4295,N_3272,N_3391);
nor U4296 (N_4296,N_3556,N_3370);
and U4297 (N_4297,N_3438,N_3637);
nor U4298 (N_4298,N_3262,N_3613);
or U4299 (N_4299,N_3521,N_3331);
and U4300 (N_4300,N_3329,N_3387);
and U4301 (N_4301,N_3712,N_3473);
nor U4302 (N_4302,N_3421,N_3467);
nor U4303 (N_4303,N_3311,N_3495);
nor U4304 (N_4304,N_3367,N_3191);
nor U4305 (N_4305,N_3341,N_3251);
nor U4306 (N_4306,N_3719,N_3265);
or U4307 (N_4307,N_3737,N_3673);
nand U4308 (N_4308,N_3181,N_3147);
and U4309 (N_4309,N_3702,N_3200);
nand U4310 (N_4310,N_3391,N_3523);
or U4311 (N_4311,N_3226,N_3049);
and U4312 (N_4312,N_3259,N_3630);
and U4313 (N_4313,N_3384,N_3480);
and U4314 (N_4314,N_3488,N_3143);
nand U4315 (N_4315,N_3434,N_3732);
nor U4316 (N_4316,N_3014,N_3248);
or U4317 (N_4317,N_3482,N_3078);
and U4318 (N_4318,N_3378,N_3224);
or U4319 (N_4319,N_3148,N_3066);
xnor U4320 (N_4320,N_3028,N_3541);
xor U4321 (N_4321,N_3383,N_3320);
nor U4322 (N_4322,N_3300,N_3335);
xor U4323 (N_4323,N_3648,N_3130);
nor U4324 (N_4324,N_3301,N_3051);
nor U4325 (N_4325,N_3005,N_3340);
nor U4326 (N_4326,N_3373,N_3184);
and U4327 (N_4327,N_3321,N_3128);
or U4328 (N_4328,N_3569,N_3453);
and U4329 (N_4329,N_3379,N_3038);
nor U4330 (N_4330,N_3387,N_3706);
or U4331 (N_4331,N_3406,N_3472);
nand U4332 (N_4332,N_3179,N_3562);
and U4333 (N_4333,N_3440,N_3377);
nand U4334 (N_4334,N_3656,N_3092);
and U4335 (N_4335,N_3084,N_3070);
nor U4336 (N_4336,N_3091,N_3364);
or U4337 (N_4337,N_3498,N_3739);
xor U4338 (N_4338,N_3356,N_3463);
nor U4339 (N_4339,N_3113,N_3452);
and U4340 (N_4340,N_3307,N_3168);
xnor U4341 (N_4341,N_3225,N_3215);
and U4342 (N_4342,N_3694,N_3467);
and U4343 (N_4343,N_3491,N_3427);
nor U4344 (N_4344,N_3162,N_3222);
or U4345 (N_4345,N_3503,N_3063);
and U4346 (N_4346,N_3109,N_3716);
nand U4347 (N_4347,N_3560,N_3729);
xor U4348 (N_4348,N_3013,N_3622);
nand U4349 (N_4349,N_3246,N_3423);
nand U4350 (N_4350,N_3542,N_3720);
or U4351 (N_4351,N_3719,N_3079);
nor U4352 (N_4352,N_3319,N_3522);
nand U4353 (N_4353,N_3059,N_3254);
nand U4354 (N_4354,N_3061,N_3715);
xor U4355 (N_4355,N_3552,N_3610);
nor U4356 (N_4356,N_3675,N_3546);
nor U4357 (N_4357,N_3271,N_3478);
nor U4358 (N_4358,N_3252,N_3377);
or U4359 (N_4359,N_3734,N_3017);
xnor U4360 (N_4360,N_3292,N_3382);
and U4361 (N_4361,N_3288,N_3357);
and U4362 (N_4362,N_3685,N_3457);
or U4363 (N_4363,N_3275,N_3069);
and U4364 (N_4364,N_3267,N_3732);
nand U4365 (N_4365,N_3500,N_3611);
or U4366 (N_4366,N_3430,N_3706);
nand U4367 (N_4367,N_3011,N_3722);
xor U4368 (N_4368,N_3318,N_3353);
xor U4369 (N_4369,N_3124,N_3434);
and U4370 (N_4370,N_3176,N_3191);
xor U4371 (N_4371,N_3186,N_3302);
and U4372 (N_4372,N_3233,N_3118);
xor U4373 (N_4373,N_3555,N_3096);
nand U4374 (N_4374,N_3251,N_3100);
nand U4375 (N_4375,N_3473,N_3322);
nor U4376 (N_4376,N_3326,N_3059);
nand U4377 (N_4377,N_3355,N_3578);
or U4378 (N_4378,N_3572,N_3695);
nor U4379 (N_4379,N_3234,N_3222);
nand U4380 (N_4380,N_3702,N_3712);
nand U4381 (N_4381,N_3300,N_3476);
and U4382 (N_4382,N_3468,N_3159);
nand U4383 (N_4383,N_3156,N_3479);
or U4384 (N_4384,N_3489,N_3532);
or U4385 (N_4385,N_3629,N_3661);
xnor U4386 (N_4386,N_3728,N_3218);
xor U4387 (N_4387,N_3085,N_3199);
and U4388 (N_4388,N_3429,N_3312);
or U4389 (N_4389,N_3126,N_3246);
or U4390 (N_4390,N_3087,N_3413);
nand U4391 (N_4391,N_3021,N_3336);
nand U4392 (N_4392,N_3660,N_3480);
xor U4393 (N_4393,N_3099,N_3355);
nor U4394 (N_4394,N_3414,N_3198);
or U4395 (N_4395,N_3461,N_3419);
and U4396 (N_4396,N_3145,N_3463);
xor U4397 (N_4397,N_3579,N_3635);
nor U4398 (N_4398,N_3121,N_3494);
xor U4399 (N_4399,N_3135,N_3229);
nand U4400 (N_4400,N_3185,N_3081);
nand U4401 (N_4401,N_3488,N_3440);
xor U4402 (N_4402,N_3171,N_3059);
nor U4403 (N_4403,N_3406,N_3435);
or U4404 (N_4404,N_3524,N_3539);
or U4405 (N_4405,N_3174,N_3473);
or U4406 (N_4406,N_3313,N_3656);
and U4407 (N_4407,N_3470,N_3194);
or U4408 (N_4408,N_3629,N_3736);
nand U4409 (N_4409,N_3370,N_3700);
and U4410 (N_4410,N_3687,N_3684);
xnor U4411 (N_4411,N_3214,N_3725);
and U4412 (N_4412,N_3414,N_3523);
nor U4413 (N_4413,N_3412,N_3018);
or U4414 (N_4414,N_3431,N_3526);
or U4415 (N_4415,N_3118,N_3322);
xor U4416 (N_4416,N_3543,N_3339);
and U4417 (N_4417,N_3165,N_3681);
and U4418 (N_4418,N_3337,N_3632);
nand U4419 (N_4419,N_3414,N_3556);
nand U4420 (N_4420,N_3679,N_3726);
nand U4421 (N_4421,N_3491,N_3659);
or U4422 (N_4422,N_3067,N_3133);
xnor U4423 (N_4423,N_3693,N_3644);
or U4424 (N_4424,N_3401,N_3286);
xnor U4425 (N_4425,N_3580,N_3231);
and U4426 (N_4426,N_3364,N_3728);
and U4427 (N_4427,N_3546,N_3537);
nand U4428 (N_4428,N_3602,N_3396);
nor U4429 (N_4429,N_3747,N_3259);
or U4430 (N_4430,N_3166,N_3678);
or U4431 (N_4431,N_3349,N_3720);
or U4432 (N_4432,N_3560,N_3056);
or U4433 (N_4433,N_3437,N_3104);
and U4434 (N_4434,N_3363,N_3013);
and U4435 (N_4435,N_3168,N_3186);
or U4436 (N_4436,N_3393,N_3353);
xor U4437 (N_4437,N_3191,N_3364);
or U4438 (N_4438,N_3277,N_3265);
and U4439 (N_4439,N_3364,N_3431);
or U4440 (N_4440,N_3130,N_3724);
xnor U4441 (N_4441,N_3679,N_3206);
nor U4442 (N_4442,N_3584,N_3437);
nor U4443 (N_4443,N_3323,N_3119);
nor U4444 (N_4444,N_3703,N_3125);
nor U4445 (N_4445,N_3146,N_3327);
nor U4446 (N_4446,N_3721,N_3459);
nand U4447 (N_4447,N_3220,N_3146);
nand U4448 (N_4448,N_3333,N_3638);
nor U4449 (N_4449,N_3218,N_3517);
or U4450 (N_4450,N_3396,N_3103);
and U4451 (N_4451,N_3669,N_3621);
xor U4452 (N_4452,N_3061,N_3495);
xor U4453 (N_4453,N_3565,N_3101);
nor U4454 (N_4454,N_3538,N_3161);
nor U4455 (N_4455,N_3700,N_3630);
nor U4456 (N_4456,N_3176,N_3741);
and U4457 (N_4457,N_3095,N_3410);
nand U4458 (N_4458,N_3258,N_3583);
xor U4459 (N_4459,N_3020,N_3286);
or U4460 (N_4460,N_3692,N_3288);
or U4461 (N_4461,N_3479,N_3343);
nand U4462 (N_4462,N_3171,N_3551);
nor U4463 (N_4463,N_3196,N_3334);
nor U4464 (N_4464,N_3449,N_3096);
and U4465 (N_4465,N_3056,N_3289);
and U4466 (N_4466,N_3096,N_3656);
and U4467 (N_4467,N_3473,N_3644);
xnor U4468 (N_4468,N_3183,N_3502);
or U4469 (N_4469,N_3187,N_3619);
nand U4470 (N_4470,N_3067,N_3503);
and U4471 (N_4471,N_3518,N_3747);
or U4472 (N_4472,N_3065,N_3189);
xor U4473 (N_4473,N_3686,N_3631);
nor U4474 (N_4474,N_3095,N_3411);
and U4475 (N_4475,N_3650,N_3741);
nor U4476 (N_4476,N_3559,N_3543);
nor U4477 (N_4477,N_3537,N_3606);
and U4478 (N_4478,N_3450,N_3218);
and U4479 (N_4479,N_3369,N_3051);
nor U4480 (N_4480,N_3329,N_3609);
and U4481 (N_4481,N_3508,N_3495);
xnor U4482 (N_4482,N_3069,N_3313);
xor U4483 (N_4483,N_3605,N_3397);
nor U4484 (N_4484,N_3039,N_3196);
nand U4485 (N_4485,N_3439,N_3452);
or U4486 (N_4486,N_3069,N_3417);
nor U4487 (N_4487,N_3077,N_3434);
xnor U4488 (N_4488,N_3139,N_3692);
xor U4489 (N_4489,N_3702,N_3519);
or U4490 (N_4490,N_3227,N_3270);
nand U4491 (N_4491,N_3165,N_3464);
or U4492 (N_4492,N_3569,N_3613);
nand U4493 (N_4493,N_3000,N_3516);
xor U4494 (N_4494,N_3443,N_3175);
nand U4495 (N_4495,N_3731,N_3436);
nand U4496 (N_4496,N_3141,N_3396);
nor U4497 (N_4497,N_3393,N_3004);
or U4498 (N_4498,N_3238,N_3147);
and U4499 (N_4499,N_3157,N_3078);
and U4500 (N_4500,N_4118,N_4014);
nor U4501 (N_4501,N_4003,N_4447);
or U4502 (N_4502,N_4377,N_3868);
nand U4503 (N_4503,N_3834,N_3801);
xnor U4504 (N_4504,N_3780,N_4052);
or U4505 (N_4505,N_4232,N_3869);
or U4506 (N_4506,N_4492,N_4170);
xnor U4507 (N_4507,N_3971,N_4060);
or U4508 (N_4508,N_3769,N_4278);
and U4509 (N_4509,N_3792,N_3836);
xor U4510 (N_4510,N_4144,N_3839);
nand U4511 (N_4511,N_4432,N_4375);
nor U4512 (N_4512,N_3948,N_3967);
nand U4513 (N_4513,N_4341,N_4050);
and U4514 (N_4514,N_4446,N_3817);
xor U4515 (N_4515,N_4015,N_4241);
xnor U4516 (N_4516,N_4450,N_3784);
nand U4517 (N_4517,N_4102,N_3988);
nor U4518 (N_4518,N_4104,N_4374);
nor U4519 (N_4519,N_3961,N_3888);
nor U4520 (N_4520,N_4113,N_4009);
nand U4521 (N_4521,N_3771,N_4087);
nand U4522 (N_4522,N_3912,N_3968);
xor U4523 (N_4523,N_4407,N_3797);
and U4524 (N_4524,N_4333,N_3918);
xor U4525 (N_4525,N_3759,N_4314);
nand U4526 (N_4526,N_4386,N_4209);
xnor U4527 (N_4527,N_4026,N_3872);
nor U4528 (N_4528,N_4169,N_3944);
xnor U4529 (N_4529,N_3881,N_4279);
nand U4530 (N_4530,N_4021,N_4331);
and U4531 (N_4531,N_4383,N_3959);
nor U4532 (N_4532,N_4205,N_4349);
or U4533 (N_4533,N_4246,N_4173);
xnor U4534 (N_4534,N_3882,N_4251);
nor U4535 (N_4535,N_3853,N_4302);
nor U4536 (N_4536,N_4280,N_3828);
nand U4537 (N_4537,N_4444,N_4031);
and U4538 (N_4538,N_4300,N_3800);
nor U4539 (N_4539,N_4426,N_4237);
or U4540 (N_4540,N_4422,N_4166);
nor U4541 (N_4541,N_4382,N_4325);
or U4542 (N_4542,N_4137,N_3983);
or U4543 (N_4543,N_3805,N_4025);
or U4544 (N_4544,N_4215,N_4041);
xnor U4545 (N_4545,N_3952,N_4451);
nor U4546 (N_4546,N_4298,N_4044);
or U4547 (N_4547,N_3902,N_4410);
xor U4548 (N_4548,N_4262,N_4002);
xor U4549 (N_4549,N_4423,N_4250);
nor U4550 (N_4550,N_3788,N_3995);
and U4551 (N_4551,N_4351,N_3806);
nand U4552 (N_4552,N_4082,N_4274);
nand U4553 (N_4553,N_3929,N_4106);
nor U4554 (N_4554,N_3826,N_4212);
nand U4555 (N_4555,N_3907,N_4380);
xor U4556 (N_4556,N_3916,N_4295);
xnor U4557 (N_4557,N_3884,N_4018);
nand U4558 (N_4558,N_3767,N_3849);
or U4559 (N_4559,N_3991,N_4271);
and U4560 (N_4560,N_4471,N_3877);
xnor U4561 (N_4561,N_4245,N_4318);
xor U4562 (N_4562,N_4477,N_4406);
nand U4563 (N_4563,N_4086,N_4072);
nand U4564 (N_4564,N_4148,N_4017);
and U4565 (N_4565,N_3871,N_4083);
nor U4566 (N_4566,N_4223,N_4490);
or U4567 (N_4567,N_3766,N_3984);
and U4568 (N_4568,N_4301,N_4191);
and U4569 (N_4569,N_4466,N_3942);
xnor U4570 (N_4570,N_4475,N_4437);
nand U4571 (N_4571,N_3950,N_4195);
and U4572 (N_4572,N_4235,N_3910);
nand U4573 (N_4573,N_3772,N_4448);
nor U4574 (N_4574,N_4114,N_3892);
nand U4575 (N_4575,N_4365,N_4270);
xor U4576 (N_4576,N_4493,N_4238);
and U4577 (N_4577,N_4421,N_4231);
xnor U4578 (N_4578,N_3996,N_4040);
nor U4579 (N_4579,N_4225,N_4263);
xnor U4580 (N_4580,N_3835,N_3799);
and U4581 (N_4581,N_3949,N_3923);
nor U4582 (N_4582,N_4109,N_3964);
nand U4583 (N_4583,N_4308,N_4327);
nor U4584 (N_4584,N_3879,N_4389);
xor U4585 (N_4585,N_4284,N_4335);
nand U4586 (N_4586,N_4126,N_3941);
xnor U4587 (N_4587,N_4277,N_4127);
nor U4588 (N_4588,N_4162,N_4188);
and U4589 (N_4589,N_4478,N_3896);
nor U4590 (N_4590,N_4061,N_4005);
or U4591 (N_4591,N_4037,N_3926);
nand U4592 (N_4592,N_4004,N_4348);
and U4593 (N_4593,N_4293,N_4056);
xnor U4594 (N_4594,N_3753,N_3885);
xor U4595 (N_4595,N_4412,N_4036);
nand U4596 (N_4596,N_4180,N_3764);
and U4597 (N_4597,N_3955,N_4417);
nand U4598 (N_4598,N_4499,N_4123);
nor U4599 (N_4599,N_4142,N_4115);
and U4600 (N_4600,N_4467,N_3813);
nor U4601 (N_4601,N_3765,N_4133);
and U4602 (N_4602,N_4100,N_3779);
or U4603 (N_4603,N_4474,N_4024);
xor U4604 (N_4604,N_4035,N_4399);
or U4605 (N_4605,N_4481,N_4268);
or U4606 (N_4606,N_4084,N_4160);
nor U4607 (N_4607,N_4273,N_3867);
nor U4608 (N_4608,N_4385,N_4292);
xor U4609 (N_4609,N_4310,N_4248);
and U4610 (N_4610,N_4364,N_3865);
nor U4611 (N_4611,N_3760,N_4343);
xor U4612 (N_4612,N_4470,N_4128);
and U4613 (N_4613,N_4071,N_3762);
nor U4614 (N_4614,N_4119,N_4355);
nor U4615 (N_4615,N_3852,N_4187);
nor U4616 (N_4616,N_4449,N_3795);
or U4617 (N_4617,N_3818,N_4424);
xnor U4618 (N_4618,N_3785,N_4189);
xnor U4619 (N_4619,N_4456,N_4255);
or U4620 (N_4620,N_4034,N_4342);
xnor U4621 (N_4621,N_4309,N_4081);
xor U4622 (N_4622,N_4054,N_3850);
or U4623 (N_4623,N_3900,N_4013);
xnor U4624 (N_4624,N_4161,N_3861);
or U4625 (N_4625,N_4266,N_4053);
or U4626 (N_4626,N_4055,N_4244);
nor U4627 (N_4627,N_4023,N_4210);
nand U4628 (N_4628,N_4392,N_4324);
nor U4629 (N_4629,N_3989,N_4108);
nand U4630 (N_4630,N_4306,N_4122);
and U4631 (N_4631,N_4125,N_3838);
and U4632 (N_4632,N_4088,N_3855);
nor U4633 (N_4633,N_4289,N_3908);
and U4634 (N_4634,N_3897,N_3927);
or U4635 (N_4635,N_4062,N_4218);
nor U4636 (N_4636,N_3775,N_4488);
nand U4637 (N_4637,N_4413,N_4479);
and U4638 (N_4638,N_4131,N_4157);
and U4639 (N_4639,N_3858,N_4214);
and U4640 (N_4640,N_4216,N_4294);
nand U4641 (N_4641,N_4336,N_4369);
or U4642 (N_4642,N_4076,N_3943);
xnor U4643 (N_4643,N_3936,N_4149);
and U4644 (N_4644,N_3893,N_3756);
and U4645 (N_4645,N_4495,N_4043);
nor U4646 (N_4646,N_4158,N_3901);
xor U4647 (N_4647,N_4316,N_4226);
nor U4648 (N_4648,N_4435,N_3829);
nor U4649 (N_4649,N_4130,N_4264);
and U4650 (N_4650,N_4443,N_4174);
nor U4651 (N_4651,N_3919,N_4372);
or U4652 (N_4652,N_4080,N_4267);
or U4653 (N_4653,N_4038,N_3928);
and U4654 (N_4654,N_4000,N_3997);
nand U4655 (N_4655,N_4473,N_4090);
xor U4656 (N_4656,N_4261,N_4346);
nor U4657 (N_4657,N_4199,N_4496);
nand U4658 (N_4658,N_4103,N_3862);
nand U4659 (N_4659,N_4096,N_3904);
nor U4660 (N_4660,N_4402,N_3794);
nor U4661 (N_4661,N_4299,N_3887);
nor U4662 (N_4662,N_4350,N_3899);
nand U4663 (N_4663,N_4340,N_3985);
and U4664 (N_4664,N_4420,N_3823);
and U4665 (N_4665,N_3906,N_4155);
nor U4666 (N_4666,N_4112,N_4176);
nor U4667 (N_4667,N_3930,N_4156);
nand U4668 (N_4668,N_4332,N_4095);
xor U4669 (N_4669,N_4051,N_3980);
and U4670 (N_4670,N_4282,N_3778);
nand U4671 (N_4671,N_4430,N_4398);
nand U4672 (N_4672,N_4193,N_4457);
nand U4673 (N_4673,N_4391,N_3898);
and U4674 (N_4674,N_4281,N_3847);
or U4675 (N_4675,N_3819,N_3856);
nor U4676 (N_4676,N_4440,N_3994);
nand U4677 (N_4677,N_4434,N_4097);
nand U4678 (N_4678,N_4204,N_3947);
nor U4679 (N_4679,N_4252,N_4227);
and U4680 (N_4680,N_4178,N_4287);
and U4681 (N_4681,N_3951,N_3832);
nor U4682 (N_4682,N_4357,N_4164);
or U4683 (N_4683,N_4269,N_4186);
nand U4684 (N_4684,N_4371,N_4482);
or U4685 (N_4685,N_3781,N_4151);
xor U4686 (N_4686,N_4453,N_4283);
nand U4687 (N_4687,N_3874,N_4116);
xor U4688 (N_4688,N_4359,N_4243);
nor U4689 (N_4689,N_3969,N_4322);
nor U4690 (N_4690,N_4405,N_3807);
xor U4691 (N_4691,N_3840,N_4361);
and U4692 (N_4692,N_3973,N_4256);
and U4693 (N_4693,N_4428,N_3821);
or U4694 (N_4694,N_4120,N_3956);
or U4695 (N_4695,N_3934,N_4312);
xor U4696 (N_4696,N_4376,N_4208);
or U4697 (N_4697,N_4338,N_3820);
and U4698 (N_4698,N_4360,N_4464);
nand U4699 (N_4699,N_4020,N_4344);
and U4700 (N_4700,N_4192,N_3808);
and U4701 (N_4701,N_4290,N_4254);
nand U4702 (N_4702,N_4319,N_3812);
nor U4703 (N_4703,N_4033,N_4249);
nand U4704 (N_4704,N_3895,N_4439);
xnor U4705 (N_4705,N_4064,N_4303);
nor U4706 (N_4706,N_4006,N_4498);
or U4707 (N_4707,N_3777,N_3886);
xor U4708 (N_4708,N_4487,N_4429);
nor U4709 (N_4709,N_3890,N_3790);
or U4710 (N_4710,N_4171,N_3889);
and U4711 (N_4711,N_4370,N_4001);
nand U4712 (N_4712,N_4105,N_3815);
and U4713 (N_4713,N_4404,N_4489);
nand U4714 (N_4714,N_3843,N_4206);
and U4715 (N_4715,N_4200,N_3851);
nor U4716 (N_4716,N_4184,N_3791);
or U4717 (N_4717,N_4030,N_3873);
nand U4718 (N_4718,N_4165,N_4461);
or U4719 (N_4719,N_4058,N_3845);
and U4720 (N_4720,N_3945,N_4468);
nand U4721 (N_4721,N_3814,N_4181);
or U4722 (N_4722,N_4177,N_4027);
or U4723 (N_4723,N_4132,N_4141);
or U4724 (N_4724,N_4194,N_4311);
nand U4725 (N_4725,N_4010,N_3848);
and U4726 (N_4726,N_4296,N_4313);
or U4727 (N_4727,N_4012,N_4046);
nor U4728 (N_4728,N_4217,N_4363);
xnor U4729 (N_4729,N_4150,N_3922);
nand U4730 (N_4730,N_4433,N_4465);
or U4731 (N_4731,N_3811,N_4134);
nor U4732 (N_4732,N_4275,N_4197);
nand U4733 (N_4733,N_3958,N_3987);
and U4734 (N_4734,N_4345,N_4168);
and U4735 (N_4735,N_4063,N_3965);
nand U4736 (N_4736,N_3963,N_4257);
nand U4737 (N_4737,N_3859,N_4354);
nor U4738 (N_4738,N_3998,N_3982);
or U4739 (N_4739,N_4032,N_4317);
or U4740 (N_4740,N_3891,N_3915);
or U4741 (N_4741,N_3875,N_3774);
nor U4742 (N_4742,N_4211,N_3905);
or U4743 (N_4743,N_4098,N_4373);
nor U4744 (N_4744,N_4390,N_3866);
or U4745 (N_4745,N_3776,N_3940);
nand U4746 (N_4746,N_4101,N_4339);
nand U4747 (N_4747,N_4207,N_4147);
and U4748 (N_4748,N_4185,N_4220);
nand U4749 (N_4749,N_4427,N_3837);
and U4750 (N_4750,N_4403,N_3757);
xor U4751 (N_4751,N_4259,N_4042);
and U4752 (N_4752,N_4078,N_4352);
xor U4753 (N_4753,N_3793,N_4089);
or U4754 (N_4754,N_3830,N_4441);
nor U4755 (N_4755,N_3880,N_3864);
nor U4756 (N_4756,N_4140,N_3782);
xnor U4757 (N_4757,N_3894,N_4458);
or U4758 (N_4758,N_3978,N_3768);
nor U4759 (N_4759,N_4276,N_3751);
or U4760 (N_4760,N_4016,N_3786);
or U4761 (N_4761,N_4085,N_3878);
nor U4762 (N_4762,N_4396,N_4222);
or U4763 (N_4763,N_3761,N_4240);
xor U4764 (N_4764,N_4362,N_3979);
xor U4765 (N_4765,N_4224,N_4272);
nor U4766 (N_4766,N_4045,N_4230);
xor U4767 (N_4767,N_4260,N_3954);
and U4768 (N_4768,N_4418,N_4154);
xnor U4769 (N_4769,N_4146,N_4400);
nand U4770 (N_4770,N_4179,N_3809);
xor U4771 (N_4771,N_4070,N_4228);
nand U4772 (N_4772,N_4288,N_4234);
nor U4773 (N_4773,N_3883,N_4347);
xnor U4774 (N_4774,N_3925,N_3846);
nor U4775 (N_4775,N_3986,N_4019);
nor U4776 (N_4776,N_3909,N_4124);
and U4777 (N_4777,N_4048,N_4039);
nor U4778 (N_4778,N_4384,N_3802);
nand U4779 (N_4779,N_4029,N_3870);
nor U4780 (N_4780,N_3977,N_3931);
xnor U4781 (N_4781,N_3816,N_4167);
or U4782 (N_4782,N_4074,N_4483);
and U4783 (N_4783,N_4455,N_4196);
nand U4784 (N_4784,N_3863,N_4379);
nand U4785 (N_4785,N_4258,N_4286);
and U4786 (N_4786,N_4408,N_4321);
nand U4787 (N_4787,N_4454,N_3924);
and U4788 (N_4788,N_4183,N_4469);
or U4789 (N_4789,N_4069,N_4476);
and U4790 (N_4790,N_4462,N_3914);
nor U4791 (N_4791,N_4011,N_4057);
and U4792 (N_4792,N_3917,N_3758);
nand U4793 (N_4793,N_3920,N_3957);
xnor U4794 (N_4794,N_3921,N_4229);
xnor U4795 (N_4795,N_3953,N_3966);
nor U4796 (N_4796,N_4121,N_3824);
xnor U4797 (N_4797,N_3796,N_3976);
and U4798 (N_4798,N_3962,N_4066);
xor U4799 (N_4799,N_4182,N_3810);
or U4800 (N_4800,N_4202,N_4239);
or U4801 (N_4801,N_3844,N_4497);
xnor U4802 (N_4802,N_3937,N_4409);
nand U4803 (N_4803,N_3773,N_3833);
xor U4804 (N_4804,N_4366,N_4425);
and U4805 (N_4805,N_4092,N_3783);
and U4806 (N_4806,N_4059,N_4247);
nand U4807 (N_4807,N_4484,N_3932);
or U4808 (N_4808,N_4485,N_3789);
or U4809 (N_4809,N_4265,N_4091);
nand U4810 (N_4810,N_4135,N_3939);
xnor U4811 (N_4811,N_4393,N_4387);
and U4812 (N_4812,N_4221,N_4337);
nor U4813 (N_4813,N_4028,N_4459);
or U4814 (N_4814,N_4094,N_4073);
xor U4815 (N_4815,N_3755,N_4494);
or U4816 (N_4816,N_4198,N_3993);
and U4817 (N_4817,N_4172,N_4065);
or U4818 (N_4818,N_4472,N_3750);
nor U4819 (N_4819,N_4145,N_4414);
nand U4820 (N_4820,N_4099,N_4323);
xnor U4821 (N_4821,N_3933,N_4397);
or U4822 (N_4822,N_4190,N_3825);
nor U4823 (N_4823,N_4008,N_4368);
and U4824 (N_4824,N_4136,N_4329);
nand U4825 (N_4825,N_3787,N_4291);
and U4826 (N_4826,N_4480,N_4242);
nor U4827 (N_4827,N_4401,N_4152);
nor U4828 (N_4828,N_4077,N_4491);
or U4829 (N_4829,N_4107,N_4236);
or U4830 (N_4830,N_4110,N_4353);
nand U4831 (N_4831,N_4326,N_4320);
nand U4832 (N_4832,N_3970,N_4419);
or U4833 (N_4833,N_3876,N_3822);
or U4834 (N_4834,N_4415,N_4139);
or U4835 (N_4835,N_4394,N_3946);
and U4836 (N_4836,N_4304,N_4388);
or U4837 (N_4837,N_3752,N_4307);
and U4838 (N_4838,N_3975,N_4143);
xor U4839 (N_4839,N_4438,N_4093);
and U4840 (N_4840,N_4378,N_4297);
xor U4841 (N_4841,N_3857,N_3841);
nand U4842 (N_4842,N_4175,N_3770);
or U4843 (N_4843,N_3903,N_3831);
and U4844 (N_4844,N_3981,N_3763);
and U4845 (N_4845,N_3911,N_4022);
and U4846 (N_4846,N_3804,N_4411);
xor U4847 (N_4847,N_4436,N_3972);
or U4848 (N_4848,N_3938,N_4007);
nor U4849 (N_4849,N_4233,N_4201);
and U4850 (N_4850,N_3798,N_4068);
nor U4851 (N_4851,N_4219,N_3974);
xor U4852 (N_4852,N_4159,N_4328);
nand U4853 (N_4853,N_4486,N_3999);
and U4854 (N_4854,N_4358,N_4047);
nand U4855 (N_4855,N_4452,N_4356);
nand U4856 (N_4856,N_3992,N_4315);
nor U4857 (N_4857,N_4111,N_4049);
or U4858 (N_4858,N_4163,N_3990);
and U4859 (N_4859,N_4075,N_4395);
nand U4860 (N_4860,N_4203,N_4117);
nor U4861 (N_4861,N_4330,N_4129);
or U4862 (N_4862,N_3854,N_4460);
nand U4863 (N_4863,N_4213,N_4153);
or U4864 (N_4864,N_4138,N_4285);
nand U4865 (N_4865,N_4431,N_4305);
and U4866 (N_4866,N_4253,N_3827);
and U4867 (N_4867,N_3754,N_4067);
nand U4868 (N_4868,N_4079,N_4416);
nor U4869 (N_4869,N_4381,N_3960);
or U4870 (N_4870,N_3913,N_4334);
nor U4871 (N_4871,N_4445,N_3935);
nand U4872 (N_4872,N_3803,N_3842);
nor U4873 (N_4873,N_4442,N_3860);
xor U4874 (N_4874,N_4367,N_4463);
nor U4875 (N_4875,N_3763,N_4246);
xor U4876 (N_4876,N_3884,N_4010);
nor U4877 (N_4877,N_3842,N_3983);
nand U4878 (N_4878,N_4376,N_3855);
and U4879 (N_4879,N_3921,N_4483);
nand U4880 (N_4880,N_4081,N_4315);
xnor U4881 (N_4881,N_3940,N_4105);
nor U4882 (N_4882,N_3965,N_3830);
xnor U4883 (N_4883,N_4055,N_4204);
xor U4884 (N_4884,N_4364,N_4272);
nor U4885 (N_4885,N_3826,N_4097);
and U4886 (N_4886,N_4356,N_4322);
or U4887 (N_4887,N_4488,N_4143);
or U4888 (N_4888,N_4205,N_4379);
xor U4889 (N_4889,N_4423,N_3761);
or U4890 (N_4890,N_4205,N_3766);
nor U4891 (N_4891,N_4361,N_4481);
xor U4892 (N_4892,N_4053,N_4103);
nand U4893 (N_4893,N_4317,N_4294);
xnor U4894 (N_4894,N_3750,N_4347);
xor U4895 (N_4895,N_4449,N_4417);
and U4896 (N_4896,N_4225,N_3762);
or U4897 (N_4897,N_3886,N_3975);
and U4898 (N_4898,N_4385,N_4048);
xnor U4899 (N_4899,N_3868,N_3843);
nand U4900 (N_4900,N_4140,N_3912);
nor U4901 (N_4901,N_3759,N_3949);
or U4902 (N_4902,N_4190,N_4293);
and U4903 (N_4903,N_4484,N_4197);
nor U4904 (N_4904,N_4012,N_3864);
nor U4905 (N_4905,N_4197,N_4177);
nand U4906 (N_4906,N_3856,N_4448);
and U4907 (N_4907,N_3906,N_3984);
and U4908 (N_4908,N_4213,N_3824);
nor U4909 (N_4909,N_4050,N_4300);
nand U4910 (N_4910,N_4116,N_4300);
and U4911 (N_4911,N_4188,N_3886);
nand U4912 (N_4912,N_4144,N_4471);
nand U4913 (N_4913,N_4138,N_4377);
nor U4914 (N_4914,N_4335,N_3803);
and U4915 (N_4915,N_3760,N_4007);
or U4916 (N_4916,N_4180,N_4433);
nand U4917 (N_4917,N_4233,N_3828);
and U4918 (N_4918,N_4415,N_4037);
xor U4919 (N_4919,N_4364,N_4396);
nand U4920 (N_4920,N_4439,N_3813);
nor U4921 (N_4921,N_4013,N_4069);
nand U4922 (N_4922,N_4263,N_4373);
nand U4923 (N_4923,N_4283,N_3756);
or U4924 (N_4924,N_4100,N_4212);
nand U4925 (N_4925,N_3814,N_3786);
and U4926 (N_4926,N_4126,N_3867);
nand U4927 (N_4927,N_3934,N_3943);
or U4928 (N_4928,N_4260,N_3753);
xnor U4929 (N_4929,N_4205,N_4108);
or U4930 (N_4930,N_4367,N_3814);
nand U4931 (N_4931,N_3812,N_4341);
or U4932 (N_4932,N_4408,N_4380);
and U4933 (N_4933,N_4487,N_4454);
or U4934 (N_4934,N_4412,N_4346);
xnor U4935 (N_4935,N_4127,N_4034);
nor U4936 (N_4936,N_4491,N_4120);
nor U4937 (N_4937,N_4215,N_4376);
nand U4938 (N_4938,N_3985,N_4393);
or U4939 (N_4939,N_3965,N_4050);
or U4940 (N_4940,N_3905,N_3762);
nor U4941 (N_4941,N_4349,N_3856);
nor U4942 (N_4942,N_4228,N_4415);
xor U4943 (N_4943,N_4027,N_4046);
nor U4944 (N_4944,N_3822,N_3777);
and U4945 (N_4945,N_3820,N_4425);
xnor U4946 (N_4946,N_3792,N_4144);
nand U4947 (N_4947,N_3856,N_4441);
xor U4948 (N_4948,N_4392,N_4234);
nand U4949 (N_4949,N_4211,N_4353);
and U4950 (N_4950,N_4042,N_4469);
xor U4951 (N_4951,N_4297,N_4488);
or U4952 (N_4952,N_4437,N_3880);
nand U4953 (N_4953,N_3902,N_4104);
and U4954 (N_4954,N_3992,N_4220);
nor U4955 (N_4955,N_3961,N_4230);
nand U4956 (N_4956,N_4477,N_4154);
xnor U4957 (N_4957,N_4363,N_4438);
or U4958 (N_4958,N_4014,N_4215);
or U4959 (N_4959,N_4079,N_4319);
xnor U4960 (N_4960,N_3971,N_4402);
nand U4961 (N_4961,N_4271,N_3935);
or U4962 (N_4962,N_4027,N_4479);
or U4963 (N_4963,N_4020,N_4084);
nor U4964 (N_4964,N_4496,N_4075);
nor U4965 (N_4965,N_3869,N_4475);
nand U4966 (N_4966,N_3826,N_4298);
and U4967 (N_4967,N_4453,N_4162);
nor U4968 (N_4968,N_3788,N_4271);
xnor U4969 (N_4969,N_3954,N_4346);
or U4970 (N_4970,N_4435,N_3940);
and U4971 (N_4971,N_4091,N_4369);
or U4972 (N_4972,N_3792,N_4254);
xor U4973 (N_4973,N_4398,N_3996);
nor U4974 (N_4974,N_3756,N_4127);
and U4975 (N_4975,N_4413,N_3969);
nor U4976 (N_4976,N_4435,N_4222);
nor U4977 (N_4977,N_3959,N_4185);
or U4978 (N_4978,N_3906,N_3864);
nand U4979 (N_4979,N_3842,N_4475);
or U4980 (N_4980,N_3822,N_4229);
xnor U4981 (N_4981,N_4226,N_3947);
xnor U4982 (N_4982,N_3890,N_4421);
or U4983 (N_4983,N_4381,N_4361);
nor U4984 (N_4984,N_4496,N_3828);
and U4985 (N_4985,N_4234,N_4199);
xnor U4986 (N_4986,N_4175,N_4154);
nor U4987 (N_4987,N_4065,N_4223);
or U4988 (N_4988,N_3983,N_4149);
nand U4989 (N_4989,N_3812,N_4383);
nor U4990 (N_4990,N_3912,N_4039);
xor U4991 (N_4991,N_3974,N_4195);
and U4992 (N_4992,N_4326,N_4184);
or U4993 (N_4993,N_3924,N_4492);
and U4994 (N_4994,N_4054,N_3805);
xnor U4995 (N_4995,N_4131,N_4321);
nand U4996 (N_4996,N_4464,N_3817);
nor U4997 (N_4997,N_3793,N_3886);
nand U4998 (N_4998,N_4466,N_4456);
xor U4999 (N_4999,N_4401,N_4112);
xnor U5000 (N_5000,N_4021,N_3791);
xnor U5001 (N_5001,N_4050,N_4279);
nor U5002 (N_5002,N_3979,N_4073);
nand U5003 (N_5003,N_3878,N_3753);
and U5004 (N_5004,N_4126,N_4258);
nand U5005 (N_5005,N_4063,N_4097);
and U5006 (N_5006,N_4182,N_4054);
xnor U5007 (N_5007,N_4004,N_3806);
nand U5008 (N_5008,N_4189,N_3793);
nand U5009 (N_5009,N_4123,N_4097);
and U5010 (N_5010,N_4225,N_4097);
or U5011 (N_5011,N_4190,N_4350);
and U5012 (N_5012,N_3984,N_4439);
xor U5013 (N_5013,N_4148,N_3834);
nor U5014 (N_5014,N_3792,N_4171);
or U5015 (N_5015,N_3861,N_4478);
or U5016 (N_5016,N_4403,N_4203);
or U5017 (N_5017,N_4370,N_3794);
nand U5018 (N_5018,N_4203,N_3965);
nor U5019 (N_5019,N_4001,N_3901);
nor U5020 (N_5020,N_3753,N_3804);
nand U5021 (N_5021,N_4164,N_4264);
nand U5022 (N_5022,N_4484,N_4087);
nor U5023 (N_5023,N_3820,N_3912);
and U5024 (N_5024,N_4403,N_4217);
xor U5025 (N_5025,N_4091,N_4242);
nand U5026 (N_5026,N_4019,N_4426);
nand U5027 (N_5027,N_3948,N_4433);
xnor U5028 (N_5028,N_3772,N_4202);
nor U5029 (N_5029,N_4128,N_4421);
or U5030 (N_5030,N_3870,N_3909);
nand U5031 (N_5031,N_3875,N_4340);
and U5032 (N_5032,N_3823,N_4147);
and U5033 (N_5033,N_4325,N_3833);
or U5034 (N_5034,N_4201,N_4194);
nor U5035 (N_5035,N_3802,N_4149);
nor U5036 (N_5036,N_3990,N_4217);
or U5037 (N_5037,N_4251,N_3877);
and U5038 (N_5038,N_4358,N_4396);
and U5039 (N_5039,N_4470,N_4212);
and U5040 (N_5040,N_4187,N_4351);
and U5041 (N_5041,N_4388,N_4478);
nor U5042 (N_5042,N_4491,N_4261);
and U5043 (N_5043,N_4240,N_4256);
xnor U5044 (N_5044,N_4310,N_4176);
nor U5045 (N_5045,N_3835,N_4394);
or U5046 (N_5046,N_4406,N_4280);
nand U5047 (N_5047,N_4333,N_4356);
and U5048 (N_5048,N_3810,N_4166);
nor U5049 (N_5049,N_4256,N_3877);
nand U5050 (N_5050,N_4023,N_3786);
nand U5051 (N_5051,N_4435,N_4475);
nor U5052 (N_5052,N_4351,N_4169);
xor U5053 (N_5053,N_4312,N_3977);
and U5054 (N_5054,N_4026,N_4231);
xnor U5055 (N_5055,N_3979,N_3823);
nor U5056 (N_5056,N_3842,N_4027);
and U5057 (N_5057,N_4332,N_3971);
xor U5058 (N_5058,N_4041,N_3938);
or U5059 (N_5059,N_4043,N_4245);
or U5060 (N_5060,N_3793,N_4455);
nor U5061 (N_5061,N_3909,N_4419);
or U5062 (N_5062,N_4223,N_3814);
and U5063 (N_5063,N_4401,N_4294);
and U5064 (N_5064,N_3850,N_4123);
or U5065 (N_5065,N_3983,N_4213);
and U5066 (N_5066,N_4077,N_3834);
or U5067 (N_5067,N_3755,N_4204);
nor U5068 (N_5068,N_4120,N_3934);
and U5069 (N_5069,N_4076,N_3808);
xor U5070 (N_5070,N_4297,N_4386);
and U5071 (N_5071,N_4135,N_3901);
and U5072 (N_5072,N_3983,N_4156);
or U5073 (N_5073,N_4353,N_3902);
nor U5074 (N_5074,N_4241,N_3871);
and U5075 (N_5075,N_4015,N_4113);
xor U5076 (N_5076,N_4228,N_4141);
and U5077 (N_5077,N_3930,N_4185);
nand U5078 (N_5078,N_3912,N_4380);
and U5079 (N_5079,N_4132,N_4101);
xor U5080 (N_5080,N_4155,N_4241);
xnor U5081 (N_5081,N_4135,N_3821);
or U5082 (N_5082,N_3970,N_4238);
nor U5083 (N_5083,N_4070,N_4221);
xor U5084 (N_5084,N_4219,N_4469);
nor U5085 (N_5085,N_4369,N_4290);
nor U5086 (N_5086,N_4170,N_4415);
nand U5087 (N_5087,N_4066,N_4301);
nor U5088 (N_5088,N_4072,N_3870);
or U5089 (N_5089,N_4200,N_4479);
xor U5090 (N_5090,N_4328,N_4442);
nand U5091 (N_5091,N_4391,N_4044);
nand U5092 (N_5092,N_4030,N_4032);
xnor U5093 (N_5093,N_4063,N_4000);
or U5094 (N_5094,N_3928,N_4047);
xor U5095 (N_5095,N_4296,N_4377);
xnor U5096 (N_5096,N_4374,N_3875);
nand U5097 (N_5097,N_4481,N_4344);
and U5098 (N_5098,N_4222,N_4218);
xor U5099 (N_5099,N_4392,N_4075);
or U5100 (N_5100,N_4174,N_4376);
or U5101 (N_5101,N_4275,N_4051);
xnor U5102 (N_5102,N_3825,N_4192);
nor U5103 (N_5103,N_4330,N_4148);
nand U5104 (N_5104,N_4196,N_4189);
nor U5105 (N_5105,N_3893,N_4382);
xnor U5106 (N_5106,N_3990,N_3915);
and U5107 (N_5107,N_3886,N_4014);
and U5108 (N_5108,N_4021,N_4046);
nand U5109 (N_5109,N_4480,N_3914);
nand U5110 (N_5110,N_4395,N_3768);
nor U5111 (N_5111,N_4205,N_4453);
xor U5112 (N_5112,N_4264,N_4402);
nand U5113 (N_5113,N_4302,N_4109);
xnor U5114 (N_5114,N_4351,N_4348);
nand U5115 (N_5115,N_3849,N_4273);
nand U5116 (N_5116,N_3952,N_4101);
nor U5117 (N_5117,N_4082,N_4282);
nor U5118 (N_5118,N_4386,N_3902);
or U5119 (N_5119,N_4227,N_4024);
xnor U5120 (N_5120,N_4295,N_4291);
nand U5121 (N_5121,N_4445,N_3823);
nand U5122 (N_5122,N_4442,N_3858);
xor U5123 (N_5123,N_3958,N_4263);
nor U5124 (N_5124,N_4351,N_3826);
xnor U5125 (N_5125,N_4160,N_4054);
nor U5126 (N_5126,N_4196,N_4146);
or U5127 (N_5127,N_4266,N_4395);
xor U5128 (N_5128,N_4239,N_4429);
and U5129 (N_5129,N_3829,N_4450);
xnor U5130 (N_5130,N_4145,N_4268);
xor U5131 (N_5131,N_4321,N_4120);
nor U5132 (N_5132,N_4071,N_3835);
xor U5133 (N_5133,N_4286,N_4232);
xnor U5134 (N_5134,N_4308,N_4183);
or U5135 (N_5135,N_4496,N_3834);
nor U5136 (N_5136,N_3885,N_4333);
nor U5137 (N_5137,N_3871,N_3961);
or U5138 (N_5138,N_4183,N_4237);
nor U5139 (N_5139,N_4014,N_4004);
nor U5140 (N_5140,N_4251,N_4303);
or U5141 (N_5141,N_4424,N_4333);
or U5142 (N_5142,N_4449,N_4332);
and U5143 (N_5143,N_3805,N_3937);
and U5144 (N_5144,N_3972,N_4294);
nand U5145 (N_5145,N_4253,N_4206);
and U5146 (N_5146,N_4064,N_3827);
nor U5147 (N_5147,N_4128,N_3875);
nand U5148 (N_5148,N_4329,N_4482);
and U5149 (N_5149,N_4029,N_4109);
or U5150 (N_5150,N_4458,N_4074);
and U5151 (N_5151,N_4463,N_4279);
nand U5152 (N_5152,N_4377,N_4331);
or U5153 (N_5153,N_3925,N_3943);
nand U5154 (N_5154,N_4144,N_3935);
nor U5155 (N_5155,N_4041,N_3953);
xor U5156 (N_5156,N_4119,N_4211);
nand U5157 (N_5157,N_4211,N_4341);
xnor U5158 (N_5158,N_4435,N_4144);
xor U5159 (N_5159,N_4154,N_4321);
and U5160 (N_5160,N_3859,N_4264);
and U5161 (N_5161,N_4191,N_3986);
nor U5162 (N_5162,N_3812,N_3750);
nand U5163 (N_5163,N_4101,N_4300);
nor U5164 (N_5164,N_4418,N_4466);
nand U5165 (N_5165,N_3983,N_3816);
xor U5166 (N_5166,N_4060,N_3773);
xor U5167 (N_5167,N_4397,N_4174);
or U5168 (N_5168,N_4034,N_4368);
xor U5169 (N_5169,N_3963,N_4244);
xor U5170 (N_5170,N_4300,N_3756);
xnor U5171 (N_5171,N_4193,N_4028);
or U5172 (N_5172,N_4001,N_4404);
nand U5173 (N_5173,N_3831,N_3775);
nand U5174 (N_5174,N_4374,N_4458);
or U5175 (N_5175,N_3800,N_3904);
nor U5176 (N_5176,N_4131,N_4293);
or U5177 (N_5177,N_4161,N_3883);
and U5178 (N_5178,N_4190,N_3937);
and U5179 (N_5179,N_3851,N_3756);
xor U5180 (N_5180,N_4092,N_4483);
and U5181 (N_5181,N_4140,N_4227);
nand U5182 (N_5182,N_3889,N_4202);
or U5183 (N_5183,N_4230,N_4170);
nor U5184 (N_5184,N_3772,N_4294);
nor U5185 (N_5185,N_4034,N_3993);
nand U5186 (N_5186,N_4212,N_4057);
nand U5187 (N_5187,N_4410,N_4088);
nor U5188 (N_5188,N_4024,N_3918);
xnor U5189 (N_5189,N_3864,N_3937);
nand U5190 (N_5190,N_3895,N_4345);
or U5191 (N_5191,N_3856,N_4419);
nor U5192 (N_5192,N_4378,N_3934);
nand U5193 (N_5193,N_3819,N_4419);
nor U5194 (N_5194,N_4280,N_4333);
and U5195 (N_5195,N_3808,N_3782);
nand U5196 (N_5196,N_4119,N_3995);
and U5197 (N_5197,N_4266,N_4179);
nor U5198 (N_5198,N_4175,N_4465);
nand U5199 (N_5199,N_3910,N_4205);
or U5200 (N_5200,N_3772,N_4098);
nand U5201 (N_5201,N_4410,N_3968);
nor U5202 (N_5202,N_4353,N_4443);
nand U5203 (N_5203,N_3906,N_4236);
nand U5204 (N_5204,N_4037,N_4252);
and U5205 (N_5205,N_4454,N_3837);
or U5206 (N_5206,N_4009,N_4116);
or U5207 (N_5207,N_3973,N_4414);
nand U5208 (N_5208,N_4240,N_4375);
nor U5209 (N_5209,N_4463,N_4100);
and U5210 (N_5210,N_4161,N_4159);
or U5211 (N_5211,N_4163,N_4248);
xnor U5212 (N_5212,N_4362,N_4298);
xor U5213 (N_5213,N_4437,N_4440);
and U5214 (N_5214,N_3756,N_3831);
or U5215 (N_5215,N_4396,N_3991);
and U5216 (N_5216,N_4230,N_4071);
or U5217 (N_5217,N_4140,N_3756);
nand U5218 (N_5218,N_3992,N_3912);
xnor U5219 (N_5219,N_3756,N_4396);
xor U5220 (N_5220,N_4234,N_4233);
nand U5221 (N_5221,N_4071,N_4459);
nand U5222 (N_5222,N_3911,N_4125);
xnor U5223 (N_5223,N_4408,N_4112);
xor U5224 (N_5224,N_4084,N_4159);
xor U5225 (N_5225,N_4143,N_4153);
and U5226 (N_5226,N_3834,N_4437);
and U5227 (N_5227,N_4211,N_3782);
xor U5228 (N_5228,N_4237,N_4294);
and U5229 (N_5229,N_3782,N_4463);
or U5230 (N_5230,N_4180,N_4080);
nand U5231 (N_5231,N_4440,N_4339);
or U5232 (N_5232,N_4100,N_3778);
or U5233 (N_5233,N_4477,N_4250);
and U5234 (N_5234,N_4444,N_3989);
xor U5235 (N_5235,N_4113,N_4106);
and U5236 (N_5236,N_4093,N_4494);
nor U5237 (N_5237,N_3916,N_4325);
nor U5238 (N_5238,N_3866,N_4472);
nand U5239 (N_5239,N_4376,N_3808);
or U5240 (N_5240,N_4449,N_3965);
nor U5241 (N_5241,N_4487,N_4025);
and U5242 (N_5242,N_4285,N_4301);
xnor U5243 (N_5243,N_4325,N_4170);
nor U5244 (N_5244,N_4083,N_4012);
nor U5245 (N_5245,N_3936,N_3755);
nor U5246 (N_5246,N_4333,N_4128);
or U5247 (N_5247,N_4191,N_4471);
nand U5248 (N_5248,N_4439,N_4044);
nand U5249 (N_5249,N_3963,N_3902);
xor U5250 (N_5250,N_4740,N_4605);
nor U5251 (N_5251,N_4987,N_4896);
nor U5252 (N_5252,N_4769,N_4720);
and U5253 (N_5253,N_4506,N_4622);
xnor U5254 (N_5254,N_4932,N_4802);
and U5255 (N_5255,N_4998,N_4598);
nand U5256 (N_5256,N_4995,N_4805);
nand U5257 (N_5257,N_4973,N_5008);
nand U5258 (N_5258,N_5144,N_5118);
xnor U5259 (N_5259,N_5157,N_5088);
xnor U5260 (N_5260,N_4825,N_4866);
nand U5261 (N_5261,N_4845,N_5188);
or U5262 (N_5262,N_5174,N_4939);
and U5263 (N_5263,N_4823,N_5029);
or U5264 (N_5264,N_4876,N_4560);
and U5265 (N_5265,N_4906,N_5190);
nand U5266 (N_5266,N_4821,N_4791);
and U5267 (N_5267,N_5241,N_4628);
or U5268 (N_5268,N_4510,N_4601);
or U5269 (N_5269,N_4798,N_4726);
nor U5270 (N_5270,N_4635,N_4661);
or U5271 (N_5271,N_5187,N_5135);
or U5272 (N_5272,N_4624,N_4859);
nand U5273 (N_5273,N_4977,N_4871);
nand U5274 (N_5274,N_4610,N_4915);
and U5275 (N_5275,N_4652,N_4651);
nor U5276 (N_5276,N_4558,N_5125);
nor U5277 (N_5277,N_4814,N_5159);
xnor U5278 (N_5278,N_4850,N_4674);
nor U5279 (N_5279,N_4929,N_5162);
xor U5280 (N_5280,N_4663,N_4618);
or U5281 (N_5281,N_4761,N_5134);
xnor U5282 (N_5282,N_4794,N_4765);
nor U5283 (N_5283,N_4826,N_4943);
nor U5284 (N_5284,N_4533,N_4971);
nor U5285 (N_5285,N_5163,N_4789);
or U5286 (N_5286,N_5039,N_4970);
nand U5287 (N_5287,N_5082,N_5120);
xor U5288 (N_5288,N_4518,N_5165);
xnor U5289 (N_5289,N_4569,N_5244);
xor U5290 (N_5290,N_4579,N_5231);
xnor U5291 (N_5291,N_4724,N_4656);
nor U5292 (N_5292,N_5110,N_5153);
or U5293 (N_5293,N_5168,N_4909);
or U5294 (N_5294,N_5073,N_5240);
nor U5295 (N_5295,N_4679,N_5161);
or U5296 (N_5296,N_5057,N_4888);
nor U5297 (N_5297,N_5107,N_4891);
and U5298 (N_5298,N_5204,N_5184);
nor U5299 (N_5299,N_5132,N_5051);
nor U5300 (N_5300,N_5084,N_5200);
nand U5301 (N_5301,N_4695,N_4937);
or U5302 (N_5302,N_5047,N_4535);
nand U5303 (N_5303,N_4701,N_4790);
nor U5304 (N_5304,N_4920,N_4702);
nand U5305 (N_5305,N_4594,N_4772);
and U5306 (N_5306,N_4684,N_5154);
and U5307 (N_5307,N_4952,N_4751);
and U5308 (N_5308,N_4875,N_4646);
xor U5309 (N_5309,N_5014,N_4557);
xor U5310 (N_5310,N_4846,N_5043);
or U5311 (N_5311,N_4827,N_5219);
or U5312 (N_5312,N_5197,N_4919);
nor U5313 (N_5313,N_4942,N_4536);
or U5314 (N_5314,N_4617,N_5237);
xor U5315 (N_5315,N_5139,N_5178);
nand U5316 (N_5316,N_4901,N_5095);
or U5317 (N_5317,N_4697,N_4596);
nor U5318 (N_5318,N_4978,N_5233);
or U5319 (N_5319,N_4689,N_4925);
nor U5320 (N_5320,N_4640,N_4815);
and U5321 (N_5321,N_5199,N_4922);
xor U5322 (N_5322,N_5045,N_5037);
xor U5323 (N_5323,N_5106,N_4949);
and U5324 (N_5324,N_4524,N_5248);
xor U5325 (N_5325,N_4575,N_4705);
and U5326 (N_5326,N_4833,N_4961);
nand U5327 (N_5327,N_4944,N_5031);
nand U5328 (N_5328,N_5097,N_5035);
and U5329 (N_5329,N_4706,N_4813);
nor U5330 (N_5330,N_4523,N_5228);
or U5331 (N_5331,N_5215,N_5185);
nand U5332 (N_5332,N_4849,N_4636);
xor U5333 (N_5333,N_5203,N_4722);
xnor U5334 (N_5334,N_5115,N_5175);
xnor U5335 (N_5335,N_5218,N_5116);
or U5336 (N_5336,N_5119,N_4566);
xnor U5337 (N_5337,N_4747,N_4621);
nand U5338 (N_5338,N_4865,N_5013);
and U5339 (N_5339,N_4568,N_5036);
xor U5340 (N_5340,N_5041,N_4658);
xor U5341 (N_5341,N_5083,N_4890);
nand U5342 (N_5342,N_5143,N_5022);
nor U5343 (N_5343,N_4779,N_4817);
nand U5344 (N_5344,N_4667,N_4629);
nor U5345 (N_5345,N_4894,N_4764);
xnor U5346 (N_5346,N_5109,N_5121);
or U5347 (N_5347,N_4728,N_4693);
xor U5348 (N_5348,N_5247,N_4811);
nand U5349 (N_5349,N_4550,N_4620);
and U5350 (N_5350,N_4732,N_5122);
nand U5351 (N_5351,N_4946,N_4976);
nor U5352 (N_5352,N_5076,N_4503);
or U5353 (N_5353,N_4967,N_5004);
nand U5354 (N_5354,N_5096,N_4545);
xor U5355 (N_5355,N_4650,N_4743);
xnor U5356 (N_5356,N_4522,N_4832);
and U5357 (N_5357,N_4672,N_4800);
xor U5358 (N_5358,N_5191,N_4861);
xnor U5359 (N_5359,N_4881,N_4889);
xnor U5360 (N_5360,N_5027,N_4512);
and U5361 (N_5361,N_4879,N_4509);
and U5362 (N_5362,N_4540,N_4838);
nand U5363 (N_5363,N_5019,N_4965);
nand U5364 (N_5364,N_4516,N_4515);
nor U5365 (N_5365,N_4588,N_4548);
or U5366 (N_5366,N_4710,N_4669);
or U5367 (N_5367,N_4599,N_4836);
xor U5368 (N_5368,N_4616,N_4854);
or U5369 (N_5369,N_5189,N_5108);
nand U5370 (N_5370,N_4912,N_4997);
xor U5371 (N_5371,N_5229,N_5001);
and U5372 (N_5372,N_5024,N_5028);
and U5373 (N_5373,N_4573,N_5018);
nand U5374 (N_5374,N_4744,N_5208);
nor U5375 (N_5375,N_4756,N_4541);
and U5376 (N_5376,N_4581,N_4553);
and U5377 (N_5377,N_5182,N_4902);
nor U5378 (N_5378,N_5183,N_4923);
xor U5379 (N_5379,N_5194,N_4947);
nor U5380 (N_5380,N_5065,N_5225);
nand U5381 (N_5381,N_4983,N_4847);
or U5382 (N_5382,N_5239,N_5113);
or U5383 (N_5383,N_4508,N_4921);
xor U5384 (N_5384,N_5046,N_4831);
and U5385 (N_5385,N_4717,N_4577);
or U5386 (N_5386,N_5025,N_4602);
and U5387 (N_5387,N_4639,N_4874);
nor U5388 (N_5388,N_5126,N_5214);
and U5389 (N_5389,N_4857,N_5243);
or U5390 (N_5390,N_4972,N_5129);
nor U5391 (N_5391,N_4547,N_4614);
nor U5392 (N_5392,N_4585,N_5246);
xor U5393 (N_5393,N_4644,N_4969);
and U5394 (N_5394,N_4883,N_4613);
or U5395 (N_5395,N_4907,N_5238);
nand U5396 (N_5396,N_4903,N_4688);
nor U5397 (N_5397,N_5091,N_4643);
xor U5398 (N_5398,N_4723,N_5005);
and U5399 (N_5399,N_5038,N_4981);
or U5400 (N_5400,N_5009,N_4609);
nor U5401 (N_5401,N_4886,N_5090);
nor U5402 (N_5402,N_4792,N_4682);
nand U5403 (N_5403,N_5150,N_4991);
nor U5404 (N_5404,N_4526,N_4955);
and U5405 (N_5405,N_4887,N_4716);
xnor U5406 (N_5406,N_5033,N_4528);
and U5407 (N_5407,N_5179,N_4637);
xnor U5408 (N_5408,N_4571,N_5207);
nor U5409 (N_5409,N_4595,N_5124);
xor U5410 (N_5410,N_4703,N_5055);
nand U5411 (N_5411,N_4694,N_4619);
nor U5412 (N_5412,N_5067,N_5054);
xor U5413 (N_5413,N_4803,N_4782);
nand U5414 (N_5414,N_5223,N_5068);
and U5415 (N_5415,N_4868,N_4659);
or U5416 (N_5416,N_5130,N_4552);
and U5417 (N_5417,N_4999,N_4911);
and U5418 (N_5418,N_4591,N_4804);
and U5419 (N_5419,N_4759,N_4908);
xnor U5420 (N_5420,N_4718,N_4530);
nand U5421 (N_5421,N_4899,N_4818);
nor U5422 (N_5422,N_4945,N_5040);
xnor U5423 (N_5423,N_4771,N_5212);
xor U5424 (N_5424,N_4727,N_4687);
nand U5425 (N_5425,N_5127,N_4627);
and U5426 (N_5426,N_5242,N_4749);
nor U5427 (N_5427,N_5145,N_4733);
or U5428 (N_5428,N_5050,N_5216);
or U5429 (N_5429,N_4529,N_4521);
and U5430 (N_5430,N_5087,N_4586);
xor U5431 (N_5431,N_4913,N_5186);
nand U5432 (N_5432,N_4835,N_4713);
and U5433 (N_5433,N_4862,N_4578);
or U5434 (N_5434,N_4918,N_4957);
nand U5435 (N_5435,N_4778,N_4707);
nand U5436 (N_5436,N_5021,N_4926);
or U5437 (N_5437,N_5117,N_5226);
or U5438 (N_5438,N_5230,N_4583);
or U5439 (N_5439,N_4870,N_4797);
nor U5440 (N_5440,N_4600,N_5104);
xor U5441 (N_5441,N_4631,N_4809);
and U5442 (N_5442,N_4653,N_4786);
nand U5443 (N_5443,N_4692,N_5151);
nor U5444 (N_5444,N_5192,N_4844);
and U5445 (N_5445,N_5052,N_4748);
xnor U5446 (N_5446,N_4954,N_4948);
or U5447 (N_5447,N_4880,N_4828);
and U5448 (N_5448,N_5099,N_4853);
nor U5449 (N_5449,N_4882,N_4917);
or U5450 (N_5450,N_4520,N_5171);
and U5451 (N_5451,N_4867,N_5114);
and U5452 (N_5452,N_5152,N_4603);
nand U5453 (N_5453,N_5170,N_4539);
or U5454 (N_5454,N_4712,N_5070);
xnor U5455 (N_5455,N_4675,N_5062);
nand U5456 (N_5456,N_4990,N_5173);
and U5457 (N_5457,N_4623,N_4670);
and U5458 (N_5458,N_4842,N_4776);
nor U5459 (N_5459,N_4615,N_5105);
or U5460 (N_5460,N_4634,N_4829);
nor U5461 (N_5461,N_4704,N_4774);
or U5462 (N_5462,N_4525,N_5042);
xnor U5463 (N_5463,N_4822,N_4690);
or U5464 (N_5464,N_5141,N_5166);
nand U5465 (N_5465,N_5101,N_4900);
xnor U5466 (N_5466,N_5049,N_5138);
xnor U5467 (N_5467,N_4505,N_4796);
and U5468 (N_5468,N_4960,N_4673);
and U5469 (N_5469,N_4940,N_5044);
and U5470 (N_5470,N_4855,N_4574);
nand U5471 (N_5471,N_5078,N_5053);
or U5472 (N_5472,N_5131,N_4914);
nand U5473 (N_5473,N_4784,N_4554);
xnor U5474 (N_5474,N_5123,N_4807);
nand U5475 (N_5475,N_5155,N_5210);
or U5476 (N_5476,N_4989,N_4768);
or U5477 (N_5477,N_4750,N_4785);
xor U5478 (N_5478,N_5072,N_5069);
nand U5479 (N_5479,N_4587,N_4546);
xnor U5480 (N_5480,N_4760,N_4916);
nand U5481 (N_5481,N_5103,N_4936);
nand U5482 (N_5482,N_4563,N_4606);
or U5483 (N_5483,N_4645,N_4576);
xor U5484 (N_5484,N_4975,N_5000);
xor U5485 (N_5485,N_4994,N_5198);
xnor U5486 (N_5486,N_4572,N_4958);
xor U5487 (N_5487,N_5222,N_4766);
and U5488 (N_5488,N_4543,N_4668);
nand U5489 (N_5489,N_4681,N_4638);
nor U5490 (N_5490,N_4513,N_4824);
nor U5491 (N_5491,N_4654,N_5202);
and U5492 (N_5492,N_4892,N_4801);
and U5493 (N_5493,N_4683,N_4993);
nand U5494 (N_5494,N_4781,N_4511);
xnor U5495 (N_5495,N_4962,N_4745);
nor U5496 (N_5496,N_4852,N_4834);
nor U5497 (N_5497,N_4755,N_5094);
nand U5498 (N_5498,N_4843,N_4597);
or U5499 (N_5499,N_5176,N_5007);
nor U5500 (N_5500,N_4795,N_5167);
or U5501 (N_5501,N_4519,N_4711);
nand U5502 (N_5502,N_4777,N_4562);
nor U5503 (N_5503,N_5011,N_5092);
or U5504 (N_5504,N_5156,N_5169);
nor U5505 (N_5505,N_4696,N_5217);
nand U5506 (N_5506,N_4934,N_4758);
nand U5507 (N_5507,N_5064,N_4708);
nand U5508 (N_5508,N_4893,N_4763);
and U5509 (N_5509,N_4762,N_5201);
or U5510 (N_5510,N_4671,N_5245);
nand U5511 (N_5511,N_5236,N_4676);
xnor U5512 (N_5512,N_4742,N_5061);
or U5513 (N_5513,N_5006,N_5158);
nor U5514 (N_5514,N_5098,N_4904);
nand U5515 (N_5515,N_5010,N_4754);
nand U5516 (N_5516,N_4974,N_5172);
nand U5517 (N_5517,N_5058,N_4746);
and U5518 (N_5518,N_5063,N_5089);
or U5519 (N_5519,N_5232,N_4664);
and U5520 (N_5520,N_4660,N_4950);
and U5521 (N_5521,N_4895,N_4561);
nand U5522 (N_5522,N_4770,N_5224);
nand U5523 (N_5523,N_4642,N_4719);
and U5524 (N_5524,N_5102,N_4632);
nand U5525 (N_5525,N_4885,N_4565);
nor U5526 (N_5526,N_4767,N_4979);
or U5527 (N_5527,N_4593,N_5079);
nand U5528 (N_5528,N_5227,N_4626);
nor U5529 (N_5529,N_5016,N_4966);
nand U5530 (N_5530,N_4641,N_4709);
and U5531 (N_5531,N_5213,N_4930);
or U5532 (N_5532,N_4819,N_5015);
nor U5533 (N_5533,N_4734,N_4992);
xor U5534 (N_5534,N_4507,N_4527);
nand U5535 (N_5535,N_4996,N_5111);
and U5536 (N_5536,N_4848,N_5209);
and U5537 (N_5537,N_4504,N_5249);
nand U5538 (N_5538,N_4570,N_5026);
nor U5539 (N_5539,N_5060,N_4538);
nor U5540 (N_5540,N_4607,N_4537);
or U5541 (N_5541,N_4856,N_4677);
or U5542 (N_5542,N_4872,N_4556);
nand U5543 (N_5543,N_5059,N_4648);
xor U5544 (N_5544,N_4869,N_4729);
or U5545 (N_5545,N_4686,N_5195);
nand U5546 (N_5546,N_5034,N_5140);
xor U5547 (N_5547,N_4927,N_5181);
and U5548 (N_5548,N_4630,N_4500);
xnor U5549 (N_5549,N_4858,N_4699);
xnor U5550 (N_5550,N_5056,N_4757);
nor U5551 (N_5551,N_4666,N_4860);
nor U5552 (N_5552,N_4982,N_4812);
nand U5553 (N_5553,N_4741,N_4788);
or U5554 (N_5554,N_4799,N_5100);
xor U5555 (N_5555,N_4730,N_4941);
xnor U5556 (N_5556,N_4532,N_4544);
nor U5557 (N_5557,N_4625,N_4780);
or U5558 (N_5558,N_4736,N_4700);
xor U5559 (N_5559,N_5128,N_5146);
nor U5560 (N_5560,N_4501,N_4938);
or U5561 (N_5561,N_5075,N_4531);
and U5562 (N_5562,N_5048,N_4584);
nand U5563 (N_5563,N_4905,N_5080);
or U5564 (N_5564,N_5112,N_4840);
nor U5565 (N_5565,N_4678,N_4897);
xnor U5566 (N_5566,N_5032,N_5177);
or U5567 (N_5567,N_4580,N_4680);
nor U5568 (N_5568,N_4910,N_5206);
xnor U5569 (N_5569,N_4551,N_4953);
nor U5570 (N_5570,N_5148,N_4808);
and U5571 (N_5571,N_5142,N_4787);
and U5572 (N_5572,N_5086,N_4898);
xnor U5573 (N_5573,N_4721,N_4737);
and U5574 (N_5574,N_4647,N_4714);
nand U5575 (N_5575,N_4933,N_4502);
or U5576 (N_5576,N_4608,N_4564);
xor U5577 (N_5577,N_4691,N_4935);
xor U5578 (N_5578,N_5211,N_4752);
nand U5579 (N_5579,N_4753,N_4884);
nand U5580 (N_5580,N_5136,N_5074);
xnor U5581 (N_5581,N_4592,N_4839);
nand U5582 (N_5582,N_5017,N_4604);
or U5583 (N_5583,N_4738,N_5030);
nor U5584 (N_5584,N_5221,N_4951);
nor U5585 (N_5585,N_5220,N_4735);
and U5586 (N_5586,N_4980,N_5180);
and U5587 (N_5587,N_4590,N_5160);
xnor U5588 (N_5588,N_4534,N_4984);
xnor U5589 (N_5589,N_4783,N_4611);
and U5590 (N_5590,N_4873,N_4924);
nor U5591 (N_5591,N_5077,N_4698);
or U5592 (N_5592,N_5023,N_4685);
or U5593 (N_5593,N_4589,N_4549);
nand U5594 (N_5594,N_4649,N_4964);
nor U5595 (N_5595,N_4662,N_4928);
and U5596 (N_5596,N_4542,N_4806);
and U5597 (N_5597,N_5235,N_5093);
xnor U5598 (N_5598,N_5133,N_4988);
nor U5599 (N_5599,N_4793,N_4739);
and U5600 (N_5600,N_4657,N_4986);
nor U5601 (N_5601,N_5012,N_5066);
xnor U5602 (N_5602,N_5147,N_4830);
nor U5603 (N_5603,N_5085,N_5205);
nor U5604 (N_5604,N_4863,N_4878);
nor U5605 (N_5605,N_4567,N_4773);
nand U5606 (N_5606,N_4864,N_5193);
nand U5607 (N_5607,N_4841,N_4851);
or U5608 (N_5608,N_5137,N_4963);
nand U5609 (N_5609,N_5020,N_4956);
nor U5610 (N_5610,N_4517,N_5071);
nor U5611 (N_5611,N_4775,N_5081);
and U5612 (N_5612,N_4837,N_4555);
nor U5613 (N_5613,N_4559,N_4715);
xor U5614 (N_5614,N_4985,N_4816);
nor U5615 (N_5615,N_4582,N_5003);
xor U5616 (N_5616,N_5002,N_4931);
xor U5617 (N_5617,N_4810,N_4514);
xor U5618 (N_5618,N_4633,N_5234);
nor U5619 (N_5619,N_4877,N_4725);
nor U5620 (N_5620,N_5164,N_5196);
or U5621 (N_5621,N_4731,N_4820);
xor U5622 (N_5622,N_5149,N_4959);
xnor U5623 (N_5623,N_4612,N_4665);
nand U5624 (N_5624,N_4655,N_4968);
nand U5625 (N_5625,N_4849,N_4748);
nor U5626 (N_5626,N_4769,N_4774);
or U5627 (N_5627,N_4565,N_4821);
and U5628 (N_5628,N_4557,N_4889);
or U5629 (N_5629,N_5222,N_5085);
nand U5630 (N_5630,N_5227,N_5209);
nand U5631 (N_5631,N_4854,N_4664);
nand U5632 (N_5632,N_4965,N_5213);
xor U5633 (N_5633,N_4989,N_4644);
nor U5634 (N_5634,N_5101,N_5084);
or U5635 (N_5635,N_4538,N_4547);
xnor U5636 (N_5636,N_4609,N_4991);
or U5637 (N_5637,N_5198,N_4633);
xor U5638 (N_5638,N_5131,N_4604);
nand U5639 (N_5639,N_5217,N_4605);
nor U5640 (N_5640,N_5175,N_4817);
nand U5641 (N_5641,N_5190,N_5214);
nor U5642 (N_5642,N_4623,N_4820);
or U5643 (N_5643,N_4945,N_4659);
and U5644 (N_5644,N_4674,N_4950);
and U5645 (N_5645,N_4805,N_4956);
and U5646 (N_5646,N_4501,N_4709);
or U5647 (N_5647,N_4559,N_4976);
xor U5648 (N_5648,N_5099,N_4564);
or U5649 (N_5649,N_4552,N_4977);
nor U5650 (N_5650,N_4890,N_4807);
nor U5651 (N_5651,N_4640,N_4846);
and U5652 (N_5652,N_4602,N_5084);
nand U5653 (N_5653,N_4742,N_4514);
nor U5654 (N_5654,N_4527,N_4818);
nand U5655 (N_5655,N_4652,N_5105);
nor U5656 (N_5656,N_5180,N_4943);
or U5657 (N_5657,N_4848,N_4559);
xor U5658 (N_5658,N_4709,N_4984);
and U5659 (N_5659,N_5150,N_5229);
or U5660 (N_5660,N_5098,N_5049);
nor U5661 (N_5661,N_4743,N_4722);
or U5662 (N_5662,N_4735,N_4948);
and U5663 (N_5663,N_4515,N_4750);
and U5664 (N_5664,N_5059,N_4733);
or U5665 (N_5665,N_4721,N_4911);
or U5666 (N_5666,N_5205,N_4600);
xor U5667 (N_5667,N_4917,N_4782);
nand U5668 (N_5668,N_4639,N_5220);
nor U5669 (N_5669,N_4928,N_5051);
or U5670 (N_5670,N_4604,N_5090);
nand U5671 (N_5671,N_5108,N_5088);
nor U5672 (N_5672,N_4857,N_4904);
xnor U5673 (N_5673,N_5098,N_4845);
or U5674 (N_5674,N_5080,N_4945);
xor U5675 (N_5675,N_4845,N_4930);
or U5676 (N_5676,N_4853,N_5094);
xnor U5677 (N_5677,N_4754,N_4845);
xnor U5678 (N_5678,N_4520,N_4905);
nor U5679 (N_5679,N_5136,N_4980);
xnor U5680 (N_5680,N_5241,N_4623);
nor U5681 (N_5681,N_5064,N_5227);
or U5682 (N_5682,N_4591,N_4993);
and U5683 (N_5683,N_4631,N_4593);
nand U5684 (N_5684,N_4634,N_4678);
xnor U5685 (N_5685,N_5132,N_4504);
nand U5686 (N_5686,N_4686,N_4524);
nand U5687 (N_5687,N_4675,N_5225);
xnor U5688 (N_5688,N_5019,N_4662);
nor U5689 (N_5689,N_4727,N_4849);
or U5690 (N_5690,N_4552,N_4724);
xnor U5691 (N_5691,N_4961,N_4742);
nand U5692 (N_5692,N_5184,N_4924);
xor U5693 (N_5693,N_5034,N_5064);
nor U5694 (N_5694,N_4923,N_5026);
nand U5695 (N_5695,N_4982,N_5146);
xor U5696 (N_5696,N_4973,N_4639);
nand U5697 (N_5697,N_4717,N_5036);
and U5698 (N_5698,N_4750,N_4532);
xnor U5699 (N_5699,N_4822,N_5049);
xnor U5700 (N_5700,N_5181,N_5006);
nor U5701 (N_5701,N_5131,N_4549);
or U5702 (N_5702,N_5204,N_4508);
and U5703 (N_5703,N_4661,N_4608);
nor U5704 (N_5704,N_5006,N_5230);
or U5705 (N_5705,N_4603,N_5138);
and U5706 (N_5706,N_4752,N_5150);
and U5707 (N_5707,N_4605,N_4721);
or U5708 (N_5708,N_4846,N_5047);
or U5709 (N_5709,N_4838,N_4587);
or U5710 (N_5710,N_5096,N_5085);
nand U5711 (N_5711,N_5115,N_4501);
xor U5712 (N_5712,N_4743,N_4569);
xor U5713 (N_5713,N_4967,N_4538);
and U5714 (N_5714,N_5211,N_4883);
or U5715 (N_5715,N_4720,N_4517);
nor U5716 (N_5716,N_4836,N_5074);
and U5717 (N_5717,N_4976,N_5140);
xnor U5718 (N_5718,N_4996,N_5235);
xor U5719 (N_5719,N_5249,N_4800);
or U5720 (N_5720,N_4846,N_4572);
and U5721 (N_5721,N_4931,N_4620);
nand U5722 (N_5722,N_4729,N_5063);
or U5723 (N_5723,N_4685,N_4568);
and U5724 (N_5724,N_4565,N_4712);
nand U5725 (N_5725,N_4749,N_4808);
nor U5726 (N_5726,N_5107,N_4676);
nor U5727 (N_5727,N_4834,N_4750);
or U5728 (N_5728,N_5225,N_4651);
xor U5729 (N_5729,N_4994,N_5179);
xor U5730 (N_5730,N_4520,N_5177);
nand U5731 (N_5731,N_4669,N_4774);
and U5732 (N_5732,N_4994,N_4854);
and U5733 (N_5733,N_4783,N_5045);
nand U5734 (N_5734,N_4525,N_4938);
nand U5735 (N_5735,N_4686,N_4703);
nor U5736 (N_5736,N_5172,N_4736);
nand U5737 (N_5737,N_5041,N_4827);
nor U5738 (N_5738,N_5202,N_5097);
nand U5739 (N_5739,N_4605,N_4922);
xor U5740 (N_5740,N_4733,N_4933);
xnor U5741 (N_5741,N_5194,N_5039);
nand U5742 (N_5742,N_5046,N_4752);
nor U5743 (N_5743,N_4572,N_5113);
or U5744 (N_5744,N_5061,N_4634);
nor U5745 (N_5745,N_4971,N_5107);
or U5746 (N_5746,N_4916,N_4667);
or U5747 (N_5747,N_5039,N_5175);
and U5748 (N_5748,N_4594,N_5142);
nor U5749 (N_5749,N_4974,N_4621);
or U5750 (N_5750,N_5063,N_5083);
nand U5751 (N_5751,N_4903,N_4822);
nand U5752 (N_5752,N_5136,N_5109);
nor U5753 (N_5753,N_4533,N_4698);
nand U5754 (N_5754,N_5126,N_4907);
xnor U5755 (N_5755,N_4861,N_5077);
and U5756 (N_5756,N_4595,N_5210);
and U5757 (N_5757,N_4688,N_4753);
or U5758 (N_5758,N_5054,N_4571);
xnor U5759 (N_5759,N_5139,N_4618);
xnor U5760 (N_5760,N_4540,N_4743);
xnor U5761 (N_5761,N_4820,N_4722);
and U5762 (N_5762,N_4710,N_4934);
or U5763 (N_5763,N_4807,N_5052);
and U5764 (N_5764,N_4847,N_4715);
nor U5765 (N_5765,N_4976,N_4514);
nand U5766 (N_5766,N_4716,N_5191);
xor U5767 (N_5767,N_4914,N_4559);
nand U5768 (N_5768,N_4683,N_5018);
nor U5769 (N_5769,N_5114,N_4614);
or U5770 (N_5770,N_4852,N_4625);
nand U5771 (N_5771,N_5188,N_4533);
and U5772 (N_5772,N_5026,N_5194);
xnor U5773 (N_5773,N_4901,N_5205);
nand U5774 (N_5774,N_4727,N_5160);
and U5775 (N_5775,N_4876,N_5218);
and U5776 (N_5776,N_4522,N_5059);
xnor U5777 (N_5777,N_4749,N_5155);
and U5778 (N_5778,N_4666,N_5049);
xor U5779 (N_5779,N_4838,N_5095);
nand U5780 (N_5780,N_5017,N_4962);
and U5781 (N_5781,N_5166,N_5104);
xnor U5782 (N_5782,N_5190,N_4919);
or U5783 (N_5783,N_4634,N_4905);
or U5784 (N_5784,N_5218,N_5213);
xnor U5785 (N_5785,N_4817,N_4607);
nor U5786 (N_5786,N_5080,N_4631);
or U5787 (N_5787,N_4973,N_4582);
nand U5788 (N_5788,N_4545,N_4977);
or U5789 (N_5789,N_4720,N_5011);
or U5790 (N_5790,N_5089,N_5218);
and U5791 (N_5791,N_5105,N_4560);
and U5792 (N_5792,N_4703,N_4935);
xor U5793 (N_5793,N_4669,N_4788);
xnor U5794 (N_5794,N_4663,N_5142);
xor U5795 (N_5795,N_4883,N_4561);
nor U5796 (N_5796,N_4958,N_5132);
and U5797 (N_5797,N_4925,N_5106);
nor U5798 (N_5798,N_4539,N_4866);
nand U5799 (N_5799,N_4530,N_5039);
xor U5800 (N_5800,N_5218,N_4513);
or U5801 (N_5801,N_4923,N_4961);
nand U5802 (N_5802,N_4697,N_5118);
nand U5803 (N_5803,N_4744,N_5094);
and U5804 (N_5804,N_5159,N_4882);
nor U5805 (N_5805,N_4694,N_5204);
nand U5806 (N_5806,N_4607,N_4794);
and U5807 (N_5807,N_4546,N_5094);
nand U5808 (N_5808,N_4840,N_5216);
xor U5809 (N_5809,N_4775,N_5020);
nor U5810 (N_5810,N_4808,N_4951);
or U5811 (N_5811,N_4979,N_5136);
and U5812 (N_5812,N_4946,N_4745);
or U5813 (N_5813,N_4530,N_4941);
nand U5814 (N_5814,N_4597,N_4715);
xor U5815 (N_5815,N_4708,N_4657);
or U5816 (N_5816,N_5156,N_4593);
xnor U5817 (N_5817,N_4871,N_4607);
xor U5818 (N_5818,N_5031,N_5027);
nand U5819 (N_5819,N_5044,N_4676);
nand U5820 (N_5820,N_5038,N_5039);
nor U5821 (N_5821,N_5000,N_5022);
and U5822 (N_5822,N_4514,N_4951);
nand U5823 (N_5823,N_4718,N_4993);
and U5824 (N_5824,N_4598,N_4889);
xnor U5825 (N_5825,N_4729,N_5090);
nand U5826 (N_5826,N_5193,N_4982);
and U5827 (N_5827,N_4660,N_4944);
nand U5828 (N_5828,N_4926,N_4985);
xor U5829 (N_5829,N_4552,N_4539);
xnor U5830 (N_5830,N_5106,N_4703);
and U5831 (N_5831,N_4857,N_4680);
xor U5832 (N_5832,N_4858,N_5216);
xor U5833 (N_5833,N_5120,N_4854);
nand U5834 (N_5834,N_4746,N_4593);
nor U5835 (N_5835,N_5098,N_4674);
and U5836 (N_5836,N_4653,N_4709);
xnor U5837 (N_5837,N_5249,N_4698);
and U5838 (N_5838,N_4635,N_4844);
nor U5839 (N_5839,N_5157,N_4828);
and U5840 (N_5840,N_4586,N_4510);
nand U5841 (N_5841,N_5173,N_4537);
nor U5842 (N_5842,N_4831,N_4926);
and U5843 (N_5843,N_5109,N_4752);
nor U5844 (N_5844,N_4816,N_5204);
xor U5845 (N_5845,N_5019,N_4553);
and U5846 (N_5846,N_4667,N_4610);
xnor U5847 (N_5847,N_4971,N_4838);
xnor U5848 (N_5848,N_4933,N_5080);
or U5849 (N_5849,N_5197,N_4941);
xnor U5850 (N_5850,N_4751,N_5217);
nand U5851 (N_5851,N_4546,N_5008);
or U5852 (N_5852,N_4595,N_4992);
xnor U5853 (N_5853,N_5117,N_5113);
nand U5854 (N_5854,N_4605,N_4726);
and U5855 (N_5855,N_5083,N_4589);
xnor U5856 (N_5856,N_5153,N_5091);
or U5857 (N_5857,N_4805,N_4933);
or U5858 (N_5858,N_5072,N_5145);
nand U5859 (N_5859,N_4536,N_4504);
or U5860 (N_5860,N_4810,N_5245);
nand U5861 (N_5861,N_5015,N_4784);
xor U5862 (N_5862,N_4596,N_4694);
nand U5863 (N_5863,N_4839,N_4786);
and U5864 (N_5864,N_4963,N_4851);
nand U5865 (N_5865,N_5160,N_4748);
nor U5866 (N_5866,N_4813,N_5216);
nor U5867 (N_5867,N_5159,N_4631);
or U5868 (N_5868,N_5047,N_4958);
or U5869 (N_5869,N_5072,N_4547);
nor U5870 (N_5870,N_4551,N_4672);
or U5871 (N_5871,N_5007,N_5077);
xor U5872 (N_5872,N_4730,N_4819);
xor U5873 (N_5873,N_4523,N_5154);
or U5874 (N_5874,N_4897,N_4916);
nor U5875 (N_5875,N_4841,N_4534);
nor U5876 (N_5876,N_5052,N_4536);
xor U5877 (N_5877,N_4656,N_4872);
xor U5878 (N_5878,N_4685,N_5058);
nor U5879 (N_5879,N_5105,N_4977);
and U5880 (N_5880,N_5132,N_5174);
or U5881 (N_5881,N_4696,N_4886);
nand U5882 (N_5882,N_4588,N_4551);
and U5883 (N_5883,N_5095,N_4918);
or U5884 (N_5884,N_4975,N_4676);
nand U5885 (N_5885,N_5161,N_4665);
and U5886 (N_5886,N_5140,N_5058);
nor U5887 (N_5887,N_4709,N_4974);
nor U5888 (N_5888,N_4738,N_4747);
nand U5889 (N_5889,N_4864,N_5138);
nand U5890 (N_5890,N_5013,N_4945);
and U5891 (N_5891,N_4584,N_4836);
nand U5892 (N_5892,N_4839,N_5221);
nand U5893 (N_5893,N_4866,N_5150);
and U5894 (N_5894,N_5218,N_4587);
and U5895 (N_5895,N_5019,N_4726);
nand U5896 (N_5896,N_5247,N_5127);
nand U5897 (N_5897,N_4798,N_4702);
nor U5898 (N_5898,N_4919,N_4501);
and U5899 (N_5899,N_4801,N_5127);
or U5900 (N_5900,N_4905,N_4731);
and U5901 (N_5901,N_4658,N_4962);
nor U5902 (N_5902,N_4735,N_4828);
and U5903 (N_5903,N_4527,N_5074);
nor U5904 (N_5904,N_4569,N_4912);
and U5905 (N_5905,N_5165,N_4919);
and U5906 (N_5906,N_5248,N_4503);
nor U5907 (N_5907,N_5057,N_5205);
or U5908 (N_5908,N_5194,N_4662);
or U5909 (N_5909,N_4950,N_4865);
xor U5910 (N_5910,N_4788,N_4844);
and U5911 (N_5911,N_4697,N_5032);
xor U5912 (N_5912,N_4919,N_4683);
and U5913 (N_5913,N_4778,N_4960);
nor U5914 (N_5914,N_4611,N_4934);
nor U5915 (N_5915,N_5242,N_4526);
nand U5916 (N_5916,N_5231,N_4852);
nand U5917 (N_5917,N_4692,N_4850);
and U5918 (N_5918,N_5182,N_4937);
or U5919 (N_5919,N_4765,N_5219);
xor U5920 (N_5920,N_4823,N_4738);
or U5921 (N_5921,N_5003,N_4616);
or U5922 (N_5922,N_4876,N_5230);
and U5923 (N_5923,N_5038,N_5212);
xor U5924 (N_5924,N_4873,N_4751);
and U5925 (N_5925,N_5004,N_5055);
or U5926 (N_5926,N_5037,N_4852);
or U5927 (N_5927,N_4688,N_4560);
and U5928 (N_5928,N_4998,N_4896);
nor U5929 (N_5929,N_5199,N_4889);
or U5930 (N_5930,N_4721,N_5192);
nand U5931 (N_5931,N_4844,N_4664);
xor U5932 (N_5932,N_5055,N_5064);
and U5933 (N_5933,N_4501,N_5241);
or U5934 (N_5934,N_4527,N_4821);
nor U5935 (N_5935,N_5198,N_4610);
xnor U5936 (N_5936,N_4728,N_4680);
and U5937 (N_5937,N_4832,N_5134);
nor U5938 (N_5938,N_5190,N_4949);
and U5939 (N_5939,N_5173,N_4716);
nor U5940 (N_5940,N_4699,N_4838);
or U5941 (N_5941,N_5138,N_4604);
nor U5942 (N_5942,N_4820,N_4522);
nor U5943 (N_5943,N_4906,N_4736);
xnor U5944 (N_5944,N_4688,N_4712);
nor U5945 (N_5945,N_5162,N_4961);
xnor U5946 (N_5946,N_5020,N_4535);
nor U5947 (N_5947,N_4833,N_4512);
xnor U5948 (N_5948,N_4536,N_4844);
xor U5949 (N_5949,N_4723,N_5044);
and U5950 (N_5950,N_5126,N_5072);
xor U5951 (N_5951,N_4909,N_4632);
nand U5952 (N_5952,N_4613,N_5064);
nand U5953 (N_5953,N_4518,N_4752);
xnor U5954 (N_5954,N_4930,N_4781);
nor U5955 (N_5955,N_4919,N_4592);
nor U5956 (N_5956,N_4578,N_4868);
xor U5957 (N_5957,N_4985,N_4907);
nor U5958 (N_5958,N_5004,N_4687);
or U5959 (N_5959,N_4911,N_4557);
nand U5960 (N_5960,N_5015,N_5188);
xor U5961 (N_5961,N_4843,N_4686);
nand U5962 (N_5962,N_5157,N_5012);
or U5963 (N_5963,N_5241,N_4980);
nor U5964 (N_5964,N_5049,N_4751);
xnor U5965 (N_5965,N_4710,N_5005);
nand U5966 (N_5966,N_5047,N_5144);
or U5967 (N_5967,N_4510,N_4544);
and U5968 (N_5968,N_4513,N_4684);
or U5969 (N_5969,N_4791,N_4611);
nand U5970 (N_5970,N_5215,N_4950);
and U5971 (N_5971,N_4726,N_5152);
nand U5972 (N_5972,N_4650,N_4740);
xor U5973 (N_5973,N_5096,N_4909);
xor U5974 (N_5974,N_4970,N_5081);
and U5975 (N_5975,N_5024,N_5179);
nand U5976 (N_5976,N_5235,N_5180);
xnor U5977 (N_5977,N_5057,N_5157);
xor U5978 (N_5978,N_4717,N_5142);
or U5979 (N_5979,N_4860,N_5190);
and U5980 (N_5980,N_5135,N_4582);
nand U5981 (N_5981,N_4590,N_4970);
or U5982 (N_5982,N_4696,N_4505);
nand U5983 (N_5983,N_4854,N_4722);
nand U5984 (N_5984,N_4753,N_4869);
or U5985 (N_5985,N_5111,N_4914);
or U5986 (N_5986,N_4580,N_4864);
nand U5987 (N_5987,N_5015,N_4540);
nor U5988 (N_5988,N_4511,N_4584);
or U5989 (N_5989,N_4514,N_5147);
or U5990 (N_5990,N_4616,N_4538);
nor U5991 (N_5991,N_5034,N_4973);
or U5992 (N_5992,N_4820,N_4777);
or U5993 (N_5993,N_4908,N_5205);
xor U5994 (N_5994,N_4634,N_4749);
xnor U5995 (N_5995,N_4653,N_4753);
or U5996 (N_5996,N_4917,N_5056);
nand U5997 (N_5997,N_4652,N_5009);
nor U5998 (N_5998,N_4932,N_4835);
or U5999 (N_5999,N_5248,N_4853);
nor U6000 (N_6000,N_5972,N_5971);
or U6001 (N_6001,N_5797,N_5687);
nor U6002 (N_6002,N_5580,N_5926);
nand U6003 (N_6003,N_5478,N_5738);
xor U6004 (N_6004,N_5425,N_5415);
xor U6005 (N_6005,N_5967,N_5944);
nor U6006 (N_6006,N_5862,N_5582);
or U6007 (N_6007,N_5808,N_5493);
nand U6008 (N_6008,N_5259,N_5308);
or U6009 (N_6009,N_5282,N_5964);
nand U6010 (N_6010,N_5515,N_5578);
nand U6011 (N_6011,N_5694,N_5433);
or U6012 (N_6012,N_5288,N_5337);
and U6013 (N_6013,N_5901,N_5417);
or U6014 (N_6014,N_5625,N_5496);
xnor U6015 (N_6015,N_5439,N_5251);
nand U6016 (N_6016,N_5869,N_5688);
and U6017 (N_6017,N_5867,N_5257);
or U6018 (N_6018,N_5511,N_5931);
xnor U6019 (N_6019,N_5342,N_5829);
or U6020 (N_6020,N_5527,N_5896);
nand U6021 (N_6021,N_5773,N_5619);
or U6022 (N_6022,N_5705,N_5655);
nor U6023 (N_6023,N_5632,N_5752);
and U6024 (N_6024,N_5995,N_5507);
or U6025 (N_6025,N_5506,N_5266);
nor U6026 (N_6026,N_5398,N_5456);
nor U6027 (N_6027,N_5691,N_5546);
and U6028 (N_6028,N_5403,N_5594);
nand U6029 (N_6029,N_5495,N_5555);
nand U6030 (N_6030,N_5316,N_5999);
nand U6031 (N_6031,N_5446,N_5737);
nor U6032 (N_6032,N_5523,N_5843);
nand U6033 (N_6033,N_5882,N_5921);
nor U6034 (N_6034,N_5922,N_5634);
xor U6035 (N_6035,N_5600,N_5871);
nor U6036 (N_6036,N_5917,N_5962);
xor U6037 (N_6037,N_5556,N_5775);
xor U6038 (N_6038,N_5286,N_5330);
or U6039 (N_6039,N_5978,N_5811);
and U6040 (N_6040,N_5492,N_5335);
nor U6041 (N_6041,N_5340,N_5874);
nand U6042 (N_6042,N_5510,N_5974);
nor U6043 (N_6043,N_5293,N_5831);
xnor U6044 (N_6044,N_5660,N_5838);
nand U6045 (N_6045,N_5327,N_5389);
nor U6046 (N_6046,N_5529,N_5501);
nor U6047 (N_6047,N_5345,N_5552);
nor U6048 (N_6048,N_5519,N_5465);
xor U6049 (N_6049,N_5814,N_5699);
nor U6050 (N_6050,N_5678,N_5535);
or U6051 (N_6051,N_5489,N_5588);
nand U6052 (N_6052,N_5416,N_5405);
nand U6053 (N_6053,N_5517,N_5540);
xnor U6054 (N_6054,N_5802,N_5386);
or U6055 (N_6055,N_5991,N_5596);
nand U6056 (N_6056,N_5778,N_5396);
nand U6057 (N_6057,N_5937,N_5509);
and U6058 (N_6058,N_5887,N_5395);
or U6059 (N_6059,N_5898,N_5852);
nand U6060 (N_6060,N_5585,N_5606);
nand U6061 (N_6061,N_5708,N_5328);
nor U6062 (N_6062,N_5363,N_5455);
and U6063 (N_6063,N_5906,N_5957);
and U6064 (N_6064,N_5640,N_5323);
nand U6065 (N_6065,N_5397,N_5790);
nand U6066 (N_6066,N_5813,N_5454);
or U6067 (N_6067,N_5980,N_5450);
and U6068 (N_6068,N_5908,N_5915);
xor U6069 (N_6069,N_5444,N_5635);
nand U6070 (N_6070,N_5449,N_5430);
nand U6071 (N_6071,N_5263,N_5740);
nand U6072 (N_6072,N_5988,N_5732);
xnor U6073 (N_6073,N_5362,N_5836);
and U6074 (N_6074,N_5782,N_5984);
and U6075 (N_6075,N_5516,N_5840);
nand U6076 (N_6076,N_5593,N_5833);
xnor U6077 (N_6077,N_5521,N_5742);
or U6078 (N_6078,N_5749,N_5365);
nand U6079 (N_6079,N_5612,N_5876);
xor U6080 (N_6080,N_5992,N_5684);
xor U6081 (N_6081,N_5562,N_5968);
and U6082 (N_6082,N_5547,N_5697);
nand U6083 (N_6083,N_5534,N_5765);
xnor U6084 (N_6084,N_5916,N_5400);
nand U6085 (N_6085,N_5716,N_5357);
or U6086 (N_6086,N_5850,N_5427);
nand U6087 (N_6087,N_5313,N_5642);
nand U6088 (N_6088,N_5322,N_5611);
and U6089 (N_6089,N_5370,N_5647);
or U6090 (N_6090,N_5318,N_5924);
and U6091 (N_6091,N_5520,N_5894);
or U6092 (N_6092,N_5324,N_5756);
xor U6093 (N_6093,N_5617,N_5380);
nand U6094 (N_6094,N_5706,N_5445);
nand U6095 (N_6095,N_5628,N_5819);
xor U6096 (N_6096,N_5630,N_5762);
or U6097 (N_6097,N_5570,N_5774);
xnor U6098 (N_6098,N_5848,N_5970);
and U6099 (N_6099,N_5277,N_5723);
nor U6100 (N_6100,N_5620,N_5950);
xor U6101 (N_6101,N_5889,N_5404);
and U6102 (N_6102,N_5973,N_5614);
nand U6103 (N_6103,N_5959,N_5820);
or U6104 (N_6104,N_5294,N_5983);
or U6105 (N_6105,N_5372,N_5822);
xor U6106 (N_6106,N_5927,N_5379);
nor U6107 (N_6107,N_5865,N_5994);
or U6108 (N_6108,N_5598,N_5763);
nor U6109 (N_6109,N_5760,N_5453);
nand U6110 (N_6110,N_5998,N_5816);
nand U6111 (N_6111,N_5720,N_5576);
or U6112 (N_6112,N_5985,N_5649);
or U6113 (N_6113,N_5408,N_5485);
xnor U6114 (N_6114,N_5584,N_5276);
nand U6115 (N_6115,N_5938,N_5609);
xor U6116 (N_6116,N_5536,N_5693);
nand U6117 (N_6117,N_5436,N_5832);
or U6118 (N_6118,N_5821,N_5668);
and U6119 (N_6119,N_5583,N_5310);
or U6120 (N_6120,N_5592,N_5332);
or U6121 (N_6121,N_5890,N_5685);
nand U6122 (N_6122,N_5626,N_5700);
and U6123 (N_6123,N_5903,N_5975);
and U6124 (N_6124,N_5928,N_5951);
xor U6125 (N_6125,N_5347,N_5573);
xor U6126 (N_6126,N_5559,N_5692);
xnor U6127 (N_6127,N_5503,N_5587);
nand U6128 (N_6128,N_5261,N_5661);
or U6129 (N_6129,N_5864,N_5548);
nor U6130 (N_6130,N_5791,N_5735);
or U6131 (N_6131,N_5344,N_5273);
nor U6132 (N_6132,N_5923,N_5383);
nand U6133 (N_6133,N_5508,N_5285);
nor U6134 (N_6134,N_5657,N_5297);
and U6135 (N_6135,N_5807,N_5961);
xor U6136 (N_6136,N_5855,N_5333);
nand U6137 (N_6137,N_5558,N_5329);
nand U6138 (N_6138,N_5267,N_5252);
nor U6139 (N_6139,N_5401,N_5488);
nor U6140 (N_6140,N_5696,N_5771);
nor U6141 (N_6141,N_5448,N_5569);
nand U6142 (N_6142,N_5525,N_5772);
nor U6143 (N_6143,N_5710,N_5304);
or U6144 (N_6144,N_5334,N_5801);
or U6145 (N_6145,N_5724,N_5679);
and U6146 (N_6146,N_5853,N_5355);
and U6147 (N_6147,N_5784,N_5377);
nor U6148 (N_6148,N_5391,N_5651);
and U6149 (N_6149,N_5296,N_5250);
nand U6150 (N_6150,N_5530,N_5891);
nor U6151 (N_6151,N_5477,N_5851);
nand U6152 (N_6152,N_5256,N_5452);
and U6153 (N_6153,N_5857,N_5940);
nand U6154 (N_6154,N_5385,N_5260);
nand U6155 (N_6155,N_5919,N_5949);
nand U6156 (N_6156,N_5868,N_5652);
and U6157 (N_6157,N_5321,N_5680);
nand U6158 (N_6158,N_5438,N_5844);
or U6159 (N_6159,N_5976,N_5522);
nand U6160 (N_6160,N_5514,N_5464);
or U6161 (N_6161,N_5567,N_5841);
or U6162 (N_6162,N_5338,N_5407);
or U6163 (N_6163,N_5788,N_5755);
nor U6164 (N_6164,N_5589,N_5990);
nand U6165 (N_6165,N_5374,N_5643);
and U6166 (N_6166,N_5714,N_5789);
nand U6167 (N_6167,N_5835,N_5645);
or U6168 (N_6168,N_5764,N_5823);
xor U6169 (N_6169,N_5390,N_5480);
and U6170 (N_6170,N_5945,N_5575);
nor U6171 (N_6171,N_5910,N_5795);
nand U6172 (N_6172,N_5892,N_5447);
and U6173 (N_6173,N_5352,N_5554);
xnor U6174 (N_6174,N_5305,N_5918);
nand U6175 (N_6175,N_5262,N_5872);
nor U6176 (N_6176,N_5796,N_5794);
nand U6177 (N_6177,N_5497,N_5930);
xor U6178 (N_6178,N_5846,N_5531);
nor U6179 (N_6179,N_5943,N_5947);
or U6180 (N_6180,N_5757,N_5902);
and U6181 (N_6181,N_5818,N_5607);
and U6182 (N_6182,N_5544,N_5353);
and U6183 (N_6183,N_5553,N_5758);
nor U6184 (N_6184,N_5331,N_5402);
nor U6185 (N_6185,N_5419,N_5603);
xor U6186 (N_6186,N_5776,N_5726);
or U6187 (N_6187,N_5900,N_5842);
xor U6188 (N_6188,N_5474,N_5644);
or U6189 (N_6189,N_5845,N_5686);
and U6190 (N_6190,N_5325,N_5608);
nor U6191 (N_6191,N_5826,N_5839);
and U6192 (N_6192,N_5925,N_5828);
nand U6193 (N_6193,N_5326,N_5675);
xor U6194 (N_6194,N_5274,N_5881);
nor U6195 (N_6195,N_5504,N_5542);
xnor U6196 (N_6196,N_5499,N_5904);
xnor U6197 (N_6197,N_5551,N_5966);
or U6198 (N_6198,N_5437,N_5728);
nand U6199 (N_6199,N_5803,N_5471);
and U6200 (N_6200,N_5715,N_5911);
nor U6201 (N_6201,N_5650,N_5309);
nand U6202 (N_6202,N_5858,N_5725);
xor U6203 (N_6203,N_5487,N_5941);
and U6204 (N_6204,N_5469,N_5690);
nor U6205 (N_6205,N_5463,N_5935);
nand U6206 (N_6206,N_5781,N_5960);
nand U6207 (N_6207,N_5289,N_5494);
or U6208 (N_6208,N_5601,N_5387);
or U6209 (N_6209,N_5793,N_5722);
nand U6210 (N_6210,N_5750,N_5615);
nand U6211 (N_6211,N_5997,N_5658);
and U6212 (N_6212,N_5572,N_5360);
or U6213 (N_6213,N_5665,N_5834);
xnor U6214 (N_6214,N_5712,N_5409);
nand U6215 (N_6215,N_5648,N_5434);
or U6216 (N_6216,N_5689,N_5761);
or U6217 (N_6217,N_5743,N_5557);
xor U6218 (N_6218,N_5669,N_5748);
or U6219 (N_6219,N_5670,N_5946);
nor U6220 (N_6220,N_5443,N_5359);
or U6221 (N_6221,N_5428,N_5932);
and U6222 (N_6222,N_5281,N_5358);
and U6223 (N_6223,N_5462,N_5641);
nand U6224 (N_6224,N_5805,N_5543);
xnor U6225 (N_6225,N_5899,N_5905);
and U6226 (N_6226,N_5989,N_5751);
or U6227 (N_6227,N_5459,N_5709);
xnor U6228 (N_6228,N_5806,N_5371);
xor U6229 (N_6229,N_5311,N_5879);
xor U6230 (N_6230,N_5613,N_5315);
nor U6231 (N_6231,N_5646,N_5351);
xnor U6232 (N_6232,N_5673,N_5539);
or U6233 (N_6233,N_5541,N_5884);
or U6234 (N_6234,N_5759,N_5627);
xor U6235 (N_6235,N_5381,N_5376);
or U6236 (N_6236,N_5320,N_5356);
nor U6237 (N_6237,N_5913,N_5431);
nor U6238 (N_6238,N_5817,N_5468);
or U6239 (N_6239,N_5629,N_5295);
nand U6240 (N_6240,N_5272,N_5981);
or U6241 (N_6241,N_5498,N_5856);
xnor U6242 (N_6242,N_5800,N_5406);
and U6243 (N_6243,N_5533,N_5590);
nor U6244 (N_6244,N_5730,N_5633);
or U6245 (N_6245,N_5280,N_5618);
or U6246 (N_6246,N_5265,N_5956);
and U6247 (N_6247,N_5963,N_5880);
nand U6248 (N_6248,N_5953,N_5271);
nand U6249 (N_6249,N_5458,N_5929);
xnor U6250 (N_6250,N_5622,N_5392);
nand U6251 (N_6251,N_5299,N_5346);
or U6252 (N_6252,N_5513,N_5369);
xor U6253 (N_6253,N_5870,N_5373);
nor U6254 (N_6254,N_5662,N_5885);
and U6255 (N_6255,N_5394,N_5287);
nand U6256 (N_6256,N_5375,N_5830);
or U6257 (N_6257,N_5432,N_5676);
nand U6258 (N_6258,N_5364,N_5664);
and U6259 (N_6259,N_5312,N_5909);
or U6260 (N_6260,N_5769,N_5269);
nand U6261 (N_6261,N_5701,N_5461);
and U6262 (N_6262,N_5528,N_5537);
and U6263 (N_6263,N_5368,N_5637);
nor U6264 (N_6264,N_5399,N_5731);
and U6265 (N_6265,N_5411,N_5258);
nor U6266 (N_6266,N_5605,N_5319);
nand U6267 (N_6267,N_5666,N_5799);
and U6268 (N_6268,N_5746,N_5502);
nand U6269 (N_6269,N_5384,N_5410);
xor U6270 (N_6270,N_5354,N_5672);
xor U6271 (N_6271,N_5659,N_5422);
and U6272 (N_6272,N_5475,N_5745);
and U6273 (N_6273,N_5704,N_5291);
or U6274 (N_6274,N_5278,N_5524);
and U6275 (N_6275,N_5421,N_5599);
xnor U6276 (N_6276,N_5307,N_5610);
or U6277 (N_6277,N_5505,N_5888);
nand U6278 (N_6278,N_5895,N_5621);
xor U6279 (N_6279,N_5873,N_5993);
and U6280 (N_6280,N_5969,N_5939);
nand U6281 (N_6281,N_5702,N_5785);
and U6282 (N_6282,N_5254,N_5302);
or U6283 (N_6283,N_5736,N_5804);
nand U6284 (N_6284,N_5866,N_5770);
and U6285 (N_6285,N_5837,N_5674);
nor U6286 (N_6286,N_5563,N_5663);
and U6287 (N_6287,N_5414,N_5275);
or U6288 (N_6288,N_5977,N_5339);
and U6289 (N_6289,N_5733,N_5579);
nand U6290 (N_6290,N_5341,N_5290);
nand U6291 (N_6291,N_5656,N_5253);
nand U6292 (N_6292,N_5825,N_5907);
nand U6293 (N_6293,N_5727,N_5695);
and U6294 (N_6294,N_5624,N_5703);
or U6295 (N_6295,N_5677,N_5718);
xor U6296 (N_6296,N_5815,N_5424);
xnor U6297 (N_6297,N_5426,N_5423);
nand U6298 (N_6298,N_5810,N_5719);
or U6299 (N_6299,N_5300,N_5314);
nand U6300 (N_6300,N_5653,N_5526);
nor U6301 (N_6301,N_5481,N_5860);
nor U6302 (N_6302,N_5739,N_5744);
nor U6303 (N_6303,N_5631,N_5717);
nand U6304 (N_6304,N_5284,N_5470);
or U6305 (N_6305,N_5255,N_5766);
xor U6306 (N_6306,N_5996,N_5671);
nor U6307 (N_6307,N_5595,N_5561);
xor U6308 (N_6308,N_5538,N_5897);
xor U6309 (N_6309,N_5859,N_5350);
xnor U6310 (N_6310,N_5483,N_5568);
and U6311 (N_6311,N_5753,N_5786);
nand U6312 (N_6312,N_5875,N_5270);
xor U6313 (N_6313,N_5591,N_5279);
and U6314 (N_6314,N_5564,N_5393);
xor U6315 (N_6315,N_5707,N_5602);
and U6316 (N_6316,N_5987,N_5729);
and U6317 (N_6317,N_5747,N_5779);
nor U6318 (N_6318,N_5886,N_5348);
or U6319 (N_6319,N_5388,N_5955);
xor U6320 (N_6320,N_5442,N_5883);
and U6321 (N_6321,N_5914,N_5549);
nand U6322 (N_6322,N_5713,N_5361);
or U6323 (N_6323,N_5451,N_5849);
xnor U6324 (N_6324,N_5378,N_5482);
nor U6325 (N_6325,N_5954,N_5979);
or U6326 (N_6326,N_5982,N_5571);
nand U6327 (N_6327,N_5780,N_5306);
nor U6328 (N_6328,N_5440,N_5566);
or U6329 (N_6329,N_5616,N_5298);
or U6330 (N_6330,N_5698,N_5777);
or U6331 (N_6331,N_5787,N_5878);
and U6332 (N_6332,N_5952,N_5479);
xor U6333 (N_6333,N_5283,N_5472);
or U6334 (N_6334,N_5264,N_5500);
and U6335 (N_6335,N_5783,N_5741);
nor U6336 (N_6336,N_5682,N_5920);
nor U6337 (N_6337,N_5303,N_5317);
and U6338 (N_6338,N_5792,N_5912);
nand U6339 (N_6339,N_5366,N_5457);
nor U6340 (N_6340,N_5577,N_5893);
xor U6341 (N_6341,N_5512,N_5560);
and U6342 (N_6342,N_5683,N_5420);
nand U6343 (N_6343,N_5429,N_5934);
nand U6344 (N_6344,N_5382,N_5604);
xnor U6345 (N_6345,N_5639,N_5809);
and U6346 (N_6346,N_5636,N_5441);
xor U6347 (N_6347,N_5550,N_5933);
xnor U6348 (N_6348,N_5476,N_5654);
nor U6349 (N_6349,N_5965,N_5292);
xnor U6350 (N_6350,N_5958,N_5367);
or U6351 (N_6351,N_5638,N_5435);
or U6352 (N_6352,N_5336,N_5473);
and U6353 (N_6353,N_5349,N_5986);
and U6354 (N_6354,N_5565,N_5268);
xnor U6355 (N_6355,N_5490,N_5767);
and U6356 (N_6356,N_5681,N_5861);
nor U6357 (N_6357,N_5597,N_5466);
xnor U6358 (N_6358,N_5721,N_5847);
xor U6359 (N_6359,N_5413,N_5623);
or U6360 (N_6360,N_5942,N_5486);
nand U6361 (N_6361,N_5418,N_5484);
xnor U6362 (N_6362,N_5667,N_5491);
or U6363 (N_6363,N_5711,N_5412);
or U6364 (N_6364,N_5532,N_5948);
nor U6365 (N_6365,N_5863,N_5768);
or U6366 (N_6366,N_5734,N_5460);
and U6367 (N_6367,N_5581,N_5467);
nand U6368 (N_6368,N_5301,N_5824);
nor U6369 (N_6369,N_5586,N_5754);
or U6370 (N_6370,N_5812,N_5518);
nor U6371 (N_6371,N_5854,N_5574);
and U6372 (N_6372,N_5343,N_5827);
and U6373 (N_6373,N_5877,N_5545);
and U6374 (N_6374,N_5798,N_5936);
nand U6375 (N_6375,N_5552,N_5656);
nand U6376 (N_6376,N_5585,N_5755);
or U6377 (N_6377,N_5588,N_5566);
nor U6378 (N_6378,N_5610,N_5827);
or U6379 (N_6379,N_5288,N_5259);
and U6380 (N_6380,N_5810,N_5306);
nand U6381 (N_6381,N_5578,N_5663);
and U6382 (N_6382,N_5788,N_5638);
nor U6383 (N_6383,N_5924,N_5732);
nor U6384 (N_6384,N_5825,N_5487);
or U6385 (N_6385,N_5616,N_5793);
nand U6386 (N_6386,N_5993,N_5500);
xor U6387 (N_6387,N_5711,N_5408);
nor U6388 (N_6388,N_5294,N_5766);
xor U6389 (N_6389,N_5786,N_5311);
and U6390 (N_6390,N_5672,N_5952);
nor U6391 (N_6391,N_5714,N_5966);
nand U6392 (N_6392,N_5368,N_5659);
or U6393 (N_6393,N_5721,N_5982);
nor U6394 (N_6394,N_5600,N_5910);
nand U6395 (N_6395,N_5261,N_5442);
and U6396 (N_6396,N_5753,N_5273);
xnor U6397 (N_6397,N_5814,N_5926);
xor U6398 (N_6398,N_5273,N_5966);
xnor U6399 (N_6399,N_5597,N_5878);
nand U6400 (N_6400,N_5399,N_5678);
nand U6401 (N_6401,N_5437,N_5883);
xor U6402 (N_6402,N_5390,N_5266);
nand U6403 (N_6403,N_5300,N_5903);
nand U6404 (N_6404,N_5449,N_5490);
nor U6405 (N_6405,N_5543,N_5936);
xor U6406 (N_6406,N_5997,N_5427);
and U6407 (N_6407,N_5522,N_5841);
nor U6408 (N_6408,N_5438,N_5888);
and U6409 (N_6409,N_5800,N_5774);
and U6410 (N_6410,N_5582,N_5422);
xnor U6411 (N_6411,N_5981,N_5942);
nor U6412 (N_6412,N_5996,N_5738);
or U6413 (N_6413,N_5473,N_5386);
nand U6414 (N_6414,N_5512,N_5625);
xnor U6415 (N_6415,N_5550,N_5878);
nor U6416 (N_6416,N_5855,N_5829);
xnor U6417 (N_6417,N_5284,N_5671);
and U6418 (N_6418,N_5792,N_5317);
and U6419 (N_6419,N_5402,N_5776);
xnor U6420 (N_6420,N_5556,N_5403);
xnor U6421 (N_6421,N_5269,N_5874);
nor U6422 (N_6422,N_5767,N_5932);
xor U6423 (N_6423,N_5572,N_5570);
nand U6424 (N_6424,N_5846,N_5458);
nand U6425 (N_6425,N_5402,N_5408);
nor U6426 (N_6426,N_5307,N_5275);
nor U6427 (N_6427,N_5386,N_5489);
nand U6428 (N_6428,N_5760,N_5566);
nor U6429 (N_6429,N_5527,N_5923);
nand U6430 (N_6430,N_5577,N_5781);
and U6431 (N_6431,N_5829,N_5590);
and U6432 (N_6432,N_5516,N_5754);
and U6433 (N_6433,N_5378,N_5557);
and U6434 (N_6434,N_5807,N_5607);
xnor U6435 (N_6435,N_5532,N_5972);
and U6436 (N_6436,N_5812,N_5579);
nor U6437 (N_6437,N_5655,N_5825);
or U6438 (N_6438,N_5574,N_5316);
nand U6439 (N_6439,N_5873,N_5260);
xor U6440 (N_6440,N_5401,N_5475);
xor U6441 (N_6441,N_5681,N_5697);
nor U6442 (N_6442,N_5955,N_5267);
nor U6443 (N_6443,N_5387,N_5422);
nand U6444 (N_6444,N_5873,N_5464);
nor U6445 (N_6445,N_5676,N_5658);
xor U6446 (N_6446,N_5755,N_5428);
nand U6447 (N_6447,N_5845,N_5681);
and U6448 (N_6448,N_5990,N_5458);
xnor U6449 (N_6449,N_5692,N_5987);
nand U6450 (N_6450,N_5704,N_5746);
and U6451 (N_6451,N_5893,N_5570);
or U6452 (N_6452,N_5751,N_5986);
nor U6453 (N_6453,N_5613,N_5270);
or U6454 (N_6454,N_5447,N_5869);
xnor U6455 (N_6455,N_5355,N_5596);
nand U6456 (N_6456,N_5939,N_5537);
or U6457 (N_6457,N_5821,N_5768);
and U6458 (N_6458,N_5664,N_5866);
xnor U6459 (N_6459,N_5636,N_5558);
and U6460 (N_6460,N_5373,N_5740);
xnor U6461 (N_6461,N_5669,N_5785);
or U6462 (N_6462,N_5392,N_5279);
or U6463 (N_6463,N_5926,N_5547);
and U6464 (N_6464,N_5405,N_5432);
or U6465 (N_6465,N_5255,N_5987);
xor U6466 (N_6466,N_5507,N_5346);
nand U6467 (N_6467,N_5993,N_5841);
and U6468 (N_6468,N_5702,N_5569);
and U6469 (N_6469,N_5543,N_5455);
nand U6470 (N_6470,N_5936,N_5857);
nor U6471 (N_6471,N_5928,N_5425);
nor U6472 (N_6472,N_5338,N_5966);
nor U6473 (N_6473,N_5530,N_5411);
xor U6474 (N_6474,N_5290,N_5549);
and U6475 (N_6475,N_5866,N_5513);
or U6476 (N_6476,N_5732,N_5684);
xor U6477 (N_6477,N_5540,N_5510);
nand U6478 (N_6478,N_5347,N_5957);
or U6479 (N_6479,N_5459,N_5790);
and U6480 (N_6480,N_5574,N_5684);
and U6481 (N_6481,N_5263,N_5456);
nor U6482 (N_6482,N_5260,N_5652);
nand U6483 (N_6483,N_5387,N_5654);
and U6484 (N_6484,N_5251,N_5437);
nor U6485 (N_6485,N_5456,N_5560);
nor U6486 (N_6486,N_5322,N_5575);
and U6487 (N_6487,N_5323,N_5728);
nor U6488 (N_6488,N_5850,N_5651);
and U6489 (N_6489,N_5523,N_5284);
and U6490 (N_6490,N_5560,N_5275);
xor U6491 (N_6491,N_5558,N_5737);
and U6492 (N_6492,N_5881,N_5549);
or U6493 (N_6493,N_5561,N_5717);
nor U6494 (N_6494,N_5979,N_5762);
nand U6495 (N_6495,N_5474,N_5831);
xnor U6496 (N_6496,N_5385,N_5543);
xor U6497 (N_6497,N_5651,N_5481);
and U6498 (N_6498,N_5425,N_5991);
nor U6499 (N_6499,N_5559,N_5848);
xor U6500 (N_6500,N_5729,N_5557);
xnor U6501 (N_6501,N_5933,N_5307);
nand U6502 (N_6502,N_5830,N_5262);
and U6503 (N_6503,N_5935,N_5956);
xor U6504 (N_6504,N_5482,N_5789);
nor U6505 (N_6505,N_5763,N_5486);
or U6506 (N_6506,N_5469,N_5849);
nand U6507 (N_6507,N_5816,N_5778);
nor U6508 (N_6508,N_5256,N_5493);
nand U6509 (N_6509,N_5446,N_5523);
xnor U6510 (N_6510,N_5895,N_5327);
xor U6511 (N_6511,N_5436,N_5303);
or U6512 (N_6512,N_5385,N_5669);
xor U6513 (N_6513,N_5385,N_5833);
xnor U6514 (N_6514,N_5951,N_5609);
or U6515 (N_6515,N_5593,N_5400);
or U6516 (N_6516,N_5286,N_5497);
xor U6517 (N_6517,N_5284,N_5869);
nand U6518 (N_6518,N_5297,N_5822);
xnor U6519 (N_6519,N_5394,N_5649);
or U6520 (N_6520,N_5585,N_5794);
xnor U6521 (N_6521,N_5439,N_5582);
or U6522 (N_6522,N_5530,N_5693);
nor U6523 (N_6523,N_5903,N_5989);
and U6524 (N_6524,N_5330,N_5839);
nand U6525 (N_6525,N_5827,N_5580);
nand U6526 (N_6526,N_5467,N_5502);
and U6527 (N_6527,N_5672,N_5807);
or U6528 (N_6528,N_5868,N_5338);
and U6529 (N_6529,N_5728,N_5930);
or U6530 (N_6530,N_5846,N_5722);
xnor U6531 (N_6531,N_5379,N_5330);
and U6532 (N_6532,N_5267,N_5301);
or U6533 (N_6533,N_5770,N_5881);
nor U6534 (N_6534,N_5500,N_5339);
nor U6535 (N_6535,N_5440,N_5559);
nand U6536 (N_6536,N_5580,N_5507);
nand U6537 (N_6537,N_5650,N_5932);
nand U6538 (N_6538,N_5485,N_5387);
xnor U6539 (N_6539,N_5265,N_5971);
xor U6540 (N_6540,N_5404,N_5546);
xor U6541 (N_6541,N_5862,N_5809);
and U6542 (N_6542,N_5981,N_5408);
xnor U6543 (N_6543,N_5719,N_5854);
nor U6544 (N_6544,N_5326,N_5781);
nor U6545 (N_6545,N_5884,N_5956);
or U6546 (N_6546,N_5406,N_5673);
nor U6547 (N_6547,N_5419,N_5569);
or U6548 (N_6548,N_5681,N_5406);
nor U6549 (N_6549,N_5305,N_5314);
or U6550 (N_6550,N_5565,N_5583);
xnor U6551 (N_6551,N_5721,N_5697);
and U6552 (N_6552,N_5715,N_5658);
or U6553 (N_6553,N_5888,N_5279);
xor U6554 (N_6554,N_5676,N_5500);
and U6555 (N_6555,N_5258,N_5779);
nor U6556 (N_6556,N_5563,N_5806);
nand U6557 (N_6557,N_5677,N_5383);
and U6558 (N_6558,N_5973,N_5438);
or U6559 (N_6559,N_5555,N_5524);
nor U6560 (N_6560,N_5328,N_5840);
and U6561 (N_6561,N_5715,N_5815);
or U6562 (N_6562,N_5257,N_5973);
nor U6563 (N_6563,N_5948,N_5882);
nor U6564 (N_6564,N_5304,N_5751);
and U6565 (N_6565,N_5792,N_5892);
xnor U6566 (N_6566,N_5644,N_5564);
nor U6567 (N_6567,N_5948,N_5578);
xnor U6568 (N_6568,N_5736,N_5905);
and U6569 (N_6569,N_5339,N_5641);
nand U6570 (N_6570,N_5909,N_5360);
or U6571 (N_6571,N_5559,N_5397);
and U6572 (N_6572,N_5956,N_5820);
nor U6573 (N_6573,N_5345,N_5703);
xnor U6574 (N_6574,N_5681,N_5959);
xnor U6575 (N_6575,N_5953,N_5556);
or U6576 (N_6576,N_5951,N_5629);
and U6577 (N_6577,N_5945,N_5812);
nand U6578 (N_6578,N_5843,N_5871);
nand U6579 (N_6579,N_5595,N_5957);
xor U6580 (N_6580,N_5844,N_5822);
and U6581 (N_6581,N_5323,N_5349);
nor U6582 (N_6582,N_5856,N_5460);
xor U6583 (N_6583,N_5835,N_5284);
nand U6584 (N_6584,N_5485,N_5266);
or U6585 (N_6585,N_5372,N_5709);
or U6586 (N_6586,N_5414,N_5429);
nor U6587 (N_6587,N_5990,N_5967);
nor U6588 (N_6588,N_5964,N_5329);
nand U6589 (N_6589,N_5946,N_5979);
and U6590 (N_6590,N_5328,N_5711);
nor U6591 (N_6591,N_5267,N_5725);
and U6592 (N_6592,N_5557,N_5417);
xnor U6593 (N_6593,N_5540,N_5290);
nand U6594 (N_6594,N_5333,N_5335);
or U6595 (N_6595,N_5481,N_5901);
nor U6596 (N_6596,N_5809,N_5382);
nand U6597 (N_6597,N_5555,N_5463);
nor U6598 (N_6598,N_5352,N_5343);
and U6599 (N_6599,N_5436,N_5589);
nor U6600 (N_6600,N_5645,N_5443);
nand U6601 (N_6601,N_5282,N_5277);
nand U6602 (N_6602,N_5666,N_5582);
or U6603 (N_6603,N_5849,N_5652);
xor U6604 (N_6604,N_5937,N_5786);
xnor U6605 (N_6605,N_5903,N_5423);
xnor U6606 (N_6606,N_5719,N_5602);
and U6607 (N_6607,N_5585,N_5987);
and U6608 (N_6608,N_5584,N_5266);
or U6609 (N_6609,N_5359,N_5725);
and U6610 (N_6610,N_5484,N_5759);
and U6611 (N_6611,N_5949,N_5253);
nand U6612 (N_6612,N_5285,N_5998);
or U6613 (N_6613,N_5435,N_5414);
and U6614 (N_6614,N_5429,N_5557);
nand U6615 (N_6615,N_5456,N_5769);
nor U6616 (N_6616,N_5549,N_5408);
and U6617 (N_6617,N_5989,N_5887);
nand U6618 (N_6618,N_5956,N_5706);
and U6619 (N_6619,N_5805,N_5931);
nand U6620 (N_6620,N_5317,N_5328);
or U6621 (N_6621,N_5886,N_5999);
xor U6622 (N_6622,N_5887,N_5473);
or U6623 (N_6623,N_5574,N_5861);
xnor U6624 (N_6624,N_5668,N_5857);
and U6625 (N_6625,N_5738,N_5404);
and U6626 (N_6626,N_5580,N_5590);
nand U6627 (N_6627,N_5348,N_5396);
and U6628 (N_6628,N_5698,N_5668);
and U6629 (N_6629,N_5841,N_5572);
nand U6630 (N_6630,N_5948,N_5646);
nand U6631 (N_6631,N_5550,N_5785);
nand U6632 (N_6632,N_5891,N_5524);
nor U6633 (N_6633,N_5811,N_5808);
or U6634 (N_6634,N_5711,N_5977);
nand U6635 (N_6635,N_5597,N_5902);
xnor U6636 (N_6636,N_5804,N_5255);
nand U6637 (N_6637,N_5500,N_5618);
and U6638 (N_6638,N_5996,N_5714);
nand U6639 (N_6639,N_5792,N_5321);
xor U6640 (N_6640,N_5912,N_5679);
xor U6641 (N_6641,N_5972,N_5941);
xnor U6642 (N_6642,N_5950,N_5474);
or U6643 (N_6643,N_5632,N_5443);
and U6644 (N_6644,N_5466,N_5446);
or U6645 (N_6645,N_5510,N_5351);
and U6646 (N_6646,N_5436,N_5969);
nand U6647 (N_6647,N_5936,N_5800);
xnor U6648 (N_6648,N_5650,N_5277);
or U6649 (N_6649,N_5843,N_5851);
or U6650 (N_6650,N_5555,N_5529);
xnor U6651 (N_6651,N_5915,N_5808);
xnor U6652 (N_6652,N_5948,N_5325);
and U6653 (N_6653,N_5329,N_5992);
and U6654 (N_6654,N_5698,N_5901);
nand U6655 (N_6655,N_5638,N_5959);
nand U6656 (N_6656,N_5957,N_5294);
or U6657 (N_6657,N_5582,N_5448);
xnor U6658 (N_6658,N_5332,N_5622);
nand U6659 (N_6659,N_5531,N_5503);
and U6660 (N_6660,N_5781,N_5682);
nand U6661 (N_6661,N_5950,N_5905);
or U6662 (N_6662,N_5258,N_5373);
and U6663 (N_6663,N_5276,N_5879);
and U6664 (N_6664,N_5647,N_5283);
and U6665 (N_6665,N_5708,N_5733);
nor U6666 (N_6666,N_5461,N_5905);
xor U6667 (N_6667,N_5878,N_5747);
xor U6668 (N_6668,N_5372,N_5388);
xor U6669 (N_6669,N_5965,N_5473);
nor U6670 (N_6670,N_5404,N_5287);
nand U6671 (N_6671,N_5984,N_5350);
or U6672 (N_6672,N_5641,N_5768);
xnor U6673 (N_6673,N_5924,N_5505);
xnor U6674 (N_6674,N_5668,N_5778);
or U6675 (N_6675,N_5346,N_5476);
nand U6676 (N_6676,N_5441,N_5965);
and U6677 (N_6677,N_5847,N_5360);
and U6678 (N_6678,N_5326,N_5903);
nor U6679 (N_6679,N_5410,N_5691);
and U6680 (N_6680,N_5509,N_5313);
or U6681 (N_6681,N_5347,N_5715);
nand U6682 (N_6682,N_5817,N_5354);
nor U6683 (N_6683,N_5902,N_5509);
nand U6684 (N_6684,N_5306,N_5620);
and U6685 (N_6685,N_5959,N_5523);
xnor U6686 (N_6686,N_5353,N_5470);
nor U6687 (N_6687,N_5424,N_5388);
and U6688 (N_6688,N_5725,N_5325);
xnor U6689 (N_6689,N_5275,N_5473);
xor U6690 (N_6690,N_5458,N_5493);
nor U6691 (N_6691,N_5975,N_5947);
or U6692 (N_6692,N_5993,N_5268);
or U6693 (N_6693,N_5694,N_5752);
or U6694 (N_6694,N_5486,N_5251);
xnor U6695 (N_6695,N_5326,N_5966);
and U6696 (N_6696,N_5624,N_5872);
xor U6697 (N_6697,N_5259,N_5380);
nor U6698 (N_6698,N_5773,N_5833);
xnor U6699 (N_6699,N_5538,N_5946);
nand U6700 (N_6700,N_5970,N_5484);
or U6701 (N_6701,N_5395,N_5684);
or U6702 (N_6702,N_5714,N_5794);
or U6703 (N_6703,N_5850,N_5995);
or U6704 (N_6704,N_5709,N_5490);
nand U6705 (N_6705,N_5843,N_5576);
nand U6706 (N_6706,N_5594,N_5988);
nand U6707 (N_6707,N_5847,N_5878);
nand U6708 (N_6708,N_5770,N_5417);
xnor U6709 (N_6709,N_5522,N_5930);
or U6710 (N_6710,N_5832,N_5382);
xnor U6711 (N_6711,N_5665,N_5342);
or U6712 (N_6712,N_5829,N_5975);
and U6713 (N_6713,N_5455,N_5659);
nand U6714 (N_6714,N_5727,N_5397);
nor U6715 (N_6715,N_5574,N_5455);
nor U6716 (N_6716,N_5832,N_5865);
nor U6717 (N_6717,N_5385,N_5577);
or U6718 (N_6718,N_5442,N_5876);
xnor U6719 (N_6719,N_5912,N_5736);
and U6720 (N_6720,N_5905,N_5351);
or U6721 (N_6721,N_5853,N_5960);
and U6722 (N_6722,N_5908,N_5914);
xor U6723 (N_6723,N_5794,N_5271);
and U6724 (N_6724,N_5541,N_5558);
nand U6725 (N_6725,N_5916,N_5708);
nand U6726 (N_6726,N_5696,N_5797);
and U6727 (N_6727,N_5387,N_5330);
or U6728 (N_6728,N_5738,N_5452);
and U6729 (N_6729,N_5264,N_5403);
and U6730 (N_6730,N_5853,N_5319);
or U6731 (N_6731,N_5478,N_5906);
or U6732 (N_6732,N_5833,N_5791);
nor U6733 (N_6733,N_5457,N_5835);
xor U6734 (N_6734,N_5505,N_5543);
or U6735 (N_6735,N_5375,N_5707);
xor U6736 (N_6736,N_5582,N_5495);
xnor U6737 (N_6737,N_5864,N_5976);
xnor U6738 (N_6738,N_5940,N_5534);
nor U6739 (N_6739,N_5986,N_5861);
xor U6740 (N_6740,N_5425,N_5744);
or U6741 (N_6741,N_5576,N_5514);
and U6742 (N_6742,N_5567,N_5358);
nor U6743 (N_6743,N_5793,N_5853);
or U6744 (N_6744,N_5989,N_5984);
or U6745 (N_6745,N_5603,N_5917);
or U6746 (N_6746,N_5281,N_5797);
nor U6747 (N_6747,N_5920,N_5664);
nand U6748 (N_6748,N_5673,N_5741);
xnor U6749 (N_6749,N_5671,N_5258);
nor U6750 (N_6750,N_6119,N_6162);
or U6751 (N_6751,N_6684,N_6478);
or U6752 (N_6752,N_6106,N_6205);
or U6753 (N_6753,N_6482,N_6117);
or U6754 (N_6754,N_6464,N_6532);
or U6755 (N_6755,N_6485,N_6191);
nor U6756 (N_6756,N_6235,N_6657);
xnor U6757 (N_6757,N_6335,N_6573);
or U6758 (N_6758,N_6500,N_6266);
and U6759 (N_6759,N_6419,N_6453);
nand U6760 (N_6760,N_6504,N_6725);
nand U6761 (N_6761,N_6655,N_6243);
nand U6762 (N_6762,N_6247,N_6240);
xnor U6763 (N_6763,N_6642,N_6654);
xnor U6764 (N_6764,N_6208,N_6249);
xnor U6765 (N_6765,N_6384,N_6696);
or U6766 (N_6766,N_6477,N_6392);
nor U6767 (N_6767,N_6302,N_6391);
or U6768 (N_6768,N_6533,N_6436);
nor U6769 (N_6769,N_6338,N_6328);
or U6770 (N_6770,N_6254,N_6256);
or U6771 (N_6771,N_6724,N_6172);
and U6772 (N_6772,N_6271,N_6300);
nand U6773 (N_6773,N_6709,N_6596);
nor U6774 (N_6774,N_6195,N_6131);
and U6775 (N_6775,N_6231,N_6171);
and U6776 (N_6776,N_6451,N_6039);
nand U6777 (N_6777,N_6074,N_6652);
and U6778 (N_6778,N_6149,N_6251);
and U6779 (N_6779,N_6364,N_6093);
and U6780 (N_6780,N_6111,N_6327);
nor U6781 (N_6781,N_6530,N_6207);
xnor U6782 (N_6782,N_6135,N_6002);
or U6783 (N_6783,N_6321,N_6013);
nor U6784 (N_6784,N_6662,N_6033);
nand U6785 (N_6785,N_6192,N_6151);
nand U6786 (N_6786,N_6287,N_6361);
xor U6787 (N_6787,N_6625,N_6520);
nor U6788 (N_6788,N_6687,N_6062);
nand U6789 (N_6789,N_6544,N_6210);
xnor U6790 (N_6790,N_6579,N_6114);
nand U6791 (N_6791,N_6692,N_6095);
nand U6792 (N_6792,N_6529,N_6649);
xnor U6793 (N_6793,N_6206,N_6682);
or U6794 (N_6794,N_6047,N_6679);
or U6795 (N_6795,N_6120,N_6020);
xnor U6796 (N_6796,N_6136,N_6517);
and U6797 (N_6797,N_6499,N_6027);
and U6798 (N_6798,N_6217,N_6648);
nand U6799 (N_6799,N_6647,N_6034);
nor U6800 (N_6800,N_6317,N_6496);
xor U6801 (N_6801,N_6351,N_6509);
or U6802 (N_6802,N_6429,N_6275);
and U6803 (N_6803,N_6422,N_6581);
or U6804 (N_6804,N_6009,N_6595);
xnor U6805 (N_6805,N_6703,N_6713);
xor U6806 (N_6806,N_6610,N_6183);
nor U6807 (N_6807,N_6615,N_6718);
or U6808 (N_6808,N_6090,N_6352);
xor U6809 (N_6809,N_6326,N_6069);
nor U6810 (N_6810,N_6267,N_6688);
xor U6811 (N_6811,N_6410,N_6345);
nand U6812 (N_6812,N_6049,N_6055);
xor U6813 (N_6813,N_6236,N_6298);
xor U6814 (N_6814,N_6105,N_6347);
or U6815 (N_6815,N_6314,N_6058);
and U6816 (N_6816,N_6148,N_6323);
xnor U6817 (N_6817,N_6081,N_6746);
xnor U6818 (N_6818,N_6346,N_6209);
nand U6819 (N_6819,N_6241,N_6639);
xor U6820 (N_6820,N_6054,N_6447);
xor U6821 (N_6821,N_6253,N_6375);
nor U6822 (N_6822,N_6014,N_6186);
or U6823 (N_6823,N_6229,N_6040);
or U6824 (N_6824,N_6094,N_6501);
nor U6825 (N_6825,N_6248,N_6582);
and U6826 (N_6826,N_6366,N_6474);
nor U6827 (N_6827,N_6194,N_6255);
xor U6828 (N_6828,N_6401,N_6045);
nor U6829 (N_6829,N_6362,N_6490);
or U6830 (N_6830,N_6001,N_6641);
or U6831 (N_6831,N_6404,N_6720);
nand U6832 (N_6832,N_6052,N_6091);
nand U6833 (N_6833,N_6580,N_6082);
or U6834 (N_6834,N_6083,N_6374);
xnor U6835 (N_6835,N_6681,N_6502);
nor U6836 (N_6836,N_6599,N_6658);
and U6837 (N_6837,N_6296,N_6279);
nand U6838 (N_6838,N_6032,N_6546);
or U6839 (N_6839,N_6733,N_6409);
nor U6840 (N_6840,N_6332,N_6378);
xor U6841 (N_6841,N_6668,N_6402);
xnor U6842 (N_6842,N_6073,N_6115);
nor U6843 (N_6843,N_6101,N_6591);
xor U6844 (N_6844,N_6683,N_6589);
and U6845 (N_6845,N_6166,N_6739);
nor U6846 (N_6846,N_6435,N_6524);
nand U6847 (N_6847,N_6437,N_6293);
or U6848 (N_6848,N_6277,N_6265);
xor U6849 (N_6849,N_6008,N_6426);
or U6850 (N_6850,N_6598,N_6356);
xnor U6851 (N_6851,N_6433,N_6350);
nand U6852 (N_6852,N_6038,N_6237);
nand U6853 (N_6853,N_6446,N_6560);
or U6854 (N_6854,N_6637,N_6165);
xnor U6855 (N_6855,N_6263,N_6694);
nor U6856 (N_6856,N_6349,N_6078);
and U6857 (N_6857,N_6489,N_6612);
nor U6858 (N_6858,N_6367,N_6479);
nor U6859 (N_6859,N_6553,N_6299);
nor U6860 (N_6860,N_6170,N_6077);
and U6861 (N_6861,N_6390,N_6487);
xnor U6862 (N_6862,N_6202,N_6548);
xnor U6863 (N_6863,N_6234,N_6449);
or U6864 (N_6864,N_6379,N_6128);
and U6865 (N_6865,N_6215,N_6528);
nor U6866 (N_6866,N_6018,N_6304);
xor U6867 (N_6867,N_6731,N_6567);
nand U6868 (N_6868,N_6159,N_6118);
and U6869 (N_6869,N_6674,N_6444);
or U6870 (N_6870,N_6512,N_6646);
xor U6871 (N_6871,N_6023,N_6605);
nand U6872 (N_6872,N_6365,N_6603);
or U6873 (N_6873,N_6129,N_6408);
nand U6874 (N_6874,N_6611,N_6188);
xnor U6875 (N_6875,N_6538,N_6656);
and U6876 (N_6876,N_6158,N_6723);
nor U6877 (N_6877,N_6664,N_6475);
and U6878 (N_6878,N_6734,N_6413);
nand U6879 (N_6879,N_6385,N_6357);
nor U6880 (N_6880,N_6221,N_6511);
xor U6881 (N_6881,N_6369,N_6308);
and U6882 (N_6882,N_6689,N_6089);
nor U6883 (N_6883,N_6130,N_6303);
nor U6884 (N_6884,N_6650,N_6334);
or U6885 (N_6885,N_6421,N_6010);
nand U6886 (N_6886,N_6565,N_6185);
or U6887 (N_6887,N_6626,N_6187);
xor U6888 (N_6888,N_6712,N_6225);
xor U6889 (N_6889,N_6693,N_6330);
nor U6890 (N_6890,N_6179,N_6109);
xnor U6891 (N_6891,N_6295,N_6643);
and U6892 (N_6892,N_6577,N_6454);
nand U6893 (N_6893,N_6415,N_6294);
nand U6894 (N_6894,N_6617,N_6706);
xor U6895 (N_6895,N_6462,N_6672);
or U6896 (N_6896,N_6306,N_6588);
and U6897 (N_6897,N_6561,N_6070);
nand U6898 (N_6898,N_6311,N_6125);
nand U6899 (N_6899,N_6666,N_6121);
nand U6900 (N_6900,N_6498,N_6678);
xnor U6901 (N_6901,N_6459,N_6284);
and U6902 (N_6902,N_6395,N_6080);
nand U6903 (N_6903,N_6383,N_6640);
or U6904 (N_6904,N_6745,N_6238);
and U6905 (N_6905,N_6259,N_6470);
nor U6906 (N_6906,N_6735,N_6196);
or U6907 (N_6907,N_6022,N_6584);
nor U6908 (N_6908,N_6432,N_6178);
xor U6909 (N_6909,N_6609,N_6406);
or U6910 (N_6910,N_6012,N_6212);
or U6911 (N_6911,N_6137,N_6430);
or U6912 (N_6912,N_6025,N_6442);
nor U6913 (N_6913,N_6086,N_6285);
and U6914 (N_6914,N_6604,N_6389);
nor U6915 (N_6915,N_6292,N_6601);
nand U6916 (N_6916,N_6585,N_6028);
or U6917 (N_6917,N_6484,N_6112);
nor U6918 (N_6918,N_6732,N_6536);
xnor U6919 (N_6919,N_6549,N_6301);
and U6920 (N_6920,N_6543,N_6157);
xnor U6921 (N_6921,N_6250,N_6239);
and U6922 (N_6922,N_6036,N_6730);
xor U6923 (N_6923,N_6164,N_6305);
nor U6924 (N_6924,N_6113,N_6452);
nand U6925 (N_6925,N_6274,N_6563);
and U6926 (N_6926,N_6515,N_6665);
xor U6927 (N_6927,N_6522,N_6198);
nand U6928 (N_6928,N_6636,N_6562);
nor U6929 (N_6929,N_6373,N_6620);
nor U6930 (N_6930,N_6331,N_6597);
nor U6931 (N_6931,N_6747,N_6525);
xnor U6932 (N_6932,N_6645,N_6261);
nor U6933 (N_6933,N_6397,N_6469);
or U6934 (N_6934,N_6246,N_6019);
and U6935 (N_6935,N_6622,N_6030);
xnor U6936 (N_6936,N_6099,N_6147);
xor U6937 (N_6937,N_6644,N_6574);
or U6938 (N_6938,N_6043,N_6486);
nand U6939 (N_6939,N_6387,N_6736);
nand U6940 (N_6940,N_6660,N_6492);
nor U6941 (N_6941,N_6100,N_6670);
nand U6942 (N_6942,N_6542,N_6476);
and U6943 (N_6943,N_6213,N_6007);
or U6944 (N_6944,N_6719,N_6051);
or U6945 (N_6945,N_6290,N_6483);
nor U6946 (N_6946,N_6439,N_6341);
and U6947 (N_6947,N_6431,N_6333);
xor U6948 (N_6948,N_6017,N_6139);
or U6949 (N_6949,N_6145,N_6363);
nand U6950 (N_6950,N_6600,N_6623);
xor U6951 (N_6951,N_6044,N_6491);
or U6952 (N_6952,N_6227,N_6613);
xnor U6953 (N_6953,N_6461,N_6150);
xor U6954 (N_6954,N_6510,N_6310);
nor U6955 (N_6955,N_6343,N_6673);
and U6956 (N_6956,N_6286,N_6571);
xor U6957 (N_6957,N_6594,N_6144);
xnor U6958 (N_6958,N_6537,N_6031);
nor U6959 (N_6959,N_6003,N_6737);
or U6960 (N_6960,N_6193,N_6228);
or U6961 (N_6961,N_6418,N_6270);
and U6962 (N_6962,N_6445,N_6506);
and U6963 (N_6963,N_6488,N_6508);
xnor U6964 (N_6964,N_6480,N_6738);
or U6965 (N_6965,N_6230,N_6152);
xnor U6966 (N_6966,N_6715,N_6184);
xnor U6967 (N_6967,N_6042,N_6060);
xnor U6968 (N_6968,N_6521,N_6315);
xnor U6969 (N_6969,N_6667,N_6110);
xnor U6970 (N_6970,N_6691,N_6201);
nand U6971 (N_6971,N_6057,N_6233);
or U6972 (N_6972,N_6319,N_6168);
or U6973 (N_6973,N_6400,N_6222);
xnor U6974 (N_6974,N_6556,N_6116);
and U6975 (N_6975,N_6122,N_6307);
or U6976 (N_6976,N_6289,N_6182);
xor U6977 (N_6977,N_6742,N_6368);
nor U6978 (N_6978,N_6214,N_6575);
or U6979 (N_6979,N_6280,N_6547);
or U6980 (N_6980,N_6721,N_6141);
and U6981 (N_6981,N_6472,N_6075);
and U6982 (N_6982,N_6348,N_6518);
nor U6983 (N_6983,N_6634,N_6695);
nor U6984 (N_6984,N_6420,N_6163);
nor U6985 (N_6985,N_6282,N_6336);
and U6986 (N_6986,N_6153,N_6393);
or U6987 (N_6987,N_6358,N_6635);
and U6988 (N_6988,N_6414,N_6108);
nand U6989 (N_6989,N_6272,N_6046);
and U6990 (N_6990,N_6329,N_6405);
xnor U6991 (N_6991,N_6748,N_6072);
nor U6992 (N_6992,N_6608,N_6219);
nand U6993 (N_6993,N_6370,N_6258);
nand U6994 (N_6994,N_6088,N_6377);
and U6995 (N_6995,N_6593,N_6539);
nand U6996 (N_6996,N_6717,N_6386);
nand U6997 (N_6997,N_6026,N_6318);
nand U6998 (N_6998,N_6388,N_6661);
nor U6999 (N_6999,N_6167,N_6450);
or U7000 (N_7000,N_6325,N_6507);
and U7001 (N_7001,N_6519,N_6606);
and U7002 (N_7002,N_6056,N_6160);
or U7003 (N_7003,N_6616,N_6382);
nor U7004 (N_7004,N_6211,N_6516);
nor U7005 (N_7005,N_6138,N_6557);
or U7006 (N_7006,N_6006,N_6079);
and U7007 (N_7007,N_6342,N_6244);
or U7008 (N_7008,N_6220,N_6276);
or U7009 (N_7009,N_6465,N_6590);
nand U7010 (N_7010,N_6704,N_6176);
xnor U7011 (N_7011,N_6197,N_6632);
and U7012 (N_7012,N_6627,N_6190);
and U7013 (N_7013,N_6558,N_6705);
nand U7014 (N_7014,N_6154,N_6523);
xor U7015 (N_7015,N_6602,N_6226);
and U7016 (N_7016,N_6570,N_6123);
and U7017 (N_7017,N_6428,N_6064);
xnor U7018 (N_7018,N_6497,N_6103);
xor U7019 (N_7019,N_6199,N_6416);
or U7020 (N_7020,N_6624,N_6068);
nand U7021 (N_7021,N_6555,N_6189);
or U7022 (N_7022,N_6540,N_6554);
or U7023 (N_7023,N_6024,N_6685);
nor U7024 (N_7024,N_6457,N_6059);
xnor U7025 (N_7025,N_6592,N_6412);
and U7026 (N_7026,N_6155,N_6638);
and U7027 (N_7027,N_6359,N_6583);
xnor U7028 (N_7028,N_6618,N_6203);
nand U7029 (N_7029,N_6252,N_6396);
nand U7030 (N_7030,N_6156,N_6360);
or U7031 (N_7031,N_6223,N_6403);
or U7032 (N_7032,N_6380,N_6578);
or U7033 (N_7033,N_6535,N_6174);
and U7034 (N_7034,N_6481,N_6743);
or U7035 (N_7035,N_6710,N_6268);
nor U7036 (N_7036,N_6092,N_6572);
xnor U7037 (N_7037,N_6514,N_6102);
and U7038 (N_7038,N_6050,N_6471);
and U7039 (N_7039,N_6067,N_6224);
xnor U7040 (N_7040,N_6607,N_6320);
nor U7041 (N_7041,N_6085,N_6216);
nor U7042 (N_7042,N_6633,N_6722);
nand U7043 (N_7043,N_6076,N_6126);
and U7044 (N_7044,N_6621,N_6353);
xnor U7045 (N_7045,N_6005,N_6425);
or U7046 (N_7046,N_6663,N_6143);
nand U7047 (N_7047,N_6564,N_6063);
or U7048 (N_7048,N_6021,N_6729);
and U7049 (N_7049,N_6440,N_6427);
or U7050 (N_7050,N_6527,N_6727);
or U7051 (N_7051,N_6140,N_6545);
nor U7052 (N_7052,N_6381,N_6041);
xor U7053 (N_7053,N_6707,N_6630);
nand U7054 (N_7054,N_6716,N_6740);
xnor U7055 (N_7055,N_6448,N_6458);
nor U7056 (N_7056,N_6702,N_6394);
and U7057 (N_7057,N_6355,N_6443);
nand U7058 (N_7058,N_6297,N_6749);
xor U7059 (N_7059,N_6503,N_6127);
xor U7060 (N_7060,N_6744,N_6177);
nand U7061 (N_7061,N_6728,N_6048);
and U7062 (N_7062,N_6455,N_6322);
xor U7063 (N_7063,N_6000,N_6467);
or U7064 (N_7064,N_6133,N_6169);
nor U7065 (N_7065,N_6411,N_6066);
nor U7066 (N_7066,N_6671,N_6653);
and U7067 (N_7067,N_6700,N_6245);
xnor U7068 (N_7068,N_6376,N_6061);
or U7069 (N_7069,N_6035,N_6354);
xor U7070 (N_7070,N_6629,N_6541);
or U7071 (N_7071,N_6407,N_6495);
or U7072 (N_7072,N_6680,N_6142);
nand U7073 (N_7073,N_6204,N_6264);
nor U7074 (N_7074,N_6424,N_6004);
xor U7075 (N_7075,N_6441,N_6741);
xnor U7076 (N_7076,N_6659,N_6493);
and U7077 (N_7077,N_6084,N_6098);
xor U7078 (N_7078,N_6631,N_6586);
or U7079 (N_7079,N_6651,N_6344);
nor U7080 (N_7080,N_6218,N_6181);
or U7081 (N_7081,N_6371,N_6260);
nor U7082 (N_7082,N_6619,N_6566);
nor U7083 (N_7083,N_6173,N_6714);
and U7084 (N_7084,N_6677,N_6242);
nand U7085 (N_7085,N_6531,N_6283);
nor U7086 (N_7086,N_6701,N_6698);
nor U7087 (N_7087,N_6016,N_6372);
or U7088 (N_7088,N_6288,N_6697);
and U7089 (N_7089,N_6398,N_6460);
and U7090 (N_7090,N_6456,N_6132);
nor U7091 (N_7091,N_6699,N_6097);
or U7092 (N_7092,N_6096,N_6124);
and U7093 (N_7093,N_6587,N_6473);
xnor U7094 (N_7094,N_6107,N_6399);
and U7095 (N_7095,N_6434,N_6676);
nor U7096 (N_7096,N_6316,N_6337);
nor U7097 (N_7097,N_6087,N_6686);
nor U7098 (N_7098,N_6065,N_6011);
nor U7099 (N_7099,N_6552,N_6313);
or U7100 (N_7100,N_6708,N_6417);
nor U7101 (N_7101,N_6463,N_6438);
xnor U7102 (N_7102,N_6614,N_6534);
or U7103 (N_7103,N_6053,N_6711);
or U7104 (N_7104,N_6161,N_6505);
and U7105 (N_7105,N_6494,N_6569);
xnor U7106 (N_7106,N_6146,N_6309);
and U7107 (N_7107,N_6273,N_6257);
xor U7108 (N_7108,N_6104,N_6726);
nor U7109 (N_7109,N_6423,N_6312);
nor U7110 (N_7110,N_6551,N_6690);
and U7111 (N_7111,N_6628,N_6550);
xnor U7112 (N_7112,N_6669,N_6559);
and U7113 (N_7113,N_6568,N_6180);
nor U7114 (N_7114,N_6269,N_6134);
and U7115 (N_7115,N_6526,N_6200);
xnor U7116 (N_7116,N_6324,N_6675);
or U7117 (N_7117,N_6029,N_6340);
nand U7118 (N_7118,N_6071,N_6281);
nor U7119 (N_7119,N_6466,N_6468);
nor U7120 (N_7120,N_6175,N_6232);
and U7121 (N_7121,N_6262,N_6037);
xor U7122 (N_7122,N_6291,N_6576);
xnor U7123 (N_7123,N_6513,N_6015);
nand U7124 (N_7124,N_6339,N_6278);
xnor U7125 (N_7125,N_6265,N_6036);
nand U7126 (N_7126,N_6077,N_6018);
nand U7127 (N_7127,N_6418,N_6728);
nand U7128 (N_7128,N_6377,N_6710);
and U7129 (N_7129,N_6524,N_6366);
nand U7130 (N_7130,N_6249,N_6006);
xor U7131 (N_7131,N_6411,N_6246);
nand U7132 (N_7132,N_6366,N_6089);
or U7133 (N_7133,N_6562,N_6453);
nand U7134 (N_7134,N_6426,N_6744);
nor U7135 (N_7135,N_6348,N_6673);
xnor U7136 (N_7136,N_6111,N_6160);
and U7137 (N_7137,N_6720,N_6484);
xor U7138 (N_7138,N_6637,N_6360);
nand U7139 (N_7139,N_6531,N_6171);
nand U7140 (N_7140,N_6001,N_6309);
or U7141 (N_7141,N_6105,N_6030);
nand U7142 (N_7142,N_6588,N_6295);
and U7143 (N_7143,N_6743,N_6517);
or U7144 (N_7144,N_6090,N_6571);
nor U7145 (N_7145,N_6083,N_6107);
and U7146 (N_7146,N_6656,N_6379);
and U7147 (N_7147,N_6059,N_6032);
and U7148 (N_7148,N_6295,N_6691);
xnor U7149 (N_7149,N_6124,N_6333);
and U7150 (N_7150,N_6439,N_6412);
and U7151 (N_7151,N_6575,N_6024);
or U7152 (N_7152,N_6726,N_6501);
or U7153 (N_7153,N_6126,N_6483);
xor U7154 (N_7154,N_6638,N_6535);
xnor U7155 (N_7155,N_6404,N_6248);
or U7156 (N_7156,N_6029,N_6674);
or U7157 (N_7157,N_6364,N_6008);
nand U7158 (N_7158,N_6275,N_6526);
nor U7159 (N_7159,N_6702,N_6701);
and U7160 (N_7160,N_6505,N_6726);
nor U7161 (N_7161,N_6067,N_6275);
nor U7162 (N_7162,N_6433,N_6011);
nor U7163 (N_7163,N_6276,N_6193);
and U7164 (N_7164,N_6460,N_6587);
and U7165 (N_7165,N_6327,N_6352);
nand U7166 (N_7166,N_6448,N_6063);
nand U7167 (N_7167,N_6550,N_6266);
and U7168 (N_7168,N_6375,N_6012);
nand U7169 (N_7169,N_6437,N_6018);
nor U7170 (N_7170,N_6480,N_6500);
and U7171 (N_7171,N_6727,N_6382);
or U7172 (N_7172,N_6663,N_6554);
nor U7173 (N_7173,N_6274,N_6176);
or U7174 (N_7174,N_6081,N_6252);
and U7175 (N_7175,N_6028,N_6681);
nor U7176 (N_7176,N_6662,N_6586);
and U7177 (N_7177,N_6042,N_6647);
and U7178 (N_7178,N_6399,N_6017);
and U7179 (N_7179,N_6260,N_6665);
nand U7180 (N_7180,N_6418,N_6726);
or U7181 (N_7181,N_6344,N_6351);
nand U7182 (N_7182,N_6198,N_6533);
or U7183 (N_7183,N_6256,N_6472);
nor U7184 (N_7184,N_6539,N_6337);
or U7185 (N_7185,N_6246,N_6730);
nor U7186 (N_7186,N_6576,N_6366);
xor U7187 (N_7187,N_6346,N_6672);
nor U7188 (N_7188,N_6142,N_6381);
xor U7189 (N_7189,N_6371,N_6110);
nor U7190 (N_7190,N_6225,N_6391);
nor U7191 (N_7191,N_6613,N_6114);
xor U7192 (N_7192,N_6071,N_6749);
xor U7193 (N_7193,N_6241,N_6426);
nor U7194 (N_7194,N_6301,N_6016);
nand U7195 (N_7195,N_6746,N_6744);
nand U7196 (N_7196,N_6625,N_6171);
nor U7197 (N_7197,N_6582,N_6276);
nor U7198 (N_7198,N_6454,N_6486);
nor U7199 (N_7199,N_6376,N_6197);
xnor U7200 (N_7200,N_6729,N_6187);
xnor U7201 (N_7201,N_6631,N_6254);
xnor U7202 (N_7202,N_6094,N_6155);
nand U7203 (N_7203,N_6271,N_6204);
nor U7204 (N_7204,N_6033,N_6292);
nand U7205 (N_7205,N_6525,N_6331);
nand U7206 (N_7206,N_6120,N_6288);
nand U7207 (N_7207,N_6073,N_6464);
and U7208 (N_7208,N_6049,N_6058);
or U7209 (N_7209,N_6122,N_6246);
or U7210 (N_7210,N_6570,N_6315);
nand U7211 (N_7211,N_6731,N_6587);
nor U7212 (N_7212,N_6306,N_6437);
xor U7213 (N_7213,N_6233,N_6230);
nor U7214 (N_7214,N_6489,N_6130);
or U7215 (N_7215,N_6417,N_6740);
or U7216 (N_7216,N_6196,N_6244);
xor U7217 (N_7217,N_6681,N_6491);
or U7218 (N_7218,N_6205,N_6447);
nor U7219 (N_7219,N_6689,N_6100);
nor U7220 (N_7220,N_6288,N_6665);
xnor U7221 (N_7221,N_6689,N_6504);
xnor U7222 (N_7222,N_6249,N_6438);
nand U7223 (N_7223,N_6200,N_6492);
and U7224 (N_7224,N_6147,N_6106);
xor U7225 (N_7225,N_6393,N_6647);
nor U7226 (N_7226,N_6252,N_6704);
nand U7227 (N_7227,N_6387,N_6012);
nor U7228 (N_7228,N_6500,N_6524);
nand U7229 (N_7229,N_6182,N_6341);
xor U7230 (N_7230,N_6254,N_6652);
and U7231 (N_7231,N_6193,N_6559);
nand U7232 (N_7232,N_6549,N_6620);
nand U7233 (N_7233,N_6206,N_6738);
or U7234 (N_7234,N_6734,N_6159);
or U7235 (N_7235,N_6712,N_6123);
or U7236 (N_7236,N_6072,N_6192);
or U7237 (N_7237,N_6615,N_6621);
nand U7238 (N_7238,N_6179,N_6746);
xor U7239 (N_7239,N_6241,N_6147);
and U7240 (N_7240,N_6651,N_6725);
and U7241 (N_7241,N_6684,N_6371);
or U7242 (N_7242,N_6628,N_6641);
and U7243 (N_7243,N_6634,N_6318);
nor U7244 (N_7244,N_6169,N_6057);
xnor U7245 (N_7245,N_6302,N_6692);
xnor U7246 (N_7246,N_6205,N_6434);
nand U7247 (N_7247,N_6243,N_6175);
and U7248 (N_7248,N_6477,N_6421);
nor U7249 (N_7249,N_6362,N_6165);
or U7250 (N_7250,N_6131,N_6566);
nand U7251 (N_7251,N_6185,N_6082);
xnor U7252 (N_7252,N_6421,N_6167);
xor U7253 (N_7253,N_6682,N_6005);
and U7254 (N_7254,N_6142,N_6263);
nand U7255 (N_7255,N_6056,N_6706);
and U7256 (N_7256,N_6494,N_6031);
or U7257 (N_7257,N_6359,N_6373);
nor U7258 (N_7258,N_6211,N_6210);
or U7259 (N_7259,N_6416,N_6196);
xnor U7260 (N_7260,N_6645,N_6426);
or U7261 (N_7261,N_6725,N_6470);
nor U7262 (N_7262,N_6478,N_6514);
and U7263 (N_7263,N_6702,N_6207);
nand U7264 (N_7264,N_6448,N_6026);
and U7265 (N_7265,N_6251,N_6698);
and U7266 (N_7266,N_6063,N_6189);
nor U7267 (N_7267,N_6084,N_6079);
or U7268 (N_7268,N_6664,N_6116);
or U7269 (N_7269,N_6346,N_6465);
nor U7270 (N_7270,N_6159,N_6642);
nand U7271 (N_7271,N_6550,N_6581);
xor U7272 (N_7272,N_6599,N_6724);
or U7273 (N_7273,N_6379,N_6544);
and U7274 (N_7274,N_6301,N_6643);
nand U7275 (N_7275,N_6215,N_6218);
or U7276 (N_7276,N_6082,N_6070);
or U7277 (N_7277,N_6272,N_6616);
and U7278 (N_7278,N_6426,N_6024);
nand U7279 (N_7279,N_6344,N_6019);
xnor U7280 (N_7280,N_6579,N_6273);
and U7281 (N_7281,N_6325,N_6556);
xor U7282 (N_7282,N_6494,N_6013);
or U7283 (N_7283,N_6122,N_6499);
nor U7284 (N_7284,N_6519,N_6695);
nor U7285 (N_7285,N_6016,N_6264);
xnor U7286 (N_7286,N_6533,N_6713);
and U7287 (N_7287,N_6039,N_6708);
nor U7288 (N_7288,N_6258,N_6219);
and U7289 (N_7289,N_6235,N_6130);
nand U7290 (N_7290,N_6538,N_6012);
and U7291 (N_7291,N_6459,N_6478);
nor U7292 (N_7292,N_6231,N_6369);
nor U7293 (N_7293,N_6010,N_6024);
nor U7294 (N_7294,N_6684,N_6571);
xor U7295 (N_7295,N_6434,N_6094);
or U7296 (N_7296,N_6405,N_6568);
and U7297 (N_7297,N_6439,N_6689);
or U7298 (N_7298,N_6064,N_6436);
nand U7299 (N_7299,N_6408,N_6621);
and U7300 (N_7300,N_6048,N_6654);
nand U7301 (N_7301,N_6439,N_6348);
and U7302 (N_7302,N_6421,N_6546);
and U7303 (N_7303,N_6659,N_6497);
or U7304 (N_7304,N_6218,N_6711);
nor U7305 (N_7305,N_6722,N_6320);
and U7306 (N_7306,N_6163,N_6309);
and U7307 (N_7307,N_6635,N_6368);
or U7308 (N_7308,N_6223,N_6745);
nand U7309 (N_7309,N_6164,N_6457);
nand U7310 (N_7310,N_6495,N_6090);
and U7311 (N_7311,N_6529,N_6297);
and U7312 (N_7312,N_6236,N_6507);
xor U7313 (N_7313,N_6330,N_6225);
nand U7314 (N_7314,N_6319,N_6231);
nand U7315 (N_7315,N_6061,N_6216);
or U7316 (N_7316,N_6144,N_6178);
and U7317 (N_7317,N_6270,N_6130);
or U7318 (N_7318,N_6719,N_6357);
and U7319 (N_7319,N_6096,N_6086);
nor U7320 (N_7320,N_6304,N_6407);
and U7321 (N_7321,N_6064,N_6479);
nand U7322 (N_7322,N_6455,N_6267);
nand U7323 (N_7323,N_6525,N_6304);
and U7324 (N_7324,N_6377,N_6143);
or U7325 (N_7325,N_6093,N_6098);
nor U7326 (N_7326,N_6501,N_6578);
or U7327 (N_7327,N_6615,N_6511);
xnor U7328 (N_7328,N_6233,N_6143);
nor U7329 (N_7329,N_6698,N_6629);
and U7330 (N_7330,N_6639,N_6308);
nor U7331 (N_7331,N_6266,N_6399);
nand U7332 (N_7332,N_6447,N_6120);
and U7333 (N_7333,N_6468,N_6348);
and U7334 (N_7334,N_6431,N_6110);
or U7335 (N_7335,N_6534,N_6009);
nand U7336 (N_7336,N_6069,N_6591);
nor U7337 (N_7337,N_6452,N_6494);
xor U7338 (N_7338,N_6069,N_6018);
and U7339 (N_7339,N_6638,N_6275);
nand U7340 (N_7340,N_6652,N_6318);
xnor U7341 (N_7341,N_6628,N_6494);
or U7342 (N_7342,N_6495,N_6574);
nor U7343 (N_7343,N_6239,N_6030);
nand U7344 (N_7344,N_6300,N_6177);
or U7345 (N_7345,N_6158,N_6489);
nand U7346 (N_7346,N_6065,N_6273);
nor U7347 (N_7347,N_6087,N_6380);
nand U7348 (N_7348,N_6539,N_6168);
nand U7349 (N_7349,N_6714,N_6512);
and U7350 (N_7350,N_6053,N_6463);
nand U7351 (N_7351,N_6393,N_6303);
and U7352 (N_7352,N_6034,N_6695);
xnor U7353 (N_7353,N_6579,N_6122);
nand U7354 (N_7354,N_6040,N_6374);
nand U7355 (N_7355,N_6634,N_6172);
and U7356 (N_7356,N_6373,N_6092);
and U7357 (N_7357,N_6169,N_6071);
and U7358 (N_7358,N_6268,N_6462);
nor U7359 (N_7359,N_6213,N_6690);
xnor U7360 (N_7360,N_6166,N_6317);
nand U7361 (N_7361,N_6749,N_6026);
and U7362 (N_7362,N_6214,N_6027);
nand U7363 (N_7363,N_6275,N_6484);
or U7364 (N_7364,N_6643,N_6736);
nor U7365 (N_7365,N_6678,N_6134);
xnor U7366 (N_7366,N_6161,N_6294);
xnor U7367 (N_7367,N_6689,N_6701);
or U7368 (N_7368,N_6381,N_6001);
or U7369 (N_7369,N_6080,N_6561);
xor U7370 (N_7370,N_6122,N_6555);
xor U7371 (N_7371,N_6031,N_6714);
or U7372 (N_7372,N_6541,N_6287);
and U7373 (N_7373,N_6652,N_6537);
or U7374 (N_7374,N_6659,N_6236);
nand U7375 (N_7375,N_6253,N_6665);
or U7376 (N_7376,N_6312,N_6407);
nor U7377 (N_7377,N_6098,N_6491);
nor U7378 (N_7378,N_6734,N_6239);
xor U7379 (N_7379,N_6522,N_6575);
or U7380 (N_7380,N_6491,N_6585);
nand U7381 (N_7381,N_6263,N_6666);
nor U7382 (N_7382,N_6511,N_6605);
and U7383 (N_7383,N_6729,N_6139);
or U7384 (N_7384,N_6313,N_6251);
nand U7385 (N_7385,N_6320,N_6043);
nor U7386 (N_7386,N_6417,N_6368);
nand U7387 (N_7387,N_6510,N_6257);
nand U7388 (N_7388,N_6326,N_6280);
xnor U7389 (N_7389,N_6411,N_6169);
xnor U7390 (N_7390,N_6067,N_6004);
nor U7391 (N_7391,N_6056,N_6088);
and U7392 (N_7392,N_6017,N_6703);
nand U7393 (N_7393,N_6535,N_6103);
or U7394 (N_7394,N_6690,N_6223);
nor U7395 (N_7395,N_6208,N_6077);
nor U7396 (N_7396,N_6691,N_6305);
nor U7397 (N_7397,N_6177,N_6235);
nor U7398 (N_7398,N_6630,N_6657);
nor U7399 (N_7399,N_6588,N_6675);
xor U7400 (N_7400,N_6161,N_6327);
and U7401 (N_7401,N_6207,N_6486);
and U7402 (N_7402,N_6480,N_6544);
or U7403 (N_7403,N_6211,N_6343);
xnor U7404 (N_7404,N_6700,N_6533);
nand U7405 (N_7405,N_6214,N_6201);
nor U7406 (N_7406,N_6337,N_6145);
xnor U7407 (N_7407,N_6166,N_6466);
nor U7408 (N_7408,N_6515,N_6152);
xor U7409 (N_7409,N_6058,N_6363);
nand U7410 (N_7410,N_6613,N_6497);
xor U7411 (N_7411,N_6719,N_6356);
nor U7412 (N_7412,N_6422,N_6384);
nor U7413 (N_7413,N_6425,N_6488);
and U7414 (N_7414,N_6157,N_6304);
xnor U7415 (N_7415,N_6132,N_6625);
nor U7416 (N_7416,N_6328,N_6539);
xnor U7417 (N_7417,N_6207,N_6433);
nor U7418 (N_7418,N_6045,N_6188);
xor U7419 (N_7419,N_6706,N_6184);
and U7420 (N_7420,N_6305,N_6675);
nand U7421 (N_7421,N_6339,N_6224);
nor U7422 (N_7422,N_6273,N_6202);
nand U7423 (N_7423,N_6120,N_6174);
nor U7424 (N_7424,N_6581,N_6676);
xor U7425 (N_7425,N_6032,N_6637);
nand U7426 (N_7426,N_6112,N_6053);
nor U7427 (N_7427,N_6447,N_6216);
or U7428 (N_7428,N_6123,N_6048);
and U7429 (N_7429,N_6450,N_6101);
and U7430 (N_7430,N_6482,N_6412);
nor U7431 (N_7431,N_6419,N_6046);
nand U7432 (N_7432,N_6064,N_6497);
nand U7433 (N_7433,N_6641,N_6163);
or U7434 (N_7434,N_6118,N_6672);
nor U7435 (N_7435,N_6703,N_6487);
xor U7436 (N_7436,N_6541,N_6004);
nor U7437 (N_7437,N_6274,N_6018);
nor U7438 (N_7438,N_6633,N_6612);
nand U7439 (N_7439,N_6397,N_6611);
nor U7440 (N_7440,N_6376,N_6166);
or U7441 (N_7441,N_6553,N_6393);
nand U7442 (N_7442,N_6074,N_6377);
nand U7443 (N_7443,N_6057,N_6567);
xnor U7444 (N_7444,N_6543,N_6458);
and U7445 (N_7445,N_6049,N_6168);
and U7446 (N_7446,N_6742,N_6513);
or U7447 (N_7447,N_6464,N_6237);
and U7448 (N_7448,N_6339,N_6523);
nor U7449 (N_7449,N_6450,N_6044);
or U7450 (N_7450,N_6113,N_6302);
or U7451 (N_7451,N_6160,N_6177);
or U7452 (N_7452,N_6197,N_6412);
nand U7453 (N_7453,N_6337,N_6095);
nor U7454 (N_7454,N_6669,N_6144);
or U7455 (N_7455,N_6060,N_6261);
and U7456 (N_7456,N_6188,N_6515);
nand U7457 (N_7457,N_6385,N_6411);
nand U7458 (N_7458,N_6222,N_6350);
nand U7459 (N_7459,N_6404,N_6006);
nand U7460 (N_7460,N_6650,N_6280);
and U7461 (N_7461,N_6148,N_6348);
and U7462 (N_7462,N_6393,N_6457);
xor U7463 (N_7463,N_6025,N_6632);
or U7464 (N_7464,N_6265,N_6298);
nand U7465 (N_7465,N_6362,N_6241);
or U7466 (N_7466,N_6396,N_6111);
and U7467 (N_7467,N_6498,N_6326);
xnor U7468 (N_7468,N_6397,N_6046);
nor U7469 (N_7469,N_6409,N_6109);
xor U7470 (N_7470,N_6418,N_6582);
or U7471 (N_7471,N_6364,N_6455);
xor U7472 (N_7472,N_6039,N_6016);
nor U7473 (N_7473,N_6336,N_6553);
nand U7474 (N_7474,N_6533,N_6482);
or U7475 (N_7475,N_6608,N_6425);
and U7476 (N_7476,N_6349,N_6266);
nor U7477 (N_7477,N_6684,N_6030);
xor U7478 (N_7478,N_6453,N_6220);
nand U7479 (N_7479,N_6138,N_6444);
nand U7480 (N_7480,N_6001,N_6407);
and U7481 (N_7481,N_6425,N_6613);
nor U7482 (N_7482,N_6533,N_6040);
or U7483 (N_7483,N_6574,N_6718);
nor U7484 (N_7484,N_6308,N_6448);
nand U7485 (N_7485,N_6260,N_6282);
nor U7486 (N_7486,N_6638,N_6072);
nand U7487 (N_7487,N_6336,N_6510);
nand U7488 (N_7488,N_6439,N_6296);
and U7489 (N_7489,N_6689,N_6215);
and U7490 (N_7490,N_6650,N_6220);
nor U7491 (N_7491,N_6475,N_6098);
or U7492 (N_7492,N_6658,N_6595);
and U7493 (N_7493,N_6554,N_6480);
nor U7494 (N_7494,N_6554,N_6128);
nor U7495 (N_7495,N_6444,N_6316);
nor U7496 (N_7496,N_6535,N_6350);
nor U7497 (N_7497,N_6225,N_6688);
xnor U7498 (N_7498,N_6476,N_6098);
nand U7499 (N_7499,N_6076,N_6583);
nand U7500 (N_7500,N_7316,N_7219);
xor U7501 (N_7501,N_6888,N_7114);
or U7502 (N_7502,N_7259,N_7199);
nor U7503 (N_7503,N_7444,N_6873);
xnor U7504 (N_7504,N_7138,N_7389);
or U7505 (N_7505,N_7058,N_6823);
xnor U7506 (N_7506,N_7481,N_6998);
nand U7507 (N_7507,N_6763,N_7127);
nand U7508 (N_7508,N_6786,N_7302);
xor U7509 (N_7509,N_7380,N_7446);
nand U7510 (N_7510,N_6951,N_7355);
xnor U7511 (N_7511,N_6826,N_7336);
and U7512 (N_7512,N_7399,N_7363);
or U7513 (N_7513,N_7436,N_6965);
and U7514 (N_7514,N_6924,N_6923);
and U7515 (N_7515,N_6794,N_6760);
or U7516 (N_7516,N_7126,N_7221);
xor U7517 (N_7517,N_7120,N_7398);
nor U7518 (N_7518,N_7434,N_7124);
or U7519 (N_7519,N_7273,N_7429);
and U7520 (N_7520,N_7395,N_7320);
xor U7521 (N_7521,N_7009,N_7404);
nor U7522 (N_7522,N_6916,N_6993);
and U7523 (N_7523,N_6845,N_7313);
nor U7524 (N_7524,N_7222,N_6982);
and U7525 (N_7525,N_7425,N_6869);
and U7526 (N_7526,N_6777,N_6911);
nor U7527 (N_7527,N_7366,N_7027);
and U7528 (N_7528,N_7098,N_7490);
nand U7529 (N_7529,N_7034,N_7240);
nand U7530 (N_7530,N_7017,N_6970);
nor U7531 (N_7531,N_7411,N_7060);
and U7532 (N_7532,N_7043,N_7076);
xor U7533 (N_7533,N_6880,N_6953);
xor U7534 (N_7534,N_7191,N_7181);
or U7535 (N_7535,N_6977,N_7385);
nor U7536 (N_7536,N_7376,N_7100);
xnor U7537 (N_7537,N_7375,N_7455);
and U7538 (N_7538,N_6939,N_7142);
nand U7539 (N_7539,N_7081,N_7397);
nand U7540 (N_7540,N_7382,N_7308);
and U7541 (N_7541,N_6824,N_6788);
xor U7542 (N_7542,N_6776,N_7052);
nand U7543 (N_7543,N_7305,N_6905);
nand U7544 (N_7544,N_7450,N_7408);
nand U7545 (N_7545,N_7431,N_7284);
or U7546 (N_7546,N_7496,N_7247);
nand U7547 (N_7547,N_7208,N_7497);
nor U7548 (N_7548,N_7440,N_7447);
nor U7549 (N_7549,N_6995,N_6866);
nand U7550 (N_7550,N_7167,N_7205);
nand U7551 (N_7551,N_6886,N_7066);
and U7552 (N_7552,N_7179,N_6972);
xnor U7553 (N_7553,N_7164,N_7326);
nand U7554 (N_7554,N_6999,N_6770);
and U7555 (N_7555,N_7456,N_6932);
nor U7556 (N_7556,N_7271,N_6986);
and U7557 (N_7557,N_6810,N_7209);
or U7558 (N_7558,N_7105,N_7140);
xor U7559 (N_7559,N_6912,N_6922);
and U7560 (N_7560,N_6811,N_6834);
xnor U7561 (N_7561,N_7274,N_7227);
nand U7562 (N_7562,N_7136,N_7262);
or U7563 (N_7563,N_7419,N_7322);
nand U7564 (N_7564,N_7256,N_7049);
nand U7565 (N_7565,N_6991,N_6971);
xnor U7566 (N_7566,N_7233,N_7359);
xnor U7567 (N_7567,N_7129,N_7372);
xnor U7568 (N_7568,N_7309,N_7001);
or U7569 (N_7569,N_7347,N_7032);
xor U7570 (N_7570,N_7261,N_7439);
nor U7571 (N_7571,N_7384,N_6917);
xnor U7572 (N_7572,N_7476,N_6839);
or U7573 (N_7573,N_7280,N_7007);
nand U7574 (N_7574,N_6825,N_6938);
or U7575 (N_7575,N_7349,N_7112);
nand U7576 (N_7576,N_7148,N_7379);
nor U7577 (N_7577,N_7119,N_7048);
xnor U7578 (N_7578,N_6781,N_7364);
and U7579 (N_7579,N_6806,N_7006);
and U7580 (N_7580,N_7213,N_6915);
or U7581 (N_7581,N_7211,N_7343);
or U7582 (N_7582,N_7108,N_7215);
nor U7583 (N_7583,N_7383,N_7184);
and U7584 (N_7584,N_7332,N_6785);
xnor U7585 (N_7585,N_7405,N_6910);
nor U7586 (N_7586,N_6840,N_7123);
and U7587 (N_7587,N_7130,N_7413);
nor U7588 (N_7588,N_7278,N_7286);
nand U7589 (N_7589,N_7055,N_7226);
and U7590 (N_7590,N_7183,N_7069);
and U7591 (N_7591,N_7403,N_6945);
and U7592 (N_7592,N_7342,N_7206);
nand U7593 (N_7593,N_7202,N_7442);
nor U7594 (N_7594,N_7248,N_6909);
nand U7595 (N_7595,N_6899,N_7462);
and U7596 (N_7596,N_7482,N_6885);
nand U7597 (N_7597,N_6882,N_7352);
nor U7598 (N_7598,N_6831,N_7082);
nand U7599 (N_7599,N_7360,N_7064);
nand U7600 (N_7600,N_7498,N_7230);
nand U7601 (N_7601,N_7021,N_6989);
and U7602 (N_7602,N_6849,N_7249);
xor U7603 (N_7603,N_7279,N_6792);
xor U7604 (N_7604,N_7203,N_6992);
nand U7605 (N_7605,N_6751,N_7428);
nand U7606 (N_7606,N_6814,N_7299);
nor U7607 (N_7607,N_7198,N_7292);
and U7608 (N_7608,N_6779,N_7294);
nand U7609 (N_7609,N_6854,N_7087);
nand U7610 (N_7610,N_6818,N_7260);
and U7611 (N_7611,N_7374,N_7472);
nand U7612 (N_7612,N_7170,N_6757);
nor U7613 (N_7613,N_6758,N_7400);
xnor U7614 (N_7614,N_7153,N_7010);
nand U7615 (N_7615,N_6904,N_7406);
or U7616 (N_7616,N_7044,N_7410);
nor U7617 (N_7617,N_6830,N_7085);
and U7618 (N_7618,N_6883,N_7441);
or U7619 (N_7619,N_6765,N_6955);
xnor U7620 (N_7620,N_7212,N_7122);
nor U7621 (N_7621,N_6796,N_7297);
xnor U7622 (N_7622,N_7451,N_7077);
or U7623 (N_7623,N_7023,N_7045);
nor U7624 (N_7624,N_7465,N_7026);
nor U7625 (N_7625,N_6907,N_6931);
or U7626 (N_7626,N_7160,N_6980);
nand U7627 (N_7627,N_7104,N_7089);
xor U7628 (N_7628,N_7031,N_7437);
xnor U7629 (N_7629,N_7004,N_7396);
and U7630 (N_7630,N_7492,N_6850);
nand U7631 (N_7631,N_7121,N_7193);
nand U7632 (N_7632,N_7362,N_7390);
or U7633 (N_7633,N_6848,N_6759);
xor U7634 (N_7634,N_7051,N_7469);
nor U7635 (N_7635,N_6877,N_6929);
xnor U7636 (N_7636,N_7288,N_7282);
nand U7637 (N_7637,N_6887,N_7168);
and U7638 (N_7638,N_7185,N_7020);
xnor U7639 (N_7639,N_6895,N_6793);
nor U7640 (N_7640,N_7432,N_6855);
and U7641 (N_7641,N_7335,N_6937);
nand U7642 (N_7642,N_7341,N_7113);
or U7643 (N_7643,N_7489,N_7196);
or U7644 (N_7644,N_7345,N_6797);
or U7645 (N_7645,N_6846,N_7139);
nor U7646 (N_7646,N_7353,N_6948);
nor U7647 (N_7647,N_6985,N_7067);
xnor U7648 (N_7648,N_7304,N_7448);
or U7649 (N_7649,N_7370,N_7296);
or U7650 (N_7650,N_7158,N_7084);
and U7651 (N_7651,N_7155,N_6889);
and U7652 (N_7652,N_7257,N_7014);
xnor U7653 (N_7653,N_7102,N_6979);
and U7654 (N_7654,N_7200,N_7417);
nor U7655 (N_7655,N_6769,N_7241);
and U7656 (N_7656,N_7463,N_7188);
and U7657 (N_7657,N_7012,N_7131);
nor U7658 (N_7658,N_6768,N_7217);
and U7659 (N_7659,N_7449,N_7330);
nor U7660 (N_7660,N_7387,N_7401);
or U7661 (N_7661,N_7315,N_7300);
nand U7662 (N_7662,N_7487,N_7042);
nor U7663 (N_7663,N_6860,N_7192);
nand U7664 (N_7664,N_7486,N_6961);
and U7665 (N_7665,N_6771,N_6802);
nor U7666 (N_7666,N_7204,N_6954);
nand U7667 (N_7667,N_7059,N_7254);
nand U7668 (N_7668,N_6946,N_6871);
and U7669 (N_7669,N_6934,N_6957);
nand U7670 (N_7670,N_6997,N_7307);
and U7671 (N_7671,N_7285,N_6842);
or U7672 (N_7672,N_7224,N_7103);
or U7673 (N_7673,N_7453,N_7331);
and U7674 (N_7674,N_7071,N_6753);
nor U7675 (N_7675,N_6851,N_6772);
nand U7676 (N_7676,N_6827,N_7426);
xnor U7677 (N_7677,N_6829,N_7176);
nand U7678 (N_7678,N_7480,N_7348);
and U7679 (N_7679,N_6975,N_7145);
and U7680 (N_7680,N_7178,N_7369);
xnor U7681 (N_7681,N_7457,N_6897);
nand U7682 (N_7682,N_7289,N_7407);
nor U7683 (N_7683,N_7133,N_7479);
nor U7684 (N_7684,N_6864,N_6981);
nand U7685 (N_7685,N_7106,N_7416);
or U7686 (N_7686,N_7061,N_7218);
nand U7687 (N_7687,N_7109,N_6767);
nor U7688 (N_7688,N_7037,N_7062);
or U7689 (N_7689,N_6919,N_6941);
and U7690 (N_7690,N_7381,N_7414);
xnor U7691 (N_7691,N_7312,N_7229);
or U7692 (N_7692,N_6890,N_7162);
xnor U7693 (N_7693,N_7454,N_7325);
and U7694 (N_7694,N_7078,N_6754);
nand U7695 (N_7695,N_7156,N_6983);
and U7696 (N_7696,N_7310,N_7466);
nor U7697 (N_7697,N_7270,N_6784);
and U7698 (N_7698,N_7146,N_7412);
xnor U7699 (N_7699,N_7295,N_7018);
xor U7700 (N_7700,N_6987,N_7187);
xnor U7701 (N_7701,N_7409,N_7107);
and U7702 (N_7702,N_7111,N_6900);
and U7703 (N_7703,N_6841,N_7371);
nand U7704 (N_7704,N_7242,N_6935);
or U7705 (N_7705,N_7475,N_7232);
nand U7706 (N_7706,N_6819,N_7137);
and U7707 (N_7707,N_7197,N_7225);
xnor U7708 (N_7708,N_6790,N_7086);
nand U7709 (N_7709,N_7022,N_6942);
nor U7710 (N_7710,N_7253,N_7019);
xnor U7711 (N_7711,N_7323,N_7277);
nor U7712 (N_7712,N_6974,N_6936);
nand U7713 (N_7713,N_6926,N_7177);
or U7714 (N_7714,N_7333,N_6833);
nor U7715 (N_7715,N_6859,N_6812);
or U7716 (N_7716,N_6807,N_7420);
and U7717 (N_7717,N_7057,N_7477);
nor U7718 (N_7718,N_7090,N_7175);
xor U7719 (N_7719,N_7207,N_6906);
and U7720 (N_7720,N_7056,N_7415);
xnor U7721 (N_7721,N_6962,N_6894);
or U7722 (N_7722,N_7287,N_6875);
and U7723 (N_7723,N_7079,N_7024);
nor U7724 (N_7724,N_7250,N_7036);
xnor U7725 (N_7725,N_7269,N_6780);
nand U7726 (N_7726,N_7161,N_7228);
or U7727 (N_7727,N_6801,N_6925);
and U7728 (N_7728,N_6950,N_6863);
xor U7729 (N_7729,N_7354,N_7378);
and U7730 (N_7730,N_7460,N_6896);
and U7731 (N_7731,N_7028,N_6847);
xor U7732 (N_7732,N_7386,N_7245);
nand U7733 (N_7733,N_7268,N_6940);
xor U7734 (N_7734,N_6973,N_7246);
nor U7735 (N_7735,N_7180,N_7306);
nor U7736 (N_7736,N_7163,N_7003);
nand U7737 (N_7737,N_6967,N_7337);
nor U7738 (N_7738,N_7340,N_7095);
nand U7739 (N_7739,N_6881,N_6870);
or U7740 (N_7740,N_7467,N_6816);
and U7741 (N_7741,N_7053,N_7314);
xnor U7742 (N_7742,N_7290,N_7135);
nand U7743 (N_7743,N_7083,N_6874);
nor U7744 (N_7744,N_6856,N_6956);
nand U7745 (N_7745,N_6861,N_7125);
nor U7746 (N_7746,N_7039,N_7195);
or U7747 (N_7747,N_6943,N_7116);
nand U7748 (N_7748,N_7471,N_7461);
nor U7749 (N_7749,N_7458,N_7361);
or U7750 (N_7750,N_7025,N_7169);
nand U7751 (N_7751,N_7117,N_7073);
or U7752 (N_7752,N_7281,N_7054);
nor U7753 (N_7753,N_6867,N_7377);
nand U7754 (N_7754,N_6817,N_7238);
nand U7755 (N_7755,N_6852,N_7258);
nand U7756 (N_7756,N_6964,N_7393);
xnor U7757 (N_7757,N_7424,N_7350);
and U7758 (N_7758,N_7499,N_7165);
xor U7759 (N_7759,N_6803,N_7275);
nor U7760 (N_7760,N_6902,N_6773);
nand U7761 (N_7761,N_7252,N_6844);
or U7762 (N_7762,N_6813,N_7174);
nand U7763 (N_7763,N_6787,N_6920);
nand U7764 (N_7764,N_7035,N_7435);
nand U7765 (N_7765,N_7339,N_6928);
and U7766 (N_7766,N_7234,N_7459);
xnor U7767 (N_7767,N_6978,N_7443);
nand U7768 (N_7768,N_7239,N_6921);
or U7769 (N_7769,N_6878,N_6774);
nand U7770 (N_7770,N_6868,N_7468);
or U7771 (N_7771,N_7172,N_6944);
nand U7772 (N_7772,N_6835,N_7488);
nand U7773 (N_7773,N_6778,N_6876);
nor U7774 (N_7774,N_7351,N_7220);
nor U7775 (N_7775,N_7484,N_6838);
and U7776 (N_7776,N_7329,N_7430);
or U7777 (N_7777,N_7016,N_7373);
xnor U7778 (N_7778,N_7283,N_6750);
xnor U7779 (N_7779,N_6843,N_6799);
nor U7780 (N_7780,N_7470,N_6798);
or U7781 (N_7781,N_7072,N_6755);
nor U7782 (N_7782,N_7091,N_7088);
nor U7783 (N_7783,N_6960,N_7324);
xnor U7784 (N_7784,N_6822,N_7096);
or U7785 (N_7785,N_7311,N_6996);
nor U7786 (N_7786,N_7029,N_6984);
nor U7787 (N_7787,N_6898,N_7301);
and U7788 (N_7788,N_7128,N_6892);
nand U7789 (N_7789,N_7423,N_7092);
nand U7790 (N_7790,N_7194,N_7147);
xor U7791 (N_7791,N_7154,N_7070);
nand U7792 (N_7792,N_7151,N_7267);
or U7793 (N_7793,N_7094,N_6958);
and U7794 (N_7794,N_7063,N_6963);
nand U7795 (N_7795,N_7473,N_7358);
nor U7796 (N_7796,N_7171,N_7464);
nor U7797 (N_7797,N_6865,N_6805);
nand U7798 (N_7798,N_7321,N_7402);
nand U7799 (N_7799,N_6988,N_7421);
nand U7800 (N_7800,N_6836,N_7266);
nor U7801 (N_7801,N_6808,N_6820);
nor U7802 (N_7802,N_7427,N_6901);
xnor U7803 (N_7803,N_6966,N_7493);
nor U7804 (N_7804,N_7236,N_7338);
nor U7805 (N_7805,N_7483,N_6804);
nor U7806 (N_7806,N_7235,N_6832);
or U7807 (N_7807,N_6968,N_7433);
or U7808 (N_7808,N_7173,N_7317);
nand U7809 (N_7809,N_6815,N_7065);
nor U7810 (N_7810,N_7075,N_7144);
and U7811 (N_7811,N_7223,N_6783);
nor U7812 (N_7812,N_7040,N_7392);
or U7813 (N_7813,N_7005,N_7182);
and U7814 (N_7814,N_6858,N_7263);
or U7815 (N_7815,N_7243,N_7365);
nand U7816 (N_7816,N_7495,N_6976);
and U7817 (N_7817,N_7159,N_6795);
and U7818 (N_7818,N_7210,N_7118);
xnor U7819 (N_7819,N_6791,N_7157);
and U7820 (N_7820,N_6821,N_7344);
xor U7821 (N_7821,N_6959,N_7186);
or U7822 (N_7822,N_7327,N_7050);
or U7823 (N_7823,N_6990,N_7150);
nor U7824 (N_7824,N_6913,N_7445);
nand U7825 (N_7825,N_7368,N_7494);
xnor U7826 (N_7826,N_7244,N_7110);
xor U7827 (N_7827,N_7002,N_7418);
xnor U7828 (N_7828,N_7041,N_7141);
or U7829 (N_7829,N_6764,N_7255);
xor U7830 (N_7830,N_6872,N_6893);
or U7831 (N_7831,N_6927,N_6947);
and U7832 (N_7832,N_7485,N_6828);
xor U7833 (N_7833,N_6789,N_6908);
xor U7834 (N_7834,N_7251,N_7190);
nor U7835 (N_7835,N_7115,N_7074);
xor U7836 (N_7836,N_6853,N_7264);
and U7837 (N_7837,N_6884,N_7189);
nor U7838 (N_7838,N_7276,N_7011);
xor U7839 (N_7839,N_6752,N_6857);
nor U7840 (N_7840,N_7149,N_7015);
nand U7841 (N_7841,N_7030,N_6914);
xnor U7842 (N_7842,N_7143,N_7356);
xor U7843 (N_7843,N_7334,N_7367);
and U7844 (N_7844,N_6782,N_6756);
and U7845 (N_7845,N_7303,N_7101);
nand U7846 (N_7846,N_7265,N_7391);
xnor U7847 (N_7847,N_7214,N_7438);
or U7848 (N_7848,N_7318,N_7099);
xor U7849 (N_7849,N_7134,N_7046);
nor U7850 (N_7850,N_7013,N_7291);
and U7851 (N_7851,N_7394,N_7237);
nor U7852 (N_7852,N_6879,N_6761);
nor U7853 (N_7853,N_7346,N_7478);
and U7854 (N_7854,N_7216,N_7491);
or U7855 (N_7855,N_7474,N_6837);
xor U7856 (N_7856,N_6952,N_7080);
nand U7857 (N_7857,N_7422,N_7328);
xor U7858 (N_7858,N_7388,N_6918);
and U7859 (N_7859,N_7132,N_6775);
and U7860 (N_7860,N_6862,N_7357);
xor U7861 (N_7861,N_6949,N_7000);
xnor U7862 (N_7862,N_6930,N_6903);
nand U7863 (N_7863,N_6762,N_6994);
nor U7864 (N_7864,N_6891,N_7319);
or U7865 (N_7865,N_6933,N_7047);
xor U7866 (N_7866,N_7166,N_7033);
nor U7867 (N_7867,N_7038,N_6969);
xnor U7868 (N_7868,N_7093,N_7231);
and U7869 (N_7869,N_6766,N_7293);
xnor U7870 (N_7870,N_7452,N_6809);
nand U7871 (N_7871,N_7008,N_7298);
and U7872 (N_7872,N_7272,N_7152);
nor U7873 (N_7873,N_6800,N_7068);
nand U7874 (N_7874,N_7201,N_7097);
xor U7875 (N_7875,N_7122,N_7050);
or U7876 (N_7876,N_7054,N_7285);
nor U7877 (N_7877,N_6832,N_6792);
nand U7878 (N_7878,N_7071,N_6949);
nand U7879 (N_7879,N_7230,N_7114);
and U7880 (N_7880,N_7444,N_7463);
xor U7881 (N_7881,N_6836,N_7172);
nor U7882 (N_7882,N_7125,N_7472);
and U7883 (N_7883,N_7323,N_7336);
xor U7884 (N_7884,N_7451,N_7494);
and U7885 (N_7885,N_7278,N_7188);
and U7886 (N_7886,N_6796,N_7372);
nand U7887 (N_7887,N_6943,N_6750);
nand U7888 (N_7888,N_7302,N_6829);
or U7889 (N_7889,N_7435,N_7329);
nor U7890 (N_7890,N_6786,N_6837);
or U7891 (N_7891,N_6822,N_6879);
and U7892 (N_7892,N_7481,N_7045);
xnor U7893 (N_7893,N_7236,N_6920);
and U7894 (N_7894,N_7222,N_7188);
nor U7895 (N_7895,N_6995,N_6986);
nand U7896 (N_7896,N_7197,N_7046);
nand U7897 (N_7897,N_7173,N_6752);
nand U7898 (N_7898,N_6779,N_7354);
xnor U7899 (N_7899,N_7171,N_7136);
nor U7900 (N_7900,N_7445,N_7478);
nor U7901 (N_7901,N_7313,N_6999);
or U7902 (N_7902,N_6763,N_7189);
xor U7903 (N_7903,N_7000,N_7020);
and U7904 (N_7904,N_7406,N_6887);
nor U7905 (N_7905,N_6962,N_6931);
nand U7906 (N_7906,N_7120,N_7349);
xor U7907 (N_7907,N_7195,N_6975);
nand U7908 (N_7908,N_6819,N_6944);
nand U7909 (N_7909,N_7207,N_7138);
or U7910 (N_7910,N_7375,N_7339);
and U7911 (N_7911,N_7063,N_7467);
xor U7912 (N_7912,N_7226,N_7225);
nand U7913 (N_7913,N_7253,N_7064);
xor U7914 (N_7914,N_7257,N_6987);
nor U7915 (N_7915,N_7257,N_6848);
nor U7916 (N_7916,N_7341,N_7210);
nand U7917 (N_7917,N_6796,N_6828);
xor U7918 (N_7918,N_7388,N_7035);
nand U7919 (N_7919,N_6960,N_7446);
xnor U7920 (N_7920,N_7415,N_7402);
and U7921 (N_7921,N_7060,N_7039);
xnor U7922 (N_7922,N_7411,N_7408);
xnor U7923 (N_7923,N_6925,N_7428);
nand U7924 (N_7924,N_7005,N_7091);
and U7925 (N_7925,N_6884,N_6919);
and U7926 (N_7926,N_6926,N_6788);
or U7927 (N_7927,N_7412,N_6822);
and U7928 (N_7928,N_7302,N_6876);
xor U7929 (N_7929,N_7400,N_7189);
nand U7930 (N_7930,N_7210,N_6979);
or U7931 (N_7931,N_7439,N_7420);
nand U7932 (N_7932,N_7412,N_7383);
nand U7933 (N_7933,N_6956,N_6779);
or U7934 (N_7934,N_7446,N_7476);
nor U7935 (N_7935,N_7321,N_6988);
nand U7936 (N_7936,N_7364,N_7408);
xor U7937 (N_7937,N_7445,N_6987);
and U7938 (N_7938,N_7246,N_7334);
or U7939 (N_7939,N_7309,N_7140);
nand U7940 (N_7940,N_6980,N_6983);
nor U7941 (N_7941,N_7228,N_7078);
nor U7942 (N_7942,N_7421,N_7495);
or U7943 (N_7943,N_6812,N_6904);
and U7944 (N_7944,N_7310,N_7399);
xor U7945 (N_7945,N_6777,N_6999);
nor U7946 (N_7946,N_7111,N_7421);
xor U7947 (N_7947,N_7253,N_7277);
nand U7948 (N_7948,N_7348,N_7089);
or U7949 (N_7949,N_7142,N_7180);
or U7950 (N_7950,N_7258,N_7152);
xor U7951 (N_7951,N_7455,N_7453);
or U7952 (N_7952,N_7024,N_6987);
and U7953 (N_7953,N_6797,N_7038);
or U7954 (N_7954,N_6908,N_7359);
xor U7955 (N_7955,N_6794,N_6814);
nand U7956 (N_7956,N_7211,N_7307);
xor U7957 (N_7957,N_7075,N_7091);
or U7958 (N_7958,N_6799,N_7169);
and U7959 (N_7959,N_7025,N_7131);
or U7960 (N_7960,N_7439,N_7328);
nand U7961 (N_7961,N_6831,N_7150);
and U7962 (N_7962,N_6769,N_7035);
and U7963 (N_7963,N_6936,N_6861);
xnor U7964 (N_7964,N_7125,N_6984);
xnor U7965 (N_7965,N_6977,N_6755);
and U7966 (N_7966,N_7466,N_6998);
or U7967 (N_7967,N_6851,N_7185);
or U7968 (N_7968,N_6769,N_7276);
nand U7969 (N_7969,N_7304,N_7051);
or U7970 (N_7970,N_7117,N_7104);
nand U7971 (N_7971,N_6812,N_7074);
nand U7972 (N_7972,N_6775,N_6859);
nand U7973 (N_7973,N_7396,N_6798);
or U7974 (N_7974,N_6750,N_7320);
or U7975 (N_7975,N_7346,N_6766);
and U7976 (N_7976,N_6996,N_6932);
nand U7977 (N_7977,N_6924,N_7034);
nand U7978 (N_7978,N_7298,N_6800);
xnor U7979 (N_7979,N_6944,N_7044);
xor U7980 (N_7980,N_7389,N_7235);
nor U7981 (N_7981,N_6979,N_6805);
nand U7982 (N_7982,N_7101,N_6915);
or U7983 (N_7983,N_7325,N_7401);
nor U7984 (N_7984,N_7177,N_7324);
or U7985 (N_7985,N_6943,N_7238);
or U7986 (N_7986,N_7443,N_7463);
and U7987 (N_7987,N_7437,N_7120);
xnor U7988 (N_7988,N_7164,N_7415);
nand U7989 (N_7989,N_6966,N_7161);
nor U7990 (N_7990,N_7461,N_7480);
nand U7991 (N_7991,N_7393,N_6897);
and U7992 (N_7992,N_7324,N_7063);
and U7993 (N_7993,N_7340,N_7226);
nor U7994 (N_7994,N_7406,N_7357);
nor U7995 (N_7995,N_6766,N_6798);
or U7996 (N_7996,N_7437,N_7191);
nand U7997 (N_7997,N_7408,N_7297);
and U7998 (N_7998,N_7037,N_7012);
and U7999 (N_7999,N_7235,N_6853);
or U8000 (N_8000,N_7008,N_7131);
nor U8001 (N_8001,N_7409,N_6928);
nor U8002 (N_8002,N_7434,N_6844);
or U8003 (N_8003,N_7468,N_6839);
nor U8004 (N_8004,N_6847,N_7238);
xor U8005 (N_8005,N_7203,N_7307);
nand U8006 (N_8006,N_7031,N_6981);
and U8007 (N_8007,N_6978,N_6848);
or U8008 (N_8008,N_7152,N_7234);
or U8009 (N_8009,N_7267,N_6764);
and U8010 (N_8010,N_7019,N_7291);
and U8011 (N_8011,N_7388,N_7366);
nand U8012 (N_8012,N_7312,N_6779);
nand U8013 (N_8013,N_7261,N_7062);
or U8014 (N_8014,N_7240,N_6901);
xor U8015 (N_8015,N_7302,N_7163);
and U8016 (N_8016,N_7194,N_7447);
nor U8017 (N_8017,N_7084,N_7400);
or U8018 (N_8018,N_6807,N_7020);
and U8019 (N_8019,N_7378,N_6898);
nand U8020 (N_8020,N_7042,N_7290);
xor U8021 (N_8021,N_7007,N_7266);
and U8022 (N_8022,N_7356,N_6813);
xor U8023 (N_8023,N_6865,N_7355);
nand U8024 (N_8024,N_7055,N_6979);
nand U8025 (N_8025,N_6900,N_7243);
nand U8026 (N_8026,N_7298,N_6824);
and U8027 (N_8027,N_7290,N_6836);
nand U8028 (N_8028,N_7026,N_7104);
xor U8029 (N_8029,N_7404,N_7198);
or U8030 (N_8030,N_7410,N_7451);
xnor U8031 (N_8031,N_7057,N_6818);
or U8032 (N_8032,N_6758,N_7396);
nand U8033 (N_8033,N_7410,N_7372);
nor U8034 (N_8034,N_7191,N_7424);
nor U8035 (N_8035,N_7161,N_7445);
xor U8036 (N_8036,N_6917,N_7374);
nand U8037 (N_8037,N_6932,N_6869);
nand U8038 (N_8038,N_7403,N_7339);
nor U8039 (N_8039,N_7006,N_7101);
or U8040 (N_8040,N_7332,N_7117);
or U8041 (N_8041,N_7275,N_7364);
nand U8042 (N_8042,N_6924,N_6775);
nand U8043 (N_8043,N_7065,N_7258);
xnor U8044 (N_8044,N_6809,N_7093);
nand U8045 (N_8045,N_7439,N_6918);
and U8046 (N_8046,N_7194,N_7123);
xor U8047 (N_8047,N_7310,N_7357);
and U8048 (N_8048,N_7073,N_7176);
and U8049 (N_8049,N_7491,N_6860);
or U8050 (N_8050,N_6819,N_7475);
nor U8051 (N_8051,N_7012,N_7296);
xnor U8052 (N_8052,N_7423,N_7343);
and U8053 (N_8053,N_7494,N_6900);
nor U8054 (N_8054,N_6841,N_7163);
nor U8055 (N_8055,N_7152,N_7303);
nand U8056 (N_8056,N_7441,N_6809);
nand U8057 (N_8057,N_7462,N_6756);
xor U8058 (N_8058,N_6993,N_7369);
or U8059 (N_8059,N_7070,N_7371);
nor U8060 (N_8060,N_6899,N_6841);
nor U8061 (N_8061,N_7235,N_6924);
and U8062 (N_8062,N_7309,N_6998);
or U8063 (N_8063,N_7408,N_7392);
xnor U8064 (N_8064,N_7266,N_6831);
nor U8065 (N_8065,N_7328,N_6991);
nand U8066 (N_8066,N_6774,N_7382);
nand U8067 (N_8067,N_7373,N_7265);
or U8068 (N_8068,N_6780,N_6758);
nand U8069 (N_8069,N_7465,N_6812);
xnor U8070 (N_8070,N_7480,N_6961);
nor U8071 (N_8071,N_6901,N_7277);
nand U8072 (N_8072,N_7169,N_7085);
or U8073 (N_8073,N_6844,N_6787);
nand U8074 (N_8074,N_7337,N_6798);
or U8075 (N_8075,N_7486,N_6850);
nand U8076 (N_8076,N_6822,N_6808);
xnor U8077 (N_8077,N_7336,N_6976);
nand U8078 (N_8078,N_7476,N_7452);
and U8079 (N_8079,N_7383,N_7355);
or U8080 (N_8080,N_7382,N_7063);
nor U8081 (N_8081,N_7352,N_7467);
nand U8082 (N_8082,N_6880,N_6910);
and U8083 (N_8083,N_6876,N_7103);
xor U8084 (N_8084,N_7328,N_7004);
and U8085 (N_8085,N_7155,N_6887);
and U8086 (N_8086,N_7424,N_6988);
nand U8087 (N_8087,N_7418,N_7097);
and U8088 (N_8088,N_6996,N_6941);
or U8089 (N_8089,N_7123,N_6759);
or U8090 (N_8090,N_7240,N_7231);
nand U8091 (N_8091,N_7020,N_7329);
and U8092 (N_8092,N_7098,N_7494);
and U8093 (N_8093,N_6772,N_6924);
or U8094 (N_8094,N_6962,N_7243);
and U8095 (N_8095,N_6889,N_7021);
or U8096 (N_8096,N_7246,N_7064);
nor U8097 (N_8097,N_7453,N_6817);
nor U8098 (N_8098,N_7268,N_7265);
nand U8099 (N_8099,N_6767,N_7247);
nor U8100 (N_8100,N_6932,N_6898);
and U8101 (N_8101,N_6780,N_7283);
nand U8102 (N_8102,N_7461,N_7457);
nand U8103 (N_8103,N_7490,N_6815);
nor U8104 (N_8104,N_6882,N_7250);
nor U8105 (N_8105,N_7272,N_7396);
and U8106 (N_8106,N_7244,N_6832);
and U8107 (N_8107,N_6929,N_7117);
xnor U8108 (N_8108,N_7456,N_7354);
nor U8109 (N_8109,N_6958,N_6825);
or U8110 (N_8110,N_7459,N_7117);
nor U8111 (N_8111,N_7448,N_6843);
nor U8112 (N_8112,N_7448,N_6874);
xnor U8113 (N_8113,N_7193,N_7369);
nand U8114 (N_8114,N_6963,N_7357);
xnor U8115 (N_8115,N_7291,N_7389);
nand U8116 (N_8116,N_6825,N_7292);
xnor U8117 (N_8117,N_6977,N_7441);
and U8118 (N_8118,N_7253,N_7406);
nor U8119 (N_8119,N_6777,N_6782);
nor U8120 (N_8120,N_7143,N_7301);
nand U8121 (N_8121,N_7175,N_7415);
nand U8122 (N_8122,N_6929,N_6807);
nand U8123 (N_8123,N_7068,N_7003);
nor U8124 (N_8124,N_7255,N_7223);
nand U8125 (N_8125,N_7470,N_6851);
nor U8126 (N_8126,N_7179,N_6960);
nor U8127 (N_8127,N_7183,N_7228);
xor U8128 (N_8128,N_7161,N_7322);
xor U8129 (N_8129,N_7449,N_6912);
nor U8130 (N_8130,N_6959,N_7283);
nand U8131 (N_8131,N_7238,N_7000);
xor U8132 (N_8132,N_6783,N_6801);
and U8133 (N_8133,N_6917,N_7468);
nor U8134 (N_8134,N_7311,N_7050);
xor U8135 (N_8135,N_6767,N_7353);
and U8136 (N_8136,N_7270,N_7108);
nand U8137 (N_8137,N_7065,N_7412);
or U8138 (N_8138,N_7416,N_6909);
xor U8139 (N_8139,N_7419,N_7336);
nor U8140 (N_8140,N_7069,N_6930);
or U8141 (N_8141,N_7011,N_7153);
and U8142 (N_8142,N_7131,N_7403);
xnor U8143 (N_8143,N_7487,N_6765);
nand U8144 (N_8144,N_6864,N_7096);
nor U8145 (N_8145,N_6887,N_6778);
xor U8146 (N_8146,N_7497,N_6878);
nor U8147 (N_8147,N_7257,N_6857);
nand U8148 (N_8148,N_7372,N_7275);
xor U8149 (N_8149,N_6887,N_7145);
and U8150 (N_8150,N_7385,N_6918);
nor U8151 (N_8151,N_7244,N_7151);
nor U8152 (N_8152,N_6822,N_7162);
and U8153 (N_8153,N_7193,N_7008);
or U8154 (N_8154,N_7176,N_7449);
nand U8155 (N_8155,N_6809,N_6812);
xor U8156 (N_8156,N_7161,N_6965);
or U8157 (N_8157,N_6951,N_6815);
and U8158 (N_8158,N_6770,N_6806);
xnor U8159 (N_8159,N_7382,N_7291);
nor U8160 (N_8160,N_7135,N_7339);
nor U8161 (N_8161,N_6988,N_7118);
xor U8162 (N_8162,N_7228,N_6773);
and U8163 (N_8163,N_6896,N_7171);
and U8164 (N_8164,N_7247,N_7218);
nand U8165 (N_8165,N_6857,N_7247);
nand U8166 (N_8166,N_6805,N_6961);
nor U8167 (N_8167,N_7061,N_7135);
nor U8168 (N_8168,N_7058,N_6837);
xnor U8169 (N_8169,N_7029,N_7070);
or U8170 (N_8170,N_7177,N_7090);
and U8171 (N_8171,N_6863,N_7168);
nor U8172 (N_8172,N_7180,N_7378);
or U8173 (N_8173,N_7299,N_7006);
nand U8174 (N_8174,N_7142,N_7012);
and U8175 (N_8175,N_7466,N_6789);
nand U8176 (N_8176,N_7200,N_7027);
or U8177 (N_8177,N_7214,N_6796);
xor U8178 (N_8178,N_7171,N_7046);
xnor U8179 (N_8179,N_7189,N_7148);
nor U8180 (N_8180,N_6826,N_6936);
nand U8181 (N_8181,N_6834,N_7247);
nor U8182 (N_8182,N_6810,N_7162);
nand U8183 (N_8183,N_7094,N_7307);
and U8184 (N_8184,N_7042,N_7048);
xnor U8185 (N_8185,N_7442,N_7059);
or U8186 (N_8186,N_7249,N_6847);
xor U8187 (N_8187,N_7424,N_7202);
nor U8188 (N_8188,N_6958,N_6764);
or U8189 (N_8189,N_7352,N_7161);
nand U8190 (N_8190,N_7345,N_7406);
xor U8191 (N_8191,N_7219,N_7050);
xor U8192 (N_8192,N_7140,N_6858);
xnor U8193 (N_8193,N_7130,N_7484);
and U8194 (N_8194,N_7180,N_6937);
and U8195 (N_8195,N_7422,N_7400);
nor U8196 (N_8196,N_7160,N_7148);
nor U8197 (N_8197,N_7292,N_7065);
nor U8198 (N_8198,N_6888,N_7118);
nor U8199 (N_8199,N_7215,N_6908);
and U8200 (N_8200,N_7423,N_7452);
or U8201 (N_8201,N_7137,N_7485);
xnor U8202 (N_8202,N_6818,N_6752);
xnor U8203 (N_8203,N_7172,N_7059);
nor U8204 (N_8204,N_7308,N_7003);
or U8205 (N_8205,N_7466,N_7267);
nor U8206 (N_8206,N_7217,N_7349);
nand U8207 (N_8207,N_6855,N_7059);
nor U8208 (N_8208,N_6962,N_7132);
xor U8209 (N_8209,N_7207,N_7250);
or U8210 (N_8210,N_6752,N_7316);
nand U8211 (N_8211,N_7055,N_6881);
xor U8212 (N_8212,N_6804,N_6803);
nor U8213 (N_8213,N_7257,N_7316);
nand U8214 (N_8214,N_6753,N_7321);
and U8215 (N_8215,N_7358,N_7164);
xor U8216 (N_8216,N_7263,N_7133);
or U8217 (N_8217,N_7263,N_7368);
nor U8218 (N_8218,N_7334,N_7312);
xor U8219 (N_8219,N_7406,N_7279);
and U8220 (N_8220,N_6911,N_6765);
nor U8221 (N_8221,N_7104,N_6979);
nor U8222 (N_8222,N_7077,N_7044);
nor U8223 (N_8223,N_6816,N_6996);
nor U8224 (N_8224,N_7016,N_7030);
and U8225 (N_8225,N_7434,N_7233);
nor U8226 (N_8226,N_7392,N_7234);
nand U8227 (N_8227,N_6977,N_7113);
or U8228 (N_8228,N_7063,N_7094);
nor U8229 (N_8229,N_7170,N_6759);
xnor U8230 (N_8230,N_7243,N_7007);
xor U8231 (N_8231,N_7284,N_7283);
nor U8232 (N_8232,N_6839,N_6823);
nor U8233 (N_8233,N_7400,N_6824);
nor U8234 (N_8234,N_7361,N_7339);
nor U8235 (N_8235,N_7022,N_7383);
xnor U8236 (N_8236,N_7306,N_7295);
xnor U8237 (N_8237,N_7049,N_6769);
nand U8238 (N_8238,N_7159,N_7007);
or U8239 (N_8239,N_6854,N_7227);
nand U8240 (N_8240,N_6857,N_7440);
nor U8241 (N_8241,N_7090,N_6845);
nand U8242 (N_8242,N_6906,N_6896);
or U8243 (N_8243,N_6790,N_7448);
xor U8244 (N_8244,N_6976,N_6927);
nand U8245 (N_8245,N_7021,N_6950);
and U8246 (N_8246,N_7294,N_6823);
and U8247 (N_8247,N_7259,N_6831);
and U8248 (N_8248,N_7255,N_7443);
and U8249 (N_8249,N_7485,N_7072);
and U8250 (N_8250,N_7508,N_7974);
and U8251 (N_8251,N_7761,N_7836);
and U8252 (N_8252,N_7783,N_7785);
nand U8253 (N_8253,N_8228,N_8179);
or U8254 (N_8254,N_7883,N_7533);
and U8255 (N_8255,N_7848,N_8238);
or U8256 (N_8256,N_8033,N_8208);
or U8257 (N_8257,N_7946,N_7617);
nand U8258 (N_8258,N_8230,N_8027);
xor U8259 (N_8259,N_7561,N_7939);
nand U8260 (N_8260,N_7959,N_8087);
nand U8261 (N_8261,N_7621,N_7715);
or U8262 (N_8262,N_7515,N_7880);
and U8263 (N_8263,N_8173,N_7638);
or U8264 (N_8264,N_8206,N_7519);
and U8265 (N_8265,N_7657,N_7948);
nor U8266 (N_8266,N_8118,N_8211);
nor U8267 (N_8267,N_7655,N_8141);
nor U8268 (N_8268,N_7516,N_7881);
nand U8269 (N_8269,N_7817,N_7906);
nand U8270 (N_8270,N_8219,N_7693);
nor U8271 (N_8271,N_8067,N_7899);
nor U8272 (N_8272,N_7903,N_7828);
xor U8273 (N_8273,N_7654,N_7667);
and U8274 (N_8274,N_7694,N_8048);
and U8275 (N_8275,N_8061,N_7915);
and U8276 (N_8276,N_7733,N_7989);
or U8277 (N_8277,N_7819,N_7581);
nor U8278 (N_8278,N_8006,N_7537);
xnor U8279 (N_8279,N_8201,N_7843);
xnor U8280 (N_8280,N_7996,N_8234);
nor U8281 (N_8281,N_7649,N_7646);
nand U8282 (N_8282,N_7928,N_7824);
and U8283 (N_8283,N_7614,N_8247);
nor U8284 (N_8284,N_8042,N_7917);
xnor U8285 (N_8285,N_7586,N_8196);
or U8286 (N_8286,N_7618,N_8032);
nand U8287 (N_8287,N_7751,N_7665);
or U8288 (N_8288,N_8138,N_7671);
and U8289 (N_8289,N_8223,N_7567);
xor U8290 (N_8290,N_8175,N_8147);
nor U8291 (N_8291,N_7668,N_8210);
nand U8292 (N_8292,N_8186,N_7776);
nand U8293 (N_8293,N_7669,N_7965);
nor U8294 (N_8294,N_7935,N_7549);
nor U8295 (N_8295,N_7923,N_7644);
nand U8296 (N_8296,N_7936,N_7979);
nand U8297 (N_8297,N_8106,N_8174);
and U8298 (N_8298,N_8188,N_7932);
nor U8299 (N_8299,N_7707,N_8189);
or U8300 (N_8300,N_8248,N_7977);
or U8301 (N_8301,N_7882,N_8080);
nor U8302 (N_8302,N_7938,N_7569);
nor U8303 (N_8303,N_7681,N_8181);
nor U8304 (N_8304,N_8028,N_7971);
and U8305 (N_8305,N_7951,N_7744);
xnor U8306 (N_8306,N_7502,N_7731);
xor U8307 (N_8307,N_7564,N_7759);
and U8308 (N_8308,N_8158,N_8246);
xnor U8309 (N_8309,N_7818,N_7807);
nor U8310 (N_8310,N_7509,N_8058);
or U8311 (N_8311,N_7978,N_8005);
xnor U8312 (N_8312,N_8224,N_7683);
xnor U8313 (N_8313,N_7827,N_7894);
nand U8314 (N_8314,N_8109,N_7780);
or U8315 (N_8315,N_7754,N_8003);
nand U8316 (N_8316,N_7760,N_7659);
nand U8317 (N_8317,N_7722,N_7726);
xor U8318 (N_8318,N_7793,N_8145);
nand U8319 (N_8319,N_8207,N_7987);
and U8320 (N_8320,N_8095,N_8114);
or U8321 (N_8321,N_7504,N_8045);
nand U8322 (N_8322,N_7629,N_8001);
and U8323 (N_8323,N_7992,N_7563);
and U8324 (N_8324,N_8044,N_7800);
and U8325 (N_8325,N_7732,N_8220);
nor U8326 (N_8326,N_7719,N_7872);
nor U8327 (N_8327,N_7797,N_7985);
or U8328 (N_8328,N_8165,N_8123);
xnor U8329 (N_8329,N_7541,N_7764);
or U8330 (N_8330,N_8101,N_8197);
or U8331 (N_8331,N_7503,N_7723);
or U8332 (N_8332,N_7565,N_7597);
and U8333 (N_8333,N_8057,N_8012);
or U8334 (N_8334,N_7860,N_7506);
nand U8335 (N_8335,N_8046,N_7670);
xnor U8336 (N_8336,N_7559,N_7749);
nor U8337 (N_8337,N_7686,N_8113);
or U8338 (N_8338,N_8093,N_7542);
or U8339 (N_8339,N_8090,N_7838);
and U8340 (N_8340,N_7769,N_7768);
nor U8341 (N_8341,N_7582,N_7627);
and U8342 (N_8342,N_8161,N_7613);
and U8343 (N_8343,N_8103,N_8085);
or U8344 (N_8344,N_7725,N_7543);
nor U8345 (N_8345,N_7823,N_7709);
xnor U8346 (N_8346,N_7610,N_8190);
nand U8347 (N_8347,N_8217,N_7849);
and U8348 (N_8348,N_7960,N_8236);
nand U8349 (N_8349,N_8185,N_7804);
nor U8350 (N_8350,N_7792,N_7990);
nand U8351 (N_8351,N_8037,N_7538);
nand U8352 (N_8352,N_8098,N_8008);
nor U8353 (N_8353,N_7689,N_8198);
xnor U8354 (N_8354,N_8105,N_7900);
nor U8355 (N_8355,N_7787,N_7607);
nand U8356 (N_8356,N_7856,N_7677);
xor U8357 (N_8357,N_7868,N_7850);
and U8358 (N_8358,N_7645,N_7877);
or U8359 (N_8359,N_8142,N_8064);
nand U8360 (N_8360,N_7835,N_8117);
nor U8361 (N_8361,N_7967,N_8083);
xnor U8362 (N_8362,N_8209,N_7808);
xnor U8363 (N_8363,N_7550,N_8014);
nand U8364 (N_8364,N_7893,N_7993);
or U8365 (N_8365,N_8244,N_8134);
nand U8366 (N_8366,N_7791,N_7529);
or U8367 (N_8367,N_8052,N_7957);
xnor U8368 (N_8368,N_7658,N_8170);
and U8369 (N_8369,N_7642,N_8034);
or U8370 (N_8370,N_7548,N_7592);
or U8371 (N_8371,N_8054,N_8183);
xor U8372 (N_8372,N_7921,N_7598);
and U8373 (N_8373,N_7690,N_7570);
nor U8374 (N_8374,N_8022,N_8212);
xnor U8375 (N_8375,N_7595,N_7666);
or U8376 (N_8376,N_7579,N_8168);
xor U8377 (N_8377,N_7984,N_7576);
nand U8378 (N_8378,N_7773,N_7520);
xor U8379 (N_8379,N_7624,N_7892);
nor U8380 (N_8380,N_8026,N_7784);
xor U8381 (N_8381,N_7730,N_8041);
and U8382 (N_8382,N_8245,N_7535);
or U8383 (N_8383,N_8097,N_7842);
nand U8384 (N_8384,N_8116,N_8227);
nand U8385 (N_8385,N_7994,N_7738);
and U8386 (N_8386,N_7640,N_7574);
and U8387 (N_8387,N_7748,N_7982);
nor U8388 (N_8388,N_8144,N_7981);
and U8389 (N_8389,N_7897,N_8136);
or U8390 (N_8390,N_7745,N_7552);
or U8391 (N_8391,N_7736,N_7844);
nor U8392 (N_8392,N_7675,N_7772);
and U8393 (N_8393,N_7558,N_7997);
nand U8394 (N_8394,N_7571,N_7933);
and U8395 (N_8395,N_8191,N_8121);
xnor U8396 (N_8396,N_7786,N_7710);
or U8397 (N_8397,N_7594,N_7554);
nor U8398 (N_8398,N_7988,N_7770);
nand U8399 (N_8399,N_8180,N_7553);
and U8400 (N_8400,N_8050,N_7833);
nor U8401 (N_8401,N_7672,N_7902);
or U8402 (N_8402,N_8009,N_7854);
xnor U8403 (N_8403,N_8192,N_8040);
and U8404 (N_8404,N_7852,N_7810);
and U8405 (N_8405,N_8135,N_8091);
and U8406 (N_8406,N_8204,N_7820);
or U8407 (N_8407,N_7815,N_7578);
and U8408 (N_8408,N_7956,N_7661);
nor U8409 (N_8409,N_7700,N_7812);
nand U8410 (N_8410,N_7679,N_7740);
nor U8411 (N_8411,N_8088,N_8108);
or U8412 (N_8412,N_7806,N_7622);
and U8413 (N_8413,N_7507,N_8218);
nand U8414 (N_8414,N_8214,N_7846);
nand U8415 (N_8415,N_7568,N_8063);
nand U8416 (N_8416,N_7931,N_8225);
and U8417 (N_8417,N_7954,N_7602);
xor U8418 (N_8418,N_8081,N_7511);
xnor U8419 (N_8419,N_7596,N_8065);
and U8420 (N_8420,N_8021,N_7631);
xor U8421 (N_8421,N_8184,N_7980);
or U8422 (N_8422,N_8166,N_7910);
nor U8423 (N_8423,N_7763,N_7692);
nand U8424 (N_8424,N_7912,N_8049);
or U8425 (N_8425,N_7867,N_7650);
and U8426 (N_8426,N_8079,N_7717);
nor U8427 (N_8427,N_8129,N_7703);
nand U8428 (N_8428,N_8231,N_7523);
or U8429 (N_8429,N_8082,N_7606);
nand U8430 (N_8430,N_7905,N_7896);
nand U8431 (N_8431,N_7826,N_7593);
and U8432 (N_8432,N_7626,N_7590);
or U8433 (N_8433,N_8243,N_7705);
xnor U8434 (N_8434,N_7534,N_7952);
nand U8435 (N_8435,N_7968,N_8120);
or U8436 (N_8436,N_7545,N_7623);
nand U8437 (N_8437,N_7628,N_8237);
nor U8438 (N_8438,N_7584,N_7876);
nand U8439 (N_8439,N_8007,N_8107);
xnor U8440 (N_8440,N_8023,N_7866);
and U8441 (N_8441,N_7963,N_7521);
and U8442 (N_8442,N_7580,N_8011);
or U8443 (N_8443,N_7781,N_7904);
xnor U8444 (N_8444,N_7857,N_7821);
nor U8445 (N_8445,N_7678,N_7653);
nand U8446 (N_8446,N_7983,N_7630);
and U8447 (N_8447,N_7739,N_7920);
and U8448 (N_8448,N_7612,N_8119);
nand U8449 (N_8449,N_8203,N_8200);
nand U8450 (N_8450,N_8020,N_8235);
and U8451 (N_8451,N_7969,N_8086);
xor U8452 (N_8452,N_7663,N_7619);
nand U8453 (N_8453,N_8039,N_8024);
nand U8454 (N_8454,N_7825,N_7701);
nor U8455 (N_8455,N_8074,N_7914);
nand U8456 (N_8456,N_7795,N_7941);
xor U8457 (N_8457,N_7609,N_8176);
nand U8458 (N_8458,N_8167,N_7636);
nor U8459 (N_8459,N_7831,N_7934);
nor U8460 (N_8460,N_8016,N_7524);
or U8461 (N_8461,N_7927,N_8143);
or U8462 (N_8462,N_7861,N_7970);
nor U8463 (N_8463,N_7855,N_7756);
nand U8464 (N_8464,N_7540,N_7514);
nand U8465 (N_8465,N_7714,N_7652);
nor U8466 (N_8466,N_7890,N_8249);
or U8467 (N_8467,N_7986,N_7958);
nor U8468 (N_8468,N_7688,N_7517);
and U8469 (N_8469,N_7615,N_8099);
xnor U8470 (N_8470,N_7699,N_7685);
xnor U8471 (N_8471,N_7556,N_8100);
nand U8472 (N_8472,N_7794,N_7706);
nor U8473 (N_8473,N_7962,N_8094);
or U8474 (N_8474,N_7746,N_8222);
or U8475 (N_8475,N_8187,N_7922);
nor U8476 (N_8476,N_7955,N_7664);
nor U8477 (N_8477,N_7729,N_7884);
and U8478 (N_8478,N_8071,N_8036);
and U8479 (N_8479,N_8029,N_8193);
or U8480 (N_8480,N_7647,N_8104);
nor U8481 (N_8481,N_7546,N_7888);
nand U8482 (N_8482,N_8110,N_7735);
nor U8483 (N_8483,N_8112,N_7839);
xor U8484 (N_8484,N_7953,N_8127);
nand U8485 (N_8485,N_7874,N_7788);
nor U8486 (N_8486,N_7811,N_7641);
nor U8487 (N_8487,N_8013,N_8051);
nand U8488 (N_8488,N_7803,N_7604);
nand U8489 (N_8489,N_8066,N_7775);
and U8490 (N_8490,N_7837,N_7637);
xor U8491 (N_8491,N_7802,N_8155);
and U8492 (N_8492,N_8139,N_8002);
xor U8493 (N_8493,N_7909,N_8171);
nand U8494 (N_8494,N_7919,N_7587);
xnor U8495 (N_8495,N_7620,N_7878);
nand U8496 (N_8496,N_7964,N_7512);
and U8497 (N_8497,N_8156,N_7782);
or U8498 (N_8498,N_8062,N_7926);
or U8499 (N_8499,N_7975,N_7885);
nand U8500 (N_8500,N_7562,N_7544);
xnor U8501 (N_8501,N_8195,N_8132);
nand U8502 (N_8502,N_7737,N_7711);
and U8503 (N_8503,N_7911,N_7510);
nor U8504 (N_8504,N_7779,N_8015);
nor U8505 (N_8505,N_7680,N_7611);
and U8506 (N_8506,N_7889,N_8150);
nand U8507 (N_8507,N_7901,N_7851);
or U8508 (N_8508,N_8169,N_7757);
and U8509 (N_8509,N_7742,N_7961);
xor U8510 (N_8510,N_8092,N_7913);
nor U8511 (N_8511,N_8163,N_7929);
and U8512 (N_8512,N_7676,N_8075);
nor U8513 (N_8513,N_8233,N_7747);
and U8514 (N_8514,N_7767,N_7765);
xor U8515 (N_8515,N_7639,N_7907);
nor U8516 (N_8516,N_7608,N_7924);
nor U8517 (N_8517,N_7859,N_7616);
nand U8518 (N_8518,N_8000,N_8154);
nand U8519 (N_8519,N_7500,N_7712);
xor U8520 (N_8520,N_7687,N_8072);
or U8521 (N_8521,N_8018,N_7832);
nor U8522 (N_8522,N_7547,N_7530);
or U8523 (N_8523,N_7741,N_8157);
or U8524 (N_8524,N_7822,N_8053);
nor U8525 (N_8525,N_7862,N_8194);
xnor U8526 (N_8526,N_8122,N_7805);
and U8527 (N_8527,N_7589,N_8164);
nor U8528 (N_8528,N_7801,N_8076);
xnor U8529 (N_8529,N_7972,N_7814);
nor U8530 (N_8530,N_7829,N_8226);
and U8531 (N_8531,N_8059,N_7845);
nor U8532 (N_8532,N_7750,N_7518);
and U8533 (N_8533,N_8035,N_7930);
or U8534 (N_8534,N_7648,N_7527);
or U8535 (N_8535,N_7771,N_7696);
nand U8536 (N_8536,N_7684,N_7753);
nand U8537 (N_8537,N_7585,N_8102);
nor U8538 (N_8538,N_8047,N_7743);
xnor U8539 (N_8539,N_8073,N_7566);
or U8540 (N_8540,N_7858,N_7716);
nand U8541 (N_8541,N_8060,N_7945);
nor U8542 (N_8542,N_7682,N_7603);
nand U8543 (N_8543,N_7673,N_8177);
and U8544 (N_8544,N_7755,N_7798);
or U8545 (N_8545,N_7999,N_7691);
nor U8546 (N_8546,N_7789,N_7816);
xnor U8547 (N_8547,N_7643,N_8149);
and U8548 (N_8548,N_7830,N_8078);
and U8549 (N_8549,N_7591,N_7708);
nand U8550 (N_8550,N_7651,N_7790);
and U8551 (N_8551,N_8140,N_7662);
nor U8552 (N_8552,N_8069,N_7976);
or U8553 (N_8553,N_7895,N_7778);
and U8554 (N_8554,N_8124,N_8056);
nand U8555 (N_8555,N_8148,N_7937);
nand U8556 (N_8556,N_7536,N_7875);
nor U8557 (N_8557,N_7601,N_7940);
xor U8558 (N_8558,N_7528,N_7752);
xor U8559 (N_8559,N_7625,N_7522);
or U8560 (N_8560,N_7766,N_7704);
or U8561 (N_8561,N_7871,N_8070);
nand U8562 (N_8562,N_7660,N_8031);
or U8563 (N_8563,N_7724,N_7777);
nor U8564 (N_8564,N_7573,N_7758);
or U8565 (N_8565,N_8159,N_7635);
nor U8566 (N_8566,N_7774,N_8232);
and U8567 (N_8567,N_7588,N_8216);
nor U8568 (N_8568,N_8240,N_7887);
nand U8569 (N_8569,N_7633,N_7555);
and U8570 (N_8570,N_7718,N_7734);
nor U8571 (N_8571,N_8178,N_7605);
nor U8572 (N_8572,N_7583,N_8151);
nand U8573 (N_8573,N_8077,N_7697);
or U8574 (N_8574,N_7600,N_7870);
and U8575 (N_8575,N_8221,N_7728);
or U8576 (N_8576,N_8017,N_8229);
nor U8577 (N_8577,N_7942,N_7656);
or U8578 (N_8578,N_8162,N_7505);
or U8579 (N_8579,N_8130,N_8172);
and U8580 (N_8580,N_8205,N_7865);
or U8581 (N_8581,N_8131,N_8213);
xnor U8582 (N_8582,N_7840,N_7713);
and U8583 (N_8583,N_7575,N_7925);
and U8584 (N_8584,N_7634,N_7947);
nand U8585 (N_8585,N_8126,N_8125);
and U8586 (N_8586,N_8241,N_8128);
or U8587 (N_8587,N_7873,N_8199);
xnor U8588 (N_8588,N_7531,N_7721);
nor U8589 (N_8589,N_7853,N_8146);
or U8590 (N_8590,N_7834,N_7513);
nand U8591 (N_8591,N_7918,N_8239);
nand U8592 (N_8592,N_8084,N_8111);
or U8593 (N_8593,N_8089,N_7632);
or U8594 (N_8594,N_8137,N_7702);
nor U8595 (N_8595,N_7557,N_7501);
and U8596 (N_8596,N_8055,N_8025);
nor U8597 (N_8597,N_7916,N_8160);
xnor U8598 (N_8598,N_8133,N_7526);
xnor U8599 (N_8599,N_8242,N_7525);
or U8600 (N_8600,N_7864,N_7944);
xnor U8601 (N_8601,N_8068,N_7577);
nor U8602 (N_8602,N_7727,N_7891);
and U8603 (N_8603,N_7973,N_7869);
and U8604 (N_8604,N_7799,N_7847);
xnor U8605 (N_8605,N_8202,N_7966);
xor U8606 (N_8606,N_7762,N_7551);
nor U8607 (N_8607,N_7950,N_7991);
nand U8608 (N_8608,N_8010,N_7796);
or U8609 (N_8609,N_7572,N_8152);
and U8610 (N_8610,N_7886,N_7695);
or U8611 (N_8611,N_7943,N_7809);
nand U8612 (N_8612,N_8182,N_8115);
nor U8613 (N_8613,N_8096,N_7949);
nand U8614 (N_8614,N_8153,N_7908);
nor U8615 (N_8615,N_7879,N_8004);
nor U8616 (N_8616,N_7898,N_7998);
xor U8617 (N_8617,N_8043,N_7560);
nor U8618 (N_8618,N_8215,N_7841);
xor U8619 (N_8619,N_7599,N_7995);
nor U8620 (N_8620,N_8038,N_7674);
nor U8621 (N_8621,N_7698,N_7813);
or U8622 (N_8622,N_7863,N_8019);
or U8623 (N_8623,N_7539,N_7532);
xor U8624 (N_8624,N_7720,N_8030);
nor U8625 (N_8625,N_7739,N_7530);
and U8626 (N_8626,N_7619,N_7869);
and U8627 (N_8627,N_7779,N_7856);
nand U8628 (N_8628,N_7743,N_8009);
nor U8629 (N_8629,N_7654,N_8147);
nor U8630 (N_8630,N_7723,N_8033);
nor U8631 (N_8631,N_8213,N_7559);
nand U8632 (N_8632,N_7647,N_7698);
xnor U8633 (N_8633,N_8026,N_7714);
and U8634 (N_8634,N_8018,N_7591);
nand U8635 (N_8635,N_8039,N_7833);
or U8636 (N_8636,N_8135,N_8233);
and U8637 (N_8637,N_7803,N_7590);
or U8638 (N_8638,N_7557,N_8177);
and U8639 (N_8639,N_7881,N_8121);
xnor U8640 (N_8640,N_7816,N_8148);
nand U8641 (N_8641,N_7701,N_8195);
nand U8642 (N_8642,N_8234,N_7773);
xor U8643 (N_8643,N_7798,N_7725);
nor U8644 (N_8644,N_7753,N_8183);
and U8645 (N_8645,N_7644,N_7702);
nand U8646 (N_8646,N_7885,N_7510);
nand U8647 (N_8647,N_8166,N_7575);
and U8648 (N_8648,N_8070,N_7836);
or U8649 (N_8649,N_7564,N_8022);
nor U8650 (N_8650,N_7642,N_7675);
or U8651 (N_8651,N_7986,N_7586);
xor U8652 (N_8652,N_7554,N_8170);
nand U8653 (N_8653,N_7935,N_7529);
and U8654 (N_8654,N_7668,N_7710);
nand U8655 (N_8655,N_8155,N_7638);
nand U8656 (N_8656,N_7960,N_8212);
or U8657 (N_8657,N_8012,N_7724);
xnor U8658 (N_8658,N_7839,N_7686);
or U8659 (N_8659,N_7684,N_8066);
nor U8660 (N_8660,N_7686,N_8234);
nand U8661 (N_8661,N_7938,N_7770);
nand U8662 (N_8662,N_7628,N_8119);
and U8663 (N_8663,N_7568,N_7992);
or U8664 (N_8664,N_8211,N_7706);
nor U8665 (N_8665,N_8024,N_7907);
nand U8666 (N_8666,N_8018,N_7959);
or U8667 (N_8667,N_8014,N_7888);
and U8668 (N_8668,N_7904,N_7750);
nand U8669 (N_8669,N_7540,N_7805);
nor U8670 (N_8670,N_7861,N_8207);
or U8671 (N_8671,N_8173,N_8174);
and U8672 (N_8672,N_7775,N_7725);
nor U8673 (N_8673,N_7945,N_7628);
xnor U8674 (N_8674,N_8076,N_7733);
nor U8675 (N_8675,N_8128,N_8230);
and U8676 (N_8676,N_7937,N_8209);
nor U8677 (N_8677,N_7719,N_7772);
xnor U8678 (N_8678,N_7763,N_7946);
xor U8679 (N_8679,N_7917,N_7957);
nand U8680 (N_8680,N_7689,N_8023);
and U8681 (N_8681,N_7530,N_7706);
or U8682 (N_8682,N_7516,N_7908);
nand U8683 (N_8683,N_7723,N_8101);
or U8684 (N_8684,N_7717,N_7877);
nand U8685 (N_8685,N_7695,N_7506);
nand U8686 (N_8686,N_7786,N_8091);
xnor U8687 (N_8687,N_8068,N_7850);
or U8688 (N_8688,N_7810,N_7780);
nor U8689 (N_8689,N_7925,N_7543);
nor U8690 (N_8690,N_7672,N_7618);
xor U8691 (N_8691,N_8108,N_7732);
nor U8692 (N_8692,N_7853,N_8151);
or U8693 (N_8693,N_8133,N_8122);
or U8694 (N_8694,N_7956,N_7800);
xor U8695 (N_8695,N_8193,N_8018);
nor U8696 (N_8696,N_7679,N_7925);
nor U8697 (N_8697,N_7615,N_8136);
xor U8698 (N_8698,N_7757,N_8211);
and U8699 (N_8699,N_7971,N_7983);
and U8700 (N_8700,N_8148,N_7944);
nor U8701 (N_8701,N_8081,N_8164);
and U8702 (N_8702,N_8097,N_8128);
and U8703 (N_8703,N_7797,N_7689);
xor U8704 (N_8704,N_7587,N_8018);
xnor U8705 (N_8705,N_7680,N_8058);
and U8706 (N_8706,N_7748,N_7777);
nor U8707 (N_8707,N_8218,N_8154);
and U8708 (N_8708,N_7818,N_7825);
xor U8709 (N_8709,N_7855,N_7744);
or U8710 (N_8710,N_7676,N_7922);
and U8711 (N_8711,N_8054,N_7591);
or U8712 (N_8712,N_8011,N_7576);
nor U8713 (N_8713,N_8121,N_8065);
nand U8714 (N_8714,N_8004,N_7996);
nor U8715 (N_8715,N_7571,N_7600);
xor U8716 (N_8716,N_7725,N_7782);
xor U8717 (N_8717,N_7869,N_7992);
nand U8718 (N_8718,N_7935,N_7843);
nand U8719 (N_8719,N_7933,N_7796);
nor U8720 (N_8720,N_7633,N_7818);
nor U8721 (N_8721,N_7963,N_8040);
nand U8722 (N_8722,N_7577,N_7908);
or U8723 (N_8723,N_7923,N_7899);
and U8724 (N_8724,N_8240,N_7959);
or U8725 (N_8725,N_7707,N_7933);
xor U8726 (N_8726,N_7952,N_8116);
nor U8727 (N_8727,N_8221,N_8073);
nand U8728 (N_8728,N_7564,N_8074);
nor U8729 (N_8729,N_7932,N_7960);
or U8730 (N_8730,N_7567,N_7599);
and U8731 (N_8731,N_8009,N_7924);
and U8732 (N_8732,N_8196,N_7616);
nand U8733 (N_8733,N_7997,N_7809);
and U8734 (N_8734,N_7942,N_7969);
nand U8735 (N_8735,N_8170,N_7527);
nand U8736 (N_8736,N_8227,N_7724);
nand U8737 (N_8737,N_7548,N_7754);
or U8738 (N_8738,N_8197,N_7531);
and U8739 (N_8739,N_8010,N_8165);
nand U8740 (N_8740,N_7524,N_7629);
xnor U8741 (N_8741,N_7941,N_7692);
and U8742 (N_8742,N_7985,N_7554);
nor U8743 (N_8743,N_7558,N_8047);
and U8744 (N_8744,N_7643,N_8002);
and U8745 (N_8745,N_7784,N_7990);
or U8746 (N_8746,N_8168,N_8063);
or U8747 (N_8747,N_8091,N_7980);
nor U8748 (N_8748,N_8127,N_8235);
xor U8749 (N_8749,N_7801,N_7813);
and U8750 (N_8750,N_7855,N_8222);
nand U8751 (N_8751,N_7841,N_7608);
xnor U8752 (N_8752,N_8095,N_8089);
xor U8753 (N_8753,N_8180,N_7602);
xnor U8754 (N_8754,N_7791,N_8191);
nor U8755 (N_8755,N_7789,N_8068);
or U8756 (N_8756,N_7683,N_7652);
nor U8757 (N_8757,N_7800,N_7542);
or U8758 (N_8758,N_7773,N_7621);
nand U8759 (N_8759,N_8157,N_7677);
nor U8760 (N_8760,N_7709,N_7699);
xnor U8761 (N_8761,N_7514,N_7904);
and U8762 (N_8762,N_8231,N_7509);
nand U8763 (N_8763,N_8129,N_7770);
nor U8764 (N_8764,N_8128,N_8012);
nand U8765 (N_8765,N_8191,N_7941);
nor U8766 (N_8766,N_7739,N_8157);
nor U8767 (N_8767,N_7606,N_7948);
and U8768 (N_8768,N_7694,N_8057);
nor U8769 (N_8769,N_7540,N_7613);
nor U8770 (N_8770,N_8214,N_7891);
or U8771 (N_8771,N_7974,N_7774);
or U8772 (N_8772,N_7583,N_7811);
or U8773 (N_8773,N_7567,N_8136);
nand U8774 (N_8774,N_7528,N_7903);
xor U8775 (N_8775,N_7890,N_8000);
xnor U8776 (N_8776,N_7578,N_7573);
nand U8777 (N_8777,N_7847,N_8229);
and U8778 (N_8778,N_7583,N_8090);
nand U8779 (N_8779,N_8212,N_7950);
and U8780 (N_8780,N_8134,N_7720);
xor U8781 (N_8781,N_7992,N_8067);
nand U8782 (N_8782,N_7652,N_8204);
and U8783 (N_8783,N_7607,N_7837);
and U8784 (N_8784,N_7751,N_8009);
xor U8785 (N_8785,N_7581,N_7630);
nand U8786 (N_8786,N_8228,N_7735);
or U8787 (N_8787,N_7828,N_7677);
or U8788 (N_8788,N_7511,N_7786);
nand U8789 (N_8789,N_8153,N_7793);
and U8790 (N_8790,N_7581,N_7732);
and U8791 (N_8791,N_8036,N_7716);
or U8792 (N_8792,N_7769,N_7649);
xnor U8793 (N_8793,N_7876,N_7576);
or U8794 (N_8794,N_7917,N_7845);
or U8795 (N_8795,N_7825,N_7634);
xnor U8796 (N_8796,N_8131,N_7887);
or U8797 (N_8797,N_7939,N_7873);
nand U8798 (N_8798,N_7851,N_7675);
xnor U8799 (N_8799,N_7816,N_7951);
or U8800 (N_8800,N_7859,N_8062);
nand U8801 (N_8801,N_7982,N_7910);
nor U8802 (N_8802,N_8179,N_7565);
nor U8803 (N_8803,N_7534,N_8132);
xor U8804 (N_8804,N_7833,N_7613);
xor U8805 (N_8805,N_8193,N_8157);
nor U8806 (N_8806,N_7516,N_8014);
and U8807 (N_8807,N_7530,N_7528);
nor U8808 (N_8808,N_8144,N_7829);
xor U8809 (N_8809,N_7717,N_8046);
and U8810 (N_8810,N_7635,N_8171);
nand U8811 (N_8811,N_8069,N_8030);
nand U8812 (N_8812,N_7796,N_7512);
or U8813 (N_8813,N_7702,N_8025);
nand U8814 (N_8814,N_8197,N_7596);
nand U8815 (N_8815,N_8122,N_8074);
nor U8816 (N_8816,N_7946,N_7914);
nand U8817 (N_8817,N_7537,N_7662);
nand U8818 (N_8818,N_7666,N_7965);
nand U8819 (N_8819,N_7883,N_7973);
nor U8820 (N_8820,N_7540,N_8142);
nand U8821 (N_8821,N_7655,N_7545);
and U8822 (N_8822,N_8227,N_8199);
nor U8823 (N_8823,N_8110,N_7662);
or U8824 (N_8824,N_7765,N_7849);
nand U8825 (N_8825,N_7864,N_8184);
or U8826 (N_8826,N_7610,N_8166);
and U8827 (N_8827,N_7961,N_7819);
nand U8828 (N_8828,N_7608,N_7609);
xor U8829 (N_8829,N_7851,N_8085);
nand U8830 (N_8830,N_7878,N_7858);
xor U8831 (N_8831,N_8192,N_8197);
or U8832 (N_8832,N_7979,N_8231);
or U8833 (N_8833,N_7768,N_7959);
xnor U8834 (N_8834,N_7982,N_7809);
xor U8835 (N_8835,N_8043,N_7899);
nor U8836 (N_8836,N_8163,N_8133);
and U8837 (N_8837,N_7515,N_7892);
xor U8838 (N_8838,N_8219,N_7798);
and U8839 (N_8839,N_8148,N_7873);
xnor U8840 (N_8840,N_7850,N_8202);
and U8841 (N_8841,N_7871,N_8150);
nand U8842 (N_8842,N_7877,N_7765);
xor U8843 (N_8843,N_7896,N_7693);
nand U8844 (N_8844,N_7810,N_7651);
nand U8845 (N_8845,N_7682,N_7997);
or U8846 (N_8846,N_7633,N_7738);
and U8847 (N_8847,N_7868,N_8178);
and U8848 (N_8848,N_8030,N_7537);
nand U8849 (N_8849,N_7749,N_8055);
xnor U8850 (N_8850,N_7865,N_8027);
or U8851 (N_8851,N_7524,N_8099);
and U8852 (N_8852,N_7631,N_7804);
nor U8853 (N_8853,N_7750,N_7951);
nand U8854 (N_8854,N_8218,N_7602);
and U8855 (N_8855,N_7919,N_7581);
or U8856 (N_8856,N_7936,N_8126);
xnor U8857 (N_8857,N_8081,N_7703);
and U8858 (N_8858,N_7574,N_7512);
and U8859 (N_8859,N_7706,N_8023);
and U8860 (N_8860,N_7636,N_7665);
nand U8861 (N_8861,N_7856,N_7831);
nand U8862 (N_8862,N_8197,N_8000);
nand U8863 (N_8863,N_7732,N_8049);
xnor U8864 (N_8864,N_7970,N_7927);
xnor U8865 (N_8865,N_8162,N_7874);
nor U8866 (N_8866,N_7704,N_7705);
or U8867 (N_8867,N_8192,N_7766);
or U8868 (N_8868,N_8087,N_8025);
and U8869 (N_8869,N_7613,N_7953);
nor U8870 (N_8870,N_7921,N_8137);
nand U8871 (N_8871,N_7782,N_7893);
nor U8872 (N_8872,N_7780,N_7773);
or U8873 (N_8873,N_7745,N_7526);
and U8874 (N_8874,N_7625,N_7763);
xor U8875 (N_8875,N_7815,N_7564);
and U8876 (N_8876,N_7583,N_8019);
nor U8877 (N_8877,N_7682,N_7720);
nor U8878 (N_8878,N_7899,N_7945);
nor U8879 (N_8879,N_8071,N_7977);
or U8880 (N_8880,N_7785,N_7510);
xor U8881 (N_8881,N_7994,N_8240);
nand U8882 (N_8882,N_7646,N_7693);
nor U8883 (N_8883,N_7860,N_7625);
xnor U8884 (N_8884,N_8056,N_7846);
or U8885 (N_8885,N_8188,N_8121);
or U8886 (N_8886,N_7821,N_7775);
nor U8887 (N_8887,N_8202,N_7829);
nand U8888 (N_8888,N_8117,N_7722);
or U8889 (N_8889,N_7502,N_7902);
and U8890 (N_8890,N_8048,N_7817);
nand U8891 (N_8891,N_8066,N_8102);
and U8892 (N_8892,N_8149,N_7934);
xor U8893 (N_8893,N_8211,N_7580);
nand U8894 (N_8894,N_8240,N_8071);
nor U8895 (N_8895,N_8128,N_8104);
or U8896 (N_8896,N_8218,N_7684);
nand U8897 (N_8897,N_8106,N_8201);
and U8898 (N_8898,N_8011,N_8151);
and U8899 (N_8899,N_8045,N_7689);
xnor U8900 (N_8900,N_7554,N_7963);
and U8901 (N_8901,N_8104,N_7873);
and U8902 (N_8902,N_7804,N_8199);
nand U8903 (N_8903,N_7814,N_7947);
nand U8904 (N_8904,N_7705,N_7529);
or U8905 (N_8905,N_7707,N_7583);
xnor U8906 (N_8906,N_8124,N_8089);
or U8907 (N_8907,N_7663,N_7691);
xor U8908 (N_8908,N_7851,N_7906);
nor U8909 (N_8909,N_7560,N_8217);
or U8910 (N_8910,N_8043,N_7933);
nand U8911 (N_8911,N_7945,N_7810);
nor U8912 (N_8912,N_8039,N_7765);
nand U8913 (N_8913,N_7616,N_8103);
xnor U8914 (N_8914,N_7829,N_8083);
nor U8915 (N_8915,N_8245,N_7963);
nand U8916 (N_8916,N_7864,N_8033);
or U8917 (N_8917,N_7936,N_7961);
or U8918 (N_8918,N_7618,N_8154);
or U8919 (N_8919,N_7798,N_7800);
xnor U8920 (N_8920,N_7596,N_8170);
or U8921 (N_8921,N_7984,N_8229);
nor U8922 (N_8922,N_7768,N_7978);
nand U8923 (N_8923,N_7727,N_8066);
and U8924 (N_8924,N_8063,N_7841);
nor U8925 (N_8925,N_7957,N_7506);
or U8926 (N_8926,N_7914,N_7775);
nor U8927 (N_8927,N_8005,N_8215);
xor U8928 (N_8928,N_8240,N_7595);
and U8929 (N_8929,N_8005,N_7504);
or U8930 (N_8930,N_7982,N_8013);
nand U8931 (N_8931,N_7871,N_8028);
nand U8932 (N_8932,N_7629,N_7791);
and U8933 (N_8933,N_7936,N_8190);
nand U8934 (N_8934,N_7639,N_7987);
nor U8935 (N_8935,N_7786,N_7585);
and U8936 (N_8936,N_7742,N_8246);
nand U8937 (N_8937,N_8142,N_7851);
or U8938 (N_8938,N_7997,N_7816);
or U8939 (N_8939,N_7815,N_8046);
xor U8940 (N_8940,N_7732,N_7813);
nor U8941 (N_8941,N_7574,N_7896);
nand U8942 (N_8942,N_7965,N_7888);
xor U8943 (N_8943,N_7776,N_7700);
and U8944 (N_8944,N_7974,N_8131);
nand U8945 (N_8945,N_7787,N_7899);
nand U8946 (N_8946,N_7704,N_8239);
xnor U8947 (N_8947,N_7707,N_7538);
or U8948 (N_8948,N_7714,N_7965);
and U8949 (N_8949,N_8011,N_7649);
xor U8950 (N_8950,N_7700,N_7550);
and U8951 (N_8951,N_7940,N_8204);
nand U8952 (N_8952,N_7983,N_7613);
or U8953 (N_8953,N_7640,N_7618);
and U8954 (N_8954,N_7922,N_7875);
nor U8955 (N_8955,N_8079,N_7684);
nand U8956 (N_8956,N_7816,N_7728);
nand U8957 (N_8957,N_8096,N_7522);
nor U8958 (N_8958,N_7822,N_8176);
nor U8959 (N_8959,N_8181,N_7594);
or U8960 (N_8960,N_7872,N_8249);
xor U8961 (N_8961,N_8008,N_7534);
nand U8962 (N_8962,N_7995,N_8240);
or U8963 (N_8963,N_7902,N_7593);
or U8964 (N_8964,N_7840,N_7660);
nand U8965 (N_8965,N_7791,N_7813);
or U8966 (N_8966,N_7879,N_7542);
and U8967 (N_8967,N_8171,N_7600);
or U8968 (N_8968,N_7842,N_8122);
and U8969 (N_8969,N_8243,N_7739);
or U8970 (N_8970,N_7657,N_7932);
or U8971 (N_8971,N_7682,N_7642);
nand U8972 (N_8972,N_7685,N_8086);
nand U8973 (N_8973,N_7820,N_7987);
or U8974 (N_8974,N_7827,N_8131);
nand U8975 (N_8975,N_7818,N_7676);
nand U8976 (N_8976,N_7601,N_7517);
and U8977 (N_8977,N_7510,N_7978);
or U8978 (N_8978,N_8063,N_7666);
nand U8979 (N_8979,N_7964,N_8187);
and U8980 (N_8980,N_7680,N_7718);
nand U8981 (N_8981,N_7825,N_8180);
nor U8982 (N_8982,N_8086,N_7771);
and U8983 (N_8983,N_7829,N_7882);
and U8984 (N_8984,N_7540,N_7749);
and U8985 (N_8985,N_7991,N_7616);
xor U8986 (N_8986,N_7778,N_7922);
xor U8987 (N_8987,N_8078,N_7927);
nand U8988 (N_8988,N_8141,N_8024);
nor U8989 (N_8989,N_7911,N_7929);
and U8990 (N_8990,N_8163,N_7800);
nand U8991 (N_8991,N_8097,N_8001);
and U8992 (N_8992,N_8076,N_8128);
xor U8993 (N_8993,N_7686,N_7965);
or U8994 (N_8994,N_7806,N_7810);
xnor U8995 (N_8995,N_7560,N_7736);
nor U8996 (N_8996,N_7720,N_8143);
nand U8997 (N_8997,N_8178,N_7771);
or U8998 (N_8998,N_7772,N_7805);
xor U8999 (N_8999,N_7542,N_7603);
nor U9000 (N_9000,N_8408,N_8284);
xor U9001 (N_9001,N_8867,N_8491);
nand U9002 (N_9002,N_8655,N_8393);
or U9003 (N_9003,N_8535,N_8870);
nand U9004 (N_9004,N_8565,N_8821);
nand U9005 (N_9005,N_8332,N_8404);
xnor U9006 (N_9006,N_8315,N_8728);
nand U9007 (N_9007,N_8878,N_8266);
xor U9008 (N_9008,N_8984,N_8989);
nor U9009 (N_9009,N_8832,N_8774);
xor U9010 (N_9010,N_8703,N_8659);
and U9011 (N_9011,N_8589,N_8440);
or U9012 (N_9012,N_8671,N_8987);
or U9013 (N_9013,N_8922,N_8667);
nand U9014 (N_9014,N_8304,N_8360);
nand U9015 (N_9015,N_8449,N_8646);
or U9016 (N_9016,N_8264,N_8926);
xnor U9017 (N_9017,N_8851,N_8390);
nand U9018 (N_9018,N_8840,N_8661);
xor U9019 (N_9019,N_8877,N_8364);
or U9020 (N_9020,N_8695,N_8379);
and U9021 (N_9021,N_8533,N_8584);
nand U9022 (N_9022,N_8442,N_8740);
and U9023 (N_9023,N_8770,N_8413);
or U9024 (N_9024,N_8674,N_8811);
nor U9025 (N_9025,N_8262,N_8638);
nor U9026 (N_9026,N_8686,N_8579);
xor U9027 (N_9027,N_8708,N_8521);
nor U9028 (N_9028,N_8791,N_8855);
xor U9029 (N_9029,N_8352,N_8267);
xnor U9030 (N_9030,N_8639,N_8810);
or U9031 (N_9031,N_8793,N_8577);
nand U9032 (N_9032,N_8309,N_8722);
xor U9033 (N_9033,N_8459,N_8316);
nand U9034 (N_9034,N_8279,N_8971);
nand U9035 (N_9035,N_8765,N_8471);
xnor U9036 (N_9036,N_8777,N_8709);
and U9037 (N_9037,N_8824,N_8961);
xor U9038 (N_9038,N_8356,N_8710);
nand U9039 (N_9039,N_8685,N_8548);
or U9040 (N_9040,N_8736,N_8788);
nor U9041 (N_9041,N_8590,N_8370);
and U9042 (N_9042,N_8907,N_8650);
xor U9043 (N_9043,N_8256,N_8976);
and U9044 (N_9044,N_8456,N_8475);
and U9045 (N_9045,N_8885,N_8813);
xnor U9046 (N_9046,N_8847,N_8787);
and U9047 (N_9047,N_8925,N_8617);
nor U9048 (N_9048,N_8322,N_8981);
xor U9049 (N_9049,N_8827,N_8918);
xor U9050 (N_9050,N_8437,N_8906);
and U9051 (N_9051,N_8883,N_8586);
nand U9052 (N_9052,N_8917,N_8994);
and U9053 (N_9053,N_8349,N_8596);
or U9054 (N_9054,N_8500,N_8758);
or U9055 (N_9055,N_8583,N_8453);
nor U9056 (N_9056,N_8476,N_8951);
xor U9057 (N_9057,N_8660,N_8553);
xnor U9058 (N_9058,N_8687,N_8371);
and U9059 (N_9059,N_8936,N_8864);
or U9060 (N_9060,N_8751,N_8959);
or U9061 (N_9061,N_8817,N_8897);
and U9062 (N_9062,N_8692,N_8572);
nand U9063 (N_9063,N_8842,N_8690);
nor U9064 (N_9064,N_8630,N_8624);
or U9065 (N_9065,N_8526,N_8465);
or U9066 (N_9066,N_8270,N_8991);
nand U9067 (N_9067,N_8537,N_8514);
or U9068 (N_9068,N_8462,N_8963);
or U9069 (N_9069,N_8620,N_8944);
nand U9070 (N_9070,N_8952,N_8560);
nor U9071 (N_9071,N_8310,N_8562);
or U9072 (N_9072,N_8990,N_8619);
nor U9073 (N_9073,N_8943,N_8454);
or U9074 (N_9074,N_8298,N_8552);
nand U9075 (N_9075,N_8445,N_8436);
and U9076 (N_9076,N_8693,N_8744);
or U9077 (N_9077,N_8752,N_8330);
nand U9078 (N_9078,N_8350,N_8326);
nand U9079 (N_9079,N_8894,N_8880);
xnor U9080 (N_9080,N_8292,N_8977);
or U9081 (N_9081,N_8490,N_8576);
nand U9082 (N_9082,N_8754,N_8282);
nand U9083 (N_9083,N_8250,N_8301);
nor U9084 (N_9084,N_8915,N_8392);
nor U9085 (N_9085,N_8458,N_8394);
nand U9086 (N_9086,N_8406,N_8988);
nand U9087 (N_9087,N_8343,N_8805);
nor U9088 (N_9088,N_8995,N_8835);
and U9089 (N_9089,N_8841,N_8644);
nor U9090 (N_9090,N_8539,N_8518);
nor U9091 (N_9091,N_8717,N_8574);
nor U9092 (N_9092,N_8732,N_8960);
or U9093 (N_9093,N_8252,N_8979);
nand U9094 (N_9094,N_8567,N_8783);
xor U9095 (N_9095,N_8724,N_8975);
nand U9096 (N_9096,N_8289,N_8320);
nand U9097 (N_9097,N_8482,N_8494);
nor U9098 (N_9098,N_8891,N_8965);
nor U9099 (N_9099,N_8499,N_8464);
and U9100 (N_9100,N_8381,N_8946);
or U9101 (N_9101,N_8798,N_8346);
nand U9102 (N_9102,N_8271,N_8358);
or U9103 (N_9103,N_8714,N_8578);
and U9104 (N_9104,N_8858,N_8697);
or U9105 (N_9105,N_8786,N_8418);
nor U9106 (N_9106,N_8654,N_8414);
and U9107 (N_9107,N_8592,N_8769);
or U9108 (N_9108,N_8524,N_8743);
and U9109 (N_9109,N_8748,N_8260);
nor U9110 (N_9110,N_8681,N_8625);
xnor U9111 (N_9111,N_8268,N_8274);
or U9112 (N_9112,N_8457,N_8919);
xor U9113 (N_9113,N_8604,N_8496);
or U9114 (N_9114,N_8269,N_8831);
or U9115 (N_9115,N_8741,N_8737);
nand U9116 (N_9116,N_8550,N_8492);
or U9117 (N_9117,N_8425,N_8334);
and U9118 (N_9118,N_8613,N_8790);
nand U9119 (N_9119,N_8280,N_8606);
nor U9120 (N_9120,N_8305,N_8512);
or U9121 (N_9121,N_8911,N_8795);
and U9122 (N_9122,N_8313,N_8410);
or U9123 (N_9123,N_8730,N_8966);
nand U9124 (N_9124,N_8816,N_8461);
xor U9125 (N_9125,N_8376,N_8347);
or U9126 (N_9126,N_8677,N_8297);
and U9127 (N_9127,N_8707,N_8747);
nor U9128 (N_9128,N_8520,N_8285);
and U9129 (N_9129,N_8557,N_8348);
nand U9130 (N_9130,N_8945,N_8649);
nor U9131 (N_9131,N_8993,N_8303);
nand U9132 (N_9132,N_8637,N_8941);
nor U9133 (N_9133,N_8780,N_8311);
nor U9134 (N_9134,N_8834,N_8389);
nand U9135 (N_9135,N_8529,N_8400);
nor U9136 (N_9136,N_8669,N_8293);
xor U9137 (N_9137,N_8399,N_8731);
nand U9138 (N_9138,N_8876,N_8433);
nor U9139 (N_9139,N_8678,N_8265);
nand U9140 (N_9140,N_8910,N_8614);
nand U9141 (N_9141,N_8366,N_8595);
nor U9142 (N_9142,N_8863,N_8713);
or U9143 (N_9143,N_8972,N_8643);
nand U9144 (N_9144,N_8628,N_8286);
and U9145 (N_9145,N_8294,N_8483);
or U9146 (N_9146,N_8931,N_8312);
nand U9147 (N_9147,N_8830,N_8575);
nand U9148 (N_9148,N_8645,N_8819);
nand U9149 (N_9149,N_8344,N_8683);
nand U9150 (N_9150,N_8386,N_8438);
nand U9151 (N_9151,N_8808,N_8853);
xnor U9152 (N_9152,N_8875,N_8856);
and U9153 (N_9153,N_8452,N_8429);
xor U9154 (N_9154,N_8964,N_8852);
nor U9155 (N_9155,N_8511,N_8278);
or U9156 (N_9156,N_8622,N_8582);
and U9157 (N_9157,N_8528,N_8460);
nand U9158 (N_9158,N_8849,N_8416);
and U9159 (N_9159,N_8684,N_8276);
or U9160 (N_9160,N_8397,N_8588);
xnor U9161 (N_9161,N_8986,N_8554);
or U9162 (N_9162,N_8869,N_8627);
nand U9163 (N_9163,N_8757,N_8942);
nand U9164 (N_9164,N_8792,N_8801);
or U9165 (N_9165,N_8339,N_8523);
nor U9166 (N_9166,N_8829,N_8663);
xnor U9167 (N_9167,N_8673,N_8776);
and U9168 (N_9168,N_8468,N_8635);
or U9169 (N_9169,N_8742,N_8314);
or U9170 (N_9170,N_8504,N_8647);
or U9171 (N_9171,N_8814,N_8680);
nand U9172 (N_9172,N_8585,N_8954);
nor U9173 (N_9173,N_8633,N_8632);
nor U9174 (N_9174,N_8750,N_8530);
nor U9175 (N_9175,N_8362,N_8275);
xor U9176 (N_9176,N_8718,N_8688);
nand U9177 (N_9177,N_8374,N_8928);
nor U9178 (N_9178,N_8825,N_8982);
xor U9179 (N_9179,N_8542,N_8525);
nor U9180 (N_9180,N_8761,N_8377);
xnor U9181 (N_9181,N_8658,N_8719);
nand U9182 (N_9182,N_8734,N_8336);
nor U9183 (N_9183,N_8721,N_8682);
xor U9184 (N_9184,N_8973,N_8306);
nor U9185 (N_9185,N_8327,N_8415);
xor U9186 (N_9186,N_8444,N_8401);
nor U9187 (N_9187,N_8365,N_8948);
xnor U9188 (N_9188,N_8898,N_8368);
xnor U9189 (N_9189,N_8342,N_8508);
nor U9190 (N_9190,N_8698,N_8921);
nor U9191 (N_9191,N_8833,N_8904);
xor U9192 (N_9192,N_8426,N_8281);
and U9193 (N_9193,N_8759,N_8920);
and U9194 (N_9194,N_8484,N_8985);
and U9195 (N_9195,N_8753,N_8321);
and U9196 (N_9196,N_8431,N_8794);
or U9197 (N_9197,N_8766,N_8570);
and U9198 (N_9198,N_8580,N_8738);
nand U9199 (N_9199,N_8258,N_8487);
xor U9200 (N_9200,N_8359,N_8725);
nand U9201 (N_9201,N_8610,N_8902);
and U9202 (N_9202,N_8479,N_8890);
or U9203 (N_9203,N_8341,N_8307);
nand U9204 (N_9204,N_8427,N_8652);
nand U9205 (N_9205,N_8493,N_8363);
nand U9206 (N_9206,N_8641,N_8317);
nor U9207 (N_9207,N_8937,N_8715);
or U9208 (N_9208,N_8527,N_8723);
or U9209 (N_9209,N_8909,N_8448);
or U9210 (N_9210,N_8519,N_8291);
xnor U9211 (N_9211,N_8727,N_8889);
or U9212 (N_9212,N_8809,N_8923);
and U9213 (N_9213,N_8749,N_8424);
and U9214 (N_9214,N_8656,N_8886);
nand U9215 (N_9215,N_8818,N_8665);
nand U9216 (N_9216,N_8802,N_8463);
and U9217 (N_9217,N_8451,N_8999);
xnor U9218 (N_9218,N_8380,N_8899);
and U9219 (N_9219,N_8544,N_8272);
nor U9220 (N_9220,N_8607,N_8323);
or U9221 (N_9221,N_8516,N_8497);
nor U9222 (N_9222,N_8324,N_8395);
or U9223 (N_9223,N_8396,N_8373);
or U9224 (N_9224,N_8300,N_8446);
and U9225 (N_9225,N_8615,N_8599);
or U9226 (N_9226,N_8308,N_8608);
nor U9227 (N_9227,N_8417,N_8908);
or U9228 (N_9228,N_8561,N_8640);
and U9229 (N_9229,N_8700,N_8779);
nor U9230 (N_9230,N_8800,N_8968);
or U9231 (N_9231,N_8563,N_8861);
or U9232 (N_9232,N_8566,N_8903);
nand U9233 (N_9233,N_8486,N_8472);
and U9234 (N_9234,N_8837,N_8419);
and U9235 (N_9235,N_8338,N_8789);
xnor U9236 (N_9236,N_8532,N_8962);
nand U9237 (N_9237,N_8935,N_8670);
nand U9238 (N_9238,N_8657,N_8916);
nor U9239 (N_9239,N_8953,N_8337);
xnor U9240 (N_9240,N_8760,N_8871);
xnor U9241 (N_9241,N_8502,N_8771);
nand U9242 (N_9242,N_8699,N_8912);
nor U9243 (N_9243,N_8277,N_8896);
or U9244 (N_9244,N_8488,N_8573);
nor U9245 (N_9245,N_8768,N_8998);
nand U9246 (N_9246,N_8679,N_8905);
xor U9247 (N_9247,N_8978,N_8611);
nor U9248 (N_9248,N_8353,N_8933);
xor U9249 (N_9249,N_8803,N_8704);
and U9250 (N_9250,N_8967,N_8259);
nand U9251 (N_9251,N_8868,N_8290);
or U9252 (N_9252,N_8781,N_8372);
xnor U9253 (N_9253,N_8545,N_8866);
and U9254 (N_9254,N_8569,N_8762);
nand U9255 (N_9255,N_8447,N_8432);
nand U9256 (N_9256,N_8295,N_8980);
nor U9257 (N_9257,N_8325,N_8631);
xor U9258 (N_9258,N_8473,N_8845);
and U9259 (N_9259,N_8318,N_8838);
nor U9260 (N_9260,N_8938,N_8505);
nand U9261 (N_9261,N_8357,N_8540);
nor U9262 (N_9262,N_8634,N_8651);
nor U9263 (N_9263,N_8756,N_8969);
nand U9264 (N_9264,N_8839,N_8434);
xnor U9265 (N_9265,N_8844,N_8836);
nand U9266 (N_9266,N_8388,N_8764);
nand U9267 (N_9267,N_8807,N_8712);
xor U9268 (N_9268,N_8273,N_8873);
or U9269 (N_9269,N_8387,N_8403);
nor U9270 (N_9270,N_8820,N_8772);
and U9271 (N_9271,N_8797,N_8559);
nor U9272 (N_9272,N_8881,N_8601);
and U9273 (N_9273,N_8331,N_8609);
and U9274 (N_9274,N_8402,N_8335);
nor U9275 (N_9275,N_8924,N_8549);
nand U9276 (N_9276,N_8299,N_8796);
and U9277 (N_9277,N_8531,N_8506);
and U9278 (N_9278,N_8913,N_8859);
or U9279 (N_9279,N_8423,N_8405);
or U9280 (N_9280,N_8329,N_8806);
or U9281 (N_9281,N_8428,N_8594);
nand U9282 (N_9282,N_8287,N_8892);
nand U9283 (N_9283,N_8857,N_8478);
or U9284 (N_9284,N_8812,N_8828);
or U9285 (N_9285,N_8927,N_8420);
xnor U9286 (N_9286,N_8662,N_8351);
nand U9287 (N_9287,N_8668,N_8412);
nand U9288 (N_9288,N_8653,N_8672);
or U9289 (N_9289,N_8354,N_8997);
nor U9290 (N_9290,N_8355,N_8739);
or U9291 (N_9291,N_8605,N_8872);
and U9292 (N_9292,N_8887,N_8664);
or U9293 (N_9293,N_8398,N_8571);
nand U9294 (N_9294,N_8782,N_8815);
and U9295 (N_9295,N_8435,N_8636);
and U9296 (N_9296,N_8253,N_8507);
nand U9297 (N_9297,N_8261,N_8450);
nand U9298 (N_9298,N_8843,N_8974);
nor U9299 (N_9299,N_8480,N_8711);
nand U9300 (N_9300,N_8591,N_8485);
nand U9301 (N_9301,N_8581,N_8558);
or U9302 (N_9302,N_8618,N_8534);
and U9303 (N_9303,N_8541,N_8407);
or U9304 (N_9304,N_8538,N_8467);
and U9305 (N_9305,N_8564,N_8513);
nor U9306 (N_9306,N_8746,N_8934);
and U9307 (N_9307,N_8701,N_8455);
nor U9308 (N_9308,N_8501,N_8983);
nand U9309 (N_9309,N_8895,N_8716);
nand U9310 (N_9310,N_8775,N_8642);
nand U9311 (N_9311,N_8726,N_8283);
nand U9312 (N_9312,N_8546,N_8375);
xor U9313 (N_9313,N_8773,N_8826);
nand U9314 (N_9314,N_8848,N_8383);
or U9315 (N_9315,N_8755,N_8555);
xnor U9316 (N_9316,N_8378,N_8430);
nor U9317 (N_9317,N_8939,N_8691);
nor U9318 (N_9318,N_8862,N_8823);
nor U9319 (N_9319,N_8495,N_8477);
nor U9320 (N_9320,N_8955,N_8391);
nor U9321 (N_9321,N_8603,N_8345);
nand U9322 (N_9322,N_8958,N_8846);
nor U9323 (N_9323,N_8850,N_8947);
nor U9324 (N_9324,N_8551,N_8257);
nor U9325 (N_9325,N_8469,N_8956);
and U9326 (N_9326,N_8503,N_8996);
and U9327 (N_9327,N_8598,N_8474);
nand U9328 (N_9328,N_8860,N_8612);
nand U9329 (N_9329,N_8706,N_8522);
and U9330 (N_9330,N_8296,N_8616);
nor U9331 (N_9331,N_8696,N_8255);
nand U9332 (N_9332,N_8421,N_8689);
xnor U9333 (N_9333,N_8992,N_8874);
xor U9334 (N_9334,N_8536,N_8914);
xor U9335 (N_9335,N_8422,N_8543);
nand U9336 (N_9336,N_8621,N_8367);
nand U9337 (N_9337,N_8510,N_8626);
nand U9338 (N_9338,N_8470,N_8932);
and U9339 (N_9339,N_8733,N_8441);
and U9340 (N_9340,N_8443,N_8593);
nand U9341 (N_9341,N_8694,N_8288);
and U9342 (N_9342,N_8369,N_8720);
and U9343 (N_9343,N_8333,N_8785);
nand U9344 (N_9344,N_8385,N_8804);
and U9345 (N_9345,N_8489,N_8778);
nor U9346 (N_9346,N_8629,N_8957);
xnor U9347 (N_9347,N_8328,N_8623);
nand U9348 (N_9348,N_8498,N_8822);
or U9349 (N_9349,N_8597,N_8745);
xor U9350 (N_9350,N_8767,N_8949);
and U9351 (N_9351,N_8854,N_8515);
or U9352 (N_9352,N_8340,N_8729);
xnor U9353 (N_9353,N_8929,N_8705);
nor U9354 (N_9354,N_8702,N_8888);
nor U9355 (N_9355,N_8600,N_8556);
nor U9356 (N_9356,N_8568,N_8882);
and U9357 (N_9357,N_8382,N_8676);
nor U9358 (N_9358,N_8466,N_8666);
and U9359 (N_9359,N_8648,N_8901);
or U9360 (N_9360,N_8251,N_8439);
and U9361 (N_9361,N_8865,N_8940);
nor U9362 (N_9362,N_8950,N_8547);
or U9363 (N_9363,N_8587,N_8302);
and U9364 (N_9364,N_8384,N_8675);
and U9365 (N_9365,N_8263,N_8254);
or U9366 (N_9366,N_8411,N_8799);
and U9367 (N_9367,N_8481,N_8900);
nand U9368 (N_9368,N_8879,N_8509);
and U9369 (N_9369,N_8784,N_8763);
or U9370 (N_9370,N_8930,N_8409);
and U9371 (N_9371,N_8602,N_8361);
and U9372 (N_9372,N_8517,N_8735);
or U9373 (N_9373,N_8970,N_8319);
or U9374 (N_9374,N_8884,N_8893);
or U9375 (N_9375,N_8381,N_8975);
and U9376 (N_9376,N_8263,N_8535);
and U9377 (N_9377,N_8770,N_8893);
and U9378 (N_9378,N_8758,N_8254);
nand U9379 (N_9379,N_8921,N_8780);
or U9380 (N_9380,N_8268,N_8400);
xor U9381 (N_9381,N_8687,N_8251);
nand U9382 (N_9382,N_8411,N_8630);
or U9383 (N_9383,N_8673,N_8377);
nor U9384 (N_9384,N_8316,N_8862);
or U9385 (N_9385,N_8359,N_8299);
and U9386 (N_9386,N_8790,N_8445);
or U9387 (N_9387,N_8844,N_8621);
or U9388 (N_9388,N_8909,N_8766);
or U9389 (N_9389,N_8291,N_8746);
or U9390 (N_9390,N_8975,N_8375);
or U9391 (N_9391,N_8352,N_8543);
nand U9392 (N_9392,N_8823,N_8735);
nand U9393 (N_9393,N_8477,N_8337);
nand U9394 (N_9394,N_8728,N_8761);
xnor U9395 (N_9395,N_8548,N_8812);
xor U9396 (N_9396,N_8497,N_8812);
and U9397 (N_9397,N_8359,N_8591);
and U9398 (N_9398,N_8758,N_8339);
and U9399 (N_9399,N_8899,N_8888);
nand U9400 (N_9400,N_8971,N_8610);
nor U9401 (N_9401,N_8750,N_8423);
nor U9402 (N_9402,N_8558,N_8430);
xor U9403 (N_9403,N_8825,N_8574);
or U9404 (N_9404,N_8709,N_8836);
or U9405 (N_9405,N_8382,N_8728);
nor U9406 (N_9406,N_8779,N_8366);
nor U9407 (N_9407,N_8626,N_8842);
nand U9408 (N_9408,N_8655,N_8789);
xnor U9409 (N_9409,N_8284,N_8398);
and U9410 (N_9410,N_8302,N_8520);
nand U9411 (N_9411,N_8791,N_8717);
nor U9412 (N_9412,N_8862,N_8837);
nand U9413 (N_9413,N_8653,N_8408);
and U9414 (N_9414,N_8396,N_8635);
nand U9415 (N_9415,N_8385,N_8846);
xor U9416 (N_9416,N_8575,N_8818);
nand U9417 (N_9417,N_8958,N_8391);
and U9418 (N_9418,N_8708,N_8358);
xor U9419 (N_9419,N_8348,N_8935);
nor U9420 (N_9420,N_8426,N_8506);
xor U9421 (N_9421,N_8576,N_8500);
and U9422 (N_9422,N_8981,N_8813);
xor U9423 (N_9423,N_8657,N_8384);
and U9424 (N_9424,N_8541,N_8567);
xor U9425 (N_9425,N_8256,N_8619);
and U9426 (N_9426,N_8895,N_8436);
nor U9427 (N_9427,N_8677,N_8735);
xor U9428 (N_9428,N_8768,N_8805);
nor U9429 (N_9429,N_8993,N_8507);
or U9430 (N_9430,N_8528,N_8284);
and U9431 (N_9431,N_8445,N_8377);
and U9432 (N_9432,N_8614,N_8744);
nor U9433 (N_9433,N_8658,N_8377);
nor U9434 (N_9434,N_8373,N_8962);
nor U9435 (N_9435,N_8664,N_8729);
nand U9436 (N_9436,N_8809,N_8864);
nor U9437 (N_9437,N_8534,N_8680);
xor U9438 (N_9438,N_8673,N_8284);
xnor U9439 (N_9439,N_8954,N_8600);
xor U9440 (N_9440,N_8804,N_8424);
xnor U9441 (N_9441,N_8700,N_8755);
nand U9442 (N_9442,N_8851,N_8526);
xnor U9443 (N_9443,N_8911,N_8946);
nor U9444 (N_9444,N_8891,N_8617);
nor U9445 (N_9445,N_8350,N_8660);
xnor U9446 (N_9446,N_8544,N_8725);
and U9447 (N_9447,N_8377,N_8534);
nand U9448 (N_9448,N_8540,N_8749);
nor U9449 (N_9449,N_8935,N_8375);
nand U9450 (N_9450,N_8586,N_8955);
or U9451 (N_9451,N_8375,N_8960);
and U9452 (N_9452,N_8479,N_8763);
and U9453 (N_9453,N_8718,N_8374);
nand U9454 (N_9454,N_8872,N_8524);
xnor U9455 (N_9455,N_8656,N_8358);
xnor U9456 (N_9456,N_8661,N_8403);
xnor U9457 (N_9457,N_8739,N_8362);
xor U9458 (N_9458,N_8325,N_8693);
and U9459 (N_9459,N_8956,N_8940);
nor U9460 (N_9460,N_8814,N_8792);
or U9461 (N_9461,N_8539,N_8514);
nor U9462 (N_9462,N_8733,N_8304);
and U9463 (N_9463,N_8974,N_8925);
or U9464 (N_9464,N_8624,N_8403);
xnor U9465 (N_9465,N_8499,N_8928);
or U9466 (N_9466,N_8877,N_8427);
xnor U9467 (N_9467,N_8544,N_8871);
xor U9468 (N_9468,N_8772,N_8354);
xor U9469 (N_9469,N_8964,N_8499);
and U9470 (N_9470,N_8293,N_8284);
or U9471 (N_9471,N_8726,N_8914);
or U9472 (N_9472,N_8323,N_8823);
or U9473 (N_9473,N_8845,N_8991);
and U9474 (N_9474,N_8421,N_8272);
xor U9475 (N_9475,N_8732,N_8747);
xor U9476 (N_9476,N_8823,N_8352);
nor U9477 (N_9477,N_8827,N_8507);
nor U9478 (N_9478,N_8431,N_8279);
or U9479 (N_9479,N_8998,N_8925);
or U9480 (N_9480,N_8476,N_8618);
nor U9481 (N_9481,N_8361,N_8670);
and U9482 (N_9482,N_8737,N_8582);
nand U9483 (N_9483,N_8588,N_8947);
xor U9484 (N_9484,N_8640,N_8383);
and U9485 (N_9485,N_8639,N_8929);
nor U9486 (N_9486,N_8250,N_8569);
nand U9487 (N_9487,N_8547,N_8643);
nand U9488 (N_9488,N_8334,N_8716);
or U9489 (N_9489,N_8790,N_8750);
nand U9490 (N_9490,N_8371,N_8336);
nand U9491 (N_9491,N_8646,N_8683);
and U9492 (N_9492,N_8803,N_8613);
nand U9493 (N_9493,N_8806,N_8766);
or U9494 (N_9494,N_8878,N_8789);
nand U9495 (N_9495,N_8409,N_8977);
xnor U9496 (N_9496,N_8660,N_8428);
and U9497 (N_9497,N_8364,N_8669);
nor U9498 (N_9498,N_8639,N_8377);
or U9499 (N_9499,N_8322,N_8819);
nor U9500 (N_9500,N_8777,N_8571);
xnor U9501 (N_9501,N_8469,N_8531);
nor U9502 (N_9502,N_8384,N_8798);
or U9503 (N_9503,N_8561,N_8366);
nand U9504 (N_9504,N_8358,N_8609);
nor U9505 (N_9505,N_8313,N_8361);
nand U9506 (N_9506,N_8537,N_8894);
nor U9507 (N_9507,N_8755,N_8880);
or U9508 (N_9508,N_8932,N_8559);
and U9509 (N_9509,N_8749,N_8607);
xnor U9510 (N_9510,N_8936,N_8552);
and U9511 (N_9511,N_8978,N_8725);
and U9512 (N_9512,N_8344,N_8366);
nor U9513 (N_9513,N_8900,N_8571);
xor U9514 (N_9514,N_8371,N_8386);
xnor U9515 (N_9515,N_8384,N_8631);
xor U9516 (N_9516,N_8881,N_8814);
nor U9517 (N_9517,N_8485,N_8537);
nor U9518 (N_9518,N_8997,N_8423);
xor U9519 (N_9519,N_8643,N_8970);
xnor U9520 (N_9520,N_8384,N_8920);
nand U9521 (N_9521,N_8822,N_8879);
nor U9522 (N_9522,N_8656,N_8675);
and U9523 (N_9523,N_8573,N_8580);
nand U9524 (N_9524,N_8800,N_8542);
and U9525 (N_9525,N_8507,N_8488);
and U9526 (N_9526,N_8776,N_8328);
xnor U9527 (N_9527,N_8745,N_8771);
or U9528 (N_9528,N_8756,N_8484);
or U9529 (N_9529,N_8820,N_8965);
nand U9530 (N_9530,N_8456,N_8932);
or U9531 (N_9531,N_8293,N_8741);
nand U9532 (N_9532,N_8723,N_8324);
or U9533 (N_9533,N_8753,N_8694);
xnor U9534 (N_9534,N_8325,N_8820);
or U9535 (N_9535,N_8671,N_8318);
nand U9536 (N_9536,N_8813,N_8292);
and U9537 (N_9537,N_8388,N_8552);
or U9538 (N_9538,N_8611,N_8937);
nand U9539 (N_9539,N_8515,N_8909);
and U9540 (N_9540,N_8478,N_8272);
and U9541 (N_9541,N_8471,N_8634);
xnor U9542 (N_9542,N_8295,N_8860);
xnor U9543 (N_9543,N_8592,N_8703);
nor U9544 (N_9544,N_8501,N_8444);
xor U9545 (N_9545,N_8776,N_8669);
or U9546 (N_9546,N_8400,N_8610);
nand U9547 (N_9547,N_8632,N_8482);
nor U9548 (N_9548,N_8471,N_8334);
nand U9549 (N_9549,N_8293,N_8757);
nor U9550 (N_9550,N_8682,N_8917);
xnor U9551 (N_9551,N_8408,N_8506);
and U9552 (N_9552,N_8490,N_8857);
nor U9553 (N_9553,N_8566,N_8578);
xnor U9554 (N_9554,N_8730,N_8595);
and U9555 (N_9555,N_8343,N_8456);
nor U9556 (N_9556,N_8838,N_8389);
nand U9557 (N_9557,N_8306,N_8718);
nand U9558 (N_9558,N_8586,N_8650);
nor U9559 (N_9559,N_8464,N_8819);
nor U9560 (N_9560,N_8264,N_8465);
nand U9561 (N_9561,N_8792,N_8494);
xnor U9562 (N_9562,N_8577,N_8365);
and U9563 (N_9563,N_8907,N_8915);
and U9564 (N_9564,N_8303,N_8865);
nor U9565 (N_9565,N_8674,N_8917);
and U9566 (N_9566,N_8410,N_8802);
nor U9567 (N_9567,N_8257,N_8763);
xor U9568 (N_9568,N_8750,N_8798);
xor U9569 (N_9569,N_8282,N_8286);
and U9570 (N_9570,N_8755,N_8720);
and U9571 (N_9571,N_8607,N_8666);
nand U9572 (N_9572,N_8850,N_8361);
nand U9573 (N_9573,N_8558,N_8413);
nor U9574 (N_9574,N_8684,N_8260);
and U9575 (N_9575,N_8284,N_8354);
and U9576 (N_9576,N_8431,N_8304);
nor U9577 (N_9577,N_8388,N_8623);
xnor U9578 (N_9578,N_8302,N_8739);
nor U9579 (N_9579,N_8637,N_8503);
nor U9580 (N_9580,N_8470,N_8720);
and U9581 (N_9581,N_8367,N_8900);
nand U9582 (N_9582,N_8781,N_8723);
and U9583 (N_9583,N_8769,N_8327);
xor U9584 (N_9584,N_8472,N_8754);
xnor U9585 (N_9585,N_8277,N_8597);
and U9586 (N_9586,N_8284,N_8579);
xor U9587 (N_9587,N_8808,N_8811);
or U9588 (N_9588,N_8776,N_8455);
nor U9589 (N_9589,N_8623,N_8777);
nor U9590 (N_9590,N_8918,N_8533);
nor U9591 (N_9591,N_8458,N_8547);
and U9592 (N_9592,N_8303,N_8397);
or U9593 (N_9593,N_8497,N_8307);
xor U9594 (N_9594,N_8807,N_8804);
and U9595 (N_9595,N_8578,N_8467);
nand U9596 (N_9596,N_8995,N_8336);
or U9597 (N_9597,N_8716,N_8392);
and U9598 (N_9598,N_8886,N_8388);
xor U9599 (N_9599,N_8885,N_8754);
nand U9600 (N_9600,N_8729,N_8840);
nand U9601 (N_9601,N_8940,N_8296);
nand U9602 (N_9602,N_8863,N_8557);
and U9603 (N_9603,N_8478,N_8316);
nand U9604 (N_9604,N_8400,N_8483);
and U9605 (N_9605,N_8408,N_8604);
or U9606 (N_9606,N_8599,N_8399);
and U9607 (N_9607,N_8760,N_8684);
nor U9608 (N_9608,N_8843,N_8727);
or U9609 (N_9609,N_8581,N_8438);
nand U9610 (N_9610,N_8963,N_8679);
and U9611 (N_9611,N_8708,N_8633);
xnor U9612 (N_9612,N_8538,N_8271);
nor U9613 (N_9613,N_8578,N_8942);
nor U9614 (N_9614,N_8388,N_8785);
nor U9615 (N_9615,N_8501,N_8515);
nor U9616 (N_9616,N_8488,N_8744);
nand U9617 (N_9617,N_8891,N_8918);
xor U9618 (N_9618,N_8572,N_8482);
and U9619 (N_9619,N_8287,N_8684);
nand U9620 (N_9620,N_8553,N_8343);
nor U9621 (N_9621,N_8516,N_8527);
or U9622 (N_9622,N_8419,N_8988);
or U9623 (N_9623,N_8359,N_8343);
nand U9624 (N_9624,N_8985,N_8849);
nor U9625 (N_9625,N_8483,N_8793);
xor U9626 (N_9626,N_8819,N_8864);
or U9627 (N_9627,N_8313,N_8272);
nor U9628 (N_9628,N_8486,N_8858);
nand U9629 (N_9629,N_8567,N_8836);
and U9630 (N_9630,N_8954,N_8925);
xnor U9631 (N_9631,N_8502,N_8907);
and U9632 (N_9632,N_8469,N_8842);
or U9633 (N_9633,N_8505,N_8625);
nand U9634 (N_9634,N_8677,N_8864);
or U9635 (N_9635,N_8637,N_8479);
nand U9636 (N_9636,N_8821,N_8392);
nor U9637 (N_9637,N_8350,N_8773);
or U9638 (N_9638,N_8615,N_8285);
nor U9639 (N_9639,N_8420,N_8414);
and U9640 (N_9640,N_8799,N_8964);
and U9641 (N_9641,N_8713,N_8779);
and U9642 (N_9642,N_8641,N_8599);
nand U9643 (N_9643,N_8414,N_8435);
nor U9644 (N_9644,N_8431,N_8704);
nor U9645 (N_9645,N_8942,N_8406);
or U9646 (N_9646,N_8523,N_8854);
nor U9647 (N_9647,N_8447,N_8458);
or U9648 (N_9648,N_8304,N_8791);
nand U9649 (N_9649,N_8345,N_8845);
nand U9650 (N_9650,N_8738,N_8523);
or U9651 (N_9651,N_8520,N_8982);
and U9652 (N_9652,N_8796,N_8715);
nor U9653 (N_9653,N_8718,N_8545);
xor U9654 (N_9654,N_8360,N_8909);
xnor U9655 (N_9655,N_8877,N_8598);
nand U9656 (N_9656,N_8826,N_8983);
and U9657 (N_9657,N_8722,N_8687);
and U9658 (N_9658,N_8331,N_8669);
nand U9659 (N_9659,N_8524,N_8968);
xor U9660 (N_9660,N_8371,N_8342);
nand U9661 (N_9661,N_8970,N_8978);
and U9662 (N_9662,N_8603,N_8353);
or U9663 (N_9663,N_8732,N_8567);
nor U9664 (N_9664,N_8565,N_8324);
nand U9665 (N_9665,N_8651,N_8746);
xor U9666 (N_9666,N_8522,N_8552);
or U9667 (N_9667,N_8936,N_8884);
xnor U9668 (N_9668,N_8647,N_8386);
nor U9669 (N_9669,N_8371,N_8465);
nand U9670 (N_9670,N_8967,N_8885);
xnor U9671 (N_9671,N_8652,N_8312);
nor U9672 (N_9672,N_8684,N_8614);
nand U9673 (N_9673,N_8371,N_8963);
nor U9674 (N_9674,N_8279,N_8802);
nand U9675 (N_9675,N_8724,N_8593);
or U9676 (N_9676,N_8931,N_8559);
or U9677 (N_9677,N_8484,N_8312);
or U9678 (N_9678,N_8287,N_8602);
nand U9679 (N_9679,N_8951,N_8955);
or U9680 (N_9680,N_8822,N_8504);
xor U9681 (N_9681,N_8661,N_8774);
xor U9682 (N_9682,N_8967,N_8844);
nor U9683 (N_9683,N_8985,N_8260);
xor U9684 (N_9684,N_8570,N_8697);
and U9685 (N_9685,N_8981,N_8603);
nand U9686 (N_9686,N_8405,N_8804);
xor U9687 (N_9687,N_8259,N_8434);
or U9688 (N_9688,N_8448,N_8590);
nand U9689 (N_9689,N_8429,N_8728);
nand U9690 (N_9690,N_8403,N_8774);
xnor U9691 (N_9691,N_8602,N_8259);
nand U9692 (N_9692,N_8802,N_8983);
or U9693 (N_9693,N_8430,N_8920);
nand U9694 (N_9694,N_8257,N_8778);
nor U9695 (N_9695,N_8891,N_8541);
xor U9696 (N_9696,N_8460,N_8255);
or U9697 (N_9697,N_8676,N_8716);
or U9698 (N_9698,N_8255,N_8714);
or U9699 (N_9699,N_8970,N_8508);
and U9700 (N_9700,N_8962,N_8673);
and U9701 (N_9701,N_8721,N_8882);
nand U9702 (N_9702,N_8593,N_8257);
or U9703 (N_9703,N_8434,N_8722);
nor U9704 (N_9704,N_8688,N_8504);
or U9705 (N_9705,N_8482,N_8750);
or U9706 (N_9706,N_8944,N_8421);
nand U9707 (N_9707,N_8432,N_8866);
xor U9708 (N_9708,N_8913,N_8662);
or U9709 (N_9709,N_8343,N_8887);
nor U9710 (N_9710,N_8485,N_8959);
xnor U9711 (N_9711,N_8262,N_8587);
and U9712 (N_9712,N_8288,N_8406);
and U9713 (N_9713,N_8393,N_8335);
xor U9714 (N_9714,N_8264,N_8664);
nor U9715 (N_9715,N_8324,N_8573);
nor U9716 (N_9716,N_8851,N_8623);
or U9717 (N_9717,N_8388,N_8539);
nand U9718 (N_9718,N_8320,N_8900);
xor U9719 (N_9719,N_8619,N_8284);
nand U9720 (N_9720,N_8362,N_8773);
nand U9721 (N_9721,N_8629,N_8274);
nand U9722 (N_9722,N_8696,N_8769);
nor U9723 (N_9723,N_8410,N_8960);
or U9724 (N_9724,N_8541,N_8901);
or U9725 (N_9725,N_8304,N_8513);
xnor U9726 (N_9726,N_8283,N_8953);
xnor U9727 (N_9727,N_8516,N_8750);
xnor U9728 (N_9728,N_8632,N_8777);
nor U9729 (N_9729,N_8546,N_8855);
nand U9730 (N_9730,N_8284,N_8660);
nor U9731 (N_9731,N_8949,N_8390);
nor U9732 (N_9732,N_8604,N_8948);
nor U9733 (N_9733,N_8585,N_8837);
nand U9734 (N_9734,N_8687,N_8680);
and U9735 (N_9735,N_8534,N_8530);
nor U9736 (N_9736,N_8520,N_8722);
xor U9737 (N_9737,N_8600,N_8691);
nand U9738 (N_9738,N_8604,N_8683);
xor U9739 (N_9739,N_8537,N_8760);
nand U9740 (N_9740,N_8705,N_8833);
and U9741 (N_9741,N_8520,N_8921);
or U9742 (N_9742,N_8811,N_8719);
nand U9743 (N_9743,N_8528,N_8588);
xor U9744 (N_9744,N_8989,N_8673);
nand U9745 (N_9745,N_8865,N_8782);
nand U9746 (N_9746,N_8596,N_8636);
xnor U9747 (N_9747,N_8397,N_8648);
and U9748 (N_9748,N_8994,N_8433);
nand U9749 (N_9749,N_8618,N_8548);
xor U9750 (N_9750,N_9569,N_9572);
xor U9751 (N_9751,N_9149,N_9407);
or U9752 (N_9752,N_9648,N_9595);
or U9753 (N_9753,N_9195,N_9730);
nor U9754 (N_9754,N_9035,N_9462);
or U9755 (N_9755,N_9282,N_9145);
and U9756 (N_9756,N_9642,N_9689);
and U9757 (N_9757,N_9535,N_9251);
and U9758 (N_9758,N_9245,N_9077);
or U9759 (N_9759,N_9290,N_9734);
xor U9760 (N_9760,N_9653,N_9682);
nor U9761 (N_9761,N_9307,N_9433);
nor U9762 (N_9762,N_9302,N_9702);
nand U9763 (N_9763,N_9122,N_9184);
and U9764 (N_9764,N_9454,N_9631);
nand U9765 (N_9765,N_9201,N_9616);
and U9766 (N_9766,N_9661,N_9691);
nand U9767 (N_9767,N_9400,N_9603);
xor U9768 (N_9768,N_9353,N_9581);
xnor U9769 (N_9769,N_9080,N_9586);
xor U9770 (N_9770,N_9651,N_9622);
nor U9771 (N_9771,N_9443,N_9376);
nor U9772 (N_9772,N_9187,N_9357);
or U9773 (N_9773,N_9529,N_9742);
nor U9774 (N_9774,N_9155,N_9150);
xor U9775 (N_9775,N_9013,N_9496);
xor U9776 (N_9776,N_9102,N_9674);
nand U9777 (N_9777,N_9512,N_9287);
or U9778 (N_9778,N_9460,N_9612);
nor U9779 (N_9779,N_9098,N_9555);
or U9780 (N_9780,N_9398,N_9303);
xnor U9781 (N_9781,N_9741,N_9470);
nand U9782 (N_9782,N_9037,N_9670);
and U9783 (N_9783,N_9254,N_9683);
xor U9784 (N_9784,N_9310,N_9226);
or U9785 (N_9785,N_9731,N_9038);
or U9786 (N_9786,N_9285,N_9534);
or U9787 (N_9787,N_9279,N_9486);
nand U9788 (N_9788,N_9000,N_9095);
xor U9789 (N_9789,N_9253,N_9543);
nand U9790 (N_9790,N_9317,N_9297);
nor U9791 (N_9791,N_9403,N_9424);
xor U9792 (N_9792,N_9503,N_9110);
xnor U9793 (N_9793,N_9343,N_9561);
xor U9794 (N_9794,N_9236,N_9594);
or U9795 (N_9795,N_9001,N_9576);
xor U9796 (N_9796,N_9606,N_9481);
xnor U9797 (N_9797,N_9719,N_9419);
or U9798 (N_9798,N_9469,N_9414);
nor U9799 (N_9799,N_9489,N_9578);
and U9800 (N_9800,N_9692,N_9560);
xor U9801 (N_9801,N_9193,N_9665);
and U9802 (N_9802,N_9428,N_9081);
or U9803 (N_9803,N_9729,N_9020);
xor U9804 (N_9804,N_9492,N_9459);
or U9805 (N_9805,N_9422,N_9521);
or U9806 (N_9806,N_9579,N_9371);
or U9807 (N_9807,N_9677,N_9427);
xor U9808 (N_9808,N_9544,N_9461);
and U9809 (N_9809,N_9699,N_9368);
xnor U9810 (N_9810,N_9620,N_9221);
or U9811 (N_9811,N_9264,N_9608);
xnor U9812 (N_9812,N_9553,N_9203);
or U9813 (N_9813,N_9412,N_9005);
nand U9814 (N_9814,N_9183,N_9749);
and U9815 (N_9815,N_9554,N_9130);
nand U9816 (N_9816,N_9585,N_9465);
and U9817 (N_9817,N_9509,N_9501);
nand U9818 (N_9818,N_9530,N_9362);
and U9819 (N_9819,N_9004,N_9637);
nor U9820 (N_9820,N_9190,N_9315);
and U9821 (N_9821,N_9152,N_9497);
and U9822 (N_9822,N_9291,N_9338);
xor U9823 (N_9823,N_9517,N_9069);
or U9824 (N_9824,N_9467,N_9344);
nor U9825 (N_9825,N_9570,N_9527);
and U9826 (N_9826,N_9507,N_9361);
or U9827 (N_9827,N_9246,N_9432);
nor U9828 (N_9828,N_9697,N_9024);
xor U9829 (N_9829,N_9619,N_9654);
or U9830 (N_9830,N_9066,N_9225);
nand U9831 (N_9831,N_9073,N_9181);
xor U9832 (N_9832,N_9533,N_9026);
or U9833 (N_9833,N_9087,N_9717);
or U9834 (N_9834,N_9546,N_9207);
nand U9835 (N_9835,N_9611,N_9289);
nand U9836 (N_9836,N_9687,N_9049);
nand U9837 (N_9837,N_9321,N_9377);
and U9838 (N_9838,N_9009,N_9593);
or U9839 (N_9839,N_9538,N_9384);
xnor U9840 (N_9840,N_9262,N_9526);
or U9841 (N_9841,N_9506,N_9390);
or U9842 (N_9842,N_9397,N_9288);
xnor U9843 (N_9843,N_9453,N_9045);
nor U9844 (N_9844,N_9350,N_9118);
xnor U9845 (N_9845,N_9278,N_9483);
nand U9846 (N_9846,N_9723,N_9513);
and U9847 (N_9847,N_9295,N_9267);
or U9848 (N_9848,N_9649,N_9093);
xor U9849 (N_9849,N_9180,N_9146);
nand U9850 (N_9850,N_9401,N_9541);
xnor U9851 (N_9851,N_9652,N_9331);
or U9852 (N_9852,N_9259,N_9205);
and U9853 (N_9853,N_9125,N_9047);
and U9854 (N_9854,N_9173,N_9564);
or U9855 (N_9855,N_9031,N_9714);
and U9856 (N_9856,N_9434,N_9456);
nand U9857 (N_9857,N_9363,N_9466);
nand U9858 (N_9858,N_9070,N_9157);
or U9859 (N_9859,N_9613,N_9010);
and U9860 (N_9860,N_9242,N_9323);
nand U9861 (N_9861,N_9524,N_9721);
nor U9862 (N_9862,N_9488,N_9003);
or U9863 (N_9863,N_9380,N_9144);
nand U9864 (N_9864,N_9219,N_9463);
nand U9865 (N_9865,N_9104,N_9588);
and U9866 (N_9866,N_9358,N_9283);
nand U9867 (N_9867,N_9332,N_9630);
nor U9868 (N_9868,N_9139,N_9249);
xor U9869 (N_9869,N_9041,N_9388);
or U9870 (N_9870,N_9737,N_9162);
nor U9871 (N_9871,N_9129,N_9393);
and U9872 (N_9872,N_9542,N_9480);
nor U9873 (N_9873,N_9235,N_9703);
and U9874 (N_9874,N_9176,N_9100);
xor U9875 (N_9875,N_9238,N_9231);
or U9876 (N_9876,N_9567,N_9710);
nor U9877 (N_9877,N_9504,N_9590);
nand U9878 (N_9878,N_9227,N_9725);
nand U9879 (N_9879,N_9266,N_9500);
and U9880 (N_9880,N_9306,N_9482);
nand U9881 (N_9881,N_9623,N_9359);
xor U9882 (N_9882,N_9743,N_9185);
xor U9883 (N_9883,N_9247,N_9114);
xor U9884 (N_9884,N_9678,N_9441);
nor U9885 (N_9885,N_9018,N_9305);
or U9886 (N_9886,N_9550,N_9575);
xor U9887 (N_9887,N_9632,N_9468);
and U9888 (N_9888,N_9105,N_9128);
and U9889 (N_9889,N_9662,N_9212);
and U9890 (N_9890,N_9381,N_9216);
and U9891 (N_9891,N_9671,N_9713);
or U9892 (N_9892,N_9327,N_9154);
xnor U9893 (N_9893,N_9349,N_9165);
or U9894 (N_9894,N_9672,N_9591);
nor U9895 (N_9895,N_9557,N_9096);
or U9896 (N_9896,N_9051,N_9293);
xor U9897 (N_9897,N_9707,N_9159);
nor U9898 (N_9898,N_9255,N_9747);
xor U9899 (N_9899,N_9402,N_9319);
or U9900 (N_9900,N_9508,N_9053);
and U9901 (N_9901,N_9086,N_9704);
and U9902 (N_9902,N_9426,N_9220);
and U9903 (N_9903,N_9164,N_9715);
xor U9904 (N_9904,N_9712,N_9573);
and U9905 (N_9905,N_9261,N_9584);
or U9906 (N_9906,N_9206,N_9726);
xor U9907 (N_9907,N_9292,N_9617);
xnor U9908 (N_9908,N_9299,N_9364);
and U9909 (N_9909,N_9369,N_9090);
nor U9910 (N_9910,N_9580,N_9431);
nand U9911 (N_9911,N_9451,N_9690);
xor U9912 (N_9912,N_9276,N_9382);
xnor U9913 (N_9913,N_9728,N_9436);
xnor U9914 (N_9914,N_9495,N_9458);
nand U9915 (N_9915,N_9511,N_9409);
or U9916 (N_9916,N_9732,N_9635);
and U9917 (N_9917,N_9065,N_9531);
or U9918 (N_9918,N_9083,N_9518);
nor U9919 (N_9919,N_9628,N_9232);
or U9920 (N_9920,N_9626,N_9106);
or U9921 (N_9921,N_9666,N_9410);
xor U9922 (N_9922,N_9634,N_9304);
and U9923 (N_9923,N_9656,N_9325);
nand U9924 (N_9924,N_9735,N_9379);
and U9925 (N_9925,N_9681,N_9539);
and U9926 (N_9926,N_9194,N_9241);
or U9927 (N_9927,N_9621,N_9693);
xor U9928 (N_9928,N_9340,N_9587);
nor U9929 (N_9929,N_9126,N_9177);
xor U9930 (N_9930,N_9598,N_9191);
xor U9931 (N_9931,N_9166,N_9525);
nor U9932 (N_9932,N_9309,N_9395);
and U9933 (N_9933,N_9519,N_9318);
and U9934 (N_9934,N_9108,N_9199);
xnor U9935 (N_9935,N_9223,N_9296);
or U9936 (N_9936,N_9660,N_9320);
xor U9937 (N_9937,N_9568,N_9650);
nand U9938 (N_9938,N_9686,N_9391);
nor U9939 (N_9939,N_9471,N_9054);
xnor U9940 (N_9940,N_9494,N_9440);
or U9941 (N_9941,N_9658,N_9345);
xnor U9942 (N_9942,N_9610,N_9447);
xor U9943 (N_9943,N_9566,N_9700);
nand U9944 (N_9944,N_9736,N_9326);
nand U9945 (N_9945,N_9655,N_9520);
nand U9946 (N_9946,N_9435,N_9464);
xor U9947 (N_9947,N_9311,N_9178);
nor U9948 (N_9948,N_9067,N_9138);
and U9949 (N_9949,N_9274,N_9657);
xor U9950 (N_9950,N_9633,N_9043);
or U9951 (N_9951,N_9498,N_9312);
nor U9952 (N_9952,N_9558,N_9015);
nor U9953 (N_9953,N_9233,N_9708);
and U9954 (N_9954,N_9059,N_9143);
nand U9955 (N_9955,N_9057,N_9646);
and U9956 (N_9956,N_9688,N_9475);
xnor U9957 (N_9957,N_9085,N_9679);
or U9958 (N_9958,N_9609,N_9367);
or U9959 (N_9959,N_9614,N_9640);
nand U9960 (N_9960,N_9445,N_9510);
or U9961 (N_9961,N_9647,N_9645);
or U9962 (N_9962,N_9473,N_9596);
nand U9963 (N_9963,N_9727,N_9006);
nand U9964 (N_9964,N_9485,N_9502);
nor U9965 (N_9965,N_9592,N_9375);
xor U9966 (N_9966,N_9421,N_9063);
nand U9967 (N_9967,N_9411,N_9600);
or U9968 (N_9968,N_9084,N_9237);
and U9969 (N_9969,N_9078,N_9416);
xor U9970 (N_9970,N_9140,N_9720);
nand U9971 (N_9971,N_9239,N_9335);
nor U9972 (N_9972,N_9457,N_9272);
or U9973 (N_9973,N_9314,N_9636);
nor U9974 (N_9974,N_9111,N_9562);
nor U9975 (N_9975,N_9167,N_9394);
and U9976 (N_9976,N_9706,N_9418);
nand U9977 (N_9977,N_9071,N_9389);
nor U9978 (N_9978,N_9685,N_9284);
nor U9979 (N_9979,N_9270,N_9605);
or U9980 (N_9980,N_9072,N_9351);
nand U9981 (N_9981,N_9156,N_9210);
xnor U9982 (N_9982,N_9629,N_9014);
xor U9983 (N_9983,N_9360,N_9387);
xor U9984 (N_9984,N_9748,N_9438);
nand U9985 (N_9985,N_9300,N_9214);
xnor U9986 (N_9986,N_9442,N_9016);
nor U9987 (N_9987,N_9244,N_9627);
and U9988 (N_9988,N_9505,N_9115);
or U9989 (N_9989,N_9491,N_9022);
xor U9990 (N_9990,N_9082,N_9034);
or U9991 (N_9991,N_9417,N_9639);
nor U9992 (N_9992,N_9171,N_9192);
or U9993 (N_9993,N_9437,N_9058);
nor U9994 (N_9994,N_9091,N_9571);
and U9995 (N_9995,N_9055,N_9039);
nand U9996 (N_9996,N_9420,N_9378);
nand U9997 (N_9997,N_9352,N_9516);
and U9998 (N_9998,N_9342,N_9204);
nor U9999 (N_9999,N_9298,N_9257);
nor U10000 (N_10000,N_9372,N_9324);
or U10001 (N_10001,N_9234,N_9316);
and U10002 (N_10002,N_9033,N_9583);
nand U10003 (N_10003,N_9709,N_9537);
or U10004 (N_10004,N_9133,N_9076);
xor U10005 (N_10005,N_9330,N_9333);
nor U10006 (N_10006,N_9365,N_9275);
and U10007 (N_10007,N_9354,N_9746);
xor U10008 (N_10008,N_9745,N_9522);
nand U10009 (N_10009,N_9313,N_9399);
nor U10010 (N_10010,N_9131,N_9452);
nor U10011 (N_10011,N_9563,N_9268);
nand U10012 (N_10012,N_9064,N_9061);
xnor U10013 (N_10013,N_9386,N_9094);
and U10014 (N_10014,N_9186,N_9029);
and U10015 (N_10015,N_9484,N_9337);
or U10016 (N_10016,N_9092,N_9487);
nor U10017 (N_10017,N_9556,N_9684);
xnor U10018 (N_10018,N_9136,N_9263);
nand U10019 (N_10019,N_9163,N_9200);
or U10020 (N_10020,N_9079,N_9449);
nor U10021 (N_10021,N_9127,N_9328);
or U10022 (N_10022,N_9673,N_9478);
or U10023 (N_10023,N_9153,N_9663);
nor U10024 (N_10024,N_9229,N_9446);
xnor U10025 (N_10025,N_9552,N_9415);
or U10026 (N_10026,N_9182,N_9137);
or U10027 (N_10027,N_9269,N_9007);
nor U10028 (N_10028,N_9701,N_9667);
and U10029 (N_10029,N_9348,N_9017);
or U10030 (N_10030,N_9230,N_9215);
nand U10031 (N_10031,N_9277,N_9252);
and U10032 (N_10032,N_9308,N_9322);
and U10033 (N_10033,N_9425,N_9392);
or U10034 (N_10034,N_9490,N_9036);
and U10035 (N_10035,N_9135,N_9021);
and U10036 (N_10036,N_9160,N_9477);
xnor U10037 (N_10037,N_9141,N_9161);
and U10038 (N_10038,N_9528,N_9675);
xor U10039 (N_10039,N_9694,N_9208);
or U10040 (N_10040,N_9032,N_9260);
or U10041 (N_10041,N_9011,N_9718);
nand U10042 (N_10042,N_9547,N_9430);
xor U10043 (N_10043,N_9281,N_9472);
nand U10044 (N_10044,N_9374,N_9448);
xor U10045 (N_10045,N_9101,N_9532);
or U10046 (N_10046,N_9341,N_9559);
nand U10047 (N_10047,N_9148,N_9025);
and U10048 (N_10048,N_9336,N_9265);
xnor U10049 (N_10049,N_9698,N_9119);
and U10050 (N_10050,N_9030,N_9103);
nand U10051 (N_10051,N_9574,N_9060);
nand U10052 (N_10052,N_9439,N_9733);
xnor U10053 (N_10053,N_9211,N_9625);
and U10054 (N_10054,N_9074,N_9582);
xnor U10055 (N_10055,N_9669,N_9548);
or U10056 (N_10056,N_9218,N_9405);
or U10057 (N_10057,N_9113,N_9540);
xnor U10058 (N_10058,N_9116,N_9565);
nor U10059 (N_10059,N_9383,N_9044);
and U10060 (N_10060,N_9722,N_9373);
xnor U10061 (N_10061,N_9189,N_9012);
nand U10062 (N_10062,N_9196,N_9062);
nor U10063 (N_10063,N_9107,N_9172);
xor U10064 (N_10064,N_9121,N_9551);
xor U10065 (N_10065,N_9696,N_9124);
or U10066 (N_10066,N_9188,N_9664);
nand U10067 (N_10067,N_9334,N_9142);
xnor U10068 (N_10068,N_9474,N_9050);
nand U10069 (N_10069,N_9068,N_9280);
nor U10070 (N_10070,N_9273,N_9450);
nand U10071 (N_10071,N_9339,N_9040);
nor U10072 (N_10072,N_9676,N_9179);
nand U10073 (N_10073,N_9329,N_9258);
or U10074 (N_10074,N_9356,N_9175);
nor U10075 (N_10075,N_9615,N_9476);
or U10076 (N_10076,N_9607,N_9641);
or U10077 (N_10077,N_9117,N_9197);
and U10078 (N_10078,N_9008,N_9147);
or U10079 (N_10079,N_9271,N_9097);
nand U10080 (N_10080,N_9346,N_9256);
nand U10081 (N_10081,N_9170,N_9695);
xor U10082 (N_10082,N_9132,N_9423);
and U10083 (N_10083,N_9042,N_9174);
nor U10084 (N_10084,N_9744,N_9740);
xnor U10085 (N_10085,N_9499,N_9738);
nor U10086 (N_10086,N_9286,N_9052);
nor U10087 (N_10087,N_9444,N_9168);
and U10088 (N_10088,N_9048,N_9347);
nor U10089 (N_10089,N_9023,N_9134);
and U10090 (N_10090,N_9222,N_9618);
or U10091 (N_10091,N_9406,N_9228);
and U10092 (N_10092,N_9240,N_9597);
nand U10093 (N_10093,N_9724,N_9370);
nand U10094 (N_10094,N_9577,N_9202);
xor U10095 (N_10095,N_9151,N_9515);
nor U10096 (N_10096,N_9599,N_9638);
or U10097 (N_10097,N_9514,N_9601);
nor U10098 (N_10098,N_9123,N_9056);
xnor U10099 (N_10099,N_9716,N_9455);
or U10100 (N_10100,N_9027,N_9366);
or U10101 (N_10101,N_9523,N_9604);
and U10102 (N_10102,N_9545,N_9429);
xnor U10103 (N_10103,N_9549,N_9120);
nand U10104 (N_10104,N_9158,N_9602);
or U10105 (N_10105,N_9089,N_9668);
and U10106 (N_10106,N_9213,N_9019);
nor U10107 (N_10107,N_9643,N_9644);
nand U10108 (N_10108,N_9659,N_9250);
xnor U10109 (N_10109,N_9479,N_9046);
nor U10110 (N_10110,N_9099,N_9209);
and U10111 (N_10111,N_9248,N_9217);
and U10112 (N_10112,N_9413,N_9169);
or U10113 (N_10113,N_9536,N_9396);
xor U10114 (N_10114,N_9739,N_9088);
and U10115 (N_10115,N_9294,N_9243);
and U10116 (N_10116,N_9224,N_9198);
nand U10117 (N_10117,N_9002,N_9680);
nand U10118 (N_10118,N_9075,N_9705);
nand U10119 (N_10119,N_9711,N_9301);
and U10120 (N_10120,N_9109,N_9624);
or U10121 (N_10121,N_9028,N_9493);
xnor U10122 (N_10122,N_9385,N_9112);
nor U10123 (N_10123,N_9404,N_9589);
nor U10124 (N_10124,N_9408,N_9355);
xnor U10125 (N_10125,N_9065,N_9173);
xor U10126 (N_10126,N_9693,N_9138);
and U10127 (N_10127,N_9340,N_9617);
xnor U10128 (N_10128,N_9150,N_9558);
xnor U10129 (N_10129,N_9665,N_9029);
nand U10130 (N_10130,N_9742,N_9101);
or U10131 (N_10131,N_9061,N_9200);
or U10132 (N_10132,N_9603,N_9479);
or U10133 (N_10133,N_9427,N_9281);
nand U10134 (N_10134,N_9137,N_9708);
nor U10135 (N_10135,N_9370,N_9018);
or U10136 (N_10136,N_9305,N_9352);
and U10137 (N_10137,N_9005,N_9258);
xor U10138 (N_10138,N_9515,N_9739);
xnor U10139 (N_10139,N_9352,N_9452);
or U10140 (N_10140,N_9376,N_9323);
xnor U10141 (N_10141,N_9329,N_9121);
and U10142 (N_10142,N_9421,N_9227);
nor U10143 (N_10143,N_9242,N_9363);
xnor U10144 (N_10144,N_9231,N_9616);
xnor U10145 (N_10145,N_9519,N_9136);
nor U10146 (N_10146,N_9634,N_9363);
and U10147 (N_10147,N_9007,N_9312);
or U10148 (N_10148,N_9120,N_9244);
or U10149 (N_10149,N_9258,N_9641);
xnor U10150 (N_10150,N_9002,N_9418);
and U10151 (N_10151,N_9055,N_9279);
nand U10152 (N_10152,N_9495,N_9251);
or U10153 (N_10153,N_9683,N_9653);
xor U10154 (N_10154,N_9083,N_9597);
or U10155 (N_10155,N_9427,N_9724);
and U10156 (N_10156,N_9516,N_9317);
xnor U10157 (N_10157,N_9706,N_9653);
nand U10158 (N_10158,N_9031,N_9203);
nor U10159 (N_10159,N_9179,N_9086);
xor U10160 (N_10160,N_9594,N_9192);
nand U10161 (N_10161,N_9663,N_9731);
and U10162 (N_10162,N_9432,N_9620);
nand U10163 (N_10163,N_9299,N_9083);
nor U10164 (N_10164,N_9226,N_9749);
xnor U10165 (N_10165,N_9645,N_9101);
nand U10166 (N_10166,N_9661,N_9671);
xor U10167 (N_10167,N_9699,N_9678);
xnor U10168 (N_10168,N_9397,N_9233);
nor U10169 (N_10169,N_9694,N_9596);
and U10170 (N_10170,N_9228,N_9110);
or U10171 (N_10171,N_9571,N_9396);
nand U10172 (N_10172,N_9015,N_9379);
nand U10173 (N_10173,N_9605,N_9515);
nor U10174 (N_10174,N_9747,N_9442);
nor U10175 (N_10175,N_9659,N_9071);
and U10176 (N_10176,N_9459,N_9154);
nand U10177 (N_10177,N_9661,N_9637);
xor U10178 (N_10178,N_9112,N_9174);
or U10179 (N_10179,N_9049,N_9396);
nor U10180 (N_10180,N_9207,N_9256);
nand U10181 (N_10181,N_9567,N_9283);
nand U10182 (N_10182,N_9179,N_9722);
and U10183 (N_10183,N_9659,N_9019);
and U10184 (N_10184,N_9124,N_9123);
and U10185 (N_10185,N_9742,N_9064);
xnor U10186 (N_10186,N_9630,N_9472);
nor U10187 (N_10187,N_9208,N_9198);
nor U10188 (N_10188,N_9351,N_9187);
and U10189 (N_10189,N_9498,N_9011);
xor U10190 (N_10190,N_9295,N_9435);
nand U10191 (N_10191,N_9317,N_9439);
xnor U10192 (N_10192,N_9374,N_9596);
or U10193 (N_10193,N_9259,N_9705);
xnor U10194 (N_10194,N_9673,N_9525);
or U10195 (N_10195,N_9529,N_9305);
and U10196 (N_10196,N_9080,N_9159);
and U10197 (N_10197,N_9080,N_9025);
and U10198 (N_10198,N_9044,N_9176);
nor U10199 (N_10199,N_9614,N_9680);
nor U10200 (N_10200,N_9572,N_9257);
nor U10201 (N_10201,N_9053,N_9194);
and U10202 (N_10202,N_9652,N_9263);
xnor U10203 (N_10203,N_9251,N_9747);
and U10204 (N_10204,N_9450,N_9593);
or U10205 (N_10205,N_9262,N_9306);
nand U10206 (N_10206,N_9147,N_9037);
nand U10207 (N_10207,N_9539,N_9361);
and U10208 (N_10208,N_9173,N_9571);
nand U10209 (N_10209,N_9613,N_9112);
xor U10210 (N_10210,N_9279,N_9310);
or U10211 (N_10211,N_9486,N_9674);
or U10212 (N_10212,N_9378,N_9075);
xor U10213 (N_10213,N_9303,N_9158);
xor U10214 (N_10214,N_9448,N_9513);
nor U10215 (N_10215,N_9173,N_9177);
nor U10216 (N_10216,N_9106,N_9683);
nor U10217 (N_10217,N_9199,N_9196);
and U10218 (N_10218,N_9202,N_9748);
nor U10219 (N_10219,N_9496,N_9108);
nor U10220 (N_10220,N_9223,N_9587);
nor U10221 (N_10221,N_9712,N_9151);
and U10222 (N_10222,N_9732,N_9195);
nor U10223 (N_10223,N_9097,N_9606);
xor U10224 (N_10224,N_9721,N_9746);
or U10225 (N_10225,N_9414,N_9669);
nand U10226 (N_10226,N_9278,N_9519);
nand U10227 (N_10227,N_9733,N_9336);
xor U10228 (N_10228,N_9425,N_9653);
nor U10229 (N_10229,N_9240,N_9301);
or U10230 (N_10230,N_9466,N_9092);
or U10231 (N_10231,N_9455,N_9700);
and U10232 (N_10232,N_9124,N_9059);
and U10233 (N_10233,N_9338,N_9453);
or U10234 (N_10234,N_9286,N_9281);
xnor U10235 (N_10235,N_9176,N_9194);
or U10236 (N_10236,N_9515,N_9071);
or U10237 (N_10237,N_9574,N_9666);
or U10238 (N_10238,N_9099,N_9326);
or U10239 (N_10239,N_9426,N_9477);
nor U10240 (N_10240,N_9208,N_9320);
nand U10241 (N_10241,N_9651,N_9236);
and U10242 (N_10242,N_9199,N_9104);
or U10243 (N_10243,N_9483,N_9126);
nor U10244 (N_10244,N_9663,N_9567);
and U10245 (N_10245,N_9343,N_9011);
and U10246 (N_10246,N_9339,N_9542);
or U10247 (N_10247,N_9261,N_9349);
xor U10248 (N_10248,N_9697,N_9084);
and U10249 (N_10249,N_9225,N_9414);
nor U10250 (N_10250,N_9660,N_9369);
xnor U10251 (N_10251,N_9645,N_9061);
xnor U10252 (N_10252,N_9074,N_9065);
and U10253 (N_10253,N_9575,N_9177);
nand U10254 (N_10254,N_9618,N_9522);
and U10255 (N_10255,N_9412,N_9663);
xnor U10256 (N_10256,N_9580,N_9717);
xnor U10257 (N_10257,N_9003,N_9265);
and U10258 (N_10258,N_9195,N_9640);
xor U10259 (N_10259,N_9591,N_9600);
xnor U10260 (N_10260,N_9216,N_9322);
and U10261 (N_10261,N_9153,N_9111);
nand U10262 (N_10262,N_9603,N_9720);
xnor U10263 (N_10263,N_9357,N_9562);
and U10264 (N_10264,N_9042,N_9101);
or U10265 (N_10265,N_9227,N_9635);
xor U10266 (N_10266,N_9467,N_9149);
xnor U10267 (N_10267,N_9014,N_9527);
and U10268 (N_10268,N_9218,N_9287);
nor U10269 (N_10269,N_9681,N_9488);
xnor U10270 (N_10270,N_9030,N_9291);
nor U10271 (N_10271,N_9422,N_9674);
or U10272 (N_10272,N_9088,N_9010);
xor U10273 (N_10273,N_9326,N_9258);
or U10274 (N_10274,N_9183,N_9424);
xnor U10275 (N_10275,N_9122,N_9697);
nand U10276 (N_10276,N_9714,N_9379);
or U10277 (N_10277,N_9460,N_9163);
and U10278 (N_10278,N_9163,N_9330);
nor U10279 (N_10279,N_9176,N_9380);
nand U10280 (N_10280,N_9294,N_9698);
nor U10281 (N_10281,N_9102,N_9262);
xor U10282 (N_10282,N_9429,N_9696);
xor U10283 (N_10283,N_9001,N_9469);
or U10284 (N_10284,N_9404,N_9087);
xor U10285 (N_10285,N_9130,N_9685);
xor U10286 (N_10286,N_9225,N_9322);
nand U10287 (N_10287,N_9079,N_9250);
nor U10288 (N_10288,N_9075,N_9348);
nand U10289 (N_10289,N_9648,N_9654);
or U10290 (N_10290,N_9348,N_9230);
nor U10291 (N_10291,N_9610,N_9291);
and U10292 (N_10292,N_9731,N_9253);
xnor U10293 (N_10293,N_9097,N_9039);
nand U10294 (N_10294,N_9301,N_9062);
and U10295 (N_10295,N_9538,N_9389);
or U10296 (N_10296,N_9641,N_9741);
and U10297 (N_10297,N_9206,N_9483);
xnor U10298 (N_10298,N_9057,N_9231);
xnor U10299 (N_10299,N_9727,N_9738);
xor U10300 (N_10300,N_9554,N_9497);
nor U10301 (N_10301,N_9417,N_9273);
and U10302 (N_10302,N_9145,N_9455);
nand U10303 (N_10303,N_9156,N_9115);
or U10304 (N_10304,N_9027,N_9509);
or U10305 (N_10305,N_9561,N_9286);
xnor U10306 (N_10306,N_9573,N_9371);
nand U10307 (N_10307,N_9296,N_9092);
nor U10308 (N_10308,N_9634,N_9658);
nor U10309 (N_10309,N_9562,N_9567);
and U10310 (N_10310,N_9330,N_9685);
nand U10311 (N_10311,N_9506,N_9345);
nor U10312 (N_10312,N_9473,N_9006);
xor U10313 (N_10313,N_9741,N_9512);
and U10314 (N_10314,N_9014,N_9271);
or U10315 (N_10315,N_9210,N_9297);
nand U10316 (N_10316,N_9304,N_9200);
xor U10317 (N_10317,N_9210,N_9657);
xor U10318 (N_10318,N_9591,N_9616);
and U10319 (N_10319,N_9161,N_9631);
or U10320 (N_10320,N_9235,N_9008);
xor U10321 (N_10321,N_9418,N_9388);
nand U10322 (N_10322,N_9668,N_9519);
nor U10323 (N_10323,N_9165,N_9491);
nor U10324 (N_10324,N_9667,N_9157);
nand U10325 (N_10325,N_9348,N_9126);
xor U10326 (N_10326,N_9533,N_9030);
nand U10327 (N_10327,N_9670,N_9572);
nand U10328 (N_10328,N_9687,N_9348);
nand U10329 (N_10329,N_9434,N_9618);
nor U10330 (N_10330,N_9367,N_9047);
nand U10331 (N_10331,N_9426,N_9659);
or U10332 (N_10332,N_9738,N_9547);
nand U10333 (N_10333,N_9613,N_9296);
nor U10334 (N_10334,N_9720,N_9349);
nor U10335 (N_10335,N_9550,N_9691);
or U10336 (N_10336,N_9472,N_9136);
and U10337 (N_10337,N_9402,N_9691);
nand U10338 (N_10338,N_9320,N_9238);
or U10339 (N_10339,N_9316,N_9221);
or U10340 (N_10340,N_9691,N_9638);
nand U10341 (N_10341,N_9192,N_9705);
or U10342 (N_10342,N_9238,N_9465);
and U10343 (N_10343,N_9104,N_9490);
nor U10344 (N_10344,N_9414,N_9066);
nor U10345 (N_10345,N_9143,N_9190);
or U10346 (N_10346,N_9484,N_9594);
xnor U10347 (N_10347,N_9060,N_9316);
or U10348 (N_10348,N_9074,N_9457);
xnor U10349 (N_10349,N_9184,N_9009);
or U10350 (N_10350,N_9050,N_9648);
nand U10351 (N_10351,N_9420,N_9374);
and U10352 (N_10352,N_9705,N_9066);
and U10353 (N_10353,N_9518,N_9392);
nor U10354 (N_10354,N_9461,N_9618);
or U10355 (N_10355,N_9370,N_9218);
or U10356 (N_10356,N_9491,N_9589);
xnor U10357 (N_10357,N_9074,N_9593);
or U10358 (N_10358,N_9639,N_9266);
nor U10359 (N_10359,N_9132,N_9347);
nand U10360 (N_10360,N_9439,N_9229);
and U10361 (N_10361,N_9658,N_9045);
xor U10362 (N_10362,N_9270,N_9355);
xnor U10363 (N_10363,N_9583,N_9171);
nand U10364 (N_10364,N_9649,N_9416);
xor U10365 (N_10365,N_9237,N_9581);
nor U10366 (N_10366,N_9014,N_9555);
xnor U10367 (N_10367,N_9290,N_9286);
nand U10368 (N_10368,N_9052,N_9253);
nand U10369 (N_10369,N_9078,N_9338);
or U10370 (N_10370,N_9672,N_9708);
nand U10371 (N_10371,N_9366,N_9014);
and U10372 (N_10372,N_9323,N_9475);
nand U10373 (N_10373,N_9279,N_9101);
nor U10374 (N_10374,N_9243,N_9592);
or U10375 (N_10375,N_9204,N_9123);
and U10376 (N_10376,N_9661,N_9669);
nor U10377 (N_10377,N_9180,N_9471);
nor U10378 (N_10378,N_9183,N_9157);
xnor U10379 (N_10379,N_9541,N_9233);
or U10380 (N_10380,N_9075,N_9061);
xnor U10381 (N_10381,N_9378,N_9564);
nand U10382 (N_10382,N_9735,N_9336);
nand U10383 (N_10383,N_9286,N_9360);
xnor U10384 (N_10384,N_9688,N_9257);
nand U10385 (N_10385,N_9180,N_9051);
xnor U10386 (N_10386,N_9519,N_9191);
nand U10387 (N_10387,N_9612,N_9017);
and U10388 (N_10388,N_9195,N_9288);
or U10389 (N_10389,N_9398,N_9415);
nand U10390 (N_10390,N_9188,N_9335);
nor U10391 (N_10391,N_9440,N_9633);
or U10392 (N_10392,N_9652,N_9410);
nand U10393 (N_10393,N_9273,N_9568);
or U10394 (N_10394,N_9310,N_9376);
and U10395 (N_10395,N_9417,N_9210);
xor U10396 (N_10396,N_9611,N_9675);
xnor U10397 (N_10397,N_9360,N_9053);
and U10398 (N_10398,N_9483,N_9323);
xor U10399 (N_10399,N_9566,N_9697);
nand U10400 (N_10400,N_9679,N_9512);
or U10401 (N_10401,N_9716,N_9517);
and U10402 (N_10402,N_9022,N_9462);
xor U10403 (N_10403,N_9174,N_9477);
xnor U10404 (N_10404,N_9523,N_9199);
nand U10405 (N_10405,N_9426,N_9215);
xnor U10406 (N_10406,N_9351,N_9160);
nor U10407 (N_10407,N_9185,N_9284);
nand U10408 (N_10408,N_9548,N_9362);
xnor U10409 (N_10409,N_9609,N_9113);
or U10410 (N_10410,N_9387,N_9697);
or U10411 (N_10411,N_9031,N_9731);
nor U10412 (N_10412,N_9249,N_9439);
and U10413 (N_10413,N_9014,N_9318);
xnor U10414 (N_10414,N_9598,N_9374);
xor U10415 (N_10415,N_9308,N_9258);
nand U10416 (N_10416,N_9197,N_9591);
or U10417 (N_10417,N_9680,N_9664);
nand U10418 (N_10418,N_9632,N_9408);
and U10419 (N_10419,N_9314,N_9749);
nor U10420 (N_10420,N_9491,N_9502);
nand U10421 (N_10421,N_9586,N_9463);
and U10422 (N_10422,N_9108,N_9484);
xnor U10423 (N_10423,N_9538,N_9087);
or U10424 (N_10424,N_9486,N_9485);
and U10425 (N_10425,N_9123,N_9555);
nor U10426 (N_10426,N_9367,N_9081);
nor U10427 (N_10427,N_9610,N_9590);
xor U10428 (N_10428,N_9470,N_9703);
or U10429 (N_10429,N_9563,N_9116);
or U10430 (N_10430,N_9328,N_9511);
nor U10431 (N_10431,N_9076,N_9226);
nand U10432 (N_10432,N_9310,N_9389);
or U10433 (N_10433,N_9652,N_9047);
and U10434 (N_10434,N_9607,N_9156);
nor U10435 (N_10435,N_9466,N_9081);
or U10436 (N_10436,N_9255,N_9015);
nor U10437 (N_10437,N_9208,N_9446);
or U10438 (N_10438,N_9599,N_9006);
xor U10439 (N_10439,N_9353,N_9503);
and U10440 (N_10440,N_9541,N_9738);
xor U10441 (N_10441,N_9469,N_9563);
nor U10442 (N_10442,N_9301,N_9031);
or U10443 (N_10443,N_9395,N_9311);
nand U10444 (N_10444,N_9649,N_9683);
nor U10445 (N_10445,N_9155,N_9044);
or U10446 (N_10446,N_9272,N_9505);
nand U10447 (N_10447,N_9167,N_9329);
nand U10448 (N_10448,N_9306,N_9252);
and U10449 (N_10449,N_9017,N_9699);
nor U10450 (N_10450,N_9373,N_9066);
and U10451 (N_10451,N_9040,N_9235);
or U10452 (N_10452,N_9166,N_9328);
nand U10453 (N_10453,N_9677,N_9641);
nand U10454 (N_10454,N_9396,N_9012);
xor U10455 (N_10455,N_9205,N_9434);
nor U10456 (N_10456,N_9161,N_9733);
nand U10457 (N_10457,N_9385,N_9152);
nor U10458 (N_10458,N_9259,N_9297);
nand U10459 (N_10459,N_9608,N_9453);
nand U10460 (N_10460,N_9502,N_9114);
or U10461 (N_10461,N_9326,N_9406);
or U10462 (N_10462,N_9305,N_9206);
and U10463 (N_10463,N_9266,N_9008);
nor U10464 (N_10464,N_9718,N_9027);
and U10465 (N_10465,N_9443,N_9071);
and U10466 (N_10466,N_9188,N_9005);
or U10467 (N_10467,N_9026,N_9051);
and U10468 (N_10468,N_9713,N_9670);
xnor U10469 (N_10469,N_9542,N_9386);
nor U10470 (N_10470,N_9444,N_9587);
nand U10471 (N_10471,N_9093,N_9228);
xor U10472 (N_10472,N_9254,N_9050);
nand U10473 (N_10473,N_9123,N_9291);
or U10474 (N_10474,N_9081,N_9187);
nor U10475 (N_10475,N_9060,N_9566);
or U10476 (N_10476,N_9395,N_9467);
xor U10477 (N_10477,N_9749,N_9129);
and U10478 (N_10478,N_9572,N_9664);
and U10479 (N_10479,N_9429,N_9662);
nand U10480 (N_10480,N_9744,N_9544);
or U10481 (N_10481,N_9406,N_9394);
xor U10482 (N_10482,N_9630,N_9245);
nor U10483 (N_10483,N_9509,N_9183);
or U10484 (N_10484,N_9365,N_9422);
nand U10485 (N_10485,N_9162,N_9448);
nand U10486 (N_10486,N_9108,N_9446);
and U10487 (N_10487,N_9320,N_9393);
or U10488 (N_10488,N_9053,N_9290);
or U10489 (N_10489,N_9667,N_9630);
xor U10490 (N_10490,N_9068,N_9414);
nand U10491 (N_10491,N_9142,N_9239);
xor U10492 (N_10492,N_9571,N_9100);
and U10493 (N_10493,N_9653,N_9151);
nor U10494 (N_10494,N_9598,N_9203);
and U10495 (N_10495,N_9107,N_9320);
nand U10496 (N_10496,N_9725,N_9259);
and U10497 (N_10497,N_9733,N_9109);
nand U10498 (N_10498,N_9273,N_9726);
nand U10499 (N_10499,N_9649,N_9268);
nand U10500 (N_10500,N_10260,N_9986);
xor U10501 (N_10501,N_10008,N_10407);
nor U10502 (N_10502,N_10478,N_9908);
or U10503 (N_10503,N_10014,N_10452);
nor U10504 (N_10504,N_10042,N_9999);
nand U10505 (N_10505,N_10132,N_10438);
and U10506 (N_10506,N_10290,N_10301);
and U10507 (N_10507,N_9782,N_9778);
nand U10508 (N_10508,N_10027,N_9849);
nor U10509 (N_10509,N_9967,N_10375);
and U10510 (N_10510,N_9913,N_10076);
nor U10511 (N_10511,N_10275,N_9870);
or U10512 (N_10512,N_10335,N_10491);
xnor U10513 (N_10513,N_9906,N_10310);
and U10514 (N_10514,N_10095,N_10046);
and U10515 (N_10515,N_10123,N_10230);
or U10516 (N_10516,N_10493,N_9979);
nor U10517 (N_10517,N_10168,N_10462);
nand U10518 (N_10518,N_9803,N_10268);
xnor U10519 (N_10519,N_10271,N_10108);
and U10520 (N_10520,N_9788,N_10004);
and U10521 (N_10521,N_10136,N_9785);
xnor U10522 (N_10522,N_10079,N_10228);
and U10523 (N_10523,N_9973,N_9848);
nand U10524 (N_10524,N_10190,N_10466);
xor U10525 (N_10525,N_9872,N_10278);
and U10526 (N_10526,N_9757,N_10455);
nand U10527 (N_10527,N_9857,N_10364);
xnor U10528 (N_10528,N_9793,N_10017);
or U10529 (N_10529,N_10142,N_10380);
xor U10530 (N_10530,N_10378,N_10138);
and U10531 (N_10531,N_9750,N_10128);
nand U10532 (N_10532,N_9844,N_10224);
and U10533 (N_10533,N_10070,N_10351);
or U10534 (N_10534,N_10253,N_10330);
xnor U10535 (N_10535,N_10398,N_10463);
and U10536 (N_10536,N_9985,N_10294);
and U10537 (N_10537,N_10293,N_10329);
xnor U10538 (N_10538,N_9899,N_9809);
nand U10539 (N_10539,N_9981,N_9772);
or U10540 (N_10540,N_9806,N_9812);
nand U10541 (N_10541,N_10192,N_9847);
and U10542 (N_10542,N_10146,N_10379);
nor U10543 (N_10543,N_10337,N_10482);
nand U10544 (N_10544,N_10494,N_10053);
nand U10545 (N_10545,N_10133,N_9895);
xnor U10546 (N_10546,N_10216,N_9992);
or U10547 (N_10547,N_10475,N_10169);
and U10548 (N_10548,N_10412,N_10094);
nand U10549 (N_10549,N_9987,N_10194);
xor U10550 (N_10550,N_10198,N_9794);
or U10551 (N_10551,N_10434,N_10113);
xnor U10552 (N_10552,N_9827,N_10315);
nor U10553 (N_10553,N_10317,N_10266);
nand U10554 (N_10554,N_10000,N_10325);
xor U10555 (N_10555,N_9854,N_9762);
xnor U10556 (N_10556,N_10223,N_10498);
xor U10557 (N_10557,N_10087,N_9774);
or U10558 (N_10558,N_9903,N_10387);
nand U10559 (N_10559,N_9896,N_9960);
and U10560 (N_10560,N_10456,N_10339);
xnor U10561 (N_10561,N_10229,N_9842);
and U10562 (N_10562,N_10469,N_9755);
or U10563 (N_10563,N_10492,N_10165);
or U10564 (N_10564,N_9974,N_10060);
and U10565 (N_10565,N_10088,N_10083);
nor U10566 (N_10566,N_9819,N_9931);
nand U10567 (N_10567,N_10447,N_10450);
xor U10568 (N_10568,N_10200,N_10309);
and U10569 (N_10569,N_10304,N_10013);
nor U10570 (N_10570,N_10193,N_9881);
xor U10571 (N_10571,N_10362,N_9802);
nand U10572 (N_10572,N_9947,N_9892);
nand U10573 (N_10573,N_10306,N_9882);
nor U10574 (N_10574,N_10020,N_10195);
nand U10575 (N_10575,N_10054,N_10189);
nand U10576 (N_10576,N_9816,N_9996);
and U10577 (N_10577,N_9912,N_10263);
or U10578 (N_10578,N_10383,N_9949);
nor U10579 (N_10579,N_10018,N_10065);
nand U10580 (N_10580,N_10444,N_9972);
or U10581 (N_10581,N_9759,N_10257);
xor U10582 (N_10582,N_9765,N_9889);
nor U10583 (N_10583,N_10041,N_10361);
nor U10584 (N_10584,N_10365,N_9826);
nor U10585 (N_10585,N_10350,N_9907);
or U10586 (N_10586,N_10021,N_10439);
and U10587 (N_10587,N_9898,N_10384);
or U10588 (N_10588,N_9779,N_9952);
or U10589 (N_10589,N_9904,N_9926);
or U10590 (N_10590,N_10254,N_10114);
xor U10591 (N_10591,N_10471,N_9879);
xor U10592 (N_10592,N_10394,N_10396);
nand U10593 (N_10593,N_9971,N_10432);
xnor U10594 (N_10594,N_10321,N_10148);
and U10595 (N_10595,N_10279,N_10281);
xor U10596 (N_10596,N_10484,N_10343);
xor U10597 (N_10597,N_9954,N_9958);
or U10598 (N_10598,N_10286,N_10251);
xor U10599 (N_10599,N_10062,N_10417);
xnor U10600 (N_10600,N_10319,N_9829);
nand U10601 (N_10601,N_10163,N_10269);
and U10602 (N_10602,N_10404,N_10393);
nand U10603 (N_10603,N_10073,N_9814);
or U10604 (N_10604,N_10408,N_10116);
xnor U10605 (N_10605,N_10388,N_10043);
xor U10606 (N_10606,N_9841,N_9965);
nand U10607 (N_10607,N_10451,N_10037);
xor U10608 (N_10608,N_10097,N_10061);
and U10609 (N_10609,N_10429,N_10006);
xor U10610 (N_10610,N_10187,N_9911);
and U10611 (N_10611,N_10312,N_9970);
and U10612 (N_10612,N_9957,N_10352);
or U10613 (N_10613,N_10129,N_10208);
or U10614 (N_10614,N_10121,N_10231);
nor U10615 (N_10615,N_10063,N_10363);
xnor U10616 (N_10616,N_10401,N_10299);
or U10617 (N_10617,N_10497,N_10470);
nor U10618 (N_10618,N_10259,N_10340);
nand U10619 (N_10619,N_10080,N_9810);
and U10620 (N_10620,N_10485,N_10139);
xnor U10621 (N_10621,N_10209,N_9867);
xnor U10622 (N_10622,N_10022,N_10460);
or U10623 (N_10623,N_10219,N_10256);
or U10624 (N_10624,N_9866,N_10112);
xnor U10625 (N_10625,N_9858,N_10207);
or U10626 (N_10626,N_9832,N_9835);
nor U10627 (N_10627,N_9871,N_10454);
nand U10628 (N_10628,N_10298,N_9824);
xor U10629 (N_10629,N_10346,N_9876);
nor U10630 (N_10630,N_10488,N_10127);
nand U10631 (N_10631,N_10368,N_10151);
nand U10632 (N_10632,N_9860,N_9886);
nor U10633 (N_10633,N_9766,N_10156);
or U10634 (N_10634,N_10249,N_10089);
nand U10635 (N_10635,N_10496,N_10359);
or U10636 (N_10636,N_10201,N_10184);
nand U10637 (N_10637,N_9781,N_10025);
xnor U10638 (N_10638,N_10377,N_10218);
nor U10639 (N_10639,N_10490,N_10212);
xor U10640 (N_10640,N_10068,N_10177);
nand U10641 (N_10641,N_10110,N_10464);
or U10642 (N_10642,N_10173,N_10395);
and U10643 (N_10643,N_9787,N_9840);
xnor U10644 (N_10644,N_10420,N_10446);
xor U10645 (N_10645,N_10338,N_10180);
nor U10646 (N_10646,N_10308,N_10082);
nor U10647 (N_10647,N_10360,N_9888);
nor U10648 (N_10648,N_9894,N_10430);
or U10649 (N_10649,N_10399,N_9795);
nand U10650 (N_10650,N_9846,N_10238);
nor U10651 (N_10651,N_9838,N_10039);
xnor U10652 (N_10652,N_10433,N_10214);
nand U10653 (N_10653,N_9820,N_9828);
and U10654 (N_10654,N_10390,N_10186);
and U10655 (N_10655,N_9964,N_10191);
nor U10656 (N_10656,N_9837,N_10235);
or U10657 (N_10657,N_10411,N_9796);
nand U10658 (N_10658,N_10197,N_9789);
and U10659 (N_10659,N_10034,N_9804);
or U10660 (N_10660,N_10147,N_10314);
nand U10661 (N_10661,N_9993,N_10001);
or U10662 (N_10662,N_10406,N_9968);
and U10663 (N_10663,N_10242,N_10204);
or U10664 (N_10664,N_10481,N_9786);
nor U10665 (N_10665,N_9753,N_10373);
nand U10666 (N_10666,N_10009,N_9900);
and U10667 (N_10667,N_10160,N_10067);
and U10668 (N_10668,N_10047,N_10426);
nor U10669 (N_10669,N_10239,N_10016);
or U10670 (N_10670,N_10297,N_9760);
xor U10671 (N_10671,N_10442,N_10284);
xor U10672 (N_10672,N_9885,N_10495);
nor U10673 (N_10673,N_9831,N_10178);
nand U10674 (N_10674,N_10479,N_10487);
or U10675 (N_10675,N_10175,N_9764);
or U10676 (N_10676,N_10354,N_10057);
nor U10677 (N_10677,N_9761,N_10171);
or U10678 (N_10678,N_10099,N_9792);
nand U10679 (N_10679,N_10386,N_10038);
nand U10680 (N_10680,N_10149,N_10066);
nor U10681 (N_10681,N_10422,N_10296);
nand U10682 (N_10682,N_10154,N_9982);
and U10683 (N_10683,N_9752,N_9853);
nand U10684 (N_10684,N_10084,N_10358);
and U10685 (N_10685,N_10369,N_10283);
nor U10686 (N_10686,N_10344,N_10115);
nor U10687 (N_10687,N_10106,N_10353);
nor U10688 (N_10688,N_9918,N_10276);
xor U10689 (N_10689,N_9945,N_9777);
nand U10690 (N_10690,N_9877,N_10356);
and U10691 (N_10691,N_9843,N_9943);
and U10692 (N_10692,N_10236,N_9955);
xor U10693 (N_10693,N_10174,N_10250);
and U10694 (N_10694,N_10397,N_10044);
and U10695 (N_10695,N_10262,N_10248);
nand U10696 (N_10696,N_9998,N_9950);
nor U10697 (N_10697,N_10217,N_10213);
or U10698 (N_10698,N_10300,N_9869);
and U10699 (N_10699,N_10141,N_10311);
and U10700 (N_10700,N_9935,N_10179);
xor U10701 (N_10701,N_10188,N_10024);
nand U10702 (N_10702,N_9780,N_10252);
xor U10703 (N_10703,N_9799,N_10211);
nor U10704 (N_10704,N_10367,N_10313);
xnor U10705 (N_10705,N_10226,N_10414);
nand U10706 (N_10706,N_9916,N_10125);
and U10707 (N_10707,N_10155,N_10270);
and U10708 (N_10708,N_10202,N_9914);
nand U10709 (N_10709,N_10458,N_9976);
nor U10710 (N_10710,N_10222,N_9944);
xor U10711 (N_10711,N_9934,N_9769);
nand U10712 (N_10712,N_10476,N_9990);
xor U10713 (N_10713,N_10145,N_9901);
nand U10714 (N_10714,N_9887,N_10302);
nor U10715 (N_10715,N_10424,N_9938);
or U10716 (N_10716,N_10258,N_10483);
nand U10717 (N_10717,N_9845,N_9797);
nor U10718 (N_10718,N_9927,N_10445);
nand U10719 (N_10719,N_9818,N_9771);
and U10720 (N_10720,N_9875,N_10419);
xnor U10721 (N_10721,N_9991,N_9798);
and U10722 (N_10722,N_10091,N_9800);
xor U10723 (N_10723,N_9989,N_9917);
xor U10724 (N_10724,N_10400,N_9836);
and U10725 (N_10725,N_9963,N_9983);
and U10726 (N_10726,N_10077,N_10051);
or U10727 (N_10727,N_10413,N_10333);
nor U10728 (N_10728,N_9940,N_10028);
nand U10729 (N_10729,N_10093,N_10135);
or U10730 (N_10730,N_9924,N_10489);
nand U10731 (N_10731,N_10172,N_9997);
nand U10732 (N_10732,N_10237,N_10410);
nor U10733 (N_10733,N_9851,N_9984);
or U10734 (N_10734,N_10161,N_10227);
nand U10735 (N_10735,N_10117,N_10098);
nor U10736 (N_10736,N_10241,N_9905);
xor U10737 (N_10737,N_10288,N_10324);
and U10738 (N_10738,N_9776,N_10280);
or U10739 (N_10739,N_10389,N_10030);
nand U10740 (N_10740,N_10264,N_9852);
nand U10741 (N_10741,N_10265,N_10307);
and U10742 (N_10742,N_10150,N_9897);
nand U10743 (N_10743,N_9859,N_9808);
or U10744 (N_10744,N_10182,N_10245);
nand U10745 (N_10745,N_10111,N_10103);
or U10746 (N_10746,N_9856,N_10385);
or U10747 (N_10747,N_9756,N_9988);
or U10748 (N_10748,N_10273,N_9770);
xnor U10749 (N_10749,N_10240,N_10015);
xnor U10750 (N_10750,N_10255,N_9929);
nor U10751 (N_10751,N_9763,N_9839);
nand U10752 (N_10752,N_10465,N_9891);
or U10753 (N_10753,N_10272,N_10473);
or U10754 (N_10754,N_9790,N_10261);
nor U10755 (N_10755,N_9953,N_10345);
nor U10756 (N_10756,N_9884,N_9937);
nor U10757 (N_10757,N_10316,N_9805);
nor U10758 (N_10758,N_10480,N_9959);
nand U10759 (N_10759,N_9948,N_9966);
xor U10760 (N_10760,N_10423,N_9933);
and U10761 (N_10761,N_10347,N_10437);
nand U10762 (N_10762,N_10167,N_9930);
or U10763 (N_10763,N_10243,N_10436);
xnor U10764 (N_10764,N_9920,N_10085);
nor U10765 (N_10765,N_10292,N_9822);
or U10766 (N_10766,N_10031,N_9880);
nand U10767 (N_10767,N_10105,N_10382);
or U10768 (N_10768,N_9823,N_10049);
nor U10769 (N_10769,N_10421,N_10233);
nand U10770 (N_10770,N_10035,N_10327);
nor U10771 (N_10771,N_10040,N_10320);
or U10772 (N_10772,N_9923,N_9863);
xnor U10773 (N_10773,N_9833,N_10086);
and U10774 (N_10774,N_10104,N_10234);
xnor U10775 (N_10775,N_9942,N_10048);
nor U10776 (N_10776,N_10277,N_10164);
xnor U10777 (N_10777,N_10402,N_9868);
and U10778 (N_10778,N_10152,N_9773);
nor U10779 (N_10779,N_10459,N_10431);
xor U10780 (N_10780,N_10303,N_9834);
nor U10781 (N_10781,N_10205,N_10059);
xor U10782 (N_10782,N_10246,N_10232);
xor U10783 (N_10783,N_9994,N_9830);
and U10784 (N_10784,N_9921,N_9815);
xor U10785 (N_10785,N_10331,N_10120);
nand U10786 (N_10786,N_10472,N_10181);
nand U10787 (N_10787,N_10416,N_10050);
and U10788 (N_10788,N_9791,N_10341);
xnor U10789 (N_10789,N_10029,N_10159);
nor U10790 (N_10790,N_10427,N_9962);
nand U10791 (N_10791,N_10449,N_10074);
nand U10792 (N_10792,N_9951,N_9801);
nand U10793 (N_10793,N_10371,N_10247);
xnor U10794 (N_10794,N_10357,N_10348);
or U10795 (N_10795,N_10033,N_9925);
xnor U10796 (N_10796,N_10267,N_10334);
and U10797 (N_10797,N_10244,N_10477);
xnor U10798 (N_10798,N_10055,N_9767);
nand U10799 (N_10799,N_10376,N_9807);
nand U10800 (N_10800,N_10326,N_10295);
nor U10801 (N_10801,N_9936,N_10019);
nor U10802 (N_10802,N_9865,N_10032);
and U10803 (N_10803,N_10131,N_10403);
nor U10804 (N_10804,N_10162,N_10101);
xnor U10805 (N_10805,N_10441,N_10096);
nor U10806 (N_10806,N_10372,N_10210);
nand U10807 (N_10807,N_10349,N_10109);
nand U10808 (N_10808,N_10415,N_10287);
nor U10809 (N_10809,N_10342,N_10468);
xor U10810 (N_10810,N_10428,N_10289);
or U10811 (N_10811,N_10448,N_10305);
and U10812 (N_10812,N_10323,N_10140);
nor U10813 (N_10813,N_9939,N_10090);
nand U10814 (N_10814,N_9821,N_10100);
nand U10815 (N_10815,N_9817,N_9775);
nor U10816 (N_10816,N_10392,N_10185);
and U10817 (N_10817,N_10036,N_10143);
or U10818 (N_10818,N_9873,N_9977);
xnor U10819 (N_10819,N_10005,N_9754);
xnor U10820 (N_10820,N_10072,N_10203);
xnor U10821 (N_10821,N_10130,N_10023);
nand U10822 (N_10822,N_9975,N_10045);
or U10823 (N_10823,N_9751,N_9878);
nand U10824 (N_10824,N_9813,N_10075);
and U10825 (N_10825,N_10206,N_10370);
xor U10826 (N_10826,N_10069,N_10467);
or U10827 (N_10827,N_10078,N_10119);
and U10828 (N_10828,N_9928,N_10010);
xnor U10829 (N_10829,N_9783,N_9915);
nand U10830 (N_10830,N_10107,N_10012);
or U10831 (N_10831,N_10064,N_10405);
and U10832 (N_10832,N_10011,N_10332);
nand U10833 (N_10833,N_10126,N_10285);
nor U10834 (N_10834,N_10443,N_10409);
xnor U10835 (N_10835,N_9864,N_10225);
or U10836 (N_10836,N_10282,N_10355);
xor U10837 (N_10837,N_9861,N_10158);
nand U10838 (N_10838,N_10052,N_10081);
nand U10839 (N_10839,N_10425,N_9919);
nand U10840 (N_10840,N_9978,N_10102);
or U10841 (N_10841,N_10220,N_10440);
and U10842 (N_10842,N_9961,N_10381);
or U10843 (N_10843,N_10007,N_10092);
or U10844 (N_10844,N_9909,N_10071);
or U10845 (N_10845,N_9850,N_10453);
xor U10846 (N_10846,N_9893,N_10056);
and U10847 (N_10847,N_10274,N_9956);
nor U10848 (N_10848,N_9902,N_10144);
xnor U10849 (N_10849,N_10166,N_9890);
and U10850 (N_10850,N_10457,N_10058);
and U10851 (N_10851,N_9784,N_10176);
nor U10852 (N_10852,N_9910,N_9941);
xor U10853 (N_10853,N_9758,N_10199);
xnor U10854 (N_10854,N_10124,N_9825);
or U10855 (N_10855,N_10153,N_10026);
xor U10856 (N_10856,N_10391,N_10122);
and U10857 (N_10857,N_10499,N_9811);
or U10858 (N_10858,N_10318,N_10374);
and U10859 (N_10859,N_10474,N_10328);
nor U10860 (N_10860,N_9922,N_9932);
or U10861 (N_10861,N_9862,N_10170);
xnor U10862 (N_10862,N_10002,N_10435);
nand U10863 (N_10863,N_10215,N_10137);
nor U10864 (N_10864,N_10291,N_9995);
nor U10865 (N_10865,N_9969,N_9768);
and U10866 (N_10866,N_10221,N_10366);
xor U10867 (N_10867,N_10336,N_10134);
xnor U10868 (N_10868,N_10418,N_10461);
or U10869 (N_10869,N_9874,N_10183);
or U10870 (N_10870,N_10003,N_9946);
or U10871 (N_10871,N_9980,N_10322);
or U10872 (N_10872,N_9855,N_10196);
nor U10873 (N_10873,N_10118,N_9883);
and U10874 (N_10874,N_10157,N_10486);
xor U10875 (N_10875,N_9978,N_10415);
nand U10876 (N_10876,N_9751,N_10038);
nand U10877 (N_10877,N_9950,N_10459);
nand U10878 (N_10878,N_10474,N_10473);
xor U10879 (N_10879,N_10026,N_10105);
or U10880 (N_10880,N_10287,N_10134);
or U10881 (N_10881,N_9901,N_10215);
and U10882 (N_10882,N_10494,N_10304);
nand U10883 (N_10883,N_9850,N_10060);
nand U10884 (N_10884,N_10180,N_10297);
nand U10885 (N_10885,N_10355,N_9893);
or U10886 (N_10886,N_10302,N_9831);
or U10887 (N_10887,N_10230,N_10177);
nand U10888 (N_10888,N_10410,N_10327);
nor U10889 (N_10889,N_10137,N_10070);
or U10890 (N_10890,N_10073,N_10493);
xor U10891 (N_10891,N_10113,N_10401);
nand U10892 (N_10892,N_10122,N_9756);
nor U10893 (N_10893,N_9760,N_10284);
xnor U10894 (N_10894,N_9964,N_10136);
nor U10895 (N_10895,N_10011,N_9818);
and U10896 (N_10896,N_10186,N_10402);
xnor U10897 (N_10897,N_10080,N_10458);
or U10898 (N_10898,N_10403,N_10204);
nand U10899 (N_10899,N_10447,N_9826);
xor U10900 (N_10900,N_9772,N_10111);
or U10901 (N_10901,N_9761,N_10095);
or U10902 (N_10902,N_9768,N_9973);
xor U10903 (N_10903,N_9990,N_10456);
or U10904 (N_10904,N_9935,N_10147);
nand U10905 (N_10905,N_10054,N_9844);
and U10906 (N_10906,N_9847,N_10104);
and U10907 (N_10907,N_10050,N_9812);
nor U10908 (N_10908,N_10050,N_9981);
nor U10909 (N_10909,N_10077,N_10009);
or U10910 (N_10910,N_10456,N_10421);
xor U10911 (N_10911,N_10159,N_9797);
and U10912 (N_10912,N_10311,N_9972);
xor U10913 (N_10913,N_10210,N_10434);
and U10914 (N_10914,N_10115,N_10148);
nor U10915 (N_10915,N_10378,N_9987);
xor U10916 (N_10916,N_10374,N_10383);
nor U10917 (N_10917,N_10083,N_9973);
nand U10918 (N_10918,N_10011,N_10034);
and U10919 (N_10919,N_10170,N_10423);
nand U10920 (N_10920,N_9758,N_10236);
or U10921 (N_10921,N_9883,N_10255);
nand U10922 (N_10922,N_10117,N_10149);
or U10923 (N_10923,N_10231,N_9803);
and U10924 (N_10924,N_9951,N_10456);
or U10925 (N_10925,N_9909,N_10058);
nand U10926 (N_10926,N_10261,N_10342);
and U10927 (N_10927,N_10407,N_10037);
nand U10928 (N_10928,N_10336,N_10414);
nor U10929 (N_10929,N_10408,N_10258);
nor U10930 (N_10930,N_10068,N_9970);
nand U10931 (N_10931,N_9993,N_9799);
nor U10932 (N_10932,N_10349,N_10018);
xnor U10933 (N_10933,N_9818,N_9858);
and U10934 (N_10934,N_9937,N_10124);
or U10935 (N_10935,N_10304,N_10064);
nor U10936 (N_10936,N_9797,N_10312);
nor U10937 (N_10937,N_10187,N_9866);
or U10938 (N_10938,N_10294,N_9758);
nor U10939 (N_10939,N_9820,N_9852);
nor U10940 (N_10940,N_10243,N_10055);
nor U10941 (N_10941,N_9797,N_10273);
nor U10942 (N_10942,N_9993,N_9959);
nor U10943 (N_10943,N_9818,N_10494);
xor U10944 (N_10944,N_10053,N_10136);
nand U10945 (N_10945,N_10235,N_10092);
and U10946 (N_10946,N_9911,N_9811);
or U10947 (N_10947,N_10416,N_9890);
xnor U10948 (N_10948,N_10347,N_10443);
or U10949 (N_10949,N_10453,N_10205);
nand U10950 (N_10950,N_10076,N_10399);
nand U10951 (N_10951,N_10317,N_9907);
xnor U10952 (N_10952,N_9890,N_10170);
and U10953 (N_10953,N_9855,N_10385);
nor U10954 (N_10954,N_9922,N_10168);
and U10955 (N_10955,N_10478,N_10256);
xnor U10956 (N_10956,N_9865,N_10449);
and U10957 (N_10957,N_10436,N_10343);
nand U10958 (N_10958,N_10461,N_10350);
or U10959 (N_10959,N_10237,N_10137);
and U10960 (N_10960,N_9932,N_10074);
xnor U10961 (N_10961,N_10309,N_10316);
and U10962 (N_10962,N_9770,N_10121);
nand U10963 (N_10963,N_10390,N_10337);
nor U10964 (N_10964,N_10025,N_10404);
nand U10965 (N_10965,N_10436,N_10479);
and U10966 (N_10966,N_9925,N_9818);
and U10967 (N_10967,N_9932,N_10169);
nor U10968 (N_10968,N_9868,N_10054);
nor U10969 (N_10969,N_9926,N_10456);
or U10970 (N_10970,N_10177,N_10219);
xnor U10971 (N_10971,N_9950,N_10380);
xnor U10972 (N_10972,N_10236,N_10428);
and U10973 (N_10973,N_10413,N_10336);
and U10974 (N_10974,N_10175,N_10450);
nor U10975 (N_10975,N_10072,N_9976);
xor U10976 (N_10976,N_10470,N_9856);
xnor U10977 (N_10977,N_9790,N_10215);
xnor U10978 (N_10978,N_10146,N_10116);
nor U10979 (N_10979,N_9795,N_10312);
or U10980 (N_10980,N_10140,N_10410);
and U10981 (N_10981,N_10291,N_9987);
and U10982 (N_10982,N_10059,N_10271);
nor U10983 (N_10983,N_10228,N_9874);
or U10984 (N_10984,N_10204,N_10197);
and U10985 (N_10985,N_10092,N_10072);
or U10986 (N_10986,N_10498,N_10317);
and U10987 (N_10987,N_9888,N_9801);
nor U10988 (N_10988,N_10395,N_10053);
nor U10989 (N_10989,N_9946,N_10300);
xnor U10990 (N_10990,N_10072,N_9760);
xor U10991 (N_10991,N_10297,N_10115);
nand U10992 (N_10992,N_9892,N_10005);
or U10993 (N_10993,N_10098,N_10324);
and U10994 (N_10994,N_10331,N_9786);
nand U10995 (N_10995,N_10219,N_10074);
and U10996 (N_10996,N_10406,N_9852);
xor U10997 (N_10997,N_10180,N_10442);
or U10998 (N_10998,N_10328,N_10457);
and U10999 (N_10999,N_10311,N_10279);
and U11000 (N_11000,N_10428,N_10058);
and U11001 (N_11001,N_10397,N_10199);
and U11002 (N_11002,N_9880,N_10489);
nor U11003 (N_11003,N_9826,N_10019);
xor U11004 (N_11004,N_10439,N_10271);
nor U11005 (N_11005,N_10003,N_10229);
and U11006 (N_11006,N_10075,N_10112);
nor U11007 (N_11007,N_10131,N_10298);
nand U11008 (N_11008,N_10353,N_9828);
or U11009 (N_11009,N_9846,N_9929);
nand U11010 (N_11010,N_10384,N_10052);
and U11011 (N_11011,N_9761,N_9971);
or U11012 (N_11012,N_9992,N_10306);
nor U11013 (N_11013,N_10227,N_10198);
nand U11014 (N_11014,N_10387,N_10087);
nand U11015 (N_11015,N_9760,N_10028);
nor U11016 (N_11016,N_10435,N_10049);
xnor U11017 (N_11017,N_9956,N_10068);
nand U11018 (N_11018,N_10005,N_9917);
nand U11019 (N_11019,N_9963,N_10445);
xor U11020 (N_11020,N_10290,N_9820);
and U11021 (N_11021,N_10425,N_10414);
or U11022 (N_11022,N_9953,N_10354);
and U11023 (N_11023,N_9892,N_9984);
and U11024 (N_11024,N_9758,N_10139);
or U11025 (N_11025,N_9856,N_10207);
and U11026 (N_11026,N_10015,N_9913);
xnor U11027 (N_11027,N_10125,N_10196);
or U11028 (N_11028,N_9895,N_9957);
nand U11029 (N_11029,N_10309,N_10439);
nor U11030 (N_11030,N_9865,N_9759);
nor U11031 (N_11031,N_10116,N_9914);
xnor U11032 (N_11032,N_10347,N_10006);
nor U11033 (N_11033,N_9891,N_9982);
xnor U11034 (N_11034,N_9873,N_10320);
or U11035 (N_11035,N_10373,N_10456);
nand U11036 (N_11036,N_9945,N_9939);
xnor U11037 (N_11037,N_9753,N_9995);
nand U11038 (N_11038,N_9802,N_9988);
and U11039 (N_11039,N_10139,N_10315);
and U11040 (N_11040,N_10026,N_9941);
nor U11041 (N_11041,N_10112,N_10495);
nor U11042 (N_11042,N_9808,N_10051);
xnor U11043 (N_11043,N_9790,N_10236);
xnor U11044 (N_11044,N_10214,N_10113);
nand U11045 (N_11045,N_10133,N_9766);
or U11046 (N_11046,N_10182,N_10075);
xnor U11047 (N_11047,N_10473,N_10372);
or U11048 (N_11048,N_10014,N_9925);
nand U11049 (N_11049,N_10021,N_10040);
nor U11050 (N_11050,N_10051,N_9892);
or U11051 (N_11051,N_10460,N_10187);
nand U11052 (N_11052,N_9814,N_10085);
and U11053 (N_11053,N_9834,N_10206);
or U11054 (N_11054,N_10422,N_10125);
or U11055 (N_11055,N_9807,N_10254);
nand U11056 (N_11056,N_10251,N_10102);
xnor U11057 (N_11057,N_9964,N_10197);
nor U11058 (N_11058,N_10472,N_10275);
nor U11059 (N_11059,N_9916,N_10227);
and U11060 (N_11060,N_10274,N_10285);
xnor U11061 (N_11061,N_9946,N_10444);
or U11062 (N_11062,N_10124,N_10389);
and U11063 (N_11063,N_10212,N_9900);
xor U11064 (N_11064,N_10101,N_10075);
nor U11065 (N_11065,N_10443,N_10482);
nand U11066 (N_11066,N_10029,N_9934);
xnor U11067 (N_11067,N_9858,N_10059);
nand U11068 (N_11068,N_9978,N_9914);
and U11069 (N_11069,N_10381,N_9812);
nor U11070 (N_11070,N_10403,N_10089);
or U11071 (N_11071,N_10246,N_9802);
and U11072 (N_11072,N_10098,N_9843);
and U11073 (N_11073,N_9853,N_10144);
and U11074 (N_11074,N_10128,N_10313);
nand U11075 (N_11075,N_10303,N_10199);
and U11076 (N_11076,N_10463,N_10413);
or U11077 (N_11077,N_9877,N_9764);
and U11078 (N_11078,N_9855,N_10090);
and U11079 (N_11079,N_10212,N_10007);
and U11080 (N_11080,N_10168,N_10217);
xor U11081 (N_11081,N_10176,N_10438);
and U11082 (N_11082,N_10113,N_10211);
xnor U11083 (N_11083,N_10432,N_9913);
or U11084 (N_11084,N_10272,N_10080);
and U11085 (N_11085,N_10057,N_10033);
and U11086 (N_11086,N_9918,N_10430);
or U11087 (N_11087,N_10192,N_10333);
nor U11088 (N_11088,N_9908,N_10278);
or U11089 (N_11089,N_10200,N_10049);
nor U11090 (N_11090,N_10022,N_10032);
nand U11091 (N_11091,N_10433,N_9788);
nand U11092 (N_11092,N_10132,N_9815);
nor U11093 (N_11093,N_9830,N_9894);
and U11094 (N_11094,N_10295,N_10304);
nor U11095 (N_11095,N_10416,N_10235);
and U11096 (N_11096,N_10472,N_10199);
xor U11097 (N_11097,N_10101,N_10438);
and U11098 (N_11098,N_10061,N_10011);
or U11099 (N_11099,N_9885,N_10198);
nor U11100 (N_11100,N_10230,N_10449);
xnor U11101 (N_11101,N_10420,N_10363);
xor U11102 (N_11102,N_10063,N_10284);
or U11103 (N_11103,N_10476,N_9976);
and U11104 (N_11104,N_10369,N_9822);
and U11105 (N_11105,N_10190,N_9974);
and U11106 (N_11106,N_10048,N_9966);
and U11107 (N_11107,N_10439,N_9823);
and U11108 (N_11108,N_10138,N_10467);
or U11109 (N_11109,N_10475,N_9910);
xor U11110 (N_11110,N_10457,N_10188);
and U11111 (N_11111,N_10168,N_10009);
or U11112 (N_11112,N_9831,N_10301);
xor U11113 (N_11113,N_10216,N_10010);
or U11114 (N_11114,N_10296,N_10405);
xnor U11115 (N_11115,N_10309,N_9920);
and U11116 (N_11116,N_9813,N_10484);
or U11117 (N_11117,N_9980,N_10246);
nand U11118 (N_11118,N_10092,N_9933);
nor U11119 (N_11119,N_10319,N_9850);
xor U11120 (N_11120,N_10366,N_10331);
and U11121 (N_11121,N_9790,N_10047);
nand U11122 (N_11122,N_9941,N_9878);
xor U11123 (N_11123,N_10001,N_9928);
and U11124 (N_11124,N_10241,N_9779);
xor U11125 (N_11125,N_10022,N_10128);
and U11126 (N_11126,N_9841,N_10205);
xnor U11127 (N_11127,N_9914,N_9925);
nor U11128 (N_11128,N_10351,N_10056);
or U11129 (N_11129,N_10143,N_10408);
xnor U11130 (N_11130,N_10201,N_9958);
or U11131 (N_11131,N_10106,N_10423);
xnor U11132 (N_11132,N_10136,N_10248);
and U11133 (N_11133,N_10464,N_10275);
nand U11134 (N_11134,N_10342,N_10054);
nor U11135 (N_11135,N_10158,N_10090);
nor U11136 (N_11136,N_9855,N_10295);
or U11137 (N_11137,N_10250,N_10475);
or U11138 (N_11138,N_10328,N_9754);
xnor U11139 (N_11139,N_10403,N_10295);
nand U11140 (N_11140,N_10012,N_9838);
nor U11141 (N_11141,N_10385,N_10325);
nand U11142 (N_11142,N_10288,N_9816);
and U11143 (N_11143,N_10292,N_10458);
and U11144 (N_11144,N_10014,N_9915);
or U11145 (N_11145,N_10398,N_10184);
or U11146 (N_11146,N_10480,N_10220);
nor U11147 (N_11147,N_10111,N_9816);
xnor U11148 (N_11148,N_9969,N_9891);
or U11149 (N_11149,N_9871,N_10135);
and U11150 (N_11150,N_10384,N_9813);
and U11151 (N_11151,N_10005,N_9901);
xnor U11152 (N_11152,N_10447,N_10421);
and U11153 (N_11153,N_10201,N_9885);
nand U11154 (N_11154,N_10347,N_10388);
xor U11155 (N_11155,N_10364,N_9863);
nor U11156 (N_11156,N_10265,N_10399);
xor U11157 (N_11157,N_10430,N_10461);
nor U11158 (N_11158,N_9807,N_10203);
nand U11159 (N_11159,N_10101,N_10343);
or U11160 (N_11160,N_9955,N_9848);
and U11161 (N_11161,N_10474,N_10220);
nor U11162 (N_11162,N_10459,N_9888);
nand U11163 (N_11163,N_9910,N_10086);
nor U11164 (N_11164,N_10046,N_9986);
xor U11165 (N_11165,N_10277,N_9848);
nor U11166 (N_11166,N_10477,N_9988);
nand U11167 (N_11167,N_10058,N_10378);
and U11168 (N_11168,N_10063,N_10434);
and U11169 (N_11169,N_10119,N_10468);
nand U11170 (N_11170,N_9801,N_10155);
or U11171 (N_11171,N_9958,N_10371);
or U11172 (N_11172,N_10323,N_10479);
xor U11173 (N_11173,N_10432,N_10171);
nand U11174 (N_11174,N_9890,N_10090);
xnor U11175 (N_11175,N_10461,N_10275);
nand U11176 (N_11176,N_10478,N_10373);
or U11177 (N_11177,N_10052,N_10193);
nor U11178 (N_11178,N_10141,N_9944);
or U11179 (N_11179,N_10283,N_9801);
xor U11180 (N_11180,N_9846,N_9938);
nand U11181 (N_11181,N_9841,N_9835);
or U11182 (N_11182,N_10184,N_10081);
and U11183 (N_11183,N_9792,N_10421);
xor U11184 (N_11184,N_9807,N_10085);
nand U11185 (N_11185,N_10235,N_10381);
and U11186 (N_11186,N_9944,N_10115);
and U11187 (N_11187,N_9962,N_10204);
nand U11188 (N_11188,N_9868,N_10277);
or U11189 (N_11189,N_10151,N_10450);
nand U11190 (N_11190,N_10169,N_9799);
nand U11191 (N_11191,N_10166,N_10149);
and U11192 (N_11192,N_9920,N_9865);
nand U11193 (N_11193,N_10369,N_10488);
nand U11194 (N_11194,N_10136,N_10174);
and U11195 (N_11195,N_10022,N_9858);
nand U11196 (N_11196,N_9880,N_10162);
nand U11197 (N_11197,N_10265,N_9955);
and U11198 (N_11198,N_9981,N_9777);
nand U11199 (N_11199,N_10047,N_10204);
and U11200 (N_11200,N_10037,N_10176);
and U11201 (N_11201,N_9778,N_9791);
xor U11202 (N_11202,N_9932,N_10252);
nor U11203 (N_11203,N_9901,N_9951);
xnor U11204 (N_11204,N_10456,N_10084);
xnor U11205 (N_11205,N_9981,N_10279);
or U11206 (N_11206,N_10155,N_9785);
nor U11207 (N_11207,N_9900,N_10434);
xor U11208 (N_11208,N_9890,N_10375);
or U11209 (N_11209,N_10236,N_10108);
or U11210 (N_11210,N_10395,N_10453);
nor U11211 (N_11211,N_10188,N_9943);
nand U11212 (N_11212,N_10365,N_10192);
xnor U11213 (N_11213,N_10022,N_10126);
xor U11214 (N_11214,N_10449,N_10359);
or U11215 (N_11215,N_9906,N_10224);
xor U11216 (N_11216,N_9864,N_10442);
xnor U11217 (N_11217,N_10372,N_9796);
and U11218 (N_11218,N_9861,N_10073);
nand U11219 (N_11219,N_9787,N_10114);
nor U11220 (N_11220,N_10356,N_10264);
or U11221 (N_11221,N_9997,N_10092);
or U11222 (N_11222,N_9994,N_10189);
nor U11223 (N_11223,N_10037,N_10131);
or U11224 (N_11224,N_10444,N_10041);
nand U11225 (N_11225,N_10059,N_9911);
or U11226 (N_11226,N_10388,N_9886);
xor U11227 (N_11227,N_10183,N_10061);
nand U11228 (N_11228,N_10462,N_10293);
xor U11229 (N_11229,N_10452,N_10366);
nand U11230 (N_11230,N_10331,N_10407);
or U11231 (N_11231,N_9805,N_10120);
or U11232 (N_11232,N_9985,N_10098);
xnor U11233 (N_11233,N_10429,N_9841);
xor U11234 (N_11234,N_10196,N_10390);
xor U11235 (N_11235,N_10328,N_10114);
nand U11236 (N_11236,N_9786,N_10368);
nand U11237 (N_11237,N_9784,N_10127);
and U11238 (N_11238,N_9996,N_10147);
and U11239 (N_11239,N_9997,N_10176);
xor U11240 (N_11240,N_10493,N_9809);
nand U11241 (N_11241,N_9888,N_10370);
and U11242 (N_11242,N_10367,N_9931);
xor U11243 (N_11243,N_10307,N_9986);
or U11244 (N_11244,N_10062,N_9758);
and U11245 (N_11245,N_10289,N_10463);
nand U11246 (N_11246,N_10160,N_9801);
or U11247 (N_11247,N_10358,N_10113);
nor U11248 (N_11248,N_10318,N_10210);
nand U11249 (N_11249,N_10009,N_9784);
nand U11250 (N_11250,N_10606,N_10927);
and U11251 (N_11251,N_10601,N_11229);
and U11252 (N_11252,N_10573,N_11081);
and U11253 (N_11253,N_10856,N_11154);
xnor U11254 (N_11254,N_10539,N_10855);
and U11255 (N_11255,N_10508,N_11069);
or U11256 (N_11256,N_10797,N_10540);
xnor U11257 (N_11257,N_10872,N_10788);
and U11258 (N_11258,N_10700,N_10627);
and U11259 (N_11259,N_11086,N_10656);
or U11260 (N_11260,N_10568,N_10911);
or U11261 (N_11261,N_10934,N_11076);
xor U11262 (N_11262,N_10860,N_10950);
xnor U11263 (N_11263,N_10883,N_10807);
or U11264 (N_11264,N_10654,N_10829);
nand U11265 (N_11265,N_10737,N_11037);
and U11266 (N_11266,N_10967,N_11056);
xor U11267 (N_11267,N_11060,N_11162);
and U11268 (N_11268,N_10873,N_10770);
and U11269 (N_11269,N_10526,N_10838);
or U11270 (N_11270,N_10703,N_10581);
xnor U11271 (N_11271,N_10789,N_10559);
and U11272 (N_11272,N_11207,N_11084);
nor U11273 (N_11273,N_11139,N_10577);
or U11274 (N_11274,N_11074,N_11015);
nor U11275 (N_11275,N_10887,N_10918);
nand U11276 (N_11276,N_10906,N_10977);
nand U11277 (N_11277,N_10739,N_10738);
and U11278 (N_11278,N_11133,N_11117);
nor U11279 (N_11279,N_10831,N_10812);
and U11280 (N_11280,N_11203,N_10956);
and U11281 (N_11281,N_11214,N_10969);
xnor U11282 (N_11282,N_10554,N_10548);
nand U11283 (N_11283,N_11205,N_11151);
nor U11284 (N_11284,N_10530,N_11095);
xor U11285 (N_11285,N_10923,N_10774);
nor U11286 (N_11286,N_10931,N_10575);
xnor U11287 (N_11287,N_11009,N_10562);
and U11288 (N_11288,N_10919,N_10979);
or U11289 (N_11289,N_10556,N_10749);
and U11290 (N_11290,N_10631,N_11067);
xor U11291 (N_11291,N_10981,N_11241);
and U11292 (N_11292,N_11247,N_11124);
and U11293 (N_11293,N_10995,N_10764);
nor U11294 (N_11294,N_11248,N_11055);
nand U11295 (N_11295,N_10946,N_11177);
or U11296 (N_11296,N_11103,N_11057);
nand U11297 (N_11297,N_10811,N_10713);
and U11298 (N_11298,N_10828,N_10620);
nor U11299 (N_11299,N_10756,N_10904);
or U11300 (N_11300,N_10718,N_10534);
and U11301 (N_11301,N_10531,N_10678);
or U11302 (N_11302,N_10507,N_10661);
xor U11303 (N_11303,N_10558,N_11190);
nand U11304 (N_11304,N_10775,N_10611);
and U11305 (N_11305,N_11080,N_10852);
or U11306 (N_11306,N_11028,N_10791);
xnor U11307 (N_11307,N_11004,N_10599);
xor U11308 (N_11308,N_10910,N_10850);
and U11309 (N_11309,N_10622,N_10624);
and U11310 (N_11310,N_10653,N_10916);
nand U11311 (N_11311,N_10961,N_10688);
or U11312 (N_11312,N_11220,N_10633);
or U11313 (N_11313,N_10869,N_10827);
nand U11314 (N_11314,N_11148,N_10999);
nor U11315 (N_11315,N_11007,N_11032);
and U11316 (N_11316,N_10900,N_10746);
or U11317 (N_11317,N_10937,N_10751);
nor U11318 (N_11318,N_11236,N_10804);
or U11319 (N_11319,N_11132,N_10663);
or U11320 (N_11320,N_10741,N_11094);
or U11321 (N_11321,N_10571,N_10816);
or U11322 (N_11322,N_11116,N_11039);
or U11323 (N_11323,N_10691,N_11199);
xnor U11324 (N_11324,N_10566,N_11170);
xor U11325 (N_11325,N_10597,N_10978);
nor U11326 (N_11326,N_10708,N_11111);
or U11327 (N_11327,N_10521,N_11156);
and U11328 (N_11328,N_11246,N_10676);
nand U11329 (N_11329,N_10520,N_10854);
xnor U11330 (N_11330,N_10564,N_10522);
xnor U11331 (N_11331,N_11054,N_10941);
xor U11332 (N_11332,N_10596,N_11138);
and U11333 (N_11333,N_11237,N_10712);
or U11334 (N_11334,N_11130,N_10859);
and U11335 (N_11335,N_10636,N_10734);
and U11336 (N_11336,N_11105,N_11106);
or U11337 (N_11337,N_10962,N_11194);
xnor U11338 (N_11338,N_11167,N_10629);
nand U11339 (N_11339,N_10996,N_11089);
or U11340 (N_11340,N_11006,N_10728);
nand U11341 (N_11341,N_10953,N_10662);
nor U11342 (N_11342,N_10879,N_10849);
xnor U11343 (N_11343,N_10871,N_10510);
nand U11344 (N_11344,N_10890,N_10716);
or U11345 (N_11345,N_10782,N_10808);
nand U11346 (N_11346,N_11046,N_11181);
nor U11347 (N_11347,N_10786,N_10701);
nor U11348 (N_11348,N_10524,N_10707);
xor U11349 (N_11349,N_11096,N_10833);
nand U11350 (N_11350,N_10635,N_10802);
nor U11351 (N_11351,N_11114,N_10655);
and U11352 (N_11352,N_11137,N_11090);
nand U11353 (N_11353,N_11019,N_10543);
nor U11354 (N_11354,N_10965,N_11200);
nor U11355 (N_11355,N_11230,N_10868);
and U11356 (N_11356,N_10652,N_10503);
or U11357 (N_11357,N_11212,N_10894);
nor U11358 (N_11358,N_10844,N_10837);
nor U11359 (N_11359,N_11008,N_10588);
and U11360 (N_11360,N_11184,N_10985);
xnor U11361 (N_11361,N_10690,N_10867);
or U11362 (N_11362,N_11213,N_10892);
and U11363 (N_11363,N_10515,N_11048);
or U11364 (N_11364,N_10974,N_10924);
and U11365 (N_11365,N_10762,N_10509);
nand U11366 (N_11366,N_10765,N_11136);
nor U11367 (N_11367,N_11208,N_10574);
nor U11368 (N_11368,N_10874,N_10563);
nor U11369 (N_11369,N_10760,N_10914);
nor U11370 (N_11370,N_10529,N_11211);
and U11371 (N_11371,N_10839,N_11066);
or U11372 (N_11372,N_11176,N_11118);
or U11373 (N_11373,N_10683,N_10517);
xnor U11374 (N_11374,N_10641,N_11159);
or U11375 (N_11375,N_10730,N_11001);
and U11376 (N_11376,N_10527,N_10818);
nor U11377 (N_11377,N_10644,N_10593);
or U11378 (N_11378,N_10901,N_10785);
or U11379 (N_11379,N_11215,N_10648);
xnor U11380 (N_11380,N_10549,N_10699);
nor U11381 (N_11381,N_11228,N_11180);
xnor U11382 (N_11382,N_10561,N_10975);
xor U11383 (N_11383,N_11204,N_10618);
xor U11384 (N_11384,N_11249,N_10799);
xnor U11385 (N_11385,N_10528,N_11003);
and U11386 (N_11386,N_10694,N_11027);
nand U11387 (N_11387,N_10815,N_10755);
nor U11388 (N_11388,N_10821,N_11239);
nor U11389 (N_11389,N_11129,N_11115);
xor U11390 (N_11390,N_10665,N_10589);
nor U11391 (N_11391,N_10915,N_10912);
nand U11392 (N_11392,N_10862,N_10537);
nor U11393 (N_11393,N_10602,N_10920);
or U11394 (N_11394,N_10922,N_11031);
and U11395 (N_11395,N_11041,N_10731);
xnor U11396 (N_11396,N_11034,N_10882);
nand U11397 (N_11397,N_11050,N_10555);
xor U11398 (N_11398,N_11023,N_10938);
nor U11399 (N_11399,N_10903,N_10584);
or U11400 (N_11400,N_10613,N_11217);
or U11401 (N_11401,N_10754,N_10902);
and U11402 (N_11402,N_10546,N_10952);
or U11403 (N_11403,N_10758,N_10949);
xor U11404 (N_11404,N_11222,N_10630);
nand U11405 (N_11405,N_10940,N_10779);
or U11406 (N_11406,N_11053,N_11134);
or U11407 (N_11407,N_11145,N_10814);
nand U11408 (N_11408,N_10777,N_10541);
and U11409 (N_11409,N_10675,N_11083);
xor U11410 (N_11410,N_10625,N_10992);
and U11411 (N_11411,N_10935,N_10616);
nand U11412 (N_11412,N_11020,N_10501);
or U11413 (N_11413,N_10553,N_10725);
nor U11414 (N_11414,N_10748,N_11146);
and U11415 (N_11415,N_10659,N_10928);
or U11416 (N_11416,N_10830,N_10710);
and U11417 (N_11417,N_11099,N_10735);
nand U11418 (N_11418,N_10970,N_10727);
and U11419 (N_11419,N_11010,N_10768);
xor U11420 (N_11420,N_11243,N_11234);
and U11421 (N_11421,N_10677,N_10997);
and U11422 (N_11422,N_11063,N_10858);
nor U11423 (N_11423,N_10796,N_10889);
or U11424 (N_11424,N_10976,N_10715);
xor U11425 (N_11425,N_10664,N_10547);
or U11426 (N_11426,N_10948,N_10790);
xor U11427 (N_11427,N_10698,N_10769);
and U11428 (N_11428,N_11172,N_10957);
nor U11429 (N_11429,N_11123,N_10702);
or U11430 (N_11430,N_10750,N_11013);
or U11431 (N_11431,N_10669,N_10542);
nand U11432 (N_11432,N_10570,N_10557);
nand U11433 (N_11433,N_10773,N_10612);
xnor U11434 (N_11434,N_10847,N_10504);
nor U11435 (N_11435,N_11153,N_10865);
or U11436 (N_11436,N_11070,N_11166);
nand U11437 (N_11437,N_10822,N_10679);
or U11438 (N_11438,N_10886,N_11065);
or U11439 (N_11439,N_11068,N_10670);
nor U11440 (N_11440,N_10836,N_11195);
nor U11441 (N_11441,N_10733,N_10704);
xor U11442 (N_11442,N_11051,N_10896);
xor U11443 (N_11443,N_11021,N_11036);
and U11444 (N_11444,N_11078,N_11127);
and U11445 (N_11445,N_11128,N_11169);
xor U11446 (N_11446,N_10650,N_10569);
and U11447 (N_11447,N_10532,N_11044);
xor U11448 (N_11448,N_10619,N_10726);
xor U11449 (N_11449,N_11072,N_11017);
xnor U11450 (N_11450,N_10697,N_10825);
nand U11451 (N_11451,N_10861,N_11045);
nand U11452 (N_11452,N_10909,N_10870);
or U11453 (N_11453,N_11058,N_11100);
and U11454 (N_11454,N_10891,N_10888);
xnor U11455 (N_11455,N_10719,N_11142);
nor U11456 (N_11456,N_11174,N_10848);
xor U11457 (N_11457,N_11087,N_11108);
xor U11458 (N_11458,N_11097,N_10955);
xnor U11459 (N_11459,N_11160,N_11149);
nor U11460 (N_11460,N_11120,N_10692);
nand U11461 (N_11461,N_10968,N_11206);
or U11462 (N_11462,N_10877,N_11125);
or U11463 (N_11463,N_10711,N_10668);
and U11464 (N_11464,N_11235,N_10876);
nand U11465 (N_11465,N_10806,N_10823);
and U11466 (N_11466,N_11155,N_11189);
nand U11467 (N_11467,N_10706,N_10745);
xor U11468 (N_11468,N_10893,N_10714);
nand U11469 (N_11469,N_10724,N_10632);
and U11470 (N_11470,N_11188,N_10983);
and U11471 (N_11471,N_10817,N_10586);
nor U11472 (N_11472,N_10533,N_10842);
nand U11473 (N_11473,N_10987,N_10638);
and U11474 (N_11474,N_10567,N_11157);
nand U11475 (N_11475,N_11164,N_10843);
or U11476 (N_11476,N_11135,N_10752);
nand U11477 (N_11477,N_10605,N_10973);
nand U11478 (N_11478,N_11071,N_11088);
and U11479 (N_11479,N_10792,N_10742);
nor U11480 (N_11480,N_10803,N_10729);
nor U11481 (N_11481,N_11043,N_10610);
nor U11482 (N_11482,N_11187,N_11052);
or U11483 (N_11483,N_10959,N_11179);
and U11484 (N_11484,N_11245,N_10998);
and U11485 (N_11485,N_11047,N_11126);
and U11486 (N_11486,N_10732,N_10971);
xnor U11487 (N_11487,N_10645,N_10932);
nand U11488 (N_11488,N_10958,N_11225);
nand U11489 (N_11489,N_11196,N_10988);
xor U11490 (N_11490,N_10525,N_11022);
xnor U11491 (N_11491,N_10693,N_10881);
or U11492 (N_11492,N_10851,N_10642);
xor U11493 (N_11493,N_10991,N_10572);
or U11494 (N_11494,N_10884,N_11091);
nand U11495 (N_11495,N_11104,N_11192);
nor U11496 (N_11496,N_10578,N_10684);
nand U11497 (N_11497,N_11026,N_11061);
and U11498 (N_11498,N_10989,N_11202);
and U11499 (N_11499,N_10846,N_11059);
or U11500 (N_11500,N_10820,N_11005);
nand U11501 (N_11501,N_10740,N_11049);
xnor U11502 (N_11502,N_11197,N_10945);
or U11503 (N_11503,N_10639,N_11121);
or U11504 (N_11504,N_10926,N_10695);
nor U11505 (N_11505,N_11101,N_11144);
nand U11506 (N_11506,N_10763,N_11062);
nand U11507 (N_11507,N_11210,N_11064);
or U11508 (N_11508,N_11098,N_10966);
and U11509 (N_11509,N_10516,N_10506);
or U11510 (N_11510,N_11079,N_10743);
or U11511 (N_11511,N_10607,N_11165);
nor U11512 (N_11512,N_10671,N_10772);
nor U11513 (N_11513,N_10594,N_11012);
nor U11514 (N_11514,N_10628,N_11143);
nor U11515 (N_11515,N_11030,N_11221);
or U11516 (N_11516,N_10864,N_11226);
and U11517 (N_11517,N_10929,N_10943);
nor U11518 (N_11518,N_10744,N_10885);
xor U11519 (N_11519,N_10917,N_11198);
nand U11520 (N_11520,N_10519,N_11182);
xor U11521 (N_11521,N_10944,N_10964);
nor U11522 (N_11522,N_11238,N_11209);
or U11523 (N_11523,N_11161,N_11040);
xnor U11524 (N_11524,N_11244,N_10897);
xnor U11525 (N_11525,N_10819,N_10853);
or U11526 (N_11526,N_10793,N_11107);
nor U11527 (N_11527,N_10895,N_11018);
nor U11528 (N_11528,N_10835,N_11109);
xnor U11529 (N_11529,N_11183,N_10657);
and U11530 (N_11530,N_10595,N_10687);
xnor U11531 (N_11531,N_10778,N_10810);
nand U11532 (N_11532,N_11158,N_10585);
nand U11533 (N_11533,N_10805,N_10936);
or U11534 (N_11534,N_11224,N_10960);
nand U11535 (N_11535,N_10809,N_10993);
nor U11536 (N_11536,N_10552,N_10544);
xnor U11537 (N_11537,N_10682,N_10640);
nor U11538 (N_11538,N_10753,N_10757);
xor U11539 (N_11539,N_10623,N_11141);
or U11540 (N_11540,N_11219,N_10560);
or U11541 (N_11541,N_10951,N_10673);
nand U11542 (N_11542,N_11216,N_10598);
nand U11543 (N_11543,N_10634,N_10505);
or U11544 (N_11544,N_10550,N_10651);
and U11545 (N_11545,N_11185,N_10681);
nor U11546 (N_11546,N_10982,N_10514);
nor U11547 (N_11547,N_10565,N_11227);
nor U11548 (N_11548,N_11150,N_10972);
and U11549 (N_11549,N_10643,N_11113);
xor U11550 (N_11550,N_11178,N_11038);
or U11551 (N_11551,N_10841,N_11186);
nor U11552 (N_11552,N_11232,N_10899);
xnor U11553 (N_11553,N_10866,N_10795);
or U11554 (N_11554,N_10579,N_10580);
nand U11555 (N_11555,N_10722,N_10600);
or U11556 (N_11556,N_10880,N_11093);
nor U11557 (N_11557,N_10603,N_11016);
xor U11558 (N_11558,N_11171,N_11131);
nor U11559 (N_11559,N_10840,N_11168);
xnor U11560 (N_11560,N_10720,N_11014);
xor U11561 (N_11561,N_11025,N_10986);
xnor U11562 (N_11562,N_10686,N_10626);
xnor U11563 (N_11563,N_10780,N_10689);
nand U11564 (N_11564,N_10857,N_10921);
nor U11565 (N_11565,N_10666,N_10512);
or U11566 (N_11566,N_10621,N_10646);
or U11567 (N_11567,N_10535,N_10609);
xor U11568 (N_11568,N_11011,N_10615);
or U11569 (N_11569,N_10604,N_11233);
xnor U11570 (N_11570,N_10908,N_11147);
or U11571 (N_11571,N_10660,N_11073);
nand U11572 (N_11572,N_10658,N_10637);
nand U11573 (N_11573,N_10747,N_10980);
xnor U11574 (N_11574,N_11119,N_10536);
or U11575 (N_11575,N_10942,N_11035);
nand U11576 (N_11576,N_10523,N_10800);
nor U11577 (N_11577,N_11092,N_10905);
nand U11578 (N_11578,N_10963,N_11163);
xnor U11579 (N_11579,N_10990,N_10717);
nand U11580 (N_11580,N_10551,N_11201);
and U11581 (N_11581,N_10590,N_10994);
or U11582 (N_11582,N_10794,N_10545);
and U11583 (N_11583,N_10592,N_10614);
and U11584 (N_11584,N_10875,N_10913);
nor U11585 (N_11585,N_10608,N_10824);
nand U11586 (N_11586,N_10781,N_11110);
xnor U11587 (N_11587,N_10518,N_10898);
or U11588 (N_11588,N_11102,N_10845);
nand U11589 (N_11589,N_11231,N_10771);
nor U11590 (N_11590,N_10705,N_10947);
nor U11591 (N_11591,N_11112,N_10767);
nor U11592 (N_11592,N_10674,N_10878);
nor U11593 (N_11593,N_11029,N_10582);
nand U11594 (N_11594,N_11085,N_10787);
nor U11595 (N_11595,N_10587,N_10925);
or U11596 (N_11596,N_10647,N_10933);
nand U11597 (N_11597,N_11002,N_10696);
xor U11598 (N_11598,N_10761,N_11223);
nand U11599 (N_11599,N_11075,N_11000);
xnor U11600 (N_11600,N_10766,N_10583);
nand U11601 (N_11601,N_10513,N_10685);
and U11602 (N_11602,N_11218,N_10776);
nor U11603 (N_11603,N_11033,N_11193);
or U11604 (N_11604,N_11077,N_10784);
xnor U11605 (N_11605,N_11122,N_10801);
nor U11606 (N_11606,N_11242,N_10511);
nand U11607 (N_11607,N_10907,N_11240);
nor U11608 (N_11608,N_10954,N_11024);
and U11609 (N_11609,N_11191,N_10649);
or U11610 (N_11610,N_11175,N_10826);
and U11611 (N_11611,N_10672,N_10721);
nand U11612 (N_11612,N_11152,N_10832);
or U11613 (N_11613,N_10798,N_10984);
and U11614 (N_11614,N_10939,N_10723);
nand U11615 (N_11615,N_11042,N_10576);
nand U11616 (N_11616,N_10680,N_11140);
and U11617 (N_11617,N_10500,N_10709);
and U11618 (N_11618,N_10538,N_10783);
nor U11619 (N_11619,N_10834,N_10502);
xnor U11620 (N_11620,N_10736,N_10813);
nand U11621 (N_11621,N_10930,N_11082);
and U11622 (N_11622,N_10617,N_10667);
or U11623 (N_11623,N_11173,N_10759);
nand U11624 (N_11624,N_10863,N_10591);
nor U11625 (N_11625,N_11199,N_10622);
or U11626 (N_11626,N_11098,N_10928);
nand U11627 (N_11627,N_10595,N_11075);
nor U11628 (N_11628,N_10918,N_11102);
nand U11629 (N_11629,N_10633,N_11073);
nand U11630 (N_11630,N_10739,N_10864);
nand U11631 (N_11631,N_10889,N_10566);
and U11632 (N_11632,N_11086,N_10522);
and U11633 (N_11633,N_10952,N_10661);
nand U11634 (N_11634,N_10916,N_10762);
nor U11635 (N_11635,N_10915,N_10948);
nor U11636 (N_11636,N_11023,N_10957);
or U11637 (N_11637,N_11158,N_11081);
xor U11638 (N_11638,N_11206,N_10864);
and U11639 (N_11639,N_10526,N_10545);
nor U11640 (N_11640,N_10746,N_11181);
nor U11641 (N_11641,N_10953,N_10882);
nand U11642 (N_11642,N_10527,N_11155);
nor U11643 (N_11643,N_10541,N_11203);
and U11644 (N_11644,N_10545,N_10940);
xor U11645 (N_11645,N_10765,N_11014);
or U11646 (N_11646,N_10917,N_10943);
nand U11647 (N_11647,N_11100,N_11066);
nor U11648 (N_11648,N_10528,N_10596);
and U11649 (N_11649,N_10851,N_10966);
nand U11650 (N_11650,N_11206,N_10635);
nand U11651 (N_11651,N_11089,N_10525);
xor U11652 (N_11652,N_10996,N_10504);
or U11653 (N_11653,N_11055,N_11038);
nor U11654 (N_11654,N_10905,N_10796);
nor U11655 (N_11655,N_11075,N_10751);
nor U11656 (N_11656,N_10534,N_11230);
and U11657 (N_11657,N_10686,N_10679);
xor U11658 (N_11658,N_10511,N_11202);
xor U11659 (N_11659,N_10704,N_11174);
nor U11660 (N_11660,N_10843,N_11017);
xnor U11661 (N_11661,N_11239,N_10710);
and U11662 (N_11662,N_11071,N_10649);
nand U11663 (N_11663,N_10914,N_10635);
nand U11664 (N_11664,N_10627,N_10793);
nand U11665 (N_11665,N_11135,N_10668);
nor U11666 (N_11666,N_10966,N_10781);
or U11667 (N_11667,N_11210,N_11029);
nor U11668 (N_11668,N_10958,N_11065);
xnor U11669 (N_11669,N_10825,N_11231);
nand U11670 (N_11670,N_10980,N_10582);
and U11671 (N_11671,N_10880,N_10844);
xor U11672 (N_11672,N_10540,N_10810);
and U11673 (N_11673,N_10769,N_11207);
or U11674 (N_11674,N_10536,N_11039);
nand U11675 (N_11675,N_10769,N_10866);
nor U11676 (N_11676,N_10931,N_10718);
or U11677 (N_11677,N_10566,N_10550);
or U11678 (N_11678,N_10616,N_10966);
and U11679 (N_11679,N_10775,N_10903);
or U11680 (N_11680,N_10665,N_10597);
xnor U11681 (N_11681,N_10810,N_10563);
nand U11682 (N_11682,N_10911,N_11067);
nand U11683 (N_11683,N_10915,N_10998);
xnor U11684 (N_11684,N_10754,N_10702);
nand U11685 (N_11685,N_10710,N_10641);
nand U11686 (N_11686,N_11045,N_10944);
or U11687 (N_11687,N_11102,N_10879);
and U11688 (N_11688,N_11042,N_10801);
nor U11689 (N_11689,N_10620,N_11153);
or U11690 (N_11690,N_10903,N_10576);
xnor U11691 (N_11691,N_10578,N_10992);
xnor U11692 (N_11692,N_10853,N_10695);
nand U11693 (N_11693,N_10929,N_10654);
nor U11694 (N_11694,N_10625,N_10513);
nand U11695 (N_11695,N_10777,N_11102);
and U11696 (N_11696,N_11001,N_11249);
nor U11697 (N_11697,N_11075,N_10573);
nand U11698 (N_11698,N_11209,N_10847);
and U11699 (N_11699,N_10630,N_11125);
or U11700 (N_11700,N_10573,N_10791);
xnor U11701 (N_11701,N_10783,N_10521);
or U11702 (N_11702,N_11147,N_10952);
and U11703 (N_11703,N_10545,N_11225);
nand U11704 (N_11704,N_10708,N_11115);
nand U11705 (N_11705,N_10822,N_10880);
nand U11706 (N_11706,N_10720,N_11166);
or U11707 (N_11707,N_11146,N_11103);
nor U11708 (N_11708,N_11165,N_10585);
nand U11709 (N_11709,N_10972,N_10617);
and U11710 (N_11710,N_11110,N_11179);
xor U11711 (N_11711,N_10662,N_10838);
xor U11712 (N_11712,N_10611,N_11193);
and U11713 (N_11713,N_10718,N_11122);
and U11714 (N_11714,N_11153,N_10830);
or U11715 (N_11715,N_10945,N_10897);
and U11716 (N_11716,N_10867,N_10604);
xnor U11717 (N_11717,N_10571,N_11114);
or U11718 (N_11718,N_11023,N_11044);
nand U11719 (N_11719,N_10630,N_10504);
and U11720 (N_11720,N_10944,N_10692);
nor U11721 (N_11721,N_10724,N_10570);
and U11722 (N_11722,N_10792,N_10590);
nand U11723 (N_11723,N_10928,N_10962);
nor U11724 (N_11724,N_10867,N_11200);
xnor U11725 (N_11725,N_11053,N_10627);
xnor U11726 (N_11726,N_10692,N_10851);
and U11727 (N_11727,N_10738,N_11113);
nand U11728 (N_11728,N_10949,N_11040);
xnor U11729 (N_11729,N_10719,N_10894);
nor U11730 (N_11730,N_10955,N_10885);
nand U11731 (N_11731,N_11175,N_10748);
nand U11732 (N_11732,N_10993,N_10945);
xor U11733 (N_11733,N_10650,N_10815);
or U11734 (N_11734,N_10669,N_10990);
nor U11735 (N_11735,N_10723,N_11029);
nand U11736 (N_11736,N_11013,N_11085);
nand U11737 (N_11737,N_10898,N_11189);
xnor U11738 (N_11738,N_11160,N_11187);
xnor U11739 (N_11739,N_11175,N_10664);
or U11740 (N_11740,N_11141,N_11038);
xnor U11741 (N_11741,N_11079,N_10814);
xor U11742 (N_11742,N_10689,N_10710);
xnor U11743 (N_11743,N_10681,N_10542);
or U11744 (N_11744,N_10527,N_10781);
and U11745 (N_11745,N_11078,N_11212);
nand U11746 (N_11746,N_10666,N_11040);
and U11747 (N_11747,N_10796,N_11050);
xor U11748 (N_11748,N_11079,N_11073);
xnor U11749 (N_11749,N_10527,N_10897);
xnor U11750 (N_11750,N_10636,N_10651);
and U11751 (N_11751,N_10757,N_11225);
or U11752 (N_11752,N_10567,N_10512);
xor U11753 (N_11753,N_10964,N_11105);
and U11754 (N_11754,N_11209,N_11105);
nor U11755 (N_11755,N_11068,N_11108);
xnor U11756 (N_11756,N_10824,N_10831);
nor U11757 (N_11757,N_11205,N_10842);
xnor U11758 (N_11758,N_11085,N_10665);
nor U11759 (N_11759,N_10883,N_11182);
nand U11760 (N_11760,N_10872,N_10653);
nor U11761 (N_11761,N_11098,N_10613);
and U11762 (N_11762,N_11123,N_11185);
xnor U11763 (N_11763,N_10690,N_11187);
or U11764 (N_11764,N_11086,N_10821);
nand U11765 (N_11765,N_10508,N_10946);
nand U11766 (N_11766,N_11185,N_11068);
nor U11767 (N_11767,N_10506,N_10835);
or U11768 (N_11768,N_10614,N_10982);
xor U11769 (N_11769,N_11131,N_10935);
nand U11770 (N_11770,N_11100,N_10556);
or U11771 (N_11771,N_10802,N_10707);
xnor U11772 (N_11772,N_11169,N_11045);
nand U11773 (N_11773,N_10653,N_11113);
xnor U11774 (N_11774,N_10563,N_10999);
xor U11775 (N_11775,N_10851,N_10545);
and U11776 (N_11776,N_10507,N_10915);
xnor U11777 (N_11777,N_11067,N_10764);
nand U11778 (N_11778,N_11099,N_10623);
or U11779 (N_11779,N_10668,N_10727);
and U11780 (N_11780,N_10515,N_10586);
and U11781 (N_11781,N_11134,N_10605);
nand U11782 (N_11782,N_10546,N_10945);
nor U11783 (N_11783,N_11169,N_11098);
xnor U11784 (N_11784,N_11101,N_11246);
nor U11785 (N_11785,N_10532,N_11007);
nand U11786 (N_11786,N_10851,N_10971);
nand U11787 (N_11787,N_11013,N_10843);
xor U11788 (N_11788,N_10514,N_11209);
and U11789 (N_11789,N_10913,N_10676);
nor U11790 (N_11790,N_11240,N_10795);
nand U11791 (N_11791,N_11077,N_11147);
nor U11792 (N_11792,N_10574,N_11051);
nand U11793 (N_11793,N_10798,N_11080);
and U11794 (N_11794,N_11244,N_11008);
or U11795 (N_11795,N_10744,N_10873);
xnor U11796 (N_11796,N_10958,N_10878);
nand U11797 (N_11797,N_10682,N_10648);
nand U11798 (N_11798,N_11167,N_11228);
nor U11799 (N_11799,N_11203,N_10879);
or U11800 (N_11800,N_10922,N_10560);
nor U11801 (N_11801,N_10785,N_10537);
or U11802 (N_11802,N_10646,N_11173);
xnor U11803 (N_11803,N_10518,N_10525);
and U11804 (N_11804,N_10549,N_11000);
nand U11805 (N_11805,N_10995,N_10509);
or U11806 (N_11806,N_10632,N_10890);
or U11807 (N_11807,N_10744,N_10677);
nor U11808 (N_11808,N_11026,N_10727);
nand U11809 (N_11809,N_10670,N_10509);
and U11810 (N_11810,N_10849,N_10963);
or U11811 (N_11811,N_10535,N_10953);
and U11812 (N_11812,N_10794,N_10520);
nand U11813 (N_11813,N_10974,N_11215);
or U11814 (N_11814,N_10548,N_10904);
nor U11815 (N_11815,N_10840,N_10773);
nand U11816 (N_11816,N_11027,N_10846);
and U11817 (N_11817,N_10527,N_11194);
nor U11818 (N_11818,N_11095,N_10645);
nand U11819 (N_11819,N_10820,N_10923);
xnor U11820 (N_11820,N_10754,N_10825);
xor U11821 (N_11821,N_11122,N_11166);
or U11822 (N_11822,N_10696,N_10555);
and U11823 (N_11823,N_11032,N_10952);
xor U11824 (N_11824,N_10602,N_10908);
nand U11825 (N_11825,N_10977,N_11153);
xnor U11826 (N_11826,N_10691,N_10780);
xor U11827 (N_11827,N_11176,N_11126);
nand U11828 (N_11828,N_10835,N_10920);
nor U11829 (N_11829,N_10955,N_11183);
nand U11830 (N_11830,N_10971,N_10948);
and U11831 (N_11831,N_10989,N_10616);
nand U11832 (N_11832,N_10618,N_10852);
and U11833 (N_11833,N_11066,N_10553);
nor U11834 (N_11834,N_10602,N_10725);
and U11835 (N_11835,N_10676,N_10542);
nand U11836 (N_11836,N_10949,N_10618);
or U11837 (N_11837,N_10567,N_10715);
nand U11838 (N_11838,N_11181,N_10921);
or U11839 (N_11839,N_11025,N_10760);
xnor U11840 (N_11840,N_10690,N_11133);
or U11841 (N_11841,N_11232,N_10690);
and U11842 (N_11842,N_10830,N_11007);
and U11843 (N_11843,N_10903,N_11169);
nor U11844 (N_11844,N_10808,N_10811);
nor U11845 (N_11845,N_10770,N_11226);
xor U11846 (N_11846,N_11112,N_11006);
xor U11847 (N_11847,N_11233,N_11018);
nor U11848 (N_11848,N_11183,N_10936);
nand U11849 (N_11849,N_10732,N_10749);
nand U11850 (N_11850,N_10823,N_10647);
nor U11851 (N_11851,N_11174,N_11193);
and U11852 (N_11852,N_10871,N_10707);
and U11853 (N_11853,N_10638,N_10944);
xnor U11854 (N_11854,N_10844,N_10980);
and U11855 (N_11855,N_10645,N_11016);
nand U11856 (N_11856,N_11183,N_10575);
and U11857 (N_11857,N_10568,N_10711);
and U11858 (N_11858,N_10594,N_10793);
and U11859 (N_11859,N_10918,N_11106);
nor U11860 (N_11860,N_10999,N_10553);
nor U11861 (N_11861,N_10932,N_10906);
or U11862 (N_11862,N_10625,N_10634);
xnor U11863 (N_11863,N_10705,N_10840);
xor U11864 (N_11864,N_10871,N_10774);
and U11865 (N_11865,N_10842,N_11069);
and U11866 (N_11866,N_11009,N_11126);
or U11867 (N_11867,N_10673,N_10725);
or U11868 (N_11868,N_10649,N_11134);
nand U11869 (N_11869,N_10810,N_10685);
or U11870 (N_11870,N_11192,N_10574);
nand U11871 (N_11871,N_11206,N_10610);
nand U11872 (N_11872,N_11003,N_10665);
and U11873 (N_11873,N_10505,N_11106);
or U11874 (N_11874,N_11028,N_10679);
and U11875 (N_11875,N_10772,N_10902);
and U11876 (N_11876,N_10849,N_11173);
xnor U11877 (N_11877,N_10748,N_10768);
and U11878 (N_11878,N_10516,N_10558);
nor U11879 (N_11879,N_10780,N_10776);
or U11880 (N_11880,N_11074,N_10989);
nor U11881 (N_11881,N_10816,N_10961);
xnor U11882 (N_11882,N_10630,N_10735);
nand U11883 (N_11883,N_10959,N_10915);
xnor U11884 (N_11884,N_10723,N_10678);
nand U11885 (N_11885,N_11031,N_10774);
and U11886 (N_11886,N_10540,N_10669);
or U11887 (N_11887,N_10835,N_10588);
nand U11888 (N_11888,N_10814,N_11137);
or U11889 (N_11889,N_10843,N_10933);
and U11890 (N_11890,N_10914,N_10789);
and U11891 (N_11891,N_11028,N_10741);
nand U11892 (N_11892,N_10903,N_10830);
nand U11893 (N_11893,N_10990,N_10848);
xnor U11894 (N_11894,N_10985,N_11074);
and U11895 (N_11895,N_11111,N_10571);
xnor U11896 (N_11896,N_10841,N_10729);
xnor U11897 (N_11897,N_11175,N_10736);
and U11898 (N_11898,N_10686,N_10777);
xor U11899 (N_11899,N_10890,N_10647);
nor U11900 (N_11900,N_10700,N_11145);
and U11901 (N_11901,N_11096,N_11175);
and U11902 (N_11902,N_10536,N_10730);
and U11903 (N_11903,N_11158,N_11165);
and U11904 (N_11904,N_11152,N_11156);
nor U11905 (N_11905,N_10518,N_10580);
nand U11906 (N_11906,N_10686,N_10612);
and U11907 (N_11907,N_10754,N_10516);
and U11908 (N_11908,N_11135,N_10940);
xnor U11909 (N_11909,N_11158,N_11200);
and U11910 (N_11910,N_11126,N_11164);
xor U11911 (N_11911,N_11095,N_10928);
xor U11912 (N_11912,N_11016,N_10744);
or U11913 (N_11913,N_11029,N_10595);
and U11914 (N_11914,N_10598,N_10920);
and U11915 (N_11915,N_10625,N_10659);
nor U11916 (N_11916,N_11031,N_11223);
and U11917 (N_11917,N_10565,N_11121);
or U11918 (N_11918,N_10748,N_10765);
nand U11919 (N_11919,N_10629,N_11068);
or U11920 (N_11920,N_11011,N_10680);
and U11921 (N_11921,N_11198,N_10715);
xnor U11922 (N_11922,N_11211,N_11226);
xnor U11923 (N_11923,N_11219,N_10950);
nand U11924 (N_11924,N_10619,N_11199);
xor U11925 (N_11925,N_11059,N_10673);
nor U11926 (N_11926,N_10576,N_10591);
and U11927 (N_11927,N_10545,N_11020);
and U11928 (N_11928,N_11230,N_11135);
xor U11929 (N_11929,N_10615,N_11000);
nand U11930 (N_11930,N_11028,N_10600);
and U11931 (N_11931,N_10838,N_10543);
and U11932 (N_11932,N_10523,N_10754);
xnor U11933 (N_11933,N_11224,N_10948);
or U11934 (N_11934,N_11012,N_11225);
nor U11935 (N_11935,N_10607,N_11072);
xor U11936 (N_11936,N_10792,N_11195);
and U11937 (N_11937,N_10540,N_10706);
xor U11938 (N_11938,N_10527,N_11055);
nand U11939 (N_11939,N_10834,N_10542);
xor U11940 (N_11940,N_10819,N_10545);
xnor U11941 (N_11941,N_11018,N_10707);
nor U11942 (N_11942,N_10781,N_11028);
nand U11943 (N_11943,N_11036,N_11076);
or U11944 (N_11944,N_10749,N_10824);
xnor U11945 (N_11945,N_10857,N_10746);
xnor U11946 (N_11946,N_10542,N_11131);
nor U11947 (N_11947,N_11042,N_10852);
and U11948 (N_11948,N_10877,N_11131);
xor U11949 (N_11949,N_10863,N_10803);
nor U11950 (N_11950,N_10886,N_10712);
and U11951 (N_11951,N_10584,N_10894);
and U11952 (N_11952,N_10967,N_10780);
nand U11953 (N_11953,N_10609,N_10922);
nor U11954 (N_11954,N_10581,N_10933);
or U11955 (N_11955,N_10811,N_10568);
xnor U11956 (N_11956,N_10933,N_10682);
nor U11957 (N_11957,N_10582,N_11071);
xnor U11958 (N_11958,N_10634,N_10875);
and U11959 (N_11959,N_10517,N_11059);
or U11960 (N_11960,N_10979,N_10574);
nor U11961 (N_11961,N_10553,N_10704);
nand U11962 (N_11962,N_10942,N_11104);
nor U11963 (N_11963,N_10774,N_10516);
xor U11964 (N_11964,N_10951,N_10597);
nand U11965 (N_11965,N_10948,N_11146);
nand U11966 (N_11966,N_10547,N_10500);
xor U11967 (N_11967,N_10944,N_11197);
or U11968 (N_11968,N_10510,N_11138);
and U11969 (N_11969,N_11245,N_10921);
nand U11970 (N_11970,N_10858,N_10697);
and U11971 (N_11971,N_10954,N_10766);
nor U11972 (N_11972,N_10873,N_11055);
and U11973 (N_11973,N_10796,N_10901);
nand U11974 (N_11974,N_10626,N_10934);
nand U11975 (N_11975,N_10996,N_10596);
nand U11976 (N_11976,N_11025,N_11135);
nor U11977 (N_11977,N_11022,N_10979);
nand U11978 (N_11978,N_11043,N_10633);
xor U11979 (N_11979,N_11004,N_11014);
and U11980 (N_11980,N_10580,N_10782);
and U11981 (N_11981,N_10682,N_11051);
and U11982 (N_11982,N_10775,N_10620);
and U11983 (N_11983,N_10699,N_10778);
nor U11984 (N_11984,N_10612,N_10924);
xor U11985 (N_11985,N_11045,N_11142);
or U11986 (N_11986,N_11030,N_11041);
or U11987 (N_11987,N_10885,N_10691);
nor U11988 (N_11988,N_11082,N_10864);
xor U11989 (N_11989,N_10536,N_10614);
and U11990 (N_11990,N_10800,N_10646);
and U11991 (N_11991,N_11189,N_11006);
nor U11992 (N_11992,N_11060,N_11038);
and U11993 (N_11993,N_10833,N_10696);
nor U11994 (N_11994,N_10824,N_10940);
nand U11995 (N_11995,N_10651,N_10648);
and U11996 (N_11996,N_11220,N_11108);
nor U11997 (N_11997,N_11235,N_11240);
nor U11998 (N_11998,N_10848,N_11033);
nor U11999 (N_11999,N_10507,N_10620);
and U12000 (N_12000,N_11634,N_11781);
xnor U12001 (N_12001,N_11320,N_11463);
and U12002 (N_12002,N_11384,N_11492);
or U12003 (N_12003,N_11616,N_11719);
nor U12004 (N_12004,N_11691,N_11410);
and U12005 (N_12005,N_11847,N_11587);
xor U12006 (N_12006,N_11987,N_11982);
or U12007 (N_12007,N_11403,N_11971);
or U12008 (N_12008,N_11339,N_11367);
nor U12009 (N_12009,N_11498,N_11763);
or U12010 (N_12010,N_11878,N_11440);
nand U12011 (N_12011,N_11362,N_11576);
nand U12012 (N_12012,N_11532,N_11623);
nor U12013 (N_12013,N_11593,N_11882);
or U12014 (N_12014,N_11448,N_11452);
xnor U12015 (N_12015,N_11352,N_11276);
nand U12016 (N_12016,N_11435,N_11891);
nor U12017 (N_12017,N_11743,N_11481);
nand U12018 (N_12018,N_11869,N_11615);
xor U12019 (N_12019,N_11581,N_11553);
nor U12020 (N_12020,N_11827,N_11852);
and U12021 (N_12021,N_11797,N_11890);
xor U12022 (N_12022,N_11810,N_11559);
nor U12023 (N_12023,N_11655,N_11744);
nor U12024 (N_12024,N_11965,N_11329);
xor U12025 (N_12025,N_11288,N_11445);
nand U12026 (N_12026,N_11796,N_11903);
xnor U12027 (N_12027,N_11280,N_11274);
xnor U12028 (N_12028,N_11383,N_11549);
nor U12029 (N_12029,N_11415,N_11446);
xnor U12030 (N_12030,N_11731,N_11281);
nor U12031 (N_12031,N_11487,N_11654);
nand U12032 (N_12032,N_11755,N_11897);
xor U12033 (N_12033,N_11318,N_11583);
nor U12034 (N_12034,N_11727,N_11506);
and U12035 (N_12035,N_11477,N_11911);
and U12036 (N_12036,N_11510,N_11692);
and U12037 (N_12037,N_11525,N_11862);
nand U12038 (N_12038,N_11718,N_11725);
and U12039 (N_12039,N_11759,N_11603);
xor U12040 (N_12040,N_11696,N_11854);
and U12041 (N_12041,N_11292,N_11282);
or U12042 (N_12042,N_11317,N_11360);
nand U12043 (N_12043,N_11838,N_11338);
xor U12044 (N_12044,N_11960,N_11877);
nand U12045 (N_12045,N_11816,N_11527);
nand U12046 (N_12046,N_11646,N_11944);
nand U12047 (N_12047,N_11625,N_11419);
or U12048 (N_12048,N_11613,N_11680);
and U12049 (N_12049,N_11257,N_11904);
or U12050 (N_12050,N_11299,N_11934);
nor U12051 (N_12051,N_11295,N_11437);
xor U12052 (N_12052,N_11704,N_11640);
nor U12053 (N_12053,N_11432,N_11678);
nor U12054 (N_12054,N_11456,N_11520);
and U12055 (N_12055,N_11518,N_11909);
xor U12056 (N_12056,N_11531,N_11547);
nor U12057 (N_12057,N_11756,N_11915);
xnor U12058 (N_12058,N_11961,N_11775);
or U12059 (N_12059,N_11660,N_11735);
and U12060 (N_12060,N_11664,N_11460);
nor U12061 (N_12061,N_11845,N_11373);
nand U12062 (N_12062,N_11426,N_11824);
nand U12063 (N_12063,N_11355,N_11331);
and U12064 (N_12064,N_11697,N_11842);
xor U12065 (N_12065,N_11279,N_11927);
nor U12066 (N_12066,N_11750,N_11289);
xor U12067 (N_12067,N_11720,N_11568);
nor U12068 (N_12068,N_11791,N_11764);
and U12069 (N_12069,N_11895,N_11730);
xnor U12070 (N_12070,N_11689,N_11939);
xnor U12071 (N_12071,N_11873,N_11284);
nand U12072 (N_12072,N_11371,N_11261);
or U12073 (N_12073,N_11267,N_11584);
and U12074 (N_12074,N_11896,N_11993);
and U12075 (N_12075,N_11602,N_11379);
nand U12076 (N_12076,N_11310,N_11918);
and U12077 (N_12077,N_11710,N_11698);
nand U12078 (N_12078,N_11539,N_11429);
and U12079 (N_12079,N_11374,N_11540);
xnor U12080 (N_12080,N_11476,N_11311);
nor U12081 (N_12081,N_11992,N_11496);
or U12082 (N_12082,N_11372,N_11974);
nand U12083 (N_12083,N_11382,N_11685);
or U12084 (N_12084,N_11538,N_11638);
nor U12085 (N_12085,N_11512,N_11332);
or U12086 (N_12086,N_11524,N_11607);
nand U12087 (N_12087,N_11575,N_11416);
nor U12088 (N_12088,N_11790,N_11760);
or U12089 (N_12089,N_11633,N_11832);
nand U12090 (N_12090,N_11434,N_11273);
nor U12091 (N_12091,N_11493,N_11973);
and U12092 (N_12092,N_11464,N_11521);
nand U12093 (N_12093,N_11682,N_11570);
nor U12094 (N_12094,N_11325,N_11666);
or U12095 (N_12095,N_11474,N_11885);
nand U12096 (N_12096,N_11639,N_11565);
and U12097 (N_12097,N_11657,N_11406);
xor U12098 (N_12098,N_11924,N_11899);
xor U12099 (N_12099,N_11359,N_11972);
or U12100 (N_12100,N_11586,N_11999);
nor U12101 (N_12101,N_11275,N_11922);
or U12102 (N_12102,N_11358,N_11344);
nor U12103 (N_12103,N_11612,N_11302);
nand U12104 (N_12104,N_11834,N_11742);
nor U12105 (N_12105,N_11647,N_11370);
nand U12106 (N_12106,N_11536,N_11589);
nor U12107 (N_12107,N_11505,N_11513);
xnor U12108 (N_12108,N_11503,N_11798);
or U12109 (N_12109,N_11622,N_11732);
nor U12110 (N_12110,N_11809,N_11703);
nand U12111 (N_12111,N_11529,N_11928);
nor U12112 (N_12112,N_11699,N_11936);
or U12113 (N_12113,N_11386,N_11541);
nand U12114 (N_12114,N_11908,N_11330);
nor U12115 (N_12115,N_11526,N_11910);
xor U12116 (N_12116,N_11788,N_11938);
nor U12117 (N_12117,N_11572,N_11392);
xnor U12118 (N_12118,N_11687,N_11844);
xnor U12119 (N_12119,N_11659,N_11390);
nand U12120 (N_12120,N_11533,N_11294);
nand U12121 (N_12121,N_11335,N_11945);
nand U12122 (N_12122,N_11876,N_11708);
xnor U12123 (N_12123,N_11767,N_11314);
nor U12124 (N_12124,N_11795,N_11500);
nor U12125 (N_12125,N_11632,N_11679);
nor U12126 (N_12126,N_11431,N_11983);
nor U12127 (N_12127,N_11327,N_11942);
nand U12128 (N_12128,N_11465,N_11511);
xnor U12129 (N_12129,N_11290,N_11480);
nand U12130 (N_12130,N_11291,N_11328);
and U12131 (N_12131,N_11418,N_11887);
nand U12132 (N_12132,N_11316,N_11745);
nand U12133 (N_12133,N_11702,N_11442);
xor U12134 (N_12134,N_11946,N_11979);
or U12135 (N_12135,N_11309,N_11479);
and U12136 (N_12136,N_11658,N_11469);
nor U12137 (N_12137,N_11770,N_11690);
xnor U12138 (N_12138,N_11849,N_11758);
or U12139 (N_12139,N_11780,N_11919);
nand U12140 (N_12140,N_11563,N_11933);
and U12141 (N_12141,N_11669,N_11253);
and U12142 (N_12142,N_11551,N_11571);
or U12143 (N_12143,N_11614,N_11864);
nand U12144 (N_12144,N_11381,N_11629);
nor U12145 (N_12145,N_11305,N_11786);
xor U12146 (N_12146,N_11930,N_11652);
nor U12147 (N_12147,N_11405,N_11557);
or U12148 (N_12148,N_11427,N_11555);
xnor U12149 (N_12149,N_11662,N_11346);
and U12150 (N_12150,N_11857,N_11734);
xnor U12151 (N_12151,N_11817,N_11747);
nor U12152 (N_12152,N_11701,N_11341);
and U12153 (N_12153,N_11969,N_11968);
or U12154 (N_12154,N_11717,N_11507);
xor U12155 (N_12155,N_11298,N_11601);
nand U12156 (N_12156,N_11430,N_11567);
and U12157 (N_12157,N_11837,N_11483);
nor U12158 (N_12158,N_11980,N_11600);
and U12159 (N_12159,N_11272,N_11322);
xnor U12160 (N_12160,N_11884,N_11535);
xnor U12161 (N_12161,N_11313,N_11648);
and U12162 (N_12162,N_11716,N_11892);
nor U12163 (N_12163,N_11765,N_11544);
nand U12164 (N_12164,N_11424,N_11729);
nor U12165 (N_12165,N_11558,N_11254);
and U12166 (N_12166,N_11627,N_11466);
nand U12167 (N_12167,N_11871,N_11843);
xnor U12168 (N_12168,N_11422,N_11604);
nor U12169 (N_12169,N_11588,N_11668);
or U12170 (N_12170,N_11439,N_11663);
and U12171 (N_12171,N_11401,N_11264);
and U12172 (N_12172,N_11619,N_11916);
nand U12173 (N_12173,N_11753,N_11950);
or U12174 (N_12174,N_11516,N_11564);
nand U12175 (N_12175,N_11932,N_11478);
nor U12176 (N_12176,N_11956,N_11994);
and U12177 (N_12177,N_11508,N_11726);
or U12178 (N_12178,N_11577,N_11552);
nor U12179 (N_12179,N_11826,N_11471);
and U12180 (N_12180,N_11265,N_11270);
or U12181 (N_12181,N_11738,N_11417);
nand U12182 (N_12182,N_11721,N_11414);
xnor U12183 (N_12183,N_11863,N_11967);
or U12184 (N_12184,N_11324,N_11262);
xnor U12185 (N_12185,N_11707,N_11782);
and U12186 (N_12186,N_11914,N_11569);
nand U12187 (N_12187,N_11686,N_11777);
nor U12188 (N_12188,N_11955,N_11671);
xor U12189 (N_12189,N_11312,N_11472);
nand U12190 (N_12190,N_11342,N_11473);
or U12191 (N_12191,N_11724,N_11580);
or U12192 (N_12192,N_11917,N_11952);
nor U12193 (N_12193,N_11462,N_11459);
nor U12194 (N_12194,N_11907,N_11772);
nor U12195 (N_12195,N_11369,N_11771);
and U12196 (N_12196,N_11349,N_11436);
nor U12197 (N_12197,N_11672,N_11957);
or U12198 (N_12198,N_11348,N_11562);
and U12199 (N_12199,N_11769,N_11441);
and U12200 (N_12200,N_11598,N_11582);
and U12201 (N_12201,N_11641,N_11811);
and U12202 (N_12202,N_11375,N_11958);
and U12203 (N_12203,N_11399,N_11741);
nand U12204 (N_12204,N_11590,N_11361);
and U12205 (N_12205,N_11684,N_11534);
or U12206 (N_12206,N_11642,N_11393);
or U12207 (N_12207,N_11566,N_11880);
nand U12208 (N_12208,N_11851,N_11398);
nand U12209 (N_12209,N_11617,N_11400);
nand U12210 (N_12210,N_11681,N_11357);
xor U12211 (N_12211,N_11898,N_11548);
nand U12212 (N_12212,N_11256,N_11605);
nand U12213 (N_12213,N_11250,N_11785);
xnor U12214 (N_12214,N_11461,N_11943);
or U12215 (N_12215,N_11740,N_11906);
xnor U12216 (N_12216,N_11776,N_11951);
nand U12217 (N_12217,N_11948,N_11509);
or U12218 (N_12218,N_11978,N_11976);
or U12219 (N_12219,N_11488,N_11902);
xnor U12220 (N_12220,N_11825,N_11920);
nor U12221 (N_12221,N_11653,N_11783);
or U12222 (N_12222,N_11709,N_11859);
and U12223 (N_12223,N_11792,N_11636);
or U12224 (N_12224,N_11395,N_11836);
nand U12225 (N_12225,N_11829,N_11501);
xnor U12226 (N_12226,N_11484,N_11964);
and U12227 (N_12227,N_11301,N_11323);
and U12228 (N_12228,N_11300,N_11304);
nand U12229 (N_12229,N_11443,N_11841);
xor U12230 (N_12230,N_11793,N_11977);
and U12231 (N_12231,N_11814,N_11807);
nor U12232 (N_12232,N_11773,N_11411);
nor U12233 (N_12233,N_11283,N_11888);
xor U12234 (N_12234,N_11347,N_11468);
nor U12235 (N_12235,N_11818,N_11271);
nor U12236 (N_12236,N_11768,N_11597);
nor U12237 (N_12237,N_11789,N_11326);
nand U12238 (N_12238,N_11447,N_11855);
or U12239 (N_12239,N_11819,N_11450);
xnor U12240 (N_12240,N_11277,N_11990);
or U12241 (N_12241,N_11364,N_11444);
xor U12242 (N_12242,N_11308,N_11475);
nor U12243 (N_12243,N_11423,N_11988);
or U12244 (N_12244,N_11428,N_11656);
or U12245 (N_12245,N_11886,N_11799);
nor U12246 (N_12246,N_11353,N_11438);
or U12247 (N_12247,N_11421,N_11365);
and U12248 (N_12248,N_11751,N_11592);
nor U12249 (N_12249,N_11561,N_11389);
nand U12250 (N_12250,N_11801,N_11453);
nor U12251 (N_12251,N_11846,N_11608);
nor U12252 (N_12252,N_11545,N_11356);
xor U12253 (N_12253,N_11947,N_11787);
xor U12254 (N_12254,N_11949,N_11839);
nand U12255 (N_12255,N_11853,N_11611);
nand U12256 (N_12256,N_11805,N_11251);
nand U12257 (N_12257,N_11591,N_11391);
nand U12258 (N_12258,N_11307,N_11490);
nor U12259 (N_12259,N_11675,N_11850);
and U12260 (N_12260,N_11560,N_11454);
nor U12261 (N_12261,N_11351,N_11865);
nor U12262 (N_12262,N_11748,N_11644);
and U12263 (N_12263,N_11645,N_11812);
nand U12264 (N_12264,N_11989,N_11778);
nor U12265 (N_12265,N_11749,N_11746);
and U12266 (N_12266,N_11766,N_11667);
xnor U12267 (N_12267,N_11806,N_11981);
nor U12268 (N_12268,N_11828,N_11676);
and U12269 (N_12269,N_11991,N_11334);
or U12270 (N_12270,N_11931,N_11624);
xor U12271 (N_12271,N_11269,N_11752);
or U12272 (N_12272,N_11861,N_11815);
nand U12273 (N_12273,N_11350,N_11550);
nor U12274 (N_12274,N_11670,N_11985);
nand U12275 (N_12275,N_11673,N_11954);
and U12276 (N_12276,N_11628,N_11574);
and U12277 (N_12277,N_11519,N_11396);
xnor U12278 (N_12278,N_11523,N_11986);
or U12279 (N_12279,N_11620,N_11883);
or U12280 (N_12280,N_11706,N_11802);
or U12281 (N_12281,N_11711,N_11820);
nand U12282 (N_12282,N_11556,N_11306);
nor U12283 (N_12283,N_11485,N_11984);
and U12284 (N_12284,N_11831,N_11366);
nand U12285 (N_12285,N_11813,N_11585);
and U12286 (N_12286,N_11333,N_11941);
nor U12287 (N_12287,N_11996,N_11926);
nand U12288 (N_12288,N_11595,N_11966);
nand U12289 (N_12289,N_11542,N_11683);
xor U12290 (N_12290,N_11925,N_11579);
or U12291 (N_12291,N_11970,N_11467);
nand U12292 (N_12292,N_11499,N_11303);
nor U12293 (N_12293,N_11998,N_11821);
nor U12294 (N_12294,N_11997,N_11959);
nand U12295 (N_12295,N_11804,N_11263);
or U12296 (N_12296,N_11975,N_11953);
and U12297 (N_12297,N_11377,N_11594);
nand U12298 (N_12298,N_11402,N_11340);
xnor U12299 (N_12299,N_11694,N_11455);
xnor U12300 (N_12300,N_11923,N_11894);
or U12301 (N_12301,N_11722,N_11693);
xnor U12302 (N_12302,N_11808,N_11266);
xnor U12303 (N_12303,N_11626,N_11757);
xnor U12304 (N_12304,N_11537,N_11268);
nand U12305 (N_12305,N_11293,N_11610);
or U12306 (N_12306,N_11433,N_11259);
nand U12307 (N_12307,N_11252,N_11762);
and U12308 (N_12308,N_11912,N_11573);
nand U12309 (N_12309,N_11995,N_11315);
nor U12310 (N_12310,N_11502,N_11631);
and U12311 (N_12311,N_11833,N_11287);
and U12312 (N_12312,N_11286,N_11700);
xnor U12313 (N_12313,N_11409,N_11387);
nor U12314 (N_12314,N_11874,N_11840);
or U12315 (N_12315,N_11354,N_11457);
or U12316 (N_12316,N_11803,N_11794);
and U12317 (N_12317,N_11866,N_11528);
xor U12318 (N_12318,N_11856,N_11630);
nand U12319 (N_12319,N_11870,N_11337);
xor U12320 (N_12320,N_11394,N_11296);
or U12321 (N_12321,N_11935,N_11345);
or U12322 (N_12322,N_11260,N_11723);
or U12323 (N_12323,N_11385,N_11258);
or U12324 (N_12324,N_11835,N_11712);
nor U12325 (N_12325,N_11578,N_11733);
xnor U12326 (N_12326,N_11449,N_11297);
and U12327 (N_12327,N_11650,N_11661);
nor U12328 (N_12328,N_11860,N_11278);
or U12329 (N_12329,N_11913,N_11368);
xnor U12330 (N_12330,N_11881,N_11522);
nor U12331 (N_12331,N_11737,N_11921);
or U12332 (N_12332,N_11889,N_11495);
nor U12333 (N_12333,N_11497,N_11517);
nand U12334 (N_12334,N_11397,N_11530);
nand U12335 (N_12335,N_11713,N_11800);
nor U12336 (N_12336,N_11875,N_11714);
and U12337 (N_12337,N_11319,N_11491);
or U12338 (N_12338,N_11482,N_11779);
and U12339 (N_12339,N_11546,N_11515);
and U12340 (N_12340,N_11425,N_11754);
nor U12341 (N_12341,N_11940,N_11867);
nor U12342 (N_12342,N_11901,N_11695);
xnor U12343 (N_12343,N_11336,N_11736);
nor U12344 (N_12344,N_11688,N_11879);
nor U12345 (N_12345,N_11774,N_11929);
nor U12346 (N_12346,N_11408,N_11677);
nor U12347 (N_12347,N_11514,N_11285);
nand U12348 (N_12348,N_11893,N_11458);
nor U12349 (N_12349,N_11413,N_11651);
nor U12350 (N_12350,N_11665,N_11380);
or U12351 (N_12351,N_11255,N_11900);
xor U12352 (N_12352,N_11376,N_11599);
or U12353 (N_12353,N_11858,N_11822);
nand U12354 (N_12354,N_11872,N_11363);
nor U12355 (N_12355,N_11962,N_11486);
or U12356 (N_12356,N_11378,N_11618);
or U12357 (N_12357,N_11470,N_11635);
and U12358 (N_12358,N_11784,N_11637);
xor U12359 (N_12359,N_11543,N_11823);
nand U12360 (N_12360,N_11905,N_11321);
nor U12361 (N_12361,N_11606,N_11848);
xor U12362 (N_12362,N_11609,N_11412);
and U12363 (N_12363,N_11404,N_11761);
or U12364 (N_12364,N_11451,N_11830);
or U12365 (N_12365,N_11504,N_11621);
nor U12366 (N_12366,N_11343,N_11937);
and U12367 (N_12367,N_11674,N_11388);
and U12368 (N_12368,N_11715,N_11649);
nand U12369 (N_12369,N_11739,N_11705);
xor U12370 (N_12370,N_11963,N_11554);
nor U12371 (N_12371,N_11407,N_11489);
or U12372 (N_12372,N_11596,N_11728);
nand U12373 (N_12373,N_11643,N_11420);
xnor U12374 (N_12374,N_11868,N_11494);
xor U12375 (N_12375,N_11713,N_11681);
nor U12376 (N_12376,N_11788,N_11342);
or U12377 (N_12377,N_11306,N_11740);
or U12378 (N_12378,N_11436,N_11583);
nor U12379 (N_12379,N_11882,N_11474);
nand U12380 (N_12380,N_11282,N_11585);
nand U12381 (N_12381,N_11806,N_11828);
xnor U12382 (N_12382,N_11259,N_11378);
nor U12383 (N_12383,N_11702,N_11342);
nand U12384 (N_12384,N_11482,N_11870);
nand U12385 (N_12385,N_11710,N_11482);
or U12386 (N_12386,N_11726,N_11500);
or U12387 (N_12387,N_11332,N_11513);
nor U12388 (N_12388,N_11631,N_11918);
xnor U12389 (N_12389,N_11679,N_11941);
and U12390 (N_12390,N_11356,N_11965);
nand U12391 (N_12391,N_11403,N_11668);
xnor U12392 (N_12392,N_11755,N_11927);
xor U12393 (N_12393,N_11762,N_11302);
nand U12394 (N_12394,N_11567,N_11309);
and U12395 (N_12395,N_11980,N_11771);
or U12396 (N_12396,N_11924,N_11942);
nor U12397 (N_12397,N_11754,N_11841);
and U12398 (N_12398,N_11476,N_11796);
and U12399 (N_12399,N_11267,N_11393);
or U12400 (N_12400,N_11901,N_11724);
nor U12401 (N_12401,N_11495,N_11917);
and U12402 (N_12402,N_11705,N_11392);
xor U12403 (N_12403,N_11594,N_11506);
nor U12404 (N_12404,N_11619,N_11466);
or U12405 (N_12405,N_11851,N_11677);
nor U12406 (N_12406,N_11672,N_11468);
nand U12407 (N_12407,N_11599,N_11809);
xnor U12408 (N_12408,N_11970,N_11950);
nor U12409 (N_12409,N_11709,N_11872);
and U12410 (N_12410,N_11754,N_11638);
and U12411 (N_12411,N_11994,N_11609);
or U12412 (N_12412,N_11361,N_11931);
nor U12413 (N_12413,N_11641,N_11474);
xor U12414 (N_12414,N_11717,N_11519);
nor U12415 (N_12415,N_11459,N_11553);
nor U12416 (N_12416,N_11791,N_11692);
and U12417 (N_12417,N_11632,N_11507);
and U12418 (N_12418,N_11937,N_11420);
nand U12419 (N_12419,N_11471,N_11735);
or U12420 (N_12420,N_11286,N_11520);
and U12421 (N_12421,N_11487,N_11941);
or U12422 (N_12422,N_11778,N_11774);
xnor U12423 (N_12423,N_11755,N_11373);
nor U12424 (N_12424,N_11984,N_11365);
or U12425 (N_12425,N_11999,N_11604);
xnor U12426 (N_12426,N_11639,N_11598);
nand U12427 (N_12427,N_11425,N_11490);
nand U12428 (N_12428,N_11645,N_11550);
or U12429 (N_12429,N_11584,N_11947);
nor U12430 (N_12430,N_11278,N_11279);
xor U12431 (N_12431,N_11990,N_11463);
xor U12432 (N_12432,N_11312,N_11988);
or U12433 (N_12433,N_11349,N_11949);
or U12434 (N_12434,N_11830,N_11711);
nand U12435 (N_12435,N_11645,N_11733);
and U12436 (N_12436,N_11624,N_11383);
nor U12437 (N_12437,N_11320,N_11605);
or U12438 (N_12438,N_11452,N_11757);
nand U12439 (N_12439,N_11757,N_11469);
nor U12440 (N_12440,N_11515,N_11993);
nand U12441 (N_12441,N_11359,N_11862);
nand U12442 (N_12442,N_11769,N_11344);
or U12443 (N_12443,N_11474,N_11338);
and U12444 (N_12444,N_11543,N_11270);
nand U12445 (N_12445,N_11688,N_11575);
or U12446 (N_12446,N_11454,N_11361);
nand U12447 (N_12447,N_11944,N_11691);
or U12448 (N_12448,N_11862,N_11841);
and U12449 (N_12449,N_11404,N_11340);
or U12450 (N_12450,N_11360,N_11616);
nor U12451 (N_12451,N_11435,N_11344);
nand U12452 (N_12452,N_11291,N_11507);
or U12453 (N_12453,N_11491,N_11966);
nor U12454 (N_12454,N_11352,N_11424);
nor U12455 (N_12455,N_11558,N_11392);
xnor U12456 (N_12456,N_11701,N_11331);
nor U12457 (N_12457,N_11277,N_11420);
nor U12458 (N_12458,N_11292,N_11665);
or U12459 (N_12459,N_11338,N_11477);
or U12460 (N_12460,N_11893,N_11767);
xor U12461 (N_12461,N_11708,N_11527);
xnor U12462 (N_12462,N_11460,N_11266);
or U12463 (N_12463,N_11751,N_11360);
nand U12464 (N_12464,N_11856,N_11783);
nor U12465 (N_12465,N_11642,N_11612);
nor U12466 (N_12466,N_11669,N_11350);
and U12467 (N_12467,N_11381,N_11791);
nand U12468 (N_12468,N_11569,N_11340);
or U12469 (N_12469,N_11665,N_11864);
xnor U12470 (N_12470,N_11270,N_11906);
or U12471 (N_12471,N_11392,N_11391);
nand U12472 (N_12472,N_11803,N_11487);
or U12473 (N_12473,N_11951,N_11372);
or U12474 (N_12474,N_11889,N_11971);
nor U12475 (N_12475,N_11773,N_11448);
or U12476 (N_12476,N_11653,N_11400);
and U12477 (N_12477,N_11473,N_11607);
xor U12478 (N_12478,N_11439,N_11710);
or U12479 (N_12479,N_11613,N_11997);
or U12480 (N_12480,N_11359,N_11282);
and U12481 (N_12481,N_11689,N_11539);
nand U12482 (N_12482,N_11966,N_11715);
nand U12483 (N_12483,N_11834,N_11580);
and U12484 (N_12484,N_11741,N_11662);
nor U12485 (N_12485,N_11859,N_11751);
nor U12486 (N_12486,N_11435,N_11661);
or U12487 (N_12487,N_11959,N_11830);
xnor U12488 (N_12488,N_11454,N_11358);
xnor U12489 (N_12489,N_11672,N_11534);
or U12490 (N_12490,N_11747,N_11304);
xnor U12491 (N_12491,N_11851,N_11692);
and U12492 (N_12492,N_11944,N_11344);
and U12493 (N_12493,N_11745,N_11449);
and U12494 (N_12494,N_11770,N_11778);
and U12495 (N_12495,N_11347,N_11388);
xnor U12496 (N_12496,N_11997,N_11589);
or U12497 (N_12497,N_11433,N_11465);
nor U12498 (N_12498,N_11618,N_11990);
nor U12499 (N_12499,N_11850,N_11659);
or U12500 (N_12500,N_11829,N_11998);
or U12501 (N_12501,N_11755,N_11578);
or U12502 (N_12502,N_11928,N_11893);
nand U12503 (N_12503,N_11337,N_11724);
or U12504 (N_12504,N_11350,N_11996);
xnor U12505 (N_12505,N_11573,N_11424);
nand U12506 (N_12506,N_11939,N_11601);
nor U12507 (N_12507,N_11932,N_11616);
nand U12508 (N_12508,N_11456,N_11429);
nor U12509 (N_12509,N_11695,N_11802);
nand U12510 (N_12510,N_11506,N_11884);
nand U12511 (N_12511,N_11492,N_11470);
xor U12512 (N_12512,N_11500,N_11355);
nor U12513 (N_12513,N_11662,N_11338);
nand U12514 (N_12514,N_11794,N_11263);
and U12515 (N_12515,N_11749,N_11479);
or U12516 (N_12516,N_11345,N_11899);
xnor U12517 (N_12517,N_11531,N_11629);
nor U12518 (N_12518,N_11292,N_11540);
xor U12519 (N_12519,N_11526,N_11485);
xor U12520 (N_12520,N_11271,N_11715);
nand U12521 (N_12521,N_11768,N_11250);
nand U12522 (N_12522,N_11399,N_11630);
nand U12523 (N_12523,N_11790,N_11649);
or U12524 (N_12524,N_11356,N_11345);
nor U12525 (N_12525,N_11349,N_11978);
xor U12526 (N_12526,N_11874,N_11331);
nor U12527 (N_12527,N_11346,N_11527);
xnor U12528 (N_12528,N_11362,N_11822);
and U12529 (N_12529,N_11736,N_11334);
and U12530 (N_12530,N_11362,N_11671);
nor U12531 (N_12531,N_11779,N_11319);
and U12532 (N_12532,N_11439,N_11732);
xor U12533 (N_12533,N_11277,N_11939);
nand U12534 (N_12534,N_11900,N_11764);
and U12535 (N_12535,N_11386,N_11844);
xnor U12536 (N_12536,N_11816,N_11656);
xnor U12537 (N_12537,N_11608,N_11814);
nor U12538 (N_12538,N_11581,N_11750);
and U12539 (N_12539,N_11517,N_11544);
nor U12540 (N_12540,N_11853,N_11808);
nand U12541 (N_12541,N_11979,N_11575);
and U12542 (N_12542,N_11873,N_11905);
nor U12543 (N_12543,N_11676,N_11613);
nor U12544 (N_12544,N_11333,N_11485);
and U12545 (N_12545,N_11380,N_11458);
and U12546 (N_12546,N_11919,N_11719);
xor U12547 (N_12547,N_11874,N_11759);
or U12548 (N_12548,N_11280,N_11739);
nor U12549 (N_12549,N_11694,N_11930);
nor U12550 (N_12550,N_11683,N_11424);
and U12551 (N_12551,N_11511,N_11471);
xor U12552 (N_12552,N_11609,N_11934);
nor U12553 (N_12553,N_11591,N_11963);
or U12554 (N_12554,N_11371,N_11825);
xnor U12555 (N_12555,N_11691,N_11829);
nand U12556 (N_12556,N_11626,N_11558);
or U12557 (N_12557,N_11279,N_11994);
xnor U12558 (N_12558,N_11509,N_11365);
nor U12559 (N_12559,N_11989,N_11549);
nand U12560 (N_12560,N_11581,N_11283);
and U12561 (N_12561,N_11877,N_11980);
or U12562 (N_12562,N_11671,N_11888);
nand U12563 (N_12563,N_11364,N_11331);
nor U12564 (N_12564,N_11961,N_11708);
xnor U12565 (N_12565,N_11495,N_11566);
nand U12566 (N_12566,N_11656,N_11996);
or U12567 (N_12567,N_11692,N_11486);
xor U12568 (N_12568,N_11358,N_11254);
and U12569 (N_12569,N_11517,N_11389);
or U12570 (N_12570,N_11310,N_11578);
or U12571 (N_12571,N_11906,N_11969);
nand U12572 (N_12572,N_11701,N_11492);
and U12573 (N_12573,N_11570,N_11906);
or U12574 (N_12574,N_11382,N_11391);
and U12575 (N_12575,N_11631,N_11822);
and U12576 (N_12576,N_11859,N_11284);
and U12577 (N_12577,N_11702,N_11767);
or U12578 (N_12578,N_11997,N_11511);
nor U12579 (N_12579,N_11930,N_11763);
and U12580 (N_12580,N_11842,N_11611);
xor U12581 (N_12581,N_11875,N_11399);
or U12582 (N_12582,N_11301,N_11489);
nor U12583 (N_12583,N_11945,N_11618);
xnor U12584 (N_12584,N_11453,N_11316);
and U12585 (N_12585,N_11636,N_11927);
xor U12586 (N_12586,N_11274,N_11256);
and U12587 (N_12587,N_11701,N_11967);
or U12588 (N_12588,N_11797,N_11253);
xnor U12589 (N_12589,N_11999,N_11667);
nor U12590 (N_12590,N_11776,N_11997);
or U12591 (N_12591,N_11638,N_11401);
nor U12592 (N_12592,N_11941,N_11940);
and U12593 (N_12593,N_11267,N_11262);
or U12594 (N_12594,N_11755,N_11253);
and U12595 (N_12595,N_11870,N_11397);
and U12596 (N_12596,N_11748,N_11554);
nand U12597 (N_12597,N_11520,N_11615);
or U12598 (N_12598,N_11740,N_11918);
and U12599 (N_12599,N_11549,N_11640);
xnor U12600 (N_12600,N_11588,N_11633);
nor U12601 (N_12601,N_11776,N_11432);
or U12602 (N_12602,N_11934,N_11787);
nand U12603 (N_12603,N_11726,N_11625);
or U12604 (N_12604,N_11702,N_11659);
nand U12605 (N_12605,N_11761,N_11377);
nand U12606 (N_12606,N_11281,N_11954);
nor U12607 (N_12607,N_11707,N_11287);
xnor U12608 (N_12608,N_11281,N_11874);
xor U12609 (N_12609,N_11475,N_11725);
or U12610 (N_12610,N_11257,N_11803);
nor U12611 (N_12611,N_11653,N_11405);
nand U12612 (N_12612,N_11870,N_11737);
or U12613 (N_12613,N_11864,N_11730);
and U12614 (N_12614,N_11307,N_11529);
and U12615 (N_12615,N_11499,N_11301);
xnor U12616 (N_12616,N_11523,N_11830);
and U12617 (N_12617,N_11332,N_11601);
and U12618 (N_12618,N_11401,N_11458);
nor U12619 (N_12619,N_11674,N_11771);
nor U12620 (N_12620,N_11714,N_11695);
nand U12621 (N_12621,N_11281,N_11633);
and U12622 (N_12622,N_11991,N_11863);
nor U12623 (N_12623,N_11303,N_11273);
or U12624 (N_12624,N_11285,N_11710);
nor U12625 (N_12625,N_11650,N_11885);
and U12626 (N_12626,N_11430,N_11621);
and U12627 (N_12627,N_11935,N_11650);
nor U12628 (N_12628,N_11536,N_11254);
and U12629 (N_12629,N_11656,N_11693);
xor U12630 (N_12630,N_11701,N_11539);
xnor U12631 (N_12631,N_11299,N_11952);
nand U12632 (N_12632,N_11868,N_11359);
nor U12633 (N_12633,N_11870,N_11253);
or U12634 (N_12634,N_11841,N_11295);
nor U12635 (N_12635,N_11749,N_11925);
nor U12636 (N_12636,N_11624,N_11491);
and U12637 (N_12637,N_11455,N_11557);
nor U12638 (N_12638,N_11289,N_11532);
xnor U12639 (N_12639,N_11684,N_11837);
and U12640 (N_12640,N_11315,N_11579);
nor U12641 (N_12641,N_11877,N_11340);
xnor U12642 (N_12642,N_11279,N_11783);
and U12643 (N_12643,N_11458,N_11574);
or U12644 (N_12644,N_11922,N_11486);
nor U12645 (N_12645,N_11473,N_11717);
and U12646 (N_12646,N_11365,N_11741);
or U12647 (N_12647,N_11488,N_11422);
nor U12648 (N_12648,N_11741,N_11714);
xnor U12649 (N_12649,N_11751,N_11911);
nor U12650 (N_12650,N_11509,N_11573);
nor U12651 (N_12651,N_11282,N_11823);
nand U12652 (N_12652,N_11743,N_11537);
and U12653 (N_12653,N_11764,N_11556);
nor U12654 (N_12654,N_11352,N_11474);
nand U12655 (N_12655,N_11878,N_11581);
nand U12656 (N_12656,N_11484,N_11726);
nand U12657 (N_12657,N_11758,N_11280);
and U12658 (N_12658,N_11518,N_11396);
or U12659 (N_12659,N_11997,N_11660);
nand U12660 (N_12660,N_11789,N_11307);
or U12661 (N_12661,N_11263,N_11452);
nor U12662 (N_12662,N_11910,N_11718);
nand U12663 (N_12663,N_11266,N_11595);
or U12664 (N_12664,N_11903,N_11729);
nand U12665 (N_12665,N_11369,N_11980);
xor U12666 (N_12666,N_11954,N_11365);
nor U12667 (N_12667,N_11343,N_11544);
nor U12668 (N_12668,N_11277,N_11599);
or U12669 (N_12669,N_11626,N_11963);
or U12670 (N_12670,N_11744,N_11822);
nand U12671 (N_12671,N_11382,N_11915);
nor U12672 (N_12672,N_11261,N_11916);
xor U12673 (N_12673,N_11627,N_11746);
nand U12674 (N_12674,N_11570,N_11900);
and U12675 (N_12675,N_11294,N_11431);
and U12676 (N_12676,N_11447,N_11838);
nor U12677 (N_12677,N_11875,N_11712);
nand U12678 (N_12678,N_11571,N_11627);
nor U12679 (N_12679,N_11914,N_11338);
or U12680 (N_12680,N_11261,N_11445);
nand U12681 (N_12681,N_11555,N_11840);
nand U12682 (N_12682,N_11423,N_11866);
xor U12683 (N_12683,N_11853,N_11541);
and U12684 (N_12684,N_11302,N_11573);
and U12685 (N_12685,N_11758,N_11888);
nor U12686 (N_12686,N_11627,N_11861);
and U12687 (N_12687,N_11843,N_11786);
or U12688 (N_12688,N_11322,N_11832);
nor U12689 (N_12689,N_11309,N_11773);
nor U12690 (N_12690,N_11670,N_11653);
and U12691 (N_12691,N_11729,N_11791);
nor U12692 (N_12692,N_11679,N_11947);
nor U12693 (N_12693,N_11344,N_11841);
nor U12694 (N_12694,N_11504,N_11934);
nor U12695 (N_12695,N_11796,N_11504);
nand U12696 (N_12696,N_11672,N_11972);
or U12697 (N_12697,N_11677,N_11672);
xor U12698 (N_12698,N_11433,N_11792);
and U12699 (N_12699,N_11329,N_11292);
nand U12700 (N_12700,N_11592,N_11782);
xor U12701 (N_12701,N_11814,N_11702);
nor U12702 (N_12702,N_11730,N_11603);
nor U12703 (N_12703,N_11418,N_11443);
nand U12704 (N_12704,N_11491,N_11533);
and U12705 (N_12705,N_11778,N_11336);
or U12706 (N_12706,N_11492,N_11733);
nor U12707 (N_12707,N_11996,N_11690);
xor U12708 (N_12708,N_11315,N_11516);
xnor U12709 (N_12709,N_11905,N_11806);
nor U12710 (N_12710,N_11513,N_11937);
xor U12711 (N_12711,N_11361,N_11919);
nand U12712 (N_12712,N_11763,N_11267);
xor U12713 (N_12713,N_11956,N_11468);
xnor U12714 (N_12714,N_11870,N_11969);
and U12715 (N_12715,N_11446,N_11400);
and U12716 (N_12716,N_11396,N_11297);
xnor U12717 (N_12717,N_11641,N_11971);
nand U12718 (N_12718,N_11331,N_11926);
nor U12719 (N_12719,N_11926,N_11862);
or U12720 (N_12720,N_11343,N_11933);
xnor U12721 (N_12721,N_11733,N_11362);
and U12722 (N_12722,N_11765,N_11285);
nor U12723 (N_12723,N_11720,N_11302);
xor U12724 (N_12724,N_11290,N_11857);
xor U12725 (N_12725,N_11271,N_11376);
or U12726 (N_12726,N_11458,N_11664);
nor U12727 (N_12727,N_11426,N_11855);
nor U12728 (N_12728,N_11913,N_11781);
nand U12729 (N_12729,N_11696,N_11978);
nand U12730 (N_12730,N_11472,N_11931);
and U12731 (N_12731,N_11393,N_11483);
nand U12732 (N_12732,N_11702,N_11480);
xnor U12733 (N_12733,N_11596,N_11646);
or U12734 (N_12734,N_11351,N_11500);
nand U12735 (N_12735,N_11717,N_11544);
nor U12736 (N_12736,N_11722,N_11532);
or U12737 (N_12737,N_11507,N_11784);
nand U12738 (N_12738,N_11600,N_11275);
or U12739 (N_12739,N_11276,N_11982);
xnor U12740 (N_12740,N_11365,N_11826);
xnor U12741 (N_12741,N_11705,N_11301);
xnor U12742 (N_12742,N_11404,N_11994);
nor U12743 (N_12743,N_11856,N_11969);
and U12744 (N_12744,N_11433,N_11575);
nor U12745 (N_12745,N_11881,N_11630);
and U12746 (N_12746,N_11745,N_11423);
nor U12747 (N_12747,N_11999,N_11600);
nor U12748 (N_12748,N_11406,N_11644);
nand U12749 (N_12749,N_11961,N_11329);
xor U12750 (N_12750,N_12345,N_12654);
and U12751 (N_12751,N_12462,N_12004);
or U12752 (N_12752,N_12367,N_12124);
xnor U12753 (N_12753,N_12439,N_12500);
nor U12754 (N_12754,N_12475,N_12363);
and U12755 (N_12755,N_12246,N_12626);
xnor U12756 (N_12756,N_12720,N_12446);
nand U12757 (N_12757,N_12185,N_12158);
nand U12758 (N_12758,N_12703,N_12073);
nand U12759 (N_12759,N_12445,N_12061);
xnor U12760 (N_12760,N_12447,N_12143);
and U12761 (N_12761,N_12564,N_12660);
and U12762 (N_12762,N_12369,N_12324);
nor U12763 (N_12763,N_12016,N_12540);
and U12764 (N_12764,N_12274,N_12681);
and U12765 (N_12765,N_12116,N_12410);
xnor U12766 (N_12766,N_12043,N_12019);
or U12767 (N_12767,N_12227,N_12258);
and U12768 (N_12768,N_12294,N_12391);
or U12769 (N_12769,N_12642,N_12068);
xnor U12770 (N_12770,N_12476,N_12286);
xor U12771 (N_12771,N_12543,N_12589);
xor U12772 (N_12772,N_12408,N_12177);
nor U12773 (N_12773,N_12449,N_12658);
nor U12774 (N_12774,N_12146,N_12747);
and U12775 (N_12775,N_12222,N_12514);
and U12776 (N_12776,N_12047,N_12269);
or U12777 (N_12777,N_12452,N_12416);
nand U12778 (N_12778,N_12678,N_12194);
xnor U12779 (N_12779,N_12189,N_12226);
xor U12780 (N_12780,N_12717,N_12080);
nor U12781 (N_12781,N_12198,N_12440);
and U12782 (N_12782,N_12022,N_12078);
nand U12783 (N_12783,N_12549,N_12238);
nand U12784 (N_12784,N_12157,N_12118);
and U12785 (N_12785,N_12620,N_12316);
nand U12786 (N_12786,N_12457,N_12516);
or U12787 (N_12787,N_12154,N_12127);
xor U12788 (N_12788,N_12507,N_12045);
and U12789 (N_12789,N_12242,N_12743);
nand U12790 (N_12790,N_12322,N_12611);
nor U12791 (N_12791,N_12663,N_12305);
and U12792 (N_12792,N_12577,N_12210);
nand U12793 (N_12793,N_12147,N_12382);
xnor U12794 (N_12794,N_12072,N_12052);
nor U12795 (N_12795,N_12539,N_12706);
xnor U12796 (N_12796,N_12314,N_12368);
or U12797 (N_12797,N_12005,N_12285);
and U12798 (N_12798,N_12437,N_12132);
nor U12799 (N_12799,N_12114,N_12737);
xnor U12800 (N_12800,N_12596,N_12380);
nor U12801 (N_12801,N_12166,N_12326);
nor U12802 (N_12802,N_12217,N_12579);
xnor U12803 (N_12803,N_12234,N_12694);
and U12804 (N_12804,N_12644,N_12599);
nand U12805 (N_12805,N_12551,N_12290);
and U12806 (N_12806,N_12035,N_12267);
nand U12807 (N_12807,N_12713,N_12602);
and U12808 (N_12808,N_12438,N_12473);
and U12809 (N_12809,N_12536,N_12104);
nor U12810 (N_12810,N_12635,N_12183);
and U12811 (N_12811,N_12586,N_12397);
and U12812 (N_12812,N_12734,N_12089);
xor U12813 (N_12813,N_12372,N_12188);
nand U12814 (N_12814,N_12745,N_12303);
or U12815 (N_12815,N_12423,N_12701);
xnor U12816 (N_12816,N_12253,N_12575);
or U12817 (N_12817,N_12548,N_12235);
or U12818 (N_12818,N_12527,N_12574);
or U12819 (N_12819,N_12361,N_12311);
or U12820 (N_12820,N_12524,N_12265);
xnor U12821 (N_12821,N_12392,N_12230);
or U12822 (N_12822,N_12174,N_12732);
nor U12823 (N_12823,N_12276,N_12386);
nor U12824 (N_12824,N_12465,N_12622);
or U12825 (N_12825,N_12101,N_12531);
and U12826 (N_12826,N_12337,N_12339);
xor U12827 (N_12827,N_12150,N_12130);
xnor U12828 (N_12828,N_12280,N_12606);
or U12829 (N_12829,N_12571,N_12010);
or U12830 (N_12830,N_12094,N_12733);
or U12831 (N_12831,N_12131,N_12590);
and U12832 (N_12832,N_12390,N_12582);
nand U12833 (N_12833,N_12149,N_12156);
or U12834 (N_12834,N_12415,N_12623);
xnor U12835 (N_12835,N_12661,N_12643);
or U12836 (N_12836,N_12155,N_12009);
nand U12837 (N_12837,N_12561,N_12618);
and U12838 (N_12838,N_12472,N_12518);
or U12839 (N_12839,N_12172,N_12133);
nand U12840 (N_12840,N_12431,N_12050);
nand U12841 (N_12841,N_12509,N_12421);
xnor U12842 (N_12842,N_12488,N_12537);
nand U12843 (N_12843,N_12323,N_12007);
or U12844 (N_12844,N_12736,N_12256);
nor U12845 (N_12845,N_12525,N_12619);
xnor U12846 (N_12846,N_12591,N_12219);
and U12847 (N_12847,N_12233,N_12293);
and U12848 (N_12848,N_12225,N_12685);
and U12849 (N_12849,N_12083,N_12262);
xnor U12850 (N_12850,N_12679,N_12749);
and U12851 (N_12851,N_12215,N_12018);
nand U12852 (N_12852,N_12639,N_12037);
nor U12853 (N_12853,N_12170,N_12729);
nand U12854 (N_12854,N_12512,N_12550);
or U12855 (N_12855,N_12142,N_12070);
nand U12856 (N_12856,N_12515,N_12134);
nand U12857 (N_12857,N_12558,N_12650);
nor U12858 (N_12858,N_12135,N_12065);
and U12859 (N_12859,N_12355,N_12604);
xor U12860 (N_12860,N_12662,N_12583);
nand U12861 (N_12861,N_12592,N_12139);
or U12862 (N_12862,N_12252,N_12381);
and U12863 (N_12863,N_12530,N_12109);
nor U12864 (N_12864,N_12562,N_12064);
nand U12865 (N_12865,N_12013,N_12640);
xnor U12866 (N_12866,N_12271,N_12502);
or U12867 (N_12867,N_12716,N_12601);
and U12868 (N_12868,N_12630,N_12029);
or U12869 (N_12869,N_12709,N_12456);
and U12870 (N_12870,N_12161,N_12433);
nor U12871 (N_12871,N_12167,N_12406);
nor U12872 (N_12872,N_12347,N_12721);
and U12873 (N_12873,N_12085,N_12165);
or U12874 (N_12874,N_12373,N_12020);
nor U12875 (N_12875,N_12015,N_12594);
nor U12876 (N_12876,N_12659,N_12557);
xor U12877 (N_12877,N_12244,N_12336);
nand U12878 (N_12878,N_12128,N_12297);
and U12879 (N_12879,N_12722,N_12148);
or U12880 (N_12880,N_12264,N_12051);
xnor U12881 (N_12881,N_12248,N_12742);
and U12882 (N_12882,N_12053,N_12478);
and U12883 (N_12883,N_12338,N_12400);
or U12884 (N_12884,N_12718,N_12168);
or U12885 (N_12885,N_12039,N_12378);
and U12886 (N_12886,N_12675,N_12647);
and U12887 (N_12887,N_12125,N_12595);
nor U12888 (N_12888,N_12434,N_12348);
nor U12889 (N_12889,N_12163,N_12444);
nor U12890 (N_12890,N_12395,N_12209);
or U12891 (N_12891,N_12261,N_12385);
or U12892 (N_12892,N_12110,N_12730);
nand U12893 (N_12893,N_12036,N_12024);
nor U12894 (N_12894,N_12028,N_12388);
xor U12895 (N_12895,N_12120,N_12625);
or U12896 (N_12896,N_12396,N_12670);
or U12897 (N_12897,N_12426,N_12689);
or U12898 (N_12898,N_12331,N_12712);
or U12899 (N_12899,N_12251,N_12714);
or U12900 (N_12900,N_12180,N_12427);
or U12901 (N_12901,N_12211,N_12404);
xnor U12902 (N_12902,N_12291,N_12542);
nor U12903 (N_12903,N_12505,N_12187);
nor U12904 (N_12904,N_12578,N_12480);
nor U12905 (N_12905,N_12376,N_12000);
xnor U12906 (N_12906,N_12432,N_12504);
xor U12907 (N_12907,N_12651,N_12182);
xor U12908 (N_12908,N_12340,N_12270);
xor U12909 (N_12909,N_12317,N_12027);
nand U12910 (N_12910,N_12186,N_12313);
and U12911 (N_12911,N_12041,N_12710);
nor U12912 (N_12912,N_12354,N_12228);
and U12913 (N_12913,N_12366,N_12184);
xor U12914 (N_12914,N_12232,N_12398);
and U12915 (N_12915,N_12484,N_12409);
nand U12916 (N_12916,N_12278,N_12048);
nand U12917 (N_12917,N_12203,N_12044);
and U12918 (N_12918,N_12699,N_12470);
or U12919 (N_12919,N_12040,N_12519);
and U12920 (N_12920,N_12741,N_12077);
and U12921 (N_12921,N_12523,N_12141);
or U12922 (N_12922,N_12201,N_12458);
nand U12923 (N_12923,N_12605,N_12614);
nand U12924 (N_12924,N_12723,N_12580);
and U12925 (N_12925,N_12247,N_12243);
xnor U12926 (N_12926,N_12422,N_12491);
nor U12927 (N_12927,N_12719,N_12236);
nor U12928 (N_12928,N_12359,N_12389);
nor U12929 (N_12929,N_12538,N_12545);
nor U12930 (N_12930,N_12451,N_12683);
nor U12931 (N_12931,N_12738,N_12668);
xnor U12932 (N_12932,N_12315,N_12076);
xor U12933 (N_12933,N_12691,N_12008);
xnor U12934 (N_12934,N_12559,N_12033);
and U12935 (N_12935,N_12613,N_12239);
nor U12936 (N_12936,N_12412,N_12673);
or U12937 (N_12937,N_12055,N_12307);
and U12938 (N_12938,N_12362,N_12063);
xor U12939 (N_12939,N_12153,N_12632);
nand U12940 (N_12940,N_12279,N_12493);
nand U12941 (N_12941,N_12138,N_12298);
xnor U12942 (N_12942,N_12062,N_12486);
nand U12943 (N_12943,N_12318,N_12707);
and U12944 (N_12944,N_12637,N_12513);
and U12945 (N_12945,N_12332,N_12306);
and U12946 (N_12946,N_12617,N_12684);
xor U12947 (N_12947,N_12205,N_12497);
xor U12948 (N_12948,N_12501,N_12726);
nor U12949 (N_12949,N_12193,N_12467);
nor U12950 (N_12950,N_12520,N_12159);
nor U12951 (N_12951,N_12636,N_12032);
or U12952 (N_12952,N_12568,N_12521);
or U12953 (N_12953,N_12490,N_12197);
nand U12954 (N_12954,N_12672,N_12697);
nand U12955 (N_12955,N_12563,N_12417);
and U12956 (N_12956,N_12325,N_12634);
xor U12957 (N_12957,N_12553,N_12459);
xnor U12958 (N_12958,N_12287,N_12555);
xor U12959 (N_12959,N_12281,N_12495);
xor U12960 (N_12960,N_12296,N_12071);
nand U12961 (N_12961,N_12546,N_12638);
and U12962 (N_12962,N_12074,N_12119);
xnor U12963 (N_12963,N_12330,N_12349);
xnor U12964 (N_12964,N_12420,N_12677);
or U12965 (N_12965,N_12383,N_12616);
nor U12966 (N_12966,N_12727,N_12711);
nand U12967 (N_12967,N_12341,N_12510);
nand U12968 (N_12968,N_12054,N_12581);
xnor U12969 (N_12969,N_12081,N_12479);
nor U12970 (N_12970,N_12384,N_12506);
xnor U12971 (N_12971,N_12454,N_12289);
and U12972 (N_12972,N_12356,N_12646);
xnor U12973 (N_12973,N_12176,N_12088);
nor U12974 (N_12974,N_12025,N_12627);
nand U12975 (N_12975,N_12231,N_12477);
and U12976 (N_12976,N_12686,N_12273);
nand U12977 (N_12977,N_12123,N_12532);
and U12978 (N_12978,N_12014,N_12221);
nand U12979 (N_12979,N_12371,N_12034);
or U12980 (N_12980,N_12192,N_12351);
or U12981 (N_12981,N_12282,N_12295);
nand U12982 (N_12982,N_12556,N_12483);
xnor U12983 (N_12983,N_12648,N_12471);
nand U12984 (N_12984,N_12666,N_12482);
and U12985 (N_12985,N_12554,N_12259);
nor U12986 (N_12986,N_12419,N_12111);
xnor U12987 (N_12987,N_12631,N_12511);
nor U12988 (N_12988,N_12607,N_12460);
or U12989 (N_12989,N_12463,N_12284);
nor U12990 (N_12990,N_12466,N_12334);
nor U12991 (N_12991,N_12600,N_12042);
or U12992 (N_12992,N_12645,N_12641);
nor U12993 (N_12993,N_12529,N_12162);
and U12994 (N_12994,N_12112,N_12704);
and U12995 (N_12995,N_12304,N_12442);
and U12996 (N_12996,N_12342,N_12405);
xnor U12997 (N_12997,N_12255,N_12402);
nor U12998 (N_12998,N_12069,N_12528);
nand U12999 (N_12999,N_12329,N_12218);
or U13000 (N_13000,N_12327,N_12012);
nand U13001 (N_13001,N_12533,N_12204);
nor U13002 (N_13002,N_12263,N_12254);
or U13003 (N_13003,N_12058,N_12740);
nor U13004 (N_13004,N_12715,N_12573);
nand U13005 (N_13005,N_12057,N_12748);
and U13006 (N_13006,N_12301,N_12430);
or U13007 (N_13007,N_12541,N_12418);
or U13008 (N_13008,N_12060,N_12098);
nand U13009 (N_13009,N_12609,N_12335);
nor U13010 (N_13010,N_12003,N_12346);
nand U13011 (N_13011,N_12312,N_12343);
xor U13012 (N_13012,N_12593,N_12202);
nand U13013 (N_13013,N_12566,N_12494);
xnor U13014 (N_13014,N_12321,N_12171);
or U13015 (N_13015,N_12690,N_12199);
nor U13016 (N_13016,N_12725,N_12240);
xor U13017 (N_13017,N_12353,N_12450);
or U13018 (N_13018,N_12669,N_12569);
nor U13019 (N_13019,N_12309,N_12079);
nor U13020 (N_13020,N_12503,N_12588);
nand U13021 (N_13021,N_12567,N_12214);
nand U13022 (N_13022,N_12492,N_12526);
and U13023 (N_13023,N_12350,N_12365);
xnor U13024 (N_13024,N_12181,N_12196);
and U13025 (N_13025,N_12744,N_12461);
nand U13026 (N_13026,N_12002,N_12612);
or U13027 (N_13027,N_12728,N_12095);
xnor U13028 (N_13028,N_12696,N_12428);
and U13029 (N_13029,N_12628,N_12633);
xor U13030 (N_13030,N_12049,N_12308);
xor U13031 (N_13031,N_12746,N_12224);
nand U13032 (N_13032,N_12046,N_12021);
nor U13033 (N_13033,N_12499,N_12319);
xnor U13034 (N_13034,N_12100,N_12653);
and U13035 (N_13035,N_12455,N_12031);
xor U13036 (N_13036,N_12216,N_12399);
nand U13037 (N_13037,N_12485,N_12195);
and U13038 (N_13038,N_12552,N_12436);
or U13039 (N_13039,N_12598,N_12310);
or U13040 (N_13040,N_12257,N_12441);
nor U13041 (N_13041,N_12207,N_12075);
xnor U13042 (N_13042,N_12629,N_12223);
nor U13043 (N_13043,N_12487,N_12245);
nand U13044 (N_13044,N_12522,N_12656);
and U13045 (N_13045,N_12137,N_12272);
and U13046 (N_13046,N_12731,N_12175);
nand U13047 (N_13047,N_12603,N_12649);
nor U13048 (N_13048,N_12249,N_12671);
and U13049 (N_13049,N_12126,N_12173);
or U13050 (N_13050,N_12059,N_12572);
or U13051 (N_13051,N_12425,N_12144);
or U13052 (N_13052,N_12011,N_12424);
or U13053 (N_13053,N_12108,N_12026);
nor U13054 (N_13054,N_12320,N_12474);
nand U13055 (N_13055,N_12692,N_12129);
or U13056 (N_13056,N_12067,N_12105);
nor U13057 (N_13057,N_12302,N_12597);
nand U13058 (N_13058,N_12414,N_12030);
nor U13059 (N_13059,N_12401,N_12164);
xnor U13060 (N_13060,N_12136,N_12664);
xor U13061 (N_13061,N_12190,N_12179);
nor U13062 (N_13062,N_12508,N_12206);
and U13063 (N_13063,N_12547,N_12375);
nand U13064 (N_13064,N_12676,N_12560);
nand U13065 (N_13065,N_12056,N_12358);
or U13066 (N_13066,N_12534,N_12535);
or U13067 (N_13067,N_12739,N_12288);
xor U13068 (N_13068,N_12565,N_12576);
and U13069 (N_13069,N_12608,N_12724);
nand U13070 (N_13070,N_12411,N_12213);
nand U13071 (N_13071,N_12407,N_12352);
nand U13072 (N_13072,N_12453,N_12364);
xor U13073 (N_13073,N_12260,N_12570);
or U13074 (N_13074,N_12096,N_12160);
and U13075 (N_13075,N_12229,N_12621);
and U13076 (N_13076,N_12448,N_12090);
or U13077 (N_13077,N_12682,N_12117);
or U13078 (N_13078,N_12212,N_12102);
nand U13079 (N_13079,N_12708,N_12082);
xor U13080 (N_13080,N_12443,N_12413);
and U13081 (N_13081,N_12145,N_12394);
nor U13082 (N_13082,N_12099,N_12106);
and U13083 (N_13083,N_12344,N_12544);
or U13084 (N_13084,N_12393,N_12333);
nor U13085 (N_13085,N_12092,N_12674);
or U13086 (N_13086,N_12374,N_12300);
and U13087 (N_13087,N_12377,N_12121);
xnor U13088 (N_13088,N_12268,N_12140);
nand U13089 (N_13089,N_12178,N_12220);
or U13090 (N_13090,N_12585,N_12292);
nand U13091 (N_13091,N_12208,N_12498);
nor U13092 (N_13092,N_12693,N_12587);
nor U13093 (N_13093,N_12169,N_12695);
nor U13094 (N_13094,N_12698,N_12496);
and U13095 (N_13095,N_12087,N_12001);
nand U13096 (N_13096,N_12093,N_12387);
nand U13097 (N_13097,N_12328,N_12091);
nor U13098 (N_13098,N_12481,N_12665);
and U13099 (N_13099,N_12237,N_12113);
or U13100 (N_13100,N_12489,N_12115);
and U13101 (N_13101,N_12429,N_12266);
nand U13102 (N_13102,N_12652,N_12624);
nand U13103 (N_13103,N_12191,N_12655);
or U13104 (N_13104,N_12657,N_12735);
nand U13105 (N_13105,N_12370,N_12667);
nand U13106 (N_13106,N_12103,N_12403);
or U13107 (N_13107,N_12151,N_12435);
or U13108 (N_13108,N_12086,N_12097);
and U13109 (N_13109,N_12517,N_12275);
nor U13110 (N_13110,N_12610,N_12584);
or U13111 (N_13111,N_12705,N_12200);
nor U13112 (N_13112,N_12084,N_12250);
nand U13113 (N_13113,N_12283,N_12017);
nand U13114 (N_13114,N_12299,N_12241);
nor U13115 (N_13115,N_12700,N_12360);
nand U13116 (N_13116,N_12006,N_12464);
nor U13117 (N_13117,N_12680,N_12122);
and U13118 (N_13118,N_12152,N_12702);
nor U13119 (N_13119,N_12023,N_12468);
and U13120 (N_13120,N_12379,N_12066);
nor U13121 (N_13121,N_12469,N_12038);
or U13122 (N_13122,N_12615,N_12688);
nand U13123 (N_13123,N_12687,N_12357);
or U13124 (N_13124,N_12277,N_12107);
nor U13125 (N_13125,N_12375,N_12655);
or U13126 (N_13126,N_12062,N_12355);
and U13127 (N_13127,N_12284,N_12315);
and U13128 (N_13128,N_12710,N_12630);
and U13129 (N_13129,N_12111,N_12071);
xnor U13130 (N_13130,N_12459,N_12352);
and U13131 (N_13131,N_12493,N_12721);
xnor U13132 (N_13132,N_12109,N_12482);
xnor U13133 (N_13133,N_12455,N_12172);
xor U13134 (N_13134,N_12420,N_12475);
or U13135 (N_13135,N_12119,N_12235);
nand U13136 (N_13136,N_12122,N_12712);
nor U13137 (N_13137,N_12362,N_12148);
or U13138 (N_13138,N_12171,N_12305);
xnor U13139 (N_13139,N_12194,N_12091);
xor U13140 (N_13140,N_12171,N_12671);
nand U13141 (N_13141,N_12349,N_12208);
and U13142 (N_13142,N_12643,N_12032);
xor U13143 (N_13143,N_12313,N_12188);
xnor U13144 (N_13144,N_12076,N_12522);
nand U13145 (N_13145,N_12749,N_12216);
xor U13146 (N_13146,N_12676,N_12411);
nand U13147 (N_13147,N_12527,N_12176);
and U13148 (N_13148,N_12248,N_12512);
and U13149 (N_13149,N_12540,N_12431);
nand U13150 (N_13150,N_12612,N_12633);
xnor U13151 (N_13151,N_12675,N_12084);
xnor U13152 (N_13152,N_12693,N_12351);
and U13153 (N_13153,N_12725,N_12730);
nor U13154 (N_13154,N_12072,N_12615);
nor U13155 (N_13155,N_12162,N_12676);
and U13156 (N_13156,N_12367,N_12461);
and U13157 (N_13157,N_12128,N_12464);
nand U13158 (N_13158,N_12092,N_12101);
xnor U13159 (N_13159,N_12131,N_12636);
and U13160 (N_13160,N_12470,N_12351);
nor U13161 (N_13161,N_12272,N_12686);
and U13162 (N_13162,N_12565,N_12057);
nor U13163 (N_13163,N_12376,N_12345);
nand U13164 (N_13164,N_12285,N_12487);
nand U13165 (N_13165,N_12347,N_12027);
and U13166 (N_13166,N_12308,N_12167);
xnor U13167 (N_13167,N_12218,N_12275);
and U13168 (N_13168,N_12512,N_12272);
nor U13169 (N_13169,N_12605,N_12609);
and U13170 (N_13170,N_12107,N_12429);
xnor U13171 (N_13171,N_12376,N_12442);
nand U13172 (N_13172,N_12125,N_12417);
and U13173 (N_13173,N_12329,N_12529);
nor U13174 (N_13174,N_12043,N_12463);
xor U13175 (N_13175,N_12575,N_12340);
nor U13176 (N_13176,N_12223,N_12178);
or U13177 (N_13177,N_12342,N_12531);
nor U13178 (N_13178,N_12226,N_12284);
nand U13179 (N_13179,N_12250,N_12403);
and U13180 (N_13180,N_12618,N_12093);
nor U13181 (N_13181,N_12123,N_12132);
or U13182 (N_13182,N_12529,N_12451);
and U13183 (N_13183,N_12423,N_12404);
nand U13184 (N_13184,N_12728,N_12064);
xnor U13185 (N_13185,N_12524,N_12260);
and U13186 (N_13186,N_12420,N_12433);
xor U13187 (N_13187,N_12568,N_12489);
and U13188 (N_13188,N_12452,N_12145);
nor U13189 (N_13189,N_12538,N_12695);
xnor U13190 (N_13190,N_12455,N_12630);
nand U13191 (N_13191,N_12719,N_12134);
and U13192 (N_13192,N_12583,N_12017);
or U13193 (N_13193,N_12520,N_12237);
nor U13194 (N_13194,N_12264,N_12374);
and U13195 (N_13195,N_12212,N_12118);
xor U13196 (N_13196,N_12306,N_12014);
xnor U13197 (N_13197,N_12570,N_12012);
or U13198 (N_13198,N_12501,N_12495);
and U13199 (N_13199,N_12310,N_12007);
or U13200 (N_13200,N_12338,N_12335);
xor U13201 (N_13201,N_12096,N_12478);
and U13202 (N_13202,N_12259,N_12342);
or U13203 (N_13203,N_12586,N_12685);
and U13204 (N_13204,N_12141,N_12572);
or U13205 (N_13205,N_12536,N_12099);
nand U13206 (N_13206,N_12046,N_12280);
and U13207 (N_13207,N_12356,N_12554);
nand U13208 (N_13208,N_12139,N_12355);
nand U13209 (N_13209,N_12536,N_12152);
nor U13210 (N_13210,N_12257,N_12689);
and U13211 (N_13211,N_12260,N_12621);
and U13212 (N_13212,N_12063,N_12593);
nor U13213 (N_13213,N_12009,N_12655);
or U13214 (N_13214,N_12341,N_12409);
and U13215 (N_13215,N_12037,N_12453);
nor U13216 (N_13216,N_12470,N_12434);
or U13217 (N_13217,N_12047,N_12682);
nand U13218 (N_13218,N_12057,N_12008);
and U13219 (N_13219,N_12424,N_12357);
nand U13220 (N_13220,N_12673,N_12748);
or U13221 (N_13221,N_12124,N_12180);
and U13222 (N_13222,N_12062,N_12674);
and U13223 (N_13223,N_12260,N_12363);
xor U13224 (N_13224,N_12021,N_12038);
or U13225 (N_13225,N_12061,N_12741);
nand U13226 (N_13226,N_12233,N_12122);
or U13227 (N_13227,N_12586,N_12346);
and U13228 (N_13228,N_12587,N_12088);
and U13229 (N_13229,N_12607,N_12184);
or U13230 (N_13230,N_12434,N_12653);
xor U13231 (N_13231,N_12498,N_12161);
nand U13232 (N_13232,N_12224,N_12494);
nor U13233 (N_13233,N_12431,N_12105);
xor U13234 (N_13234,N_12597,N_12059);
or U13235 (N_13235,N_12619,N_12276);
or U13236 (N_13236,N_12018,N_12037);
nand U13237 (N_13237,N_12746,N_12586);
and U13238 (N_13238,N_12730,N_12049);
or U13239 (N_13239,N_12528,N_12248);
and U13240 (N_13240,N_12749,N_12285);
or U13241 (N_13241,N_12052,N_12032);
and U13242 (N_13242,N_12639,N_12077);
nor U13243 (N_13243,N_12511,N_12315);
nor U13244 (N_13244,N_12284,N_12338);
nor U13245 (N_13245,N_12254,N_12727);
nand U13246 (N_13246,N_12549,N_12459);
nand U13247 (N_13247,N_12263,N_12358);
nor U13248 (N_13248,N_12418,N_12182);
xnor U13249 (N_13249,N_12607,N_12407);
nand U13250 (N_13250,N_12190,N_12502);
xnor U13251 (N_13251,N_12738,N_12108);
or U13252 (N_13252,N_12364,N_12435);
nand U13253 (N_13253,N_12102,N_12220);
nor U13254 (N_13254,N_12690,N_12275);
or U13255 (N_13255,N_12600,N_12244);
xor U13256 (N_13256,N_12596,N_12270);
nor U13257 (N_13257,N_12698,N_12569);
xor U13258 (N_13258,N_12739,N_12318);
xor U13259 (N_13259,N_12572,N_12627);
nand U13260 (N_13260,N_12346,N_12100);
nor U13261 (N_13261,N_12414,N_12017);
nor U13262 (N_13262,N_12451,N_12195);
nor U13263 (N_13263,N_12648,N_12710);
xnor U13264 (N_13264,N_12008,N_12471);
xnor U13265 (N_13265,N_12038,N_12273);
xnor U13266 (N_13266,N_12096,N_12030);
or U13267 (N_13267,N_12171,N_12610);
nand U13268 (N_13268,N_12539,N_12008);
nor U13269 (N_13269,N_12671,N_12265);
xor U13270 (N_13270,N_12490,N_12495);
or U13271 (N_13271,N_12748,N_12575);
nor U13272 (N_13272,N_12324,N_12224);
nand U13273 (N_13273,N_12433,N_12305);
or U13274 (N_13274,N_12021,N_12659);
and U13275 (N_13275,N_12302,N_12350);
or U13276 (N_13276,N_12047,N_12247);
and U13277 (N_13277,N_12297,N_12284);
nand U13278 (N_13278,N_12249,N_12385);
nor U13279 (N_13279,N_12059,N_12517);
nor U13280 (N_13280,N_12103,N_12072);
xnor U13281 (N_13281,N_12169,N_12303);
and U13282 (N_13282,N_12326,N_12045);
nor U13283 (N_13283,N_12591,N_12212);
xnor U13284 (N_13284,N_12169,N_12563);
or U13285 (N_13285,N_12684,N_12254);
nand U13286 (N_13286,N_12654,N_12391);
nor U13287 (N_13287,N_12742,N_12173);
nor U13288 (N_13288,N_12586,N_12635);
xnor U13289 (N_13289,N_12285,N_12632);
nor U13290 (N_13290,N_12423,N_12616);
xor U13291 (N_13291,N_12236,N_12071);
nand U13292 (N_13292,N_12194,N_12642);
nor U13293 (N_13293,N_12450,N_12408);
nor U13294 (N_13294,N_12264,N_12353);
nor U13295 (N_13295,N_12158,N_12004);
or U13296 (N_13296,N_12640,N_12234);
or U13297 (N_13297,N_12375,N_12683);
nand U13298 (N_13298,N_12549,N_12146);
or U13299 (N_13299,N_12030,N_12061);
or U13300 (N_13300,N_12386,N_12232);
nand U13301 (N_13301,N_12212,N_12473);
and U13302 (N_13302,N_12713,N_12055);
nor U13303 (N_13303,N_12070,N_12430);
and U13304 (N_13304,N_12310,N_12113);
or U13305 (N_13305,N_12388,N_12651);
and U13306 (N_13306,N_12499,N_12218);
xnor U13307 (N_13307,N_12598,N_12148);
or U13308 (N_13308,N_12138,N_12445);
xor U13309 (N_13309,N_12566,N_12163);
and U13310 (N_13310,N_12468,N_12084);
nand U13311 (N_13311,N_12606,N_12339);
nor U13312 (N_13312,N_12661,N_12363);
nor U13313 (N_13313,N_12537,N_12423);
or U13314 (N_13314,N_12443,N_12650);
xnor U13315 (N_13315,N_12679,N_12635);
nor U13316 (N_13316,N_12492,N_12078);
nor U13317 (N_13317,N_12080,N_12514);
nand U13318 (N_13318,N_12095,N_12483);
nand U13319 (N_13319,N_12654,N_12578);
nand U13320 (N_13320,N_12476,N_12336);
xor U13321 (N_13321,N_12267,N_12067);
xnor U13322 (N_13322,N_12726,N_12116);
nand U13323 (N_13323,N_12079,N_12424);
nor U13324 (N_13324,N_12621,N_12327);
nand U13325 (N_13325,N_12430,N_12734);
and U13326 (N_13326,N_12047,N_12271);
or U13327 (N_13327,N_12714,N_12367);
and U13328 (N_13328,N_12645,N_12247);
xnor U13329 (N_13329,N_12290,N_12250);
and U13330 (N_13330,N_12004,N_12328);
nand U13331 (N_13331,N_12071,N_12273);
or U13332 (N_13332,N_12419,N_12334);
nand U13333 (N_13333,N_12285,N_12449);
nand U13334 (N_13334,N_12608,N_12384);
nand U13335 (N_13335,N_12113,N_12589);
nor U13336 (N_13336,N_12110,N_12205);
xor U13337 (N_13337,N_12567,N_12394);
and U13338 (N_13338,N_12022,N_12447);
and U13339 (N_13339,N_12661,N_12222);
or U13340 (N_13340,N_12400,N_12616);
or U13341 (N_13341,N_12678,N_12256);
nor U13342 (N_13342,N_12651,N_12285);
xnor U13343 (N_13343,N_12098,N_12123);
and U13344 (N_13344,N_12323,N_12114);
or U13345 (N_13345,N_12121,N_12340);
xor U13346 (N_13346,N_12358,N_12333);
or U13347 (N_13347,N_12226,N_12358);
or U13348 (N_13348,N_12518,N_12437);
or U13349 (N_13349,N_12723,N_12160);
xnor U13350 (N_13350,N_12429,N_12558);
nor U13351 (N_13351,N_12586,N_12532);
and U13352 (N_13352,N_12081,N_12568);
nand U13353 (N_13353,N_12561,N_12423);
nand U13354 (N_13354,N_12492,N_12031);
nor U13355 (N_13355,N_12736,N_12642);
or U13356 (N_13356,N_12719,N_12671);
and U13357 (N_13357,N_12603,N_12507);
and U13358 (N_13358,N_12125,N_12714);
nand U13359 (N_13359,N_12510,N_12084);
and U13360 (N_13360,N_12741,N_12528);
or U13361 (N_13361,N_12025,N_12214);
and U13362 (N_13362,N_12709,N_12480);
nor U13363 (N_13363,N_12300,N_12242);
or U13364 (N_13364,N_12593,N_12162);
and U13365 (N_13365,N_12331,N_12585);
nand U13366 (N_13366,N_12478,N_12744);
nand U13367 (N_13367,N_12346,N_12144);
or U13368 (N_13368,N_12319,N_12235);
and U13369 (N_13369,N_12001,N_12414);
or U13370 (N_13370,N_12652,N_12114);
xnor U13371 (N_13371,N_12121,N_12108);
xor U13372 (N_13372,N_12058,N_12506);
or U13373 (N_13373,N_12460,N_12054);
nand U13374 (N_13374,N_12494,N_12260);
xnor U13375 (N_13375,N_12626,N_12552);
nor U13376 (N_13376,N_12352,N_12440);
nor U13377 (N_13377,N_12193,N_12470);
and U13378 (N_13378,N_12682,N_12377);
nand U13379 (N_13379,N_12480,N_12251);
xor U13380 (N_13380,N_12462,N_12502);
or U13381 (N_13381,N_12075,N_12714);
nor U13382 (N_13382,N_12129,N_12550);
nor U13383 (N_13383,N_12082,N_12620);
nand U13384 (N_13384,N_12172,N_12106);
or U13385 (N_13385,N_12189,N_12044);
or U13386 (N_13386,N_12152,N_12061);
and U13387 (N_13387,N_12533,N_12325);
xor U13388 (N_13388,N_12271,N_12108);
and U13389 (N_13389,N_12449,N_12332);
nand U13390 (N_13390,N_12574,N_12456);
nand U13391 (N_13391,N_12282,N_12058);
xor U13392 (N_13392,N_12588,N_12744);
nor U13393 (N_13393,N_12504,N_12206);
xor U13394 (N_13394,N_12690,N_12589);
nor U13395 (N_13395,N_12671,N_12605);
xor U13396 (N_13396,N_12037,N_12486);
nor U13397 (N_13397,N_12733,N_12087);
or U13398 (N_13398,N_12235,N_12746);
and U13399 (N_13399,N_12318,N_12136);
or U13400 (N_13400,N_12382,N_12088);
or U13401 (N_13401,N_12455,N_12440);
and U13402 (N_13402,N_12400,N_12183);
nand U13403 (N_13403,N_12463,N_12099);
nor U13404 (N_13404,N_12324,N_12027);
and U13405 (N_13405,N_12336,N_12367);
or U13406 (N_13406,N_12163,N_12054);
or U13407 (N_13407,N_12569,N_12641);
xor U13408 (N_13408,N_12441,N_12442);
xor U13409 (N_13409,N_12179,N_12531);
and U13410 (N_13410,N_12074,N_12356);
xor U13411 (N_13411,N_12045,N_12673);
nand U13412 (N_13412,N_12412,N_12055);
nand U13413 (N_13413,N_12375,N_12304);
or U13414 (N_13414,N_12105,N_12294);
nand U13415 (N_13415,N_12061,N_12056);
or U13416 (N_13416,N_12281,N_12355);
or U13417 (N_13417,N_12151,N_12621);
xnor U13418 (N_13418,N_12243,N_12300);
xnor U13419 (N_13419,N_12200,N_12396);
nor U13420 (N_13420,N_12222,N_12474);
nor U13421 (N_13421,N_12227,N_12639);
nand U13422 (N_13422,N_12135,N_12591);
nor U13423 (N_13423,N_12146,N_12534);
or U13424 (N_13424,N_12185,N_12384);
xnor U13425 (N_13425,N_12118,N_12395);
and U13426 (N_13426,N_12019,N_12633);
and U13427 (N_13427,N_12554,N_12272);
and U13428 (N_13428,N_12745,N_12482);
or U13429 (N_13429,N_12550,N_12460);
and U13430 (N_13430,N_12189,N_12743);
and U13431 (N_13431,N_12705,N_12075);
nand U13432 (N_13432,N_12718,N_12199);
nand U13433 (N_13433,N_12019,N_12374);
and U13434 (N_13434,N_12440,N_12194);
xor U13435 (N_13435,N_12319,N_12244);
nand U13436 (N_13436,N_12745,N_12346);
nand U13437 (N_13437,N_12465,N_12476);
or U13438 (N_13438,N_12094,N_12442);
nor U13439 (N_13439,N_12032,N_12498);
nand U13440 (N_13440,N_12601,N_12297);
and U13441 (N_13441,N_12311,N_12082);
nand U13442 (N_13442,N_12088,N_12704);
and U13443 (N_13443,N_12739,N_12623);
or U13444 (N_13444,N_12744,N_12233);
xor U13445 (N_13445,N_12409,N_12179);
or U13446 (N_13446,N_12267,N_12708);
and U13447 (N_13447,N_12619,N_12572);
and U13448 (N_13448,N_12695,N_12458);
or U13449 (N_13449,N_12708,N_12099);
nand U13450 (N_13450,N_12365,N_12065);
nor U13451 (N_13451,N_12694,N_12544);
nand U13452 (N_13452,N_12368,N_12469);
nand U13453 (N_13453,N_12177,N_12008);
nand U13454 (N_13454,N_12708,N_12076);
nor U13455 (N_13455,N_12142,N_12301);
or U13456 (N_13456,N_12724,N_12403);
xor U13457 (N_13457,N_12584,N_12244);
and U13458 (N_13458,N_12530,N_12141);
or U13459 (N_13459,N_12556,N_12601);
xor U13460 (N_13460,N_12344,N_12278);
xnor U13461 (N_13461,N_12749,N_12474);
xor U13462 (N_13462,N_12450,N_12414);
and U13463 (N_13463,N_12744,N_12679);
nand U13464 (N_13464,N_12530,N_12517);
and U13465 (N_13465,N_12639,N_12184);
nand U13466 (N_13466,N_12143,N_12657);
and U13467 (N_13467,N_12576,N_12179);
or U13468 (N_13468,N_12498,N_12433);
xnor U13469 (N_13469,N_12013,N_12617);
and U13470 (N_13470,N_12695,N_12065);
xor U13471 (N_13471,N_12273,N_12666);
nor U13472 (N_13472,N_12131,N_12606);
nor U13473 (N_13473,N_12587,N_12525);
and U13474 (N_13474,N_12062,N_12207);
nand U13475 (N_13475,N_12328,N_12446);
nand U13476 (N_13476,N_12527,N_12146);
nor U13477 (N_13477,N_12238,N_12171);
or U13478 (N_13478,N_12627,N_12106);
and U13479 (N_13479,N_12141,N_12086);
xnor U13480 (N_13480,N_12108,N_12387);
and U13481 (N_13481,N_12335,N_12127);
nor U13482 (N_13482,N_12352,N_12437);
nand U13483 (N_13483,N_12044,N_12649);
or U13484 (N_13484,N_12041,N_12194);
nor U13485 (N_13485,N_12568,N_12189);
nand U13486 (N_13486,N_12492,N_12403);
nand U13487 (N_13487,N_12543,N_12580);
nor U13488 (N_13488,N_12253,N_12025);
nor U13489 (N_13489,N_12132,N_12090);
and U13490 (N_13490,N_12448,N_12349);
nand U13491 (N_13491,N_12453,N_12178);
and U13492 (N_13492,N_12536,N_12702);
or U13493 (N_13493,N_12404,N_12446);
or U13494 (N_13494,N_12225,N_12119);
nand U13495 (N_13495,N_12576,N_12585);
xnor U13496 (N_13496,N_12420,N_12370);
and U13497 (N_13497,N_12493,N_12028);
xor U13498 (N_13498,N_12628,N_12748);
nand U13499 (N_13499,N_12231,N_12748);
or U13500 (N_13500,N_12779,N_13250);
or U13501 (N_13501,N_12817,N_13065);
xor U13502 (N_13502,N_13432,N_12933);
xor U13503 (N_13503,N_13187,N_12774);
and U13504 (N_13504,N_13229,N_12828);
nor U13505 (N_13505,N_13411,N_13087);
nor U13506 (N_13506,N_12784,N_12822);
or U13507 (N_13507,N_12985,N_13167);
nand U13508 (N_13508,N_13104,N_13365);
or U13509 (N_13509,N_12994,N_13484);
nor U13510 (N_13510,N_13429,N_12962);
xnor U13511 (N_13511,N_13311,N_12764);
nor U13512 (N_13512,N_12860,N_12954);
or U13513 (N_13513,N_13348,N_13122);
or U13514 (N_13514,N_13426,N_12757);
xor U13515 (N_13515,N_13218,N_13401);
or U13516 (N_13516,N_12857,N_12937);
nor U13517 (N_13517,N_13391,N_12815);
and U13518 (N_13518,N_12751,N_13333);
and U13519 (N_13519,N_13388,N_12928);
nand U13520 (N_13520,N_13350,N_13019);
or U13521 (N_13521,N_13143,N_13375);
nand U13522 (N_13522,N_13406,N_12889);
nor U13523 (N_13523,N_12943,N_13112);
nor U13524 (N_13524,N_13277,N_12785);
and U13525 (N_13525,N_13370,N_12795);
and U13526 (N_13526,N_13231,N_13307);
nand U13527 (N_13527,N_12931,N_13466);
nor U13528 (N_13528,N_12995,N_13496);
or U13529 (N_13529,N_13319,N_13085);
nand U13530 (N_13530,N_12959,N_13376);
and U13531 (N_13531,N_13062,N_13114);
and U13532 (N_13532,N_12821,N_13073);
or U13533 (N_13533,N_13165,N_13237);
and U13534 (N_13534,N_12909,N_12776);
nand U13535 (N_13535,N_12819,N_13436);
and U13536 (N_13536,N_13223,N_12914);
and U13537 (N_13537,N_12976,N_13485);
nand U13538 (N_13538,N_13280,N_12899);
nand U13539 (N_13539,N_13068,N_13448);
xnor U13540 (N_13540,N_12855,N_12811);
nand U13541 (N_13541,N_13259,N_13089);
and U13542 (N_13542,N_13139,N_13385);
nor U13543 (N_13543,N_13027,N_13442);
nand U13544 (N_13544,N_13458,N_13208);
or U13545 (N_13545,N_13434,N_13278);
or U13546 (N_13546,N_13053,N_13393);
nand U13547 (N_13547,N_13449,N_12788);
and U13548 (N_13548,N_13238,N_13312);
and U13549 (N_13549,N_13140,N_13047);
nor U13550 (N_13550,N_13362,N_12812);
and U13551 (N_13551,N_13135,N_13182);
nor U13552 (N_13552,N_12966,N_12881);
and U13553 (N_13553,N_13324,N_13467);
and U13554 (N_13554,N_13265,N_13121);
nand U13555 (N_13555,N_13258,N_13013);
nor U13556 (N_13556,N_13389,N_13244);
or U13557 (N_13557,N_13402,N_13322);
nand U13558 (N_13558,N_12946,N_13042);
or U13559 (N_13559,N_12756,N_13300);
xor U13560 (N_13560,N_12871,N_13005);
nor U13561 (N_13561,N_12830,N_12953);
or U13562 (N_13562,N_13180,N_13001);
xor U13563 (N_13563,N_12856,N_13146);
and U13564 (N_13564,N_13220,N_13248);
and U13565 (N_13565,N_12964,N_12957);
nor U13566 (N_13566,N_12772,N_12965);
and U13567 (N_13567,N_13025,N_12932);
nand U13568 (N_13568,N_12865,N_12872);
xor U13569 (N_13569,N_13334,N_12910);
or U13570 (N_13570,N_13346,N_13067);
nor U13571 (N_13571,N_12798,N_13310);
nor U13572 (N_13572,N_12980,N_13308);
nand U13573 (N_13573,N_12921,N_13166);
nand U13574 (N_13574,N_13291,N_12903);
xor U13575 (N_13575,N_13292,N_12926);
xor U13576 (N_13576,N_13041,N_13373);
or U13577 (N_13577,N_12977,N_12864);
nor U13578 (N_13578,N_13188,N_13261);
nor U13579 (N_13579,N_13183,N_12752);
and U13580 (N_13580,N_13021,N_12758);
xnor U13581 (N_13581,N_13460,N_13301);
nand U13582 (N_13582,N_13046,N_12929);
or U13583 (N_13583,N_13342,N_13274);
xnor U13584 (N_13584,N_13245,N_13396);
nor U13585 (N_13585,N_13490,N_13051);
and U13586 (N_13586,N_13256,N_12908);
xnor U13587 (N_13587,N_13164,N_13195);
nand U13588 (N_13588,N_12942,N_12882);
nand U13589 (N_13589,N_13133,N_13029);
xnor U13590 (N_13590,N_12922,N_13058);
xnor U13591 (N_13591,N_13205,N_12952);
nor U13592 (N_13592,N_12923,N_12898);
xor U13593 (N_13593,N_12963,N_12790);
and U13594 (N_13594,N_12939,N_13414);
nor U13595 (N_13595,N_12997,N_13254);
xor U13596 (N_13596,N_12941,N_13197);
and U13597 (N_13597,N_13323,N_12802);
or U13598 (N_13598,N_13387,N_12984);
nand U13599 (N_13599,N_12917,N_12777);
and U13600 (N_13600,N_13384,N_13214);
or U13601 (N_13601,N_13476,N_12971);
and U13602 (N_13602,N_13149,N_13359);
nand U13603 (N_13603,N_13050,N_13453);
or U13604 (N_13604,N_12835,N_12780);
nand U13605 (N_13605,N_12991,N_13398);
or U13606 (N_13606,N_12750,N_12841);
or U13607 (N_13607,N_13433,N_12905);
or U13608 (N_13608,N_12759,N_12753);
and U13609 (N_13609,N_12891,N_13262);
xnor U13610 (N_13610,N_13289,N_12924);
xnor U13611 (N_13611,N_12775,N_12869);
and U13612 (N_13612,N_13239,N_13386);
or U13613 (N_13613,N_13036,N_13459);
nand U13614 (N_13614,N_12988,N_13209);
nor U13615 (N_13615,N_13427,N_13022);
nand U13616 (N_13616,N_13253,N_13006);
nor U13617 (N_13617,N_12766,N_12816);
nand U13618 (N_13618,N_13355,N_13227);
nand U13619 (N_13619,N_13107,N_13321);
nand U13620 (N_13620,N_13132,N_13158);
nand U13621 (N_13621,N_12993,N_13482);
or U13622 (N_13622,N_12810,N_13263);
or U13623 (N_13623,N_12918,N_13086);
nand U13624 (N_13624,N_13399,N_12862);
xnor U13625 (N_13625,N_13251,N_12916);
nor U13626 (N_13626,N_13286,N_13240);
nor U13627 (N_13627,N_13198,N_13040);
nand U13628 (N_13628,N_12875,N_12883);
nor U13629 (N_13629,N_13488,N_13230);
xnor U13630 (N_13630,N_13381,N_13232);
and U13631 (N_13631,N_13106,N_12934);
or U13632 (N_13632,N_13163,N_12996);
nand U13633 (N_13633,N_13331,N_12840);
xnor U13634 (N_13634,N_13222,N_13079);
xnor U13635 (N_13635,N_13294,N_13002);
xor U13636 (N_13636,N_12806,N_12796);
nand U13637 (N_13637,N_13302,N_12803);
xor U13638 (N_13638,N_13445,N_12868);
and U13639 (N_13639,N_12832,N_13236);
nor U13640 (N_13640,N_13093,N_13160);
nand U13641 (N_13641,N_12853,N_12833);
xor U13642 (N_13642,N_13416,N_12854);
or U13643 (N_13643,N_13423,N_12925);
and U13644 (N_13644,N_12808,N_12878);
xnor U13645 (N_13645,N_13216,N_13055);
nand U13646 (N_13646,N_13012,N_13113);
xor U13647 (N_13647,N_12814,N_13407);
and U13648 (N_13648,N_13337,N_13366);
or U13649 (N_13649,N_12986,N_13039);
or U13650 (N_13650,N_13336,N_13465);
and U13651 (N_13651,N_13455,N_13276);
xnor U13652 (N_13652,N_13137,N_12896);
nor U13653 (N_13653,N_13059,N_13363);
nor U13654 (N_13654,N_13155,N_13226);
nand U13655 (N_13655,N_13437,N_13264);
or U13656 (N_13656,N_13344,N_13268);
and U13657 (N_13657,N_12754,N_12846);
xnor U13658 (N_13658,N_13456,N_13494);
or U13659 (N_13659,N_13123,N_12907);
or U13660 (N_13660,N_12786,N_13234);
and U13661 (N_13661,N_12763,N_12804);
or U13662 (N_13662,N_12900,N_13428);
nand U13663 (N_13663,N_12992,N_13493);
nor U13664 (N_13664,N_13127,N_12970);
and U13665 (N_13665,N_13179,N_12894);
or U13666 (N_13666,N_13446,N_13097);
xor U13667 (N_13667,N_13316,N_13405);
or U13668 (N_13668,N_13215,N_12904);
or U13669 (N_13669,N_12800,N_13266);
and U13670 (N_13670,N_13211,N_13242);
nor U13671 (N_13671,N_13260,N_13017);
nand U13672 (N_13672,N_13033,N_13201);
nor U13673 (N_13673,N_13147,N_12998);
or U13674 (N_13674,N_12760,N_13142);
nor U13675 (N_13675,N_13473,N_13210);
nand U13676 (N_13676,N_13094,N_13221);
or U13677 (N_13677,N_12902,N_12972);
nand U13678 (N_13678,N_12771,N_12887);
and U13679 (N_13679,N_12919,N_13084);
or U13680 (N_13680,N_12895,N_13247);
and U13681 (N_13681,N_13326,N_13091);
nand U13682 (N_13682,N_12765,N_12809);
nor U13683 (N_13683,N_13119,N_13361);
nand U13684 (N_13684,N_13270,N_12967);
xnor U13685 (N_13685,N_13194,N_13438);
nor U13686 (N_13686,N_12866,N_13054);
or U13687 (N_13687,N_13471,N_13475);
nand U13688 (N_13688,N_12911,N_13109);
nand U13689 (N_13689,N_12936,N_13374);
or U13690 (N_13690,N_12982,N_13469);
xnor U13691 (N_13691,N_13076,N_13349);
xnor U13692 (N_13692,N_13477,N_12886);
nor U13693 (N_13693,N_12888,N_12787);
nand U13694 (N_13694,N_12901,N_13128);
nor U13695 (N_13695,N_13024,N_13000);
nor U13696 (N_13696,N_13172,N_12935);
and U13697 (N_13697,N_13287,N_13313);
xor U13698 (N_13698,N_13367,N_13358);
nor U13699 (N_13699,N_13305,N_13273);
and U13700 (N_13700,N_13202,N_13169);
nand U13701 (N_13701,N_13392,N_12949);
nor U13702 (N_13702,N_13173,N_13070);
nand U13703 (N_13703,N_12892,N_13424);
xnor U13704 (N_13704,N_12973,N_12990);
xnor U13705 (N_13705,N_12893,N_12768);
nand U13706 (N_13706,N_13196,N_13463);
or U13707 (N_13707,N_13329,N_13083);
xor U13708 (N_13708,N_13332,N_13299);
nand U13709 (N_13709,N_13110,N_12851);
xor U13710 (N_13710,N_12770,N_13031);
xor U13711 (N_13711,N_12940,N_12791);
nand U13712 (N_13712,N_12838,N_12829);
and U13713 (N_13713,N_13372,N_13452);
and U13714 (N_13714,N_12844,N_13281);
xnor U13715 (N_13715,N_13327,N_13498);
nand U13716 (N_13716,N_13175,N_12979);
nor U13717 (N_13717,N_12879,N_13212);
xnor U13718 (N_13718,N_13383,N_13082);
xnor U13719 (N_13719,N_12792,N_12825);
or U13720 (N_13720,N_13296,N_13295);
or U13721 (N_13721,N_13454,N_12861);
or U13722 (N_13722,N_13315,N_12850);
or U13723 (N_13723,N_12870,N_13081);
and U13724 (N_13724,N_12987,N_13092);
xnor U13725 (N_13725,N_12824,N_12805);
nor U13726 (N_13726,N_13074,N_13144);
or U13727 (N_13727,N_13377,N_13397);
nor U13728 (N_13728,N_13224,N_12843);
xor U13729 (N_13729,N_13447,N_13161);
xor U13730 (N_13730,N_13404,N_13102);
xor U13731 (N_13731,N_12955,N_12890);
nor U13732 (N_13732,N_12769,N_13048);
and U13733 (N_13733,N_12961,N_12818);
or U13734 (N_13734,N_12852,N_12797);
xor U13735 (N_13735,N_12960,N_12793);
and U13736 (N_13736,N_13479,N_12983);
and U13737 (N_13737,N_13297,N_13152);
xor U13738 (N_13738,N_13283,N_12858);
and U13739 (N_13739,N_13497,N_13072);
nor U13740 (N_13740,N_13007,N_13368);
and U13741 (N_13741,N_12826,N_13421);
or U13742 (N_13742,N_13200,N_13468);
xor U13743 (N_13743,N_13157,N_13257);
and U13744 (N_13744,N_13118,N_12767);
and U13745 (N_13745,N_13255,N_13035);
or U13746 (N_13746,N_13117,N_12874);
xnor U13747 (N_13747,N_12873,N_13444);
xnor U13748 (N_13748,N_13353,N_13489);
nand U13749 (N_13749,N_12956,N_12950);
nor U13750 (N_13750,N_13400,N_12978);
and U13751 (N_13751,N_13462,N_12969);
nand U13752 (N_13752,N_13271,N_13450);
xor U13753 (N_13753,N_12755,N_12876);
or U13754 (N_13754,N_13116,N_12778);
xnor U13755 (N_13755,N_13413,N_13009);
nand U13756 (N_13756,N_12948,N_13395);
and U13757 (N_13757,N_13306,N_13330);
xor U13758 (N_13758,N_13233,N_13063);
and U13759 (N_13759,N_13343,N_13145);
and U13760 (N_13760,N_13481,N_13379);
or U13761 (N_13761,N_13192,N_13335);
nand U13762 (N_13762,N_13243,N_13235);
and U13763 (N_13763,N_12842,N_13320);
and U13764 (N_13764,N_13408,N_13185);
or U13765 (N_13765,N_13241,N_12944);
nor U13766 (N_13766,N_13246,N_13478);
nor U13767 (N_13767,N_13080,N_13115);
nor U13768 (N_13768,N_13181,N_12807);
nand U13769 (N_13769,N_13045,N_13440);
nor U13770 (N_13770,N_13105,N_13282);
xor U13771 (N_13771,N_12999,N_13325);
nand U13772 (N_13772,N_13154,N_12863);
xnor U13773 (N_13773,N_13430,N_13483);
and U13774 (N_13774,N_13038,N_12968);
or U13775 (N_13775,N_13288,N_13345);
nand U13776 (N_13776,N_12927,N_12915);
nand U13777 (N_13777,N_13425,N_13225);
or U13778 (N_13778,N_12813,N_13049);
xor U13779 (N_13779,N_13124,N_12782);
xor U13780 (N_13780,N_13153,N_13360);
xor U13781 (N_13781,N_13011,N_12794);
or U13782 (N_13782,N_12789,N_13150);
nor U13783 (N_13783,N_12958,N_13004);
nand U13784 (N_13784,N_13390,N_12930);
and U13785 (N_13785,N_13409,N_13159);
nand U13786 (N_13786,N_13491,N_13298);
xnor U13787 (N_13787,N_13023,N_12989);
nand U13788 (N_13788,N_12847,N_13010);
or U13789 (N_13789,N_13472,N_13364);
and U13790 (N_13790,N_12761,N_13394);
xor U13791 (N_13791,N_13439,N_13304);
and U13792 (N_13792,N_13131,N_13317);
xnor U13793 (N_13793,N_13136,N_13129);
and U13794 (N_13794,N_12837,N_13219);
and U13795 (N_13795,N_13037,N_13470);
xnor U13796 (N_13796,N_13486,N_13269);
nand U13797 (N_13797,N_13203,N_13206);
and U13798 (N_13798,N_13191,N_13030);
and U13799 (N_13799,N_13412,N_13156);
and U13800 (N_13800,N_13026,N_13020);
xnor U13801 (N_13801,N_13267,N_13126);
nand U13802 (N_13802,N_13352,N_13151);
nand U13803 (N_13803,N_12897,N_13184);
or U13804 (N_13804,N_13347,N_13016);
nand U13805 (N_13805,N_13495,N_13303);
xor U13806 (N_13806,N_13043,N_13314);
and U13807 (N_13807,N_13419,N_13060);
or U13808 (N_13808,N_12827,N_13189);
nor U13809 (N_13809,N_13103,N_13417);
and U13810 (N_13810,N_12884,N_13285);
nor U13811 (N_13811,N_13293,N_12762);
xnor U13812 (N_13812,N_13499,N_13141);
or U13813 (N_13813,N_12848,N_12947);
nor U13814 (N_13814,N_13382,N_12913);
or U13815 (N_13815,N_13461,N_13171);
nor U13816 (N_13816,N_13369,N_13170);
or U13817 (N_13817,N_13357,N_13275);
xnor U13818 (N_13818,N_13108,N_13410);
or U13819 (N_13819,N_13088,N_13052);
or U13820 (N_13820,N_12938,N_13014);
nand U13821 (N_13821,N_13101,N_13371);
nand U13822 (N_13822,N_12783,N_13069);
or U13823 (N_13823,N_12880,N_13061);
or U13824 (N_13824,N_12845,N_13190);
xnor U13825 (N_13825,N_12823,N_13028);
nand U13826 (N_13826,N_13431,N_12975);
and U13827 (N_13827,N_12820,N_13207);
nand U13828 (N_13828,N_13178,N_13217);
nand U13829 (N_13829,N_12981,N_13015);
xor U13830 (N_13830,N_13176,N_13044);
nand U13831 (N_13831,N_13125,N_12834);
and U13832 (N_13832,N_12867,N_13090);
nand U13833 (N_13833,N_13457,N_13018);
nand U13834 (N_13834,N_12885,N_13378);
nor U13835 (N_13835,N_13099,N_12951);
xnor U13836 (N_13836,N_13443,N_13422);
nor U13837 (N_13837,N_13077,N_13279);
xnor U13838 (N_13838,N_13193,N_13354);
and U13839 (N_13839,N_13100,N_13204);
nand U13840 (N_13840,N_13351,N_13403);
or U13841 (N_13841,N_13098,N_13148);
and U13842 (N_13842,N_13056,N_13492);
xor U13843 (N_13843,N_13464,N_12801);
nand U13844 (N_13844,N_12906,N_12836);
xor U13845 (N_13845,N_13420,N_13078);
xor U13846 (N_13846,N_13034,N_13415);
nand U13847 (N_13847,N_13451,N_13138);
xnor U13848 (N_13848,N_13380,N_12839);
or U13849 (N_13849,N_13309,N_12877);
xnor U13850 (N_13850,N_13066,N_13213);
xor U13851 (N_13851,N_12945,N_13356);
nand U13852 (N_13852,N_13418,N_13487);
or U13853 (N_13853,N_12781,N_12974);
nor U13854 (N_13854,N_13474,N_13057);
or U13855 (N_13855,N_13328,N_12859);
or U13856 (N_13856,N_13177,N_13272);
or U13857 (N_13857,N_13318,N_13096);
xnor U13858 (N_13858,N_13120,N_12912);
nand U13859 (N_13859,N_13008,N_13111);
nor U13860 (N_13860,N_13168,N_13071);
nor U13861 (N_13861,N_13095,N_12831);
xnor U13862 (N_13862,N_13064,N_13480);
nor U13863 (N_13863,N_13340,N_13032);
nor U13864 (N_13864,N_13338,N_13003);
xor U13865 (N_13865,N_13199,N_13130);
nor U13866 (N_13866,N_13290,N_13252);
or U13867 (N_13867,N_13186,N_12849);
xnor U13868 (N_13868,N_13441,N_13435);
xnor U13869 (N_13869,N_13284,N_12920);
xnor U13870 (N_13870,N_13249,N_13162);
and U13871 (N_13871,N_13075,N_13134);
nor U13872 (N_13872,N_13228,N_13174);
and U13873 (N_13873,N_13339,N_12773);
and U13874 (N_13874,N_12799,N_13341);
nor U13875 (N_13875,N_13357,N_12893);
nand U13876 (N_13876,N_12952,N_13187);
or U13877 (N_13877,N_13274,N_12944);
nor U13878 (N_13878,N_13029,N_13249);
nor U13879 (N_13879,N_13152,N_12843);
nor U13880 (N_13880,N_12889,N_13382);
or U13881 (N_13881,N_13152,N_13322);
nor U13882 (N_13882,N_13397,N_12786);
nor U13883 (N_13883,N_13397,N_13155);
nand U13884 (N_13884,N_13303,N_13301);
nand U13885 (N_13885,N_13004,N_12898);
and U13886 (N_13886,N_12823,N_12955);
and U13887 (N_13887,N_13383,N_12936);
nor U13888 (N_13888,N_13121,N_13115);
xor U13889 (N_13889,N_13040,N_13338);
and U13890 (N_13890,N_13124,N_13027);
and U13891 (N_13891,N_12939,N_13272);
xnor U13892 (N_13892,N_12841,N_13457);
nor U13893 (N_13893,N_13354,N_13189);
xnor U13894 (N_13894,N_13144,N_12900);
or U13895 (N_13895,N_13328,N_12811);
xnor U13896 (N_13896,N_13245,N_13393);
nor U13897 (N_13897,N_13080,N_13122);
nor U13898 (N_13898,N_13132,N_12899);
or U13899 (N_13899,N_13014,N_13488);
nand U13900 (N_13900,N_13107,N_13080);
xor U13901 (N_13901,N_13061,N_13476);
and U13902 (N_13902,N_13164,N_13336);
xnor U13903 (N_13903,N_13141,N_13008);
nand U13904 (N_13904,N_12799,N_13157);
and U13905 (N_13905,N_13264,N_13422);
and U13906 (N_13906,N_12909,N_13398);
nand U13907 (N_13907,N_13075,N_13117);
or U13908 (N_13908,N_13069,N_12828);
or U13909 (N_13909,N_12792,N_13369);
nor U13910 (N_13910,N_13105,N_12869);
and U13911 (N_13911,N_13051,N_12855);
nand U13912 (N_13912,N_12903,N_12984);
nand U13913 (N_13913,N_12862,N_13128);
nand U13914 (N_13914,N_12976,N_13272);
xor U13915 (N_13915,N_13088,N_12941);
or U13916 (N_13916,N_13467,N_13391);
and U13917 (N_13917,N_13325,N_13473);
nor U13918 (N_13918,N_12899,N_13340);
nand U13919 (N_13919,N_13337,N_13245);
or U13920 (N_13920,N_13324,N_13048);
or U13921 (N_13921,N_13173,N_12866);
nand U13922 (N_13922,N_13426,N_13299);
or U13923 (N_13923,N_13188,N_13441);
xor U13924 (N_13924,N_12969,N_12846);
or U13925 (N_13925,N_12758,N_12863);
and U13926 (N_13926,N_13342,N_13108);
nand U13927 (N_13927,N_13139,N_12899);
and U13928 (N_13928,N_13356,N_12901);
or U13929 (N_13929,N_12937,N_13462);
and U13930 (N_13930,N_12922,N_13350);
and U13931 (N_13931,N_12798,N_13164);
nor U13932 (N_13932,N_13244,N_13413);
nand U13933 (N_13933,N_12817,N_13329);
nor U13934 (N_13934,N_13426,N_13498);
xor U13935 (N_13935,N_13054,N_13471);
and U13936 (N_13936,N_12802,N_13310);
and U13937 (N_13937,N_13078,N_13019);
and U13938 (N_13938,N_13409,N_13396);
xnor U13939 (N_13939,N_13473,N_12839);
and U13940 (N_13940,N_13149,N_13018);
nand U13941 (N_13941,N_13293,N_13183);
nor U13942 (N_13942,N_13294,N_12869);
and U13943 (N_13943,N_13245,N_13304);
nand U13944 (N_13944,N_12847,N_12750);
and U13945 (N_13945,N_12813,N_12904);
xnor U13946 (N_13946,N_13466,N_13237);
nand U13947 (N_13947,N_13213,N_12968);
nor U13948 (N_13948,N_13271,N_13128);
and U13949 (N_13949,N_13079,N_13011);
and U13950 (N_13950,N_13072,N_12810);
xnor U13951 (N_13951,N_13107,N_13006);
nor U13952 (N_13952,N_12817,N_13176);
nor U13953 (N_13953,N_13121,N_13213);
nor U13954 (N_13954,N_13177,N_13452);
and U13955 (N_13955,N_13312,N_13176);
xor U13956 (N_13956,N_13315,N_13298);
nand U13957 (N_13957,N_13265,N_13043);
nand U13958 (N_13958,N_13424,N_13475);
and U13959 (N_13959,N_13173,N_12844);
nor U13960 (N_13960,N_13159,N_12901);
nand U13961 (N_13961,N_13224,N_13400);
xnor U13962 (N_13962,N_13243,N_13470);
nand U13963 (N_13963,N_12779,N_12892);
xnor U13964 (N_13964,N_13174,N_13442);
xnor U13965 (N_13965,N_13075,N_12957);
nor U13966 (N_13966,N_13086,N_12867);
or U13967 (N_13967,N_13059,N_13010);
nand U13968 (N_13968,N_13227,N_13225);
nand U13969 (N_13969,N_12798,N_13404);
and U13970 (N_13970,N_12857,N_12943);
or U13971 (N_13971,N_12924,N_13030);
nor U13972 (N_13972,N_12764,N_13260);
and U13973 (N_13973,N_13478,N_13147);
xor U13974 (N_13974,N_12963,N_13332);
xnor U13975 (N_13975,N_13168,N_13399);
nor U13976 (N_13976,N_13138,N_13048);
nor U13977 (N_13977,N_12788,N_12760);
and U13978 (N_13978,N_13461,N_12965);
or U13979 (N_13979,N_13410,N_13185);
xor U13980 (N_13980,N_13124,N_12800);
nand U13981 (N_13981,N_13037,N_12856);
nor U13982 (N_13982,N_13417,N_13363);
and U13983 (N_13983,N_12753,N_12968);
and U13984 (N_13984,N_13105,N_13200);
xor U13985 (N_13985,N_12860,N_12939);
and U13986 (N_13986,N_12836,N_13170);
nor U13987 (N_13987,N_12867,N_13266);
nand U13988 (N_13988,N_13101,N_13124);
xor U13989 (N_13989,N_13156,N_12943);
nor U13990 (N_13990,N_12783,N_12833);
nand U13991 (N_13991,N_13333,N_13441);
nor U13992 (N_13992,N_13462,N_12834);
xnor U13993 (N_13993,N_13369,N_13284);
nand U13994 (N_13994,N_13192,N_13066);
and U13995 (N_13995,N_12930,N_12789);
or U13996 (N_13996,N_13361,N_13451);
nand U13997 (N_13997,N_13015,N_13130);
or U13998 (N_13998,N_13338,N_12807);
nor U13999 (N_13999,N_12940,N_13167);
nor U14000 (N_14000,N_12842,N_12988);
and U14001 (N_14001,N_12990,N_13316);
xnor U14002 (N_14002,N_13178,N_13257);
nand U14003 (N_14003,N_13005,N_12758);
nor U14004 (N_14004,N_13434,N_13191);
nand U14005 (N_14005,N_13135,N_13083);
xnor U14006 (N_14006,N_13261,N_13098);
nor U14007 (N_14007,N_13405,N_13441);
xor U14008 (N_14008,N_12853,N_13029);
nor U14009 (N_14009,N_12994,N_13264);
or U14010 (N_14010,N_13412,N_13123);
and U14011 (N_14011,N_13158,N_12910);
and U14012 (N_14012,N_13275,N_12864);
nand U14013 (N_14013,N_12858,N_13032);
or U14014 (N_14014,N_13449,N_13237);
and U14015 (N_14015,N_13156,N_13076);
nor U14016 (N_14016,N_13457,N_13454);
xor U14017 (N_14017,N_12757,N_12930);
or U14018 (N_14018,N_13442,N_13326);
nor U14019 (N_14019,N_13396,N_13248);
xor U14020 (N_14020,N_13320,N_13069);
and U14021 (N_14021,N_12923,N_13034);
or U14022 (N_14022,N_13008,N_13308);
nor U14023 (N_14023,N_13481,N_12988);
and U14024 (N_14024,N_13494,N_13262);
xor U14025 (N_14025,N_12754,N_13384);
nand U14026 (N_14026,N_13298,N_13329);
and U14027 (N_14027,N_13095,N_13246);
xnor U14028 (N_14028,N_13039,N_13179);
nor U14029 (N_14029,N_12795,N_13032);
nor U14030 (N_14030,N_12906,N_13265);
and U14031 (N_14031,N_13443,N_12836);
and U14032 (N_14032,N_12784,N_12907);
xnor U14033 (N_14033,N_13343,N_13424);
nor U14034 (N_14034,N_13156,N_12883);
or U14035 (N_14035,N_13067,N_13031);
and U14036 (N_14036,N_13260,N_13418);
xor U14037 (N_14037,N_12964,N_12921);
xor U14038 (N_14038,N_13411,N_12822);
nand U14039 (N_14039,N_12806,N_13003);
or U14040 (N_14040,N_12937,N_13208);
nor U14041 (N_14041,N_13389,N_13382);
xor U14042 (N_14042,N_13368,N_13382);
or U14043 (N_14043,N_13371,N_13477);
nor U14044 (N_14044,N_13105,N_13428);
or U14045 (N_14045,N_13196,N_13314);
and U14046 (N_14046,N_13282,N_12912);
nor U14047 (N_14047,N_13463,N_13353);
and U14048 (N_14048,N_13316,N_13483);
and U14049 (N_14049,N_12771,N_13015);
or U14050 (N_14050,N_13178,N_13013);
or U14051 (N_14051,N_13248,N_13386);
xnor U14052 (N_14052,N_13436,N_13421);
or U14053 (N_14053,N_13116,N_12806);
and U14054 (N_14054,N_13354,N_13192);
nand U14055 (N_14055,N_13291,N_13383);
and U14056 (N_14056,N_13425,N_13192);
nor U14057 (N_14057,N_13061,N_12938);
or U14058 (N_14058,N_13010,N_13340);
and U14059 (N_14059,N_12992,N_13125);
xor U14060 (N_14060,N_13391,N_13070);
or U14061 (N_14061,N_13373,N_13310);
nand U14062 (N_14062,N_13223,N_12818);
xor U14063 (N_14063,N_13394,N_13103);
xnor U14064 (N_14064,N_12960,N_13194);
nand U14065 (N_14065,N_13382,N_12991);
or U14066 (N_14066,N_12981,N_13256);
nor U14067 (N_14067,N_13115,N_13208);
xnor U14068 (N_14068,N_13355,N_12963);
xnor U14069 (N_14069,N_13282,N_12766);
and U14070 (N_14070,N_13130,N_13308);
xor U14071 (N_14071,N_12764,N_12926);
xor U14072 (N_14072,N_13331,N_13393);
or U14073 (N_14073,N_13332,N_13085);
and U14074 (N_14074,N_12891,N_13364);
nor U14075 (N_14075,N_12907,N_13422);
nand U14076 (N_14076,N_12816,N_13343);
xnor U14077 (N_14077,N_12794,N_13263);
nand U14078 (N_14078,N_12909,N_13053);
xor U14079 (N_14079,N_13068,N_12890);
nor U14080 (N_14080,N_13270,N_13140);
nand U14081 (N_14081,N_13192,N_12755);
and U14082 (N_14082,N_13255,N_13266);
or U14083 (N_14083,N_12825,N_13040);
xor U14084 (N_14084,N_13384,N_12990);
or U14085 (N_14085,N_13379,N_13097);
or U14086 (N_14086,N_12832,N_12781);
xnor U14087 (N_14087,N_13324,N_12952);
and U14088 (N_14088,N_12962,N_13498);
nand U14089 (N_14089,N_13419,N_13112);
xnor U14090 (N_14090,N_13450,N_12854);
nor U14091 (N_14091,N_12908,N_12814);
and U14092 (N_14092,N_13082,N_12860);
or U14093 (N_14093,N_13090,N_13454);
nand U14094 (N_14094,N_13162,N_13476);
nand U14095 (N_14095,N_13159,N_12962);
nand U14096 (N_14096,N_13017,N_13028);
xnor U14097 (N_14097,N_12860,N_13381);
xnor U14098 (N_14098,N_13273,N_13402);
and U14099 (N_14099,N_13192,N_12840);
xor U14100 (N_14100,N_12794,N_12808);
or U14101 (N_14101,N_12879,N_12909);
or U14102 (N_14102,N_12853,N_12943);
nor U14103 (N_14103,N_13203,N_13016);
or U14104 (N_14104,N_13058,N_12805);
nand U14105 (N_14105,N_13044,N_13457);
or U14106 (N_14106,N_13147,N_12896);
or U14107 (N_14107,N_13020,N_13168);
and U14108 (N_14108,N_13380,N_13371);
and U14109 (N_14109,N_13238,N_13365);
or U14110 (N_14110,N_13039,N_13384);
and U14111 (N_14111,N_12938,N_13054);
nand U14112 (N_14112,N_12843,N_12754);
xor U14113 (N_14113,N_12757,N_12828);
xor U14114 (N_14114,N_13013,N_13286);
and U14115 (N_14115,N_12893,N_12971);
or U14116 (N_14116,N_13265,N_13193);
nand U14117 (N_14117,N_13367,N_12858);
or U14118 (N_14118,N_12888,N_13003);
nor U14119 (N_14119,N_12823,N_12987);
and U14120 (N_14120,N_12995,N_12756);
or U14121 (N_14121,N_13017,N_13446);
or U14122 (N_14122,N_12865,N_13136);
xnor U14123 (N_14123,N_13184,N_13216);
nor U14124 (N_14124,N_13257,N_13122);
and U14125 (N_14125,N_12799,N_12812);
xnor U14126 (N_14126,N_13472,N_13117);
xor U14127 (N_14127,N_13255,N_12977);
nor U14128 (N_14128,N_13000,N_13210);
and U14129 (N_14129,N_13264,N_13468);
xor U14130 (N_14130,N_12795,N_13189);
or U14131 (N_14131,N_12753,N_12984);
and U14132 (N_14132,N_13413,N_13494);
or U14133 (N_14133,N_13171,N_13257);
and U14134 (N_14134,N_13454,N_12892);
nand U14135 (N_14135,N_13155,N_13065);
nor U14136 (N_14136,N_12760,N_13383);
or U14137 (N_14137,N_13302,N_13340);
nand U14138 (N_14138,N_13189,N_13011);
xnor U14139 (N_14139,N_12926,N_12947);
xor U14140 (N_14140,N_13115,N_12793);
and U14141 (N_14141,N_12834,N_13467);
and U14142 (N_14142,N_13033,N_13232);
xnor U14143 (N_14143,N_13242,N_13403);
and U14144 (N_14144,N_13115,N_13419);
xor U14145 (N_14145,N_13198,N_13324);
and U14146 (N_14146,N_13335,N_13417);
nor U14147 (N_14147,N_12885,N_13458);
nand U14148 (N_14148,N_12908,N_13184);
nor U14149 (N_14149,N_13436,N_13111);
nand U14150 (N_14150,N_13474,N_12821);
xor U14151 (N_14151,N_12887,N_13224);
or U14152 (N_14152,N_12890,N_13249);
and U14153 (N_14153,N_13490,N_13130);
or U14154 (N_14154,N_13116,N_12868);
xor U14155 (N_14155,N_12844,N_13399);
and U14156 (N_14156,N_13356,N_13146);
nor U14157 (N_14157,N_13221,N_12865);
and U14158 (N_14158,N_13068,N_12951);
xnor U14159 (N_14159,N_12807,N_13438);
nand U14160 (N_14160,N_13487,N_13309);
nor U14161 (N_14161,N_13454,N_13004);
nor U14162 (N_14162,N_13279,N_13053);
xnor U14163 (N_14163,N_13489,N_13066);
and U14164 (N_14164,N_12947,N_13303);
nor U14165 (N_14165,N_12939,N_13217);
and U14166 (N_14166,N_12831,N_13202);
nor U14167 (N_14167,N_13125,N_13469);
nand U14168 (N_14168,N_13427,N_13141);
nand U14169 (N_14169,N_13196,N_12752);
nand U14170 (N_14170,N_12752,N_12855);
nand U14171 (N_14171,N_13380,N_13490);
xor U14172 (N_14172,N_13252,N_13416);
xor U14173 (N_14173,N_13366,N_13134);
nand U14174 (N_14174,N_12849,N_12946);
and U14175 (N_14175,N_12971,N_12847);
or U14176 (N_14176,N_13277,N_13292);
nand U14177 (N_14177,N_12812,N_13499);
nand U14178 (N_14178,N_13286,N_13464);
or U14179 (N_14179,N_13435,N_13094);
nor U14180 (N_14180,N_13182,N_13470);
or U14181 (N_14181,N_13450,N_12786);
or U14182 (N_14182,N_13469,N_13236);
nand U14183 (N_14183,N_12929,N_12905);
nor U14184 (N_14184,N_12897,N_13258);
nand U14185 (N_14185,N_12941,N_13469);
xor U14186 (N_14186,N_12942,N_13111);
nor U14187 (N_14187,N_13298,N_13202);
xor U14188 (N_14188,N_13050,N_13315);
nor U14189 (N_14189,N_13269,N_13227);
xor U14190 (N_14190,N_12902,N_12943);
xor U14191 (N_14191,N_12940,N_13218);
nor U14192 (N_14192,N_13090,N_13023);
or U14193 (N_14193,N_13057,N_13257);
nor U14194 (N_14194,N_13261,N_13007);
nor U14195 (N_14195,N_13260,N_12824);
xnor U14196 (N_14196,N_13357,N_12795);
nor U14197 (N_14197,N_13100,N_12990);
nand U14198 (N_14198,N_13246,N_13016);
or U14199 (N_14199,N_13270,N_13260);
or U14200 (N_14200,N_13161,N_13498);
xor U14201 (N_14201,N_13030,N_13418);
and U14202 (N_14202,N_13060,N_12855);
xor U14203 (N_14203,N_13294,N_12878);
or U14204 (N_14204,N_12934,N_12819);
xnor U14205 (N_14205,N_13196,N_13474);
xor U14206 (N_14206,N_13422,N_13441);
nor U14207 (N_14207,N_12958,N_12816);
nand U14208 (N_14208,N_13179,N_12853);
nor U14209 (N_14209,N_13445,N_12938);
or U14210 (N_14210,N_12949,N_13010);
nand U14211 (N_14211,N_12839,N_13139);
or U14212 (N_14212,N_13010,N_13219);
nor U14213 (N_14213,N_12970,N_13334);
nor U14214 (N_14214,N_13277,N_12913);
nor U14215 (N_14215,N_13431,N_12880);
nand U14216 (N_14216,N_12759,N_13225);
and U14217 (N_14217,N_13341,N_12898);
nand U14218 (N_14218,N_13243,N_13346);
nor U14219 (N_14219,N_13407,N_13317);
and U14220 (N_14220,N_13312,N_12817);
or U14221 (N_14221,N_12910,N_12852);
or U14222 (N_14222,N_13154,N_13009);
nor U14223 (N_14223,N_13173,N_13433);
or U14224 (N_14224,N_13452,N_12912);
xor U14225 (N_14225,N_13081,N_12959);
nand U14226 (N_14226,N_12808,N_12903);
nor U14227 (N_14227,N_12966,N_13210);
nand U14228 (N_14228,N_13031,N_13356);
nor U14229 (N_14229,N_13406,N_13156);
or U14230 (N_14230,N_13343,N_13022);
and U14231 (N_14231,N_12942,N_12973);
nand U14232 (N_14232,N_13337,N_13463);
xor U14233 (N_14233,N_13440,N_13405);
nor U14234 (N_14234,N_13480,N_13177);
or U14235 (N_14235,N_13311,N_13221);
nor U14236 (N_14236,N_12878,N_13050);
xor U14237 (N_14237,N_13189,N_13096);
and U14238 (N_14238,N_13077,N_12821);
or U14239 (N_14239,N_13254,N_13054);
nor U14240 (N_14240,N_13326,N_12798);
xor U14241 (N_14241,N_13398,N_13491);
and U14242 (N_14242,N_13284,N_13324);
or U14243 (N_14243,N_12965,N_12828);
nor U14244 (N_14244,N_13377,N_13150);
xor U14245 (N_14245,N_13167,N_12777);
or U14246 (N_14246,N_13453,N_13402);
or U14247 (N_14247,N_13012,N_12945);
nand U14248 (N_14248,N_13247,N_12964);
or U14249 (N_14249,N_12799,N_13317);
nor U14250 (N_14250,N_13965,N_14141);
and U14251 (N_14251,N_13794,N_14108);
or U14252 (N_14252,N_14102,N_13847);
nor U14253 (N_14253,N_13906,N_13845);
or U14254 (N_14254,N_14233,N_13797);
and U14255 (N_14255,N_14076,N_14061);
or U14256 (N_14256,N_13534,N_13935);
nor U14257 (N_14257,N_13814,N_14099);
nor U14258 (N_14258,N_14094,N_13866);
and U14259 (N_14259,N_14023,N_13701);
nand U14260 (N_14260,N_13816,N_13551);
or U14261 (N_14261,N_13919,N_13944);
nor U14262 (N_14262,N_14179,N_14161);
or U14263 (N_14263,N_13564,N_13711);
or U14264 (N_14264,N_13672,N_13954);
and U14265 (N_14265,N_13864,N_13706);
xnor U14266 (N_14266,N_13992,N_13779);
nor U14267 (N_14267,N_13913,N_13710);
or U14268 (N_14268,N_14009,N_13898);
nand U14269 (N_14269,N_13752,N_13975);
and U14270 (N_14270,N_14034,N_14190);
xor U14271 (N_14271,N_13940,N_14126);
nand U14272 (N_14272,N_13652,N_13715);
nor U14273 (N_14273,N_14085,N_14000);
or U14274 (N_14274,N_14051,N_13638);
and U14275 (N_14275,N_14014,N_14056);
nand U14276 (N_14276,N_13695,N_13583);
or U14277 (N_14277,N_13812,N_14052);
xor U14278 (N_14278,N_13744,N_13501);
and U14279 (N_14279,N_13737,N_14055);
and U14280 (N_14280,N_14020,N_13681);
nand U14281 (N_14281,N_14174,N_14155);
or U14282 (N_14282,N_14154,N_13663);
and U14283 (N_14283,N_13854,N_13735);
nor U14284 (N_14284,N_13575,N_13838);
xor U14285 (N_14285,N_14064,N_13630);
and U14286 (N_14286,N_14185,N_13951);
nor U14287 (N_14287,N_13956,N_14027);
or U14288 (N_14288,N_14216,N_14240);
and U14289 (N_14289,N_13559,N_13754);
nor U14290 (N_14290,N_14069,N_13668);
nor U14291 (N_14291,N_14160,N_13861);
xor U14292 (N_14292,N_14109,N_13932);
and U14293 (N_14293,N_14077,N_13660);
xnor U14294 (N_14294,N_14128,N_13768);
nor U14295 (N_14295,N_13871,N_13533);
nor U14296 (N_14296,N_13820,N_13922);
xor U14297 (N_14297,N_13863,N_13772);
or U14298 (N_14298,N_13662,N_13896);
and U14299 (N_14299,N_13811,N_13617);
and U14300 (N_14300,N_13916,N_14175);
or U14301 (N_14301,N_14138,N_13709);
and U14302 (N_14302,N_13707,N_13817);
nor U14303 (N_14303,N_13742,N_13597);
and U14304 (N_14304,N_13540,N_13565);
and U14305 (N_14305,N_13923,N_13795);
nor U14306 (N_14306,N_14242,N_13598);
nor U14307 (N_14307,N_14123,N_13560);
and U14308 (N_14308,N_13552,N_14247);
or U14309 (N_14309,N_13719,N_14049);
nor U14310 (N_14310,N_13542,N_14137);
xor U14311 (N_14311,N_13971,N_13949);
or U14312 (N_14312,N_13897,N_13846);
and U14313 (N_14313,N_13569,N_13986);
nor U14314 (N_14314,N_14186,N_13982);
xnor U14315 (N_14315,N_13958,N_13642);
xor U14316 (N_14316,N_13925,N_14196);
xor U14317 (N_14317,N_13733,N_13789);
and U14318 (N_14318,N_13646,N_14237);
nor U14319 (N_14319,N_13624,N_13556);
nand U14320 (N_14320,N_14243,N_13786);
or U14321 (N_14321,N_13953,N_13902);
xor U14322 (N_14322,N_14088,N_14101);
nor U14323 (N_14323,N_13836,N_13834);
xor U14324 (N_14324,N_13527,N_13582);
or U14325 (N_14325,N_14112,N_13833);
nor U14326 (N_14326,N_14072,N_13558);
or U14327 (N_14327,N_13800,N_13623);
xnor U14328 (N_14328,N_13568,N_13592);
nand U14329 (N_14329,N_13764,N_13978);
and U14330 (N_14330,N_13718,N_13887);
and U14331 (N_14331,N_14092,N_14036);
or U14332 (N_14332,N_14035,N_14012);
or U14333 (N_14333,N_13792,N_13507);
nand U14334 (N_14334,N_13543,N_13665);
or U14335 (N_14335,N_14083,N_13815);
and U14336 (N_14336,N_14145,N_13591);
nand U14337 (N_14337,N_14231,N_14060);
and U14338 (N_14338,N_13872,N_14223);
xnor U14339 (N_14339,N_13536,N_14227);
xor U14340 (N_14340,N_14224,N_14149);
nand U14341 (N_14341,N_13673,N_14037);
nor U14342 (N_14342,N_13831,N_14024);
nor U14343 (N_14343,N_14229,N_13875);
xor U14344 (N_14344,N_14158,N_13827);
nand U14345 (N_14345,N_13850,N_14093);
nor U14346 (N_14346,N_13927,N_13911);
nor U14347 (N_14347,N_13757,N_14080);
nor U14348 (N_14348,N_13849,N_13553);
nor U14349 (N_14349,N_14122,N_13621);
xor U14350 (N_14350,N_14063,N_13717);
or U14351 (N_14351,N_14022,N_14147);
or U14352 (N_14352,N_13513,N_13781);
nor U14353 (N_14353,N_14095,N_13545);
xnor U14354 (N_14354,N_14048,N_14188);
or U14355 (N_14355,N_13622,N_13539);
xor U14356 (N_14356,N_14198,N_13566);
nand U14357 (N_14357,N_13918,N_14235);
nand U14358 (N_14358,N_13793,N_13782);
nand U14359 (N_14359,N_13937,N_14065);
xor U14360 (N_14360,N_13889,N_14004);
nand U14361 (N_14361,N_13899,N_14070);
or U14362 (N_14362,N_13685,N_13712);
nor U14363 (N_14363,N_13761,N_13508);
nor U14364 (N_14364,N_13878,N_13810);
nor U14365 (N_14365,N_13999,N_13941);
or U14366 (N_14366,N_13517,N_14038);
nor U14367 (N_14367,N_13968,N_14017);
nand U14368 (N_14368,N_14210,N_13704);
or U14369 (N_14369,N_13518,N_14135);
nand U14370 (N_14370,N_13577,N_13868);
or U14371 (N_14371,N_13851,N_13914);
xor U14372 (N_14372,N_14238,N_13607);
nand U14373 (N_14373,N_13938,N_13778);
xor U14374 (N_14374,N_14183,N_13599);
or U14375 (N_14375,N_14218,N_13874);
nand U14376 (N_14376,N_13516,N_13666);
or U14377 (N_14377,N_14166,N_13555);
and U14378 (N_14378,N_13580,N_13505);
and U14379 (N_14379,N_14002,N_13741);
and U14380 (N_14380,N_13691,N_13588);
nor U14381 (N_14381,N_14184,N_13759);
or U14382 (N_14382,N_14140,N_13586);
nand U14383 (N_14383,N_14221,N_13842);
xor U14384 (N_14384,N_14200,N_14030);
and U14385 (N_14385,N_14234,N_13581);
and U14386 (N_14386,N_13809,N_13824);
and U14387 (N_14387,N_13546,N_13694);
xnor U14388 (N_14388,N_13578,N_13618);
and U14389 (N_14389,N_13912,N_13979);
or U14390 (N_14390,N_13869,N_13720);
nand U14391 (N_14391,N_13983,N_14236);
nor U14392 (N_14392,N_13561,N_13512);
nand U14393 (N_14393,N_14195,N_14084);
nand U14394 (N_14394,N_13819,N_13880);
nor U14395 (N_14395,N_14033,N_13727);
or U14396 (N_14396,N_14119,N_13848);
xor U14397 (N_14397,N_13736,N_13840);
nand U14398 (N_14398,N_13526,N_13893);
xor U14399 (N_14399,N_13593,N_14150);
nor U14400 (N_14400,N_13960,N_13945);
and U14401 (N_14401,N_13544,N_13799);
xor U14402 (N_14402,N_13659,N_14098);
or U14403 (N_14403,N_13500,N_14040);
and U14404 (N_14404,N_13749,N_13620);
and U14405 (N_14405,N_13760,N_13901);
and U14406 (N_14406,N_13839,N_13557);
nand U14407 (N_14407,N_13683,N_14073);
nand U14408 (N_14408,N_14205,N_14230);
xnor U14409 (N_14409,N_13957,N_13947);
nor U14410 (N_14410,N_14213,N_14097);
nand U14411 (N_14411,N_13867,N_14197);
nand U14412 (N_14412,N_13939,N_13686);
xor U14413 (N_14413,N_14136,N_13969);
or U14414 (N_14414,N_14071,N_13931);
xor U14415 (N_14415,N_13521,N_13802);
and U14416 (N_14416,N_13791,N_13762);
and U14417 (N_14417,N_13567,N_14127);
nand U14418 (N_14418,N_13699,N_13635);
nor U14419 (N_14419,N_13651,N_13787);
nand U14420 (N_14420,N_14054,N_13855);
nor U14421 (N_14421,N_14181,N_14176);
xnor U14422 (N_14422,N_14110,N_14103);
xor U14423 (N_14423,N_13783,N_13502);
nor U14424 (N_14424,N_13882,N_13900);
nor U14425 (N_14425,N_14209,N_13728);
nor U14426 (N_14426,N_13770,N_13675);
xor U14427 (N_14427,N_14042,N_13628);
or U14428 (N_14428,N_14228,N_13693);
and U14429 (N_14429,N_13860,N_13589);
xnor U14430 (N_14430,N_14182,N_13639);
and U14431 (N_14431,N_13818,N_13780);
nand U14432 (N_14432,N_13645,N_13637);
or U14433 (N_14433,N_13773,N_13790);
xnor U14434 (N_14434,N_13682,N_13529);
nand U14435 (N_14435,N_13629,N_14162);
nor U14436 (N_14436,N_13511,N_13751);
xor U14437 (N_14437,N_14146,N_14019);
or U14438 (N_14438,N_13977,N_13532);
nor U14439 (N_14439,N_13857,N_14118);
xnor U14440 (N_14440,N_13808,N_13933);
nor U14441 (N_14441,N_14001,N_14194);
nor U14442 (N_14442,N_13837,N_13876);
nor U14443 (N_14443,N_14131,N_13509);
and U14444 (N_14444,N_14082,N_14178);
and U14445 (N_14445,N_13649,N_13822);
or U14446 (N_14446,N_13655,N_13604);
or U14447 (N_14447,N_14245,N_13995);
xor U14448 (N_14448,N_13547,N_13677);
or U14449 (N_14449,N_14057,N_13626);
xor U14450 (N_14450,N_13929,N_13858);
nand U14451 (N_14451,N_13585,N_13667);
nor U14452 (N_14452,N_13510,N_14116);
xnor U14453 (N_14453,N_14005,N_13627);
and U14454 (N_14454,N_13571,N_13826);
or U14455 (N_14455,N_13664,N_14003);
xnor U14456 (N_14456,N_14173,N_13894);
and U14457 (N_14457,N_14089,N_13881);
and U14458 (N_14458,N_13961,N_14217);
or U14459 (N_14459,N_13739,N_13714);
nand U14460 (N_14460,N_13550,N_13636);
or U14461 (N_14461,N_13669,N_14164);
nand U14462 (N_14462,N_13974,N_13616);
xor U14463 (N_14463,N_13563,N_13909);
or U14464 (N_14464,N_14171,N_13554);
nand U14465 (N_14465,N_13796,N_13807);
nand U14466 (N_14466,N_13753,N_14100);
nor U14467 (N_14467,N_13997,N_13688);
nand U14468 (N_14468,N_14239,N_14011);
nand U14469 (N_14469,N_13702,N_14091);
xor U14470 (N_14470,N_13985,N_13803);
nor U14471 (N_14471,N_13926,N_14177);
nand U14472 (N_14472,N_13633,N_13967);
or U14473 (N_14473,N_13562,N_13724);
nor U14474 (N_14474,N_13679,N_13703);
nor U14475 (N_14475,N_14244,N_14151);
or U14476 (N_14476,N_13804,N_14029);
nor U14477 (N_14477,N_13687,N_13530);
nand U14478 (N_14478,N_13943,N_14081);
and U14479 (N_14479,N_13998,N_13613);
nand U14480 (N_14480,N_14222,N_13601);
and U14481 (N_14481,N_13784,N_13722);
xnor U14482 (N_14482,N_13531,N_13734);
nand U14483 (N_14483,N_13619,N_13924);
or U14484 (N_14484,N_13747,N_14220);
or U14485 (N_14485,N_14246,N_13821);
nor U14486 (N_14486,N_13595,N_14066);
and U14487 (N_14487,N_14139,N_14006);
or U14488 (N_14488,N_13600,N_14191);
nand U14489 (N_14489,N_13689,N_13934);
and U14490 (N_14490,N_13692,N_14044);
nor U14491 (N_14491,N_14053,N_14189);
nand U14492 (N_14492,N_14248,N_13964);
nor U14493 (N_14493,N_13523,N_14045);
nor U14494 (N_14494,N_13989,N_13657);
nand U14495 (N_14495,N_14168,N_13859);
and U14496 (N_14496,N_13972,N_13862);
xor U14497 (N_14497,N_13920,N_14018);
or U14498 (N_14498,N_13708,N_13548);
and U14499 (N_14499,N_13603,N_14013);
xor U14500 (N_14500,N_13643,N_13769);
nand U14501 (N_14501,N_13541,N_14021);
nor U14502 (N_14502,N_13654,N_14062);
nor U14503 (N_14503,N_13835,N_13713);
nand U14504 (N_14504,N_14193,N_14047);
or U14505 (N_14505,N_13515,N_14159);
nand U14506 (N_14506,N_13765,N_14219);
xnor U14507 (N_14507,N_14152,N_14132);
or U14508 (N_14508,N_14167,N_14199);
nor U14509 (N_14509,N_13806,N_13885);
xor U14510 (N_14510,N_14212,N_14117);
or U14511 (N_14511,N_13584,N_14153);
xnor U14512 (N_14512,N_13525,N_13519);
xor U14513 (N_14513,N_13825,N_13886);
and U14514 (N_14514,N_13955,N_13549);
nand U14515 (N_14515,N_13930,N_14039);
and U14516 (N_14516,N_14043,N_13748);
and U14517 (N_14517,N_13981,N_13873);
or U14518 (N_14518,N_14165,N_13767);
or U14519 (N_14519,N_14113,N_13573);
or U14520 (N_14520,N_13883,N_14106);
nor U14521 (N_14521,N_14215,N_13608);
and U14522 (N_14522,N_13731,N_13705);
or U14523 (N_14523,N_14249,N_13606);
xnor U14524 (N_14524,N_13884,N_14031);
and U14525 (N_14525,N_14026,N_13579);
xnor U14526 (N_14526,N_13776,N_13987);
nor U14527 (N_14527,N_13750,N_14107);
and U14528 (N_14528,N_14096,N_14015);
nand U14529 (N_14529,N_13805,N_14226);
and U14530 (N_14530,N_13631,N_14008);
nor U14531 (N_14531,N_14058,N_13976);
xor U14532 (N_14532,N_13504,N_13970);
nand U14533 (N_14533,N_13538,N_13828);
and U14534 (N_14534,N_13832,N_14121);
and U14535 (N_14535,N_13950,N_13890);
or U14536 (N_14536,N_13936,N_13946);
nand U14537 (N_14537,N_13766,N_13948);
or U14538 (N_14538,N_13853,N_14090);
nor U14539 (N_14539,N_13910,N_14124);
and U14540 (N_14540,N_14208,N_13865);
xnor U14541 (N_14541,N_13678,N_13605);
or U14542 (N_14542,N_14211,N_13590);
xor U14543 (N_14543,N_14105,N_13777);
nand U14544 (N_14544,N_14010,N_13506);
nand U14545 (N_14545,N_14144,N_13907);
nor U14546 (N_14546,N_13915,N_14115);
nor U14547 (N_14547,N_14079,N_14202);
and U14548 (N_14548,N_13729,N_14046);
xnor U14549 (N_14549,N_13723,N_14059);
and U14550 (N_14550,N_13917,N_13756);
and U14551 (N_14551,N_13813,N_14163);
and U14552 (N_14552,N_13537,N_13574);
nand U14553 (N_14553,N_13632,N_13661);
and U14554 (N_14554,N_13801,N_13676);
and U14555 (N_14555,N_13830,N_14130);
nand U14556 (N_14556,N_13746,N_13587);
or U14557 (N_14557,N_14111,N_13908);
nor U14558 (N_14558,N_13829,N_14204);
xnor U14559 (N_14559,N_14169,N_13647);
and U14560 (N_14560,N_13697,N_13528);
xor U14561 (N_14561,N_13973,N_13641);
and U14562 (N_14562,N_13634,N_13743);
and U14563 (N_14563,N_14087,N_14068);
nor U14564 (N_14564,N_13658,N_14125);
xnor U14565 (N_14565,N_13966,N_14086);
or U14566 (N_14566,N_13841,N_13520);
or U14567 (N_14567,N_13503,N_13903);
xor U14568 (N_14568,N_13596,N_13905);
or U14569 (N_14569,N_13962,N_13670);
nand U14570 (N_14570,N_14133,N_14157);
nand U14571 (N_14571,N_14120,N_13514);
and U14572 (N_14572,N_13730,N_13798);
nand U14573 (N_14573,N_13644,N_13877);
nand U14574 (N_14574,N_14032,N_13648);
nor U14575 (N_14575,N_13844,N_14025);
nand U14576 (N_14576,N_13892,N_14075);
or U14577 (N_14577,N_14192,N_13653);
xnor U14578 (N_14578,N_13696,N_14241);
nand U14579 (N_14579,N_13610,N_14074);
nand U14580 (N_14580,N_13888,N_13674);
xor U14581 (N_14581,N_14225,N_13640);
and U14582 (N_14582,N_13959,N_13785);
or U14583 (N_14583,N_14007,N_13843);
xor U14584 (N_14584,N_13984,N_13602);
and U14585 (N_14585,N_14041,N_13726);
and U14586 (N_14586,N_13522,N_13576);
xor U14587 (N_14587,N_13725,N_13993);
or U14588 (N_14588,N_13952,N_13721);
or U14589 (N_14589,N_13614,N_14016);
or U14590 (N_14590,N_13771,N_14187);
nand U14591 (N_14591,N_13921,N_13788);
and U14592 (N_14592,N_13996,N_13856);
and U14593 (N_14593,N_13775,N_14172);
nor U14594 (N_14594,N_13570,N_13904);
or U14595 (N_14595,N_13716,N_14143);
or U14596 (N_14596,N_14104,N_13680);
and U14597 (N_14597,N_14142,N_14180);
xor U14598 (N_14598,N_14214,N_14067);
and U14599 (N_14599,N_14203,N_13732);
xor U14600 (N_14600,N_13870,N_13758);
and U14601 (N_14601,N_13942,N_14050);
and U14602 (N_14602,N_13594,N_13990);
or U14603 (N_14603,N_13994,N_13738);
nand U14604 (N_14604,N_13891,N_13988);
or U14605 (N_14605,N_13625,N_13852);
xnor U14606 (N_14606,N_13612,N_14232);
and U14607 (N_14607,N_13609,N_13963);
nor U14608 (N_14608,N_13895,N_13740);
or U14609 (N_14609,N_14114,N_13671);
xor U14610 (N_14610,N_14201,N_13684);
xnor U14611 (N_14611,N_13980,N_13572);
nor U14612 (N_14612,N_14129,N_14206);
nand U14613 (N_14613,N_13823,N_14028);
xor U14614 (N_14614,N_13879,N_13991);
and U14615 (N_14615,N_14078,N_13928);
xnor U14616 (N_14616,N_13611,N_14148);
nor U14617 (N_14617,N_13615,N_13763);
nor U14618 (N_14618,N_14207,N_14170);
nor U14619 (N_14619,N_13774,N_13755);
nor U14620 (N_14620,N_13700,N_14156);
and U14621 (N_14621,N_13535,N_13698);
or U14622 (N_14622,N_13745,N_13524);
xnor U14623 (N_14623,N_13656,N_13650);
nand U14624 (N_14624,N_14134,N_13690);
xnor U14625 (N_14625,N_14004,N_13648);
or U14626 (N_14626,N_13787,N_13865);
nor U14627 (N_14627,N_13897,N_13549);
or U14628 (N_14628,N_14184,N_13966);
nor U14629 (N_14629,N_13587,N_13525);
nor U14630 (N_14630,N_13631,N_14185);
xor U14631 (N_14631,N_13602,N_13720);
or U14632 (N_14632,N_13603,N_13931);
or U14633 (N_14633,N_13902,N_14194);
nand U14634 (N_14634,N_13915,N_14014);
and U14635 (N_14635,N_13974,N_13694);
nor U14636 (N_14636,N_13743,N_13575);
or U14637 (N_14637,N_13876,N_13902);
nor U14638 (N_14638,N_14095,N_13870);
and U14639 (N_14639,N_13502,N_14154);
and U14640 (N_14640,N_13634,N_14128);
and U14641 (N_14641,N_13805,N_13689);
xor U14642 (N_14642,N_13525,N_13957);
nand U14643 (N_14643,N_13909,N_13794);
or U14644 (N_14644,N_14198,N_13876);
nand U14645 (N_14645,N_14131,N_14093);
nand U14646 (N_14646,N_13955,N_14094);
nor U14647 (N_14647,N_14097,N_14027);
and U14648 (N_14648,N_13856,N_13683);
and U14649 (N_14649,N_13541,N_13562);
and U14650 (N_14650,N_13631,N_13867);
or U14651 (N_14651,N_14073,N_14027);
and U14652 (N_14652,N_13728,N_13915);
xor U14653 (N_14653,N_13823,N_13881);
xnor U14654 (N_14654,N_13793,N_13670);
nor U14655 (N_14655,N_13953,N_14024);
nand U14656 (N_14656,N_14027,N_14183);
xor U14657 (N_14657,N_14221,N_13990);
nand U14658 (N_14658,N_13647,N_13640);
or U14659 (N_14659,N_14164,N_13748);
or U14660 (N_14660,N_13861,N_14079);
xor U14661 (N_14661,N_13607,N_13611);
xnor U14662 (N_14662,N_13684,N_13929);
nand U14663 (N_14663,N_14134,N_13568);
or U14664 (N_14664,N_13585,N_13615);
and U14665 (N_14665,N_14154,N_14145);
nor U14666 (N_14666,N_13921,N_13937);
nand U14667 (N_14667,N_13844,N_13859);
nand U14668 (N_14668,N_13802,N_14051);
nand U14669 (N_14669,N_13662,N_13535);
xor U14670 (N_14670,N_14239,N_13967);
nand U14671 (N_14671,N_14012,N_13831);
or U14672 (N_14672,N_13832,N_14027);
and U14673 (N_14673,N_13551,N_14157);
xnor U14674 (N_14674,N_13757,N_13799);
and U14675 (N_14675,N_13528,N_13633);
nor U14676 (N_14676,N_14195,N_13703);
or U14677 (N_14677,N_13988,N_13554);
and U14678 (N_14678,N_13758,N_14121);
xor U14679 (N_14679,N_14196,N_13619);
nand U14680 (N_14680,N_14099,N_14052);
or U14681 (N_14681,N_13582,N_13913);
nand U14682 (N_14682,N_13616,N_14142);
nor U14683 (N_14683,N_13876,N_13985);
and U14684 (N_14684,N_13738,N_13700);
nor U14685 (N_14685,N_13712,N_14220);
nand U14686 (N_14686,N_13785,N_14183);
nand U14687 (N_14687,N_13565,N_13996);
or U14688 (N_14688,N_14226,N_13706);
and U14689 (N_14689,N_13766,N_13706);
nor U14690 (N_14690,N_13701,N_14014);
xor U14691 (N_14691,N_13691,N_13805);
nand U14692 (N_14692,N_13901,N_13910);
or U14693 (N_14693,N_14249,N_14100);
xnor U14694 (N_14694,N_13528,N_14022);
nand U14695 (N_14695,N_14021,N_14146);
or U14696 (N_14696,N_13522,N_13818);
or U14697 (N_14697,N_13832,N_13805);
and U14698 (N_14698,N_14249,N_14026);
nor U14699 (N_14699,N_13892,N_13771);
and U14700 (N_14700,N_13792,N_13820);
nor U14701 (N_14701,N_14215,N_14109);
and U14702 (N_14702,N_13535,N_13809);
nand U14703 (N_14703,N_13568,N_13930);
xor U14704 (N_14704,N_13641,N_13954);
nand U14705 (N_14705,N_13951,N_14219);
xor U14706 (N_14706,N_13646,N_14099);
nand U14707 (N_14707,N_13701,N_14056);
nand U14708 (N_14708,N_13509,N_13967);
nor U14709 (N_14709,N_14108,N_13523);
or U14710 (N_14710,N_13621,N_13885);
and U14711 (N_14711,N_13628,N_14061);
nand U14712 (N_14712,N_14015,N_13621);
xnor U14713 (N_14713,N_14124,N_13768);
and U14714 (N_14714,N_14134,N_14031);
and U14715 (N_14715,N_13705,N_13503);
xnor U14716 (N_14716,N_14178,N_13554);
and U14717 (N_14717,N_14124,N_13601);
or U14718 (N_14718,N_13668,N_13503);
nor U14719 (N_14719,N_13699,N_14174);
nand U14720 (N_14720,N_13911,N_13912);
or U14721 (N_14721,N_13747,N_13517);
xor U14722 (N_14722,N_13746,N_13801);
or U14723 (N_14723,N_13734,N_13525);
or U14724 (N_14724,N_13671,N_13798);
nand U14725 (N_14725,N_13857,N_13695);
nor U14726 (N_14726,N_14087,N_13729);
nor U14727 (N_14727,N_13917,N_13806);
and U14728 (N_14728,N_13704,N_14009);
xor U14729 (N_14729,N_14224,N_13712);
nor U14730 (N_14730,N_13716,N_13960);
or U14731 (N_14731,N_14191,N_14187);
xnor U14732 (N_14732,N_13885,N_13565);
and U14733 (N_14733,N_13860,N_13661);
nand U14734 (N_14734,N_13712,N_13737);
nor U14735 (N_14735,N_13656,N_14123);
nand U14736 (N_14736,N_13851,N_13668);
nand U14737 (N_14737,N_14231,N_13615);
and U14738 (N_14738,N_14083,N_14223);
nand U14739 (N_14739,N_13615,N_13880);
or U14740 (N_14740,N_13703,N_13875);
xnor U14741 (N_14741,N_14001,N_13735);
xor U14742 (N_14742,N_13798,N_13555);
nor U14743 (N_14743,N_13858,N_13735);
or U14744 (N_14744,N_13898,N_14166);
nand U14745 (N_14745,N_14203,N_14024);
and U14746 (N_14746,N_13846,N_13874);
or U14747 (N_14747,N_13603,N_14056);
nor U14748 (N_14748,N_14026,N_14047);
and U14749 (N_14749,N_13896,N_13768);
nand U14750 (N_14750,N_13538,N_14234);
and U14751 (N_14751,N_13874,N_13895);
nor U14752 (N_14752,N_14130,N_13503);
or U14753 (N_14753,N_13919,N_13789);
nor U14754 (N_14754,N_13976,N_13665);
nand U14755 (N_14755,N_13579,N_14131);
xor U14756 (N_14756,N_13793,N_13750);
xor U14757 (N_14757,N_14201,N_13786);
or U14758 (N_14758,N_13822,N_13500);
xor U14759 (N_14759,N_13546,N_13630);
nand U14760 (N_14760,N_13528,N_13644);
nand U14761 (N_14761,N_13545,N_13513);
nand U14762 (N_14762,N_13791,N_13672);
nand U14763 (N_14763,N_13553,N_13877);
nor U14764 (N_14764,N_13869,N_13762);
or U14765 (N_14765,N_13663,N_13704);
or U14766 (N_14766,N_13817,N_13599);
or U14767 (N_14767,N_13838,N_13655);
and U14768 (N_14768,N_13614,N_14218);
or U14769 (N_14769,N_13540,N_13632);
or U14770 (N_14770,N_14169,N_14139);
or U14771 (N_14771,N_13775,N_14206);
xnor U14772 (N_14772,N_14106,N_14170);
and U14773 (N_14773,N_14053,N_13654);
and U14774 (N_14774,N_13885,N_14069);
or U14775 (N_14775,N_13814,N_13549);
xor U14776 (N_14776,N_13878,N_13674);
or U14777 (N_14777,N_13622,N_13997);
xor U14778 (N_14778,N_13853,N_14233);
xnor U14779 (N_14779,N_14224,N_14031);
nor U14780 (N_14780,N_13769,N_13596);
xor U14781 (N_14781,N_13587,N_13872);
nor U14782 (N_14782,N_13726,N_13604);
nor U14783 (N_14783,N_13834,N_13548);
xor U14784 (N_14784,N_13780,N_14110);
xnor U14785 (N_14785,N_13934,N_14155);
nand U14786 (N_14786,N_13955,N_14106);
xnor U14787 (N_14787,N_13942,N_13848);
nand U14788 (N_14788,N_14130,N_13859);
nand U14789 (N_14789,N_13647,N_13959);
nor U14790 (N_14790,N_14014,N_14136);
xor U14791 (N_14791,N_14124,N_13702);
nand U14792 (N_14792,N_13797,N_14009);
and U14793 (N_14793,N_14235,N_14169);
or U14794 (N_14794,N_13532,N_13524);
or U14795 (N_14795,N_13798,N_13847);
and U14796 (N_14796,N_13832,N_13972);
and U14797 (N_14797,N_13528,N_13588);
nand U14798 (N_14798,N_14215,N_13669);
and U14799 (N_14799,N_13566,N_13588);
nand U14800 (N_14800,N_14099,N_14167);
and U14801 (N_14801,N_13862,N_13552);
or U14802 (N_14802,N_13867,N_13844);
and U14803 (N_14803,N_14060,N_13824);
or U14804 (N_14804,N_13523,N_14077);
or U14805 (N_14805,N_14172,N_13938);
xnor U14806 (N_14806,N_14077,N_13907);
or U14807 (N_14807,N_13648,N_14111);
nor U14808 (N_14808,N_13871,N_13777);
or U14809 (N_14809,N_14157,N_13706);
xor U14810 (N_14810,N_14040,N_14134);
nand U14811 (N_14811,N_14118,N_13711);
or U14812 (N_14812,N_13716,N_13978);
or U14813 (N_14813,N_13575,N_13760);
and U14814 (N_14814,N_14246,N_13511);
nor U14815 (N_14815,N_13604,N_14171);
nor U14816 (N_14816,N_13782,N_13834);
or U14817 (N_14817,N_13508,N_13707);
and U14818 (N_14818,N_13667,N_13589);
nand U14819 (N_14819,N_13755,N_13915);
nand U14820 (N_14820,N_13860,N_13856);
or U14821 (N_14821,N_13837,N_14031);
nor U14822 (N_14822,N_13705,N_13897);
xor U14823 (N_14823,N_14020,N_13868);
xnor U14824 (N_14824,N_13651,N_14119);
nand U14825 (N_14825,N_14116,N_14065);
xnor U14826 (N_14826,N_13780,N_13744);
nor U14827 (N_14827,N_14148,N_13918);
and U14828 (N_14828,N_13613,N_13770);
and U14829 (N_14829,N_13797,N_14139);
xor U14830 (N_14830,N_14022,N_13523);
nor U14831 (N_14831,N_14074,N_14115);
xnor U14832 (N_14832,N_14142,N_14192);
nor U14833 (N_14833,N_13656,N_13784);
nor U14834 (N_14834,N_14158,N_14216);
nand U14835 (N_14835,N_14162,N_13586);
xnor U14836 (N_14836,N_13931,N_14242);
nand U14837 (N_14837,N_13533,N_13757);
xor U14838 (N_14838,N_13842,N_14181);
nand U14839 (N_14839,N_13702,N_14247);
xor U14840 (N_14840,N_14150,N_14080);
and U14841 (N_14841,N_13569,N_13897);
and U14842 (N_14842,N_14246,N_13958);
nor U14843 (N_14843,N_13757,N_13596);
xor U14844 (N_14844,N_13743,N_14123);
or U14845 (N_14845,N_14238,N_13653);
nand U14846 (N_14846,N_13687,N_13893);
and U14847 (N_14847,N_13502,N_13835);
nor U14848 (N_14848,N_13812,N_14108);
nor U14849 (N_14849,N_13645,N_13664);
and U14850 (N_14850,N_13626,N_14198);
xor U14851 (N_14851,N_14246,N_13778);
xor U14852 (N_14852,N_13519,N_13886);
xnor U14853 (N_14853,N_14071,N_13850);
nand U14854 (N_14854,N_13960,N_13963);
xor U14855 (N_14855,N_14046,N_13716);
and U14856 (N_14856,N_14073,N_13763);
or U14857 (N_14857,N_13823,N_13743);
xor U14858 (N_14858,N_14101,N_13629);
xnor U14859 (N_14859,N_14033,N_13958);
nand U14860 (N_14860,N_13932,N_13831);
or U14861 (N_14861,N_13867,N_13790);
nand U14862 (N_14862,N_13628,N_13825);
or U14863 (N_14863,N_13769,N_13652);
xor U14864 (N_14864,N_13638,N_13699);
nor U14865 (N_14865,N_13821,N_13862);
xor U14866 (N_14866,N_13718,N_13804);
nand U14867 (N_14867,N_14199,N_13601);
nor U14868 (N_14868,N_13768,N_13847);
nor U14869 (N_14869,N_13527,N_13911);
nand U14870 (N_14870,N_13579,N_14197);
and U14871 (N_14871,N_14105,N_13686);
xor U14872 (N_14872,N_13532,N_14116);
nand U14873 (N_14873,N_14148,N_14014);
xor U14874 (N_14874,N_13918,N_13981);
nor U14875 (N_14875,N_13992,N_13920);
xor U14876 (N_14876,N_14021,N_14218);
or U14877 (N_14877,N_13748,N_14107);
nor U14878 (N_14878,N_14141,N_13960);
xnor U14879 (N_14879,N_14000,N_14115);
nand U14880 (N_14880,N_14099,N_13797);
xnor U14881 (N_14881,N_13937,N_13587);
nor U14882 (N_14882,N_13828,N_13551);
and U14883 (N_14883,N_13604,N_14032);
nor U14884 (N_14884,N_13980,N_13840);
and U14885 (N_14885,N_14243,N_14010);
nand U14886 (N_14886,N_13961,N_14045);
nor U14887 (N_14887,N_14071,N_13620);
nor U14888 (N_14888,N_13642,N_13921);
xor U14889 (N_14889,N_13714,N_13841);
xor U14890 (N_14890,N_14040,N_13552);
xnor U14891 (N_14891,N_14081,N_13801);
xnor U14892 (N_14892,N_13745,N_13753);
xor U14893 (N_14893,N_14169,N_14069);
xor U14894 (N_14894,N_13602,N_13523);
nand U14895 (N_14895,N_13659,N_13619);
nand U14896 (N_14896,N_14038,N_14135);
or U14897 (N_14897,N_13696,N_14049);
or U14898 (N_14898,N_13625,N_13819);
xnor U14899 (N_14899,N_13959,N_14191);
nor U14900 (N_14900,N_13579,N_13613);
and U14901 (N_14901,N_14162,N_13507);
nor U14902 (N_14902,N_14144,N_14041);
and U14903 (N_14903,N_13928,N_14005);
and U14904 (N_14904,N_13647,N_14173);
nor U14905 (N_14905,N_13759,N_14091);
xor U14906 (N_14906,N_13542,N_13848);
and U14907 (N_14907,N_13860,N_13745);
nand U14908 (N_14908,N_13614,N_13934);
xnor U14909 (N_14909,N_14214,N_14110);
xnor U14910 (N_14910,N_13566,N_13907);
or U14911 (N_14911,N_13794,N_13801);
nor U14912 (N_14912,N_14168,N_13804);
nand U14913 (N_14913,N_13761,N_13831);
nand U14914 (N_14914,N_13692,N_13815);
nand U14915 (N_14915,N_13725,N_13721);
xor U14916 (N_14916,N_14180,N_13664);
nor U14917 (N_14917,N_13514,N_13521);
xnor U14918 (N_14918,N_13763,N_13834);
and U14919 (N_14919,N_14105,N_13933);
and U14920 (N_14920,N_14221,N_13775);
or U14921 (N_14921,N_13649,N_14013);
or U14922 (N_14922,N_13895,N_13582);
and U14923 (N_14923,N_13675,N_14222);
and U14924 (N_14924,N_13780,N_14122);
nor U14925 (N_14925,N_13587,N_13854);
xor U14926 (N_14926,N_13913,N_13580);
xor U14927 (N_14927,N_14058,N_13857);
and U14928 (N_14928,N_13884,N_14062);
or U14929 (N_14929,N_13576,N_13907);
nor U14930 (N_14930,N_14043,N_13763);
nor U14931 (N_14931,N_14021,N_13691);
and U14932 (N_14932,N_13983,N_14161);
xnor U14933 (N_14933,N_13575,N_13660);
nand U14934 (N_14934,N_13817,N_13732);
nor U14935 (N_14935,N_13679,N_14236);
xor U14936 (N_14936,N_14055,N_14092);
xnor U14937 (N_14937,N_13995,N_13977);
nor U14938 (N_14938,N_13939,N_14104);
nor U14939 (N_14939,N_13783,N_13813);
xor U14940 (N_14940,N_14144,N_13529);
or U14941 (N_14941,N_13612,N_14080);
nor U14942 (N_14942,N_13814,N_14062);
nor U14943 (N_14943,N_13853,N_13743);
nor U14944 (N_14944,N_13794,N_14203);
nor U14945 (N_14945,N_14212,N_14014);
or U14946 (N_14946,N_13651,N_13824);
or U14947 (N_14947,N_13867,N_14069);
xor U14948 (N_14948,N_14211,N_13858);
and U14949 (N_14949,N_13609,N_13853);
xnor U14950 (N_14950,N_13857,N_13763);
and U14951 (N_14951,N_14089,N_14116);
and U14952 (N_14952,N_14167,N_13895);
nor U14953 (N_14953,N_14218,N_13604);
nand U14954 (N_14954,N_13836,N_13689);
xor U14955 (N_14955,N_13693,N_13803);
and U14956 (N_14956,N_13970,N_14005);
nand U14957 (N_14957,N_13806,N_13899);
nor U14958 (N_14958,N_14224,N_13657);
and U14959 (N_14959,N_13665,N_13547);
and U14960 (N_14960,N_13543,N_14086);
or U14961 (N_14961,N_13673,N_13721);
and U14962 (N_14962,N_13525,N_13608);
and U14963 (N_14963,N_13655,N_13771);
or U14964 (N_14964,N_14135,N_13894);
xor U14965 (N_14965,N_14168,N_14004);
or U14966 (N_14966,N_13551,N_13679);
and U14967 (N_14967,N_13963,N_14034);
xor U14968 (N_14968,N_13575,N_14233);
nor U14969 (N_14969,N_13893,N_13967);
and U14970 (N_14970,N_14089,N_14095);
nand U14971 (N_14971,N_13721,N_13906);
xnor U14972 (N_14972,N_13528,N_13518);
and U14973 (N_14973,N_13712,N_13568);
nor U14974 (N_14974,N_14150,N_13965);
or U14975 (N_14975,N_13606,N_14003);
or U14976 (N_14976,N_14110,N_13619);
or U14977 (N_14977,N_13693,N_13958);
and U14978 (N_14978,N_13773,N_13587);
nor U14979 (N_14979,N_13924,N_14137);
or U14980 (N_14980,N_13655,N_14139);
nand U14981 (N_14981,N_13864,N_13850);
xor U14982 (N_14982,N_13627,N_13555);
xnor U14983 (N_14983,N_14128,N_13840);
and U14984 (N_14984,N_13873,N_13982);
or U14985 (N_14985,N_13576,N_13774);
or U14986 (N_14986,N_13675,N_13905);
xor U14987 (N_14987,N_13708,N_13596);
and U14988 (N_14988,N_13946,N_13761);
or U14989 (N_14989,N_13834,N_13788);
and U14990 (N_14990,N_13640,N_13892);
and U14991 (N_14991,N_13712,N_13608);
nor U14992 (N_14992,N_13673,N_13872);
nor U14993 (N_14993,N_14214,N_13879);
nor U14994 (N_14994,N_13529,N_14083);
xnor U14995 (N_14995,N_13740,N_13614);
or U14996 (N_14996,N_14203,N_13846);
or U14997 (N_14997,N_14237,N_13511);
and U14998 (N_14998,N_13626,N_13795);
xnor U14999 (N_14999,N_13655,N_14178);
nand UO_0 (O_0,N_14444,N_14637);
nor UO_1 (O_1,N_14481,N_14964);
nand UO_2 (O_2,N_14610,N_14615);
nor UO_3 (O_3,N_14310,N_14771);
nand UO_4 (O_4,N_14435,N_14507);
nor UO_5 (O_5,N_14387,N_14355);
or UO_6 (O_6,N_14763,N_14775);
or UO_7 (O_7,N_14886,N_14519);
xnor UO_8 (O_8,N_14393,N_14357);
and UO_9 (O_9,N_14417,N_14450);
xnor UO_10 (O_10,N_14384,N_14822);
xnor UO_11 (O_11,N_14431,N_14858);
or UO_12 (O_12,N_14328,N_14787);
xor UO_13 (O_13,N_14604,N_14550);
and UO_14 (O_14,N_14506,N_14252);
or UO_15 (O_15,N_14802,N_14844);
or UO_16 (O_16,N_14380,N_14841);
xnor UO_17 (O_17,N_14962,N_14358);
nand UO_18 (O_18,N_14305,N_14752);
and UO_19 (O_19,N_14884,N_14260);
or UO_20 (O_20,N_14650,N_14491);
or UO_21 (O_21,N_14809,N_14983);
and UO_22 (O_22,N_14793,N_14979);
xnor UO_23 (O_23,N_14633,N_14508);
nand UO_24 (O_24,N_14390,N_14784);
or UO_25 (O_25,N_14535,N_14927);
and UO_26 (O_26,N_14383,N_14897);
xnor UO_27 (O_27,N_14833,N_14302);
or UO_28 (O_28,N_14422,N_14411);
nand UO_29 (O_29,N_14798,N_14915);
or UO_30 (O_30,N_14812,N_14902);
xnor UO_31 (O_31,N_14338,N_14482);
or UO_32 (O_32,N_14466,N_14708);
and UO_33 (O_33,N_14363,N_14926);
nor UO_34 (O_34,N_14746,N_14285);
nor UO_35 (O_35,N_14297,N_14627);
or UO_36 (O_36,N_14909,N_14683);
xnor UO_37 (O_37,N_14255,N_14547);
xor UO_38 (O_38,N_14301,N_14287);
nor UO_39 (O_39,N_14498,N_14726);
xnor UO_40 (O_40,N_14942,N_14439);
xor UO_41 (O_41,N_14666,N_14656);
nand UO_42 (O_42,N_14861,N_14665);
nor UO_43 (O_43,N_14334,N_14776);
or UO_44 (O_44,N_14441,N_14382);
xor UO_45 (O_45,N_14770,N_14894);
or UO_46 (O_46,N_14832,N_14376);
nand UO_47 (O_47,N_14663,N_14325);
or UO_48 (O_48,N_14349,N_14674);
nor UO_49 (O_49,N_14308,N_14572);
nor UO_50 (O_50,N_14702,N_14361);
and UO_51 (O_51,N_14473,N_14279);
nand UO_52 (O_52,N_14699,N_14531);
and UO_53 (O_53,N_14740,N_14961);
xor UO_54 (O_54,N_14596,N_14972);
nand UO_55 (O_55,N_14854,N_14324);
xnor UO_56 (O_56,N_14924,N_14703);
nand UO_57 (O_57,N_14658,N_14678);
or UO_58 (O_58,N_14944,N_14865);
xnor UO_59 (O_59,N_14590,N_14912);
nand UO_60 (O_60,N_14286,N_14456);
nand UO_61 (O_61,N_14985,N_14515);
or UO_62 (O_62,N_14753,N_14395);
nand UO_63 (O_63,N_14921,N_14373);
and UO_64 (O_64,N_14419,N_14354);
xor UO_65 (O_65,N_14367,N_14681);
xnor UO_66 (O_66,N_14957,N_14996);
nor UO_67 (O_67,N_14584,N_14513);
nor UO_68 (O_68,N_14738,N_14360);
nand UO_69 (O_69,N_14394,N_14309);
or UO_70 (O_70,N_14359,N_14953);
and UO_71 (O_71,N_14459,N_14404);
nand UO_72 (O_72,N_14322,N_14635);
nor UO_73 (O_73,N_14631,N_14789);
nor UO_74 (O_74,N_14568,N_14928);
nand UO_75 (O_75,N_14520,N_14378);
and UO_76 (O_76,N_14811,N_14407);
or UO_77 (O_77,N_14774,N_14552);
xnor UO_78 (O_78,N_14406,N_14478);
or UO_79 (O_79,N_14769,N_14619);
or UO_80 (O_80,N_14808,N_14867);
and UO_81 (O_81,N_14856,N_14881);
or UO_82 (O_82,N_14379,N_14689);
or UO_83 (O_83,N_14303,N_14267);
xnor UO_84 (O_84,N_14530,N_14644);
or UO_85 (O_85,N_14850,N_14313);
nand UO_86 (O_86,N_14791,N_14671);
nor UO_87 (O_87,N_14842,N_14602);
and UO_88 (O_88,N_14454,N_14721);
or UO_89 (O_89,N_14370,N_14931);
nor UO_90 (O_90,N_14722,N_14503);
xor UO_91 (O_91,N_14561,N_14609);
nor UO_92 (O_92,N_14877,N_14340);
or UO_93 (O_93,N_14668,N_14563);
nand UO_94 (O_94,N_14554,N_14480);
nor UO_95 (O_95,N_14460,N_14718);
and UO_96 (O_96,N_14262,N_14428);
or UO_97 (O_97,N_14664,N_14667);
or UO_98 (O_98,N_14589,N_14720);
nand UO_99 (O_99,N_14256,N_14599);
or UO_100 (O_100,N_14748,N_14709);
or UO_101 (O_101,N_14558,N_14846);
or UO_102 (O_102,N_14662,N_14622);
and UO_103 (O_103,N_14283,N_14581);
nand UO_104 (O_104,N_14801,N_14749);
nand UO_105 (O_105,N_14870,N_14710);
or UO_106 (O_106,N_14300,N_14875);
and UO_107 (O_107,N_14392,N_14880);
and UO_108 (O_108,N_14617,N_14320);
nand UO_109 (O_109,N_14879,N_14461);
nand UO_110 (O_110,N_14495,N_14465);
nand UO_111 (O_111,N_14505,N_14551);
nand UO_112 (O_112,N_14999,N_14691);
xnor UO_113 (O_113,N_14778,N_14706);
nand UO_114 (O_114,N_14990,N_14878);
xnor UO_115 (O_115,N_14938,N_14892);
xor UO_116 (O_116,N_14537,N_14396);
nor UO_117 (O_117,N_14479,N_14825);
nor UO_118 (O_118,N_14306,N_14760);
nor UO_119 (O_119,N_14786,N_14295);
and UO_120 (O_120,N_14933,N_14831);
nor UO_121 (O_121,N_14475,N_14732);
and UO_122 (O_122,N_14862,N_14982);
xnor UO_123 (O_123,N_14275,N_14352);
nand UO_124 (O_124,N_14591,N_14343);
nor UO_125 (O_125,N_14974,N_14860);
xnor UO_126 (O_126,N_14315,N_14647);
nand UO_127 (O_127,N_14342,N_14487);
xor UO_128 (O_128,N_14420,N_14911);
nor UO_129 (O_129,N_14987,N_14564);
and UO_130 (O_130,N_14823,N_14268);
xor UO_131 (O_131,N_14939,N_14333);
xor UO_132 (O_132,N_14969,N_14646);
xnor UO_133 (O_133,N_14486,N_14745);
nor UO_134 (O_134,N_14731,N_14937);
nor UO_135 (O_135,N_14981,N_14484);
or UO_136 (O_136,N_14579,N_14282);
and UO_137 (O_137,N_14694,N_14369);
or UO_138 (O_138,N_14546,N_14814);
or UO_139 (O_139,N_14274,N_14735);
or UO_140 (O_140,N_14652,N_14578);
and UO_141 (O_141,N_14574,N_14330);
and UO_142 (O_142,N_14336,N_14251);
xnor UO_143 (O_143,N_14253,N_14254);
nand UO_144 (O_144,N_14686,N_14800);
or UO_145 (O_145,N_14829,N_14815);
nand UO_146 (O_146,N_14936,N_14810);
nor UO_147 (O_147,N_14522,N_14945);
nand UO_148 (O_148,N_14761,N_14366);
nand UO_149 (O_149,N_14571,N_14669);
and UO_150 (O_150,N_14597,N_14679);
and UO_151 (O_151,N_14430,N_14742);
xor UO_152 (O_152,N_14687,N_14273);
nor UO_153 (O_153,N_14777,N_14941);
nand UO_154 (O_154,N_14673,N_14575);
or UO_155 (O_155,N_14818,N_14541);
nand UO_156 (O_156,N_14605,N_14529);
or UO_157 (O_157,N_14292,N_14835);
nand UO_158 (O_158,N_14331,N_14885);
and UO_159 (O_159,N_14446,N_14954);
nand UO_160 (O_160,N_14840,N_14293);
or UO_161 (O_161,N_14701,N_14291);
xnor UO_162 (O_162,N_14913,N_14405);
nor UO_163 (O_163,N_14872,N_14418);
nor UO_164 (O_164,N_14783,N_14612);
nand UO_165 (O_165,N_14526,N_14695);
or UO_166 (O_166,N_14826,N_14278);
and UO_167 (O_167,N_14448,N_14950);
or UO_168 (O_168,N_14754,N_14511);
nor UO_169 (O_169,N_14925,N_14704);
or UO_170 (O_170,N_14501,N_14773);
and UO_171 (O_171,N_14271,N_14432);
or UO_172 (O_172,N_14470,N_14449);
nor UO_173 (O_173,N_14766,N_14688);
nor UO_174 (O_174,N_14966,N_14995);
or UO_175 (O_175,N_14607,N_14437);
nand UO_176 (O_176,N_14368,N_14423);
nor UO_177 (O_177,N_14410,N_14845);
or UO_178 (O_178,N_14797,N_14611);
nor UO_179 (O_179,N_14457,N_14318);
nand UO_180 (O_180,N_14534,N_14264);
or UO_181 (O_181,N_14518,N_14524);
xnor UO_182 (O_182,N_14289,N_14426);
or UO_183 (O_183,N_14757,N_14716);
xnor UO_184 (O_184,N_14932,N_14724);
nand UO_185 (O_185,N_14493,N_14277);
or UO_186 (O_186,N_14920,N_14952);
or UO_187 (O_187,N_14582,N_14468);
nand UO_188 (O_188,N_14490,N_14916);
xor UO_189 (O_189,N_14903,N_14341);
nor UO_190 (O_190,N_14959,N_14692);
nand UO_191 (O_191,N_14623,N_14586);
and UO_192 (O_192,N_14447,N_14288);
nand UO_193 (O_193,N_14796,N_14890);
xnor UO_194 (O_194,N_14477,N_14569);
or UO_195 (O_195,N_14559,N_14976);
nand UO_196 (O_196,N_14259,N_14620);
nand UO_197 (O_197,N_14528,N_14907);
xor UO_198 (O_198,N_14712,N_14270);
nand UO_199 (O_199,N_14970,N_14307);
nor UO_200 (O_200,N_14837,N_14819);
nand UO_201 (O_201,N_14836,N_14374);
xnor UO_202 (O_202,N_14891,N_14398);
or UO_203 (O_203,N_14463,N_14824);
xor UO_204 (O_204,N_14648,N_14523);
and UO_205 (O_205,N_14940,N_14804);
nor UO_206 (O_206,N_14639,N_14852);
or UO_207 (O_207,N_14958,N_14723);
or UO_208 (O_208,N_14794,N_14764);
nor UO_209 (O_209,N_14863,N_14905);
nor UO_210 (O_210,N_14311,N_14853);
nor UO_211 (O_211,N_14409,N_14497);
nand UO_212 (O_212,N_14467,N_14504);
or UO_213 (O_213,N_14883,N_14377);
xor UO_214 (O_214,N_14616,N_14855);
and UO_215 (O_215,N_14641,N_14690);
nand UO_216 (O_216,N_14968,N_14284);
or UO_217 (O_217,N_14553,N_14888);
nor UO_218 (O_218,N_14889,N_14427);
nand UO_219 (O_219,N_14848,N_14910);
nor UO_220 (O_220,N_14603,N_14567);
nand UO_221 (O_221,N_14988,N_14592);
or UO_222 (O_222,N_14266,N_14896);
xnor UO_223 (O_223,N_14759,N_14476);
nand UO_224 (O_224,N_14464,N_14556);
or UO_225 (O_225,N_14971,N_14536);
xor UO_226 (O_226,N_14626,N_14828);
or UO_227 (O_227,N_14951,N_14587);
or UO_228 (O_228,N_14628,N_14304);
and UO_229 (O_229,N_14657,N_14645);
nand UO_230 (O_230,N_14733,N_14901);
nand UO_231 (O_231,N_14272,N_14827);
xnor UO_232 (O_232,N_14820,N_14294);
and UO_233 (O_233,N_14728,N_14682);
nor UO_234 (O_234,N_14643,N_14344);
nor UO_235 (O_235,N_14651,N_14290);
nor UO_236 (O_236,N_14545,N_14280);
nor UO_237 (O_237,N_14576,N_14817);
and UO_238 (O_238,N_14312,N_14514);
and UO_239 (O_239,N_14714,N_14594);
nand UO_240 (O_240,N_14795,N_14421);
xnor UO_241 (O_241,N_14562,N_14350);
nor UO_242 (O_242,N_14805,N_14734);
and UO_243 (O_243,N_14621,N_14655);
or UO_244 (O_244,N_14887,N_14472);
and UO_245 (O_245,N_14371,N_14434);
and UO_246 (O_246,N_14517,N_14483);
xnor UO_247 (O_247,N_14632,N_14510);
nand UO_248 (O_248,N_14685,N_14781);
xor UO_249 (O_249,N_14765,N_14598);
xnor UO_250 (O_250,N_14269,N_14401);
nand UO_251 (O_251,N_14593,N_14918);
and UO_252 (O_252,N_14843,N_14717);
and UO_253 (O_253,N_14725,N_14986);
nor UO_254 (O_254,N_14298,N_14250);
nor UO_255 (O_255,N_14462,N_14339);
nor UO_256 (O_256,N_14895,N_14263);
and UO_257 (O_257,N_14696,N_14496);
and UO_258 (O_258,N_14549,N_14744);
and UO_259 (O_259,N_14653,N_14555);
nor UO_260 (O_260,N_14873,N_14543);
nor UO_261 (O_261,N_14661,N_14413);
nand UO_262 (O_262,N_14337,N_14351);
nor UO_263 (O_263,N_14365,N_14739);
and UO_264 (O_264,N_14527,N_14600);
nand UO_265 (O_265,N_14672,N_14321);
nor UO_266 (O_266,N_14992,N_14741);
nand UO_267 (O_267,N_14525,N_14601);
and UO_268 (O_268,N_14967,N_14806);
and UO_269 (O_269,N_14730,N_14698);
xnor UO_270 (O_270,N_14747,N_14458);
or UO_271 (O_271,N_14700,N_14750);
and UO_272 (O_272,N_14542,N_14412);
and UO_273 (O_273,N_14323,N_14919);
nor UO_274 (O_274,N_14566,N_14512);
nand UO_275 (O_275,N_14906,N_14984);
nor UO_276 (O_276,N_14914,N_14606);
nand UO_277 (O_277,N_14613,N_14538);
or UO_278 (O_278,N_14400,N_14485);
nor UO_279 (O_279,N_14630,N_14711);
or UO_280 (O_280,N_14675,N_14385);
and UO_281 (O_281,N_14327,N_14898);
xor UO_282 (O_282,N_14577,N_14847);
nor UO_283 (O_283,N_14329,N_14790);
nor UO_284 (O_284,N_14839,N_14834);
xnor UO_285 (O_285,N_14314,N_14346);
nand UO_286 (O_286,N_14676,N_14509);
or UO_287 (O_287,N_14634,N_14372);
xnor UO_288 (O_288,N_14882,N_14494);
or UO_289 (O_289,N_14381,N_14816);
and UO_290 (O_290,N_14859,N_14474);
nor UO_291 (O_291,N_14397,N_14993);
and UO_292 (O_292,N_14636,N_14532);
nor UO_293 (O_293,N_14857,N_14489);
nor UO_294 (O_294,N_14317,N_14414);
xnor UO_295 (O_295,N_14874,N_14416);
nor UO_296 (O_296,N_14743,N_14642);
and UO_297 (O_297,N_14965,N_14670);
xor UO_298 (O_298,N_14719,N_14963);
xor UO_299 (O_299,N_14955,N_14684);
and UO_300 (O_300,N_14585,N_14779);
nand UO_301 (O_301,N_14727,N_14391);
nand UO_302 (O_302,N_14948,N_14680);
or UO_303 (O_303,N_14991,N_14614);
xnor UO_304 (O_304,N_14960,N_14539);
nand UO_305 (O_305,N_14402,N_14943);
or UO_306 (O_306,N_14989,N_14893);
or UO_307 (O_307,N_14443,N_14540);
nor UO_308 (O_308,N_14438,N_14756);
nor UO_309 (O_309,N_14580,N_14565);
xnor UO_310 (O_310,N_14977,N_14316);
xnor UO_311 (O_311,N_14455,N_14356);
xor UO_312 (O_312,N_14751,N_14980);
xor UO_313 (O_313,N_14640,N_14469);
xor UO_314 (O_314,N_14649,N_14364);
xor UO_315 (O_315,N_14908,N_14348);
nor UO_316 (O_316,N_14715,N_14929);
nor UO_317 (O_317,N_14319,N_14595);
nand UO_318 (O_318,N_14713,N_14707);
or UO_319 (O_319,N_14930,N_14737);
and UO_320 (O_320,N_14386,N_14705);
nor UO_321 (O_321,N_14935,N_14471);
nand UO_322 (O_322,N_14326,N_14624);
nand UO_323 (O_323,N_14299,N_14768);
and UO_324 (O_324,N_14573,N_14799);
nand UO_325 (O_325,N_14767,N_14425);
nand UO_326 (O_326,N_14399,N_14502);
nor UO_327 (O_327,N_14629,N_14265);
nor UO_328 (O_328,N_14257,N_14500);
and UO_329 (O_329,N_14869,N_14258);
nor UO_330 (O_330,N_14362,N_14557);
xnor UO_331 (O_331,N_14946,N_14917);
or UO_332 (O_332,N_14973,N_14762);
nand UO_333 (O_333,N_14947,N_14451);
nor UO_334 (O_334,N_14923,N_14868);
and UO_335 (O_335,N_14548,N_14900);
nor UO_336 (O_336,N_14588,N_14975);
and UO_337 (O_337,N_14871,N_14608);
and UO_338 (O_338,N_14436,N_14560);
xor UO_339 (O_339,N_14533,N_14956);
xnor UO_340 (O_340,N_14492,N_14788);
xnor UO_341 (O_341,N_14583,N_14830);
nor UO_342 (O_342,N_14453,N_14433);
xnor UO_343 (O_343,N_14660,N_14838);
and UO_344 (O_344,N_14347,N_14618);
or UO_345 (O_345,N_14570,N_14922);
nand UO_346 (O_346,N_14807,N_14353);
and UO_347 (O_347,N_14654,N_14736);
xnor UO_348 (O_348,N_14403,N_14375);
nor UO_349 (O_349,N_14261,N_14785);
nor UO_350 (O_350,N_14445,N_14997);
nand UO_351 (O_351,N_14904,N_14693);
nor UO_352 (O_352,N_14949,N_14408);
nor UO_353 (O_353,N_14345,N_14296);
and UO_354 (O_354,N_14780,N_14876);
and UO_355 (O_355,N_14697,N_14442);
xnor UO_356 (O_356,N_14388,N_14281);
or UO_357 (O_357,N_14758,N_14544);
and UO_358 (O_358,N_14389,N_14782);
and UO_359 (O_359,N_14803,N_14998);
nor UO_360 (O_360,N_14488,N_14625);
or UO_361 (O_361,N_14516,N_14429);
and UO_362 (O_362,N_14638,N_14934);
nor UO_363 (O_363,N_14899,N_14813);
or UO_364 (O_364,N_14792,N_14821);
nand UO_365 (O_365,N_14755,N_14849);
and UO_366 (O_366,N_14415,N_14729);
or UO_367 (O_367,N_14440,N_14452);
nor UO_368 (O_368,N_14521,N_14499);
or UO_369 (O_369,N_14851,N_14659);
or UO_370 (O_370,N_14864,N_14978);
or UO_371 (O_371,N_14772,N_14276);
or UO_372 (O_372,N_14677,N_14866);
and UO_373 (O_373,N_14424,N_14335);
nand UO_374 (O_374,N_14994,N_14332);
or UO_375 (O_375,N_14501,N_14252);
or UO_376 (O_376,N_14524,N_14636);
or UO_377 (O_377,N_14796,N_14765);
nor UO_378 (O_378,N_14761,N_14354);
and UO_379 (O_379,N_14429,N_14253);
nand UO_380 (O_380,N_14492,N_14603);
and UO_381 (O_381,N_14336,N_14569);
nand UO_382 (O_382,N_14457,N_14972);
or UO_383 (O_383,N_14879,N_14858);
or UO_384 (O_384,N_14820,N_14847);
nand UO_385 (O_385,N_14875,N_14908);
nor UO_386 (O_386,N_14735,N_14738);
and UO_387 (O_387,N_14576,N_14778);
and UO_388 (O_388,N_14620,N_14577);
or UO_389 (O_389,N_14570,N_14298);
nor UO_390 (O_390,N_14426,N_14556);
nor UO_391 (O_391,N_14676,N_14929);
and UO_392 (O_392,N_14678,N_14460);
nor UO_393 (O_393,N_14551,N_14915);
and UO_394 (O_394,N_14925,N_14727);
nor UO_395 (O_395,N_14614,N_14252);
nor UO_396 (O_396,N_14496,N_14493);
and UO_397 (O_397,N_14299,N_14898);
and UO_398 (O_398,N_14666,N_14724);
nor UO_399 (O_399,N_14568,N_14845);
or UO_400 (O_400,N_14484,N_14899);
or UO_401 (O_401,N_14870,N_14399);
xor UO_402 (O_402,N_14327,N_14926);
nand UO_403 (O_403,N_14903,N_14460);
or UO_404 (O_404,N_14980,N_14776);
nand UO_405 (O_405,N_14373,N_14456);
or UO_406 (O_406,N_14313,N_14263);
or UO_407 (O_407,N_14482,N_14833);
xnor UO_408 (O_408,N_14282,N_14917);
xnor UO_409 (O_409,N_14753,N_14653);
and UO_410 (O_410,N_14961,N_14734);
nand UO_411 (O_411,N_14562,N_14459);
and UO_412 (O_412,N_14350,N_14346);
and UO_413 (O_413,N_14820,N_14737);
and UO_414 (O_414,N_14388,N_14870);
xnor UO_415 (O_415,N_14758,N_14268);
or UO_416 (O_416,N_14812,N_14464);
and UO_417 (O_417,N_14414,N_14726);
nor UO_418 (O_418,N_14882,N_14346);
and UO_419 (O_419,N_14656,N_14279);
and UO_420 (O_420,N_14647,N_14253);
and UO_421 (O_421,N_14849,N_14393);
nand UO_422 (O_422,N_14874,N_14730);
and UO_423 (O_423,N_14955,N_14857);
xor UO_424 (O_424,N_14317,N_14895);
xor UO_425 (O_425,N_14795,N_14267);
xnor UO_426 (O_426,N_14550,N_14487);
xnor UO_427 (O_427,N_14893,N_14377);
and UO_428 (O_428,N_14540,N_14278);
or UO_429 (O_429,N_14264,N_14731);
and UO_430 (O_430,N_14877,N_14283);
xnor UO_431 (O_431,N_14278,N_14892);
and UO_432 (O_432,N_14982,N_14359);
and UO_433 (O_433,N_14410,N_14684);
xor UO_434 (O_434,N_14587,N_14366);
or UO_435 (O_435,N_14368,N_14930);
xor UO_436 (O_436,N_14916,N_14924);
nand UO_437 (O_437,N_14733,N_14774);
or UO_438 (O_438,N_14737,N_14445);
nor UO_439 (O_439,N_14573,N_14361);
nor UO_440 (O_440,N_14411,N_14290);
xnor UO_441 (O_441,N_14469,N_14523);
or UO_442 (O_442,N_14516,N_14994);
and UO_443 (O_443,N_14769,N_14537);
or UO_444 (O_444,N_14955,N_14540);
xnor UO_445 (O_445,N_14270,N_14833);
or UO_446 (O_446,N_14488,N_14465);
nor UO_447 (O_447,N_14524,N_14349);
or UO_448 (O_448,N_14505,N_14398);
xnor UO_449 (O_449,N_14797,N_14501);
nand UO_450 (O_450,N_14435,N_14451);
and UO_451 (O_451,N_14619,N_14793);
or UO_452 (O_452,N_14518,N_14997);
xor UO_453 (O_453,N_14302,N_14751);
nor UO_454 (O_454,N_14958,N_14387);
nor UO_455 (O_455,N_14480,N_14644);
nor UO_456 (O_456,N_14932,N_14878);
nor UO_457 (O_457,N_14695,N_14394);
xnor UO_458 (O_458,N_14958,N_14855);
nor UO_459 (O_459,N_14418,N_14685);
nand UO_460 (O_460,N_14549,N_14678);
and UO_461 (O_461,N_14943,N_14611);
nand UO_462 (O_462,N_14929,N_14862);
nor UO_463 (O_463,N_14518,N_14471);
and UO_464 (O_464,N_14519,N_14325);
and UO_465 (O_465,N_14882,N_14359);
and UO_466 (O_466,N_14600,N_14627);
nor UO_467 (O_467,N_14772,N_14472);
or UO_468 (O_468,N_14950,N_14659);
xnor UO_469 (O_469,N_14769,N_14856);
nand UO_470 (O_470,N_14575,N_14413);
and UO_471 (O_471,N_14925,N_14658);
and UO_472 (O_472,N_14913,N_14250);
xor UO_473 (O_473,N_14610,N_14563);
xnor UO_474 (O_474,N_14775,N_14302);
xnor UO_475 (O_475,N_14312,N_14638);
or UO_476 (O_476,N_14824,N_14404);
nand UO_477 (O_477,N_14511,N_14824);
or UO_478 (O_478,N_14393,N_14458);
or UO_479 (O_479,N_14484,N_14580);
xnor UO_480 (O_480,N_14802,N_14787);
or UO_481 (O_481,N_14302,N_14477);
or UO_482 (O_482,N_14448,N_14778);
xnor UO_483 (O_483,N_14319,N_14724);
xnor UO_484 (O_484,N_14302,N_14271);
nand UO_485 (O_485,N_14852,N_14354);
and UO_486 (O_486,N_14771,N_14360);
nand UO_487 (O_487,N_14617,N_14458);
and UO_488 (O_488,N_14394,N_14745);
and UO_489 (O_489,N_14624,N_14253);
xnor UO_490 (O_490,N_14391,N_14435);
nor UO_491 (O_491,N_14418,N_14903);
xor UO_492 (O_492,N_14770,N_14936);
nand UO_493 (O_493,N_14971,N_14811);
or UO_494 (O_494,N_14758,N_14702);
nand UO_495 (O_495,N_14741,N_14753);
or UO_496 (O_496,N_14402,N_14749);
nor UO_497 (O_497,N_14969,N_14958);
nand UO_498 (O_498,N_14581,N_14893);
or UO_499 (O_499,N_14429,N_14369);
or UO_500 (O_500,N_14319,N_14661);
nand UO_501 (O_501,N_14265,N_14267);
nand UO_502 (O_502,N_14611,N_14522);
or UO_503 (O_503,N_14826,N_14823);
nand UO_504 (O_504,N_14888,N_14785);
nor UO_505 (O_505,N_14504,N_14379);
or UO_506 (O_506,N_14656,N_14972);
nand UO_507 (O_507,N_14843,N_14649);
or UO_508 (O_508,N_14402,N_14973);
nor UO_509 (O_509,N_14485,N_14398);
or UO_510 (O_510,N_14465,N_14288);
nand UO_511 (O_511,N_14556,N_14620);
xor UO_512 (O_512,N_14662,N_14934);
or UO_513 (O_513,N_14288,N_14581);
xor UO_514 (O_514,N_14342,N_14473);
or UO_515 (O_515,N_14648,N_14388);
or UO_516 (O_516,N_14402,N_14925);
and UO_517 (O_517,N_14453,N_14458);
nand UO_518 (O_518,N_14892,N_14457);
or UO_519 (O_519,N_14418,N_14434);
and UO_520 (O_520,N_14557,N_14805);
or UO_521 (O_521,N_14741,N_14852);
nand UO_522 (O_522,N_14698,N_14680);
xnor UO_523 (O_523,N_14690,N_14636);
nand UO_524 (O_524,N_14787,N_14362);
nand UO_525 (O_525,N_14789,N_14397);
and UO_526 (O_526,N_14308,N_14457);
xor UO_527 (O_527,N_14435,N_14550);
nand UO_528 (O_528,N_14685,N_14484);
xnor UO_529 (O_529,N_14517,N_14421);
or UO_530 (O_530,N_14825,N_14679);
or UO_531 (O_531,N_14450,N_14337);
nor UO_532 (O_532,N_14406,N_14887);
or UO_533 (O_533,N_14250,N_14671);
nor UO_534 (O_534,N_14348,N_14932);
xor UO_535 (O_535,N_14557,N_14552);
xor UO_536 (O_536,N_14614,N_14870);
or UO_537 (O_537,N_14915,N_14817);
nand UO_538 (O_538,N_14416,N_14696);
or UO_539 (O_539,N_14333,N_14857);
nand UO_540 (O_540,N_14928,N_14285);
and UO_541 (O_541,N_14644,N_14780);
nor UO_542 (O_542,N_14404,N_14742);
nand UO_543 (O_543,N_14894,N_14250);
nor UO_544 (O_544,N_14488,N_14393);
nand UO_545 (O_545,N_14263,N_14793);
and UO_546 (O_546,N_14762,N_14856);
nor UO_547 (O_547,N_14643,N_14753);
xor UO_548 (O_548,N_14762,N_14774);
nand UO_549 (O_549,N_14853,N_14940);
nand UO_550 (O_550,N_14912,N_14614);
or UO_551 (O_551,N_14698,N_14747);
xnor UO_552 (O_552,N_14862,N_14934);
nor UO_553 (O_553,N_14695,N_14484);
nand UO_554 (O_554,N_14408,N_14647);
nor UO_555 (O_555,N_14447,N_14369);
nand UO_556 (O_556,N_14274,N_14934);
and UO_557 (O_557,N_14873,N_14707);
nand UO_558 (O_558,N_14260,N_14898);
xnor UO_559 (O_559,N_14772,N_14251);
xnor UO_560 (O_560,N_14361,N_14712);
nand UO_561 (O_561,N_14916,N_14303);
nand UO_562 (O_562,N_14961,N_14665);
nand UO_563 (O_563,N_14682,N_14291);
or UO_564 (O_564,N_14329,N_14321);
or UO_565 (O_565,N_14744,N_14932);
nor UO_566 (O_566,N_14884,N_14317);
xnor UO_567 (O_567,N_14879,N_14352);
and UO_568 (O_568,N_14503,N_14450);
nand UO_569 (O_569,N_14308,N_14634);
nor UO_570 (O_570,N_14277,N_14698);
nor UO_571 (O_571,N_14274,N_14506);
and UO_572 (O_572,N_14579,N_14804);
nor UO_573 (O_573,N_14270,N_14960);
or UO_574 (O_574,N_14538,N_14824);
xor UO_575 (O_575,N_14594,N_14624);
nand UO_576 (O_576,N_14331,N_14475);
or UO_577 (O_577,N_14499,N_14291);
nor UO_578 (O_578,N_14464,N_14871);
nor UO_579 (O_579,N_14271,N_14719);
nor UO_580 (O_580,N_14973,N_14867);
nor UO_581 (O_581,N_14585,N_14627);
nor UO_582 (O_582,N_14976,N_14338);
or UO_583 (O_583,N_14762,N_14915);
nor UO_584 (O_584,N_14831,N_14903);
or UO_585 (O_585,N_14530,N_14705);
xnor UO_586 (O_586,N_14972,N_14943);
nor UO_587 (O_587,N_14639,N_14333);
nand UO_588 (O_588,N_14551,N_14721);
nor UO_589 (O_589,N_14357,N_14296);
nand UO_590 (O_590,N_14278,N_14515);
and UO_591 (O_591,N_14910,N_14890);
xnor UO_592 (O_592,N_14833,N_14822);
xnor UO_593 (O_593,N_14649,N_14266);
and UO_594 (O_594,N_14845,N_14869);
xor UO_595 (O_595,N_14980,N_14392);
xnor UO_596 (O_596,N_14910,N_14579);
and UO_597 (O_597,N_14804,N_14616);
nand UO_598 (O_598,N_14349,N_14687);
or UO_599 (O_599,N_14290,N_14528);
xor UO_600 (O_600,N_14431,N_14954);
and UO_601 (O_601,N_14909,N_14948);
and UO_602 (O_602,N_14532,N_14692);
and UO_603 (O_603,N_14682,N_14388);
nor UO_604 (O_604,N_14687,N_14827);
nand UO_605 (O_605,N_14545,N_14829);
nand UO_606 (O_606,N_14527,N_14499);
nor UO_607 (O_607,N_14547,N_14454);
nand UO_608 (O_608,N_14937,N_14875);
or UO_609 (O_609,N_14733,N_14758);
or UO_610 (O_610,N_14665,N_14733);
xor UO_611 (O_611,N_14750,N_14978);
nand UO_612 (O_612,N_14663,N_14832);
nor UO_613 (O_613,N_14718,N_14551);
xnor UO_614 (O_614,N_14696,N_14759);
nor UO_615 (O_615,N_14705,N_14552);
nand UO_616 (O_616,N_14356,N_14508);
nand UO_617 (O_617,N_14775,N_14339);
nand UO_618 (O_618,N_14392,N_14488);
xnor UO_619 (O_619,N_14948,N_14899);
xor UO_620 (O_620,N_14737,N_14888);
nor UO_621 (O_621,N_14366,N_14611);
xnor UO_622 (O_622,N_14843,N_14741);
or UO_623 (O_623,N_14892,N_14379);
or UO_624 (O_624,N_14482,N_14264);
nor UO_625 (O_625,N_14890,N_14813);
nand UO_626 (O_626,N_14325,N_14846);
or UO_627 (O_627,N_14571,N_14885);
nor UO_628 (O_628,N_14979,N_14850);
and UO_629 (O_629,N_14582,N_14731);
xor UO_630 (O_630,N_14770,N_14823);
xor UO_631 (O_631,N_14633,N_14534);
nand UO_632 (O_632,N_14544,N_14701);
nand UO_633 (O_633,N_14833,N_14841);
xor UO_634 (O_634,N_14921,N_14953);
or UO_635 (O_635,N_14954,N_14919);
nand UO_636 (O_636,N_14760,N_14251);
and UO_637 (O_637,N_14839,N_14851);
xor UO_638 (O_638,N_14654,N_14413);
xor UO_639 (O_639,N_14792,N_14400);
xnor UO_640 (O_640,N_14744,N_14362);
and UO_641 (O_641,N_14947,N_14298);
and UO_642 (O_642,N_14839,N_14458);
xnor UO_643 (O_643,N_14921,N_14316);
xnor UO_644 (O_644,N_14557,N_14830);
or UO_645 (O_645,N_14768,N_14640);
nor UO_646 (O_646,N_14703,N_14312);
nand UO_647 (O_647,N_14397,N_14684);
xor UO_648 (O_648,N_14341,N_14714);
and UO_649 (O_649,N_14418,N_14504);
xnor UO_650 (O_650,N_14378,N_14300);
xnor UO_651 (O_651,N_14508,N_14765);
nor UO_652 (O_652,N_14385,N_14333);
and UO_653 (O_653,N_14918,N_14727);
and UO_654 (O_654,N_14582,N_14545);
and UO_655 (O_655,N_14367,N_14636);
nand UO_656 (O_656,N_14467,N_14527);
xor UO_657 (O_657,N_14354,N_14394);
or UO_658 (O_658,N_14949,N_14637);
or UO_659 (O_659,N_14300,N_14537);
nand UO_660 (O_660,N_14276,N_14375);
or UO_661 (O_661,N_14902,N_14709);
nor UO_662 (O_662,N_14424,N_14953);
or UO_663 (O_663,N_14567,N_14324);
xnor UO_664 (O_664,N_14697,N_14314);
xor UO_665 (O_665,N_14692,N_14931);
nand UO_666 (O_666,N_14504,N_14304);
nand UO_667 (O_667,N_14575,N_14615);
and UO_668 (O_668,N_14394,N_14541);
nand UO_669 (O_669,N_14285,N_14957);
xnor UO_670 (O_670,N_14264,N_14536);
nor UO_671 (O_671,N_14879,N_14932);
xor UO_672 (O_672,N_14621,N_14328);
nor UO_673 (O_673,N_14452,N_14325);
xor UO_674 (O_674,N_14388,N_14752);
nor UO_675 (O_675,N_14785,N_14384);
nand UO_676 (O_676,N_14604,N_14707);
or UO_677 (O_677,N_14800,N_14562);
or UO_678 (O_678,N_14917,N_14694);
nand UO_679 (O_679,N_14951,N_14799);
xnor UO_680 (O_680,N_14675,N_14324);
or UO_681 (O_681,N_14928,N_14807);
and UO_682 (O_682,N_14313,N_14360);
nand UO_683 (O_683,N_14995,N_14740);
or UO_684 (O_684,N_14676,N_14901);
or UO_685 (O_685,N_14298,N_14863);
xnor UO_686 (O_686,N_14612,N_14354);
nand UO_687 (O_687,N_14774,N_14434);
and UO_688 (O_688,N_14353,N_14511);
xor UO_689 (O_689,N_14449,N_14505);
nor UO_690 (O_690,N_14895,N_14497);
nor UO_691 (O_691,N_14447,N_14406);
nand UO_692 (O_692,N_14842,N_14259);
xnor UO_693 (O_693,N_14977,N_14840);
and UO_694 (O_694,N_14373,N_14881);
nor UO_695 (O_695,N_14975,N_14493);
xor UO_696 (O_696,N_14502,N_14293);
or UO_697 (O_697,N_14370,N_14481);
nor UO_698 (O_698,N_14770,N_14901);
xor UO_699 (O_699,N_14344,N_14391);
xnor UO_700 (O_700,N_14326,N_14764);
and UO_701 (O_701,N_14459,N_14498);
and UO_702 (O_702,N_14444,N_14453);
or UO_703 (O_703,N_14592,N_14846);
and UO_704 (O_704,N_14676,N_14990);
or UO_705 (O_705,N_14314,N_14384);
and UO_706 (O_706,N_14916,N_14318);
xnor UO_707 (O_707,N_14995,N_14873);
nor UO_708 (O_708,N_14981,N_14338);
nand UO_709 (O_709,N_14505,N_14441);
nor UO_710 (O_710,N_14429,N_14979);
or UO_711 (O_711,N_14973,N_14728);
and UO_712 (O_712,N_14621,N_14304);
and UO_713 (O_713,N_14796,N_14670);
xnor UO_714 (O_714,N_14697,N_14567);
nor UO_715 (O_715,N_14522,N_14880);
or UO_716 (O_716,N_14816,N_14658);
nor UO_717 (O_717,N_14441,N_14509);
nand UO_718 (O_718,N_14498,N_14469);
or UO_719 (O_719,N_14327,N_14260);
nor UO_720 (O_720,N_14918,N_14741);
nor UO_721 (O_721,N_14444,N_14456);
and UO_722 (O_722,N_14262,N_14922);
nand UO_723 (O_723,N_14644,N_14482);
nor UO_724 (O_724,N_14855,N_14739);
nor UO_725 (O_725,N_14568,N_14678);
nand UO_726 (O_726,N_14891,N_14950);
nor UO_727 (O_727,N_14366,N_14433);
nor UO_728 (O_728,N_14642,N_14643);
nand UO_729 (O_729,N_14747,N_14467);
or UO_730 (O_730,N_14528,N_14791);
and UO_731 (O_731,N_14783,N_14881);
and UO_732 (O_732,N_14593,N_14868);
and UO_733 (O_733,N_14554,N_14698);
xnor UO_734 (O_734,N_14439,N_14810);
and UO_735 (O_735,N_14918,N_14904);
nand UO_736 (O_736,N_14593,N_14434);
or UO_737 (O_737,N_14561,N_14737);
and UO_738 (O_738,N_14485,N_14663);
and UO_739 (O_739,N_14713,N_14289);
nand UO_740 (O_740,N_14565,N_14258);
nor UO_741 (O_741,N_14253,N_14957);
nand UO_742 (O_742,N_14391,N_14642);
and UO_743 (O_743,N_14988,N_14726);
nor UO_744 (O_744,N_14689,N_14996);
xnor UO_745 (O_745,N_14546,N_14644);
or UO_746 (O_746,N_14908,N_14784);
xor UO_747 (O_747,N_14697,N_14869);
and UO_748 (O_748,N_14739,N_14860);
nor UO_749 (O_749,N_14635,N_14646);
nand UO_750 (O_750,N_14896,N_14711);
nand UO_751 (O_751,N_14934,N_14250);
or UO_752 (O_752,N_14558,N_14269);
nand UO_753 (O_753,N_14758,N_14978);
or UO_754 (O_754,N_14970,N_14807);
xnor UO_755 (O_755,N_14705,N_14681);
xor UO_756 (O_756,N_14518,N_14652);
nor UO_757 (O_757,N_14819,N_14505);
nor UO_758 (O_758,N_14525,N_14463);
and UO_759 (O_759,N_14598,N_14489);
nand UO_760 (O_760,N_14603,N_14288);
nand UO_761 (O_761,N_14497,N_14730);
nor UO_762 (O_762,N_14380,N_14926);
nand UO_763 (O_763,N_14917,N_14891);
xnor UO_764 (O_764,N_14749,N_14944);
nand UO_765 (O_765,N_14792,N_14445);
and UO_766 (O_766,N_14282,N_14562);
or UO_767 (O_767,N_14774,N_14991);
or UO_768 (O_768,N_14254,N_14519);
or UO_769 (O_769,N_14545,N_14435);
nand UO_770 (O_770,N_14341,N_14271);
and UO_771 (O_771,N_14425,N_14871);
or UO_772 (O_772,N_14898,N_14292);
or UO_773 (O_773,N_14402,N_14420);
nor UO_774 (O_774,N_14649,N_14866);
and UO_775 (O_775,N_14731,N_14476);
and UO_776 (O_776,N_14271,N_14402);
and UO_777 (O_777,N_14388,N_14485);
or UO_778 (O_778,N_14975,N_14454);
nor UO_779 (O_779,N_14341,N_14883);
nor UO_780 (O_780,N_14546,N_14409);
xnor UO_781 (O_781,N_14649,N_14363);
or UO_782 (O_782,N_14940,N_14946);
nor UO_783 (O_783,N_14629,N_14517);
and UO_784 (O_784,N_14559,N_14409);
nand UO_785 (O_785,N_14698,N_14918);
or UO_786 (O_786,N_14951,N_14426);
or UO_787 (O_787,N_14599,N_14909);
or UO_788 (O_788,N_14945,N_14352);
nor UO_789 (O_789,N_14265,N_14474);
nor UO_790 (O_790,N_14841,N_14675);
or UO_791 (O_791,N_14925,N_14954);
and UO_792 (O_792,N_14711,N_14498);
or UO_793 (O_793,N_14310,N_14809);
or UO_794 (O_794,N_14720,N_14256);
or UO_795 (O_795,N_14927,N_14696);
nand UO_796 (O_796,N_14377,N_14988);
nand UO_797 (O_797,N_14389,N_14492);
or UO_798 (O_798,N_14401,N_14557);
nand UO_799 (O_799,N_14584,N_14666);
and UO_800 (O_800,N_14901,N_14751);
xnor UO_801 (O_801,N_14860,N_14284);
nand UO_802 (O_802,N_14347,N_14456);
and UO_803 (O_803,N_14540,N_14315);
nor UO_804 (O_804,N_14491,N_14567);
xnor UO_805 (O_805,N_14564,N_14405);
xor UO_806 (O_806,N_14654,N_14721);
and UO_807 (O_807,N_14899,N_14435);
nor UO_808 (O_808,N_14635,N_14686);
xnor UO_809 (O_809,N_14620,N_14507);
or UO_810 (O_810,N_14881,N_14968);
or UO_811 (O_811,N_14987,N_14615);
nor UO_812 (O_812,N_14833,N_14665);
and UO_813 (O_813,N_14356,N_14421);
nand UO_814 (O_814,N_14450,N_14702);
or UO_815 (O_815,N_14695,N_14848);
and UO_816 (O_816,N_14540,N_14581);
or UO_817 (O_817,N_14337,N_14478);
nand UO_818 (O_818,N_14790,N_14745);
nor UO_819 (O_819,N_14561,N_14858);
nor UO_820 (O_820,N_14857,N_14913);
and UO_821 (O_821,N_14436,N_14993);
nand UO_822 (O_822,N_14815,N_14353);
and UO_823 (O_823,N_14581,N_14832);
nor UO_824 (O_824,N_14632,N_14626);
nand UO_825 (O_825,N_14631,N_14544);
or UO_826 (O_826,N_14444,N_14337);
xor UO_827 (O_827,N_14268,N_14496);
nor UO_828 (O_828,N_14869,N_14565);
nor UO_829 (O_829,N_14512,N_14599);
and UO_830 (O_830,N_14900,N_14793);
nor UO_831 (O_831,N_14376,N_14881);
or UO_832 (O_832,N_14343,N_14874);
nand UO_833 (O_833,N_14778,N_14377);
xnor UO_834 (O_834,N_14307,N_14890);
and UO_835 (O_835,N_14316,N_14404);
xor UO_836 (O_836,N_14356,N_14795);
and UO_837 (O_837,N_14420,N_14760);
nor UO_838 (O_838,N_14567,N_14693);
and UO_839 (O_839,N_14331,N_14449);
xnor UO_840 (O_840,N_14476,N_14372);
nor UO_841 (O_841,N_14398,N_14517);
nand UO_842 (O_842,N_14497,N_14595);
nand UO_843 (O_843,N_14620,N_14292);
nand UO_844 (O_844,N_14667,N_14349);
xnor UO_845 (O_845,N_14770,N_14540);
nor UO_846 (O_846,N_14974,N_14942);
nor UO_847 (O_847,N_14640,N_14741);
and UO_848 (O_848,N_14258,N_14817);
or UO_849 (O_849,N_14648,N_14799);
and UO_850 (O_850,N_14960,N_14993);
nand UO_851 (O_851,N_14957,N_14870);
and UO_852 (O_852,N_14703,N_14394);
or UO_853 (O_853,N_14822,N_14731);
nor UO_854 (O_854,N_14822,N_14279);
or UO_855 (O_855,N_14855,N_14743);
nand UO_856 (O_856,N_14473,N_14570);
and UO_857 (O_857,N_14454,N_14607);
xnor UO_858 (O_858,N_14426,N_14566);
nand UO_859 (O_859,N_14416,N_14780);
and UO_860 (O_860,N_14863,N_14467);
nor UO_861 (O_861,N_14588,N_14847);
or UO_862 (O_862,N_14680,N_14549);
nor UO_863 (O_863,N_14530,N_14646);
nand UO_864 (O_864,N_14871,N_14477);
nor UO_865 (O_865,N_14985,N_14910);
xnor UO_866 (O_866,N_14353,N_14716);
or UO_867 (O_867,N_14490,N_14250);
nor UO_868 (O_868,N_14590,N_14697);
nor UO_869 (O_869,N_14547,N_14854);
and UO_870 (O_870,N_14959,N_14803);
nor UO_871 (O_871,N_14382,N_14636);
or UO_872 (O_872,N_14704,N_14528);
or UO_873 (O_873,N_14335,N_14350);
nor UO_874 (O_874,N_14670,N_14306);
or UO_875 (O_875,N_14826,N_14922);
nand UO_876 (O_876,N_14355,N_14468);
or UO_877 (O_877,N_14481,N_14812);
and UO_878 (O_878,N_14932,N_14387);
nor UO_879 (O_879,N_14366,N_14763);
nor UO_880 (O_880,N_14577,N_14675);
xor UO_881 (O_881,N_14361,N_14721);
xnor UO_882 (O_882,N_14259,N_14434);
and UO_883 (O_883,N_14768,N_14796);
or UO_884 (O_884,N_14599,N_14800);
nor UO_885 (O_885,N_14862,N_14301);
nor UO_886 (O_886,N_14888,N_14364);
xnor UO_887 (O_887,N_14426,N_14682);
nor UO_888 (O_888,N_14525,N_14540);
and UO_889 (O_889,N_14322,N_14593);
and UO_890 (O_890,N_14921,N_14973);
xnor UO_891 (O_891,N_14772,N_14922);
and UO_892 (O_892,N_14468,N_14571);
nor UO_893 (O_893,N_14809,N_14491);
nand UO_894 (O_894,N_14735,N_14695);
nand UO_895 (O_895,N_14804,N_14442);
and UO_896 (O_896,N_14524,N_14643);
nor UO_897 (O_897,N_14250,N_14418);
nor UO_898 (O_898,N_14690,N_14740);
nor UO_899 (O_899,N_14746,N_14523);
xnor UO_900 (O_900,N_14787,N_14480);
nor UO_901 (O_901,N_14754,N_14617);
nand UO_902 (O_902,N_14421,N_14796);
xor UO_903 (O_903,N_14365,N_14656);
nand UO_904 (O_904,N_14876,N_14451);
xnor UO_905 (O_905,N_14861,N_14655);
or UO_906 (O_906,N_14413,N_14816);
nor UO_907 (O_907,N_14850,N_14803);
xnor UO_908 (O_908,N_14929,N_14347);
nor UO_909 (O_909,N_14939,N_14960);
nor UO_910 (O_910,N_14765,N_14480);
nor UO_911 (O_911,N_14671,N_14838);
nand UO_912 (O_912,N_14918,N_14358);
xor UO_913 (O_913,N_14349,N_14403);
nand UO_914 (O_914,N_14973,N_14852);
or UO_915 (O_915,N_14364,N_14546);
and UO_916 (O_916,N_14933,N_14854);
nand UO_917 (O_917,N_14912,N_14522);
or UO_918 (O_918,N_14434,N_14294);
xnor UO_919 (O_919,N_14352,N_14659);
and UO_920 (O_920,N_14791,N_14438);
or UO_921 (O_921,N_14636,N_14996);
xor UO_922 (O_922,N_14783,N_14851);
nor UO_923 (O_923,N_14708,N_14404);
xnor UO_924 (O_924,N_14406,N_14855);
or UO_925 (O_925,N_14544,N_14866);
xnor UO_926 (O_926,N_14397,N_14829);
xnor UO_927 (O_927,N_14975,N_14718);
nand UO_928 (O_928,N_14309,N_14487);
and UO_929 (O_929,N_14265,N_14791);
nor UO_930 (O_930,N_14880,N_14379);
nor UO_931 (O_931,N_14459,N_14813);
nor UO_932 (O_932,N_14700,N_14279);
xor UO_933 (O_933,N_14668,N_14917);
nand UO_934 (O_934,N_14452,N_14688);
or UO_935 (O_935,N_14791,N_14659);
or UO_936 (O_936,N_14407,N_14485);
and UO_937 (O_937,N_14966,N_14313);
and UO_938 (O_938,N_14663,N_14833);
and UO_939 (O_939,N_14489,N_14663);
nand UO_940 (O_940,N_14840,N_14861);
xnor UO_941 (O_941,N_14581,N_14392);
or UO_942 (O_942,N_14364,N_14942);
nor UO_943 (O_943,N_14858,N_14757);
and UO_944 (O_944,N_14486,N_14501);
and UO_945 (O_945,N_14276,N_14398);
nand UO_946 (O_946,N_14630,N_14923);
or UO_947 (O_947,N_14420,N_14741);
and UO_948 (O_948,N_14481,N_14383);
nor UO_949 (O_949,N_14477,N_14443);
or UO_950 (O_950,N_14663,N_14968);
and UO_951 (O_951,N_14789,N_14650);
nand UO_952 (O_952,N_14369,N_14903);
nor UO_953 (O_953,N_14646,N_14971);
nand UO_954 (O_954,N_14315,N_14801);
or UO_955 (O_955,N_14308,N_14469);
nand UO_956 (O_956,N_14622,N_14943);
nor UO_957 (O_957,N_14782,N_14327);
or UO_958 (O_958,N_14501,N_14627);
nor UO_959 (O_959,N_14616,N_14451);
and UO_960 (O_960,N_14254,N_14462);
and UO_961 (O_961,N_14588,N_14824);
nand UO_962 (O_962,N_14903,N_14635);
nand UO_963 (O_963,N_14558,N_14421);
and UO_964 (O_964,N_14852,N_14796);
nor UO_965 (O_965,N_14878,N_14510);
nand UO_966 (O_966,N_14701,N_14493);
or UO_967 (O_967,N_14322,N_14972);
xor UO_968 (O_968,N_14804,N_14505);
or UO_969 (O_969,N_14483,N_14532);
nor UO_970 (O_970,N_14441,N_14266);
or UO_971 (O_971,N_14299,N_14370);
xor UO_972 (O_972,N_14489,N_14789);
and UO_973 (O_973,N_14881,N_14552);
xnor UO_974 (O_974,N_14950,N_14500);
and UO_975 (O_975,N_14818,N_14503);
nand UO_976 (O_976,N_14933,N_14801);
nor UO_977 (O_977,N_14555,N_14947);
or UO_978 (O_978,N_14600,N_14808);
nor UO_979 (O_979,N_14682,N_14452);
nand UO_980 (O_980,N_14300,N_14251);
nor UO_981 (O_981,N_14393,N_14904);
nand UO_982 (O_982,N_14434,N_14255);
or UO_983 (O_983,N_14316,N_14343);
or UO_984 (O_984,N_14895,N_14844);
nand UO_985 (O_985,N_14661,N_14754);
nand UO_986 (O_986,N_14663,N_14424);
or UO_987 (O_987,N_14824,N_14769);
nor UO_988 (O_988,N_14490,N_14485);
nor UO_989 (O_989,N_14255,N_14754);
xnor UO_990 (O_990,N_14626,N_14471);
and UO_991 (O_991,N_14476,N_14725);
or UO_992 (O_992,N_14988,N_14253);
nor UO_993 (O_993,N_14916,N_14375);
or UO_994 (O_994,N_14617,N_14436);
nand UO_995 (O_995,N_14560,N_14635);
nand UO_996 (O_996,N_14875,N_14523);
and UO_997 (O_997,N_14612,N_14269);
nand UO_998 (O_998,N_14909,N_14944);
xnor UO_999 (O_999,N_14322,N_14490);
nand UO_1000 (O_1000,N_14654,N_14573);
nor UO_1001 (O_1001,N_14314,N_14711);
nand UO_1002 (O_1002,N_14708,N_14675);
xor UO_1003 (O_1003,N_14400,N_14791);
nor UO_1004 (O_1004,N_14354,N_14959);
and UO_1005 (O_1005,N_14391,N_14646);
xnor UO_1006 (O_1006,N_14383,N_14540);
or UO_1007 (O_1007,N_14708,N_14961);
or UO_1008 (O_1008,N_14480,N_14451);
nand UO_1009 (O_1009,N_14866,N_14553);
and UO_1010 (O_1010,N_14271,N_14487);
and UO_1011 (O_1011,N_14429,N_14820);
nand UO_1012 (O_1012,N_14666,N_14963);
and UO_1013 (O_1013,N_14587,N_14911);
xnor UO_1014 (O_1014,N_14606,N_14423);
nand UO_1015 (O_1015,N_14466,N_14827);
and UO_1016 (O_1016,N_14997,N_14649);
and UO_1017 (O_1017,N_14878,N_14646);
or UO_1018 (O_1018,N_14982,N_14736);
nand UO_1019 (O_1019,N_14945,N_14854);
nor UO_1020 (O_1020,N_14826,N_14474);
nand UO_1021 (O_1021,N_14415,N_14645);
nand UO_1022 (O_1022,N_14633,N_14310);
and UO_1023 (O_1023,N_14870,N_14453);
nor UO_1024 (O_1024,N_14533,N_14550);
or UO_1025 (O_1025,N_14442,N_14581);
nand UO_1026 (O_1026,N_14301,N_14310);
and UO_1027 (O_1027,N_14352,N_14547);
nor UO_1028 (O_1028,N_14897,N_14815);
nand UO_1029 (O_1029,N_14253,N_14946);
and UO_1030 (O_1030,N_14363,N_14568);
nor UO_1031 (O_1031,N_14437,N_14837);
xor UO_1032 (O_1032,N_14572,N_14740);
nor UO_1033 (O_1033,N_14774,N_14315);
nand UO_1034 (O_1034,N_14606,N_14342);
nor UO_1035 (O_1035,N_14297,N_14927);
or UO_1036 (O_1036,N_14911,N_14357);
xor UO_1037 (O_1037,N_14250,N_14459);
nor UO_1038 (O_1038,N_14821,N_14513);
or UO_1039 (O_1039,N_14860,N_14259);
or UO_1040 (O_1040,N_14522,N_14956);
and UO_1041 (O_1041,N_14801,N_14453);
and UO_1042 (O_1042,N_14900,N_14457);
or UO_1043 (O_1043,N_14736,N_14996);
xnor UO_1044 (O_1044,N_14992,N_14748);
or UO_1045 (O_1045,N_14602,N_14571);
nand UO_1046 (O_1046,N_14961,N_14412);
nor UO_1047 (O_1047,N_14700,N_14818);
xor UO_1048 (O_1048,N_14901,N_14314);
xnor UO_1049 (O_1049,N_14430,N_14762);
xnor UO_1050 (O_1050,N_14557,N_14443);
nor UO_1051 (O_1051,N_14799,N_14997);
nand UO_1052 (O_1052,N_14433,N_14692);
xnor UO_1053 (O_1053,N_14911,N_14693);
nand UO_1054 (O_1054,N_14425,N_14993);
xnor UO_1055 (O_1055,N_14786,N_14609);
and UO_1056 (O_1056,N_14803,N_14636);
nand UO_1057 (O_1057,N_14250,N_14644);
nor UO_1058 (O_1058,N_14479,N_14275);
xor UO_1059 (O_1059,N_14914,N_14529);
and UO_1060 (O_1060,N_14885,N_14493);
and UO_1061 (O_1061,N_14635,N_14518);
or UO_1062 (O_1062,N_14683,N_14429);
xor UO_1063 (O_1063,N_14442,N_14340);
and UO_1064 (O_1064,N_14882,N_14928);
nand UO_1065 (O_1065,N_14658,N_14694);
or UO_1066 (O_1066,N_14955,N_14522);
or UO_1067 (O_1067,N_14748,N_14708);
xnor UO_1068 (O_1068,N_14709,N_14473);
nor UO_1069 (O_1069,N_14331,N_14263);
nor UO_1070 (O_1070,N_14439,N_14443);
and UO_1071 (O_1071,N_14615,N_14695);
nand UO_1072 (O_1072,N_14416,N_14761);
or UO_1073 (O_1073,N_14697,N_14612);
xnor UO_1074 (O_1074,N_14288,N_14826);
xor UO_1075 (O_1075,N_14296,N_14905);
xnor UO_1076 (O_1076,N_14287,N_14737);
and UO_1077 (O_1077,N_14391,N_14871);
or UO_1078 (O_1078,N_14681,N_14381);
or UO_1079 (O_1079,N_14787,N_14784);
xnor UO_1080 (O_1080,N_14272,N_14707);
xor UO_1081 (O_1081,N_14642,N_14794);
or UO_1082 (O_1082,N_14529,N_14524);
nor UO_1083 (O_1083,N_14645,N_14848);
nor UO_1084 (O_1084,N_14720,N_14505);
and UO_1085 (O_1085,N_14348,N_14801);
nor UO_1086 (O_1086,N_14979,N_14866);
or UO_1087 (O_1087,N_14463,N_14424);
nand UO_1088 (O_1088,N_14900,N_14522);
and UO_1089 (O_1089,N_14627,N_14798);
xnor UO_1090 (O_1090,N_14410,N_14731);
nand UO_1091 (O_1091,N_14940,N_14733);
xnor UO_1092 (O_1092,N_14589,N_14934);
and UO_1093 (O_1093,N_14423,N_14431);
xnor UO_1094 (O_1094,N_14625,N_14336);
or UO_1095 (O_1095,N_14255,N_14771);
and UO_1096 (O_1096,N_14504,N_14724);
or UO_1097 (O_1097,N_14977,N_14464);
nand UO_1098 (O_1098,N_14381,N_14996);
and UO_1099 (O_1099,N_14873,N_14661);
nand UO_1100 (O_1100,N_14645,N_14833);
nand UO_1101 (O_1101,N_14889,N_14608);
nand UO_1102 (O_1102,N_14713,N_14441);
and UO_1103 (O_1103,N_14886,N_14629);
and UO_1104 (O_1104,N_14809,N_14843);
nand UO_1105 (O_1105,N_14425,N_14325);
nor UO_1106 (O_1106,N_14484,N_14508);
nor UO_1107 (O_1107,N_14270,N_14905);
and UO_1108 (O_1108,N_14274,N_14366);
and UO_1109 (O_1109,N_14534,N_14453);
nor UO_1110 (O_1110,N_14986,N_14594);
or UO_1111 (O_1111,N_14986,N_14904);
nor UO_1112 (O_1112,N_14293,N_14559);
or UO_1113 (O_1113,N_14673,N_14556);
and UO_1114 (O_1114,N_14423,N_14706);
nor UO_1115 (O_1115,N_14789,N_14864);
and UO_1116 (O_1116,N_14957,N_14667);
and UO_1117 (O_1117,N_14886,N_14594);
or UO_1118 (O_1118,N_14479,N_14578);
nor UO_1119 (O_1119,N_14987,N_14538);
nor UO_1120 (O_1120,N_14948,N_14625);
xnor UO_1121 (O_1121,N_14648,N_14840);
nor UO_1122 (O_1122,N_14773,N_14549);
nand UO_1123 (O_1123,N_14441,N_14854);
and UO_1124 (O_1124,N_14376,N_14276);
xor UO_1125 (O_1125,N_14705,N_14767);
nand UO_1126 (O_1126,N_14617,N_14582);
nor UO_1127 (O_1127,N_14573,N_14349);
nand UO_1128 (O_1128,N_14517,N_14813);
xor UO_1129 (O_1129,N_14535,N_14325);
or UO_1130 (O_1130,N_14873,N_14478);
nand UO_1131 (O_1131,N_14817,N_14731);
nand UO_1132 (O_1132,N_14951,N_14316);
nand UO_1133 (O_1133,N_14941,N_14415);
or UO_1134 (O_1134,N_14386,N_14761);
or UO_1135 (O_1135,N_14869,N_14883);
nand UO_1136 (O_1136,N_14955,N_14870);
or UO_1137 (O_1137,N_14669,N_14873);
nor UO_1138 (O_1138,N_14907,N_14627);
or UO_1139 (O_1139,N_14706,N_14879);
or UO_1140 (O_1140,N_14411,N_14273);
xnor UO_1141 (O_1141,N_14551,N_14555);
and UO_1142 (O_1142,N_14594,N_14430);
nor UO_1143 (O_1143,N_14792,N_14959);
nor UO_1144 (O_1144,N_14718,N_14468);
nand UO_1145 (O_1145,N_14739,N_14492);
and UO_1146 (O_1146,N_14572,N_14835);
or UO_1147 (O_1147,N_14608,N_14868);
nor UO_1148 (O_1148,N_14503,N_14251);
nand UO_1149 (O_1149,N_14982,N_14568);
nor UO_1150 (O_1150,N_14620,N_14655);
nor UO_1151 (O_1151,N_14491,N_14678);
and UO_1152 (O_1152,N_14943,N_14841);
nor UO_1153 (O_1153,N_14540,N_14892);
or UO_1154 (O_1154,N_14432,N_14740);
or UO_1155 (O_1155,N_14970,N_14293);
xnor UO_1156 (O_1156,N_14537,N_14420);
xnor UO_1157 (O_1157,N_14584,N_14346);
xor UO_1158 (O_1158,N_14462,N_14605);
xor UO_1159 (O_1159,N_14454,N_14472);
xor UO_1160 (O_1160,N_14871,N_14624);
and UO_1161 (O_1161,N_14473,N_14566);
xnor UO_1162 (O_1162,N_14876,N_14764);
and UO_1163 (O_1163,N_14458,N_14873);
xnor UO_1164 (O_1164,N_14659,N_14433);
nand UO_1165 (O_1165,N_14758,N_14717);
nor UO_1166 (O_1166,N_14952,N_14635);
or UO_1167 (O_1167,N_14388,N_14478);
and UO_1168 (O_1168,N_14801,N_14508);
nor UO_1169 (O_1169,N_14500,N_14666);
or UO_1170 (O_1170,N_14533,N_14783);
and UO_1171 (O_1171,N_14941,N_14462);
xor UO_1172 (O_1172,N_14436,N_14275);
and UO_1173 (O_1173,N_14918,N_14980);
nand UO_1174 (O_1174,N_14653,N_14793);
and UO_1175 (O_1175,N_14290,N_14274);
nand UO_1176 (O_1176,N_14337,N_14622);
or UO_1177 (O_1177,N_14479,N_14796);
nand UO_1178 (O_1178,N_14838,N_14376);
nand UO_1179 (O_1179,N_14562,N_14811);
nand UO_1180 (O_1180,N_14414,N_14920);
nand UO_1181 (O_1181,N_14648,N_14711);
or UO_1182 (O_1182,N_14937,N_14433);
nor UO_1183 (O_1183,N_14710,N_14718);
xor UO_1184 (O_1184,N_14459,N_14576);
nand UO_1185 (O_1185,N_14799,N_14738);
nor UO_1186 (O_1186,N_14478,N_14786);
nor UO_1187 (O_1187,N_14700,N_14574);
xnor UO_1188 (O_1188,N_14798,N_14957);
or UO_1189 (O_1189,N_14738,N_14629);
and UO_1190 (O_1190,N_14998,N_14719);
nand UO_1191 (O_1191,N_14588,N_14458);
nand UO_1192 (O_1192,N_14261,N_14615);
or UO_1193 (O_1193,N_14623,N_14417);
and UO_1194 (O_1194,N_14341,N_14482);
nor UO_1195 (O_1195,N_14424,N_14871);
or UO_1196 (O_1196,N_14757,N_14551);
nor UO_1197 (O_1197,N_14437,N_14585);
xnor UO_1198 (O_1198,N_14402,N_14472);
nand UO_1199 (O_1199,N_14380,N_14556);
or UO_1200 (O_1200,N_14900,N_14914);
nor UO_1201 (O_1201,N_14612,N_14467);
nand UO_1202 (O_1202,N_14744,N_14660);
and UO_1203 (O_1203,N_14778,N_14633);
xor UO_1204 (O_1204,N_14351,N_14471);
and UO_1205 (O_1205,N_14387,N_14875);
nor UO_1206 (O_1206,N_14574,N_14379);
xor UO_1207 (O_1207,N_14284,N_14530);
nand UO_1208 (O_1208,N_14356,N_14494);
nor UO_1209 (O_1209,N_14255,N_14698);
nor UO_1210 (O_1210,N_14734,N_14494);
nor UO_1211 (O_1211,N_14928,N_14343);
and UO_1212 (O_1212,N_14387,N_14625);
nor UO_1213 (O_1213,N_14507,N_14994);
nand UO_1214 (O_1214,N_14789,N_14524);
and UO_1215 (O_1215,N_14337,N_14505);
or UO_1216 (O_1216,N_14515,N_14904);
and UO_1217 (O_1217,N_14913,N_14502);
or UO_1218 (O_1218,N_14448,N_14687);
or UO_1219 (O_1219,N_14687,N_14876);
and UO_1220 (O_1220,N_14298,N_14957);
and UO_1221 (O_1221,N_14497,N_14909);
and UO_1222 (O_1222,N_14904,N_14437);
xor UO_1223 (O_1223,N_14417,N_14937);
and UO_1224 (O_1224,N_14563,N_14423);
nor UO_1225 (O_1225,N_14941,N_14749);
and UO_1226 (O_1226,N_14556,N_14345);
nor UO_1227 (O_1227,N_14904,N_14583);
nand UO_1228 (O_1228,N_14570,N_14491);
xor UO_1229 (O_1229,N_14840,N_14536);
nand UO_1230 (O_1230,N_14841,N_14820);
xor UO_1231 (O_1231,N_14913,N_14524);
nand UO_1232 (O_1232,N_14961,N_14504);
xor UO_1233 (O_1233,N_14446,N_14958);
and UO_1234 (O_1234,N_14408,N_14279);
and UO_1235 (O_1235,N_14586,N_14938);
nor UO_1236 (O_1236,N_14375,N_14397);
or UO_1237 (O_1237,N_14656,N_14691);
xor UO_1238 (O_1238,N_14589,N_14968);
and UO_1239 (O_1239,N_14581,N_14712);
and UO_1240 (O_1240,N_14950,N_14727);
or UO_1241 (O_1241,N_14769,N_14658);
or UO_1242 (O_1242,N_14528,N_14984);
and UO_1243 (O_1243,N_14548,N_14788);
nor UO_1244 (O_1244,N_14362,N_14368);
or UO_1245 (O_1245,N_14279,N_14740);
xor UO_1246 (O_1246,N_14797,N_14826);
xor UO_1247 (O_1247,N_14874,N_14275);
nor UO_1248 (O_1248,N_14451,N_14702);
nor UO_1249 (O_1249,N_14735,N_14797);
xor UO_1250 (O_1250,N_14283,N_14747);
nand UO_1251 (O_1251,N_14828,N_14907);
or UO_1252 (O_1252,N_14926,N_14347);
xnor UO_1253 (O_1253,N_14960,N_14353);
nor UO_1254 (O_1254,N_14467,N_14517);
and UO_1255 (O_1255,N_14697,N_14905);
and UO_1256 (O_1256,N_14685,N_14429);
or UO_1257 (O_1257,N_14272,N_14603);
or UO_1258 (O_1258,N_14873,N_14974);
nor UO_1259 (O_1259,N_14684,N_14959);
nor UO_1260 (O_1260,N_14515,N_14621);
nand UO_1261 (O_1261,N_14775,N_14653);
or UO_1262 (O_1262,N_14659,N_14668);
xnor UO_1263 (O_1263,N_14695,N_14961);
nand UO_1264 (O_1264,N_14520,N_14949);
and UO_1265 (O_1265,N_14498,N_14564);
nor UO_1266 (O_1266,N_14462,N_14609);
or UO_1267 (O_1267,N_14516,N_14828);
and UO_1268 (O_1268,N_14530,N_14428);
nand UO_1269 (O_1269,N_14376,N_14446);
and UO_1270 (O_1270,N_14637,N_14847);
xor UO_1271 (O_1271,N_14771,N_14997);
xor UO_1272 (O_1272,N_14263,N_14350);
or UO_1273 (O_1273,N_14559,N_14970);
nor UO_1274 (O_1274,N_14783,N_14762);
xnor UO_1275 (O_1275,N_14376,N_14425);
or UO_1276 (O_1276,N_14847,N_14409);
or UO_1277 (O_1277,N_14613,N_14738);
or UO_1278 (O_1278,N_14852,N_14309);
nand UO_1279 (O_1279,N_14431,N_14454);
and UO_1280 (O_1280,N_14866,N_14343);
nand UO_1281 (O_1281,N_14576,N_14426);
nor UO_1282 (O_1282,N_14256,N_14329);
or UO_1283 (O_1283,N_14351,N_14701);
nand UO_1284 (O_1284,N_14703,N_14922);
nor UO_1285 (O_1285,N_14662,N_14676);
xor UO_1286 (O_1286,N_14658,N_14625);
or UO_1287 (O_1287,N_14306,N_14445);
nor UO_1288 (O_1288,N_14784,N_14578);
nor UO_1289 (O_1289,N_14811,N_14571);
nor UO_1290 (O_1290,N_14726,N_14671);
and UO_1291 (O_1291,N_14753,N_14340);
and UO_1292 (O_1292,N_14796,N_14594);
nor UO_1293 (O_1293,N_14623,N_14576);
nand UO_1294 (O_1294,N_14623,N_14532);
xnor UO_1295 (O_1295,N_14726,N_14619);
or UO_1296 (O_1296,N_14665,N_14805);
and UO_1297 (O_1297,N_14901,N_14260);
nor UO_1298 (O_1298,N_14588,N_14439);
and UO_1299 (O_1299,N_14788,N_14880);
or UO_1300 (O_1300,N_14829,N_14620);
or UO_1301 (O_1301,N_14995,N_14827);
nor UO_1302 (O_1302,N_14729,N_14632);
nand UO_1303 (O_1303,N_14620,N_14711);
xnor UO_1304 (O_1304,N_14466,N_14862);
xor UO_1305 (O_1305,N_14372,N_14482);
nor UO_1306 (O_1306,N_14390,N_14981);
or UO_1307 (O_1307,N_14734,N_14648);
nand UO_1308 (O_1308,N_14850,N_14729);
nand UO_1309 (O_1309,N_14657,N_14478);
or UO_1310 (O_1310,N_14673,N_14257);
nand UO_1311 (O_1311,N_14394,N_14683);
or UO_1312 (O_1312,N_14801,N_14520);
and UO_1313 (O_1313,N_14994,N_14765);
nor UO_1314 (O_1314,N_14577,N_14967);
or UO_1315 (O_1315,N_14324,N_14571);
or UO_1316 (O_1316,N_14519,N_14477);
nor UO_1317 (O_1317,N_14872,N_14877);
and UO_1318 (O_1318,N_14856,N_14630);
or UO_1319 (O_1319,N_14598,N_14672);
nand UO_1320 (O_1320,N_14401,N_14391);
or UO_1321 (O_1321,N_14916,N_14465);
and UO_1322 (O_1322,N_14837,N_14672);
xnor UO_1323 (O_1323,N_14776,N_14357);
or UO_1324 (O_1324,N_14358,N_14488);
or UO_1325 (O_1325,N_14806,N_14860);
xnor UO_1326 (O_1326,N_14400,N_14863);
or UO_1327 (O_1327,N_14284,N_14254);
xor UO_1328 (O_1328,N_14409,N_14374);
xor UO_1329 (O_1329,N_14531,N_14320);
nand UO_1330 (O_1330,N_14357,N_14917);
and UO_1331 (O_1331,N_14882,N_14757);
xnor UO_1332 (O_1332,N_14939,N_14415);
and UO_1333 (O_1333,N_14590,N_14846);
or UO_1334 (O_1334,N_14823,N_14454);
or UO_1335 (O_1335,N_14643,N_14714);
nor UO_1336 (O_1336,N_14553,N_14395);
nor UO_1337 (O_1337,N_14526,N_14788);
xor UO_1338 (O_1338,N_14481,N_14646);
and UO_1339 (O_1339,N_14511,N_14970);
nor UO_1340 (O_1340,N_14720,N_14470);
and UO_1341 (O_1341,N_14925,N_14431);
or UO_1342 (O_1342,N_14849,N_14854);
nor UO_1343 (O_1343,N_14250,N_14304);
nand UO_1344 (O_1344,N_14698,N_14872);
or UO_1345 (O_1345,N_14465,N_14434);
xor UO_1346 (O_1346,N_14898,N_14885);
or UO_1347 (O_1347,N_14328,N_14949);
or UO_1348 (O_1348,N_14788,N_14765);
and UO_1349 (O_1349,N_14569,N_14810);
nand UO_1350 (O_1350,N_14645,N_14382);
nor UO_1351 (O_1351,N_14321,N_14355);
and UO_1352 (O_1352,N_14296,N_14597);
or UO_1353 (O_1353,N_14982,N_14971);
or UO_1354 (O_1354,N_14283,N_14992);
nor UO_1355 (O_1355,N_14306,N_14789);
nor UO_1356 (O_1356,N_14737,N_14413);
nand UO_1357 (O_1357,N_14820,N_14444);
nand UO_1358 (O_1358,N_14597,N_14933);
nand UO_1359 (O_1359,N_14651,N_14619);
and UO_1360 (O_1360,N_14859,N_14748);
and UO_1361 (O_1361,N_14930,N_14831);
or UO_1362 (O_1362,N_14656,N_14334);
nor UO_1363 (O_1363,N_14626,N_14580);
and UO_1364 (O_1364,N_14383,N_14566);
nor UO_1365 (O_1365,N_14440,N_14441);
nor UO_1366 (O_1366,N_14936,N_14928);
nor UO_1367 (O_1367,N_14312,N_14415);
nand UO_1368 (O_1368,N_14478,N_14499);
xnor UO_1369 (O_1369,N_14883,N_14313);
nand UO_1370 (O_1370,N_14325,N_14442);
nand UO_1371 (O_1371,N_14672,N_14730);
nor UO_1372 (O_1372,N_14255,N_14859);
or UO_1373 (O_1373,N_14857,N_14616);
xor UO_1374 (O_1374,N_14969,N_14802);
or UO_1375 (O_1375,N_14691,N_14926);
and UO_1376 (O_1376,N_14574,N_14582);
and UO_1377 (O_1377,N_14772,N_14400);
or UO_1378 (O_1378,N_14991,N_14363);
or UO_1379 (O_1379,N_14421,N_14746);
nand UO_1380 (O_1380,N_14484,N_14675);
and UO_1381 (O_1381,N_14517,N_14468);
xor UO_1382 (O_1382,N_14540,N_14866);
and UO_1383 (O_1383,N_14786,N_14934);
and UO_1384 (O_1384,N_14977,N_14972);
xor UO_1385 (O_1385,N_14266,N_14840);
nor UO_1386 (O_1386,N_14855,N_14274);
and UO_1387 (O_1387,N_14450,N_14302);
nand UO_1388 (O_1388,N_14654,N_14600);
xor UO_1389 (O_1389,N_14889,N_14329);
nor UO_1390 (O_1390,N_14904,N_14914);
nor UO_1391 (O_1391,N_14939,N_14422);
nand UO_1392 (O_1392,N_14884,N_14822);
or UO_1393 (O_1393,N_14423,N_14470);
and UO_1394 (O_1394,N_14397,N_14774);
or UO_1395 (O_1395,N_14566,N_14265);
nand UO_1396 (O_1396,N_14319,N_14745);
or UO_1397 (O_1397,N_14756,N_14590);
nand UO_1398 (O_1398,N_14342,N_14819);
xor UO_1399 (O_1399,N_14984,N_14962);
nand UO_1400 (O_1400,N_14529,N_14385);
xor UO_1401 (O_1401,N_14597,N_14430);
and UO_1402 (O_1402,N_14629,N_14408);
xor UO_1403 (O_1403,N_14524,N_14749);
nor UO_1404 (O_1404,N_14439,N_14537);
or UO_1405 (O_1405,N_14760,N_14731);
or UO_1406 (O_1406,N_14575,N_14549);
xnor UO_1407 (O_1407,N_14277,N_14971);
xor UO_1408 (O_1408,N_14416,N_14985);
or UO_1409 (O_1409,N_14701,N_14843);
nand UO_1410 (O_1410,N_14979,N_14638);
nand UO_1411 (O_1411,N_14715,N_14762);
xor UO_1412 (O_1412,N_14558,N_14648);
or UO_1413 (O_1413,N_14904,N_14667);
xor UO_1414 (O_1414,N_14741,N_14600);
and UO_1415 (O_1415,N_14331,N_14796);
xnor UO_1416 (O_1416,N_14611,N_14900);
xnor UO_1417 (O_1417,N_14830,N_14659);
and UO_1418 (O_1418,N_14674,N_14335);
and UO_1419 (O_1419,N_14794,N_14703);
nand UO_1420 (O_1420,N_14302,N_14443);
xor UO_1421 (O_1421,N_14611,N_14416);
or UO_1422 (O_1422,N_14561,N_14413);
xnor UO_1423 (O_1423,N_14512,N_14864);
or UO_1424 (O_1424,N_14511,N_14814);
nor UO_1425 (O_1425,N_14993,N_14270);
or UO_1426 (O_1426,N_14540,N_14682);
and UO_1427 (O_1427,N_14767,N_14343);
xnor UO_1428 (O_1428,N_14810,N_14769);
or UO_1429 (O_1429,N_14458,N_14462);
nand UO_1430 (O_1430,N_14789,N_14367);
nor UO_1431 (O_1431,N_14799,N_14415);
nor UO_1432 (O_1432,N_14397,N_14285);
nand UO_1433 (O_1433,N_14458,N_14945);
xor UO_1434 (O_1434,N_14759,N_14477);
xor UO_1435 (O_1435,N_14689,N_14709);
or UO_1436 (O_1436,N_14832,N_14607);
or UO_1437 (O_1437,N_14469,N_14935);
xor UO_1438 (O_1438,N_14601,N_14787);
nor UO_1439 (O_1439,N_14971,N_14451);
nand UO_1440 (O_1440,N_14924,N_14803);
nand UO_1441 (O_1441,N_14326,N_14632);
nand UO_1442 (O_1442,N_14353,N_14674);
or UO_1443 (O_1443,N_14917,N_14559);
and UO_1444 (O_1444,N_14942,N_14583);
nor UO_1445 (O_1445,N_14744,N_14780);
or UO_1446 (O_1446,N_14498,N_14697);
xor UO_1447 (O_1447,N_14705,N_14711);
and UO_1448 (O_1448,N_14567,N_14653);
and UO_1449 (O_1449,N_14265,N_14974);
xor UO_1450 (O_1450,N_14708,N_14406);
nand UO_1451 (O_1451,N_14556,N_14644);
nor UO_1452 (O_1452,N_14337,N_14497);
or UO_1453 (O_1453,N_14431,N_14523);
xor UO_1454 (O_1454,N_14632,N_14967);
and UO_1455 (O_1455,N_14721,N_14525);
xnor UO_1456 (O_1456,N_14544,N_14436);
or UO_1457 (O_1457,N_14473,N_14879);
nand UO_1458 (O_1458,N_14658,N_14818);
nor UO_1459 (O_1459,N_14599,N_14782);
and UO_1460 (O_1460,N_14615,N_14668);
or UO_1461 (O_1461,N_14788,N_14394);
nor UO_1462 (O_1462,N_14410,N_14993);
or UO_1463 (O_1463,N_14573,N_14522);
xnor UO_1464 (O_1464,N_14816,N_14577);
nor UO_1465 (O_1465,N_14609,N_14949);
nor UO_1466 (O_1466,N_14565,N_14688);
and UO_1467 (O_1467,N_14466,N_14366);
xor UO_1468 (O_1468,N_14917,N_14299);
and UO_1469 (O_1469,N_14254,N_14887);
and UO_1470 (O_1470,N_14333,N_14361);
nand UO_1471 (O_1471,N_14595,N_14630);
xnor UO_1472 (O_1472,N_14907,N_14995);
and UO_1473 (O_1473,N_14529,N_14947);
or UO_1474 (O_1474,N_14652,N_14495);
and UO_1475 (O_1475,N_14695,N_14459);
nor UO_1476 (O_1476,N_14780,N_14466);
xnor UO_1477 (O_1477,N_14339,N_14429);
nand UO_1478 (O_1478,N_14517,N_14274);
and UO_1479 (O_1479,N_14365,N_14564);
or UO_1480 (O_1480,N_14323,N_14790);
or UO_1481 (O_1481,N_14283,N_14989);
and UO_1482 (O_1482,N_14528,N_14301);
nor UO_1483 (O_1483,N_14998,N_14529);
nand UO_1484 (O_1484,N_14670,N_14674);
xnor UO_1485 (O_1485,N_14456,N_14745);
nor UO_1486 (O_1486,N_14336,N_14794);
or UO_1487 (O_1487,N_14555,N_14784);
nor UO_1488 (O_1488,N_14644,N_14657);
nor UO_1489 (O_1489,N_14965,N_14468);
or UO_1490 (O_1490,N_14943,N_14375);
and UO_1491 (O_1491,N_14842,N_14873);
nor UO_1492 (O_1492,N_14583,N_14413);
nor UO_1493 (O_1493,N_14545,N_14594);
xnor UO_1494 (O_1494,N_14817,N_14384);
and UO_1495 (O_1495,N_14490,N_14786);
xnor UO_1496 (O_1496,N_14423,N_14394);
nor UO_1497 (O_1497,N_14763,N_14741);
nor UO_1498 (O_1498,N_14597,N_14755);
nand UO_1499 (O_1499,N_14737,N_14799);
nand UO_1500 (O_1500,N_14565,N_14379);
xnor UO_1501 (O_1501,N_14264,N_14326);
or UO_1502 (O_1502,N_14895,N_14695);
or UO_1503 (O_1503,N_14883,N_14862);
nand UO_1504 (O_1504,N_14357,N_14973);
nor UO_1505 (O_1505,N_14934,N_14527);
nand UO_1506 (O_1506,N_14411,N_14941);
or UO_1507 (O_1507,N_14807,N_14597);
xor UO_1508 (O_1508,N_14804,N_14293);
nor UO_1509 (O_1509,N_14253,N_14775);
nor UO_1510 (O_1510,N_14630,N_14752);
nor UO_1511 (O_1511,N_14829,N_14993);
and UO_1512 (O_1512,N_14512,N_14914);
xnor UO_1513 (O_1513,N_14425,N_14251);
or UO_1514 (O_1514,N_14672,N_14308);
or UO_1515 (O_1515,N_14633,N_14853);
nor UO_1516 (O_1516,N_14561,N_14541);
nor UO_1517 (O_1517,N_14504,N_14917);
nor UO_1518 (O_1518,N_14544,N_14335);
nor UO_1519 (O_1519,N_14444,N_14632);
xnor UO_1520 (O_1520,N_14873,N_14983);
and UO_1521 (O_1521,N_14341,N_14484);
or UO_1522 (O_1522,N_14716,N_14446);
or UO_1523 (O_1523,N_14806,N_14455);
nor UO_1524 (O_1524,N_14784,N_14946);
and UO_1525 (O_1525,N_14839,N_14335);
xor UO_1526 (O_1526,N_14515,N_14391);
xor UO_1527 (O_1527,N_14789,N_14571);
or UO_1528 (O_1528,N_14358,N_14448);
xnor UO_1529 (O_1529,N_14666,N_14417);
nor UO_1530 (O_1530,N_14892,N_14310);
xnor UO_1531 (O_1531,N_14687,N_14602);
nor UO_1532 (O_1532,N_14884,N_14824);
or UO_1533 (O_1533,N_14985,N_14650);
nand UO_1534 (O_1534,N_14730,N_14268);
and UO_1535 (O_1535,N_14650,N_14321);
nand UO_1536 (O_1536,N_14992,N_14409);
xnor UO_1537 (O_1537,N_14514,N_14648);
or UO_1538 (O_1538,N_14947,N_14995);
and UO_1539 (O_1539,N_14309,N_14990);
or UO_1540 (O_1540,N_14814,N_14295);
or UO_1541 (O_1541,N_14663,N_14772);
nor UO_1542 (O_1542,N_14699,N_14296);
or UO_1543 (O_1543,N_14322,N_14916);
nand UO_1544 (O_1544,N_14662,N_14530);
nor UO_1545 (O_1545,N_14625,N_14306);
nor UO_1546 (O_1546,N_14869,N_14735);
or UO_1547 (O_1547,N_14478,N_14885);
or UO_1548 (O_1548,N_14894,N_14932);
nor UO_1549 (O_1549,N_14945,N_14503);
nor UO_1550 (O_1550,N_14354,N_14353);
or UO_1551 (O_1551,N_14251,N_14411);
nor UO_1552 (O_1552,N_14619,N_14609);
or UO_1553 (O_1553,N_14547,N_14879);
nand UO_1554 (O_1554,N_14846,N_14738);
nor UO_1555 (O_1555,N_14320,N_14940);
or UO_1556 (O_1556,N_14778,N_14511);
xor UO_1557 (O_1557,N_14826,N_14959);
nor UO_1558 (O_1558,N_14803,N_14632);
nand UO_1559 (O_1559,N_14835,N_14391);
and UO_1560 (O_1560,N_14689,N_14877);
xnor UO_1561 (O_1561,N_14343,N_14504);
nor UO_1562 (O_1562,N_14398,N_14534);
or UO_1563 (O_1563,N_14843,N_14324);
and UO_1564 (O_1564,N_14908,N_14533);
nand UO_1565 (O_1565,N_14417,N_14949);
xor UO_1566 (O_1566,N_14436,N_14978);
xnor UO_1567 (O_1567,N_14509,N_14290);
or UO_1568 (O_1568,N_14938,N_14666);
or UO_1569 (O_1569,N_14536,N_14641);
nor UO_1570 (O_1570,N_14417,N_14818);
and UO_1571 (O_1571,N_14359,N_14520);
nand UO_1572 (O_1572,N_14587,N_14926);
xnor UO_1573 (O_1573,N_14435,N_14358);
xnor UO_1574 (O_1574,N_14304,N_14924);
nand UO_1575 (O_1575,N_14569,N_14723);
or UO_1576 (O_1576,N_14583,N_14901);
nand UO_1577 (O_1577,N_14833,N_14916);
nand UO_1578 (O_1578,N_14362,N_14711);
xor UO_1579 (O_1579,N_14912,N_14532);
nor UO_1580 (O_1580,N_14496,N_14544);
or UO_1581 (O_1581,N_14543,N_14704);
nor UO_1582 (O_1582,N_14508,N_14707);
xor UO_1583 (O_1583,N_14678,N_14613);
nor UO_1584 (O_1584,N_14365,N_14945);
or UO_1585 (O_1585,N_14889,N_14956);
nor UO_1586 (O_1586,N_14827,N_14718);
or UO_1587 (O_1587,N_14860,N_14906);
and UO_1588 (O_1588,N_14400,N_14368);
nor UO_1589 (O_1589,N_14495,N_14493);
nor UO_1590 (O_1590,N_14303,N_14717);
or UO_1591 (O_1591,N_14340,N_14627);
xor UO_1592 (O_1592,N_14748,N_14534);
xor UO_1593 (O_1593,N_14845,N_14924);
xnor UO_1594 (O_1594,N_14900,N_14295);
xnor UO_1595 (O_1595,N_14596,N_14402);
nand UO_1596 (O_1596,N_14740,N_14569);
xor UO_1597 (O_1597,N_14763,N_14420);
and UO_1598 (O_1598,N_14680,N_14660);
or UO_1599 (O_1599,N_14599,N_14482);
and UO_1600 (O_1600,N_14900,N_14287);
and UO_1601 (O_1601,N_14843,N_14574);
or UO_1602 (O_1602,N_14729,N_14465);
or UO_1603 (O_1603,N_14531,N_14344);
xnor UO_1604 (O_1604,N_14997,N_14829);
xnor UO_1605 (O_1605,N_14370,N_14705);
nand UO_1606 (O_1606,N_14570,N_14497);
nor UO_1607 (O_1607,N_14641,N_14464);
nand UO_1608 (O_1608,N_14324,N_14646);
or UO_1609 (O_1609,N_14316,N_14784);
nand UO_1610 (O_1610,N_14807,N_14816);
or UO_1611 (O_1611,N_14491,N_14901);
nor UO_1612 (O_1612,N_14953,N_14814);
nor UO_1613 (O_1613,N_14871,N_14663);
or UO_1614 (O_1614,N_14706,N_14509);
or UO_1615 (O_1615,N_14806,N_14420);
and UO_1616 (O_1616,N_14353,N_14428);
nand UO_1617 (O_1617,N_14474,N_14751);
and UO_1618 (O_1618,N_14959,N_14362);
xor UO_1619 (O_1619,N_14867,N_14463);
xor UO_1620 (O_1620,N_14726,N_14254);
and UO_1621 (O_1621,N_14989,N_14322);
nor UO_1622 (O_1622,N_14431,N_14350);
or UO_1623 (O_1623,N_14825,N_14743);
nor UO_1624 (O_1624,N_14819,N_14294);
and UO_1625 (O_1625,N_14948,N_14669);
nand UO_1626 (O_1626,N_14617,N_14797);
xor UO_1627 (O_1627,N_14651,N_14274);
or UO_1628 (O_1628,N_14334,N_14944);
or UO_1629 (O_1629,N_14540,N_14975);
nor UO_1630 (O_1630,N_14542,N_14671);
nand UO_1631 (O_1631,N_14572,N_14604);
and UO_1632 (O_1632,N_14901,N_14594);
or UO_1633 (O_1633,N_14723,N_14885);
and UO_1634 (O_1634,N_14353,N_14736);
nor UO_1635 (O_1635,N_14855,N_14629);
nand UO_1636 (O_1636,N_14415,N_14566);
nand UO_1637 (O_1637,N_14401,N_14615);
xnor UO_1638 (O_1638,N_14527,N_14522);
xnor UO_1639 (O_1639,N_14817,N_14644);
or UO_1640 (O_1640,N_14270,N_14672);
nand UO_1641 (O_1641,N_14892,N_14632);
or UO_1642 (O_1642,N_14750,N_14601);
and UO_1643 (O_1643,N_14705,N_14759);
or UO_1644 (O_1644,N_14409,N_14315);
and UO_1645 (O_1645,N_14367,N_14811);
xnor UO_1646 (O_1646,N_14930,N_14418);
or UO_1647 (O_1647,N_14417,N_14324);
xor UO_1648 (O_1648,N_14393,N_14638);
nor UO_1649 (O_1649,N_14541,N_14891);
or UO_1650 (O_1650,N_14265,N_14592);
xor UO_1651 (O_1651,N_14654,N_14254);
or UO_1652 (O_1652,N_14396,N_14585);
nor UO_1653 (O_1653,N_14675,N_14808);
nor UO_1654 (O_1654,N_14434,N_14537);
or UO_1655 (O_1655,N_14336,N_14524);
xnor UO_1656 (O_1656,N_14848,N_14606);
xor UO_1657 (O_1657,N_14829,N_14897);
or UO_1658 (O_1658,N_14757,N_14621);
or UO_1659 (O_1659,N_14501,N_14443);
and UO_1660 (O_1660,N_14969,N_14955);
xor UO_1661 (O_1661,N_14739,N_14822);
xnor UO_1662 (O_1662,N_14600,N_14449);
nor UO_1663 (O_1663,N_14352,N_14834);
nor UO_1664 (O_1664,N_14758,N_14780);
nand UO_1665 (O_1665,N_14480,N_14424);
xnor UO_1666 (O_1666,N_14496,N_14619);
xnor UO_1667 (O_1667,N_14564,N_14725);
xor UO_1668 (O_1668,N_14737,N_14390);
nand UO_1669 (O_1669,N_14913,N_14472);
or UO_1670 (O_1670,N_14693,N_14927);
nand UO_1671 (O_1671,N_14646,N_14667);
and UO_1672 (O_1672,N_14300,N_14678);
or UO_1673 (O_1673,N_14395,N_14758);
and UO_1674 (O_1674,N_14948,N_14640);
xnor UO_1675 (O_1675,N_14955,N_14451);
nor UO_1676 (O_1676,N_14840,N_14639);
and UO_1677 (O_1677,N_14788,N_14264);
and UO_1678 (O_1678,N_14883,N_14900);
xor UO_1679 (O_1679,N_14370,N_14257);
or UO_1680 (O_1680,N_14992,N_14555);
or UO_1681 (O_1681,N_14921,N_14657);
or UO_1682 (O_1682,N_14336,N_14439);
nor UO_1683 (O_1683,N_14641,N_14995);
xnor UO_1684 (O_1684,N_14481,N_14253);
nand UO_1685 (O_1685,N_14764,N_14974);
or UO_1686 (O_1686,N_14321,N_14886);
xnor UO_1687 (O_1687,N_14795,N_14902);
nor UO_1688 (O_1688,N_14262,N_14577);
or UO_1689 (O_1689,N_14649,N_14335);
nor UO_1690 (O_1690,N_14936,N_14630);
xnor UO_1691 (O_1691,N_14742,N_14839);
nand UO_1692 (O_1692,N_14616,N_14314);
or UO_1693 (O_1693,N_14886,N_14806);
or UO_1694 (O_1694,N_14356,N_14757);
or UO_1695 (O_1695,N_14317,N_14859);
and UO_1696 (O_1696,N_14364,N_14685);
nor UO_1697 (O_1697,N_14366,N_14696);
nor UO_1698 (O_1698,N_14523,N_14721);
xor UO_1699 (O_1699,N_14275,N_14295);
xor UO_1700 (O_1700,N_14473,N_14795);
xor UO_1701 (O_1701,N_14536,N_14684);
or UO_1702 (O_1702,N_14983,N_14556);
nor UO_1703 (O_1703,N_14330,N_14727);
nor UO_1704 (O_1704,N_14651,N_14945);
nand UO_1705 (O_1705,N_14935,N_14836);
nor UO_1706 (O_1706,N_14959,N_14272);
xnor UO_1707 (O_1707,N_14428,N_14878);
and UO_1708 (O_1708,N_14304,N_14682);
xor UO_1709 (O_1709,N_14480,N_14641);
xnor UO_1710 (O_1710,N_14265,N_14666);
nand UO_1711 (O_1711,N_14679,N_14321);
or UO_1712 (O_1712,N_14809,N_14411);
xor UO_1713 (O_1713,N_14861,N_14795);
nand UO_1714 (O_1714,N_14269,N_14470);
and UO_1715 (O_1715,N_14963,N_14569);
nor UO_1716 (O_1716,N_14838,N_14824);
nor UO_1717 (O_1717,N_14491,N_14978);
nand UO_1718 (O_1718,N_14842,N_14650);
and UO_1719 (O_1719,N_14744,N_14959);
and UO_1720 (O_1720,N_14736,N_14635);
nand UO_1721 (O_1721,N_14818,N_14490);
and UO_1722 (O_1722,N_14764,N_14436);
xnor UO_1723 (O_1723,N_14508,N_14294);
nor UO_1724 (O_1724,N_14440,N_14901);
nor UO_1725 (O_1725,N_14797,N_14800);
and UO_1726 (O_1726,N_14453,N_14692);
nand UO_1727 (O_1727,N_14487,N_14444);
xor UO_1728 (O_1728,N_14408,N_14808);
or UO_1729 (O_1729,N_14815,N_14345);
nand UO_1730 (O_1730,N_14551,N_14309);
xor UO_1731 (O_1731,N_14785,N_14665);
nor UO_1732 (O_1732,N_14947,N_14777);
nor UO_1733 (O_1733,N_14418,N_14771);
and UO_1734 (O_1734,N_14959,N_14341);
nor UO_1735 (O_1735,N_14520,N_14583);
nand UO_1736 (O_1736,N_14340,N_14383);
or UO_1737 (O_1737,N_14439,N_14398);
or UO_1738 (O_1738,N_14832,N_14635);
and UO_1739 (O_1739,N_14645,N_14408);
and UO_1740 (O_1740,N_14958,N_14944);
or UO_1741 (O_1741,N_14439,N_14507);
and UO_1742 (O_1742,N_14541,N_14696);
nor UO_1743 (O_1743,N_14370,N_14436);
and UO_1744 (O_1744,N_14714,N_14679);
nand UO_1745 (O_1745,N_14750,N_14676);
and UO_1746 (O_1746,N_14389,N_14378);
xor UO_1747 (O_1747,N_14625,N_14675);
or UO_1748 (O_1748,N_14934,N_14859);
nor UO_1749 (O_1749,N_14437,N_14382);
nor UO_1750 (O_1750,N_14672,N_14857);
nor UO_1751 (O_1751,N_14505,N_14306);
xor UO_1752 (O_1752,N_14993,N_14959);
nand UO_1753 (O_1753,N_14296,N_14942);
nand UO_1754 (O_1754,N_14603,N_14664);
and UO_1755 (O_1755,N_14288,N_14917);
and UO_1756 (O_1756,N_14687,N_14931);
xor UO_1757 (O_1757,N_14416,N_14484);
xnor UO_1758 (O_1758,N_14826,N_14770);
and UO_1759 (O_1759,N_14979,N_14789);
nor UO_1760 (O_1760,N_14433,N_14355);
xnor UO_1761 (O_1761,N_14821,N_14726);
xnor UO_1762 (O_1762,N_14676,N_14760);
xor UO_1763 (O_1763,N_14791,N_14482);
nand UO_1764 (O_1764,N_14687,N_14637);
nor UO_1765 (O_1765,N_14265,N_14320);
nor UO_1766 (O_1766,N_14331,N_14928);
nand UO_1767 (O_1767,N_14644,N_14552);
xnor UO_1768 (O_1768,N_14411,N_14560);
nand UO_1769 (O_1769,N_14634,N_14326);
nand UO_1770 (O_1770,N_14662,N_14663);
nand UO_1771 (O_1771,N_14721,N_14997);
nand UO_1772 (O_1772,N_14370,N_14646);
xor UO_1773 (O_1773,N_14554,N_14751);
and UO_1774 (O_1774,N_14649,N_14730);
nand UO_1775 (O_1775,N_14782,N_14477);
and UO_1776 (O_1776,N_14645,N_14677);
nand UO_1777 (O_1777,N_14518,N_14962);
or UO_1778 (O_1778,N_14971,N_14963);
or UO_1779 (O_1779,N_14425,N_14884);
and UO_1780 (O_1780,N_14679,N_14840);
xor UO_1781 (O_1781,N_14697,N_14746);
nor UO_1782 (O_1782,N_14937,N_14662);
and UO_1783 (O_1783,N_14857,N_14277);
and UO_1784 (O_1784,N_14473,N_14497);
or UO_1785 (O_1785,N_14649,N_14967);
and UO_1786 (O_1786,N_14366,N_14939);
nand UO_1787 (O_1787,N_14824,N_14806);
nor UO_1788 (O_1788,N_14974,N_14448);
nand UO_1789 (O_1789,N_14657,N_14590);
and UO_1790 (O_1790,N_14771,N_14683);
and UO_1791 (O_1791,N_14275,N_14894);
nand UO_1792 (O_1792,N_14969,N_14459);
nor UO_1793 (O_1793,N_14522,N_14922);
nand UO_1794 (O_1794,N_14586,N_14676);
nor UO_1795 (O_1795,N_14354,N_14974);
and UO_1796 (O_1796,N_14775,N_14336);
nand UO_1797 (O_1797,N_14641,N_14585);
nand UO_1798 (O_1798,N_14868,N_14846);
xor UO_1799 (O_1799,N_14933,N_14858);
nand UO_1800 (O_1800,N_14965,N_14873);
nand UO_1801 (O_1801,N_14892,N_14471);
xnor UO_1802 (O_1802,N_14525,N_14809);
and UO_1803 (O_1803,N_14974,N_14499);
nand UO_1804 (O_1804,N_14670,N_14475);
or UO_1805 (O_1805,N_14868,N_14751);
nand UO_1806 (O_1806,N_14765,N_14445);
nor UO_1807 (O_1807,N_14821,N_14316);
and UO_1808 (O_1808,N_14977,N_14283);
and UO_1809 (O_1809,N_14487,N_14266);
nand UO_1810 (O_1810,N_14932,N_14516);
xor UO_1811 (O_1811,N_14900,N_14461);
nor UO_1812 (O_1812,N_14383,N_14741);
nor UO_1813 (O_1813,N_14552,N_14986);
nor UO_1814 (O_1814,N_14327,N_14415);
xnor UO_1815 (O_1815,N_14867,N_14639);
and UO_1816 (O_1816,N_14258,N_14376);
and UO_1817 (O_1817,N_14272,N_14358);
nor UO_1818 (O_1818,N_14970,N_14617);
xor UO_1819 (O_1819,N_14542,N_14270);
nand UO_1820 (O_1820,N_14664,N_14562);
or UO_1821 (O_1821,N_14351,N_14844);
and UO_1822 (O_1822,N_14598,N_14872);
or UO_1823 (O_1823,N_14845,N_14740);
nor UO_1824 (O_1824,N_14797,N_14762);
or UO_1825 (O_1825,N_14709,N_14309);
nor UO_1826 (O_1826,N_14252,N_14636);
or UO_1827 (O_1827,N_14318,N_14268);
or UO_1828 (O_1828,N_14706,N_14590);
xor UO_1829 (O_1829,N_14988,N_14836);
or UO_1830 (O_1830,N_14698,N_14691);
and UO_1831 (O_1831,N_14593,N_14606);
nor UO_1832 (O_1832,N_14728,N_14558);
xor UO_1833 (O_1833,N_14786,N_14919);
nor UO_1834 (O_1834,N_14680,N_14399);
or UO_1835 (O_1835,N_14714,N_14372);
xor UO_1836 (O_1836,N_14787,N_14618);
xor UO_1837 (O_1837,N_14761,N_14929);
or UO_1838 (O_1838,N_14725,N_14280);
nand UO_1839 (O_1839,N_14627,N_14390);
nand UO_1840 (O_1840,N_14572,N_14541);
xor UO_1841 (O_1841,N_14615,N_14829);
and UO_1842 (O_1842,N_14618,N_14423);
and UO_1843 (O_1843,N_14326,N_14736);
and UO_1844 (O_1844,N_14889,N_14825);
nand UO_1845 (O_1845,N_14451,N_14655);
xor UO_1846 (O_1846,N_14709,N_14466);
nor UO_1847 (O_1847,N_14458,N_14388);
and UO_1848 (O_1848,N_14614,N_14282);
nand UO_1849 (O_1849,N_14874,N_14554);
and UO_1850 (O_1850,N_14356,N_14384);
nand UO_1851 (O_1851,N_14937,N_14302);
and UO_1852 (O_1852,N_14263,N_14982);
nor UO_1853 (O_1853,N_14450,N_14938);
nand UO_1854 (O_1854,N_14849,N_14684);
nand UO_1855 (O_1855,N_14833,N_14481);
and UO_1856 (O_1856,N_14949,N_14741);
xor UO_1857 (O_1857,N_14384,N_14574);
nor UO_1858 (O_1858,N_14823,N_14352);
xor UO_1859 (O_1859,N_14612,N_14635);
nand UO_1860 (O_1860,N_14980,N_14701);
nand UO_1861 (O_1861,N_14501,N_14421);
or UO_1862 (O_1862,N_14478,N_14453);
and UO_1863 (O_1863,N_14587,N_14878);
nor UO_1864 (O_1864,N_14763,N_14498);
xnor UO_1865 (O_1865,N_14396,N_14756);
nand UO_1866 (O_1866,N_14696,N_14627);
xnor UO_1867 (O_1867,N_14753,N_14739);
or UO_1868 (O_1868,N_14532,N_14358);
xnor UO_1869 (O_1869,N_14776,N_14895);
and UO_1870 (O_1870,N_14623,N_14875);
nor UO_1871 (O_1871,N_14583,N_14563);
and UO_1872 (O_1872,N_14860,N_14445);
nand UO_1873 (O_1873,N_14923,N_14706);
xnor UO_1874 (O_1874,N_14703,N_14802);
nand UO_1875 (O_1875,N_14861,N_14617);
xor UO_1876 (O_1876,N_14615,N_14820);
nor UO_1877 (O_1877,N_14756,N_14808);
or UO_1878 (O_1878,N_14691,N_14437);
and UO_1879 (O_1879,N_14719,N_14279);
nand UO_1880 (O_1880,N_14360,N_14309);
nand UO_1881 (O_1881,N_14571,N_14715);
nand UO_1882 (O_1882,N_14356,N_14665);
or UO_1883 (O_1883,N_14630,N_14984);
nand UO_1884 (O_1884,N_14812,N_14561);
and UO_1885 (O_1885,N_14596,N_14916);
xor UO_1886 (O_1886,N_14518,N_14529);
nor UO_1887 (O_1887,N_14798,N_14367);
or UO_1888 (O_1888,N_14663,N_14427);
nor UO_1889 (O_1889,N_14498,N_14315);
xnor UO_1890 (O_1890,N_14707,N_14296);
or UO_1891 (O_1891,N_14287,N_14293);
and UO_1892 (O_1892,N_14854,N_14815);
nor UO_1893 (O_1893,N_14584,N_14601);
and UO_1894 (O_1894,N_14372,N_14458);
nor UO_1895 (O_1895,N_14330,N_14864);
nor UO_1896 (O_1896,N_14263,N_14586);
nor UO_1897 (O_1897,N_14689,N_14559);
nand UO_1898 (O_1898,N_14624,N_14855);
xnor UO_1899 (O_1899,N_14491,N_14697);
and UO_1900 (O_1900,N_14497,N_14309);
xor UO_1901 (O_1901,N_14582,N_14889);
nor UO_1902 (O_1902,N_14692,N_14743);
nor UO_1903 (O_1903,N_14922,N_14610);
xnor UO_1904 (O_1904,N_14551,N_14603);
and UO_1905 (O_1905,N_14896,N_14540);
nand UO_1906 (O_1906,N_14805,N_14587);
or UO_1907 (O_1907,N_14736,N_14516);
and UO_1908 (O_1908,N_14432,N_14436);
or UO_1909 (O_1909,N_14259,N_14930);
nor UO_1910 (O_1910,N_14843,N_14707);
nor UO_1911 (O_1911,N_14772,N_14649);
nand UO_1912 (O_1912,N_14812,N_14910);
and UO_1913 (O_1913,N_14596,N_14859);
and UO_1914 (O_1914,N_14350,N_14898);
xor UO_1915 (O_1915,N_14454,N_14939);
xnor UO_1916 (O_1916,N_14724,N_14570);
nand UO_1917 (O_1917,N_14886,N_14614);
and UO_1918 (O_1918,N_14906,N_14928);
nand UO_1919 (O_1919,N_14825,N_14752);
xnor UO_1920 (O_1920,N_14265,N_14431);
xnor UO_1921 (O_1921,N_14458,N_14471);
nand UO_1922 (O_1922,N_14717,N_14912);
and UO_1923 (O_1923,N_14502,N_14635);
nor UO_1924 (O_1924,N_14576,N_14356);
or UO_1925 (O_1925,N_14308,N_14999);
or UO_1926 (O_1926,N_14694,N_14806);
nand UO_1927 (O_1927,N_14679,N_14447);
and UO_1928 (O_1928,N_14803,N_14289);
xor UO_1929 (O_1929,N_14695,N_14290);
nand UO_1930 (O_1930,N_14329,N_14319);
nand UO_1931 (O_1931,N_14662,N_14965);
xor UO_1932 (O_1932,N_14305,N_14488);
xor UO_1933 (O_1933,N_14479,N_14650);
and UO_1934 (O_1934,N_14250,N_14942);
and UO_1935 (O_1935,N_14456,N_14956);
xnor UO_1936 (O_1936,N_14857,N_14503);
or UO_1937 (O_1937,N_14401,N_14585);
nand UO_1938 (O_1938,N_14351,N_14990);
xnor UO_1939 (O_1939,N_14656,N_14946);
nand UO_1940 (O_1940,N_14369,N_14570);
nand UO_1941 (O_1941,N_14843,N_14268);
xnor UO_1942 (O_1942,N_14328,N_14370);
nand UO_1943 (O_1943,N_14305,N_14935);
and UO_1944 (O_1944,N_14533,N_14914);
nor UO_1945 (O_1945,N_14931,N_14363);
xor UO_1946 (O_1946,N_14607,N_14887);
nand UO_1947 (O_1947,N_14723,N_14721);
nor UO_1948 (O_1948,N_14864,N_14322);
or UO_1949 (O_1949,N_14835,N_14477);
or UO_1950 (O_1950,N_14252,N_14400);
or UO_1951 (O_1951,N_14549,N_14261);
nor UO_1952 (O_1952,N_14537,N_14590);
or UO_1953 (O_1953,N_14369,N_14655);
nor UO_1954 (O_1954,N_14299,N_14685);
and UO_1955 (O_1955,N_14769,N_14867);
or UO_1956 (O_1956,N_14641,N_14875);
or UO_1957 (O_1957,N_14944,N_14533);
nand UO_1958 (O_1958,N_14675,N_14434);
nor UO_1959 (O_1959,N_14419,N_14976);
or UO_1960 (O_1960,N_14793,N_14253);
nor UO_1961 (O_1961,N_14415,N_14325);
xor UO_1962 (O_1962,N_14387,N_14469);
nor UO_1963 (O_1963,N_14572,N_14688);
or UO_1964 (O_1964,N_14636,N_14992);
nor UO_1965 (O_1965,N_14253,N_14873);
and UO_1966 (O_1966,N_14314,N_14916);
nor UO_1967 (O_1967,N_14602,N_14995);
nor UO_1968 (O_1968,N_14781,N_14428);
or UO_1969 (O_1969,N_14934,N_14669);
nand UO_1970 (O_1970,N_14397,N_14336);
or UO_1971 (O_1971,N_14911,N_14882);
xor UO_1972 (O_1972,N_14502,N_14887);
and UO_1973 (O_1973,N_14640,N_14368);
nor UO_1974 (O_1974,N_14326,N_14270);
nor UO_1975 (O_1975,N_14637,N_14520);
nand UO_1976 (O_1976,N_14935,N_14591);
nor UO_1977 (O_1977,N_14479,N_14421);
nand UO_1978 (O_1978,N_14383,N_14452);
and UO_1979 (O_1979,N_14759,N_14305);
or UO_1980 (O_1980,N_14556,N_14553);
xnor UO_1981 (O_1981,N_14276,N_14730);
nand UO_1982 (O_1982,N_14950,N_14730);
xnor UO_1983 (O_1983,N_14953,N_14775);
nor UO_1984 (O_1984,N_14322,N_14719);
or UO_1985 (O_1985,N_14492,N_14658);
xnor UO_1986 (O_1986,N_14914,N_14557);
nand UO_1987 (O_1987,N_14846,N_14774);
nand UO_1988 (O_1988,N_14698,N_14899);
xnor UO_1989 (O_1989,N_14426,N_14895);
and UO_1990 (O_1990,N_14802,N_14542);
and UO_1991 (O_1991,N_14284,N_14727);
xor UO_1992 (O_1992,N_14695,N_14421);
and UO_1993 (O_1993,N_14466,N_14359);
nand UO_1994 (O_1994,N_14504,N_14775);
nor UO_1995 (O_1995,N_14278,N_14874);
and UO_1996 (O_1996,N_14472,N_14448);
nand UO_1997 (O_1997,N_14386,N_14536);
xnor UO_1998 (O_1998,N_14835,N_14260);
nand UO_1999 (O_1999,N_14540,N_14445);
endmodule